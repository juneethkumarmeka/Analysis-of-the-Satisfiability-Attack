module basic_5000_50000_5000_10_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
and U0 (N_0,In_4616,In_4281);
and U1 (N_1,In_1519,In_2167);
nand U2 (N_2,In_3738,In_2468);
nand U3 (N_3,In_3180,In_2161);
or U4 (N_4,In_1734,In_57);
nor U5 (N_5,In_3177,In_2143);
or U6 (N_6,In_4465,In_624);
or U7 (N_7,In_2830,In_3515);
nand U8 (N_8,In_658,In_104);
xnor U9 (N_9,In_662,In_1493);
xor U10 (N_10,In_4963,In_1797);
or U11 (N_11,In_967,In_479);
xor U12 (N_12,In_2461,In_577);
or U13 (N_13,In_892,In_3365);
and U14 (N_14,In_1154,In_2436);
nand U15 (N_15,In_4974,In_1149);
and U16 (N_16,In_2101,In_3498);
xor U17 (N_17,In_1349,In_1117);
or U18 (N_18,In_4991,In_4431);
nand U19 (N_19,In_4858,In_3794);
and U20 (N_20,In_3776,In_2431);
and U21 (N_21,In_3345,In_2601);
nor U22 (N_22,In_3882,In_1173);
nor U23 (N_23,In_4178,In_220);
xor U24 (N_24,In_2607,In_3868);
and U25 (N_25,In_847,In_3876);
or U26 (N_26,In_1219,In_1762);
nor U27 (N_27,In_4481,In_4749);
or U28 (N_28,In_1062,In_4631);
or U29 (N_29,In_3624,In_3096);
nand U30 (N_30,In_1524,In_619);
nor U31 (N_31,In_4012,In_3148);
or U32 (N_32,In_2994,In_4862);
xnor U33 (N_33,In_4493,In_1268);
or U34 (N_34,In_79,In_1472);
xnor U35 (N_35,In_3470,In_2875);
or U36 (N_36,In_2706,In_3815);
or U37 (N_37,In_4747,In_1764);
xor U38 (N_38,In_4022,In_2);
or U39 (N_39,In_3424,In_990);
xnor U40 (N_40,In_4180,In_1082);
or U41 (N_41,In_396,In_958);
xnor U42 (N_42,In_935,In_2139);
or U43 (N_43,In_2929,In_2338);
or U44 (N_44,In_1435,In_4921);
or U45 (N_45,In_4225,In_1412);
nor U46 (N_46,In_3136,In_1107);
xnor U47 (N_47,In_4418,In_947);
or U48 (N_48,In_767,In_3203);
xnor U49 (N_49,In_3128,In_3328);
nand U50 (N_50,In_1186,In_2464);
or U51 (N_51,In_1758,In_2515);
nor U52 (N_52,In_2681,In_38);
or U53 (N_53,In_3621,In_1692);
and U54 (N_54,In_39,In_3113);
nand U55 (N_55,In_2459,In_1247);
nor U56 (N_56,In_4855,In_4803);
xnor U57 (N_57,In_2068,In_4321);
xnor U58 (N_58,In_1943,In_572);
xnor U59 (N_59,In_2734,In_696);
nand U60 (N_60,In_4655,In_2888);
nand U61 (N_61,In_4039,In_2320);
and U62 (N_62,In_91,In_4625);
and U63 (N_63,In_1682,In_3332);
nand U64 (N_64,In_4877,In_2259);
or U65 (N_65,In_2597,In_1482);
and U66 (N_66,In_668,In_3909);
and U67 (N_67,In_4863,In_1452);
nand U68 (N_68,In_2121,In_4918);
and U69 (N_69,In_1877,In_3510);
xor U70 (N_70,In_3719,In_3667);
nand U71 (N_71,In_4259,In_4739);
nand U72 (N_72,In_394,In_4816);
and U73 (N_73,In_639,In_2268);
xor U74 (N_74,In_1122,In_1458);
and U75 (N_75,In_46,In_747);
or U76 (N_76,In_1688,In_4154);
nor U77 (N_77,In_1230,In_2294);
xor U78 (N_78,In_1779,In_4675);
or U79 (N_79,In_2744,In_1495);
nor U80 (N_80,In_4235,In_2614);
nand U81 (N_81,In_675,In_1893);
or U82 (N_82,In_4490,In_3171);
and U83 (N_83,In_1376,In_3573);
nand U84 (N_84,In_3795,In_326);
and U85 (N_85,In_4685,In_571);
nand U86 (N_86,In_2424,In_3756);
and U87 (N_87,In_3712,In_3578);
nand U88 (N_88,In_4046,In_1578);
and U89 (N_89,In_3778,In_646);
or U90 (N_90,In_4577,In_2066);
and U91 (N_91,In_4289,In_2708);
nand U92 (N_92,In_1052,In_4884);
and U93 (N_93,In_2947,In_4860);
nor U94 (N_94,In_918,In_1539);
nor U95 (N_95,In_3351,In_1799);
xnor U96 (N_96,In_2185,In_4204);
xnor U97 (N_97,In_2403,In_2998);
or U98 (N_98,In_921,In_1743);
nor U99 (N_99,In_1293,In_3052);
nand U100 (N_100,In_2979,In_2444);
nor U101 (N_101,In_4854,In_3438);
nor U102 (N_102,In_3494,In_4732);
xnor U103 (N_103,In_4116,In_1379);
and U104 (N_104,In_1403,In_1803);
nor U105 (N_105,In_3408,In_4314);
nor U106 (N_106,In_1141,In_2524);
and U107 (N_107,In_3919,In_4946);
nand U108 (N_108,In_2132,In_727);
nand U109 (N_109,In_4993,In_93);
and U110 (N_110,In_1862,In_1777);
nor U111 (N_111,In_36,In_3064);
and U112 (N_112,In_928,In_1419);
or U113 (N_113,In_965,In_688);
nor U114 (N_114,In_1928,In_3822);
nor U115 (N_115,In_1248,In_4920);
nand U116 (N_116,In_3459,In_355);
and U117 (N_117,In_2800,In_2663);
xor U118 (N_118,In_2946,In_4642);
or U119 (N_119,In_2102,In_4724);
xor U120 (N_120,In_3143,In_2650);
and U121 (N_121,In_995,In_2784);
nor U122 (N_122,In_4410,In_1182);
xor U123 (N_123,In_2545,In_4442);
and U124 (N_124,In_4443,In_1297);
nand U125 (N_125,In_1469,In_3561);
or U126 (N_126,In_638,In_72);
and U127 (N_127,In_2322,In_217);
or U128 (N_128,In_2127,In_3629);
nand U129 (N_129,In_4379,In_3486);
nor U130 (N_130,In_1146,In_4069);
or U131 (N_131,In_1430,In_1597);
or U132 (N_132,In_3854,In_3541);
nor U133 (N_133,In_4663,In_3651);
nor U134 (N_134,In_3090,In_1063);
nor U135 (N_135,In_327,In_4602);
or U136 (N_136,In_3635,In_4793);
or U137 (N_137,In_2756,In_2973);
xnor U138 (N_138,In_2125,In_2120);
or U139 (N_139,In_3964,In_2260);
nor U140 (N_140,In_4590,In_286);
nand U141 (N_141,In_3114,In_524);
and U142 (N_142,In_835,In_922);
nand U143 (N_143,In_4233,In_1974);
xnor U144 (N_144,In_2060,In_3791);
nor U145 (N_145,In_1548,In_1038);
and U146 (N_146,In_4859,In_2200);
nand U147 (N_147,In_1627,In_779);
nand U148 (N_148,In_1262,In_4640);
and U149 (N_149,In_3285,In_4010);
nor U150 (N_150,In_651,In_765);
xor U151 (N_151,In_4215,In_4436);
nand U152 (N_152,In_301,In_2608);
xnor U153 (N_153,In_3511,In_3352);
or U154 (N_154,In_1410,In_3263);
xor U155 (N_155,In_2350,In_4997);
nor U156 (N_156,In_2171,In_4825);
xor U157 (N_157,In_3230,In_756);
or U158 (N_158,In_989,In_2703);
nand U159 (N_159,In_609,In_813);
xnor U160 (N_160,In_3767,In_1355);
or U161 (N_161,In_2212,In_889);
nand U162 (N_162,In_595,In_4444);
xnor U163 (N_163,In_2218,In_3249);
xnor U164 (N_164,In_3082,In_2346);
nand U165 (N_165,In_3048,In_4341);
nor U166 (N_166,In_810,In_2225);
or U167 (N_167,In_1610,In_1947);
nand U168 (N_168,In_1282,In_2899);
and U169 (N_169,In_3679,In_4193);
or U170 (N_170,In_1654,In_2027);
nand U171 (N_171,In_478,In_2670);
and U172 (N_172,In_1973,In_1044);
and U173 (N_173,In_4274,In_1331);
nor U174 (N_174,In_4250,In_1089);
nand U175 (N_175,In_681,In_2540);
nand U176 (N_176,In_1833,In_1908);
xor U177 (N_177,In_1914,In_2053);
nand U178 (N_178,In_339,In_1480);
or U179 (N_179,In_4307,In_1424);
nand U180 (N_180,In_4750,In_1522);
or U181 (N_181,In_8,In_4578);
nand U182 (N_182,In_415,In_4714);
and U183 (N_183,In_2882,In_4683);
nor U184 (N_184,In_2932,In_1967);
or U185 (N_185,In_771,In_3466);
and U186 (N_186,In_3562,In_443);
nand U187 (N_187,In_1948,In_3922);
nor U188 (N_188,In_130,In_3808);
xnor U189 (N_189,In_1924,In_4780);
xnor U190 (N_190,In_485,In_1401);
xor U191 (N_191,In_1949,In_4807);
or U192 (N_192,In_2592,In_1715);
nand U193 (N_193,In_4645,In_1673);
nor U194 (N_194,In_1638,In_2668);
xnor U195 (N_195,In_1371,In_4832);
or U196 (N_196,In_246,In_2737);
nand U197 (N_197,In_3613,In_566);
nand U198 (N_198,In_1712,In_976);
or U199 (N_199,In_4820,In_3897);
nand U200 (N_200,In_3540,In_2581);
nor U201 (N_201,In_393,In_1783);
and U202 (N_202,In_1237,In_527);
xor U203 (N_203,In_4025,In_3967);
nand U204 (N_204,In_3106,In_3769);
nor U205 (N_205,In_1164,In_2775);
nor U206 (N_206,In_1716,In_4870);
and U207 (N_207,In_334,In_290);
or U208 (N_208,In_4659,In_161);
or U209 (N_209,In_1813,In_4298);
nand U210 (N_210,In_3229,In_4387);
xor U211 (N_211,In_731,In_2666);
nor U212 (N_212,In_2187,In_4679);
and U213 (N_213,In_773,In_3824);
or U214 (N_214,In_1547,In_2988);
or U215 (N_215,In_784,In_3902);
and U216 (N_216,In_3780,In_742);
nor U217 (N_217,In_3444,In_4762);
xor U218 (N_218,In_4909,In_1115);
nand U219 (N_219,In_4463,In_4575);
xnor U220 (N_220,In_1285,In_1781);
or U221 (N_221,In_3432,In_1582);
nor U222 (N_222,In_1301,In_4893);
nor U223 (N_223,In_4474,In_1213);
and U224 (N_224,In_185,In_4834);
nor U225 (N_225,In_1546,In_4285);
nor U226 (N_226,In_3088,In_833);
nor U227 (N_227,In_37,In_4030);
nor U228 (N_228,In_1347,In_1123);
xnor U229 (N_229,In_3924,In_2921);
nand U230 (N_230,In_1827,In_1459);
nor U231 (N_231,In_4149,In_2859);
xor U232 (N_232,In_3724,In_4435);
and U233 (N_233,In_4252,In_2164);
nor U234 (N_234,In_4302,In_3007);
or U235 (N_235,In_1793,In_4172);
xnor U236 (N_236,In_776,In_2684);
xnor U237 (N_237,In_4579,In_1380);
and U238 (N_238,In_151,In_2748);
nand U239 (N_239,In_1859,In_2504);
nand U240 (N_240,In_23,In_399);
xnor U241 (N_241,In_1405,In_3147);
nand U242 (N_242,In_2099,In_1809);
nand U243 (N_243,In_3931,In_4766);
or U244 (N_244,In_2502,In_1315);
nand U245 (N_245,In_1385,In_3454);
nor U246 (N_246,In_163,In_3832);
nor U247 (N_247,In_1589,In_2385);
xnor U248 (N_248,In_514,In_1303);
and U249 (N_249,In_1216,In_3025);
nand U250 (N_250,In_2747,In_1151);
nor U251 (N_251,In_1953,In_3517);
nor U252 (N_252,In_1966,In_2626);
or U253 (N_253,In_991,In_2525);
xnor U254 (N_254,In_3903,In_4557);
nand U255 (N_255,In_2713,In_2443);
nand U256 (N_256,In_3698,In_2889);
xor U257 (N_257,In_735,In_1921);
nor U258 (N_258,In_542,In_769);
and U259 (N_259,In_3349,In_3845);
nor U260 (N_260,In_3550,In_3284);
nand U261 (N_261,In_4571,In_1572);
nand U262 (N_262,In_245,In_1475);
xor U263 (N_263,In_1614,In_1003);
or U264 (N_264,In_4282,In_3786);
nand U265 (N_265,In_2850,In_4197);
or U266 (N_266,In_3032,In_4491);
nor U267 (N_267,In_1969,In_895);
or U268 (N_268,In_2588,In_3890);
xor U269 (N_269,In_3084,In_2300);
nand U270 (N_270,In_1902,In_3783);
nor U271 (N_271,In_715,In_2825);
xnor U272 (N_272,In_2559,In_4420);
xnor U273 (N_273,In_67,In_2216);
nor U274 (N_274,In_1681,In_351);
and U275 (N_275,In_3848,In_437);
or U276 (N_276,In_4191,In_1917);
nor U277 (N_277,In_348,In_2495);
xor U278 (N_278,In_1940,In_2590);
or U279 (N_279,In_4156,In_1552);
nor U280 (N_280,In_1897,In_3563);
nor U281 (N_281,In_1497,In_4488);
and U282 (N_282,In_4139,In_3857);
or U283 (N_283,In_3010,In_1790);
and U284 (N_284,In_4222,In_2827);
or U285 (N_285,In_1810,In_2657);
xor U286 (N_286,In_3525,In_3900);
nor U287 (N_287,In_1901,In_4853);
nand U288 (N_288,In_2571,In_678);
and U289 (N_289,In_2206,In_796);
xnor U290 (N_290,In_2849,In_3601);
and U291 (N_291,In_753,In_4323);
nor U292 (N_292,In_2142,In_2846);
nor U293 (N_293,In_1135,In_2586);
and U294 (N_294,In_350,In_4665);
or U295 (N_295,In_4413,In_4547);
or U296 (N_296,In_1359,In_4623);
nor U297 (N_297,In_4620,In_208);
nor U298 (N_298,In_3279,In_4704);
or U299 (N_299,In_3233,In_3571);
nand U300 (N_300,In_2238,In_3990);
nor U301 (N_301,In_3535,In_317);
nand U302 (N_302,In_1880,In_710);
nand U303 (N_303,In_4981,In_4260);
nand U304 (N_304,In_3181,In_4707);
and U305 (N_305,In_1343,In_2520);
and U306 (N_306,In_4868,In_2742);
nor U307 (N_307,In_3210,In_353);
nand U308 (N_308,In_3384,In_4389);
and U309 (N_309,In_1163,In_3929);
nor U310 (N_310,In_674,In_2088);
and U311 (N_311,In_48,In_235);
and U312 (N_312,In_1402,In_2126);
xor U313 (N_313,In_4367,In_2430);
or U314 (N_314,In_3893,In_2730);
xnor U315 (N_315,In_1570,In_2304);
nor U316 (N_316,In_3245,In_938);
or U317 (N_317,In_4541,In_4753);
and U318 (N_318,In_559,In_4350);
nand U319 (N_319,In_243,In_2579);
and U320 (N_320,In_728,In_3140);
nor U321 (N_321,In_1772,In_2278);
and U322 (N_322,In_3252,In_4654);
xnor U323 (N_323,In_581,In_1253);
and U324 (N_324,In_3669,In_3717);
xor U325 (N_325,In_386,In_4908);
nand U326 (N_326,In_4839,In_585);
nor U327 (N_327,In_3544,In_1363);
nor U328 (N_328,In_2337,In_3178);
xor U329 (N_329,In_3984,In_3539);
and U330 (N_330,In_794,In_439);
and U331 (N_331,In_1291,In_3907);
nor U332 (N_332,In_2675,In_4374);
and U333 (N_333,In_3527,In_1700);
nand U334 (N_334,In_692,In_2378);
nand U335 (N_335,In_377,In_318);
xor U336 (N_336,In_171,In_2492);
and U337 (N_337,In_2149,In_540);
and U338 (N_338,In_2572,In_4040);
or U339 (N_339,In_2632,In_512);
xor U340 (N_340,In_2890,In_3130);
nor U341 (N_341,In_4245,In_2363);
or U342 (N_342,In_2642,In_4689);
nand U343 (N_343,In_3366,In_1321);
or U344 (N_344,In_461,In_466);
nor U345 (N_345,In_1795,In_2479);
nor U346 (N_346,In_590,In_374);
xor U347 (N_347,In_854,In_2544);
nand U348 (N_348,In_240,In_4630);
nor U349 (N_349,In_1330,In_0);
xnor U350 (N_350,In_1312,In_2437);
and U351 (N_351,In_3315,In_3939);
and U352 (N_352,In_809,In_1982);
xor U353 (N_353,In_3702,In_4668);
nand U354 (N_354,In_3191,In_2037);
or U355 (N_355,In_4947,In_2871);
or U356 (N_356,In_2458,In_844);
nand U357 (N_357,In_4822,In_2814);
or U358 (N_358,In_1538,In_225);
nand U359 (N_359,In_4660,In_4105);
nor U360 (N_360,In_1605,In_495);
or U361 (N_361,In_1602,In_3456);
xnor U362 (N_362,In_2123,In_1626);
or U363 (N_363,In_4896,In_1776);
nand U364 (N_364,In_837,In_1370);
or U365 (N_365,In_2878,In_3912);
nor U366 (N_366,In_849,In_2274);
nor U367 (N_367,In_1250,In_1300);
xnor U368 (N_368,In_2348,In_1218);
nor U369 (N_369,In_4574,In_234);
nand U370 (N_370,In_1968,In_1275);
and U371 (N_371,In_3138,In_1986);
and U372 (N_372,In_3666,In_4228);
xor U373 (N_373,In_222,In_2381);
nand U374 (N_374,In_2094,In_4459);
xnor U375 (N_375,In_1110,In_2330);
or U376 (N_376,In_565,In_421);
nor U377 (N_377,In_4009,In_4375);
xor U378 (N_378,In_997,In_346);
or U379 (N_379,In_3219,In_550);
xor U380 (N_380,In_1494,In_2506);
xnor U381 (N_381,In_3436,In_1634);
nor U382 (N_382,In_3676,In_3913);
or U383 (N_383,In_2289,In_683);
or U384 (N_384,In_4552,In_2508);
nand U385 (N_385,In_2992,In_4455);
or U386 (N_386,In_1478,In_1389);
xor U387 (N_387,In_2858,In_4475);
or U388 (N_388,In_763,In_4824);
xnor U389 (N_389,In_2232,In_4721);
xnor U390 (N_390,In_1018,In_4889);
xnor U391 (N_391,In_1143,In_4477);
nand U392 (N_392,In_3251,In_2604);
nor U393 (N_393,In_4220,In_3194);
nand U394 (N_394,In_179,In_3940);
or U395 (N_395,In_836,In_3699);
xnor U396 (N_396,In_3974,In_1575);
nor U397 (N_397,In_3448,In_2145);
and U398 (N_398,In_4351,In_3329);
nand U399 (N_399,In_1514,In_1223);
and U400 (N_400,In_2439,In_4429);
and U401 (N_401,In_3516,In_3162);
nor U402 (N_402,In_3412,In_3086);
nand U403 (N_403,In_2595,In_2175);
nand U404 (N_404,In_2774,In_498);
or U405 (N_405,In_4174,In_3326);
xnor U406 (N_406,In_4984,In_4754);
nand U407 (N_407,In_4800,In_966);
xor U408 (N_408,In_3265,In_3642);
and U409 (N_409,In_108,In_2453);
or U410 (N_410,In_2549,In_2168);
or U411 (N_411,In_2533,In_3434);
and U412 (N_412,In_1442,In_939);
or U413 (N_413,In_2897,In_4564);
and U414 (N_414,In_4534,In_1709);
nand U415 (N_415,In_4062,In_1856);
nand U416 (N_416,In_4155,In_10);
xor U417 (N_417,In_1368,In_409);
and U418 (N_418,In_1705,In_4271);
or U419 (N_419,In_424,In_418);
xor U420 (N_420,In_4267,In_3672);
nand U421 (N_421,In_73,In_1574);
nand U422 (N_422,In_3886,In_4597);
nand U423 (N_423,In_2205,In_1946);
or U424 (N_424,In_912,In_3925);
and U425 (N_425,In_2686,In_2964);
nand U426 (N_426,In_3611,In_459);
and U427 (N_427,In_119,In_3906);
nand U428 (N_428,In_1188,In_4037);
or U429 (N_429,In_1227,In_4954);
nand U430 (N_430,In_2327,In_1890);
and U431 (N_431,In_4347,In_2059);
or U432 (N_432,In_4052,In_2812);
nor U433 (N_433,In_1782,In_3376);
or U434 (N_434,In_1453,In_262);
or U435 (N_435,In_3999,In_631);
or U436 (N_436,In_2408,In_3121);
xnor U437 (N_437,In_4656,In_3830);
xor U438 (N_438,In_2917,In_2315);
or U439 (N_439,In_2521,In_1704);
or U440 (N_440,In_4923,In_4546);
xnor U441 (N_441,In_2012,In_2065);
and U442 (N_442,In_3866,In_3819);
or U443 (N_443,In_3789,In_2823);
and U444 (N_444,In_507,In_63);
nor U445 (N_445,In_3149,In_2317);
nand U446 (N_446,In_3861,In_2951);
nand U447 (N_447,In_821,In_2165);
and U448 (N_448,In_3443,In_3644);
nor U449 (N_449,In_3125,In_1719);
nand U450 (N_450,In_1422,In_3617);
nor U451 (N_451,In_21,In_337);
xnor U452 (N_452,In_3641,In_3221);
or U453 (N_453,In_4523,In_896);
nand U454 (N_454,In_3051,In_4967);
xnor U455 (N_455,In_3093,In_3986);
nor U456 (N_456,In_3942,In_1831);
or U457 (N_457,In_3850,In_4018);
nand U458 (N_458,In_2990,In_2537);
nand U459 (N_459,In_948,In_3610);
nand U460 (N_460,In_2518,In_3943);
nand U461 (N_461,In_4061,In_2199);
nand U462 (N_462,In_3319,In_4091);
xnor U463 (N_463,In_2332,In_3640);
and U464 (N_464,In_1148,In_3379);
and U465 (N_465,In_2954,In_453);
xnor U466 (N_466,In_4035,In_2213);
nand U467 (N_467,In_1222,In_2934);
or U468 (N_468,In_3422,In_3634);
and U469 (N_469,In_4764,In_4497);
or U470 (N_470,In_2630,In_4412);
xnor U471 (N_471,In_711,In_2301);
and U472 (N_472,In_2637,In_4473);
and U473 (N_473,In_1283,In_1544);
and U474 (N_474,In_3735,In_2024);
nor U475 (N_475,In_2894,In_2722);
xnor U476 (N_476,In_1729,In_3318);
nand U477 (N_477,In_2781,In_1642);
or U478 (N_478,In_4958,In_297);
and U479 (N_479,In_4338,In_2420);
xor U480 (N_480,In_2486,In_3190);
or U481 (N_481,In_4084,In_1333);
nor U482 (N_482,In_1249,In_70);
nand U483 (N_483,In_2901,In_919);
nor U484 (N_484,In_2564,In_2451);
and U485 (N_485,In_4142,In_1741);
nand U486 (N_486,In_471,In_1980);
nand U487 (N_487,In_2032,In_2879);
or U488 (N_488,In_253,In_2982);
xor U489 (N_489,In_1996,In_69);
xor U490 (N_490,In_218,In_32);
nand U491 (N_491,In_3117,In_2654);
or U492 (N_492,In_2252,In_3399);
xor U493 (N_493,In_2217,In_444);
or U494 (N_494,In_3739,In_920);
and U495 (N_495,In_1278,In_2360);
nand U496 (N_496,In_3325,In_3585);
and U497 (N_497,In_2705,In_3748);
nor U498 (N_498,In_3732,In_1077);
nor U499 (N_499,In_1925,In_2215);
nor U500 (N_500,In_4880,In_3846);
nand U501 (N_501,In_2151,In_4945);
or U502 (N_502,In_400,In_1096);
nor U503 (N_503,In_4275,In_2691);
nand U504 (N_504,In_258,In_3445);
nor U505 (N_505,In_1245,In_85);
and U506 (N_506,In_3948,In_3950);
nor U507 (N_507,In_4499,In_3395);
xnor U508 (N_508,In_1543,In_3975);
nor U509 (N_509,In_3529,In_1745);
or U510 (N_510,In_3281,In_118);
or U511 (N_511,In_3323,In_4633);
xor U512 (N_512,In_3295,In_3650);
or U513 (N_513,In_1395,In_3195);
nor U514 (N_514,In_1034,In_140);
and U515 (N_515,In_3526,In_3873);
and U516 (N_516,In_4583,In_4306);
nor U517 (N_517,In_628,In_4171);
xnor U518 (N_518,In_943,In_1920);
and U519 (N_519,In_2098,In_955);
or U520 (N_520,In_1104,In_135);
xor U521 (N_521,In_1130,In_4518);
and U522 (N_522,In_3881,In_3170);
xor U523 (N_523,In_2071,In_2644);
xnor U524 (N_524,In_875,In_3107);
nand U525 (N_525,In_3556,In_4266);
and U526 (N_526,In_4134,In_2778);
xnor U527 (N_527,In_4417,In_3409);
nor U528 (N_528,In_3670,In_3680);
nor U529 (N_529,In_4622,In_3904);
or U530 (N_530,In_3752,In_4598);
nand U531 (N_531,In_2843,In_4636);
nand U532 (N_532,In_4368,In_2625);
and U533 (N_533,In_4295,In_4118);
nand U534 (N_534,In_113,In_1759);
nor U535 (N_535,In_3992,In_3167);
and U536 (N_536,In_3065,In_4555);
xor U537 (N_537,In_3473,In_2908);
or U538 (N_538,In_2399,In_926);
and U539 (N_539,In_3760,In_4028);
nor U540 (N_540,In_3116,In_1952);
and U541 (N_541,In_2247,In_4089);
and U542 (N_542,In_852,In_420);
and U543 (N_543,In_1,In_3728);
nor U544 (N_544,In_3759,In_3471);
nor U545 (N_545,In_548,In_4408);
nand U546 (N_546,In_1760,In_2272);
xnor U547 (N_547,In_2280,In_3154);
xnor U548 (N_548,In_1336,In_4354);
nor U549 (N_549,In_923,In_2860);
and U550 (N_550,In_4876,In_626);
nand U551 (N_551,In_517,In_899);
and U552 (N_552,In_2826,In_4183);
or U553 (N_553,In_506,In_376);
nand U554 (N_554,In_788,In_3447);
nand U555 (N_555,In_4309,In_4544);
nor U556 (N_556,In_3311,In_4986);
and U557 (N_557,In_3347,In_1464);
nand U558 (N_558,In_3962,In_4470);
xor U559 (N_559,In_2928,In_1069);
nand U560 (N_560,In_3996,In_1780);
nor U561 (N_561,In_614,In_1257);
or U562 (N_562,In_4162,In_2531);
nand U563 (N_563,In_4044,In_1733);
and U564 (N_564,In_4680,In_2963);
and U565 (N_565,In_2207,In_4643);
nand U566 (N_566,In_3380,In_4828);
and U567 (N_567,In_4242,In_1023);
or U568 (N_568,In_263,In_3308);
or U569 (N_569,In_4738,In_2835);
and U570 (N_570,In_2128,In_30);
nand U571 (N_571,In_3733,In_642);
and U572 (N_572,In_473,In_1346);
and U573 (N_573,In_1721,In_978);
nor U574 (N_574,In_1592,In_3689);
nor U575 (N_575,In_2851,In_3031);
nand U576 (N_576,In_1449,In_2903);
or U577 (N_577,In_1997,In_3983);
nor U578 (N_578,In_3009,In_504);
nor U579 (N_579,In_1279,In_797);
xnor U580 (N_580,In_557,In_3407);
and U581 (N_581,In_2924,In_4254);
and U582 (N_582,In_31,In_764);
nor U583 (N_583,In_4894,In_4219);
nand U584 (N_584,In_4005,In_1364);
nand U585 (N_585,In_1964,In_3937);
nand U586 (N_586,In_3020,In_1033);
nand U587 (N_587,In_413,In_3623);
xnor U588 (N_588,In_1977,In_3665);
or U589 (N_589,In_795,In_3901);
nand U590 (N_590,In_4533,In_1039);
or U591 (N_591,In_867,In_2499);
nor U592 (N_592,In_4530,In_4416);
nor U593 (N_593,In_723,In_4769);
and U594 (N_594,In_2428,In_4352);
nand U595 (N_595,In_1569,In_3357);
xor U596 (N_596,In_1837,In_4294);
xnor U597 (N_597,In_2589,In_4122);
nor U598 (N_598,In_2347,In_607);
xor U599 (N_599,In_3860,In_164);
or U600 (N_600,In_945,In_4189);
nand U601 (N_601,In_4126,In_2249);
and U602 (N_602,In_4987,In_685);
or U603 (N_603,In_3889,In_1471);
and U604 (N_604,In_4553,In_3716);
xor U605 (N_605,In_3997,In_2214);
nor U606 (N_606,In_307,In_724);
nand U607 (N_607,In_914,In_215);
xor U608 (N_608,In_1652,In_4449);
nor U609 (N_609,In_474,In_308);
nor U610 (N_610,In_1177,In_14);
nand U611 (N_611,In_1407,In_3145);
or U612 (N_612,In_2080,In_824);
xor U613 (N_613,In_2967,In_1307);
nor U614 (N_614,In_62,In_1428);
nor U615 (N_615,In_4403,In_1298);
or U616 (N_616,In_1933,In_3417);
and U617 (N_617,In_2299,In_1987);
nand U618 (N_618,In_3455,In_1391);
xnor U619 (N_619,In_2466,In_1600);
nor U620 (N_620,In_1515,In_2824);
nor U621 (N_621,In_3478,In_4453);
xor U622 (N_622,In_4340,In_4814);
nor U623 (N_623,In_1097,In_3095);
xnor U624 (N_624,In_1630,In_3371);
or U625 (N_625,In_1255,In_3797);
or U626 (N_626,In_304,In_500);
or U627 (N_627,In_3092,In_4344);
nor U628 (N_628,In_2271,In_4264);
and U629 (N_629,In_4634,In_383);
or U630 (N_630,In_961,In_3122);
nor U631 (N_631,In_391,In_4796);
nor U632 (N_632,In_2834,In_2489);
nor U633 (N_633,In_1171,In_1903);
nand U634 (N_634,In_4396,In_4919);
nand U635 (N_635,In_4904,In_3420);
or U636 (N_636,In_4941,In_4141);
nand U637 (N_637,In_3021,In_1983);
nor U638 (N_638,In_3260,In_4014);
xnor U639 (N_639,In_1773,In_4372);
or U640 (N_640,In_275,In_1120);
nand U641 (N_641,In_4725,In_547);
or U642 (N_642,In_1679,In_673);
nand U643 (N_643,In_4482,In_4194);
or U644 (N_644,In_2288,In_1697);
nor U645 (N_645,In_289,In_4406);
xnor U646 (N_646,In_3362,In_2556);
nand U647 (N_647,In_3419,In_906);
or U648 (N_648,In_2432,In_120);
nor U649 (N_649,In_1621,In_3450);
nand U650 (N_650,In_4959,In_1577);
or U651 (N_651,In_980,In_4329);
or U652 (N_652,In_3500,In_1489);
and U653 (N_653,In_4070,In_4838);
xnor U654 (N_654,In_616,In_925);
and U655 (N_655,In_184,In_4844);
xnor U656 (N_656,In_3859,In_1579);
or U657 (N_657,In_3076,In_1789);
and U658 (N_658,In_4311,In_3898);
and U659 (N_659,In_1246,In_1613);
or U660 (N_660,In_4569,In_755);
xor U661 (N_661,In_1317,In_1839);
and U662 (N_662,In_754,In_4976);
xor U663 (N_663,In_830,In_3189);
nor U664 (N_664,In_1649,In_1103);
xnor U665 (N_665,In_3877,In_4939);
xnor U666 (N_666,In_2961,In_4962);
and U667 (N_667,In_2405,In_3183);
or U668 (N_668,In_78,In_1690);
or U669 (N_669,In_2805,In_47);
or U670 (N_670,In_1868,In_1179);
or U671 (N_671,In_3003,In_1046);
or U672 (N_672,In_1785,In_3870);
and U673 (N_673,In_1528,In_2627);
and U674 (N_674,In_4415,In_182);
xor U675 (N_675,In_1226,In_3820);
or U676 (N_676,In_3928,In_3591);
or U677 (N_677,In_789,In_4639);
xor U678 (N_678,In_3440,In_3439);
xor U679 (N_679,In_4223,In_4911);
nor U680 (N_680,In_1236,In_843);
nor U681 (N_681,In_313,In_1944);
nand U682 (N_682,In_2269,In_4072);
xnor U683 (N_683,In_2390,In_1158);
or U684 (N_684,In_3368,In_2078);
nor U685 (N_685,In_2821,In_2538);
nand U686 (N_686,In_1792,In_2612);
and U687 (N_687,In_3994,In_2364);
nand U688 (N_688,In_1923,In_2202);
and U689 (N_689,In_2661,In_2010);
and U690 (N_690,In_1205,In_630);
nand U691 (N_691,In_2984,In_2029);
xnor U692 (N_692,In_591,In_1121);
nand U693 (N_693,In_4407,In_1109);
nor U694 (N_694,In_277,In_917);
nor U695 (N_695,In_4888,In_2462);
nor U696 (N_696,In_3155,In_4185);
nand U697 (N_697,In_1479,In_251);
xnor U698 (N_698,In_4953,In_381);
xnor U699 (N_699,In_956,In_352);
xnor U700 (N_700,In_3891,In_4117);
and U701 (N_701,In_1994,In_1185);
xnor U702 (N_702,In_2221,In_2234);
or U703 (N_703,In_1558,In_4867);
nor U704 (N_704,In_2448,In_1562);
nand U705 (N_705,In_2869,In_3333);
nand U706 (N_706,In_3111,In_3961);
nor U707 (N_707,In_741,In_3656);
xnor U708 (N_708,In_4673,In_1564);
nor U709 (N_709,In_977,In_4288);
xor U710 (N_710,In_1157,In_4424);
or U711 (N_711,In_4479,In_3973);
nor U712 (N_712,In_3131,In_2422);
xnor U713 (N_713,In_546,In_1843);
nand U714 (N_714,In_3098,In_3182);
or U715 (N_715,In_1020,In_1010);
nand U716 (N_716,In_1926,In_680);
xor U717 (N_717,In_3754,In_3206);
and U718 (N_718,In_942,In_553);
and U719 (N_719,In_223,In_4610);
or U720 (N_720,In_2023,In_1127);
and U721 (N_721,In_1070,In_3246);
nor U722 (N_722,In_4937,In_864);
and U723 (N_723,In_1686,In_2115);
and U724 (N_724,In_180,In_3835);
nor U725 (N_725,In_3741,In_3798);
nand U726 (N_726,In_1970,In_3934);
and U727 (N_727,In_2255,In_176);
nor U728 (N_728,In_682,In_1751);
xor U729 (N_729,In_1061,In_195);
or U730 (N_730,In_650,In_4886);
or U731 (N_731,In_575,In_4767);
xnor U732 (N_732,In_112,In_2900);
and U733 (N_733,In_4719,In_3257);
nand U734 (N_734,In_3375,In_2845);
nor U735 (N_735,In_2456,In_4055);
nand U736 (N_736,In_911,In_1517);
xnor U737 (N_737,In_2539,In_3490);
nor U738 (N_738,In_2047,In_1507);
or U739 (N_739,In_1756,In_1074);
nand U740 (N_740,In_1670,In_1563);
nand U741 (N_741,In_2336,In_4734);
or U742 (N_742,In_3411,In_2353);
nor U743 (N_743,In_4038,In_2876);
and U744 (N_744,In_2324,In_3283);
and U745 (N_745,In_2935,In_670);
and U746 (N_746,In_3856,In_2368);
nor U747 (N_747,In_4777,In_3792);
nand U748 (N_748,In_4891,In_2971);
xnor U749 (N_749,In_4075,In_4545);
and U750 (N_750,In_1805,In_3268);
and U751 (N_751,In_2154,In_4973);
nand U752 (N_752,In_1685,In_934);
nor U753 (N_753,In_3564,In_186);
and U754 (N_754,In_831,In_232);
or U755 (N_755,In_145,In_1505);
xor U756 (N_756,In_2780,In_1026);
nor U757 (N_757,In_2359,In_4811);
nand U758 (N_758,In_1669,In_3041);
or U759 (N_759,In_2575,In_483);
nand U760 (N_760,In_2086,In_3734);
xor U761 (N_761,In_1542,In_236);
xor U762 (N_762,In_1386,In_2427);
and U763 (N_763,In_3463,In_3070);
or U764 (N_764,In_4078,In_3273);
nor U765 (N_765,In_3572,In_4505);
or U766 (N_766,In_3616,In_4226);
nand U767 (N_767,In_2404,In_4815);
and U768 (N_768,In_3811,In_395);
xor U769 (N_769,In_143,In_2633);
nor U770 (N_770,In_4461,In_4079);
and U771 (N_771,In_2035,In_2514);
xnor U772 (N_772,In_803,In_1348);
or U773 (N_773,In_102,In_4948);
or U774 (N_774,In_2551,In_4708);
nand U775 (N_775,In_4212,In_3686);
xnor U776 (N_776,In_1888,In_2155);
xnor U777 (N_777,In_1876,In_2811);
or U778 (N_778,In_1209,In_293);
or U779 (N_779,In_4273,In_2648);
xor U780 (N_780,In_2472,In_3955);
nand U781 (N_781,In_1090,In_2968);
xnor U782 (N_782,In_1643,In_1863);
and U783 (N_783,In_1339,In_3701);
nor U784 (N_784,In_1882,In_2754);
or U785 (N_785,In_2342,In_419);
xor U786 (N_786,In_4509,In_278);
nor U787 (N_787,In_3694,In_3648);
nand U788 (N_788,In_4916,In_2482);
xor U789 (N_789,In_451,In_1027);
xnor U790 (N_790,In_3176,In_95);
or U791 (N_791,In_4132,In_3757);
nand U792 (N_792,In_3337,In_2726);
nand U793 (N_793,In_1210,In_333);
or U794 (N_794,In_2716,In_433);
nor U795 (N_795,In_2152,In_3458);
nor U796 (N_796,In_1861,In_3546);
nand U797 (N_797,In_4187,In_4153);
xor U798 (N_798,In_1932,In_3324);
or U799 (N_799,In_3481,In_4914);
or U800 (N_800,In_3046,In_2717);
nor U801 (N_801,In_3519,In_4011);
nor U802 (N_802,In_2138,In_700);
nor U803 (N_803,In_3580,In_3394);
or U804 (N_804,In_698,In_26);
and U805 (N_805,In_3618,In_3742);
nor U806 (N_806,In_1394,In_1849);
nand U807 (N_807,In_1162,In_3560);
or U808 (N_808,In_826,In_898);
and U809 (N_809,In_3899,In_3530);
nor U810 (N_810,In_661,In_3441);
xor U811 (N_811,In_3374,In_916);
xor U812 (N_812,In_1231,In_2817);
nor U813 (N_813,In_175,In_97);
nand U814 (N_814,In_1999,In_1942);
nor U815 (N_815,In_4637,In_1280);
and U816 (N_816,In_3202,In_1000);
or U817 (N_817,In_3039,In_2194);
and U818 (N_818,In_3242,In_4454);
or U819 (N_819,In_2308,In_1739);
and U820 (N_820,In_4320,In_4237);
nand U821 (N_821,In_264,In_168);
xor U822 (N_822,In_3119,In_2618);
or U823 (N_823,In_4658,In_3826);
or U824 (N_824,In_4357,In_1426);
nand U825 (N_825,In_3491,In_736);
or U826 (N_826,In_1763,In_4200);
or U827 (N_827,In_606,In_3159);
nand U828 (N_828,In_1319,In_405);
and U829 (N_829,In_1267,In_3508);
and U830 (N_830,In_3552,In_3274);
nand U831 (N_831,In_2914,In_4971);
or U832 (N_832,In_4398,In_3024);
nor U833 (N_833,In_3755,In_2972);
and U834 (N_834,In_777,In_862);
xnor U835 (N_835,In_2980,In_2694);
or U836 (N_836,In_3631,In_4771);
xnor U837 (N_837,In_3684,In_528);
and U838 (N_838,In_4626,In_273);
nand U839 (N_839,In_4020,In_3071);
nand U840 (N_840,In_4111,In_4706);
xnor U841 (N_841,In_385,In_2500);
and U842 (N_842,In_1334,In_544);
or U843 (N_843,In_4649,In_2991);
and U844 (N_844,In_4566,In_2230);
and U845 (N_845,In_4077,In_1022);
and U846 (N_846,In_3123,In_148);
xnor U847 (N_847,In_2782,In_3872);
and U848 (N_848,In_1381,In_2558);
xnor U849 (N_849,In_2110,In_2100);
xor U850 (N_850,In_3749,In_4524);
xnor U851 (N_851,In_165,In_770);
nor U852 (N_852,In_940,In_702);
nand U853 (N_853,In_6,In_3157);
or U854 (N_854,In_1316,In_1147);
or U855 (N_855,In_4127,In_2256);
or U856 (N_856,In_3918,In_4730);
nand U857 (N_857,In_4992,In_2772);
or U858 (N_858,In_4504,In_3713);
nand U859 (N_859,In_969,In_1466);
or U860 (N_860,In_3397,In_1841);
xnor U861 (N_861,In_1308,In_1978);
nor U862 (N_862,In_3321,In_778);
nor U863 (N_863,In_622,In_2773);
nor U864 (N_864,In_2316,In_3288);
nand U865 (N_865,In_1661,In_3224);
xor U866 (N_866,In_68,In_1956);
nor U867 (N_867,In_4592,In_2475);
nand U868 (N_868,In_20,In_3812);
nor U869 (N_869,In_3895,In_3880);
and U870 (N_870,In_2755,In_2512);
nand U871 (N_871,In_3382,In_1775);
and U872 (N_872,In_1054,In_1624);
nor U873 (N_873,In_4106,In_2329);
and U874 (N_874,In_4301,In_3097);
and U875 (N_875,In_2113,In_1031);
nand U876 (N_876,In_1737,In_2494);
xnor U877 (N_877,In_4588,In_3278);
nand U878 (N_878,In_55,In_979);
xnor U879 (N_879,In_3377,In_2055);
nand U880 (N_880,In_2119,In_4021);
and U881 (N_881,In_4526,In_2503);
xor U882 (N_882,In_1501,In_4548);
or U883 (N_883,In_2383,In_4297);
xnor U884 (N_884,In_3993,In_4878);
nor U885 (N_885,In_105,In_2891);
xnor U886 (N_886,In_2672,In_2292);
or U887 (N_887,In_4023,In_3534);
nand U888 (N_888,In_300,In_212);
xnor U889 (N_889,In_4421,In_1606);
and U890 (N_890,In_781,In_1718);
nor U891 (N_891,In_4378,In_2323);
xor U892 (N_892,In_3737,In_56);
and U893 (N_893,In_3696,In_4098);
nand U894 (N_894,In_1008,In_635);
xor U895 (N_895,In_460,In_4678);
and U896 (N_896,In_3484,In_750);
xor U897 (N_897,In_4460,In_1754);
nand U898 (N_898,In_4361,In_2885);
nand U899 (N_899,In_502,In_4019);
xor U900 (N_900,In_3920,In_516);
and U901 (N_901,In_3428,In_4348);
nand U902 (N_902,In_2818,In_2033);
and U903 (N_903,In_4064,In_3805);
or U904 (N_904,In_1094,In_1633);
xnor U905 (N_905,In_1029,In_677);
and U906 (N_906,In_2605,In_859);
nand U907 (N_907,In_3674,In_1536);
nand U908 (N_908,In_3522,In_1016);
nand U909 (N_909,In_4990,In_3951);
and U910 (N_910,In_3664,In_4808);
or U911 (N_911,In_3991,In_2162);
or U912 (N_912,In_2395,In_1771);
xor U913 (N_913,In_3570,In_2501);
and U914 (N_914,In_4360,In_410);
or U915 (N_915,In_3567,In_4615);
nand U916 (N_916,In_4928,In_2286);
nor U917 (N_917,In_2887,In_4305);
xnor U918 (N_918,In_726,In_4699);
or U919 (N_919,In_1111,In_4686);
nand U920 (N_920,In_2739,In_4439);
xnor U921 (N_921,In_1042,In_629);
nor U922 (N_922,In_2886,In_1683);
and U923 (N_923,In_4898,In_4925);
and U924 (N_924,In_4670,In_3341);
xor U925 (N_925,In_2623,In_4558);
or U926 (N_926,In_1511,In_1907);
nor U927 (N_927,In_3637,In_1593);
nand U928 (N_928,In_1484,In_2070);
nor U929 (N_929,In_1093,In_373);
nand U930 (N_930,In_2902,In_3537);
or U931 (N_931,In_4768,In_1720);
xnor U932 (N_932,In_1503,In_2015);
nor U933 (N_933,In_3286,In_2679);
nor U934 (N_934,In_3193,In_4299);
xnor U935 (N_935,In_2389,In_1637);
nor U936 (N_936,In_4536,In_4000);
nor U937 (N_937,In_4746,In_4772);
xnor U938 (N_938,In_4083,In_3028);
or U939 (N_939,In_667,In_1204);
nor U940 (N_940,In_3435,In_2282);
or U941 (N_941,In_1641,In_3063);
or U942 (N_942,In_3259,In_601);
or U943 (N_943,In_2233,In_4395);
xor U944 (N_944,In_1975,In_4008);
or U945 (N_945,In_4865,In_1879);
nand U946 (N_946,In_96,In_2339);
and U947 (N_947,In_2417,In_303);
and U948 (N_948,In_4745,In_4752);
nor U949 (N_949,In_4096,In_910);
or U950 (N_950,In_3429,In_4248);
nor U951 (N_951,In_4080,In_2406);
nand U952 (N_952,In_887,In_134);
xor U953 (N_953,In_2305,In_3468);
nand U954 (N_954,In_1072,In_3683);
xnor U955 (N_955,In_964,In_4045);
and U956 (N_956,In_4205,In_3276);
nor U957 (N_957,In_3910,In_431);
or U958 (N_958,In_4291,In_1768);
nor U959 (N_959,In_2349,In_1815);
nor U960 (N_960,In_1159,In_42);
nor U961 (N_961,In_3059,In_487);
nand U962 (N_962,In_2372,In_1655);
and U963 (N_963,In_1636,In_4255);
nand U964 (N_964,In_2530,In_2435);
and U965 (N_965,In_4929,In_4053);
xnor U966 (N_966,In_1328,In_4097);
nand U967 (N_967,In_3446,In_4727);
xor U968 (N_968,In_3588,In_1098);
xor U969 (N_969,In_1382,In_2938);
and U970 (N_970,In_740,In_4628);
nor U971 (N_971,In_3012,In_1108);
and U972 (N_972,In_1425,In_4326);
xor U973 (N_973,In_1383,In_2011);
and U974 (N_974,In_1680,In_970);
xor U975 (N_975,In_2532,In_4784);
nand U976 (N_976,In_556,In_3163);
or U977 (N_977,In_3514,In_462);
and U978 (N_978,In_2108,In_4995);
and U979 (N_979,In_509,In_4907);
xnor U980 (N_980,In_2854,In_2895);
or U981 (N_981,In_4394,In_3788);
and U982 (N_982,In_2683,In_1106);
or U983 (N_983,In_4480,In_3280);
xor U984 (N_984,In_3077,In_196);
and U985 (N_985,In_1028,In_4542);
xnor U986 (N_986,In_4296,In_4676);
and U987 (N_987,In_4231,In_82);
nor U988 (N_988,In_3110,In_3988);
and U989 (N_989,In_2596,In_1747);
nor U990 (N_990,In_4845,In_636);
and U991 (N_991,In_535,In_3040);
and U992 (N_992,In_1532,In_2808);
or U993 (N_993,In_2852,In_2021);
or U994 (N_994,In_3725,In_4864);
xor U995 (N_995,In_3289,In_99);
and U996 (N_996,In_4206,In_4093);
and U997 (N_997,In_4970,In_3381);
or U998 (N_998,In_2552,In_4492);
nor U999 (N_999,In_3387,In_1835);
nor U1000 (N_1000,In_1894,In_1571);
or U1001 (N_1001,In_2725,In_384);
nor U1002 (N_1002,In_4591,In_446);
xor U1003 (N_1003,In_3677,In_1962);
or U1004 (N_1004,In_4478,In_90);
nand U1005 (N_1005,In_3705,In_3232);
nand U1006 (N_1006,In_3512,In_3547);
xnor U1007 (N_1007,In_4114,In_230);
xnor U1008 (N_1008,In_428,In_3237);
nor U1009 (N_1009,In_2248,In_3354);
and U1010 (N_1010,In_3198,In_298);
xor U1011 (N_1011,In_3709,In_1198);
nand U1012 (N_1012,In_2109,In_2429);
xnor U1013 (N_1013,In_3972,In_1050);
xnor U1014 (N_1014,In_493,In_1668);
or U1015 (N_1015,In_3501,In_3793);
xor U1016 (N_1016,In_1796,In_1819);
or U1017 (N_1017,In_932,In_3017);
or U1018 (N_1018,In_1728,In_4573);
nor U1019 (N_1019,In_202,In_4451);
and U1020 (N_1020,In_725,In_1695);
nand U1021 (N_1021,In_292,In_4841);
or U1022 (N_1022,In_1445,In_2792);
nand U1023 (N_1023,In_1252,In_127);
and U1024 (N_1024,In_1595,In_359);
nor U1025 (N_1025,In_2477,In_790);
or U1026 (N_1026,In_2487,In_3628);
and U1027 (N_1027,In_880,In_124);
or U1028 (N_1028,In_3005,In_4996);
nor U1029 (N_1029,In_1266,In_4840);
nand U1030 (N_1030,In_121,In_1904);
nor U1031 (N_1031,In_3390,In_999);
and U1032 (N_1032,In_3774,In_3941);
nand U1033 (N_1033,In_3884,In_191);
nand U1034 (N_1034,In_3335,In_1663);
nor U1035 (N_1035,In_3209,In_1342);
or U1036 (N_1036,In_759,In_4056);
xnor U1037 (N_1037,In_2129,In_4074);
nor U1038 (N_1038,In_447,In_1116);
nor U1039 (N_1039,In_1058,In_2051);
xnor U1040 (N_1040,In_3744,In_3372);
and U1041 (N_1041,In_3497,In_2591);
or U1042 (N_1042,In_4195,In_3050);
xor U1043 (N_1043,In_4930,In_3000);
xnor U1044 (N_1044,In_687,In_3022);
nand U1045 (N_1045,In_4585,In_4969);
nor U1046 (N_1046,In_3087,In_876);
xnor U1047 (N_1047,In_4842,In_4198);
xor U1048 (N_1048,In_1881,In_3655);
or U1049 (N_1049,In_525,In_4627);
xor U1050 (N_1050,In_1129,In_2836);
or U1051 (N_1051,In_3223,In_1590);
or U1052 (N_1052,In_4787,In_2471);
nand U1053 (N_1053,In_131,In_4890);
or U1054 (N_1054,In_768,In_1520);
nand U1055 (N_1055,In_1744,In_3115);
nor U1056 (N_1056,In_3079,In_3026);
or U1057 (N_1057,In_4177,In_4874);
xor U1058 (N_1058,In_952,In_4316);
or U1059 (N_1059,In_1456,In_122);
xor U1060 (N_1060,In_3451,In_3874);
and U1061 (N_1061,In_3344,In_1523);
nor U1062 (N_1062,In_2673,In_1059);
xor U1063 (N_1063,In_4217,In_4798);
or U1064 (N_1064,In_1585,In_4809);
xnor U1065 (N_1065,In_3228,In_1015);
nand U1066 (N_1066,In_4184,In_950);
or U1067 (N_1067,In_3216,In_2457);
nor U1068 (N_1068,In_1084,In_1457);
and U1069 (N_1069,In_1788,In_3204);
nand U1070 (N_1070,In_1195,In_584);
nor U1071 (N_1071,In_2203,In_4049);
and U1072 (N_1072,In_4414,In_3401);
xor U1073 (N_1073,In_2553,In_3437);
xor U1074 (N_1074,In_379,In_174);
and U1075 (N_1075,In_4036,In_1874);
xor U1076 (N_1076,In_1736,In_694);
nor U1077 (N_1077,In_4456,In_1527);
xor U1078 (N_1078,In_1071,In_1400);
nand U1079 (N_1079,In_4684,In_3645);
or U1080 (N_1080,In_1240,In_3244);
nand U1081 (N_1081,In_2764,In_3594);
or U1082 (N_1082,In_2351,In_1338);
nor U1083 (N_1083,In_4467,In_2794);
nand U1084 (N_1084,In_4400,In_2244);
and U1085 (N_1085,In_4050,In_1260);
nand U1086 (N_1086,In_894,In_4687);
xnor U1087 (N_1087,In_1635,In_156);
and U1088 (N_1088,In_1553,In_807);
xor U1089 (N_1089,In_801,In_594);
nand U1090 (N_1090,In_4362,In_4489);
xor U1091 (N_1091,In_3277,In_288);
xor U1092 (N_1092,In_387,In_281);
nor U1093 (N_1093,In_2635,In_3592);
and U1094 (N_1094,In_1707,In_4160);
xnor U1095 (N_1095,In_2328,In_2546);
and U1096 (N_1096,In_3442,In_244);
nand U1097 (N_1097,In_705,In_814);
or U1098 (N_1098,In_1529,In_3453);
nand U1099 (N_1099,In_4605,In_1327);
xnor U1100 (N_1100,In_454,In_522);
xnor U1101 (N_1101,In_476,In_1440);
and U1102 (N_1102,In_2942,In_88);
nor U1103 (N_1103,In_3350,In_4163);
xor U1104 (N_1104,In_204,In_3551);
xor U1105 (N_1105,In_2554,In_12);
xor U1106 (N_1106,In_1053,In_4356);
xnor U1107 (N_1107,In_2646,In_4209);
nor U1108 (N_1108,In_2741,In_2557);
and U1109 (N_1109,In_4383,In_666);
nand U1110 (N_1110,In_3049,In_2925);
xor U1111 (N_1111,In_2535,In_1864);
xor U1112 (N_1112,In_1842,In_2295);
nand U1113 (N_1113,In_166,In_593);
nor U1114 (N_1114,In_83,In_4457);
nand U1115 (N_1115,In_1325,In_4742);
or U1116 (N_1116,In_16,In_4330);
or U1117 (N_1117,In_457,In_2048);
and U1118 (N_1118,In_4452,In_4910);
or U1119 (N_1119,In_3055,In_2084);
and U1120 (N_1120,In_2093,In_1048);
and U1121 (N_1121,In_1431,In_2583);
and U1122 (N_1122,In_802,In_4384);
or U1123 (N_1123,In_1192,In_2062);
or U1124 (N_1124,In_2729,In_4755);
and U1125 (N_1125,In_412,In_570);
xnor U1126 (N_1126,In_2141,In_749);
and U1127 (N_1127,In_1496,In_2246);
or U1128 (N_1128,In_4718,In_1439);
xnor U1129 (N_1129,In_2883,In_1420);
nor U1130 (N_1130,In_545,In_3091);
xor U1131 (N_1131,In_3804,In_4756);
nor U1132 (N_1132,In_2529,In_1207);
nand U1133 (N_1133,In_3916,In_1454);
or U1134 (N_1134,In_2441,In_1153);
xnor U1135 (N_1135,In_4029,In_1512);
nand U1136 (N_1136,In_2680,In_2958);
nor U1137 (N_1137,In_2617,In_4551);
nand U1138 (N_1138,In_521,In_974);
or U1139 (N_1139,In_1508,In_2896);
xor U1140 (N_1140,In_3060,In_321);
and U1141 (N_1141,In_2582,In_2038);
nand U1142 (N_1142,In_3067,In_3598);
nand U1143 (N_1143,In_2117,In_640);
and U1144 (N_1144,In_2402,In_365);
xnor U1145 (N_1145,In_3761,In_3472);
and U1146 (N_1146,In_2727,In_1567);
xnor U1147 (N_1147,In_4726,In_4024);
and U1148 (N_1148,In_3313,In_2776);
xnor U1149 (N_1149,In_3296,In_1488);
nand U1150 (N_1150,In_267,In_4112);
or U1151 (N_1151,In_1133,In_2455);
xor U1152 (N_1152,In_349,In_3885);
xor U1153 (N_1153,In_2414,In_1398);
nor U1154 (N_1154,In_2220,In_272);
nand U1155 (N_1155,In_981,In_2334);
xnor U1156 (N_1156,In_2995,In_61);
and U1157 (N_1157,In_3502,In_3426);
nor U1158 (N_1158,In_1826,In_3896);
or U1159 (N_1159,In_3129,In_4131);
or U1160 (N_1160,In_2916,In_2276);
or U1161 (N_1161,In_2374,In_3207);
or U1162 (N_1162,In_937,In_4119);
nor U1163 (N_1163,In_820,In_1504);
nor U1164 (N_1164,In_2146,In_2412);
nand U1165 (N_1165,In_829,In_893);
nand U1166 (N_1166,In_2795,In_4797);
xnor U1167 (N_1167,In_2816,In_2018);
and U1168 (N_1168,In_800,In_2191);
or U1169 (N_1169,In_737,In_1617);
nor U1170 (N_1170,In_3892,In_1105);
and U1171 (N_1171,In_3391,In_819);
nor U1172 (N_1172,In_197,In_2158);
xor U1173 (N_1173,In_4312,In_1290);
or U1174 (N_1174,In_2733,In_3094);
nand U1175 (N_1175,In_2311,In_2237);
nor U1176 (N_1176,In_2045,In_227);
nor U1177 (N_1177,In_2388,In_1865);
nand U1178 (N_1178,In_4681,In_2807);
nand U1179 (N_1179,In_3359,In_4582);
xor U1180 (N_1180,In_2279,In_1992);
and U1181 (N_1181,In_2452,In_2058);
xnor U1182 (N_1182,In_2674,In_3322);
nand U1183 (N_1183,In_371,In_1628);
or U1184 (N_1184,In_4783,In_282);
xor U1185 (N_1185,In_4263,In_721);
and U1186 (N_1186,In_2718,In_3287);
nand U1187 (N_1187,In_441,In_2970);
xnor U1188 (N_1188,In_4871,In_4760);
xor U1189 (N_1189,In_4364,In_2868);
nor U1190 (N_1190,In_4781,In_3214);
nand U1191 (N_1191,In_2701,In_649);
nand U1192 (N_1192,In_1619,In_3118);
or U1193 (N_1193,In_1599,In_2509);
or U1194 (N_1194,In_4713,In_531);
or U1195 (N_1195,In_2285,In_2296);
nor U1196 (N_1196,In_2091,In_1832);
xor U1197 (N_1197,In_177,In_4535);
nand U1198 (N_1198,In_3765,In_4370);
or U1199 (N_1199,In_126,In_1264);
xor U1200 (N_1200,In_780,In_4924);
nand U1201 (N_1201,In_3938,In_3);
or U1202 (N_1202,In_861,In_4001);
and U1203 (N_1203,In_2382,In_1244);
or U1204 (N_1204,In_3911,In_4068);
and U1205 (N_1205,In_247,In_3888);
nand U1206 (N_1206,In_1950,In_366);
xor U1207 (N_1207,In_2013,In_3615);
nand U1208 (N_1208,In_3188,In_1510);
and U1209 (N_1209,In_4968,In_4795);
or U1210 (N_1210,In_2750,In_1409);
and U1211 (N_1211,In_2563,In_2087);
xnor U1212 (N_1212,In_564,In_4373);
or U1213 (N_1213,In_3587,In_3970);
or U1214 (N_1214,In_4241,In_2959);
nor U1215 (N_1215,In_1672,In_2697);
nand U1216 (N_1216,In_4698,In_2939);
nor U1217 (N_1217,In_689,In_1131);
or U1218 (N_1218,In_3671,In_4041);
and U1219 (N_1219,In_1939,In_1483);
nor U1220 (N_1220,In_1432,In_342);
and U1221 (N_1221,In_231,In_2711);
xnor U1222 (N_1222,In_1448,In_2687);
nand U1223 (N_1223,In_2262,In_2927);
nor U1224 (N_1224,In_825,In_946);
nor U1225 (N_1225,In_2097,In_4094);
nand U1226 (N_1226,In_3496,In_3054);
nand U1227 (N_1227,In_1417,In_1873);
nand U1228 (N_1228,In_448,In_2783);
nand U1229 (N_1229,In_752,In_2189);
nor U1230 (N_1230,In_1765,In_3649);
xor U1231 (N_1231,In_1142,In_2193);
nor U1232 (N_1232,In_75,In_3781);
nor U1233 (N_1233,In_2467,In_1434);
nor U1234 (N_1234,In_475,In_2989);
or U1235 (N_1235,In_4801,In_1139);
nand U1236 (N_1236,In_2547,In_1079);
and U1237 (N_1237,In_2923,In_2354);
or U1238 (N_1238,In_4527,In_3736);
nand U1239 (N_1239,In_1269,In_43);
xor U1240 (N_1240,In_4487,In_2621);
xor U1241 (N_1241,In_207,In_2423);
nand U1242 (N_1242,In_908,In_1993);
or U1243 (N_1243,In_2665,In_4901);
nand U1244 (N_1244,In_883,In_1937);
nor U1245 (N_1245,In_2075,In_4063);
and U1246 (N_1246,In_3361,In_2275);
and U1247 (N_1247,In_2746,In_60);
or U1248 (N_1248,In_878,In_1156);
nand U1249 (N_1249,In_2160,In_4051);
nand U1250 (N_1250,In_3935,In_4758);
nor U1251 (N_1251,In_4774,In_1443);
xnor U1252 (N_1252,In_4159,In_347);
nor U1253 (N_1253,In_2698,In_4614);
or U1254 (N_1254,In_3235,In_4437);
or U1255 (N_1255,In_4617,In_1989);
or U1256 (N_1256,In_1878,In_4221);
xnor U1257 (N_1257,In_2076,In_149);
nand U1258 (N_1258,In_2677,In_2077);
and U1259 (N_1259,In_3264,In_2948);
or U1260 (N_1260,In_2195,In_2724);
or U1261 (N_1261,In_1491,In_4736);
nand U1262 (N_1262,In_4887,In_1243);
xor U1263 (N_1263,In_4335,In_417);
nand U1264 (N_1264,In_2576,In_4938);
or U1265 (N_1265,In_18,In_2560);
nor U1266 (N_1266,In_3878,In_2209);
and U1267 (N_1267,In_1166,In_3731);
nand U1268 (N_1268,In_4458,In_4342);
nor U1269 (N_1269,In_3241,In_128);
or U1270 (N_1270,In_1896,In_4007);
or U1271 (N_1271,In_4812,In_3864);
or U1272 (N_1272,In_392,In_3599);
nand U1273 (N_1273,In_4561,In_229);
nor U1274 (N_1274,In_4618,In_656);
nand U1275 (N_1275,In_3367,In_3275);
nand U1276 (N_1276,In_4635,In_11);
xor U1277 (N_1277,In_2006,In_1032);
xor U1278 (N_1278,In_973,In_791);
or U1279 (N_1279,In_1556,In_760);
nand U1280 (N_1280,In_900,In_1073);
nand U1281 (N_1281,In_193,In_3723);
nand U1282 (N_1282,In_4512,In_882);
nor U1283 (N_1283,In_2190,In_2786);
and U1284 (N_1284,In_2358,In_3270);
nand U1285 (N_1285,In_3566,In_329);
nor U1286 (N_1286,In_3800,In_4560);
and U1287 (N_1287,In_1455,In_3827);
and U1288 (N_1288,In_3604,In_3431);
xnor U1289 (N_1289,In_957,In_2645);
nand U1290 (N_1290,In_621,In_1675);
nand U1291 (N_1291,In_4353,In_3840);
nor U1292 (N_1292,In_2229,In_587);
nor U1293 (N_1293,In_3652,In_1774);
or U1294 (N_1294,In_3388,In_3852);
nor U1295 (N_1295,In_4595,In_357);
or U1296 (N_1296,In_2922,In_3927);
or U1297 (N_1297,In_3238,In_213);
nand U1298 (N_1298,In_3467,In_4765);
nor U1299 (N_1299,In_663,In_3465);
or U1300 (N_1300,In_2853,In_4175);
nor U1301 (N_1301,In_4017,In_4902);
or U1302 (N_1302,In_647,In_1055);
xnor U1303 (N_1303,In_378,In_4792);
or U1304 (N_1304,In_54,In_3421);
or U1305 (N_1305,In_1884,In_2136);
xnor U1306 (N_1306,In_1509,In_1311);
or U1307 (N_1307,In_573,In_637);
nand U1308 (N_1308,In_3011,In_2177);
nand U1309 (N_1309,In_4333,In_1265);
or U1310 (N_1310,In_4169,In_2019);
nor U1311 (N_1311,In_3336,In_971);
and U1312 (N_1312,In_3981,In_3403);
xor U1313 (N_1313,In_4763,In_5);
nor U1314 (N_1314,In_2577,In_709);
nand U1315 (N_1315,In_2842,In_2721);
nor U1316 (N_1316,In_2106,In_2587);
nor U1317 (N_1317,In_445,In_1199);
nor U1318 (N_1318,In_4,In_4912);
and U1319 (N_1319,In_3751,In_1326);
nor U1320 (N_1320,In_3946,In_4802);
nand U1321 (N_1321,In_1492,In_2361);
and U1322 (N_1322,In_1551,In_284);
xor U1323 (N_1323,In_51,In_2223);
or U1324 (N_1324,In_3056,In_4508);
and U1325 (N_1325,In_929,In_1891);
xnor U1326 (N_1326,In_1804,In_3777);
nor U1327 (N_1327,In_4385,In_2877);
nor U1328 (N_1328,In_3659,In_1664);
and U1329 (N_1329,In_271,In_4203);
xor U1330 (N_1330,In_3073,In_4411);
nand U1331 (N_1331,In_1866,In_3393);
and U1332 (N_1332,In_2610,In_717);
and U1333 (N_1333,In_2251,In_4712);
nand U1334 (N_1334,In_4915,In_1041);
xnor U1335 (N_1335,In_4562,In_4935);
and U1336 (N_1336,In_4715,In_1261);
or U1337 (N_1337,In_2392,In_4540);
or U1338 (N_1338,In_2647,In_4164);
nor U1339 (N_1339,In_2752,In_4317);
or U1340 (N_1340,In_4757,In_3099);
nor U1341 (N_1341,In_3400,In_3558);
xnor U1342 (N_1342,In_1187,In_2239);
nor U1343 (N_1343,In_1915,In_1976);
nand U1344 (N_1344,In_1545,In_1981);
or U1345 (N_1345,In_4735,In_458);
and U1346 (N_1346,In_2767,In_3853);
nand U1347 (N_1347,In_4897,In_1794);
nor U1348 (N_1348,In_1900,In_2344);
or U1349 (N_1349,In_2598,In_713);
or U1350 (N_1350,In_362,In_1611);
nand U1351 (N_1351,In_3127,In_2658);
nor U1352 (N_1352,In_1305,In_2016);
nand U1353 (N_1353,In_603,In_3773);
nand U1354 (N_1354,In_4964,In_76);
and U1355 (N_1355,In_4247,In_4393);
nor U1356 (N_1356,In_4940,In_623);
or U1357 (N_1357,In_52,In_1242);
nor U1358 (N_1358,In_4058,In_4722);
nand U1359 (N_1359,In_975,In_4528);
or U1360 (N_1360,In_706,In_1320);
and U1361 (N_1361,In_1134,In_2312);
or U1362 (N_1362,In_2950,In_4448);
nand U1363 (N_1363,In_2920,In_729);
nor U1364 (N_1364,In_1555,In_115);
or U1365 (N_1365,In_4942,In_4818);
and U1366 (N_1366,In_1825,In_429);
and U1367 (N_1367,In_2986,In_913);
or U1368 (N_1368,In_3627,In_2224);
and U1369 (N_1369,In_1753,In_2394);
nor U1370 (N_1370,In_1374,In_1360);
and U1371 (N_1371,In_1858,In_4833);
xor U1372 (N_1372,In_665,In_15);
or U1373 (N_1373,In_369,In_4835);
or U1374 (N_1374,In_4165,In_4688);
and U1375 (N_1375,In_1276,In_2227);
or U1376 (N_1376,In_994,In_101);
and U1377 (N_1377,In_3282,In_4549);
nor U1378 (N_1378,In_2931,In_4705);
nand U1379 (N_1379,In_1114,In_4476);
or U1380 (N_1380,In_3243,In_425);
or U1381 (N_1381,In_3687,In_874);
xor U1382 (N_1382,In_3987,In_3553);
xor U1383 (N_1383,In_3386,In_2073);
xnor U1384 (N_1384,In_3433,In_2173);
or U1385 (N_1385,In_4293,In_933);
and U1386 (N_1386,In_3707,In_3584);
or U1387 (N_1387,In_1885,In_291);
and U1388 (N_1388,In_2367,In_1640);
or U1389 (N_1389,In_2092,In_4943);
nand U1390 (N_1390,In_1887,In_1238);
nand U1391 (N_1391,In_822,In_1911);
or U1392 (N_1392,In_2636,In_1184);
nor U1393 (N_1393,In_3137,In_2693);
or U1394 (N_1394,In_3695,In_3775);
and U1395 (N_1395,In_4799,In_2204);
or U1396 (N_1396,In_116,In_4147);
and U1397 (N_1397,In_3536,In_3146);
xor U1398 (N_1398,In_4520,In_3980);
or U1399 (N_1399,In_907,In_4115);
nor U1400 (N_1400,In_1708,In_1373);
xor U1401 (N_1401,In_1190,In_2999);
and U1402 (N_1402,In_2555,In_2365);
and U1403 (N_1403,In_3579,In_221);
nand U1404 (N_1404,In_4133,In_2656);
and U1405 (N_1405,In_1299,In_3415);
xnor U1406 (N_1406,In_4308,In_538);
nor U1407 (N_1407,In_2600,In_1554);
and U1408 (N_1408,In_1830,In_511);
and U1409 (N_1409,In_4148,In_3839);
xnor U1410 (N_1410,In_2912,In_941);
xnor U1411 (N_1411,In_336,In_205);
nor U1412 (N_1412,In_4048,In_2759);
xnor U1413 (N_1413,In_390,In_2651);
or U1414 (N_1414,In_1499,In_3018);
nor U1415 (N_1415,In_2425,In_3703);
or U1416 (N_1416,In_4550,In_397);
nand U1417 (N_1417,In_4851,In_2857);
nor U1418 (N_1418,In_1586,In_1375);
xor U1419 (N_1419,In_2450,In_2491);
xor U1420 (N_1420,In_3817,In_1087);
nand U1421 (N_1421,In_3169,In_92);
or U1422 (N_1422,In_3661,In_4358);
nand U1423 (N_1423,In_361,In_3743);
nand U1424 (N_1424,In_2208,In_4525);
nand U1425 (N_1425,In_657,In_1724);
nor U1426 (N_1426,In_2615,In_250);
nand U1427 (N_1427,In_4328,In_1126);
xnor U1428 (N_1428,In_872,In_1767);
and U1429 (N_1429,In_3538,In_2240);
nor U1430 (N_1430,In_664,In_3905);
nand U1431 (N_1431,In_1892,In_2031);
nand U1432 (N_1432,In_3565,In_519);
nand U1433 (N_1433,In_1588,In_2283);
nor U1434 (N_1434,In_4613,In_851);
and U1435 (N_1435,In_897,In_3001);
or U1436 (N_1436,In_89,In_1128);
nand U1437 (N_1437,In_1007,In_4949);
or U1438 (N_1438,In_146,In_3917);
nor U1439 (N_1439,In_1625,In_1201);
xnor U1440 (N_1440,In_1487,In_3215);
and U1441 (N_1441,In_49,In_1013);
nand U1442 (N_1442,In_4430,In_2505);
or U1443 (N_1443,In_4653,In_3609);
and U1444 (N_1444,In_3256,In_3596);
and U1445 (N_1445,In_2293,In_817);
nand U1446 (N_1446,In_2469,In_187);
nand U1447 (N_1447,In_4827,In_2619);
nor U1448 (N_1448,In_2940,In_505);
xor U1449 (N_1449,In_1324,In_3762);
or U1450 (N_1450,In_1965,In_2996);
nand U1451 (N_1451,In_4188,In_1168);
and U1452 (N_1452,In_526,In_2918);
xor U1453 (N_1453,In_4744,In_2440);
or U1454 (N_1454,In_4359,In_2040);
or U1455 (N_1455,In_2804,In_2898);
nand U1456 (N_1456,In_4593,In_4346);
xor U1457 (N_1457,In_4258,In_905);
or U1458 (N_1458,In_1271,In_3405);
nand U1459 (N_1459,In_58,In_4711);
xnor U1460 (N_1460,In_4857,In_612);
or U1461 (N_1461,In_3504,In_2534);
nand U1462 (N_1462,In_2682,In_3492);
nand U1463 (N_1463,In_1418,In_1631);
nor U1464 (N_1464,In_3105,In_490);
and U1465 (N_1465,In_4152,In_4531);
nand U1466 (N_1466,In_1427,In_3262);
nand U1467 (N_1467,In_2562,In_2219);
and U1468 (N_1468,In_2542,In_2096);
nor U1469 (N_1469,In_1935,In_4179);
nand U1470 (N_1470,In_1284,In_7);
nand U1471 (N_1471,In_2977,In_1731);
nand U1472 (N_1472,In_1671,In_2386);
or U1473 (N_1473,In_1659,In_2135);
and U1474 (N_1474,In_1867,In_4674);
nor U1475 (N_1475,In_2166,In_3894);
xor U1476 (N_1476,In_1372,In_4790);
nand U1477 (N_1477,In_743,In_793);
nand U1478 (N_1478,In_4107,In_4695);
xor U1479 (N_1479,In_2785,In_4054);
and U1480 (N_1480,In_335,In_2366);
and U1481 (N_1481,In_877,In_3768);
nand U1482 (N_1482,In_686,In_3675);
xnor U1483 (N_1483,In_582,In_2707);
nand U1484 (N_1484,In_4057,In_4376);
and U1485 (N_1485,In_4927,In_3179);
xnor U1486 (N_1486,In_3858,In_1506);
or U1487 (N_1487,In_1344,In_2089);
nor U1488 (N_1488,In_2867,In_4016);
xnor U1489 (N_1489,In_4199,In_1537);
or U1490 (N_1490,In_503,In_2044);
xor U1491 (N_1491,In_4386,In_1883);
and U1492 (N_1492,In_210,In_1931);
or U1493 (N_1493,In_4110,In_4951);
or U1494 (N_1494,In_4979,In_1451);
xnor U1495 (N_1495,In_610,In_4279);
nand U1496 (N_1496,In_3248,In_3608);
nor U1497 (N_1497,In_2580,In_3636);
or U1498 (N_1498,In_2669,In_2837);
nand U1499 (N_1499,In_312,In_3327);
xnor U1500 (N_1500,In_3545,In_1847);
nand U1501 (N_1501,In_2356,In_722);
and U1502 (N_1502,In_1581,In_1202);
or U1503 (N_1503,In_3926,In_2880);
xor U1504 (N_1504,In_4829,In_3965);
xor U1505 (N_1505,In_3457,In_4717);
nor U1506 (N_1506,In_2235,In_25);
nor U1507 (N_1507,In_3693,In_2298);
and U1508 (N_1508,In_1941,In_718);
nand U1509 (N_1509,In_2433,In_4539);
nor U1510 (N_1510,In_2987,In_1051);
or U1511 (N_1511,In_1036,In_4272);
nand U1512 (N_1512,In_4380,In_2643);
and U1513 (N_1513,In_1323,In_2652);
nor U1514 (N_1514,In_4496,In_1174);
nor U1515 (N_1515,In_4922,In_2766);
nand U1516 (N_1516,In_2319,In_3103);
xnor U1517 (N_1517,In_1502,In_2156);
nand U1518 (N_1518,In_615,In_233);
nand U1519 (N_1519,In_1500,In_4109);
nor U1520 (N_1520,In_3006,In_3132);
nand U1521 (N_1521,In_1584,In_3654);
or U1522 (N_1522,In_1698,In_265);
xnor U1523 (N_1523,In_209,In_2265);
or U1524 (N_1524,In_2090,In_3036);
nand U1525 (N_1525,In_4761,In_4672);
nor U1526 (N_1526,In_3915,In_1421);
or U1527 (N_1527,In_1886,In_1854);
nor U1528 (N_1528,In_3414,In_325);
nor U1529 (N_1529,In_422,In_1521);
xor U1530 (N_1530,In_2819,In_4446);
xor U1531 (N_1531,In_3161,In_879);
xor U1532 (N_1532,In_4709,In_4600);
xor U1533 (N_1533,In_4125,In_1304);
nand U1534 (N_1534,In_4931,In_4224);
xor U1535 (N_1535,In_1152,In_959);
and U1536 (N_1536,In_625,In_1438);
nor U1537 (N_1537,In_2192,In_2133);
nor U1538 (N_1538,In_1470,In_3151);
nor U1539 (N_1539,In_3373,In_3075);
or U1540 (N_1540,In_1791,In_123);
xor U1541 (N_1541,In_972,In_2926);
xnor U1542 (N_1542,In_627,In_178);
xnor U1543 (N_1543,In_4251,In_3452);
or U1544 (N_1544,In_3258,In_751);
and U1545 (N_1545,In_2281,In_4280);
nor U1546 (N_1546,In_855,In_4310);
or U1547 (N_1547,In_1954,In_4723);
or U1548 (N_1548,In_3971,In_3160);
xnor U1549 (N_1549,In_4076,In_2700);
nor U1550 (N_1550,In_580,In_469);
or U1551 (N_1551,In_1169,In_3058);
xor U1552 (N_1552,In_3555,In_4140);
xnor U1553 (N_1553,In_554,In_3104);
xnor U1554 (N_1554,In_3461,In_2676);
nor U1555 (N_1555,In_1229,In_1468);
or U1556 (N_1556,In_107,In_1711);
nor U1557 (N_1557,In_4782,In_3053);
or U1558 (N_1558,In_4848,In_106);
nor U1559 (N_1559,In_2054,In_4866);
nor U1560 (N_1560,In_643,In_1329);
nor U1561 (N_1561,In_4604,In_3989);
nand U1562 (N_1562,In_2522,In_732);
or U1563 (N_1563,In_2122,In_3622);
nand U1564 (N_1564,In_309,In_1005);
nand U1565 (N_1565,In_2480,In_1752);
or U1566 (N_1566,In_1197,In_4246);
or U1567 (N_1567,In_2022,In_189);
nor U1568 (N_1568,In_840,In_552);
and U1569 (N_1569,In_1693,In_2838);
or U1570 (N_1570,In_3141,In_2809);
or U1571 (N_1571,In_4243,In_4703);
or U1572 (N_1572,In_4494,In_3185);
nand U1573 (N_1573,In_320,In_3309);
and U1574 (N_1574,In_4092,In_2226);
nand U1575 (N_1575,In_1985,In_3212);
and U1576 (N_1576,In_3014,In_3509);
nand U1577 (N_1577,In_172,In_1871);
xor U1578 (N_1578,In_2641,In_1318);
and U1579 (N_1579,In_3745,In_241);
xor U1580 (N_1580,In_3865,In_316);
xnor U1581 (N_1581,In_532,In_3150);
nor U1582 (N_1582,In_1714,In_3691);
nor U1583 (N_1583,In_1656,In_1004);
xnor U1584 (N_1584,In_3378,In_1387);
xnor U1585 (N_1585,In_4047,In_1254);
and U1586 (N_1586,In_1583,In_3101);
or U1587 (N_1587,In_2978,In_4464);
xnor U1588 (N_1588,In_4849,In_4881);
nor U1589 (N_1589,In_2829,In_4576);
nand U1590 (N_1590,In_617,In_2069);
and U1591 (N_1591,In_1021,In_1607);
nor U1592 (N_1592,In_3506,In_4355);
or U1593 (N_1593,In_1165,In_4819);
xor U1594 (N_1594,In_1183,In_435);
or U1595 (N_1595,In_2474,In_2355);
nand U1596 (N_1596,In_98,In_1594);
and U1597 (N_1597,In_3979,In_2478);
xnor U1598 (N_1598,In_3966,In_438);
nand U1599 (N_1599,In_4956,In_782);
nor U1600 (N_1600,In_3722,In_3607);
xnor U1601 (N_1601,In_1362,In_1807);
xnor U1602 (N_1602,In_885,In_194);
nand U1603 (N_1603,In_3606,In_4751);
or U1604 (N_1604,In_785,In_3952);
nand U1605 (N_1605,In_2735,In_1938);
nor U1606 (N_1606,In_4789,In_2517);
and U1607 (N_1607,In_4960,In_2690);
xnor U1608 (N_1608,In_3348,In_4872);
and U1609 (N_1609,In_430,In_1930);
nor U1610 (N_1610,In_2258,In_4440);
or U1611 (N_1611,In_1397,In_1851);
nand U1612 (N_1612,In_1001,In_3726);
nor U1613 (N_1613,In_2969,In_41);
or U1614 (N_1614,In_1658,In_1228);
nand U1615 (N_1615,In_489,In_1388);
and U1616 (N_1616,In_1869,In_4883);
xnor U1617 (N_1617,In_3225,In_2180);
nand U1618 (N_1618,In_4846,In_2401);
nor U1619 (N_1619,In_4409,In_962);
nand U1620 (N_1620,In_3038,In_508);
nand U1621 (N_1621,In_4982,In_2380);
nor U1622 (N_1622,In_1848,In_4201);
and U1623 (N_1623,In_1963,In_676);
nor U1624 (N_1624,In_2481,In_1961);
nor U1625 (N_1625,In_2357,In_4104);
or U1626 (N_1626,In_1399,In_1194);
nand U1627 (N_1627,In_249,In_3083);
and U1628 (N_1628,In_2302,In_3542);
or U1629 (N_1629,In_4515,In_1844);
xor U1630 (N_1630,In_2307,In_915);
nand U1631 (N_1631,In_276,In_4031);
nor U1632 (N_1632,In_2321,In_951);
nand U1633 (N_1633,In_2254,In_1232);
or U1634 (N_1634,In_1898,In_239);
nand U1635 (N_1635,In_2941,In_998);
nand U1636 (N_1636,In_1918,In_1078);
and U1637 (N_1637,In_3883,In_744);
nor U1638 (N_1638,In_4138,In_3505);
and U1639 (N_1639,In_3002,In_285);
nand U1640 (N_1640,In_4345,In_1665);
or U1641 (N_1641,In_4495,In_1351);
nand U1642 (N_1642,In_1650,In_2892);
nand U1643 (N_1643,In_4733,In_2624);
or U1644 (N_1644,In_4936,In_4895);
nand U1645 (N_1645,In_1273,In_734);
nor U1646 (N_1646,In_3520,In_3619);
nand U1647 (N_1647,In_4043,In_2839);
nand U1648 (N_1648,In_1091,In_3355);
xnor U1649 (N_1649,In_1045,In_1991);
nor U1650 (N_1650,In_2985,In_2370);
xnor U1651 (N_1651,In_1936,In_4580);
xnor U1652 (N_1652,In_1356,In_539);
and U1653 (N_1653,In_968,In_4202);
or U1654 (N_1654,In_2473,In_255);
xnor U1655 (N_1655,In_4570,In_3842);
nand U1656 (N_1656,In_169,In_80);
and U1657 (N_1657,In_1392,In_4662);
and U1658 (N_1658,In_2181,In_3475);
nand U1659 (N_1659,In_3045,In_3923);
and U1660 (N_1660,In_2788,In_3620);
nand U1661 (N_1661,In_671,In_4227);
xor U1662 (N_1662,In_1694,In_2416);
or U1663 (N_1663,In_4606,In_2848);
or U1664 (N_1664,In_34,In_1477);
nand U1665 (N_1665,In_4425,In_4146);
xor U1666 (N_1666,In_3706,In_4332);
and U1667 (N_1667,In_4522,In_4211);
nand U1668 (N_1668,In_652,In_902);
nand U1669 (N_1669,In_1088,In_4852);
nor U1670 (N_1670,In_963,In_1212);
nor U1671 (N_1671,In_2081,In_375);
and U1672 (N_1672,In_322,In_3660);
nor U1673 (N_1673,In_2910,In_2446);
nor U1674 (N_1674,In_4661,In_3710);
or U1675 (N_1675,In_1644,In_2198);
xnor U1676 (N_1676,In_3590,In_1929);
xnor U1677 (N_1677,In_690,In_888);
and U1678 (N_1678,In_2379,In_1821);
xor U1679 (N_1679,In_360,In_53);
nand U1680 (N_1680,In_3727,In_1345);
nand U1681 (N_1681,In_4810,In_4324);
or U1682 (N_1682,In_1498,In_3771);
and U1683 (N_1683,In_3487,In_2864);
nand U1684 (N_1684,In_3479,In_1561);
or U1685 (N_1685,In_2434,In_3810);
nand U1686 (N_1686,In_3430,In_3513);
or U1687 (N_1687,In_644,In_3688);
nand U1688 (N_1688,In_4955,In_1732);
xnor U1689 (N_1689,In_2667,In_1770);
xor U1690 (N_1690,In_3869,In_3124);
nor U1691 (N_1691,In_1287,In_3995);
nand U1692 (N_1692,In_294,In_2659);
nand U1693 (N_1693,In_3821,In_2043);
nand U1694 (N_1694,In_1350,In_2345);
xnor U1695 (N_1695,In_3597,In_2454);
or U1696 (N_1696,In_242,In_846);
and U1697 (N_1697,In_1905,In_588);
nor U1698 (N_1698,In_224,In_2421);
and U1699 (N_1699,In_2137,In_3269);
nor U1700 (N_1700,In_3061,In_3518);
nand U1701 (N_1701,In_1800,In_364);
nand U1702 (N_1702,In_4086,In_4638);
xnor U1703 (N_1703,In_4253,In_1012);
nor U1704 (N_1704,In_4269,In_1384);
or U1705 (N_1705,In_3196,In_1340);
nand U1706 (N_1706,In_4181,In_3605);
nor U1707 (N_1707,In_870,In_3843);
xor U1708 (N_1708,In_1748,In_1281);
nor U1709 (N_1709,In_4216,In_2170);
xor U1710 (N_1710,In_4073,In_838);
nor U1711 (N_1711,In_238,In_328);
and U1712 (N_1712,In_3543,In_2653);
xnor U1713 (N_1713,In_3963,In_1132);
and U1714 (N_1714,In_4042,In_199);
nand U1715 (N_1715,In_4405,In_4059);
or U1716 (N_1716,In_4785,In_1019);
and U1717 (N_1717,In_1934,In_3764);
or U1718 (N_1718,In_2079,In_4101);
or U1719 (N_1719,In_3072,In_1875);
or U1720 (N_1720,In_2172,In_1988);
xor U1721 (N_1721,In_3416,In_1822);
xnor U1722 (N_1722,In_3718,In_4349);
nand U1723 (N_1723,In_520,In_1660);
nand U1724 (N_1724,In_2470,In_3027);
xnor U1725 (N_1725,In_4434,In_3253);
nor U1726 (N_1726,In_2841,In_2465);
xor U1727 (N_1727,In_3369,In_3837);
xor U1728 (N_1728,In_3801,In_691);
xor U1729 (N_1729,In_111,In_839);
nand U1730 (N_1730,In_1025,In_1241);
or U1731 (N_1731,In_3528,In_1703);
nor U1732 (N_1732,In_704,In_2004);
nor U1733 (N_1733,In_4401,In_4740);
nand U1734 (N_1734,In_2796,In_2769);
and U1735 (N_1735,In_2797,In_3364);
nor U1736 (N_1736,In_1099,In_804);
or U1737 (N_1737,In_1167,In_4261);
xnor U1738 (N_1738,In_94,In_2393);
or U1739 (N_1739,In_2085,In_287);
nand U1740 (N_1740,In_4856,In_1423);
or U1741 (N_1741,In_4466,In_4423);
nand U1742 (N_1742,In_406,In_17);
nand U1743 (N_1743,In_608,In_4696);
xor U1744 (N_1744,In_4026,In_4315);
or U1745 (N_1745,In_533,In_983);
and U1746 (N_1746,In_470,In_4218);
and U1747 (N_1747,In_2287,In_1645);
and U1748 (N_1748,In_2241,In_3841);
and U1749 (N_1749,In_1889,In_901);
xor U1750 (N_1750,In_818,In_3770);
and U1751 (N_1751,In_1221,In_2042);
nand U1752 (N_1752,In_408,In_1817);
nor U1753 (N_1753,In_1060,In_4629);
nand U1754 (N_1754,In_3306,In_1870);
nor U1755 (N_1755,In_3985,In_401);
and U1756 (N_1756,In_2284,In_2245);
nor U1757 (N_1757,In_153,In_3272);
or U1758 (N_1758,In_842,In_4568);
or U1759 (N_1759,In_3982,In_310);
nor U1760 (N_1760,In_3133,In_2067);
xnor U1761 (N_1761,In_1951,In_3495);
xnor U1762 (N_1762,In_3968,In_1196);
and U1763 (N_1763,In_4847,In_4692);
nand U1764 (N_1764,In_3485,In_1798);
nor U1765 (N_1765,In_3304,In_574);
and U1766 (N_1766,In_1909,In_2184);
and U1767 (N_1767,In_440,In_719);
nand U1768 (N_1768,In_2710,In_1224);
and U1769 (N_1769,In_4899,In_2270);
or U1770 (N_1770,In_4151,In_2407);
or U1771 (N_1771,In_2105,In_2569);
nor U1772 (N_1772,In_3271,In_2660);
xor U1773 (N_1773,In_1446,In_2904);
nor U1774 (N_1774,In_1609,In_3932);
nor U1775 (N_1775,In_2732,In_2009);
and U1776 (N_1776,In_84,In_3142);
xnor U1777 (N_1777,In_4143,In_2565);
or U1778 (N_1778,In_1140,In_4102);
xor U1779 (N_1779,In_841,In_1390);
nand U1780 (N_1780,In_3293,In_3480);
xor U1781 (N_1781,In_192,In_477);
nor U1782 (N_1782,In_510,In_684);
and U1783 (N_1783,In_4366,In_3192);
nor U1784 (N_1784,In_3772,In_3630);
and U1785 (N_1785,In_259,In_1251);
and U1786 (N_1786,In_2116,In_4469);
nand U1787 (N_1787,In_1286,In_2815);
or U1788 (N_1788,In_2498,In_2768);
xnor U1789 (N_1789,In_2306,In_4926);
nand U1790 (N_1790,In_2638,In_2488);
nor U1791 (N_1791,In_4565,In_1612);
xnor U1792 (N_1792,In_19,In_1738);
or U1793 (N_1793,In_2277,In_137);
or U1794 (N_1794,In_579,In_2376);
nand U1795 (N_1795,In_2993,In_482);
nor U1796 (N_1796,In_602,In_890);
and U1797 (N_1797,In_167,In_1006);
nor U1798 (N_1798,In_4900,In_1534);
nand U1799 (N_1799,In_3267,In_2975);
nand U1800 (N_1800,In_2753,In_3109);
xnor U1801 (N_1801,In_3568,In_2072);
xnor U1802 (N_1802,In_3647,In_1814);
xor U1803 (N_1803,In_2745,In_4419);
xor U1804 (N_1804,In_3035,In_206);
and U1805 (N_1805,In_501,In_3998);
nor U1806 (N_1806,In_1239,In_903);
nor U1807 (N_1807,In_2112,In_3340);
nor U1808 (N_1808,In_536,In_426);
or U1809 (N_1809,In_2749,In_2153);
nand U1810 (N_1810,In_28,In_3829);
xor U1811 (N_1811,In_659,In_4503);
or U1812 (N_1812,In_1377,In_2196);
nand U1813 (N_1813,In_129,In_2397);
and U1814 (N_1814,In_2118,In_4933);
nand U1815 (N_1815,In_597,In_1337);
and U1816 (N_1816,In_2613,In_2884);
or U1817 (N_1817,In_2523,In_2150);
xor U1818 (N_1818,In_3711,In_1995);
or U1819 (N_1819,In_1852,In_2409);
and U1820 (N_1820,In_1603,In_295);
nor U1821 (N_1821,In_4608,In_2936);
and U1822 (N_1822,In_733,In_1066);
nand U1823 (N_1823,In_1687,In_2695);
and U1824 (N_1824,In_4510,In_1486);
and U1825 (N_1825,In_4697,In_600);
nand U1826 (N_1826,In_1203,In_4190);
nor U1827 (N_1827,In_2692,In_4371);
and U1828 (N_1828,In_4690,In_274);
or U1829 (N_1829,In_2688,In_815);
nand U1830 (N_1830,In_344,In_319);
xor U1831 (N_1831,In_2685,In_4325);
nand U1832 (N_1832,In_1541,In_3307);
nand U1833 (N_1833,In_1957,In_3639);
nor U1834 (N_1834,In_4027,In_555);
and U1835 (N_1835,In_4278,In_4067);
or U1836 (N_1836,In_2561,In_1587);
nor U1837 (N_1837,In_1749,In_4130);
nand U1838 (N_1838,In_35,In_3254);
or U1839 (N_1839,In_3483,In_2639);
nor U1840 (N_1840,In_1393,In_3346);
and U1841 (N_1841,In_1778,In_4952);
or U1842 (N_1842,In_3085,In_1750);
nand U1843 (N_1843,In_1085,In_3953);
xor U1844 (N_1844,In_3044,In_3503);
xnor U1845 (N_1845,In_3220,In_279);
xor U1846 (N_1846,In_4514,In_1971);
xor U1847 (N_1847,In_1872,In_4975);
or U1848 (N_1848,In_1354,In_1313);
or U1849 (N_1849,In_3168,In_1441);
and U1850 (N_1850,In_1727,In_3921);
nand U1851 (N_1851,In_4213,In_3750);
nor U1852 (N_1852,In_4060,In_228);
xnor U1853 (N_1853,In_1295,In_3402);
nand U1854 (N_1854,In_3042,In_827);
and U1855 (N_1855,In_3126,In_2655);
xnor U1856 (N_1856,In_29,In_4821);
nand U1857 (N_1857,In_848,In_2445);
and U1858 (N_1858,In_3312,In_1632);
nor U1859 (N_1859,In_3164,In_1413);
xnor U1860 (N_1860,In_4486,In_237);
and U1861 (N_1861,In_3301,In_3949);
or U1862 (N_1862,In_1742,In_3474);
nor U1863 (N_1863,In_1598,In_4135);
nand U1864 (N_1864,In_669,In_4377);
or U1865 (N_1865,In_1124,In_2007);
or U1866 (N_1866,In_632,In_2159);
and U1867 (N_1867,In_4988,In_3908);
or U1868 (N_1868,In_3135,In_2543);
and U1869 (N_1869,In_4399,In_712);
and U1870 (N_1870,In_2373,In_1411);
nor U1871 (N_1871,In_4129,In_2186);
and U1872 (N_1872,In_2411,In_3201);
nor U1873 (N_1873,In_157,In_4232);
or U1874 (N_1874,In_3226,In_340);
nand U1875 (N_1875,In_3849,In_1808);
nor U1876 (N_1876,In_1811,In_3222);
nand U1877 (N_1877,In_2790,In_1710);
and U1878 (N_1878,In_537,In_2738);
xnor U1879 (N_1879,In_2313,In_1014);
and U1880 (N_1880,In_4120,In_758);
and U1881 (N_1881,In_1691,In_2541);
nand U1882 (N_1882,In_4989,In_4176);
nor U1883 (N_1883,In_3969,In_2130);
nand U1884 (N_1884,In_2865,In_2909);
nand U1885 (N_1885,In_1047,In_984);
nand U1886 (N_1886,In_543,In_3700);
nand U1887 (N_1887,In_3586,In_3343);
xor U1888 (N_1888,In_2758,In_2014);
xor U1889 (N_1889,In_3152,In_2763);
or U1890 (N_1890,In_1666,In_1137);
and U1891 (N_1891,In_3425,In_3977);
xnor U1892 (N_1892,In_2261,In_4773);
xor U1893 (N_1893,In_3685,In_1310);
nand U1894 (N_1894,In_3247,In_4234);
xor U1895 (N_1895,In_3600,In_4521);
nor U1896 (N_1896,In_3342,In_960);
nand U1897 (N_1897,In_4484,In_4472);
nand U1898 (N_1898,In_2634,In_634);
or U1899 (N_1899,In_269,In_183);
nand U1900 (N_1900,In_613,In_4170);
nor U1901 (N_1901,In_1416,In_4192);
nand U1902 (N_1902,In_4830,In_4994);
or U1903 (N_1903,In_4826,In_3316);
nor U1904 (N_1904,In_4327,In_2762);
nand U1905 (N_1905,In_4240,In_9);
nand U1906 (N_1906,In_853,In_1002);
and U1907 (N_1907,In_1214,In_936);
or U1908 (N_1908,In_3029,In_2689);
nand U1909 (N_1909,In_44,In_2855);
and U1910 (N_1910,In_1518,In_3533);
nor U1911 (N_1911,In_3844,In_1366);
nor U1912 (N_1912,In_4587,In_1696);
nand U1913 (N_1913,In_1101,In_1080);
nor U1914 (N_1914,In_1717,In_4776);
and U1915 (N_1915,In_1526,In_1296);
nor U1916 (N_1916,In_50,In_2791);
and U1917 (N_1917,In_3144,In_1820);
nor U1918 (N_1918,In_738,In_4563);
and U1919 (N_1919,In_3062,In_3554);
xor U1920 (N_1920,In_1919,In_4770);
nand U1921 (N_1921,In_3385,In_4292);
or U1922 (N_1922,In_4669,In_1309);
nor U1923 (N_1923,In_2507,In_3069);
nand U1924 (N_1924,In_332,In_3589);
or U1925 (N_1925,In_745,In_2516);
or U1926 (N_1926,In_203,In_3851);
nand U1927 (N_1927,In_3120,In_1206);
and U1928 (N_1928,In_2034,In_3524);
nand U1929 (N_1929,In_1178,In_2114);
nor U1930 (N_1930,In_1984,In_3410);
or U1931 (N_1931,In_432,In_806);
or U1932 (N_1932,In_3016,In_3266);
and U1933 (N_1933,In_2483,In_211);
xor U1934 (N_1934,In_2719,In_562);
or U1935 (N_1935,In_1369,In_3646);
nor U1936 (N_1936,In_4390,In_2919);
nor U1937 (N_1937,In_1622,In_1181);
xor U1938 (N_1938,In_2002,In_423);
xor U1939 (N_1939,In_2570,In_2447);
nand U1940 (N_1940,In_772,In_4999);
and U1941 (N_1941,In_173,In_372);
nand U1942 (N_1942,In_2960,In_3303);
or U1943 (N_1943,In_816,In_4167);
nand U1944 (N_1944,In_4741,In_2799);
nand U1945 (N_1945,In_4244,In_1292);
nor U1946 (N_1946,In_1068,In_2264);
or U1947 (N_1947,In_1618,In_3715);
nor U1948 (N_1948,In_3317,In_1648);
and U1949 (N_1949,In_181,In_2384);
nor U1950 (N_1950,In_1927,In_2957);
and U1951 (N_1951,In_2493,In_404);
nand U1952 (N_1952,In_3217,In_2709);
nand U1953 (N_1953,In_1270,In_4300);
or U1954 (N_1954,In_4737,In_4624);
or U1955 (N_1955,In_2622,In_1824);
nand U1956 (N_1956,In_1604,In_4664);
and U1957 (N_1957,In_427,In_1761);
and U1958 (N_1958,In_436,In_2526);
nor U1959 (N_1959,In_2616,In_3614);
nor U1960 (N_1960,In_4671,In_2671);
xor U1961 (N_1961,In_2144,In_3339);
and U1962 (N_1962,In_949,In_2362);
xor U1963 (N_1963,In_3030,In_4794);
xnor U1964 (N_1964,In_492,In_1533);
or U1965 (N_1965,In_2074,In_3960);
and U1966 (N_1966,In_4823,In_2490);
and U1967 (N_1967,In_4214,In_1444);
xnor U1968 (N_1968,In_4978,In_3595);
nor U1969 (N_1969,In_4869,In_518);
nor U1970 (N_1970,In_22,In_4879);
or U1971 (N_1971,In_370,In_3782);
and U1972 (N_1972,In_953,In_3153);
nand U1973 (N_1973,In_954,In_109);
nand U1974 (N_1974,In_1838,In_2371);
xnor U1975 (N_1975,In_4256,In_2566);
xor U1976 (N_1976,In_2611,In_2369);
and U1977 (N_1977,In_1225,In_2770);
or U1978 (N_1978,In_3806,In_1274);
nor U1979 (N_1979,In_1272,In_2046);
nand U1980 (N_1980,In_1676,In_2242);
xor U1981 (N_1981,In_3175,In_1787);
nor U1982 (N_1982,In_2201,In_3499);
xor U1983 (N_1983,In_3643,In_1211);
and U1984 (N_1984,In_808,In_1485);
or U1985 (N_1985,In_1335,In_930);
and U1986 (N_1986,In_2050,In_2485);
nor U1987 (N_1987,In_1473,In_3823);
and U1988 (N_1988,In_4432,In_4612);
or U1989 (N_1989,In_775,In_2178);
nand U1990 (N_1990,In_541,In_3427);
xor U1991 (N_1991,In_2266,In_3460);
xnor U1992 (N_1992,In_3657,In_4513);
nor U1993 (N_1993,In_3807,In_226);
or U1994 (N_1994,In_654,In_1530);
nand U1995 (N_1995,In_1730,In_160);
nor U1996 (N_1996,In_87,In_3747);
and U1997 (N_1997,In_1850,In_3729);
nor U1998 (N_1998,In_2418,In_4980);
nand U1999 (N_1999,In_2510,In_3834);
and U2000 (N_2000,In_4150,In_792);
nor U2001 (N_2001,In_2820,In_3493);
or U2002 (N_2002,In_1049,In_598);
and U2003 (N_2003,In_798,In_4123);
nor U2004 (N_2004,In_3261,In_4778);
or U2005 (N_2005,In_3575,In_3875);
nand U2006 (N_2006,In_280,In_4483);
and U2007 (N_2007,In_323,In_4290);
and U2008 (N_2008,In_3583,In_2157);
nand U2009 (N_2009,In_2976,In_3423);
nor U2010 (N_2010,In_4082,In_4873);
and U2011 (N_2011,In_4369,In_1263);
xor U2012 (N_2012,In_3255,In_2662);
nand U2013 (N_2013,In_2937,In_3831);
and U2014 (N_2014,In_2802,In_2182);
nor U2015 (N_2015,In_3574,In_162);
or U2016 (N_2016,In_1234,In_2318);
or U2017 (N_2017,In_604,In_3234);
nor U2018 (N_2018,In_4471,In_858);
and U2019 (N_2019,In_4647,In_3353);
and U2020 (N_2020,In_558,In_1361);
and U2021 (N_2021,In_730,In_2148);
nor U2022 (N_2022,In_2030,In_2893);
nand U2023 (N_2023,In_2426,In_464);
nand U2024 (N_2024,In_4584,In_2267);
and U2025 (N_2025,In_1040,In_1353);
xor U2026 (N_2026,In_4950,In_761);
nor U2027 (N_2027,In_2704,In_1535);
xor U2028 (N_2028,In_1357,In_523);
or U2029 (N_2029,In_114,In_4422);
xnor U2030 (N_2030,In_2375,In_3023);
xor U2031 (N_2031,In_1215,In_2352);
and U2032 (N_2032,In_2715,In_2649);
nor U2033 (N_2033,In_3320,In_2905);
nor U2034 (N_2034,In_2751,In_1406);
or U2035 (N_2035,In_633,In_2008);
and U2036 (N_2036,In_1378,In_2856);
and U2037 (N_2037,In_4532,In_1302);
xor U2038 (N_2038,In_4168,In_2396);
and U2039 (N_2039,In_1217,In_596);
or U2040 (N_2040,In_4507,In_3799);
or U2041 (N_2041,In_4501,In_4331);
and U2042 (N_2042,In_3033,In_2083);
or U2043 (N_2043,In_4085,In_40);
nor U2044 (N_2044,In_1601,In_4090);
and U2045 (N_2045,In_4196,In_1560);
xor U2046 (N_2046,In_3531,In_3577);
nor U2047 (N_2047,In_757,In_2331);
and U2048 (N_2048,In_3730,In_257);
or U2049 (N_2049,In_4882,In_452);
nand U2050 (N_2050,In_529,In_3158);
xor U2051 (N_2051,In_155,In_1860);
xor U2052 (N_2052,In_4701,In_2949);
nand U2053 (N_2053,In_4905,In_1855);
and U2054 (N_2054,In_1396,In_2511);
and U2055 (N_2055,In_3945,In_3300);
or U2056 (N_2056,In_1910,In_256);
nand U2057 (N_2057,In_2810,In_1701);
nor U2058 (N_2058,In_248,In_2603);
xor U2059 (N_2059,In_4065,In_3790);
and U2060 (N_2060,In_2056,In_24);
nand U2061 (N_2061,In_3593,In_4287);
nor U2062 (N_2062,In_4498,In_3418);
nor U2063 (N_2063,In_3389,In_1623);
and U2064 (N_2064,In_1191,In_1550);
and U2065 (N_2065,In_2956,In_3576);
or U2066 (N_2066,In_2183,In_1460);
nor U2067 (N_2067,In_3690,In_1651);
or U2068 (N_2068,In_695,In_2771);
or U2069 (N_2069,In_77,In_924);
nor U2070 (N_2070,In_3802,In_468);
nand U2071 (N_2071,In_4071,In_1913);
xor U2072 (N_2072,In_2210,In_2513);
nand U2073 (N_2073,In_2911,In_2822);
xnor U2074 (N_2074,In_3954,In_1056);
nand U2075 (N_2075,In_4677,In_1125);
nand U2076 (N_2076,In_2723,In_71);
nand U2077 (N_2077,In_2974,In_3360);
nor U2078 (N_2078,In_927,In_3187);
nand U2079 (N_2079,In_1653,In_1699);
nand U2080 (N_2080,In_1629,In_1024);
and U2081 (N_2081,In_641,In_2442);
nor U2082 (N_2082,In_3034,In_2236);
or U2083 (N_2083,In_1706,In_1746);
or U2084 (N_2084,In_1481,In_455);
and U2085 (N_2085,In_472,In_2952);
nor U2086 (N_2086,In_4343,In_2609);
or U2087 (N_2087,In_4594,In_3302);
nand U2088 (N_2088,In_1100,In_4805);
xnor U2089 (N_2089,In_3310,In_1306);
nand U2090 (N_2090,In_620,In_3936);
or U2091 (N_2091,In_3947,In_4066);
and U2092 (N_2092,In_3803,In_4166);
and U2093 (N_2093,In_4611,In_1193);
nand U2094 (N_2094,In_2906,In_823);
and U2095 (N_2095,In_1678,In_1955);
nor U2096 (N_2096,In_3697,In_3004);
xor U2097 (N_2097,In_2728,In_4427);
xnor U2098 (N_2098,In_3582,In_4032);
and U2099 (N_2099,In_2057,In_2678);
and U2100 (N_2100,In_2714,In_2064);
and U2101 (N_2101,In_1256,In_3746);
nand U2102 (N_2102,In_4651,In_865);
nor U2103 (N_2103,In_3112,In_589);
nand U2104 (N_2104,In_4099,In_2107);
nor U2105 (N_2105,In_1806,In_1755);
or U2106 (N_2106,In_2962,In_1723);
nand U2107 (N_2107,In_4468,In_1990);
or U2108 (N_2108,In_3758,In_3682);
nor U2109 (N_2109,In_1972,In_3632);
nand U2110 (N_2110,In_4033,In_3507);
xor U2111 (N_2111,In_3787,In_480);
xnor U2112 (N_2112,In_3043,In_857);
nor U2113 (N_2113,In_4917,In_3383);
and U2114 (N_2114,In_3603,In_481);
and U2115 (N_2115,In_2847,In_1998);
and U2116 (N_2116,In_354,In_3134);
nand U2117 (N_2117,In_1677,In_402);
or U2118 (N_2118,In_2573,In_891);
xnor U2119 (N_2119,In_1119,In_1834);
and U2120 (N_2120,In_3019,In_2061);
xnor U2121 (N_2121,In_154,In_3958);
nand U2122 (N_2122,In_1922,In_2881);
nor U2123 (N_2123,In_2052,In_403);
xnor U2124 (N_2124,In_136,In_398);
xor U2125 (N_2125,In_931,In_4268);
or U2126 (N_2126,In_1367,In_1846);
or U2127 (N_2127,In_45,In_2832);
nand U2128 (N_2128,In_219,In_496);
nor U2129 (N_2129,In_3828,In_216);
and U2130 (N_2130,In_3488,In_4644);
xnor U2131 (N_2131,In_3370,In_2134);
xnor U2132 (N_2132,In_2640,In_2231);
nor U2133 (N_2133,In_2528,In_1436);
nand U2134 (N_2134,In_4363,In_3186);
and U2135 (N_2135,In_2387,In_2844);
nor U2136 (N_2136,In_2997,In_2291);
nor U2137 (N_2137,In_4207,In_845);
xor U2138 (N_2138,In_1180,In_1095);
nor U2139 (N_2139,In_2026,In_4572);
nor U2140 (N_2140,In_2863,In_467);
xor U2141 (N_2141,In_1035,In_4652);
or U2142 (N_2142,In_3363,In_2179);
nor U2143 (N_2143,In_2779,In_4441);
nand U2144 (N_2144,In_4445,In_3626);
or U2145 (N_2145,In_578,In_3174);
nand U2146 (N_2146,In_1565,In_4004);
or U2147 (N_2147,In_4667,In_1566);
nand U2148 (N_2148,In_4391,In_4788);
or U2149 (N_2149,In_1559,In_3753);
xor U2150 (N_2150,In_3930,In_3521);
nand U2151 (N_2151,In_407,In_886);
or U2152 (N_2152,In_4257,In_1067);
nor U2153 (N_2153,In_2944,In_583);
xor U2154 (N_2154,In_2761,In_4903);
or U2155 (N_2155,In_133,In_2197);
xnor U2156 (N_2156,In_4603,In_1516);
xor U2157 (N_2157,In_2777,In_4128);
nor U2158 (N_2158,In_2593,In_1945);
nand U2159 (N_2159,In_4731,In_2628);
xnor U2160 (N_2160,In_1113,In_4161);
and U2161 (N_2161,In_494,In_4337);
xnor U2162 (N_2162,In_2861,In_4543);
xor U2163 (N_2163,In_762,In_4609);
nor U2164 (N_2164,In_4720,In_1786);
or U2165 (N_2165,In_1639,In_834);
nor U2166 (N_2166,In_986,In_4861);
nor U2167 (N_2167,In_3548,In_2955);
nand U2168 (N_2168,In_567,In_3240);
and U2169 (N_2169,In_1259,In_2874);
nor U2170 (N_2170,In_201,In_611);
and U2171 (N_2171,In_832,In_3638);
xnor U2172 (N_2172,In_4682,In_324);
or U2173 (N_2173,In_302,In_4382);
nand U2174 (N_2174,In_513,In_3396);
or U2175 (N_2175,In_4088,In_4710);
and U2176 (N_2176,In_2297,In_152);
nor U2177 (N_2177,In_693,In_110);
and U2178 (N_2178,In_4836,In_198);
nand U2179 (N_2179,In_1172,In_3663);
xnor U2180 (N_2180,In_141,In_2548);
nor U2181 (N_2181,In_787,In_2257);
and U2182 (N_2182,In_117,In_2806);
nand U2183 (N_2183,In_4283,In_2415);
and U2184 (N_2184,In_4519,In_1414);
or U2185 (N_2185,In_884,In_270);
or U2186 (N_2186,In_1404,In_4506);
nand U2187 (N_2187,In_4276,In_1462);
and U2188 (N_2188,In_569,In_33);
nor U2189 (N_2189,In_3208,In_4817);
nor U2190 (N_2190,In_4775,In_2095);
nor U2191 (N_2191,In_1568,In_463);
or U2192 (N_2192,In_3305,In_1647);
or U2193 (N_2193,In_158,In_283);
nor U2194 (N_2194,In_1288,In_3205);
or U2195 (N_2195,In_1160,In_1289);
or U2196 (N_2196,In_338,In_4319);
nand U2197 (N_2197,In_645,In_2629);
and U2198 (N_2198,In_1836,In_1447);
nor U2199 (N_2199,In_380,In_739);
xnor U2200 (N_2200,In_3398,In_388);
or U2201 (N_2201,In_4388,In_2862);
nand U2202 (N_2202,In_618,In_2965);
xor U2203 (N_2203,In_4462,In_2211);
nand U2204 (N_2204,In_4806,In_828);
or U2205 (N_2205,In_2036,In_3625);
and U2206 (N_2206,In_3290,In_2419);
nor U2207 (N_2207,In_1549,In_1450);
or U2208 (N_2208,In_3213,In_1017);
nor U2209 (N_2209,In_1083,In_1801);
nor U2210 (N_2210,In_3809,In_4837);
xnor U2211 (N_2211,In_701,In_4691);
nor U2212 (N_2212,In_3197,In_4402);
or U2213 (N_2213,In_1030,In_4265);
nor U2214 (N_2214,In_3978,In_3047);
or U2215 (N_2215,In_4322,In_4779);
nand U2216 (N_2216,In_982,In_2377);
xnor U2217 (N_2217,In_491,In_4913);
and U2218 (N_2218,In_4404,In_3211);
or U2219 (N_2219,In_416,In_1845);
or U2220 (N_2220,In_2335,In_3080);
nor U2221 (N_2221,In_4103,In_2273);
nand U2222 (N_2222,In_1667,In_1615);
nor U2223 (N_2223,In_568,In_3173);
and U2224 (N_2224,In_1573,In_330);
and U2225 (N_2225,In_2720,In_2410);
nand U2226 (N_2226,In_4485,In_4318);
or U2227 (N_2227,In_1646,In_3008);
or U2228 (N_2228,In_299,In_4158);
or U2229 (N_2229,In_465,In_3156);
nor U2230 (N_2230,In_2731,In_530);
nor U2231 (N_2231,In_2111,In_3956);
xnor U2232 (N_2232,In_4621,In_3294);
nor U2233 (N_2233,In_592,In_1144);
xor U2234 (N_2234,In_1057,In_1725);
xor U2235 (N_2235,In_1591,In_147);
nor U2236 (N_2236,In_442,In_2740);
xnor U2237 (N_2237,In_1959,In_1620);
nand U2238 (N_2238,In_3779,In_4843);
nor U2239 (N_2239,In_3469,In_3239);
xnor U2240 (N_2240,In_3658,In_389);
nand U2241 (N_2241,In_551,In_4157);
and U2242 (N_2242,In_449,In_2020);
or U2243 (N_2243,In_59,In_2326);
and U2244 (N_2244,In_3871,In_672);
nor U2245 (N_2245,In_2163,In_1823);
and U2246 (N_2246,In_4236,In_144);
xor U2247 (N_2247,In_3236,In_356);
and U2248 (N_2248,In_988,In_904);
xor U2249 (N_2249,In_992,In_866);
nor U2250 (N_2250,In_2664,In_305);
and U2251 (N_2251,In_4182,In_3581);
nand U2252 (N_2252,In_4743,In_746);
or U2253 (N_2253,In_799,In_3633);
nor U2254 (N_2254,In_4759,In_2915);
nor U2255 (N_2255,In_1314,In_3358);
nor U2256 (N_2256,In_2188,In_3763);
nand U2257 (N_2257,In_81,In_4081);
nand U2258 (N_2258,In_1150,In_3813);
nand U2259 (N_2259,In_4002,In_2222);
xor U2260 (N_2260,In_2063,In_714);
or U2261 (N_2261,In_3476,In_860);
or U2262 (N_2262,In_3720,In_1043);
nand U2263 (N_2263,In_4095,In_1828);
and U2264 (N_2264,In_805,In_2003);
nor U2265 (N_2265,In_100,In_2340);
nand U2266 (N_2266,In_1735,In_1899);
or U2267 (N_2267,In_4875,In_331);
nand U2268 (N_2268,In_3184,In_2174);
nand U2269 (N_2269,In_2314,In_2484);
or U2270 (N_2270,In_2147,In_1818);
nand U2271 (N_2271,In_3297,In_2702);
nand U2272 (N_2272,In_3914,In_4589);
xor U2273 (N_2273,In_560,In_1233);
nand U2274 (N_2274,In_4397,In_2438);
nor U2275 (N_2275,In_3218,In_2813);
and U2276 (N_2276,In_4270,In_3678);
xor U2277 (N_2277,In_1757,In_3172);
or U2278 (N_2278,In_1189,In_1802);
and U2279 (N_2279,In_3464,In_4303);
or U2280 (N_2280,In_268,In_4173);
or U2281 (N_2281,In_414,In_132);
xor U2282 (N_2282,In_306,In_2250);
xnor U2283 (N_2283,In_1853,In_3569);
nand U2284 (N_2284,In_1674,In_2333);
nor U2285 (N_2285,In_3404,In_2341);
nand U2286 (N_2286,In_3825,In_1415);
nor U2287 (N_2287,In_74,In_3227);
xor U2288 (N_2288,In_3338,In_2831);
xor U2289 (N_2289,In_1513,In_2082);
nand U2290 (N_2290,In_3863,In_2699);
nand U2291 (N_2291,In_868,In_1235);
xor U2292 (N_2292,In_13,In_4694);
xnor U2293 (N_2293,In_1960,In_2343);
xor U2294 (N_2294,In_4100,In_4517);
nand U2295 (N_2295,In_2833,In_2049);
and U2296 (N_2296,In_4932,In_170);
xnor U2297 (N_2297,In_1076,In_3959);
nor U2298 (N_2298,In_4700,In_1102);
xor U2299 (N_2299,In_3796,In_3057);
nor U2300 (N_2300,In_3862,In_382);
xor U2301 (N_2301,In_64,In_314);
or U2302 (N_2302,In_1463,In_987);
and U2303 (N_2303,In_484,In_27);
nor U2304 (N_2304,In_2620,In_2696);
and U2305 (N_2305,In_3708,In_2585);
xnor U2306 (N_2306,In_3944,In_3413);
xnor U2307 (N_2307,In_774,In_707);
or U2308 (N_2308,In_3066,In_2567);
or U2309 (N_2309,In_4586,In_3673);
or U2310 (N_2310,In_2712,In_4648);
nor U2311 (N_2311,In_3879,In_4977);
nand U2312 (N_2312,In_3449,In_1596);
and U2313 (N_2313,In_1490,In_2584);
nor U2314 (N_2314,In_1713,In_3933);
nor U2315 (N_2315,In_311,In_1176);
nor U2316 (N_2316,In_2933,In_4693);
or U2317 (N_2317,In_996,In_850);
xor U2318 (N_2318,In_1365,In_3078);
nand U2319 (N_2319,In_3532,In_486);
nand U2320 (N_2320,In_3406,In_586);
xnor U2321 (N_2321,In_3250,In_1540);
xnor U2322 (N_2322,In_4124,In_4516);
or U2323 (N_2323,In_4262,In_3549);
xor U2324 (N_2324,In_1138,In_3291);
xnor U2325 (N_2325,In_4554,In_2017);
xor U2326 (N_2326,In_103,In_4428);
nand U2327 (N_2327,In_1769,In_716);
and U2328 (N_2328,In_4641,In_4392);
xnor U2329 (N_2329,In_4646,In_4365);
or U2330 (N_2330,In_4702,In_4556);
or U2331 (N_2331,In_1208,In_3784);
and U2332 (N_2332,In_3557,In_150);
nand U2333 (N_2333,In_1011,In_4972);
nor U2334 (N_2334,In_3477,In_2460);
and U2335 (N_2335,In_1220,In_2290);
and U2336 (N_2336,In_4831,In_1906);
and U2337 (N_2337,In_139,In_4748);
nor U2338 (N_2338,In_1465,In_3037);
or U2339 (N_2339,In_871,In_4728);
or U2340 (N_2340,In_1112,In_1161);
or U2341 (N_2341,In_4015,In_4985);
or U2342 (N_2342,In_1145,In_2760);
or U2343 (N_2343,In_748,In_2228);
and U2344 (N_2344,In_1155,In_2606);
and U2345 (N_2345,In_1912,In_2945);
nand U2346 (N_2346,In_3668,In_4965);
nand U2347 (N_2347,In_1766,In_65);
and U2348 (N_2348,In_3704,In_3887);
or U2349 (N_2349,In_1979,In_3833);
or U2350 (N_2350,In_2463,In_1857);
or U2351 (N_2351,In_2840,In_4502);
nor U2352 (N_2352,In_1065,In_3766);
nand U2353 (N_2353,In_2309,In_3653);
and U2354 (N_2354,In_4144,In_1474);
or U2355 (N_2355,In_873,In_2787);
nor U2356 (N_2356,In_2496,In_1332);
or U2357 (N_2357,In_2519,In_1608);
nor U2358 (N_2358,In_138,In_3814);
nand U2359 (N_2359,In_450,In_341);
xnor U2360 (N_2360,In_1277,In_4944);
nor U2361 (N_2361,In_3299,In_4716);
nand U2362 (N_2362,In_4277,In_2391);
and U2363 (N_2363,In_4447,In_4137);
or U2364 (N_2364,In_3314,In_3714);
and U2365 (N_2365,In_766,In_254);
nand U2366 (N_2366,In_1576,In_3089);
and U2367 (N_2367,In_411,In_3462);
nor U2368 (N_2368,In_599,In_3165);
and U2369 (N_2369,In_2497,In_3166);
and U2370 (N_2370,In_4113,In_2001);
xnor U2371 (N_2371,In_2798,In_1722);
nand U2372 (N_2372,In_2131,In_1662);
and U2373 (N_2373,In_4596,In_2169);
xor U2374 (N_2374,In_4087,In_2310);
and U2375 (N_2375,In_2743,In_2803);
nand U2376 (N_2376,In_1702,In_4601);
nand U2377 (N_2377,In_2966,In_2793);
nand U2378 (N_2378,In_4230,In_2550);
and U2379 (N_2379,In_2025,In_1294);
or U2380 (N_2380,In_2568,In_2005);
or U2381 (N_2381,In_3847,In_4003);
and U2382 (N_2382,In_4121,In_3392);
xnor U2383 (N_2383,In_363,In_1118);
nor U2384 (N_2384,In_4961,In_488);
and U2385 (N_2385,In_3523,In_3356);
nand U2386 (N_2386,In_786,In_2000);
and U2387 (N_2387,In_563,In_1684);
or U2388 (N_2388,In_4210,In_2757);
xor U2389 (N_2389,In_811,In_4666);
xor U2390 (N_2390,In_3334,In_881);
or U2391 (N_2391,In_3785,In_4438);
nand U2392 (N_2392,In_4983,In_1829);
and U2393 (N_2393,In_944,In_1086);
nand U2394 (N_2394,In_4729,In_2028);
nand U2395 (N_2395,In_3836,In_1557);
nand U2396 (N_2396,In_4650,In_296);
xor U2397 (N_2397,In_190,In_909);
nand U2398 (N_2398,In_200,In_534);
and U2399 (N_2399,In_2828,In_1958);
xor U2400 (N_2400,In_3818,In_2253);
xnor U2401 (N_2401,In_4529,In_2039);
and U2402 (N_2402,In_86,In_2103);
and U2403 (N_2403,In_3681,In_4657);
or U2404 (N_2404,In_2140,In_2124);
and U2405 (N_2405,In_1916,In_1341);
nand U2406 (N_2406,In_4433,In_3692);
and U2407 (N_2407,In_4966,In_2930);
nor U2408 (N_2408,In_2953,In_4313);
nand U2409 (N_2409,In_2631,In_456);
nand U2410 (N_2410,In_4284,In_679);
nor U2411 (N_2411,In_4336,In_2602);
and U2412 (N_2412,In_2303,In_2913);
nand U2413 (N_2413,In_4238,In_648);
or U2414 (N_2414,In_4537,In_1037);
xnor U2415 (N_2415,In_3612,In_367);
nand U2416 (N_2416,In_3331,In_4249);
nand U2417 (N_2417,In_697,In_1064);
xor U2418 (N_2418,In_993,In_358);
nor U2419 (N_2419,In_4145,In_1657);
or U2420 (N_2420,In_703,In_1175);
and U2421 (N_2421,In_4304,In_783);
xor U2422 (N_2422,In_3298,In_142);
and U2423 (N_2423,In_1616,In_159);
or U2424 (N_2424,In_4339,In_2594);
nand U2425 (N_2425,In_985,In_3330);
xor U2426 (N_2426,In_4538,In_345);
and U2427 (N_2427,In_4450,In_869);
xor U2428 (N_2428,In_605,In_660);
or U2429 (N_2429,In_561,In_3139);
nor U2430 (N_2430,In_4034,In_66);
and U2431 (N_2431,In_4013,In_4229);
and U2432 (N_2432,In_1358,In_3976);
nor U2433 (N_2433,In_3074,In_3199);
nor U2434 (N_2434,In_4791,In_2981);
xor U2435 (N_2435,In_655,In_4286);
or U2436 (N_2436,In_4804,In_4892);
and U2437 (N_2437,In_4108,In_1812);
and U2438 (N_2438,In_4186,In_3662);
or U2439 (N_2439,In_1075,In_3015);
xnor U2440 (N_2440,In_4581,In_1136);
xnor U2441 (N_2441,In_1689,In_2449);
or U2442 (N_2442,In_343,In_2041);
nor U2443 (N_2443,In_4786,In_2536);
nor U2444 (N_2444,In_549,In_1531);
xor U2445 (N_2445,In_3102,In_515);
xor U2446 (N_2446,In_125,In_2873);
nor U2447 (N_2447,In_1437,In_2574);
and U2448 (N_2448,In_699,In_2578);
or U2449 (N_2449,In_2907,In_2870);
nand U2450 (N_2450,In_4632,In_3292);
nor U2451 (N_2451,In_4934,In_3489);
and U2452 (N_2452,In_2263,In_260);
xor U2453 (N_2453,In_4957,In_3108);
or U2454 (N_2454,In_2789,In_3816);
nor U2455 (N_2455,In_266,In_3740);
and U2456 (N_2456,In_1726,In_3602);
nor U2457 (N_2457,In_1429,In_1009);
nand U2458 (N_2458,In_261,In_4006);
nor U2459 (N_2459,In_1092,In_1433);
or U2460 (N_2460,In_188,In_2104);
or U2461 (N_2461,In_2736,In_3200);
or U2462 (N_2462,In_4208,In_2413);
or U2463 (N_2463,In_1258,In_1322);
and U2464 (N_2464,In_1525,In_4559);
or U2465 (N_2465,In_1476,In_2325);
nand U2466 (N_2466,In_2801,In_4239);
or U2467 (N_2467,In_1580,In_4381);
or U2468 (N_2468,In_3482,In_2527);
nand U2469 (N_2469,In_3957,In_3867);
and U2470 (N_2470,In_4813,In_720);
xor U2471 (N_2471,In_2476,In_4511);
and U2472 (N_2472,In_4998,In_3231);
nand U2473 (N_2473,In_1170,In_708);
xnor U2474 (N_2474,In_1467,In_4500);
or U2475 (N_2475,In_4426,In_3068);
xor U2476 (N_2476,In_3100,In_4599);
and U2477 (N_2477,In_2983,In_1840);
and U2478 (N_2478,In_1895,In_2872);
nor U2479 (N_2479,In_1740,In_2176);
or U2480 (N_2480,In_4619,In_1081);
nand U2481 (N_2481,In_3721,In_2400);
or U2482 (N_2482,In_2243,In_214);
and U2483 (N_2483,In_812,In_653);
or U2484 (N_2484,In_252,In_3081);
and U2485 (N_2485,In_3838,In_4334);
or U2486 (N_2486,In_4607,In_863);
and U2487 (N_2487,In_4906,In_2765);
or U2488 (N_2488,In_2866,In_4136);
and U2489 (N_2489,In_315,In_368);
or U2490 (N_2490,In_1200,In_3559);
nor U2491 (N_2491,In_856,In_3855);
nor U2492 (N_2492,In_1461,In_3013);
or U2493 (N_2493,In_2398,In_2943);
xnor U2494 (N_2494,In_576,In_434);
and U2495 (N_2495,In_499,In_1816);
and U2496 (N_2496,In_4567,In_4850);
nand U2497 (N_2497,In_1352,In_1408);
nor U2498 (N_2498,In_497,In_1784);
nand U2499 (N_2499,In_2599,In_4885);
or U2500 (N_2500,In_3925,In_4092);
nand U2501 (N_2501,In_4134,In_2841);
nand U2502 (N_2502,In_3824,In_4368);
nand U2503 (N_2503,In_3980,In_3000);
xor U2504 (N_2504,In_902,In_3573);
and U2505 (N_2505,In_2637,In_567);
nand U2506 (N_2506,In_2740,In_2778);
or U2507 (N_2507,In_4540,In_3247);
nand U2508 (N_2508,In_248,In_2462);
and U2509 (N_2509,In_820,In_1478);
nand U2510 (N_2510,In_4486,In_4201);
xor U2511 (N_2511,In_3899,In_2990);
and U2512 (N_2512,In_3414,In_1193);
nor U2513 (N_2513,In_2866,In_156);
and U2514 (N_2514,In_2644,In_3527);
and U2515 (N_2515,In_4875,In_4506);
nand U2516 (N_2516,In_1025,In_273);
xor U2517 (N_2517,In_477,In_970);
nand U2518 (N_2518,In_3501,In_1388);
and U2519 (N_2519,In_986,In_2264);
or U2520 (N_2520,In_264,In_1429);
xnor U2521 (N_2521,In_4740,In_3929);
nor U2522 (N_2522,In_2352,In_4577);
nor U2523 (N_2523,In_225,In_356);
nand U2524 (N_2524,In_2753,In_3382);
or U2525 (N_2525,In_4365,In_958);
and U2526 (N_2526,In_3075,In_2922);
nor U2527 (N_2527,In_2715,In_4620);
nand U2528 (N_2528,In_140,In_3967);
xnor U2529 (N_2529,In_3484,In_2036);
xnor U2530 (N_2530,In_4317,In_1032);
and U2531 (N_2531,In_4462,In_2746);
xor U2532 (N_2532,In_4506,In_1879);
nand U2533 (N_2533,In_4783,In_1009);
and U2534 (N_2534,In_4030,In_639);
and U2535 (N_2535,In_969,In_1307);
nand U2536 (N_2536,In_4768,In_2391);
and U2537 (N_2537,In_2902,In_2491);
xnor U2538 (N_2538,In_699,In_619);
nand U2539 (N_2539,In_3493,In_3151);
or U2540 (N_2540,In_2712,In_1542);
or U2541 (N_2541,In_351,In_3920);
xor U2542 (N_2542,In_437,In_4013);
nand U2543 (N_2543,In_672,In_886);
or U2544 (N_2544,In_3378,In_3801);
nand U2545 (N_2545,In_951,In_1565);
nor U2546 (N_2546,In_2508,In_3674);
or U2547 (N_2547,In_4537,In_4244);
nand U2548 (N_2548,In_2618,In_2680);
nor U2549 (N_2549,In_98,In_722);
nand U2550 (N_2550,In_2732,In_4800);
xnor U2551 (N_2551,In_4334,In_2552);
and U2552 (N_2552,In_3388,In_4973);
or U2553 (N_2553,In_2102,In_333);
or U2554 (N_2554,In_3927,In_2132);
xnor U2555 (N_2555,In_435,In_2155);
nor U2556 (N_2556,In_1524,In_4003);
xnor U2557 (N_2557,In_516,In_3897);
nor U2558 (N_2558,In_3222,In_3803);
xnor U2559 (N_2559,In_1312,In_3738);
nand U2560 (N_2560,In_543,In_2004);
or U2561 (N_2561,In_774,In_686);
nor U2562 (N_2562,In_3067,In_2472);
nand U2563 (N_2563,In_1098,In_4851);
nor U2564 (N_2564,In_1862,In_536);
and U2565 (N_2565,In_2274,In_2421);
xor U2566 (N_2566,In_4017,In_663);
nand U2567 (N_2567,In_2507,In_867);
or U2568 (N_2568,In_3349,In_3671);
and U2569 (N_2569,In_3485,In_4056);
xnor U2570 (N_2570,In_1924,In_1840);
nor U2571 (N_2571,In_182,In_2425);
nand U2572 (N_2572,In_1703,In_650);
xor U2573 (N_2573,In_1210,In_2611);
or U2574 (N_2574,In_4313,In_2473);
xnor U2575 (N_2575,In_3360,In_4785);
and U2576 (N_2576,In_455,In_658);
xnor U2577 (N_2577,In_3713,In_2433);
nor U2578 (N_2578,In_1021,In_3364);
and U2579 (N_2579,In_2689,In_741);
and U2580 (N_2580,In_3858,In_704);
or U2581 (N_2581,In_2521,In_1681);
nor U2582 (N_2582,In_4443,In_31);
nand U2583 (N_2583,In_574,In_4827);
xor U2584 (N_2584,In_2746,In_2658);
and U2585 (N_2585,In_4647,In_525);
and U2586 (N_2586,In_432,In_2114);
and U2587 (N_2587,In_4496,In_491);
or U2588 (N_2588,In_2907,In_167);
nor U2589 (N_2589,In_53,In_453);
nor U2590 (N_2590,In_4356,In_2114);
and U2591 (N_2591,In_2752,In_2050);
or U2592 (N_2592,In_2129,In_4826);
xnor U2593 (N_2593,In_2379,In_3033);
nor U2594 (N_2594,In_1353,In_4120);
xor U2595 (N_2595,In_3594,In_2916);
or U2596 (N_2596,In_2889,In_3131);
nor U2597 (N_2597,In_3941,In_2890);
nor U2598 (N_2598,In_42,In_784);
and U2599 (N_2599,In_4271,In_2776);
nor U2600 (N_2600,In_4484,In_1249);
or U2601 (N_2601,In_2251,In_3891);
nor U2602 (N_2602,In_4063,In_2886);
nor U2603 (N_2603,In_4216,In_4149);
nor U2604 (N_2604,In_1245,In_1174);
or U2605 (N_2605,In_2858,In_3025);
xnor U2606 (N_2606,In_4590,In_3232);
xor U2607 (N_2607,In_3926,In_519);
nand U2608 (N_2608,In_4549,In_1446);
and U2609 (N_2609,In_3479,In_2443);
nor U2610 (N_2610,In_4014,In_3868);
and U2611 (N_2611,In_3864,In_2257);
and U2612 (N_2612,In_2823,In_2592);
nor U2613 (N_2613,In_72,In_979);
and U2614 (N_2614,In_960,In_1576);
nand U2615 (N_2615,In_671,In_884);
nand U2616 (N_2616,In_4553,In_4018);
nand U2617 (N_2617,In_2210,In_57);
and U2618 (N_2618,In_4558,In_760);
and U2619 (N_2619,In_4096,In_3328);
and U2620 (N_2620,In_1613,In_114);
nor U2621 (N_2621,In_3749,In_551);
nor U2622 (N_2622,In_893,In_3297);
or U2623 (N_2623,In_2405,In_4716);
and U2624 (N_2624,In_88,In_284);
nor U2625 (N_2625,In_4693,In_3202);
nand U2626 (N_2626,In_308,In_3696);
nor U2627 (N_2627,In_644,In_4821);
nor U2628 (N_2628,In_3836,In_996);
xor U2629 (N_2629,In_3568,In_4296);
and U2630 (N_2630,In_1256,In_1635);
nor U2631 (N_2631,In_2311,In_2226);
and U2632 (N_2632,In_203,In_4664);
nand U2633 (N_2633,In_2982,In_2918);
and U2634 (N_2634,In_1241,In_3414);
and U2635 (N_2635,In_3720,In_4570);
and U2636 (N_2636,In_4402,In_2517);
nand U2637 (N_2637,In_4831,In_4995);
and U2638 (N_2638,In_4268,In_4871);
and U2639 (N_2639,In_3390,In_2317);
xor U2640 (N_2640,In_4959,In_3992);
xor U2641 (N_2641,In_2487,In_4942);
nor U2642 (N_2642,In_2375,In_1255);
nor U2643 (N_2643,In_3373,In_461);
nor U2644 (N_2644,In_2993,In_3896);
xor U2645 (N_2645,In_827,In_3096);
xor U2646 (N_2646,In_435,In_4751);
nand U2647 (N_2647,In_3185,In_2919);
nand U2648 (N_2648,In_2902,In_916);
xnor U2649 (N_2649,In_1228,In_3220);
xnor U2650 (N_2650,In_761,In_2987);
and U2651 (N_2651,In_1311,In_2420);
or U2652 (N_2652,In_947,In_1173);
nand U2653 (N_2653,In_418,In_1056);
nand U2654 (N_2654,In_3446,In_1363);
xor U2655 (N_2655,In_1521,In_2362);
and U2656 (N_2656,In_259,In_2383);
nor U2657 (N_2657,In_3002,In_1444);
nor U2658 (N_2658,In_2414,In_2872);
and U2659 (N_2659,In_2200,In_269);
xnor U2660 (N_2660,In_4422,In_2587);
or U2661 (N_2661,In_623,In_3661);
xor U2662 (N_2662,In_82,In_1928);
xnor U2663 (N_2663,In_551,In_3938);
nor U2664 (N_2664,In_2341,In_3147);
nor U2665 (N_2665,In_2265,In_193);
xnor U2666 (N_2666,In_4120,In_115);
nand U2667 (N_2667,In_3212,In_1304);
xnor U2668 (N_2668,In_1643,In_866);
nand U2669 (N_2669,In_1066,In_4892);
and U2670 (N_2670,In_1670,In_4377);
nand U2671 (N_2671,In_195,In_3727);
nor U2672 (N_2672,In_3641,In_1);
nor U2673 (N_2673,In_3603,In_1535);
nand U2674 (N_2674,In_32,In_4273);
or U2675 (N_2675,In_2262,In_4272);
or U2676 (N_2676,In_657,In_4202);
xnor U2677 (N_2677,In_2261,In_1354);
and U2678 (N_2678,In_2286,In_642);
nand U2679 (N_2679,In_1488,In_720);
nand U2680 (N_2680,In_3235,In_17);
xor U2681 (N_2681,In_3074,In_3753);
xor U2682 (N_2682,In_3537,In_934);
and U2683 (N_2683,In_14,In_2752);
nor U2684 (N_2684,In_2325,In_4294);
or U2685 (N_2685,In_0,In_17);
or U2686 (N_2686,In_1122,In_3172);
and U2687 (N_2687,In_1811,In_2794);
nand U2688 (N_2688,In_3150,In_130);
nand U2689 (N_2689,In_4896,In_1124);
xor U2690 (N_2690,In_2690,In_1400);
nand U2691 (N_2691,In_670,In_2298);
nor U2692 (N_2692,In_3605,In_3981);
and U2693 (N_2693,In_1440,In_4548);
or U2694 (N_2694,In_4124,In_3235);
nand U2695 (N_2695,In_1675,In_548);
or U2696 (N_2696,In_793,In_3896);
nor U2697 (N_2697,In_2331,In_3623);
nor U2698 (N_2698,In_485,In_3030);
nand U2699 (N_2699,In_1140,In_936);
or U2700 (N_2700,In_808,In_2058);
or U2701 (N_2701,In_4803,In_372);
and U2702 (N_2702,In_1843,In_4504);
nand U2703 (N_2703,In_43,In_4473);
and U2704 (N_2704,In_4688,In_4344);
nand U2705 (N_2705,In_2188,In_4140);
nand U2706 (N_2706,In_2302,In_1708);
nand U2707 (N_2707,In_1493,In_4162);
nand U2708 (N_2708,In_1651,In_2980);
or U2709 (N_2709,In_4857,In_553);
or U2710 (N_2710,In_1350,In_2814);
nor U2711 (N_2711,In_4226,In_2119);
and U2712 (N_2712,In_1101,In_4407);
xnor U2713 (N_2713,In_524,In_3726);
and U2714 (N_2714,In_3130,In_352);
or U2715 (N_2715,In_881,In_4268);
and U2716 (N_2716,In_832,In_2992);
or U2717 (N_2717,In_1989,In_4636);
or U2718 (N_2718,In_1632,In_4344);
and U2719 (N_2719,In_2479,In_3053);
or U2720 (N_2720,In_2216,In_249);
and U2721 (N_2721,In_1741,In_954);
and U2722 (N_2722,In_1805,In_2146);
nor U2723 (N_2723,In_3655,In_1034);
nand U2724 (N_2724,In_344,In_4345);
or U2725 (N_2725,In_3601,In_4129);
nor U2726 (N_2726,In_2957,In_1250);
nor U2727 (N_2727,In_2705,In_4930);
xnor U2728 (N_2728,In_3536,In_2312);
and U2729 (N_2729,In_3087,In_3132);
xnor U2730 (N_2730,In_30,In_2990);
nor U2731 (N_2731,In_4468,In_2184);
and U2732 (N_2732,In_1763,In_1497);
nand U2733 (N_2733,In_4573,In_256);
xnor U2734 (N_2734,In_2101,In_3126);
nand U2735 (N_2735,In_414,In_3110);
nand U2736 (N_2736,In_3651,In_4927);
xor U2737 (N_2737,In_2826,In_1125);
and U2738 (N_2738,In_3797,In_2014);
nand U2739 (N_2739,In_4276,In_1004);
and U2740 (N_2740,In_4375,In_2389);
and U2741 (N_2741,In_4690,In_442);
nand U2742 (N_2742,In_1281,In_941);
nor U2743 (N_2743,In_2840,In_1930);
xnor U2744 (N_2744,In_4917,In_2419);
and U2745 (N_2745,In_2999,In_3375);
and U2746 (N_2746,In_4558,In_2859);
or U2747 (N_2747,In_4606,In_1081);
nor U2748 (N_2748,In_29,In_4741);
and U2749 (N_2749,In_4153,In_196);
nand U2750 (N_2750,In_4525,In_4371);
and U2751 (N_2751,In_2642,In_586);
nor U2752 (N_2752,In_3808,In_3870);
or U2753 (N_2753,In_2052,In_3899);
and U2754 (N_2754,In_2853,In_3394);
xor U2755 (N_2755,In_3133,In_2485);
and U2756 (N_2756,In_3214,In_4351);
nor U2757 (N_2757,In_1971,In_33);
or U2758 (N_2758,In_49,In_2466);
nand U2759 (N_2759,In_604,In_1051);
xnor U2760 (N_2760,In_1359,In_3689);
xor U2761 (N_2761,In_4610,In_4133);
nand U2762 (N_2762,In_4080,In_3007);
and U2763 (N_2763,In_1282,In_3504);
nor U2764 (N_2764,In_4857,In_351);
and U2765 (N_2765,In_4736,In_1546);
nand U2766 (N_2766,In_3836,In_2378);
or U2767 (N_2767,In_1596,In_1038);
nand U2768 (N_2768,In_950,In_1604);
xor U2769 (N_2769,In_2364,In_2416);
nor U2770 (N_2770,In_552,In_397);
nor U2771 (N_2771,In_270,In_4418);
nor U2772 (N_2772,In_3870,In_509);
or U2773 (N_2773,In_1020,In_757);
nand U2774 (N_2774,In_817,In_1498);
nor U2775 (N_2775,In_235,In_4063);
nor U2776 (N_2776,In_217,In_385);
xnor U2777 (N_2777,In_4873,In_2871);
nand U2778 (N_2778,In_2732,In_3567);
nor U2779 (N_2779,In_2449,In_2972);
nor U2780 (N_2780,In_1943,In_1901);
nand U2781 (N_2781,In_779,In_118);
and U2782 (N_2782,In_2345,In_2295);
or U2783 (N_2783,In_1797,In_840);
and U2784 (N_2784,In_3432,In_3478);
nor U2785 (N_2785,In_4444,In_631);
and U2786 (N_2786,In_4539,In_4523);
or U2787 (N_2787,In_2973,In_4082);
or U2788 (N_2788,In_4304,In_3813);
nor U2789 (N_2789,In_4827,In_333);
or U2790 (N_2790,In_864,In_4457);
and U2791 (N_2791,In_1841,In_4394);
or U2792 (N_2792,In_4827,In_352);
or U2793 (N_2793,In_4315,In_4478);
or U2794 (N_2794,In_776,In_1384);
xor U2795 (N_2795,In_2986,In_4364);
or U2796 (N_2796,In_3549,In_1780);
nor U2797 (N_2797,In_1244,In_1428);
or U2798 (N_2798,In_3462,In_1997);
or U2799 (N_2799,In_4471,In_3814);
xor U2800 (N_2800,In_1626,In_2431);
nor U2801 (N_2801,In_78,In_4375);
or U2802 (N_2802,In_4527,In_4688);
xor U2803 (N_2803,In_2737,In_902);
nor U2804 (N_2804,In_3328,In_1004);
or U2805 (N_2805,In_4141,In_1612);
and U2806 (N_2806,In_4443,In_3848);
nand U2807 (N_2807,In_1226,In_4766);
or U2808 (N_2808,In_3134,In_708);
nand U2809 (N_2809,In_637,In_2047);
or U2810 (N_2810,In_569,In_2347);
or U2811 (N_2811,In_3399,In_3691);
nand U2812 (N_2812,In_1253,In_294);
nand U2813 (N_2813,In_4759,In_753);
nor U2814 (N_2814,In_4744,In_2399);
nand U2815 (N_2815,In_1797,In_1412);
nand U2816 (N_2816,In_3070,In_1243);
or U2817 (N_2817,In_4766,In_3455);
nand U2818 (N_2818,In_4829,In_930);
nand U2819 (N_2819,In_972,In_1351);
nand U2820 (N_2820,In_3582,In_2225);
nand U2821 (N_2821,In_868,In_321);
and U2822 (N_2822,In_2263,In_1604);
or U2823 (N_2823,In_964,In_1860);
or U2824 (N_2824,In_1277,In_4662);
nand U2825 (N_2825,In_4352,In_4244);
xor U2826 (N_2826,In_4384,In_3270);
nor U2827 (N_2827,In_3965,In_3308);
xnor U2828 (N_2828,In_3728,In_3892);
nor U2829 (N_2829,In_3809,In_1116);
nor U2830 (N_2830,In_2927,In_1717);
xor U2831 (N_2831,In_4181,In_3618);
and U2832 (N_2832,In_4754,In_1744);
xnor U2833 (N_2833,In_4865,In_3812);
xor U2834 (N_2834,In_1812,In_291);
xor U2835 (N_2835,In_1697,In_2644);
and U2836 (N_2836,In_1999,In_4390);
or U2837 (N_2837,In_3121,In_3700);
and U2838 (N_2838,In_2627,In_3805);
or U2839 (N_2839,In_3194,In_3954);
xnor U2840 (N_2840,In_4798,In_1356);
xor U2841 (N_2841,In_443,In_993);
nor U2842 (N_2842,In_2270,In_3455);
xor U2843 (N_2843,In_1446,In_3027);
and U2844 (N_2844,In_1583,In_310);
nand U2845 (N_2845,In_3901,In_4714);
and U2846 (N_2846,In_2197,In_2521);
and U2847 (N_2847,In_1311,In_4927);
nand U2848 (N_2848,In_1451,In_4302);
or U2849 (N_2849,In_3194,In_174);
nor U2850 (N_2850,In_2465,In_1635);
nor U2851 (N_2851,In_3,In_1906);
nand U2852 (N_2852,In_2455,In_1430);
xnor U2853 (N_2853,In_4022,In_262);
nand U2854 (N_2854,In_141,In_473);
xor U2855 (N_2855,In_4385,In_2337);
nor U2856 (N_2856,In_2669,In_469);
nand U2857 (N_2857,In_2490,In_4064);
or U2858 (N_2858,In_2905,In_280);
nand U2859 (N_2859,In_1239,In_701);
or U2860 (N_2860,In_3254,In_1606);
or U2861 (N_2861,In_1005,In_4529);
xnor U2862 (N_2862,In_4356,In_2748);
or U2863 (N_2863,In_3164,In_910);
and U2864 (N_2864,In_2974,In_3242);
or U2865 (N_2865,In_2791,In_403);
nor U2866 (N_2866,In_4255,In_4078);
nor U2867 (N_2867,In_3608,In_3921);
xor U2868 (N_2868,In_4685,In_3531);
and U2869 (N_2869,In_169,In_617);
xnor U2870 (N_2870,In_334,In_3803);
or U2871 (N_2871,In_2622,In_4127);
and U2872 (N_2872,In_1966,In_1955);
xnor U2873 (N_2873,In_2586,In_4705);
or U2874 (N_2874,In_636,In_3762);
nand U2875 (N_2875,In_2268,In_1536);
or U2876 (N_2876,In_2145,In_27);
xor U2877 (N_2877,In_890,In_3299);
or U2878 (N_2878,In_2124,In_4297);
nand U2879 (N_2879,In_4880,In_2997);
or U2880 (N_2880,In_927,In_2373);
nor U2881 (N_2881,In_231,In_2049);
xnor U2882 (N_2882,In_2480,In_3791);
nor U2883 (N_2883,In_2234,In_677);
xnor U2884 (N_2884,In_1642,In_4880);
and U2885 (N_2885,In_3069,In_4218);
xor U2886 (N_2886,In_3652,In_1158);
and U2887 (N_2887,In_894,In_4383);
xnor U2888 (N_2888,In_2859,In_414);
nand U2889 (N_2889,In_58,In_4098);
nor U2890 (N_2890,In_1528,In_4014);
nor U2891 (N_2891,In_1571,In_1713);
nand U2892 (N_2892,In_3034,In_849);
nand U2893 (N_2893,In_118,In_1089);
nand U2894 (N_2894,In_2458,In_1897);
and U2895 (N_2895,In_4344,In_4963);
or U2896 (N_2896,In_1908,In_4787);
xor U2897 (N_2897,In_4588,In_197);
or U2898 (N_2898,In_4231,In_844);
nor U2899 (N_2899,In_3781,In_1847);
xnor U2900 (N_2900,In_3149,In_3118);
and U2901 (N_2901,In_1221,In_1500);
nor U2902 (N_2902,In_2589,In_4953);
nor U2903 (N_2903,In_153,In_1832);
xor U2904 (N_2904,In_2678,In_1546);
or U2905 (N_2905,In_1490,In_1771);
and U2906 (N_2906,In_1880,In_3521);
xnor U2907 (N_2907,In_1766,In_4278);
or U2908 (N_2908,In_3026,In_3238);
and U2909 (N_2909,In_4855,In_971);
and U2910 (N_2910,In_734,In_1843);
nand U2911 (N_2911,In_2375,In_3527);
or U2912 (N_2912,In_2537,In_4956);
or U2913 (N_2913,In_3858,In_4149);
nand U2914 (N_2914,In_4921,In_1564);
and U2915 (N_2915,In_3385,In_3928);
nand U2916 (N_2916,In_4790,In_1168);
and U2917 (N_2917,In_3821,In_933);
xnor U2918 (N_2918,In_3529,In_2890);
nand U2919 (N_2919,In_4683,In_4895);
and U2920 (N_2920,In_4334,In_813);
nor U2921 (N_2921,In_2187,In_1799);
nor U2922 (N_2922,In_2873,In_1603);
and U2923 (N_2923,In_3314,In_3894);
and U2924 (N_2924,In_1986,In_1473);
or U2925 (N_2925,In_3709,In_4029);
nor U2926 (N_2926,In_477,In_219);
xor U2927 (N_2927,In_452,In_4991);
xnor U2928 (N_2928,In_4340,In_3030);
nor U2929 (N_2929,In_540,In_1859);
and U2930 (N_2930,In_2005,In_4395);
and U2931 (N_2931,In_343,In_2051);
nor U2932 (N_2932,In_2082,In_147);
nand U2933 (N_2933,In_226,In_4733);
xnor U2934 (N_2934,In_4918,In_1231);
nand U2935 (N_2935,In_556,In_4496);
xor U2936 (N_2936,In_3610,In_562);
and U2937 (N_2937,In_1138,In_1024);
and U2938 (N_2938,In_493,In_4616);
and U2939 (N_2939,In_4146,In_880);
xnor U2940 (N_2940,In_673,In_3574);
xor U2941 (N_2941,In_4070,In_1710);
nand U2942 (N_2942,In_669,In_1803);
or U2943 (N_2943,In_746,In_4063);
nor U2944 (N_2944,In_4228,In_2056);
and U2945 (N_2945,In_1210,In_3478);
nor U2946 (N_2946,In_1295,In_4399);
nor U2947 (N_2947,In_638,In_2338);
nor U2948 (N_2948,In_3962,In_1602);
or U2949 (N_2949,In_3169,In_2139);
nor U2950 (N_2950,In_2616,In_591);
nand U2951 (N_2951,In_3575,In_523);
nor U2952 (N_2952,In_4971,In_4076);
nor U2953 (N_2953,In_1835,In_1428);
or U2954 (N_2954,In_2003,In_1005);
nand U2955 (N_2955,In_478,In_2195);
xor U2956 (N_2956,In_4481,In_4614);
and U2957 (N_2957,In_612,In_4182);
or U2958 (N_2958,In_2781,In_3171);
nor U2959 (N_2959,In_1421,In_1254);
or U2960 (N_2960,In_651,In_4646);
nand U2961 (N_2961,In_3825,In_816);
nand U2962 (N_2962,In_3279,In_2364);
nand U2963 (N_2963,In_601,In_4058);
xnor U2964 (N_2964,In_667,In_195);
or U2965 (N_2965,In_52,In_3169);
and U2966 (N_2966,In_443,In_340);
nor U2967 (N_2967,In_4279,In_2354);
or U2968 (N_2968,In_3690,In_4494);
or U2969 (N_2969,In_829,In_285);
or U2970 (N_2970,In_338,In_2517);
nand U2971 (N_2971,In_4789,In_289);
or U2972 (N_2972,In_1323,In_3012);
or U2973 (N_2973,In_4694,In_326);
nand U2974 (N_2974,In_4077,In_2238);
and U2975 (N_2975,In_4408,In_581);
nor U2976 (N_2976,In_1900,In_4008);
or U2977 (N_2977,In_2034,In_4788);
nand U2978 (N_2978,In_2431,In_4676);
or U2979 (N_2979,In_4008,In_3642);
and U2980 (N_2980,In_2662,In_2591);
and U2981 (N_2981,In_3182,In_133);
nor U2982 (N_2982,In_2380,In_4089);
xor U2983 (N_2983,In_2221,In_2119);
or U2984 (N_2984,In_2212,In_78);
nor U2985 (N_2985,In_3905,In_1359);
xor U2986 (N_2986,In_908,In_4660);
nand U2987 (N_2987,In_2637,In_859);
nand U2988 (N_2988,In_2937,In_2993);
and U2989 (N_2989,In_2951,In_4006);
or U2990 (N_2990,In_463,In_3091);
nor U2991 (N_2991,In_1987,In_935);
or U2992 (N_2992,In_3374,In_1315);
and U2993 (N_2993,In_737,In_1212);
xor U2994 (N_2994,In_3057,In_4339);
nor U2995 (N_2995,In_3343,In_4501);
and U2996 (N_2996,In_2766,In_3000);
nor U2997 (N_2997,In_3334,In_1672);
and U2998 (N_2998,In_4433,In_1975);
and U2999 (N_2999,In_3535,In_3872);
nand U3000 (N_3000,In_1453,In_3207);
nor U3001 (N_3001,In_3866,In_1621);
xnor U3002 (N_3002,In_3629,In_198);
xnor U3003 (N_3003,In_3613,In_3869);
or U3004 (N_3004,In_3848,In_2189);
nor U3005 (N_3005,In_1186,In_987);
and U3006 (N_3006,In_1008,In_603);
xor U3007 (N_3007,In_3755,In_2419);
nor U3008 (N_3008,In_3992,In_2195);
nor U3009 (N_3009,In_3125,In_1561);
nor U3010 (N_3010,In_408,In_2786);
nor U3011 (N_3011,In_2352,In_4937);
nor U3012 (N_3012,In_1603,In_4969);
nand U3013 (N_3013,In_2825,In_1282);
nand U3014 (N_3014,In_4802,In_822);
xnor U3015 (N_3015,In_4737,In_4943);
or U3016 (N_3016,In_4457,In_4255);
nand U3017 (N_3017,In_354,In_3857);
nor U3018 (N_3018,In_2320,In_834);
nand U3019 (N_3019,In_3875,In_2177);
or U3020 (N_3020,In_943,In_1836);
nor U3021 (N_3021,In_2196,In_1286);
or U3022 (N_3022,In_1141,In_2899);
nor U3023 (N_3023,In_2422,In_2840);
xor U3024 (N_3024,In_144,In_2105);
and U3025 (N_3025,In_4823,In_1153);
xnor U3026 (N_3026,In_4715,In_4300);
xor U3027 (N_3027,In_508,In_2648);
nor U3028 (N_3028,In_517,In_4564);
and U3029 (N_3029,In_2638,In_3435);
or U3030 (N_3030,In_3858,In_2073);
and U3031 (N_3031,In_2275,In_1898);
or U3032 (N_3032,In_92,In_3718);
or U3033 (N_3033,In_342,In_2162);
or U3034 (N_3034,In_922,In_770);
and U3035 (N_3035,In_2233,In_755);
and U3036 (N_3036,In_46,In_3080);
xor U3037 (N_3037,In_785,In_3625);
and U3038 (N_3038,In_2434,In_703);
and U3039 (N_3039,In_1237,In_2695);
or U3040 (N_3040,In_2683,In_4620);
nor U3041 (N_3041,In_4131,In_1750);
or U3042 (N_3042,In_4817,In_12);
nor U3043 (N_3043,In_938,In_3022);
xor U3044 (N_3044,In_3410,In_1924);
nand U3045 (N_3045,In_3130,In_2874);
or U3046 (N_3046,In_190,In_4058);
xor U3047 (N_3047,In_4136,In_2944);
nor U3048 (N_3048,In_91,In_1992);
or U3049 (N_3049,In_369,In_1287);
nor U3050 (N_3050,In_772,In_2209);
nand U3051 (N_3051,In_4337,In_1151);
nor U3052 (N_3052,In_4479,In_99);
or U3053 (N_3053,In_311,In_2932);
and U3054 (N_3054,In_4385,In_390);
nor U3055 (N_3055,In_676,In_411);
nand U3056 (N_3056,In_1770,In_2265);
and U3057 (N_3057,In_3508,In_1685);
xor U3058 (N_3058,In_2806,In_4511);
nor U3059 (N_3059,In_4596,In_1136);
nand U3060 (N_3060,In_3808,In_4817);
nand U3061 (N_3061,In_2584,In_2762);
and U3062 (N_3062,In_3656,In_573);
xnor U3063 (N_3063,In_4084,In_1308);
and U3064 (N_3064,In_2633,In_1855);
xnor U3065 (N_3065,In_4469,In_582);
and U3066 (N_3066,In_4584,In_3085);
nand U3067 (N_3067,In_4686,In_4030);
xor U3068 (N_3068,In_3649,In_2028);
nor U3069 (N_3069,In_1347,In_3932);
xnor U3070 (N_3070,In_2868,In_110);
or U3071 (N_3071,In_1916,In_1020);
and U3072 (N_3072,In_238,In_2828);
and U3073 (N_3073,In_2991,In_3199);
and U3074 (N_3074,In_3431,In_4065);
nor U3075 (N_3075,In_3392,In_2751);
xnor U3076 (N_3076,In_4898,In_256);
or U3077 (N_3077,In_4339,In_964);
nor U3078 (N_3078,In_1192,In_2415);
xor U3079 (N_3079,In_627,In_4695);
and U3080 (N_3080,In_3634,In_872);
nor U3081 (N_3081,In_711,In_4865);
or U3082 (N_3082,In_1038,In_3112);
and U3083 (N_3083,In_2665,In_647);
nand U3084 (N_3084,In_4151,In_2435);
and U3085 (N_3085,In_4931,In_4250);
nor U3086 (N_3086,In_304,In_1224);
or U3087 (N_3087,In_3977,In_1787);
and U3088 (N_3088,In_1080,In_3015);
xnor U3089 (N_3089,In_3555,In_1254);
xnor U3090 (N_3090,In_1988,In_3321);
nand U3091 (N_3091,In_3546,In_1802);
and U3092 (N_3092,In_1126,In_1286);
and U3093 (N_3093,In_668,In_492);
xor U3094 (N_3094,In_2864,In_2578);
or U3095 (N_3095,In_2369,In_509);
and U3096 (N_3096,In_3641,In_3908);
nand U3097 (N_3097,In_2873,In_1796);
nand U3098 (N_3098,In_2772,In_4680);
or U3099 (N_3099,In_729,In_527);
and U3100 (N_3100,In_1041,In_2046);
xor U3101 (N_3101,In_1391,In_747);
and U3102 (N_3102,In_4017,In_2653);
nand U3103 (N_3103,In_3033,In_3354);
nand U3104 (N_3104,In_2898,In_3140);
and U3105 (N_3105,In_3961,In_3596);
nor U3106 (N_3106,In_138,In_2137);
nand U3107 (N_3107,In_667,In_1110);
xor U3108 (N_3108,In_1245,In_761);
nor U3109 (N_3109,In_3457,In_3145);
nor U3110 (N_3110,In_709,In_172);
and U3111 (N_3111,In_2016,In_2673);
and U3112 (N_3112,In_2895,In_2331);
xnor U3113 (N_3113,In_1342,In_1406);
or U3114 (N_3114,In_1336,In_1829);
xor U3115 (N_3115,In_313,In_3597);
nor U3116 (N_3116,In_409,In_3697);
or U3117 (N_3117,In_898,In_176);
and U3118 (N_3118,In_4554,In_1467);
nand U3119 (N_3119,In_4678,In_3695);
nand U3120 (N_3120,In_4113,In_231);
and U3121 (N_3121,In_3593,In_3880);
nand U3122 (N_3122,In_2221,In_318);
xnor U3123 (N_3123,In_3106,In_4138);
nor U3124 (N_3124,In_2775,In_4572);
nand U3125 (N_3125,In_4088,In_4135);
nand U3126 (N_3126,In_4154,In_2166);
nand U3127 (N_3127,In_411,In_4880);
xor U3128 (N_3128,In_4766,In_590);
nor U3129 (N_3129,In_527,In_4175);
nor U3130 (N_3130,In_1668,In_4060);
nor U3131 (N_3131,In_4858,In_4900);
or U3132 (N_3132,In_4817,In_117);
nand U3133 (N_3133,In_2838,In_4168);
or U3134 (N_3134,In_3136,In_4393);
nand U3135 (N_3135,In_3229,In_3290);
nand U3136 (N_3136,In_3488,In_4914);
xor U3137 (N_3137,In_4682,In_2889);
xor U3138 (N_3138,In_2910,In_4827);
and U3139 (N_3139,In_352,In_1563);
xnor U3140 (N_3140,In_4809,In_3766);
and U3141 (N_3141,In_2136,In_1075);
and U3142 (N_3142,In_4844,In_2116);
or U3143 (N_3143,In_4297,In_4661);
nor U3144 (N_3144,In_4255,In_1739);
xor U3145 (N_3145,In_1513,In_1896);
xnor U3146 (N_3146,In_2148,In_4964);
xor U3147 (N_3147,In_3783,In_861);
and U3148 (N_3148,In_4504,In_3466);
nand U3149 (N_3149,In_1793,In_1203);
nor U3150 (N_3150,In_4207,In_2142);
nor U3151 (N_3151,In_1923,In_49);
xor U3152 (N_3152,In_3639,In_4555);
and U3153 (N_3153,In_3726,In_2585);
xor U3154 (N_3154,In_445,In_1047);
or U3155 (N_3155,In_1901,In_3331);
or U3156 (N_3156,In_1592,In_3238);
nor U3157 (N_3157,In_2003,In_4218);
and U3158 (N_3158,In_385,In_284);
nor U3159 (N_3159,In_2907,In_4240);
nand U3160 (N_3160,In_3911,In_1943);
and U3161 (N_3161,In_1491,In_2769);
nor U3162 (N_3162,In_647,In_3782);
or U3163 (N_3163,In_4467,In_3250);
nand U3164 (N_3164,In_3206,In_3353);
nand U3165 (N_3165,In_4333,In_2648);
nor U3166 (N_3166,In_3153,In_2457);
or U3167 (N_3167,In_3925,In_1164);
or U3168 (N_3168,In_4159,In_469);
nor U3169 (N_3169,In_3763,In_733);
or U3170 (N_3170,In_4596,In_4649);
or U3171 (N_3171,In_4816,In_891);
and U3172 (N_3172,In_868,In_1921);
xnor U3173 (N_3173,In_2639,In_3780);
or U3174 (N_3174,In_3959,In_1347);
xnor U3175 (N_3175,In_3358,In_4378);
xnor U3176 (N_3176,In_3258,In_3731);
nor U3177 (N_3177,In_1224,In_4234);
nand U3178 (N_3178,In_3430,In_1706);
xor U3179 (N_3179,In_2844,In_1889);
nand U3180 (N_3180,In_967,In_4662);
xnor U3181 (N_3181,In_4001,In_2486);
nand U3182 (N_3182,In_290,In_1938);
and U3183 (N_3183,In_177,In_564);
and U3184 (N_3184,In_1168,In_2661);
nand U3185 (N_3185,In_1596,In_4504);
or U3186 (N_3186,In_1528,In_2992);
and U3187 (N_3187,In_785,In_784);
nand U3188 (N_3188,In_2987,In_16);
xnor U3189 (N_3189,In_4798,In_596);
and U3190 (N_3190,In_116,In_4970);
or U3191 (N_3191,In_893,In_548);
and U3192 (N_3192,In_850,In_546);
or U3193 (N_3193,In_1710,In_1794);
xor U3194 (N_3194,In_789,In_450);
and U3195 (N_3195,In_4309,In_2552);
nor U3196 (N_3196,In_4765,In_2642);
nor U3197 (N_3197,In_305,In_4970);
and U3198 (N_3198,In_2718,In_4653);
nor U3199 (N_3199,In_2806,In_4059);
or U3200 (N_3200,In_2926,In_167);
xnor U3201 (N_3201,In_4570,In_4439);
xnor U3202 (N_3202,In_3579,In_1452);
and U3203 (N_3203,In_147,In_2161);
nor U3204 (N_3204,In_3847,In_1879);
nor U3205 (N_3205,In_1267,In_1844);
xnor U3206 (N_3206,In_833,In_4919);
and U3207 (N_3207,In_4199,In_3891);
and U3208 (N_3208,In_708,In_2421);
xor U3209 (N_3209,In_487,In_3783);
nand U3210 (N_3210,In_2529,In_2401);
and U3211 (N_3211,In_3681,In_4789);
xor U3212 (N_3212,In_544,In_4746);
nor U3213 (N_3213,In_2193,In_2825);
and U3214 (N_3214,In_3598,In_4536);
nor U3215 (N_3215,In_4170,In_4702);
nor U3216 (N_3216,In_406,In_1636);
nor U3217 (N_3217,In_4431,In_1991);
and U3218 (N_3218,In_4499,In_455);
xnor U3219 (N_3219,In_3331,In_2351);
nand U3220 (N_3220,In_488,In_797);
xor U3221 (N_3221,In_2717,In_1341);
nor U3222 (N_3222,In_3145,In_1790);
xor U3223 (N_3223,In_4218,In_1888);
xor U3224 (N_3224,In_59,In_543);
nand U3225 (N_3225,In_4388,In_4216);
nor U3226 (N_3226,In_967,In_391);
nand U3227 (N_3227,In_4051,In_4058);
and U3228 (N_3228,In_2408,In_4626);
or U3229 (N_3229,In_1695,In_4087);
and U3230 (N_3230,In_3494,In_2145);
nor U3231 (N_3231,In_4826,In_4195);
or U3232 (N_3232,In_2937,In_3818);
nand U3233 (N_3233,In_1346,In_2216);
nand U3234 (N_3234,In_3727,In_2758);
xor U3235 (N_3235,In_3720,In_1817);
or U3236 (N_3236,In_794,In_3250);
xnor U3237 (N_3237,In_4807,In_3459);
and U3238 (N_3238,In_2429,In_3122);
nand U3239 (N_3239,In_337,In_2871);
or U3240 (N_3240,In_1467,In_3913);
nor U3241 (N_3241,In_3728,In_3971);
nand U3242 (N_3242,In_2961,In_4796);
nand U3243 (N_3243,In_1335,In_3513);
nor U3244 (N_3244,In_1974,In_323);
nand U3245 (N_3245,In_3076,In_3298);
nand U3246 (N_3246,In_840,In_4563);
or U3247 (N_3247,In_3804,In_3249);
xnor U3248 (N_3248,In_2589,In_2775);
nand U3249 (N_3249,In_4393,In_963);
nand U3250 (N_3250,In_4583,In_1001);
nor U3251 (N_3251,In_4509,In_3739);
xnor U3252 (N_3252,In_3839,In_3709);
nor U3253 (N_3253,In_2019,In_1152);
nand U3254 (N_3254,In_3645,In_664);
nor U3255 (N_3255,In_1004,In_2579);
nand U3256 (N_3256,In_3689,In_2726);
or U3257 (N_3257,In_1799,In_2899);
nor U3258 (N_3258,In_4846,In_1589);
xnor U3259 (N_3259,In_238,In_4848);
and U3260 (N_3260,In_2769,In_364);
xor U3261 (N_3261,In_2991,In_2161);
or U3262 (N_3262,In_3133,In_3950);
xnor U3263 (N_3263,In_1568,In_2989);
xnor U3264 (N_3264,In_4630,In_4014);
nand U3265 (N_3265,In_3877,In_706);
nor U3266 (N_3266,In_1768,In_3764);
and U3267 (N_3267,In_1150,In_2457);
nand U3268 (N_3268,In_281,In_4730);
nor U3269 (N_3269,In_22,In_4003);
or U3270 (N_3270,In_4416,In_3556);
xor U3271 (N_3271,In_3868,In_1090);
nand U3272 (N_3272,In_2567,In_719);
nand U3273 (N_3273,In_1663,In_4719);
nand U3274 (N_3274,In_4985,In_216);
or U3275 (N_3275,In_2985,In_4902);
xor U3276 (N_3276,In_1137,In_2554);
nand U3277 (N_3277,In_3924,In_2939);
nor U3278 (N_3278,In_3789,In_1045);
xor U3279 (N_3279,In_4165,In_1692);
nand U3280 (N_3280,In_383,In_4186);
or U3281 (N_3281,In_2512,In_2853);
nand U3282 (N_3282,In_3852,In_2049);
and U3283 (N_3283,In_2700,In_3755);
nor U3284 (N_3284,In_3796,In_4143);
xor U3285 (N_3285,In_3748,In_1750);
nor U3286 (N_3286,In_2800,In_2216);
or U3287 (N_3287,In_1206,In_2606);
or U3288 (N_3288,In_3216,In_941);
nor U3289 (N_3289,In_4755,In_1125);
xor U3290 (N_3290,In_322,In_216);
and U3291 (N_3291,In_1923,In_804);
and U3292 (N_3292,In_555,In_4651);
xor U3293 (N_3293,In_1928,In_3834);
nor U3294 (N_3294,In_774,In_1165);
nor U3295 (N_3295,In_3099,In_85);
and U3296 (N_3296,In_3330,In_4693);
nand U3297 (N_3297,In_4595,In_450);
nand U3298 (N_3298,In_287,In_946);
xor U3299 (N_3299,In_937,In_936);
and U3300 (N_3300,In_3100,In_4584);
and U3301 (N_3301,In_2352,In_1513);
nor U3302 (N_3302,In_2822,In_1173);
xnor U3303 (N_3303,In_2142,In_2114);
nor U3304 (N_3304,In_848,In_3681);
nand U3305 (N_3305,In_3066,In_1175);
nor U3306 (N_3306,In_1999,In_873);
nand U3307 (N_3307,In_1308,In_753);
xnor U3308 (N_3308,In_3208,In_1852);
nand U3309 (N_3309,In_352,In_3388);
xor U3310 (N_3310,In_4720,In_3532);
and U3311 (N_3311,In_1425,In_4260);
nor U3312 (N_3312,In_4751,In_37);
or U3313 (N_3313,In_2123,In_1830);
or U3314 (N_3314,In_946,In_1422);
nor U3315 (N_3315,In_3592,In_3037);
nand U3316 (N_3316,In_2149,In_3249);
xor U3317 (N_3317,In_4071,In_2217);
nor U3318 (N_3318,In_3778,In_2336);
and U3319 (N_3319,In_2473,In_4064);
or U3320 (N_3320,In_1410,In_1023);
nor U3321 (N_3321,In_1834,In_952);
and U3322 (N_3322,In_1490,In_2693);
nand U3323 (N_3323,In_2116,In_3098);
nor U3324 (N_3324,In_2085,In_4362);
or U3325 (N_3325,In_3299,In_3356);
and U3326 (N_3326,In_2423,In_4497);
xor U3327 (N_3327,In_1917,In_2248);
nor U3328 (N_3328,In_70,In_4266);
or U3329 (N_3329,In_3600,In_4116);
or U3330 (N_3330,In_18,In_322);
and U3331 (N_3331,In_1510,In_1613);
xor U3332 (N_3332,In_3253,In_3491);
nor U3333 (N_3333,In_2629,In_23);
xnor U3334 (N_3334,In_1042,In_1227);
nand U3335 (N_3335,In_517,In_3877);
or U3336 (N_3336,In_4034,In_2525);
xnor U3337 (N_3337,In_858,In_4350);
or U3338 (N_3338,In_330,In_1804);
or U3339 (N_3339,In_4630,In_2842);
or U3340 (N_3340,In_111,In_1683);
nand U3341 (N_3341,In_2172,In_4905);
nor U3342 (N_3342,In_2336,In_253);
nand U3343 (N_3343,In_3382,In_3166);
and U3344 (N_3344,In_3301,In_4025);
or U3345 (N_3345,In_4115,In_3461);
or U3346 (N_3346,In_67,In_4455);
or U3347 (N_3347,In_1964,In_2482);
nand U3348 (N_3348,In_3821,In_1440);
nor U3349 (N_3349,In_1501,In_3084);
and U3350 (N_3350,In_1341,In_2683);
and U3351 (N_3351,In_1570,In_670);
nor U3352 (N_3352,In_1849,In_4960);
nor U3353 (N_3353,In_2237,In_2336);
or U3354 (N_3354,In_111,In_3647);
nor U3355 (N_3355,In_1727,In_2926);
nor U3356 (N_3356,In_1330,In_1555);
or U3357 (N_3357,In_1437,In_860);
nor U3358 (N_3358,In_3431,In_2457);
or U3359 (N_3359,In_4866,In_3320);
and U3360 (N_3360,In_2292,In_683);
nor U3361 (N_3361,In_413,In_1141);
nand U3362 (N_3362,In_306,In_1283);
or U3363 (N_3363,In_3004,In_2699);
nor U3364 (N_3364,In_3892,In_2117);
nor U3365 (N_3365,In_3676,In_3674);
xor U3366 (N_3366,In_1126,In_1536);
xnor U3367 (N_3367,In_818,In_4673);
xnor U3368 (N_3368,In_3957,In_2006);
or U3369 (N_3369,In_985,In_859);
or U3370 (N_3370,In_2669,In_4201);
nand U3371 (N_3371,In_1823,In_2257);
nand U3372 (N_3372,In_402,In_694);
nand U3373 (N_3373,In_717,In_2932);
and U3374 (N_3374,In_434,In_4738);
or U3375 (N_3375,In_564,In_2240);
xnor U3376 (N_3376,In_916,In_3609);
nand U3377 (N_3377,In_206,In_680);
and U3378 (N_3378,In_4363,In_429);
or U3379 (N_3379,In_645,In_3499);
xnor U3380 (N_3380,In_4205,In_3154);
xor U3381 (N_3381,In_2994,In_1106);
nor U3382 (N_3382,In_4282,In_978);
nor U3383 (N_3383,In_326,In_1059);
xnor U3384 (N_3384,In_1157,In_2643);
xnor U3385 (N_3385,In_4357,In_2438);
and U3386 (N_3386,In_4838,In_3781);
xor U3387 (N_3387,In_2651,In_2161);
nand U3388 (N_3388,In_4465,In_2072);
xor U3389 (N_3389,In_1326,In_645);
nor U3390 (N_3390,In_1899,In_4339);
and U3391 (N_3391,In_2796,In_166);
or U3392 (N_3392,In_1049,In_1293);
and U3393 (N_3393,In_3901,In_359);
nand U3394 (N_3394,In_1952,In_351);
xor U3395 (N_3395,In_4073,In_2100);
nand U3396 (N_3396,In_1192,In_2443);
nor U3397 (N_3397,In_3096,In_2640);
nand U3398 (N_3398,In_3527,In_350);
nor U3399 (N_3399,In_671,In_4301);
nor U3400 (N_3400,In_2655,In_2108);
or U3401 (N_3401,In_1243,In_29);
xnor U3402 (N_3402,In_732,In_207);
nor U3403 (N_3403,In_4281,In_1181);
and U3404 (N_3404,In_3470,In_1243);
xor U3405 (N_3405,In_1945,In_3626);
nor U3406 (N_3406,In_4522,In_4337);
and U3407 (N_3407,In_1088,In_1945);
xnor U3408 (N_3408,In_4,In_3961);
and U3409 (N_3409,In_3669,In_3841);
or U3410 (N_3410,In_680,In_3063);
or U3411 (N_3411,In_2463,In_4132);
or U3412 (N_3412,In_3188,In_4065);
and U3413 (N_3413,In_36,In_2618);
or U3414 (N_3414,In_66,In_1999);
xor U3415 (N_3415,In_628,In_3275);
nor U3416 (N_3416,In_1412,In_592);
or U3417 (N_3417,In_2938,In_2647);
xnor U3418 (N_3418,In_1734,In_2067);
xor U3419 (N_3419,In_1187,In_4224);
nand U3420 (N_3420,In_1125,In_3567);
nor U3421 (N_3421,In_2049,In_4796);
and U3422 (N_3422,In_637,In_977);
and U3423 (N_3423,In_4955,In_1196);
nor U3424 (N_3424,In_3990,In_1255);
and U3425 (N_3425,In_1868,In_1907);
nand U3426 (N_3426,In_3298,In_3240);
xor U3427 (N_3427,In_1819,In_2310);
and U3428 (N_3428,In_3685,In_1858);
or U3429 (N_3429,In_3296,In_1008);
or U3430 (N_3430,In_4863,In_2723);
nand U3431 (N_3431,In_3357,In_905);
and U3432 (N_3432,In_2339,In_3206);
nor U3433 (N_3433,In_1625,In_3924);
xnor U3434 (N_3434,In_4832,In_2555);
and U3435 (N_3435,In_517,In_4089);
or U3436 (N_3436,In_1825,In_4289);
nor U3437 (N_3437,In_3182,In_3503);
xor U3438 (N_3438,In_325,In_3834);
nand U3439 (N_3439,In_3815,In_3072);
and U3440 (N_3440,In_55,In_1786);
or U3441 (N_3441,In_2584,In_2801);
nor U3442 (N_3442,In_359,In_2825);
nor U3443 (N_3443,In_892,In_4047);
or U3444 (N_3444,In_4534,In_124);
nor U3445 (N_3445,In_513,In_4483);
nor U3446 (N_3446,In_453,In_2472);
and U3447 (N_3447,In_3583,In_4935);
xor U3448 (N_3448,In_2468,In_1703);
nor U3449 (N_3449,In_4765,In_3447);
and U3450 (N_3450,In_3631,In_4089);
nand U3451 (N_3451,In_222,In_4304);
and U3452 (N_3452,In_513,In_1881);
nor U3453 (N_3453,In_1070,In_3765);
and U3454 (N_3454,In_3213,In_2723);
nor U3455 (N_3455,In_4495,In_3391);
and U3456 (N_3456,In_2447,In_468);
or U3457 (N_3457,In_1928,In_3344);
or U3458 (N_3458,In_4060,In_813);
nand U3459 (N_3459,In_1933,In_1500);
nor U3460 (N_3460,In_1021,In_2605);
and U3461 (N_3461,In_1145,In_2982);
nand U3462 (N_3462,In_2389,In_1135);
and U3463 (N_3463,In_1388,In_976);
nand U3464 (N_3464,In_4544,In_3630);
or U3465 (N_3465,In_13,In_3170);
nor U3466 (N_3466,In_3389,In_1236);
nand U3467 (N_3467,In_3112,In_3525);
or U3468 (N_3468,In_3597,In_1468);
xnor U3469 (N_3469,In_4772,In_4303);
nor U3470 (N_3470,In_4490,In_3041);
nor U3471 (N_3471,In_1681,In_475);
nor U3472 (N_3472,In_3552,In_876);
or U3473 (N_3473,In_3275,In_746);
and U3474 (N_3474,In_4618,In_3374);
nand U3475 (N_3475,In_4040,In_284);
xor U3476 (N_3476,In_1818,In_2077);
or U3477 (N_3477,In_3727,In_561);
nand U3478 (N_3478,In_4037,In_3531);
nand U3479 (N_3479,In_3852,In_3370);
nor U3480 (N_3480,In_3752,In_3553);
or U3481 (N_3481,In_3799,In_114);
nor U3482 (N_3482,In_4347,In_2842);
nor U3483 (N_3483,In_4276,In_2709);
or U3484 (N_3484,In_2024,In_112);
nor U3485 (N_3485,In_3909,In_4193);
nand U3486 (N_3486,In_4506,In_1260);
and U3487 (N_3487,In_4588,In_4887);
nor U3488 (N_3488,In_1953,In_4240);
nor U3489 (N_3489,In_1708,In_15);
nand U3490 (N_3490,In_2249,In_2948);
nor U3491 (N_3491,In_2101,In_2636);
and U3492 (N_3492,In_4768,In_2929);
or U3493 (N_3493,In_97,In_2987);
or U3494 (N_3494,In_3341,In_163);
nor U3495 (N_3495,In_3570,In_1280);
and U3496 (N_3496,In_4060,In_3665);
and U3497 (N_3497,In_2297,In_4401);
nand U3498 (N_3498,In_2083,In_429);
and U3499 (N_3499,In_125,In_3583);
and U3500 (N_3500,In_731,In_1238);
or U3501 (N_3501,In_1588,In_192);
nand U3502 (N_3502,In_2301,In_21);
xnor U3503 (N_3503,In_628,In_3778);
or U3504 (N_3504,In_0,In_1371);
nand U3505 (N_3505,In_393,In_1648);
xor U3506 (N_3506,In_4944,In_4990);
or U3507 (N_3507,In_726,In_4316);
xnor U3508 (N_3508,In_137,In_4495);
xnor U3509 (N_3509,In_4483,In_1374);
nor U3510 (N_3510,In_845,In_1570);
nand U3511 (N_3511,In_3004,In_1005);
nand U3512 (N_3512,In_1773,In_1717);
xnor U3513 (N_3513,In_216,In_1164);
xor U3514 (N_3514,In_3277,In_939);
nand U3515 (N_3515,In_977,In_340);
and U3516 (N_3516,In_229,In_2379);
or U3517 (N_3517,In_230,In_591);
nand U3518 (N_3518,In_1795,In_1438);
or U3519 (N_3519,In_1699,In_3320);
or U3520 (N_3520,In_2821,In_2808);
and U3521 (N_3521,In_2318,In_517);
xor U3522 (N_3522,In_3778,In_4418);
or U3523 (N_3523,In_342,In_3077);
or U3524 (N_3524,In_1096,In_3086);
nor U3525 (N_3525,In_2635,In_1477);
xor U3526 (N_3526,In_1884,In_4040);
xnor U3527 (N_3527,In_4331,In_3157);
and U3528 (N_3528,In_798,In_4003);
or U3529 (N_3529,In_3661,In_1472);
nand U3530 (N_3530,In_2270,In_1660);
nand U3531 (N_3531,In_3576,In_4015);
and U3532 (N_3532,In_2176,In_4000);
and U3533 (N_3533,In_1782,In_2782);
xor U3534 (N_3534,In_2707,In_1814);
xor U3535 (N_3535,In_725,In_844);
or U3536 (N_3536,In_3403,In_4590);
and U3537 (N_3537,In_1775,In_4530);
nor U3538 (N_3538,In_2401,In_67);
xor U3539 (N_3539,In_2285,In_4538);
or U3540 (N_3540,In_3367,In_129);
and U3541 (N_3541,In_4573,In_2792);
nor U3542 (N_3542,In_1772,In_1473);
or U3543 (N_3543,In_4397,In_0);
or U3544 (N_3544,In_4734,In_4132);
xnor U3545 (N_3545,In_1672,In_3704);
nor U3546 (N_3546,In_1397,In_2719);
nor U3547 (N_3547,In_4459,In_1740);
or U3548 (N_3548,In_585,In_394);
and U3549 (N_3549,In_1231,In_2130);
or U3550 (N_3550,In_3537,In_4762);
nand U3551 (N_3551,In_1531,In_2714);
or U3552 (N_3552,In_3468,In_3248);
and U3553 (N_3553,In_4527,In_651);
xor U3554 (N_3554,In_1248,In_983);
xnor U3555 (N_3555,In_3920,In_549);
or U3556 (N_3556,In_3701,In_1049);
xnor U3557 (N_3557,In_111,In_1097);
xor U3558 (N_3558,In_82,In_503);
xor U3559 (N_3559,In_2083,In_2805);
nand U3560 (N_3560,In_2827,In_3675);
or U3561 (N_3561,In_4757,In_3634);
and U3562 (N_3562,In_1418,In_2526);
and U3563 (N_3563,In_4568,In_4593);
nand U3564 (N_3564,In_348,In_2449);
nand U3565 (N_3565,In_456,In_2268);
nand U3566 (N_3566,In_798,In_3282);
nand U3567 (N_3567,In_4730,In_2800);
or U3568 (N_3568,In_1442,In_3890);
or U3569 (N_3569,In_3657,In_4605);
and U3570 (N_3570,In_2269,In_3350);
nand U3571 (N_3571,In_3163,In_1081);
or U3572 (N_3572,In_623,In_4459);
or U3573 (N_3573,In_439,In_1989);
or U3574 (N_3574,In_3688,In_717);
nor U3575 (N_3575,In_3210,In_491);
nand U3576 (N_3576,In_3212,In_3022);
nand U3577 (N_3577,In_2071,In_1547);
nor U3578 (N_3578,In_3614,In_963);
and U3579 (N_3579,In_4283,In_4922);
nor U3580 (N_3580,In_4811,In_1482);
or U3581 (N_3581,In_715,In_2552);
or U3582 (N_3582,In_406,In_1531);
or U3583 (N_3583,In_4310,In_2443);
nor U3584 (N_3584,In_2638,In_4043);
nor U3585 (N_3585,In_4391,In_2634);
nand U3586 (N_3586,In_74,In_3895);
nand U3587 (N_3587,In_3915,In_515);
nand U3588 (N_3588,In_2855,In_2269);
nor U3589 (N_3589,In_1678,In_4173);
nand U3590 (N_3590,In_197,In_4633);
nor U3591 (N_3591,In_1674,In_3889);
nand U3592 (N_3592,In_1357,In_731);
and U3593 (N_3593,In_3297,In_4738);
and U3594 (N_3594,In_1776,In_1348);
or U3595 (N_3595,In_2096,In_3252);
and U3596 (N_3596,In_2719,In_3609);
nand U3597 (N_3597,In_3028,In_2687);
xor U3598 (N_3598,In_2044,In_182);
and U3599 (N_3599,In_1162,In_4755);
or U3600 (N_3600,In_3205,In_4529);
nor U3601 (N_3601,In_4079,In_2769);
or U3602 (N_3602,In_2096,In_3577);
nand U3603 (N_3603,In_2647,In_2020);
nor U3604 (N_3604,In_997,In_944);
and U3605 (N_3605,In_2147,In_3471);
or U3606 (N_3606,In_3464,In_1661);
nor U3607 (N_3607,In_2913,In_2427);
and U3608 (N_3608,In_3953,In_3666);
nor U3609 (N_3609,In_4296,In_3490);
nor U3610 (N_3610,In_3056,In_3104);
xor U3611 (N_3611,In_2261,In_4041);
xor U3612 (N_3612,In_1382,In_221);
and U3613 (N_3613,In_2483,In_4154);
nand U3614 (N_3614,In_4538,In_1621);
xor U3615 (N_3615,In_2238,In_2197);
xor U3616 (N_3616,In_342,In_549);
or U3617 (N_3617,In_3543,In_997);
nor U3618 (N_3618,In_4068,In_4174);
and U3619 (N_3619,In_2850,In_4424);
nand U3620 (N_3620,In_891,In_2479);
nor U3621 (N_3621,In_1654,In_1765);
or U3622 (N_3622,In_4455,In_125);
or U3623 (N_3623,In_890,In_490);
nand U3624 (N_3624,In_4576,In_520);
or U3625 (N_3625,In_4675,In_1958);
and U3626 (N_3626,In_4856,In_2462);
and U3627 (N_3627,In_452,In_3136);
xnor U3628 (N_3628,In_688,In_760);
nand U3629 (N_3629,In_2008,In_4120);
nand U3630 (N_3630,In_3062,In_381);
and U3631 (N_3631,In_3004,In_855);
and U3632 (N_3632,In_1314,In_2982);
and U3633 (N_3633,In_1426,In_1741);
or U3634 (N_3634,In_626,In_952);
nand U3635 (N_3635,In_3914,In_3295);
and U3636 (N_3636,In_4525,In_2577);
xor U3637 (N_3637,In_4615,In_4608);
xnor U3638 (N_3638,In_3693,In_915);
or U3639 (N_3639,In_3642,In_1456);
xnor U3640 (N_3640,In_4747,In_3407);
and U3641 (N_3641,In_4079,In_4609);
or U3642 (N_3642,In_1862,In_2219);
xor U3643 (N_3643,In_3825,In_702);
xor U3644 (N_3644,In_3273,In_1446);
and U3645 (N_3645,In_2944,In_2081);
nor U3646 (N_3646,In_1451,In_1196);
nor U3647 (N_3647,In_4669,In_1750);
xnor U3648 (N_3648,In_2526,In_1908);
or U3649 (N_3649,In_1995,In_3284);
nor U3650 (N_3650,In_4462,In_3137);
nand U3651 (N_3651,In_2877,In_1619);
nand U3652 (N_3652,In_3423,In_2746);
nor U3653 (N_3653,In_3549,In_910);
nand U3654 (N_3654,In_3015,In_1019);
and U3655 (N_3655,In_4603,In_3433);
nand U3656 (N_3656,In_1720,In_972);
and U3657 (N_3657,In_3016,In_3366);
nand U3658 (N_3658,In_3695,In_2586);
nor U3659 (N_3659,In_1362,In_1131);
nand U3660 (N_3660,In_3976,In_2247);
and U3661 (N_3661,In_2887,In_524);
xor U3662 (N_3662,In_4917,In_3462);
xor U3663 (N_3663,In_2467,In_4497);
nor U3664 (N_3664,In_2217,In_3535);
or U3665 (N_3665,In_3963,In_2722);
nand U3666 (N_3666,In_2572,In_4264);
xor U3667 (N_3667,In_3844,In_254);
nor U3668 (N_3668,In_2805,In_957);
xor U3669 (N_3669,In_1214,In_1456);
or U3670 (N_3670,In_2360,In_2224);
or U3671 (N_3671,In_163,In_1224);
and U3672 (N_3672,In_1501,In_230);
or U3673 (N_3673,In_1345,In_115);
nand U3674 (N_3674,In_521,In_854);
or U3675 (N_3675,In_4822,In_3327);
xor U3676 (N_3676,In_523,In_3316);
xnor U3677 (N_3677,In_2649,In_2864);
or U3678 (N_3678,In_455,In_3253);
or U3679 (N_3679,In_2340,In_3240);
nor U3680 (N_3680,In_3999,In_58);
nand U3681 (N_3681,In_241,In_4427);
or U3682 (N_3682,In_4785,In_1056);
and U3683 (N_3683,In_910,In_4142);
and U3684 (N_3684,In_2074,In_1612);
and U3685 (N_3685,In_903,In_3704);
or U3686 (N_3686,In_4396,In_3313);
and U3687 (N_3687,In_1789,In_17);
xor U3688 (N_3688,In_1565,In_490);
and U3689 (N_3689,In_2632,In_899);
and U3690 (N_3690,In_489,In_2351);
nor U3691 (N_3691,In_3682,In_4326);
nand U3692 (N_3692,In_469,In_1868);
and U3693 (N_3693,In_1070,In_1300);
nor U3694 (N_3694,In_3102,In_1111);
nor U3695 (N_3695,In_3069,In_3691);
or U3696 (N_3696,In_2474,In_4259);
or U3697 (N_3697,In_2180,In_2684);
nor U3698 (N_3698,In_3482,In_4226);
nor U3699 (N_3699,In_477,In_1590);
and U3700 (N_3700,In_4035,In_4652);
xnor U3701 (N_3701,In_4047,In_3679);
and U3702 (N_3702,In_2822,In_4097);
nor U3703 (N_3703,In_4414,In_4223);
and U3704 (N_3704,In_1989,In_4460);
nand U3705 (N_3705,In_1247,In_3357);
or U3706 (N_3706,In_1162,In_818);
nand U3707 (N_3707,In_649,In_3593);
nand U3708 (N_3708,In_3416,In_2360);
and U3709 (N_3709,In_3317,In_4013);
nor U3710 (N_3710,In_468,In_3423);
xor U3711 (N_3711,In_828,In_2810);
and U3712 (N_3712,In_89,In_4522);
xnor U3713 (N_3713,In_2085,In_1582);
nor U3714 (N_3714,In_2401,In_533);
nand U3715 (N_3715,In_2958,In_1901);
or U3716 (N_3716,In_2245,In_1153);
and U3717 (N_3717,In_1650,In_1463);
xnor U3718 (N_3718,In_2480,In_4108);
and U3719 (N_3719,In_54,In_352);
nor U3720 (N_3720,In_4708,In_3415);
or U3721 (N_3721,In_4459,In_3491);
and U3722 (N_3722,In_1515,In_4457);
or U3723 (N_3723,In_4726,In_2880);
and U3724 (N_3724,In_4233,In_245);
and U3725 (N_3725,In_2540,In_865);
or U3726 (N_3726,In_3606,In_4097);
xnor U3727 (N_3727,In_1737,In_861);
or U3728 (N_3728,In_3745,In_3449);
xor U3729 (N_3729,In_2158,In_691);
nor U3730 (N_3730,In_919,In_3861);
nand U3731 (N_3731,In_4503,In_3914);
and U3732 (N_3732,In_4308,In_4000);
xnor U3733 (N_3733,In_60,In_4812);
and U3734 (N_3734,In_1591,In_4538);
or U3735 (N_3735,In_1702,In_4273);
nand U3736 (N_3736,In_546,In_1647);
nand U3737 (N_3737,In_631,In_4129);
and U3738 (N_3738,In_1188,In_3798);
nor U3739 (N_3739,In_951,In_3516);
nand U3740 (N_3740,In_1795,In_3742);
or U3741 (N_3741,In_3388,In_4142);
xnor U3742 (N_3742,In_4540,In_289);
and U3743 (N_3743,In_2658,In_575);
xor U3744 (N_3744,In_891,In_569);
nor U3745 (N_3745,In_2310,In_702);
nor U3746 (N_3746,In_4522,In_1947);
nand U3747 (N_3747,In_2919,In_4166);
nand U3748 (N_3748,In_2355,In_3415);
nand U3749 (N_3749,In_2757,In_4998);
nor U3750 (N_3750,In_1831,In_3588);
xnor U3751 (N_3751,In_2342,In_1456);
nor U3752 (N_3752,In_421,In_1387);
or U3753 (N_3753,In_188,In_604);
nand U3754 (N_3754,In_3070,In_1068);
or U3755 (N_3755,In_1765,In_2882);
nor U3756 (N_3756,In_3879,In_3126);
nand U3757 (N_3757,In_1556,In_4677);
or U3758 (N_3758,In_174,In_1354);
nand U3759 (N_3759,In_4036,In_715);
nand U3760 (N_3760,In_4178,In_382);
nor U3761 (N_3761,In_3766,In_2121);
and U3762 (N_3762,In_1393,In_1599);
or U3763 (N_3763,In_4685,In_205);
nor U3764 (N_3764,In_4698,In_2234);
nand U3765 (N_3765,In_2200,In_4832);
and U3766 (N_3766,In_2132,In_3389);
nand U3767 (N_3767,In_453,In_3453);
or U3768 (N_3768,In_3314,In_2229);
and U3769 (N_3769,In_1353,In_374);
and U3770 (N_3770,In_3394,In_4947);
or U3771 (N_3771,In_2972,In_3255);
nor U3772 (N_3772,In_3133,In_2963);
xnor U3773 (N_3773,In_3814,In_4437);
and U3774 (N_3774,In_4754,In_773);
nor U3775 (N_3775,In_688,In_364);
and U3776 (N_3776,In_4154,In_1323);
and U3777 (N_3777,In_3999,In_2405);
nor U3778 (N_3778,In_3529,In_46);
nor U3779 (N_3779,In_3547,In_2232);
nor U3780 (N_3780,In_3388,In_3179);
xor U3781 (N_3781,In_862,In_4209);
nand U3782 (N_3782,In_933,In_967);
xor U3783 (N_3783,In_444,In_300);
nor U3784 (N_3784,In_310,In_4040);
nand U3785 (N_3785,In_1317,In_1266);
xor U3786 (N_3786,In_231,In_2017);
xnor U3787 (N_3787,In_1023,In_2741);
nor U3788 (N_3788,In_3443,In_3893);
xor U3789 (N_3789,In_937,In_211);
nor U3790 (N_3790,In_1182,In_2583);
or U3791 (N_3791,In_2996,In_2245);
xor U3792 (N_3792,In_1761,In_2352);
or U3793 (N_3793,In_2801,In_1194);
xnor U3794 (N_3794,In_41,In_1253);
nor U3795 (N_3795,In_1068,In_2596);
xor U3796 (N_3796,In_1996,In_2232);
xnor U3797 (N_3797,In_2841,In_4912);
or U3798 (N_3798,In_1732,In_2244);
nor U3799 (N_3799,In_3257,In_1183);
xor U3800 (N_3800,In_444,In_165);
xnor U3801 (N_3801,In_1371,In_1273);
nor U3802 (N_3802,In_2396,In_2346);
and U3803 (N_3803,In_1242,In_1653);
and U3804 (N_3804,In_2582,In_4736);
nand U3805 (N_3805,In_2056,In_1168);
nand U3806 (N_3806,In_3766,In_3874);
nand U3807 (N_3807,In_1465,In_1434);
nand U3808 (N_3808,In_863,In_3920);
or U3809 (N_3809,In_4555,In_2501);
nor U3810 (N_3810,In_4843,In_1094);
nor U3811 (N_3811,In_2308,In_2179);
xnor U3812 (N_3812,In_2491,In_4573);
nor U3813 (N_3813,In_1805,In_3418);
and U3814 (N_3814,In_1434,In_4585);
nor U3815 (N_3815,In_1290,In_1596);
or U3816 (N_3816,In_4119,In_2618);
nor U3817 (N_3817,In_2871,In_2701);
nor U3818 (N_3818,In_2662,In_412);
nor U3819 (N_3819,In_1465,In_530);
nand U3820 (N_3820,In_4490,In_2301);
nand U3821 (N_3821,In_840,In_1713);
nand U3822 (N_3822,In_3937,In_3099);
or U3823 (N_3823,In_2188,In_4851);
or U3824 (N_3824,In_3696,In_4078);
xnor U3825 (N_3825,In_2372,In_1810);
or U3826 (N_3826,In_857,In_1159);
nand U3827 (N_3827,In_1351,In_3939);
and U3828 (N_3828,In_3829,In_645);
nand U3829 (N_3829,In_1588,In_1519);
and U3830 (N_3830,In_2037,In_2280);
or U3831 (N_3831,In_2556,In_4777);
nor U3832 (N_3832,In_1809,In_1083);
or U3833 (N_3833,In_543,In_4851);
or U3834 (N_3834,In_2052,In_42);
nor U3835 (N_3835,In_2925,In_2891);
nor U3836 (N_3836,In_3035,In_557);
xor U3837 (N_3837,In_4245,In_3278);
nor U3838 (N_3838,In_2649,In_1846);
and U3839 (N_3839,In_346,In_4965);
nor U3840 (N_3840,In_3124,In_2124);
nand U3841 (N_3841,In_1544,In_3519);
and U3842 (N_3842,In_2402,In_3074);
or U3843 (N_3843,In_1644,In_193);
or U3844 (N_3844,In_3592,In_2929);
nand U3845 (N_3845,In_3008,In_4246);
nand U3846 (N_3846,In_880,In_1331);
xor U3847 (N_3847,In_3764,In_3065);
or U3848 (N_3848,In_4653,In_2118);
or U3849 (N_3849,In_2157,In_2519);
or U3850 (N_3850,In_2259,In_1059);
nand U3851 (N_3851,In_1757,In_329);
or U3852 (N_3852,In_2405,In_2576);
xnor U3853 (N_3853,In_4392,In_1068);
xnor U3854 (N_3854,In_4060,In_2984);
nor U3855 (N_3855,In_2279,In_4100);
or U3856 (N_3856,In_573,In_4045);
nand U3857 (N_3857,In_3453,In_3578);
nor U3858 (N_3858,In_719,In_3561);
nand U3859 (N_3859,In_3418,In_1048);
xnor U3860 (N_3860,In_4956,In_1269);
and U3861 (N_3861,In_996,In_3029);
nand U3862 (N_3862,In_3960,In_2103);
or U3863 (N_3863,In_43,In_4712);
nand U3864 (N_3864,In_4103,In_884);
xor U3865 (N_3865,In_4285,In_884);
or U3866 (N_3866,In_424,In_3069);
nand U3867 (N_3867,In_898,In_1726);
nand U3868 (N_3868,In_1249,In_2354);
and U3869 (N_3869,In_231,In_2494);
and U3870 (N_3870,In_4957,In_1753);
xor U3871 (N_3871,In_4014,In_1894);
and U3872 (N_3872,In_4599,In_1692);
or U3873 (N_3873,In_222,In_729);
and U3874 (N_3874,In_1024,In_3138);
or U3875 (N_3875,In_784,In_3663);
or U3876 (N_3876,In_2904,In_2175);
or U3877 (N_3877,In_4899,In_4029);
nand U3878 (N_3878,In_1637,In_3984);
xnor U3879 (N_3879,In_51,In_4685);
or U3880 (N_3880,In_2168,In_3484);
and U3881 (N_3881,In_2626,In_2587);
and U3882 (N_3882,In_90,In_1699);
nand U3883 (N_3883,In_3202,In_2407);
xnor U3884 (N_3884,In_159,In_4308);
nand U3885 (N_3885,In_1687,In_363);
xnor U3886 (N_3886,In_1386,In_109);
xor U3887 (N_3887,In_2646,In_254);
xnor U3888 (N_3888,In_3427,In_1673);
xor U3889 (N_3889,In_1190,In_2150);
nand U3890 (N_3890,In_2380,In_850);
nor U3891 (N_3891,In_3039,In_3104);
xnor U3892 (N_3892,In_3474,In_1243);
nand U3893 (N_3893,In_1016,In_1679);
and U3894 (N_3894,In_4564,In_3120);
or U3895 (N_3895,In_4246,In_1362);
nor U3896 (N_3896,In_4110,In_2321);
nor U3897 (N_3897,In_4634,In_3382);
nor U3898 (N_3898,In_2015,In_4701);
xor U3899 (N_3899,In_4568,In_1139);
nand U3900 (N_3900,In_1063,In_779);
and U3901 (N_3901,In_2807,In_1852);
nand U3902 (N_3902,In_1326,In_2404);
or U3903 (N_3903,In_2891,In_3743);
nor U3904 (N_3904,In_3618,In_3961);
and U3905 (N_3905,In_1445,In_3482);
nor U3906 (N_3906,In_4086,In_817);
nor U3907 (N_3907,In_4968,In_448);
nand U3908 (N_3908,In_190,In_2499);
or U3909 (N_3909,In_2609,In_4972);
nand U3910 (N_3910,In_4822,In_943);
xor U3911 (N_3911,In_3701,In_4678);
nor U3912 (N_3912,In_1758,In_797);
and U3913 (N_3913,In_4360,In_1602);
nand U3914 (N_3914,In_1881,In_4531);
nand U3915 (N_3915,In_1437,In_2758);
nor U3916 (N_3916,In_3211,In_191);
and U3917 (N_3917,In_4163,In_2942);
and U3918 (N_3918,In_2754,In_3054);
nand U3919 (N_3919,In_684,In_2258);
nand U3920 (N_3920,In_4433,In_4157);
xnor U3921 (N_3921,In_1429,In_4158);
nand U3922 (N_3922,In_4202,In_1654);
or U3923 (N_3923,In_4111,In_3413);
xor U3924 (N_3924,In_1256,In_3486);
xor U3925 (N_3925,In_3065,In_2022);
or U3926 (N_3926,In_2083,In_2220);
and U3927 (N_3927,In_3363,In_2536);
xor U3928 (N_3928,In_181,In_1797);
and U3929 (N_3929,In_384,In_2882);
or U3930 (N_3930,In_2032,In_1677);
and U3931 (N_3931,In_3135,In_2015);
and U3932 (N_3932,In_1852,In_1868);
or U3933 (N_3933,In_2274,In_2183);
nor U3934 (N_3934,In_4510,In_3986);
nand U3935 (N_3935,In_3194,In_1352);
xnor U3936 (N_3936,In_4483,In_4314);
nand U3937 (N_3937,In_63,In_3554);
nand U3938 (N_3938,In_1763,In_524);
and U3939 (N_3939,In_2722,In_3712);
nand U3940 (N_3940,In_4505,In_4171);
nor U3941 (N_3941,In_4567,In_3065);
and U3942 (N_3942,In_1802,In_4071);
and U3943 (N_3943,In_3892,In_178);
xor U3944 (N_3944,In_2297,In_1127);
or U3945 (N_3945,In_4716,In_4928);
nor U3946 (N_3946,In_4235,In_3179);
xnor U3947 (N_3947,In_937,In_254);
or U3948 (N_3948,In_4771,In_830);
xnor U3949 (N_3949,In_1670,In_1480);
and U3950 (N_3950,In_1612,In_3511);
nor U3951 (N_3951,In_4232,In_1770);
xor U3952 (N_3952,In_2681,In_2112);
xnor U3953 (N_3953,In_104,In_3145);
or U3954 (N_3954,In_1124,In_4657);
or U3955 (N_3955,In_2197,In_934);
nand U3956 (N_3956,In_1513,In_1707);
and U3957 (N_3957,In_2029,In_3502);
and U3958 (N_3958,In_3511,In_2220);
nand U3959 (N_3959,In_3595,In_3312);
xnor U3960 (N_3960,In_2909,In_2362);
and U3961 (N_3961,In_3480,In_76);
or U3962 (N_3962,In_4258,In_599);
nor U3963 (N_3963,In_4236,In_4708);
xor U3964 (N_3964,In_1907,In_2759);
and U3965 (N_3965,In_1110,In_3139);
nor U3966 (N_3966,In_401,In_4069);
and U3967 (N_3967,In_4027,In_4675);
or U3968 (N_3968,In_3925,In_4835);
and U3969 (N_3969,In_3587,In_1506);
nand U3970 (N_3970,In_1302,In_951);
or U3971 (N_3971,In_4199,In_2325);
or U3972 (N_3972,In_4404,In_1342);
xor U3973 (N_3973,In_438,In_4582);
nand U3974 (N_3974,In_4383,In_4614);
or U3975 (N_3975,In_2387,In_1685);
nand U3976 (N_3976,In_4688,In_2843);
and U3977 (N_3977,In_4153,In_2730);
xor U3978 (N_3978,In_2535,In_916);
nand U3979 (N_3979,In_2253,In_411);
nand U3980 (N_3980,In_654,In_4341);
and U3981 (N_3981,In_3936,In_2141);
xor U3982 (N_3982,In_3455,In_713);
and U3983 (N_3983,In_2050,In_3575);
or U3984 (N_3984,In_777,In_3236);
xor U3985 (N_3985,In_4235,In_4601);
xor U3986 (N_3986,In_2146,In_1857);
nor U3987 (N_3987,In_920,In_2354);
nor U3988 (N_3988,In_2267,In_3168);
xor U3989 (N_3989,In_1756,In_4198);
and U3990 (N_3990,In_914,In_3432);
nor U3991 (N_3991,In_1303,In_4199);
and U3992 (N_3992,In_3131,In_817);
and U3993 (N_3993,In_2850,In_3252);
nand U3994 (N_3994,In_4973,In_1053);
or U3995 (N_3995,In_4219,In_2145);
or U3996 (N_3996,In_2044,In_853);
nor U3997 (N_3997,In_509,In_304);
xnor U3998 (N_3998,In_510,In_2505);
or U3999 (N_3999,In_3589,In_2804);
nor U4000 (N_4000,In_2237,In_1448);
nor U4001 (N_4001,In_939,In_2100);
and U4002 (N_4002,In_1984,In_2569);
and U4003 (N_4003,In_1970,In_3449);
and U4004 (N_4004,In_4379,In_2105);
nor U4005 (N_4005,In_4235,In_558);
xnor U4006 (N_4006,In_170,In_2251);
or U4007 (N_4007,In_4418,In_336);
and U4008 (N_4008,In_1589,In_3117);
xnor U4009 (N_4009,In_2966,In_4139);
xnor U4010 (N_4010,In_4738,In_4714);
nor U4011 (N_4011,In_3891,In_4693);
xor U4012 (N_4012,In_4524,In_101);
nand U4013 (N_4013,In_4108,In_4956);
xnor U4014 (N_4014,In_344,In_389);
xnor U4015 (N_4015,In_2955,In_4287);
nand U4016 (N_4016,In_126,In_2495);
and U4017 (N_4017,In_4055,In_2251);
nor U4018 (N_4018,In_1996,In_2629);
or U4019 (N_4019,In_4231,In_311);
nand U4020 (N_4020,In_3409,In_1337);
nor U4021 (N_4021,In_946,In_3573);
and U4022 (N_4022,In_4194,In_3084);
and U4023 (N_4023,In_182,In_4977);
or U4024 (N_4024,In_2083,In_4234);
or U4025 (N_4025,In_1581,In_2249);
nor U4026 (N_4026,In_4259,In_2980);
nand U4027 (N_4027,In_1160,In_2908);
nor U4028 (N_4028,In_2718,In_4002);
xor U4029 (N_4029,In_1327,In_2943);
nor U4030 (N_4030,In_1291,In_1208);
nand U4031 (N_4031,In_3164,In_1939);
nand U4032 (N_4032,In_4387,In_3543);
nand U4033 (N_4033,In_1779,In_1925);
nand U4034 (N_4034,In_4715,In_3625);
nand U4035 (N_4035,In_3873,In_837);
and U4036 (N_4036,In_3081,In_1746);
nand U4037 (N_4037,In_100,In_4062);
xor U4038 (N_4038,In_4649,In_233);
and U4039 (N_4039,In_364,In_4918);
or U4040 (N_4040,In_610,In_4728);
xnor U4041 (N_4041,In_3685,In_589);
xnor U4042 (N_4042,In_3239,In_16);
and U4043 (N_4043,In_580,In_3245);
and U4044 (N_4044,In_4633,In_3792);
xnor U4045 (N_4045,In_1299,In_1230);
nand U4046 (N_4046,In_4165,In_156);
and U4047 (N_4047,In_2163,In_1850);
and U4048 (N_4048,In_4338,In_1671);
and U4049 (N_4049,In_118,In_1145);
nand U4050 (N_4050,In_3158,In_4711);
xnor U4051 (N_4051,In_113,In_458);
nand U4052 (N_4052,In_4221,In_3356);
nor U4053 (N_4053,In_3100,In_2514);
nand U4054 (N_4054,In_2863,In_905);
or U4055 (N_4055,In_2018,In_4017);
or U4056 (N_4056,In_852,In_3950);
nor U4057 (N_4057,In_2311,In_3768);
and U4058 (N_4058,In_1528,In_4159);
or U4059 (N_4059,In_1592,In_3025);
and U4060 (N_4060,In_3963,In_782);
xor U4061 (N_4061,In_2440,In_4118);
nand U4062 (N_4062,In_368,In_1545);
or U4063 (N_4063,In_3011,In_1148);
or U4064 (N_4064,In_3200,In_945);
xor U4065 (N_4065,In_4443,In_2203);
nor U4066 (N_4066,In_2775,In_559);
nor U4067 (N_4067,In_1771,In_4170);
or U4068 (N_4068,In_3396,In_268);
and U4069 (N_4069,In_468,In_4408);
and U4070 (N_4070,In_113,In_1137);
or U4071 (N_4071,In_3292,In_127);
or U4072 (N_4072,In_4352,In_4869);
nor U4073 (N_4073,In_2088,In_1071);
and U4074 (N_4074,In_3092,In_2477);
xnor U4075 (N_4075,In_902,In_1159);
or U4076 (N_4076,In_4166,In_3256);
nand U4077 (N_4077,In_534,In_3234);
nand U4078 (N_4078,In_1746,In_2187);
xor U4079 (N_4079,In_1476,In_705);
xor U4080 (N_4080,In_3710,In_3390);
nor U4081 (N_4081,In_1920,In_2013);
xnor U4082 (N_4082,In_1717,In_1038);
nor U4083 (N_4083,In_3380,In_1787);
xor U4084 (N_4084,In_1849,In_2510);
and U4085 (N_4085,In_3674,In_3096);
xnor U4086 (N_4086,In_4759,In_3822);
nor U4087 (N_4087,In_1055,In_976);
nor U4088 (N_4088,In_3858,In_969);
nor U4089 (N_4089,In_1037,In_1118);
nor U4090 (N_4090,In_1860,In_2495);
nand U4091 (N_4091,In_3979,In_4967);
nor U4092 (N_4092,In_1338,In_4674);
nor U4093 (N_4093,In_1886,In_2958);
and U4094 (N_4094,In_4968,In_363);
nor U4095 (N_4095,In_1388,In_1990);
or U4096 (N_4096,In_2811,In_3325);
xnor U4097 (N_4097,In_2192,In_2231);
or U4098 (N_4098,In_4867,In_4990);
xnor U4099 (N_4099,In_917,In_2873);
nand U4100 (N_4100,In_3036,In_1800);
nor U4101 (N_4101,In_1788,In_4075);
and U4102 (N_4102,In_1398,In_3687);
nor U4103 (N_4103,In_4533,In_79);
or U4104 (N_4104,In_3791,In_4351);
or U4105 (N_4105,In_861,In_2289);
nand U4106 (N_4106,In_2062,In_3505);
nor U4107 (N_4107,In_2172,In_1781);
nand U4108 (N_4108,In_4503,In_3233);
xor U4109 (N_4109,In_4487,In_4476);
nor U4110 (N_4110,In_1464,In_4257);
xor U4111 (N_4111,In_3522,In_4647);
and U4112 (N_4112,In_3727,In_3762);
nand U4113 (N_4113,In_4422,In_27);
and U4114 (N_4114,In_3233,In_89);
and U4115 (N_4115,In_3768,In_4277);
and U4116 (N_4116,In_4227,In_2318);
nor U4117 (N_4117,In_1454,In_181);
nand U4118 (N_4118,In_3263,In_3762);
nand U4119 (N_4119,In_2649,In_2272);
nor U4120 (N_4120,In_3712,In_3852);
and U4121 (N_4121,In_4629,In_637);
nor U4122 (N_4122,In_1726,In_3689);
nand U4123 (N_4123,In_4606,In_2733);
xnor U4124 (N_4124,In_71,In_2452);
and U4125 (N_4125,In_2228,In_1038);
or U4126 (N_4126,In_3598,In_131);
nand U4127 (N_4127,In_1853,In_3359);
nand U4128 (N_4128,In_4998,In_4010);
xnor U4129 (N_4129,In_3873,In_4213);
nand U4130 (N_4130,In_4016,In_2929);
or U4131 (N_4131,In_1980,In_3838);
or U4132 (N_4132,In_4355,In_118);
xnor U4133 (N_4133,In_3036,In_275);
nor U4134 (N_4134,In_3325,In_2546);
and U4135 (N_4135,In_2928,In_952);
xnor U4136 (N_4136,In_2873,In_4044);
or U4137 (N_4137,In_1461,In_1365);
nand U4138 (N_4138,In_3525,In_4523);
nor U4139 (N_4139,In_3532,In_2310);
nor U4140 (N_4140,In_79,In_3315);
and U4141 (N_4141,In_955,In_126);
nor U4142 (N_4142,In_2971,In_4208);
nand U4143 (N_4143,In_3882,In_903);
and U4144 (N_4144,In_4473,In_2804);
and U4145 (N_4145,In_1261,In_1612);
nor U4146 (N_4146,In_1869,In_355);
xnor U4147 (N_4147,In_585,In_354);
or U4148 (N_4148,In_3843,In_1260);
or U4149 (N_4149,In_1358,In_1472);
nand U4150 (N_4150,In_2202,In_3262);
or U4151 (N_4151,In_4048,In_2411);
xor U4152 (N_4152,In_203,In_4143);
nor U4153 (N_4153,In_4224,In_3318);
and U4154 (N_4154,In_3456,In_3020);
and U4155 (N_4155,In_9,In_3014);
nand U4156 (N_4156,In_3964,In_4380);
xnor U4157 (N_4157,In_4102,In_104);
nor U4158 (N_4158,In_412,In_3128);
xnor U4159 (N_4159,In_381,In_1917);
xor U4160 (N_4160,In_3678,In_3535);
nor U4161 (N_4161,In_1701,In_1651);
or U4162 (N_4162,In_3944,In_2109);
or U4163 (N_4163,In_131,In_1665);
xor U4164 (N_4164,In_370,In_40);
nand U4165 (N_4165,In_2977,In_1833);
xor U4166 (N_4166,In_2571,In_4565);
nor U4167 (N_4167,In_2394,In_773);
xnor U4168 (N_4168,In_2888,In_1457);
or U4169 (N_4169,In_3568,In_2822);
nand U4170 (N_4170,In_2764,In_4839);
nor U4171 (N_4171,In_3944,In_4572);
xnor U4172 (N_4172,In_4207,In_136);
xnor U4173 (N_4173,In_3421,In_2735);
xor U4174 (N_4174,In_1797,In_4259);
xnor U4175 (N_4175,In_1672,In_3567);
or U4176 (N_4176,In_3798,In_2062);
nand U4177 (N_4177,In_215,In_607);
nand U4178 (N_4178,In_1478,In_4426);
and U4179 (N_4179,In_335,In_1971);
nand U4180 (N_4180,In_315,In_3579);
nor U4181 (N_4181,In_1550,In_1159);
nand U4182 (N_4182,In_1018,In_4849);
or U4183 (N_4183,In_2445,In_310);
and U4184 (N_4184,In_3324,In_1650);
or U4185 (N_4185,In_2346,In_2991);
or U4186 (N_4186,In_4275,In_4685);
nand U4187 (N_4187,In_4272,In_4522);
nor U4188 (N_4188,In_1088,In_2144);
or U4189 (N_4189,In_2042,In_1775);
or U4190 (N_4190,In_3584,In_2403);
nor U4191 (N_4191,In_2797,In_3032);
nand U4192 (N_4192,In_38,In_1631);
xor U4193 (N_4193,In_4240,In_1924);
xor U4194 (N_4194,In_4688,In_4237);
nand U4195 (N_4195,In_504,In_898);
xnor U4196 (N_4196,In_1028,In_3264);
or U4197 (N_4197,In_4100,In_3113);
nor U4198 (N_4198,In_3993,In_315);
nand U4199 (N_4199,In_2817,In_2846);
or U4200 (N_4200,In_4236,In_4234);
or U4201 (N_4201,In_4681,In_2586);
nor U4202 (N_4202,In_3781,In_3492);
nand U4203 (N_4203,In_2447,In_555);
xor U4204 (N_4204,In_2975,In_4959);
nor U4205 (N_4205,In_1762,In_3243);
xnor U4206 (N_4206,In_5,In_3681);
or U4207 (N_4207,In_286,In_3244);
or U4208 (N_4208,In_1716,In_1415);
nand U4209 (N_4209,In_905,In_1258);
or U4210 (N_4210,In_2699,In_3349);
nand U4211 (N_4211,In_4017,In_2695);
nor U4212 (N_4212,In_3908,In_4845);
nor U4213 (N_4213,In_1813,In_1372);
nand U4214 (N_4214,In_812,In_3898);
or U4215 (N_4215,In_3983,In_395);
xor U4216 (N_4216,In_2589,In_3818);
or U4217 (N_4217,In_513,In_3779);
or U4218 (N_4218,In_177,In_1979);
nor U4219 (N_4219,In_726,In_3154);
or U4220 (N_4220,In_2012,In_1033);
or U4221 (N_4221,In_1698,In_1890);
nand U4222 (N_4222,In_49,In_4244);
or U4223 (N_4223,In_3862,In_1075);
xor U4224 (N_4224,In_90,In_2082);
nand U4225 (N_4225,In_4152,In_2173);
nor U4226 (N_4226,In_3941,In_1435);
or U4227 (N_4227,In_2162,In_992);
or U4228 (N_4228,In_583,In_4198);
nand U4229 (N_4229,In_1528,In_376);
or U4230 (N_4230,In_3866,In_4757);
nand U4231 (N_4231,In_4759,In_4412);
or U4232 (N_4232,In_3455,In_207);
or U4233 (N_4233,In_596,In_1575);
nand U4234 (N_4234,In_428,In_3769);
and U4235 (N_4235,In_2749,In_394);
or U4236 (N_4236,In_617,In_4360);
nor U4237 (N_4237,In_4895,In_2895);
and U4238 (N_4238,In_3245,In_774);
and U4239 (N_4239,In_3135,In_619);
and U4240 (N_4240,In_3549,In_2826);
nor U4241 (N_4241,In_2273,In_219);
and U4242 (N_4242,In_4155,In_2583);
nand U4243 (N_4243,In_4987,In_1334);
or U4244 (N_4244,In_3884,In_622);
nand U4245 (N_4245,In_1952,In_2438);
xnor U4246 (N_4246,In_3809,In_438);
nand U4247 (N_4247,In_411,In_2859);
nand U4248 (N_4248,In_1740,In_226);
nor U4249 (N_4249,In_2398,In_1490);
nand U4250 (N_4250,In_3170,In_1756);
or U4251 (N_4251,In_3263,In_661);
nand U4252 (N_4252,In_4641,In_11);
xnor U4253 (N_4253,In_2329,In_3084);
xnor U4254 (N_4254,In_2912,In_36);
and U4255 (N_4255,In_4990,In_2021);
xnor U4256 (N_4256,In_141,In_3120);
nand U4257 (N_4257,In_4295,In_2663);
nor U4258 (N_4258,In_4317,In_3130);
nor U4259 (N_4259,In_865,In_4309);
nor U4260 (N_4260,In_3568,In_1117);
xnor U4261 (N_4261,In_1435,In_4758);
xor U4262 (N_4262,In_1092,In_4314);
nor U4263 (N_4263,In_864,In_1171);
nor U4264 (N_4264,In_2185,In_4860);
or U4265 (N_4265,In_4927,In_3174);
and U4266 (N_4266,In_682,In_4952);
xnor U4267 (N_4267,In_4400,In_4553);
and U4268 (N_4268,In_1199,In_4102);
xnor U4269 (N_4269,In_390,In_2665);
nand U4270 (N_4270,In_271,In_629);
nand U4271 (N_4271,In_3255,In_2795);
nand U4272 (N_4272,In_3199,In_1703);
nor U4273 (N_4273,In_2800,In_2330);
nor U4274 (N_4274,In_3615,In_2976);
and U4275 (N_4275,In_1197,In_3664);
xnor U4276 (N_4276,In_1868,In_929);
and U4277 (N_4277,In_2803,In_4649);
nand U4278 (N_4278,In_529,In_1774);
nand U4279 (N_4279,In_4402,In_4240);
and U4280 (N_4280,In_1822,In_1821);
nor U4281 (N_4281,In_3979,In_2353);
xor U4282 (N_4282,In_4968,In_218);
xor U4283 (N_4283,In_3278,In_4583);
nand U4284 (N_4284,In_267,In_4545);
nand U4285 (N_4285,In_1039,In_2048);
nand U4286 (N_4286,In_1222,In_4047);
or U4287 (N_4287,In_2550,In_2374);
nand U4288 (N_4288,In_1540,In_2779);
xnor U4289 (N_4289,In_2539,In_2204);
nor U4290 (N_4290,In_2954,In_1178);
and U4291 (N_4291,In_83,In_3596);
nor U4292 (N_4292,In_2716,In_3227);
xnor U4293 (N_4293,In_696,In_114);
xor U4294 (N_4294,In_3170,In_865);
and U4295 (N_4295,In_2218,In_4624);
nor U4296 (N_4296,In_4633,In_1735);
and U4297 (N_4297,In_4952,In_2203);
nand U4298 (N_4298,In_1629,In_2733);
nor U4299 (N_4299,In_992,In_642);
nor U4300 (N_4300,In_3264,In_177);
and U4301 (N_4301,In_3390,In_3775);
nand U4302 (N_4302,In_3860,In_3939);
nor U4303 (N_4303,In_780,In_3028);
xnor U4304 (N_4304,In_1724,In_137);
xor U4305 (N_4305,In_4950,In_3690);
and U4306 (N_4306,In_1703,In_1287);
or U4307 (N_4307,In_1327,In_4588);
and U4308 (N_4308,In_4515,In_120);
nand U4309 (N_4309,In_3729,In_3828);
nand U4310 (N_4310,In_3686,In_994);
xor U4311 (N_4311,In_300,In_1623);
nand U4312 (N_4312,In_1788,In_4296);
nor U4313 (N_4313,In_4214,In_1250);
or U4314 (N_4314,In_2410,In_276);
and U4315 (N_4315,In_2,In_1626);
xor U4316 (N_4316,In_2357,In_4203);
xnor U4317 (N_4317,In_883,In_3626);
or U4318 (N_4318,In_42,In_845);
nand U4319 (N_4319,In_1329,In_308);
xor U4320 (N_4320,In_3859,In_1795);
or U4321 (N_4321,In_289,In_3599);
and U4322 (N_4322,In_4353,In_1078);
nand U4323 (N_4323,In_4739,In_4592);
or U4324 (N_4324,In_2428,In_1031);
or U4325 (N_4325,In_2160,In_2109);
or U4326 (N_4326,In_531,In_2815);
nand U4327 (N_4327,In_1924,In_4175);
xnor U4328 (N_4328,In_2554,In_2950);
nor U4329 (N_4329,In_1443,In_2406);
and U4330 (N_4330,In_3615,In_245);
or U4331 (N_4331,In_3762,In_852);
or U4332 (N_4332,In_4071,In_1834);
or U4333 (N_4333,In_3943,In_504);
nor U4334 (N_4334,In_4550,In_3847);
or U4335 (N_4335,In_439,In_3615);
and U4336 (N_4336,In_3980,In_1048);
xnor U4337 (N_4337,In_3821,In_1250);
nor U4338 (N_4338,In_225,In_2989);
xnor U4339 (N_4339,In_3238,In_4401);
and U4340 (N_4340,In_4700,In_3947);
nor U4341 (N_4341,In_4146,In_2752);
nor U4342 (N_4342,In_1552,In_1934);
or U4343 (N_4343,In_1760,In_3147);
nor U4344 (N_4344,In_1754,In_1229);
and U4345 (N_4345,In_4922,In_1521);
xnor U4346 (N_4346,In_2124,In_3422);
nor U4347 (N_4347,In_2828,In_2371);
nor U4348 (N_4348,In_1740,In_1492);
or U4349 (N_4349,In_1686,In_3751);
xnor U4350 (N_4350,In_1968,In_1182);
and U4351 (N_4351,In_2962,In_2353);
xor U4352 (N_4352,In_3854,In_1478);
xor U4353 (N_4353,In_1408,In_3985);
or U4354 (N_4354,In_3096,In_120);
xor U4355 (N_4355,In_205,In_732);
nor U4356 (N_4356,In_556,In_652);
and U4357 (N_4357,In_4916,In_192);
nand U4358 (N_4358,In_3101,In_2995);
and U4359 (N_4359,In_3396,In_728);
nor U4360 (N_4360,In_3519,In_492);
nor U4361 (N_4361,In_3859,In_1456);
or U4362 (N_4362,In_1518,In_1418);
xnor U4363 (N_4363,In_3327,In_1816);
xnor U4364 (N_4364,In_4718,In_3485);
or U4365 (N_4365,In_2771,In_4356);
nor U4366 (N_4366,In_1923,In_3978);
and U4367 (N_4367,In_4091,In_2787);
and U4368 (N_4368,In_3981,In_4682);
or U4369 (N_4369,In_2130,In_3775);
nor U4370 (N_4370,In_3578,In_3240);
or U4371 (N_4371,In_2336,In_131);
and U4372 (N_4372,In_1039,In_190);
nand U4373 (N_4373,In_992,In_30);
nand U4374 (N_4374,In_93,In_376);
and U4375 (N_4375,In_4351,In_2685);
or U4376 (N_4376,In_2867,In_4497);
and U4377 (N_4377,In_2551,In_4551);
and U4378 (N_4378,In_4892,In_1848);
and U4379 (N_4379,In_4335,In_455);
or U4380 (N_4380,In_1820,In_4305);
or U4381 (N_4381,In_4631,In_43);
xnor U4382 (N_4382,In_2305,In_2052);
xor U4383 (N_4383,In_4509,In_1898);
and U4384 (N_4384,In_2497,In_4351);
xor U4385 (N_4385,In_3382,In_2279);
or U4386 (N_4386,In_4315,In_44);
nor U4387 (N_4387,In_2705,In_4378);
and U4388 (N_4388,In_1125,In_2286);
nor U4389 (N_4389,In_2994,In_3459);
and U4390 (N_4390,In_1588,In_1521);
and U4391 (N_4391,In_2650,In_89);
nor U4392 (N_4392,In_3163,In_1620);
nor U4393 (N_4393,In_3038,In_4167);
and U4394 (N_4394,In_2181,In_4500);
or U4395 (N_4395,In_4084,In_3979);
nand U4396 (N_4396,In_2504,In_514);
or U4397 (N_4397,In_881,In_2869);
nor U4398 (N_4398,In_4664,In_754);
nor U4399 (N_4399,In_2666,In_1442);
or U4400 (N_4400,In_4386,In_122);
nor U4401 (N_4401,In_1831,In_3088);
or U4402 (N_4402,In_3761,In_4834);
nand U4403 (N_4403,In_1085,In_486);
and U4404 (N_4404,In_3025,In_3076);
and U4405 (N_4405,In_826,In_2980);
nand U4406 (N_4406,In_3410,In_1137);
nor U4407 (N_4407,In_512,In_3191);
nor U4408 (N_4408,In_4303,In_463);
xor U4409 (N_4409,In_2938,In_1967);
and U4410 (N_4410,In_1884,In_3780);
xnor U4411 (N_4411,In_4016,In_3600);
nand U4412 (N_4412,In_327,In_3236);
nor U4413 (N_4413,In_4883,In_2962);
xnor U4414 (N_4414,In_1161,In_1745);
and U4415 (N_4415,In_1985,In_3848);
nor U4416 (N_4416,In_1076,In_1754);
nand U4417 (N_4417,In_2707,In_2086);
nor U4418 (N_4418,In_270,In_4702);
nor U4419 (N_4419,In_4792,In_280);
and U4420 (N_4420,In_2627,In_1896);
nand U4421 (N_4421,In_3591,In_152);
xnor U4422 (N_4422,In_2287,In_653);
nand U4423 (N_4423,In_4738,In_3033);
nand U4424 (N_4424,In_2657,In_1419);
nand U4425 (N_4425,In_2886,In_3471);
nand U4426 (N_4426,In_2807,In_1591);
and U4427 (N_4427,In_1063,In_1927);
nor U4428 (N_4428,In_2878,In_4176);
nor U4429 (N_4429,In_3093,In_4274);
and U4430 (N_4430,In_1091,In_4570);
or U4431 (N_4431,In_3115,In_533);
or U4432 (N_4432,In_1335,In_858);
and U4433 (N_4433,In_3651,In_1573);
nand U4434 (N_4434,In_3625,In_121);
or U4435 (N_4435,In_1277,In_1698);
nor U4436 (N_4436,In_1832,In_1402);
or U4437 (N_4437,In_4547,In_1992);
nand U4438 (N_4438,In_3069,In_4541);
or U4439 (N_4439,In_427,In_4022);
nand U4440 (N_4440,In_475,In_963);
or U4441 (N_4441,In_1325,In_2133);
xor U4442 (N_4442,In_4754,In_2920);
xnor U4443 (N_4443,In_1017,In_3319);
xnor U4444 (N_4444,In_4135,In_4814);
xor U4445 (N_4445,In_619,In_894);
and U4446 (N_4446,In_3507,In_3349);
nand U4447 (N_4447,In_1170,In_1238);
nand U4448 (N_4448,In_276,In_193);
nor U4449 (N_4449,In_2292,In_4251);
or U4450 (N_4450,In_4711,In_2795);
and U4451 (N_4451,In_2148,In_1496);
xnor U4452 (N_4452,In_2122,In_2342);
xor U4453 (N_4453,In_2660,In_3733);
nor U4454 (N_4454,In_3847,In_4619);
nand U4455 (N_4455,In_2840,In_1974);
and U4456 (N_4456,In_979,In_3171);
and U4457 (N_4457,In_1190,In_2466);
xor U4458 (N_4458,In_2407,In_2437);
and U4459 (N_4459,In_4556,In_3984);
nor U4460 (N_4460,In_905,In_1494);
nor U4461 (N_4461,In_4981,In_1066);
and U4462 (N_4462,In_4337,In_3261);
or U4463 (N_4463,In_658,In_3530);
or U4464 (N_4464,In_2025,In_3036);
and U4465 (N_4465,In_276,In_2556);
and U4466 (N_4466,In_4620,In_2186);
or U4467 (N_4467,In_1048,In_422);
or U4468 (N_4468,In_1988,In_3191);
or U4469 (N_4469,In_2180,In_1808);
and U4470 (N_4470,In_2855,In_187);
nor U4471 (N_4471,In_21,In_4418);
nand U4472 (N_4472,In_2487,In_1106);
or U4473 (N_4473,In_4863,In_271);
xor U4474 (N_4474,In_2788,In_2772);
or U4475 (N_4475,In_1295,In_1714);
xor U4476 (N_4476,In_4789,In_428);
xnor U4477 (N_4477,In_3609,In_3382);
or U4478 (N_4478,In_2972,In_2872);
nand U4479 (N_4479,In_581,In_1878);
or U4480 (N_4480,In_4746,In_4781);
or U4481 (N_4481,In_3808,In_1395);
xor U4482 (N_4482,In_62,In_629);
nor U4483 (N_4483,In_4187,In_4125);
nor U4484 (N_4484,In_3039,In_3999);
nor U4485 (N_4485,In_4731,In_1278);
nor U4486 (N_4486,In_4242,In_447);
or U4487 (N_4487,In_3593,In_4779);
nand U4488 (N_4488,In_335,In_4383);
and U4489 (N_4489,In_3891,In_2237);
or U4490 (N_4490,In_4245,In_4816);
nor U4491 (N_4491,In_3959,In_2024);
or U4492 (N_4492,In_1868,In_1821);
nand U4493 (N_4493,In_4386,In_4898);
nand U4494 (N_4494,In_1153,In_2863);
and U4495 (N_4495,In_180,In_3396);
and U4496 (N_4496,In_4624,In_955);
or U4497 (N_4497,In_2070,In_125);
nand U4498 (N_4498,In_4109,In_2870);
xor U4499 (N_4499,In_2081,In_1209);
nand U4500 (N_4500,In_4005,In_3093);
and U4501 (N_4501,In_1805,In_3135);
nor U4502 (N_4502,In_1039,In_765);
xor U4503 (N_4503,In_864,In_4091);
or U4504 (N_4504,In_1222,In_4429);
and U4505 (N_4505,In_2104,In_3950);
nor U4506 (N_4506,In_4567,In_385);
nor U4507 (N_4507,In_4146,In_866);
and U4508 (N_4508,In_488,In_4406);
xor U4509 (N_4509,In_3724,In_2116);
nor U4510 (N_4510,In_3931,In_2065);
nand U4511 (N_4511,In_3639,In_4572);
nor U4512 (N_4512,In_1186,In_1219);
and U4513 (N_4513,In_622,In_1517);
or U4514 (N_4514,In_110,In_2357);
nor U4515 (N_4515,In_333,In_2272);
nand U4516 (N_4516,In_136,In_1071);
and U4517 (N_4517,In_986,In_4549);
and U4518 (N_4518,In_3917,In_1392);
nor U4519 (N_4519,In_2900,In_1207);
xnor U4520 (N_4520,In_2189,In_2208);
nand U4521 (N_4521,In_2198,In_3983);
and U4522 (N_4522,In_4196,In_1998);
or U4523 (N_4523,In_3130,In_981);
xor U4524 (N_4524,In_1498,In_2134);
nor U4525 (N_4525,In_1260,In_2304);
and U4526 (N_4526,In_1325,In_3508);
or U4527 (N_4527,In_3113,In_4136);
nand U4528 (N_4528,In_3262,In_2374);
nand U4529 (N_4529,In_850,In_4221);
nor U4530 (N_4530,In_303,In_3290);
nor U4531 (N_4531,In_1675,In_1777);
nand U4532 (N_4532,In_2669,In_4250);
nor U4533 (N_4533,In_270,In_2033);
xor U4534 (N_4534,In_738,In_3295);
xnor U4535 (N_4535,In_1122,In_1470);
nand U4536 (N_4536,In_1720,In_1711);
nor U4537 (N_4537,In_691,In_3816);
nor U4538 (N_4538,In_163,In_4288);
or U4539 (N_4539,In_4162,In_1561);
xnor U4540 (N_4540,In_1905,In_120);
and U4541 (N_4541,In_4744,In_756);
nand U4542 (N_4542,In_1967,In_154);
and U4543 (N_4543,In_68,In_151);
nor U4544 (N_4544,In_2020,In_1763);
and U4545 (N_4545,In_1653,In_2853);
or U4546 (N_4546,In_4710,In_3880);
xor U4547 (N_4547,In_2602,In_1105);
nor U4548 (N_4548,In_123,In_1783);
nand U4549 (N_4549,In_3462,In_2916);
nor U4550 (N_4550,In_3103,In_128);
and U4551 (N_4551,In_3174,In_3823);
nor U4552 (N_4552,In_479,In_4390);
nand U4553 (N_4553,In_2428,In_1967);
or U4554 (N_4554,In_2297,In_756);
nor U4555 (N_4555,In_391,In_2661);
nor U4556 (N_4556,In_4212,In_3844);
xor U4557 (N_4557,In_1751,In_4085);
xor U4558 (N_4558,In_3592,In_3119);
xor U4559 (N_4559,In_4534,In_1663);
xor U4560 (N_4560,In_4996,In_2832);
nor U4561 (N_4561,In_1189,In_3807);
nand U4562 (N_4562,In_30,In_2753);
and U4563 (N_4563,In_3515,In_1020);
nand U4564 (N_4564,In_4561,In_240);
nand U4565 (N_4565,In_265,In_3526);
or U4566 (N_4566,In_1516,In_3117);
and U4567 (N_4567,In_4582,In_3063);
xor U4568 (N_4568,In_1403,In_1062);
xnor U4569 (N_4569,In_3665,In_1048);
or U4570 (N_4570,In_2479,In_1083);
nand U4571 (N_4571,In_3509,In_1484);
or U4572 (N_4572,In_2674,In_1568);
nor U4573 (N_4573,In_176,In_1386);
nand U4574 (N_4574,In_2969,In_4603);
xor U4575 (N_4575,In_2500,In_978);
or U4576 (N_4576,In_3003,In_167);
and U4577 (N_4577,In_3195,In_487);
xnor U4578 (N_4578,In_3684,In_3463);
xor U4579 (N_4579,In_2452,In_4717);
and U4580 (N_4580,In_2619,In_4053);
nor U4581 (N_4581,In_2347,In_4727);
or U4582 (N_4582,In_1429,In_1973);
and U4583 (N_4583,In_1370,In_1342);
and U4584 (N_4584,In_2287,In_674);
nor U4585 (N_4585,In_1091,In_2452);
nand U4586 (N_4586,In_4965,In_4206);
nand U4587 (N_4587,In_1842,In_3718);
and U4588 (N_4588,In_787,In_1256);
or U4589 (N_4589,In_604,In_3567);
xor U4590 (N_4590,In_3076,In_996);
or U4591 (N_4591,In_22,In_1379);
nand U4592 (N_4592,In_2766,In_2142);
nand U4593 (N_4593,In_2660,In_1817);
xnor U4594 (N_4594,In_3933,In_67);
nand U4595 (N_4595,In_2081,In_12);
nand U4596 (N_4596,In_3476,In_4745);
xor U4597 (N_4597,In_1431,In_310);
nand U4598 (N_4598,In_1510,In_2243);
nand U4599 (N_4599,In_1167,In_457);
and U4600 (N_4600,In_2484,In_3854);
nor U4601 (N_4601,In_2600,In_2475);
and U4602 (N_4602,In_1364,In_2501);
nor U4603 (N_4603,In_1401,In_4019);
nand U4604 (N_4604,In_2240,In_3438);
nand U4605 (N_4605,In_4980,In_2522);
nor U4606 (N_4606,In_110,In_354);
nand U4607 (N_4607,In_3134,In_582);
and U4608 (N_4608,In_1193,In_2867);
and U4609 (N_4609,In_4105,In_1392);
xnor U4610 (N_4610,In_2100,In_2285);
and U4611 (N_4611,In_186,In_3273);
or U4612 (N_4612,In_4176,In_4875);
nor U4613 (N_4613,In_196,In_370);
nor U4614 (N_4614,In_3421,In_2752);
xnor U4615 (N_4615,In_4837,In_2706);
xor U4616 (N_4616,In_4798,In_2613);
and U4617 (N_4617,In_1045,In_3786);
nand U4618 (N_4618,In_3827,In_4148);
and U4619 (N_4619,In_2974,In_2294);
or U4620 (N_4620,In_2326,In_1818);
or U4621 (N_4621,In_4036,In_4083);
nor U4622 (N_4622,In_112,In_3986);
nor U4623 (N_4623,In_584,In_623);
nor U4624 (N_4624,In_4303,In_4305);
nor U4625 (N_4625,In_4906,In_1970);
xor U4626 (N_4626,In_152,In_1953);
or U4627 (N_4627,In_2401,In_1676);
and U4628 (N_4628,In_3989,In_2703);
nand U4629 (N_4629,In_4867,In_1522);
and U4630 (N_4630,In_3731,In_519);
nand U4631 (N_4631,In_4570,In_2021);
nand U4632 (N_4632,In_648,In_3614);
nor U4633 (N_4633,In_4160,In_704);
nand U4634 (N_4634,In_644,In_2042);
nand U4635 (N_4635,In_4,In_2586);
or U4636 (N_4636,In_2637,In_3302);
or U4637 (N_4637,In_1741,In_4168);
nand U4638 (N_4638,In_716,In_1105);
nor U4639 (N_4639,In_4904,In_1895);
nor U4640 (N_4640,In_4480,In_1110);
nand U4641 (N_4641,In_4695,In_1032);
xor U4642 (N_4642,In_4861,In_3266);
nand U4643 (N_4643,In_111,In_4907);
nor U4644 (N_4644,In_1594,In_3093);
or U4645 (N_4645,In_444,In_3303);
or U4646 (N_4646,In_2426,In_3610);
nor U4647 (N_4647,In_1352,In_3940);
nor U4648 (N_4648,In_2939,In_3614);
or U4649 (N_4649,In_4770,In_4726);
or U4650 (N_4650,In_4333,In_143);
or U4651 (N_4651,In_2389,In_3359);
or U4652 (N_4652,In_681,In_4109);
nand U4653 (N_4653,In_2523,In_2785);
and U4654 (N_4654,In_4263,In_3636);
nor U4655 (N_4655,In_4119,In_2242);
and U4656 (N_4656,In_2149,In_2203);
xor U4657 (N_4657,In_1941,In_3859);
nor U4658 (N_4658,In_1567,In_239);
nor U4659 (N_4659,In_2911,In_3367);
nand U4660 (N_4660,In_1855,In_2113);
nor U4661 (N_4661,In_273,In_112);
nor U4662 (N_4662,In_779,In_1869);
and U4663 (N_4663,In_3347,In_1784);
nor U4664 (N_4664,In_31,In_163);
xnor U4665 (N_4665,In_52,In_4755);
xnor U4666 (N_4666,In_2870,In_494);
and U4667 (N_4667,In_3799,In_1750);
nor U4668 (N_4668,In_227,In_974);
and U4669 (N_4669,In_789,In_2337);
nand U4670 (N_4670,In_4700,In_4474);
nor U4671 (N_4671,In_650,In_4228);
nand U4672 (N_4672,In_337,In_4106);
nor U4673 (N_4673,In_2753,In_2739);
xor U4674 (N_4674,In_2556,In_2803);
nand U4675 (N_4675,In_2668,In_2581);
xor U4676 (N_4676,In_2424,In_4781);
nor U4677 (N_4677,In_3450,In_2892);
nor U4678 (N_4678,In_545,In_2721);
and U4679 (N_4679,In_3996,In_3154);
or U4680 (N_4680,In_3119,In_2566);
xnor U4681 (N_4681,In_1744,In_2772);
and U4682 (N_4682,In_4507,In_1121);
or U4683 (N_4683,In_2316,In_1506);
xor U4684 (N_4684,In_2972,In_2280);
or U4685 (N_4685,In_4979,In_2381);
xor U4686 (N_4686,In_2670,In_3376);
and U4687 (N_4687,In_3363,In_2643);
and U4688 (N_4688,In_4797,In_3469);
nand U4689 (N_4689,In_1354,In_643);
or U4690 (N_4690,In_1712,In_3401);
or U4691 (N_4691,In_3908,In_3429);
and U4692 (N_4692,In_2017,In_772);
nor U4693 (N_4693,In_3133,In_4303);
and U4694 (N_4694,In_3222,In_1477);
nor U4695 (N_4695,In_251,In_1206);
nor U4696 (N_4696,In_419,In_1542);
and U4697 (N_4697,In_1541,In_3391);
nand U4698 (N_4698,In_3131,In_1859);
xor U4699 (N_4699,In_2886,In_1629);
xnor U4700 (N_4700,In_2419,In_4921);
xnor U4701 (N_4701,In_4459,In_3642);
nor U4702 (N_4702,In_1337,In_1412);
nor U4703 (N_4703,In_2534,In_1612);
nand U4704 (N_4704,In_3048,In_1332);
or U4705 (N_4705,In_4549,In_2173);
nor U4706 (N_4706,In_2766,In_2381);
xor U4707 (N_4707,In_2376,In_175);
or U4708 (N_4708,In_2429,In_2482);
nand U4709 (N_4709,In_3136,In_4356);
or U4710 (N_4710,In_2109,In_1692);
nor U4711 (N_4711,In_434,In_3666);
xor U4712 (N_4712,In_2612,In_2175);
xor U4713 (N_4713,In_1036,In_625);
and U4714 (N_4714,In_238,In_1054);
and U4715 (N_4715,In_4094,In_3611);
xor U4716 (N_4716,In_2290,In_493);
or U4717 (N_4717,In_2204,In_3216);
xor U4718 (N_4718,In_3598,In_3363);
nand U4719 (N_4719,In_377,In_1766);
or U4720 (N_4720,In_4439,In_3396);
nand U4721 (N_4721,In_1673,In_476);
and U4722 (N_4722,In_80,In_413);
or U4723 (N_4723,In_4544,In_886);
nor U4724 (N_4724,In_1207,In_4830);
nand U4725 (N_4725,In_3520,In_962);
xnor U4726 (N_4726,In_3461,In_3085);
xor U4727 (N_4727,In_2104,In_1232);
or U4728 (N_4728,In_4381,In_2673);
and U4729 (N_4729,In_3064,In_1240);
or U4730 (N_4730,In_1323,In_2153);
and U4731 (N_4731,In_993,In_1986);
or U4732 (N_4732,In_3182,In_2755);
and U4733 (N_4733,In_2629,In_4879);
and U4734 (N_4734,In_3667,In_386);
nor U4735 (N_4735,In_897,In_3604);
or U4736 (N_4736,In_4691,In_2424);
nand U4737 (N_4737,In_477,In_4552);
nand U4738 (N_4738,In_524,In_4745);
xnor U4739 (N_4739,In_1531,In_3267);
nor U4740 (N_4740,In_589,In_378);
or U4741 (N_4741,In_120,In_2196);
nand U4742 (N_4742,In_209,In_2251);
nor U4743 (N_4743,In_3877,In_2093);
and U4744 (N_4744,In_2422,In_982);
nor U4745 (N_4745,In_2595,In_4524);
and U4746 (N_4746,In_219,In_1604);
or U4747 (N_4747,In_3269,In_1143);
nor U4748 (N_4748,In_1735,In_258);
and U4749 (N_4749,In_2729,In_4923);
and U4750 (N_4750,In_2369,In_1753);
and U4751 (N_4751,In_2577,In_1831);
and U4752 (N_4752,In_2061,In_4080);
or U4753 (N_4753,In_1290,In_3825);
nor U4754 (N_4754,In_3295,In_1775);
nor U4755 (N_4755,In_1736,In_493);
nor U4756 (N_4756,In_4754,In_1594);
or U4757 (N_4757,In_3252,In_3420);
xnor U4758 (N_4758,In_1987,In_1307);
nand U4759 (N_4759,In_4722,In_1267);
or U4760 (N_4760,In_2726,In_253);
xnor U4761 (N_4761,In_165,In_4321);
and U4762 (N_4762,In_218,In_2809);
nor U4763 (N_4763,In_4653,In_1840);
and U4764 (N_4764,In_1371,In_3803);
or U4765 (N_4765,In_4251,In_2941);
or U4766 (N_4766,In_3183,In_1479);
nor U4767 (N_4767,In_3110,In_4898);
nand U4768 (N_4768,In_745,In_4589);
or U4769 (N_4769,In_202,In_847);
and U4770 (N_4770,In_4024,In_2070);
nor U4771 (N_4771,In_1862,In_2977);
nand U4772 (N_4772,In_1670,In_4133);
or U4773 (N_4773,In_1143,In_4433);
xnor U4774 (N_4774,In_3707,In_3601);
nor U4775 (N_4775,In_4819,In_1280);
or U4776 (N_4776,In_2130,In_1294);
xor U4777 (N_4777,In_476,In_3824);
nor U4778 (N_4778,In_1172,In_2900);
nand U4779 (N_4779,In_1778,In_2555);
xnor U4780 (N_4780,In_2846,In_2821);
or U4781 (N_4781,In_4475,In_4536);
and U4782 (N_4782,In_2872,In_2769);
or U4783 (N_4783,In_4535,In_3271);
and U4784 (N_4784,In_358,In_4359);
nor U4785 (N_4785,In_274,In_2219);
nand U4786 (N_4786,In_2823,In_1465);
xnor U4787 (N_4787,In_1563,In_3237);
xor U4788 (N_4788,In_3301,In_3321);
xnor U4789 (N_4789,In_3804,In_2581);
or U4790 (N_4790,In_4308,In_2190);
nor U4791 (N_4791,In_1550,In_46);
nand U4792 (N_4792,In_1154,In_488);
nor U4793 (N_4793,In_4228,In_3281);
nor U4794 (N_4794,In_2780,In_3812);
or U4795 (N_4795,In_3618,In_4508);
nand U4796 (N_4796,In_1649,In_6);
or U4797 (N_4797,In_912,In_1401);
and U4798 (N_4798,In_1652,In_955);
xor U4799 (N_4799,In_3639,In_504);
nor U4800 (N_4800,In_3138,In_2818);
xnor U4801 (N_4801,In_926,In_2594);
and U4802 (N_4802,In_2734,In_4148);
nor U4803 (N_4803,In_682,In_3490);
xnor U4804 (N_4804,In_1775,In_3263);
nand U4805 (N_4805,In_123,In_1585);
nand U4806 (N_4806,In_2330,In_103);
and U4807 (N_4807,In_4697,In_3635);
nor U4808 (N_4808,In_1083,In_3832);
nor U4809 (N_4809,In_570,In_3961);
and U4810 (N_4810,In_2438,In_2786);
or U4811 (N_4811,In_100,In_2520);
xnor U4812 (N_4812,In_4219,In_1448);
nand U4813 (N_4813,In_3541,In_4010);
nand U4814 (N_4814,In_4305,In_4351);
xnor U4815 (N_4815,In_2145,In_3609);
and U4816 (N_4816,In_1957,In_2546);
nor U4817 (N_4817,In_1982,In_210);
or U4818 (N_4818,In_890,In_2465);
or U4819 (N_4819,In_2909,In_4070);
or U4820 (N_4820,In_99,In_4324);
or U4821 (N_4821,In_2129,In_4960);
xor U4822 (N_4822,In_1552,In_4246);
or U4823 (N_4823,In_2340,In_1627);
xnor U4824 (N_4824,In_2386,In_162);
or U4825 (N_4825,In_2425,In_4226);
and U4826 (N_4826,In_921,In_4800);
and U4827 (N_4827,In_2241,In_813);
and U4828 (N_4828,In_4377,In_1652);
and U4829 (N_4829,In_1320,In_595);
or U4830 (N_4830,In_1929,In_2048);
and U4831 (N_4831,In_317,In_2992);
nor U4832 (N_4832,In_103,In_1927);
nor U4833 (N_4833,In_815,In_1122);
nor U4834 (N_4834,In_645,In_2777);
nand U4835 (N_4835,In_2413,In_4400);
xnor U4836 (N_4836,In_2527,In_2239);
and U4837 (N_4837,In_67,In_4521);
and U4838 (N_4838,In_3756,In_2913);
and U4839 (N_4839,In_4056,In_1209);
xnor U4840 (N_4840,In_93,In_1595);
nand U4841 (N_4841,In_1398,In_2612);
or U4842 (N_4842,In_3870,In_3427);
or U4843 (N_4843,In_4239,In_1985);
and U4844 (N_4844,In_1026,In_3901);
or U4845 (N_4845,In_4541,In_2456);
and U4846 (N_4846,In_814,In_357);
nor U4847 (N_4847,In_8,In_882);
nor U4848 (N_4848,In_4840,In_2077);
nand U4849 (N_4849,In_53,In_2337);
or U4850 (N_4850,In_3555,In_347);
or U4851 (N_4851,In_148,In_3833);
nor U4852 (N_4852,In_289,In_3308);
nand U4853 (N_4853,In_309,In_2189);
xnor U4854 (N_4854,In_3972,In_3414);
and U4855 (N_4855,In_1202,In_4294);
xor U4856 (N_4856,In_2013,In_4687);
nor U4857 (N_4857,In_3698,In_1631);
or U4858 (N_4858,In_1247,In_4733);
nor U4859 (N_4859,In_853,In_2456);
nand U4860 (N_4860,In_2396,In_2416);
nor U4861 (N_4861,In_1276,In_2118);
or U4862 (N_4862,In_3353,In_3876);
xnor U4863 (N_4863,In_4065,In_2276);
and U4864 (N_4864,In_563,In_2271);
xor U4865 (N_4865,In_2058,In_1900);
nand U4866 (N_4866,In_891,In_3097);
and U4867 (N_4867,In_1257,In_1743);
and U4868 (N_4868,In_1022,In_1917);
xnor U4869 (N_4869,In_4595,In_4545);
and U4870 (N_4870,In_2707,In_2599);
xnor U4871 (N_4871,In_3559,In_283);
nor U4872 (N_4872,In_1842,In_4894);
xor U4873 (N_4873,In_823,In_618);
or U4874 (N_4874,In_2096,In_3668);
and U4875 (N_4875,In_4862,In_4986);
xor U4876 (N_4876,In_2577,In_4385);
nor U4877 (N_4877,In_3535,In_1250);
or U4878 (N_4878,In_1634,In_3423);
nor U4879 (N_4879,In_4354,In_2459);
or U4880 (N_4880,In_976,In_4303);
xnor U4881 (N_4881,In_954,In_2446);
xnor U4882 (N_4882,In_2618,In_3763);
nor U4883 (N_4883,In_174,In_4826);
xnor U4884 (N_4884,In_2446,In_346);
xor U4885 (N_4885,In_3948,In_1252);
nand U4886 (N_4886,In_763,In_3684);
nand U4887 (N_4887,In_1468,In_4060);
nor U4888 (N_4888,In_3795,In_2071);
nor U4889 (N_4889,In_904,In_4225);
nand U4890 (N_4890,In_91,In_2501);
and U4891 (N_4891,In_4307,In_4304);
nand U4892 (N_4892,In_816,In_404);
or U4893 (N_4893,In_3707,In_1977);
and U4894 (N_4894,In_4804,In_1738);
nor U4895 (N_4895,In_1516,In_622);
and U4896 (N_4896,In_4402,In_816);
or U4897 (N_4897,In_4515,In_4674);
nor U4898 (N_4898,In_2215,In_1794);
xnor U4899 (N_4899,In_1629,In_4321);
xor U4900 (N_4900,In_462,In_3968);
nand U4901 (N_4901,In_3585,In_3384);
nor U4902 (N_4902,In_2155,In_2501);
and U4903 (N_4903,In_2567,In_2167);
xor U4904 (N_4904,In_2982,In_3884);
nand U4905 (N_4905,In_3192,In_2814);
or U4906 (N_4906,In_4459,In_1125);
nand U4907 (N_4907,In_2097,In_4492);
nand U4908 (N_4908,In_1599,In_736);
nand U4909 (N_4909,In_3670,In_340);
or U4910 (N_4910,In_1881,In_1950);
or U4911 (N_4911,In_4979,In_1593);
nor U4912 (N_4912,In_1991,In_6);
xnor U4913 (N_4913,In_563,In_4852);
xnor U4914 (N_4914,In_2512,In_4277);
nand U4915 (N_4915,In_1592,In_1238);
and U4916 (N_4916,In_1219,In_1197);
nor U4917 (N_4917,In_1224,In_4816);
nor U4918 (N_4918,In_3881,In_3230);
xor U4919 (N_4919,In_4766,In_1406);
and U4920 (N_4920,In_3980,In_3933);
and U4921 (N_4921,In_2165,In_4538);
and U4922 (N_4922,In_4080,In_1490);
nor U4923 (N_4923,In_2800,In_127);
or U4924 (N_4924,In_2178,In_433);
xor U4925 (N_4925,In_142,In_834);
or U4926 (N_4926,In_1557,In_2225);
xnor U4927 (N_4927,In_1392,In_1839);
nor U4928 (N_4928,In_192,In_3727);
nand U4929 (N_4929,In_188,In_568);
nand U4930 (N_4930,In_1902,In_3027);
nor U4931 (N_4931,In_1942,In_236);
xnor U4932 (N_4932,In_4542,In_3007);
or U4933 (N_4933,In_4310,In_254);
nand U4934 (N_4934,In_288,In_4278);
and U4935 (N_4935,In_4780,In_4442);
or U4936 (N_4936,In_4830,In_544);
nand U4937 (N_4937,In_1363,In_4903);
nor U4938 (N_4938,In_4707,In_2365);
nor U4939 (N_4939,In_1890,In_1195);
or U4940 (N_4940,In_3179,In_4752);
or U4941 (N_4941,In_4071,In_1352);
and U4942 (N_4942,In_1210,In_770);
or U4943 (N_4943,In_1956,In_643);
xor U4944 (N_4944,In_910,In_4821);
and U4945 (N_4945,In_513,In_1347);
nor U4946 (N_4946,In_1001,In_3899);
or U4947 (N_4947,In_899,In_1474);
or U4948 (N_4948,In_3712,In_2095);
xnor U4949 (N_4949,In_3904,In_692);
and U4950 (N_4950,In_19,In_4163);
or U4951 (N_4951,In_1239,In_1723);
or U4952 (N_4952,In_2299,In_4007);
and U4953 (N_4953,In_925,In_2987);
or U4954 (N_4954,In_4049,In_4414);
nor U4955 (N_4955,In_2031,In_2603);
and U4956 (N_4956,In_4067,In_4264);
or U4957 (N_4957,In_52,In_665);
or U4958 (N_4958,In_315,In_3339);
nor U4959 (N_4959,In_4426,In_1886);
or U4960 (N_4960,In_1267,In_1652);
nor U4961 (N_4961,In_3019,In_3799);
nand U4962 (N_4962,In_365,In_1779);
nand U4963 (N_4963,In_3719,In_4438);
and U4964 (N_4964,In_2649,In_2103);
nor U4965 (N_4965,In_717,In_1762);
and U4966 (N_4966,In_4936,In_3444);
or U4967 (N_4967,In_2022,In_30);
xor U4968 (N_4968,In_862,In_984);
and U4969 (N_4969,In_2784,In_3153);
nand U4970 (N_4970,In_1145,In_544);
xnor U4971 (N_4971,In_1013,In_2757);
nand U4972 (N_4972,In_829,In_3500);
nand U4973 (N_4973,In_2978,In_610);
or U4974 (N_4974,In_656,In_595);
or U4975 (N_4975,In_2316,In_749);
nor U4976 (N_4976,In_4313,In_447);
and U4977 (N_4977,In_2345,In_472);
nand U4978 (N_4978,In_282,In_1448);
nand U4979 (N_4979,In_916,In_3542);
and U4980 (N_4980,In_1347,In_876);
or U4981 (N_4981,In_2854,In_1885);
and U4982 (N_4982,In_89,In_68);
and U4983 (N_4983,In_65,In_2936);
xor U4984 (N_4984,In_958,In_446);
and U4985 (N_4985,In_346,In_1399);
and U4986 (N_4986,In_3463,In_2509);
and U4987 (N_4987,In_3801,In_1189);
and U4988 (N_4988,In_2836,In_376);
or U4989 (N_4989,In_4113,In_1686);
nor U4990 (N_4990,In_1651,In_3191);
or U4991 (N_4991,In_2788,In_506);
nor U4992 (N_4992,In_3989,In_1744);
nand U4993 (N_4993,In_785,In_2154);
nor U4994 (N_4994,In_1047,In_3700);
nand U4995 (N_4995,In_1282,In_4952);
and U4996 (N_4996,In_970,In_483);
and U4997 (N_4997,In_3714,In_4121);
nand U4998 (N_4998,In_1697,In_211);
xor U4999 (N_4999,In_743,In_4048);
or U5000 (N_5000,N_3516,N_2806);
nand U5001 (N_5001,N_2775,N_2837);
nor U5002 (N_5002,N_3711,N_538);
nand U5003 (N_5003,N_3382,N_4016);
xor U5004 (N_5004,N_2980,N_2194);
nand U5005 (N_5005,N_1810,N_3432);
or U5006 (N_5006,N_1530,N_3807);
nor U5007 (N_5007,N_3222,N_3143);
nand U5008 (N_5008,N_3286,N_1599);
or U5009 (N_5009,N_3799,N_4536);
or U5010 (N_5010,N_2645,N_256);
xnor U5011 (N_5011,N_2848,N_1964);
nand U5012 (N_5012,N_136,N_3842);
nor U5013 (N_5013,N_2091,N_923);
and U5014 (N_5014,N_1186,N_2389);
xor U5015 (N_5015,N_3440,N_194);
nand U5016 (N_5016,N_2922,N_232);
nor U5017 (N_5017,N_4030,N_3874);
nor U5018 (N_5018,N_4229,N_3820);
and U5019 (N_5019,N_1280,N_4240);
or U5020 (N_5020,N_779,N_4054);
xor U5021 (N_5021,N_1603,N_3801);
or U5022 (N_5022,N_4864,N_824);
or U5023 (N_5023,N_1840,N_11);
and U5024 (N_5024,N_1566,N_752);
nor U5025 (N_5025,N_1904,N_2513);
nand U5026 (N_5026,N_1938,N_4755);
nand U5027 (N_5027,N_2363,N_4938);
nor U5028 (N_5028,N_3224,N_4799);
and U5029 (N_5029,N_32,N_2051);
nor U5030 (N_5030,N_2063,N_2540);
xor U5031 (N_5031,N_1540,N_3893);
xnor U5032 (N_5032,N_203,N_2706);
nor U5033 (N_5033,N_1570,N_1272);
nor U5034 (N_5034,N_205,N_3275);
and U5035 (N_5035,N_2155,N_3967);
or U5036 (N_5036,N_518,N_2012);
nor U5037 (N_5037,N_4092,N_3024);
and U5038 (N_5038,N_755,N_3168);
or U5039 (N_5039,N_1204,N_743);
xor U5040 (N_5040,N_3529,N_1290);
and U5041 (N_5041,N_1562,N_3839);
xor U5042 (N_5042,N_551,N_1177);
or U5043 (N_5043,N_651,N_1620);
nor U5044 (N_5044,N_4070,N_3954);
and U5045 (N_5045,N_2867,N_3646);
nor U5046 (N_5046,N_855,N_1198);
nor U5047 (N_5047,N_856,N_4301);
xor U5048 (N_5048,N_1278,N_4180);
nand U5049 (N_5049,N_994,N_2139);
and U5050 (N_5050,N_993,N_153);
nor U5051 (N_5051,N_4825,N_570);
nand U5052 (N_5052,N_863,N_312);
xor U5053 (N_5053,N_2360,N_789);
nand U5054 (N_5054,N_4945,N_4298);
xor U5055 (N_5055,N_2106,N_1803);
nand U5056 (N_5056,N_2748,N_2141);
nor U5057 (N_5057,N_2102,N_2392);
and U5058 (N_5058,N_4225,N_2696);
nand U5059 (N_5059,N_3554,N_2662);
nor U5060 (N_5060,N_2167,N_2997);
nand U5061 (N_5061,N_676,N_2142);
nor U5062 (N_5062,N_2314,N_1427);
nand U5063 (N_5063,N_1179,N_2163);
and U5064 (N_5064,N_2116,N_4367);
nand U5065 (N_5065,N_688,N_323);
nor U5066 (N_5066,N_1346,N_3251);
xnor U5067 (N_5067,N_541,N_1705);
xnor U5068 (N_5068,N_4119,N_757);
xnor U5069 (N_5069,N_2971,N_1273);
nor U5070 (N_5070,N_2929,N_4280);
nand U5071 (N_5071,N_395,N_2214);
xor U5072 (N_5072,N_1002,N_14);
xnor U5073 (N_5073,N_3145,N_1515);
nand U5074 (N_5074,N_1792,N_420);
and U5075 (N_5075,N_868,N_4625);
or U5076 (N_5076,N_4918,N_2871);
and U5077 (N_5077,N_1622,N_902);
nor U5078 (N_5078,N_2824,N_4144);
xor U5079 (N_5079,N_2518,N_3634);
nand U5080 (N_5080,N_2726,N_3482);
and U5081 (N_5081,N_35,N_3218);
or U5082 (N_5082,N_2897,N_3715);
nor U5083 (N_5083,N_4838,N_1788);
and U5084 (N_5084,N_707,N_1499);
xnor U5085 (N_5085,N_2455,N_4137);
nand U5086 (N_5086,N_3565,N_2376);
nor U5087 (N_5087,N_4546,N_1460);
and U5088 (N_5088,N_4985,N_1136);
nand U5089 (N_5089,N_3136,N_1604);
nand U5090 (N_5090,N_3696,N_1385);
or U5091 (N_5091,N_796,N_1312);
xnor U5092 (N_5092,N_761,N_1818);
xor U5093 (N_5093,N_2860,N_3741);
or U5094 (N_5094,N_3320,N_4849);
and U5095 (N_5095,N_748,N_507);
and U5096 (N_5096,N_4692,N_614);
nor U5097 (N_5097,N_1434,N_4896);
or U5098 (N_5098,N_1369,N_1423);
or U5099 (N_5099,N_4707,N_1078);
or U5100 (N_5100,N_1138,N_1642);
nor U5101 (N_5101,N_1597,N_3325);
nor U5102 (N_5102,N_1781,N_1697);
nor U5103 (N_5103,N_238,N_4745);
nor U5104 (N_5104,N_3392,N_826);
or U5105 (N_5105,N_2820,N_4005);
or U5106 (N_5106,N_4636,N_1421);
and U5107 (N_5107,N_1924,N_2138);
nand U5108 (N_5108,N_2781,N_3614);
and U5109 (N_5109,N_3819,N_1174);
nand U5110 (N_5110,N_984,N_4680);
xnor U5111 (N_5111,N_3683,N_596);
or U5112 (N_5112,N_1183,N_4894);
nor U5113 (N_5113,N_869,N_3973);
nand U5114 (N_5114,N_3597,N_1378);
nor U5115 (N_5115,N_3705,N_525);
or U5116 (N_5116,N_894,N_3399);
or U5117 (N_5117,N_2803,N_643);
xnor U5118 (N_5118,N_961,N_3099);
xor U5119 (N_5119,N_1744,N_3075);
nand U5120 (N_5120,N_2898,N_652);
and U5121 (N_5121,N_4758,N_1428);
or U5122 (N_5122,N_2839,N_3074);
and U5123 (N_5123,N_1758,N_3528);
and U5124 (N_5124,N_990,N_3864);
nor U5125 (N_5125,N_831,N_4722);
or U5126 (N_5126,N_3598,N_432);
or U5127 (N_5127,N_3602,N_4174);
nand U5128 (N_5128,N_3905,N_3285);
xor U5129 (N_5129,N_2219,N_34);
or U5130 (N_5130,N_2632,N_4423);
nand U5131 (N_5131,N_4014,N_1898);
and U5132 (N_5132,N_2182,N_4669);
nor U5133 (N_5133,N_2725,N_849);
or U5134 (N_5134,N_1891,N_2996);
or U5135 (N_5135,N_331,N_1981);
xor U5136 (N_5136,N_2197,N_292);
and U5137 (N_5137,N_4658,N_3794);
xnor U5138 (N_5138,N_1234,N_3913);
xor U5139 (N_5139,N_3412,N_513);
and U5140 (N_5140,N_368,N_3685);
xnor U5141 (N_5141,N_3497,N_3613);
nand U5142 (N_5142,N_1324,N_2737);
nor U5143 (N_5143,N_3311,N_2157);
nor U5144 (N_5144,N_883,N_781);
or U5145 (N_5145,N_29,N_1381);
nand U5146 (N_5146,N_4798,N_1111);
nand U5147 (N_5147,N_731,N_3235);
nand U5148 (N_5148,N_4528,N_3501);
nand U5149 (N_5149,N_3771,N_1621);
and U5150 (N_5150,N_759,N_3126);
nand U5151 (N_5151,N_3479,N_4740);
and U5152 (N_5152,N_1229,N_1316);
nor U5153 (N_5153,N_644,N_2491);
nand U5154 (N_5154,N_3548,N_1587);
nor U5155 (N_5155,N_4618,N_2066);
nand U5156 (N_5156,N_1940,N_3828);
nand U5157 (N_5157,N_1257,N_4125);
or U5158 (N_5158,N_2093,N_2624);
or U5159 (N_5159,N_1197,N_2836);
or U5160 (N_5160,N_2653,N_3978);
xnor U5161 (N_5161,N_907,N_3826);
nor U5162 (N_5162,N_3784,N_172);
or U5163 (N_5163,N_1220,N_3225);
xor U5164 (N_5164,N_1990,N_2186);
and U5165 (N_5165,N_243,N_2739);
and U5166 (N_5166,N_3393,N_2944);
xnor U5167 (N_5167,N_3322,N_2162);
nor U5168 (N_5168,N_2549,N_3612);
xor U5169 (N_5169,N_3180,N_4565);
or U5170 (N_5170,N_615,N_4580);
nand U5171 (N_5171,N_3474,N_4322);
and U5172 (N_5172,N_934,N_1471);
and U5173 (N_5173,N_3005,N_4404);
xnor U5174 (N_5174,N_1255,N_545);
and U5175 (N_5175,N_4900,N_4357);
nor U5176 (N_5176,N_4492,N_2904);
xor U5177 (N_5177,N_2807,N_2418);
nand U5178 (N_5178,N_542,N_4791);
and U5179 (N_5179,N_805,N_1976);
nand U5180 (N_5180,N_4866,N_4169);
xnor U5181 (N_5181,N_4397,N_106);
nand U5182 (N_5182,N_3464,N_957);
and U5183 (N_5183,N_1484,N_784);
xor U5184 (N_5184,N_4993,N_566);
or U5185 (N_5185,N_4624,N_341);
and U5186 (N_5186,N_3241,N_2232);
xor U5187 (N_5187,N_4364,N_1349);
nor U5188 (N_5188,N_2691,N_2057);
nor U5189 (N_5189,N_1582,N_1038);
and U5190 (N_5190,N_4205,N_4428);
or U5191 (N_5191,N_2069,N_641);
xnor U5192 (N_5192,N_386,N_574);
or U5193 (N_5193,N_3526,N_2723);
nand U5194 (N_5194,N_2667,N_2893);
nor U5195 (N_5195,N_2500,N_4507);
nand U5196 (N_5196,N_3456,N_1413);
and U5197 (N_5197,N_2067,N_1624);
or U5198 (N_5198,N_601,N_810);
and U5199 (N_5199,N_879,N_898);
or U5200 (N_5200,N_160,N_4813);
nor U5201 (N_5201,N_1106,N_1087);
nand U5202 (N_5202,N_1768,N_744);
or U5203 (N_5203,N_938,N_335);
or U5204 (N_5204,N_4365,N_4575);
xnor U5205 (N_5205,N_1206,N_773);
or U5206 (N_5206,N_964,N_3427);
nor U5207 (N_5207,N_587,N_2296);
and U5208 (N_5208,N_771,N_239);
or U5209 (N_5209,N_1655,N_2629);
nor U5210 (N_5210,N_4915,N_1497);
nand U5211 (N_5211,N_358,N_3390);
or U5212 (N_5212,N_3712,N_4858);
or U5213 (N_5213,N_556,N_3971);
xor U5214 (N_5214,N_4065,N_2841);
nand U5215 (N_5215,N_3453,N_2778);
or U5216 (N_5216,N_76,N_4292);
or U5217 (N_5217,N_1927,N_4186);
and U5218 (N_5218,N_2939,N_4673);
or U5219 (N_5219,N_4973,N_1634);
xnor U5220 (N_5220,N_1590,N_3909);
nor U5221 (N_5221,N_3237,N_924);
nor U5222 (N_5222,N_1814,N_971);
xnor U5223 (N_5223,N_111,N_2364);
nand U5224 (N_5224,N_4188,N_3611);
or U5225 (N_5225,N_770,N_3883);
or U5226 (N_5226,N_227,N_4192);
xor U5227 (N_5227,N_4376,N_2432);
nand U5228 (N_5228,N_1490,N_1779);
xor U5229 (N_5229,N_1693,N_2006);
xor U5230 (N_5230,N_502,N_1609);
nand U5231 (N_5231,N_355,N_1059);
nor U5232 (N_5232,N_307,N_144);
nand U5233 (N_5233,N_2011,N_2238);
xor U5234 (N_5234,N_1881,N_3994);
nand U5235 (N_5235,N_460,N_2615);
or U5236 (N_5236,N_3762,N_1580);
nand U5237 (N_5237,N_2796,N_3965);
and U5238 (N_5238,N_741,N_4141);
nor U5239 (N_5239,N_3633,N_2179);
nor U5240 (N_5240,N_860,N_4668);
nand U5241 (N_5241,N_4793,N_1920);
or U5242 (N_5242,N_612,N_148);
and U5243 (N_5243,N_2150,N_2253);
or U5244 (N_5244,N_778,N_3106);
or U5245 (N_5245,N_4777,N_4541);
and U5246 (N_5246,N_983,N_288);
and U5247 (N_5247,N_819,N_2354);
nor U5248 (N_5248,N_4530,N_2474);
and U5249 (N_5249,N_3146,N_2669);
or U5250 (N_5250,N_4111,N_582);
or U5251 (N_5251,N_378,N_3525);
and U5252 (N_5252,N_499,N_413);
xor U5253 (N_5253,N_3092,N_2041);
nor U5254 (N_5254,N_569,N_270);
nor U5255 (N_5255,N_762,N_2398);
nand U5256 (N_5256,N_4456,N_3498);
or U5257 (N_5257,N_4004,N_2265);
and U5258 (N_5258,N_1332,N_1928);
or U5259 (N_5259,N_4461,N_3162);
nor U5260 (N_5260,N_665,N_4075);
nor U5261 (N_5261,N_303,N_1856);
and U5262 (N_5262,N_2813,N_1752);
xnor U5263 (N_5263,N_4374,N_445);
xor U5264 (N_5264,N_2908,N_1209);
nand U5265 (N_5265,N_274,N_1438);
or U5266 (N_5266,N_1035,N_2936);
xor U5267 (N_5267,N_89,N_2703);
xor U5268 (N_5268,N_4071,N_1284);
and U5269 (N_5269,N_3844,N_1857);
and U5270 (N_5270,N_3221,N_1995);
or U5271 (N_5271,N_2925,N_1345);
and U5272 (N_5272,N_456,N_428);
xor U5273 (N_5273,N_366,N_4809);
nand U5274 (N_5274,N_969,N_2889);
or U5275 (N_5275,N_423,N_3128);
nand U5276 (N_5276,N_4060,N_4018);
or U5277 (N_5277,N_3449,N_2923);
or U5278 (N_5278,N_2911,N_1973);
xnor U5279 (N_5279,N_1151,N_843);
xor U5280 (N_5280,N_3191,N_1246);
or U5281 (N_5281,N_2484,N_324);
xor U5282 (N_5282,N_1951,N_1550);
nor U5283 (N_5283,N_154,N_163);
nand U5284 (N_5284,N_4421,N_3764);
nor U5285 (N_5285,N_371,N_2494);
nand U5286 (N_5286,N_3103,N_4287);
or U5287 (N_5287,N_1980,N_3273);
xor U5288 (N_5288,N_3307,N_1672);
and U5289 (N_5289,N_4744,N_1314);
nand U5290 (N_5290,N_4366,N_2178);
nand U5291 (N_5291,N_4262,N_3022);
or U5292 (N_5292,N_3077,N_3381);
and U5293 (N_5293,N_53,N_3278);
and U5294 (N_5294,N_613,N_2466);
and U5295 (N_5295,N_2810,N_404);
and U5296 (N_5296,N_4852,N_2207);
nand U5297 (N_5297,N_58,N_4406);
nor U5298 (N_5298,N_1532,N_997);
nor U5299 (N_5299,N_2794,N_2187);
xor U5300 (N_5300,N_1911,N_686);
or U5301 (N_5301,N_897,N_2597);
or U5302 (N_5302,N_215,N_3398);
nor U5303 (N_5303,N_4316,N_2853);
xor U5304 (N_5304,N_4664,N_4170);
and U5305 (N_5305,N_1780,N_3493);
nor U5306 (N_5306,N_1236,N_1508);
nand U5307 (N_5307,N_4941,N_4089);
nand U5308 (N_5308,N_1707,N_1537);
xor U5309 (N_5309,N_4485,N_91);
nand U5310 (N_5310,N_1491,N_2708);
nand U5311 (N_5311,N_311,N_3429);
or U5312 (N_5312,N_291,N_605);
xor U5313 (N_5313,N_334,N_1359);
and U5314 (N_5314,N_4402,N_623);
xor U5315 (N_5315,N_4264,N_1353);
nand U5316 (N_5316,N_2920,N_4245);
or U5317 (N_5317,N_580,N_1786);
or U5318 (N_5318,N_1579,N_462);
nand U5319 (N_5319,N_3009,N_1401);
and U5320 (N_5320,N_4455,N_3034);
nand U5321 (N_5321,N_4390,N_186);
and U5322 (N_5322,N_1101,N_852);
xnor U5323 (N_5323,N_717,N_2267);
and U5324 (N_5324,N_749,N_3047);
or U5325 (N_5325,N_2899,N_4677);
or U5326 (N_5326,N_2188,N_1119);
xor U5327 (N_5327,N_39,N_2246);
and U5328 (N_5328,N_3886,N_1041);
xnor U5329 (N_5329,N_1083,N_1800);
or U5330 (N_5330,N_3013,N_4066);
xnor U5331 (N_5331,N_1504,N_4251);
and U5332 (N_5332,N_3818,N_4597);
and U5333 (N_5333,N_3450,N_4290);
or U5334 (N_5334,N_2200,N_1261);
or U5335 (N_5335,N_1252,N_4401);
nor U5336 (N_5336,N_4459,N_913);
xor U5337 (N_5337,N_2673,N_4749);
nand U5338 (N_5338,N_1102,N_1551);
and U5339 (N_5339,N_2013,N_650);
or U5340 (N_5340,N_1966,N_581);
nand U5341 (N_5341,N_1009,N_1380);
or U5342 (N_5342,N_4465,N_760);
nand U5343 (N_5343,N_3197,N_108);
nand U5344 (N_5344,N_1948,N_2617);
xor U5345 (N_5345,N_105,N_4679);
or U5346 (N_5346,N_955,N_2528);
nand U5347 (N_5347,N_281,N_3433);
and U5348 (N_5348,N_740,N_68);
and U5349 (N_5349,N_3186,N_164);
and U5350 (N_5350,N_2568,N_2875);
nand U5351 (N_5351,N_2507,N_4796);
or U5352 (N_5352,N_1137,N_681);
or U5353 (N_5353,N_197,N_2674);
xnor U5354 (N_5354,N_3740,N_1836);
and U5355 (N_5355,N_3882,N_2647);
nor U5356 (N_5356,N_1367,N_787);
and U5357 (N_5357,N_3804,N_562);
and U5358 (N_5358,N_4183,N_4487);
or U5359 (N_5359,N_3253,N_280);
and U5360 (N_5360,N_1266,N_703);
nand U5361 (N_5361,N_2019,N_851);
nor U5362 (N_5362,N_3137,N_123);
or U5363 (N_5363,N_2514,N_2438);
or U5364 (N_5364,N_2872,N_906);
and U5365 (N_5365,N_3256,N_2124);
nor U5366 (N_5366,N_440,N_2329);
xnor U5367 (N_5367,N_113,N_3364);
nor U5368 (N_5368,N_2955,N_2924);
and U5369 (N_5369,N_3063,N_4439);
nor U5370 (N_5370,N_628,N_3451);
nor U5371 (N_5371,N_3060,N_1825);
and U5372 (N_5372,N_2270,N_479);
nor U5373 (N_5373,N_2605,N_2917);
nor U5374 (N_5374,N_3488,N_1157);
or U5375 (N_5375,N_3508,N_3161);
or U5376 (N_5376,N_4691,N_2385);
nand U5377 (N_5377,N_4425,N_3182);
nor U5378 (N_5378,N_2834,N_301);
nor U5379 (N_5379,N_689,N_2791);
and U5380 (N_5380,N_3265,N_4368);
nor U5381 (N_5381,N_3543,N_3366);
nand U5382 (N_5382,N_1320,N_1325);
or U5383 (N_5383,N_4931,N_486);
nand U5384 (N_5384,N_604,N_4810);
and U5385 (N_5385,N_3689,N_2025);
nand U5386 (N_5386,N_3607,N_2879);
nor U5387 (N_5387,N_1171,N_3987);
or U5388 (N_5388,N_1931,N_1987);
xor U5389 (N_5389,N_3347,N_4898);
nand U5390 (N_5390,N_2797,N_3862);
nand U5391 (N_5391,N_3968,N_3416);
nand U5392 (N_5392,N_1961,N_453);
or U5393 (N_5393,N_1044,N_4353);
nand U5394 (N_5394,N_2761,N_121);
xor U5395 (N_5395,N_975,N_2490);
nor U5396 (N_5396,N_880,N_4458);
and U5397 (N_5397,N_4874,N_3386);
nor U5398 (N_5398,N_2445,N_308);
nand U5399 (N_5399,N_3231,N_4248);
or U5400 (N_5400,N_3732,N_3838);
or U5401 (N_5401,N_3,N_4164);
nand U5402 (N_5402,N_3343,N_573);
xnor U5403 (N_5403,N_1014,N_1318);
nand U5404 (N_5404,N_3644,N_4362);
xnor U5405 (N_5405,N_3591,N_3044);
and U5406 (N_5406,N_692,N_4380);
and U5407 (N_5407,N_572,N_1328);
nor U5408 (N_5408,N_4077,N_1949);
or U5409 (N_5409,N_2016,N_2847);
nand U5410 (N_5410,N_2552,N_1999);
nor U5411 (N_5411,N_3108,N_374);
nor U5412 (N_5412,N_4410,N_4579);
nor U5413 (N_5413,N_87,N_3439);
xor U5414 (N_5414,N_1555,N_2998);
or U5415 (N_5415,N_2574,N_1790);
or U5416 (N_5416,N_625,N_4808);
xnor U5417 (N_5417,N_1929,N_1013);
and U5418 (N_5418,N_261,N_4836);
xor U5419 (N_5419,N_4925,N_2566);
nand U5420 (N_5420,N_1190,N_2874);
and U5421 (N_5421,N_1667,N_4539);
xor U5422 (N_5422,N_4942,N_4592);
xor U5423 (N_5423,N_3217,N_2685);
and U5424 (N_5424,N_3487,N_4662);
nand U5425 (N_5425,N_409,N_3463);
nand U5426 (N_5426,N_4695,N_2712);
xor U5427 (N_5427,N_1215,N_2564);
or U5428 (N_5428,N_2121,N_3491);
and U5429 (N_5429,N_618,N_2961);
or U5430 (N_5430,N_2830,N_1224);
xnor U5431 (N_5431,N_2580,N_1558);
or U5432 (N_5432,N_3867,N_3691);
or U5433 (N_5433,N_4643,N_3116);
nor U5434 (N_5434,N_2992,N_3514);
nand U5435 (N_5435,N_795,N_1068);
nand U5436 (N_5436,N_553,N_157);
or U5437 (N_5437,N_908,N_2895);
or U5438 (N_5438,N_1945,N_1592);
nand U5439 (N_5439,N_1776,N_1680);
xor U5440 (N_5440,N_3769,N_3720);
nand U5441 (N_5441,N_543,N_3139);
nand U5442 (N_5442,N_1439,N_477);
xor U5443 (N_5443,N_3869,N_255);
and U5444 (N_5444,N_454,N_2312);
nor U5445 (N_5445,N_664,N_901);
or U5446 (N_5446,N_196,N_2419);
or U5447 (N_5447,N_490,N_687);
xnor U5448 (N_5448,N_3518,N_4746);
nor U5449 (N_5449,N_2988,N_4827);
xor U5450 (N_5450,N_3816,N_1660);
nand U5451 (N_5451,N_1307,N_4675);
and U5452 (N_5452,N_2821,N_1548);
and U5453 (N_5453,N_2517,N_4951);
xnor U5454 (N_5454,N_1057,N_2918);
nand U5455 (N_5455,N_647,N_2914);
or U5456 (N_5456,N_4355,N_1598);
nand U5457 (N_5457,N_2391,N_3735);
and U5458 (N_5458,N_1860,N_1983);
xor U5459 (N_5459,N_4232,N_1889);
or U5460 (N_5460,N_4626,N_4286);
and U5461 (N_5461,N_1795,N_3353);
nor U5462 (N_5462,N_3761,N_3890);
nor U5463 (N_5463,N_4129,N_2560);
nor U5464 (N_5464,N_4068,N_4552);
xnor U5465 (N_5465,N_4094,N_2581);
or U5466 (N_5466,N_3444,N_3173);
and U5467 (N_5467,N_790,N_4860);
nor U5468 (N_5468,N_3248,N_234);
or U5469 (N_5469,N_4202,N_4992);
nor U5470 (N_5470,N_704,N_4194);
xor U5471 (N_5471,N_3561,N_1559);
and U5472 (N_5472,N_2680,N_658);
nor U5473 (N_5473,N_1109,N_3308);
xnor U5474 (N_5474,N_1180,N_3317);
or U5475 (N_5475,N_377,N_2711);
or U5476 (N_5476,N_1631,N_617);
or U5477 (N_5477,N_4314,N_4467);
or U5478 (N_5478,N_1042,N_2047);
nand U5479 (N_5479,N_3425,N_4504);
nand U5480 (N_5480,N_364,N_4215);
and U5481 (N_5481,N_2159,N_626);
xnor U5482 (N_5482,N_3421,N_3927);
xnor U5483 (N_5483,N_4613,N_3292);
and U5484 (N_5484,N_2442,N_3797);
or U5485 (N_5485,N_184,N_1478);
nand U5486 (N_5486,N_2417,N_2263);
nand U5487 (N_5487,N_1214,N_989);
nand U5488 (N_5488,N_2381,N_3000);
or U5489 (N_5489,N_903,N_3375);
or U5490 (N_5490,N_3345,N_2147);
and U5491 (N_5491,N_786,N_2592);
or U5492 (N_5492,N_3981,N_2695);
nand U5493 (N_5493,N_2681,N_970);
nor U5494 (N_5494,N_2509,N_259);
nand U5495 (N_5495,N_461,N_4820);
and U5496 (N_5496,N_2910,N_724);
nor U5497 (N_5497,N_1746,N_2690);
or U5498 (N_5498,N_812,N_2291);
and U5499 (N_5499,N_4157,N_2994);
or U5500 (N_5500,N_954,N_3558);
nand U5501 (N_5501,N_4757,N_4763);
xor U5502 (N_5502,N_591,N_742);
nand U5503 (N_5503,N_2152,N_356);
or U5504 (N_5504,N_3389,N_4438);
or U5505 (N_5505,N_2003,N_3076);
nor U5506 (N_5506,N_4817,N_3262);
nor U5507 (N_5507,N_4142,N_2809);
or U5508 (N_5508,N_2584,N_1392);
nand U5509 (N_5509,N_1384,N_791);
or U5510 (N_5510,N_3023,N_2370);
xor U5511 (N_5511,N_3664,N_4025);
or U5512 (N_5512,N_2416,N_2294);
or U5513 (N_5513,N_3605,N_3172);
nand U5514 (N_5514,N_2359,N_3590);
or U5515 (N_5515,N_2477,N_4317);
and U5516 (N_5516,N_1016,N_1944);
nand U5517 (N_5517,N_1837,N_2262);
xnor U5518 (N_5518,N_2702,N_532);
or U5519 (N_5519,N_1017,N_2423);
nand U5520 (N_5520,N_4551,N_862);
or U5521 (N_5521,N_3411,N_275);
nor U5522 (N_5522,N_2991,N_4484);
or U5523 (N_5523,N_1123,N_895);
nand U5524 (N_5524,N_1391,N_4855);
and U5525 (N_5525,N_1716,N_1118);
xnor U5526 (N_5526,N_2909,N_1309);
nor U5527 (N_5527,N_4462,N_4720);
nand U5528 (N_5528,N_2610,N_523);
and U5529 (N_5529,N_3750,N_1750);
nor U5530 (N_5530,N_1237,N_3208);
and U5531 (N_5531,N_1601,N_2465);
xor U5532 (N_5532,N_1658,N_3171);
nand U5533 (N_5533,N_2334,N_2402);
nand U5534 (N_5534,N_2343,N_4501);
xor U5535 (N_5535,N_4705,N_2499);
nor U5536 (N_5536,N_251,N_41);
and U5537 (N_5537,N_3144,N_2603);
or U5538 (N_5538,N_3545,N_2604);
and U5539 (N_5539,N_4429,N_1105);
nand U5540 (N_5540,N_1015,N_2295);
nand U5541 (N_5541,N_2833,N_3587);
nor U5542 (N_5542,N_180,N_4538);
nand U5543 (N_5543,N_3368,N_4482);
nor U5544 (N_5544,N_2114,N_3223);
and U5545 (N_5545,N_1383,N_2932);
nor U5546 (N_5546,N_536,N_3585);
nor U5547 (N_5547,N_4189,N_4034);
xor U5548 (N_5548,N_702,N_2169);
nand U5549 (N_5549,N_110,N_4486);
nand U5550 (N_5550,N_1643,N_2868);
xnor U5551 (N_5551,N_3852,N_2733);
nor U5552 (N_5552,N_4250,N_2520);
and U5553 (N_5553,N_1146,N_2349);
and U5554 (N_5554,N_3532,N_1757);
and U5555 (N_5555,N_1028,N_1355);
xor U5556 (N_5556,N_3378,N_4372);
and U5557 (N_5557,N_190,N_2181);
nor U5558 (N_5558,N_3854,N_1503);
xnor U5559 (N_5559,N_2264,N_1285);
nor U5560 (N_5560,N_3277,N_2213);
or U5561 (N_5561,N_827,N_3454);
and U5562 (N_5562,N_4247,N_842);
and U5563 (N_5563,N_3007,N_2488);
nor U5564 (N_5564,N_3656,N_447);
xor U5565 (N_5565,N_431,N_2043);
nor U5566 (N_5566,N_4646,N_4922);
nor U5567 (N_5567,N_1851,N_133);
nand U5568 (N_5568,N_1748,N_2081);
or U5569 (N_5569,N_3635,N_733);
xnor U5570 (N_5570,N_4399,N_3885);
xor U5571 (N_5571,N_4097,N_4683);
nor U5572 (N_5572,N_1242,N_1571);
xor U5573 (N_5573,N_1751,N_2);
xor U5574 (N_5574,N_119,N_2954);
xor U5575 (N_5575,N_1791,N_3374);
and U5576 (N_5576,N_4804,N_3782);
nor U5577 (N_5577,N_398,N_4446);
nor U5578 (N_5578,N_2982,N_829);
nand U5579 (N_5579,N_3845,N_915);
nand U5580 (N_5580,N_2745,N_185);
xnor U5581 (N_5581,N_977,N_2134);
nand U5582 (N_5582,N_2223,N_4979);
xnor U5583 (N_5583,N_2230,N_3944);
nor U5584 (N_5584,N_2059,N_4490);
nand U5585 (N_5585,N_3876,N_3859);
and U5586 (N_5586,N_670,N_156);
and U5587 (N_5587,N_4952,N_426);
nand U5588 (N_5588,N_3541,N_2896);
xnor U5589 (N_5589,N_427,N_400);
xnor U5590 (N_5590,N_4426,N_4223);
nor U5591 (N_5591,N_1483,N_1093);
nor U5592 (N_5592,N_4811,N_4771);
and U5593 (N_5593,N_4787,N_2963);
and U5594 (N_5594,N_4656,N_1049);
or U5595 (N_5595,N_3901,N_2229);
xor U5596 (N_5596,N_3661,N_1441);
and U5597 (N_5597,N_4831,N_3070);
nand U5598 (N_5598,N_1583,N_2611);
and U5599 (N_5599,N_974,N_1420);
nand U5600 (N_5600,N_4064,N_273);
nand U5601 (N_5601,N_2964,N_3228);
xnor U5602 (N_5602,N_340,N_2462);
nand U5603 (N_5603,N_2736,N_3894);
and U5604 (N_5604,N_2248,N_3174);
or U5605 (N_5605,N_4956,N_1430);
nand U5606 (N_5606,N_3069,N_3053);
or U5607 (N_5607,N_4468,N_2710);
nand U5608 (N_5608,N_1262,N_3288);
xor U5609 (N_5609,N_1143,N_4469);
nor U5610 (N_5610,N_1694,N_4328);
xnor U5611 (N_5611,N_3693,N_735);
or U5612 (N_5612,N_1816,N_1591);
nor U5613 (N_5613,N_266,N_691);
or U5614 (N_5614,N_383,N_804);
nand U5615 (N_5615,N_2765,N_1341);
or U5616 (N_5616,N_2731,N_3962);
nor U5617 (N_5617,N_1670,N_4405);
xnor U5618 (N_5618,N_3485,N_3998);
and U5619 (N_5619,N_2793,N_1866);
xnor U5620 (N_5620,N_4038,N_4233);
nor U5621 (N_5621,N_2974,N_1544);
nor U5622 (N_5622,N_1389,N_813);
nor U5623 (N_5623,N_1572,N_4448);
xnor U5624 (N_5624,N_2826,N_1379);
or U5625 (N_5625,N_2709,N_4761);
nor U5626 (N_5626,N_4647,N_1227);
nor U5627 (N_5627,N_4637,N_4252);
and U5628 (N_5628,N_2539,N_3743);
or U5629 (N_5629,N_1424,N_3388);
xnor U5630 (N_5630,N_1398,N_3932);
and U5631 (N_5631,N_4214,N_2656);
and U5632 (N_5632,N_3800,N_3673);
and U5633 (N_5633,N_2087,N_1573);
nand U5634 (N_5634,N_510,N_1947);
nand U5635 (N_5635,N_4253,N_4570);
xor U5636 (N_5636,N_682,N_1249);
nand U5637 (N_5637,N_1095,N_1577);
nor U5638 (N_5638,N_4550,N_4865);
and U5639 (N_5639,N_1772,N_2422);
and U5640 (N_5640,N_526,N_4553);
and U5641 (N_5641,N_2023,N_3997);
or U5642 (N_5642,N_1809,N_963);
nand U5643 (N_5643,N_4713,N_4434);
nor U5644 (N_5644,N_756,N_3097);
xnor U5645 (N_5645,N_2070,N_2271);
nor U5646 (N_5646,N_3287,N_3610);
or U5647 (N_5647,N_968,N_2355);
and U5648 (N_5648,N_2947,N_2430);
nand U5649 (N_5649,N_2628,N_4574);
xnor U5650 (N_5650,N_4464,N_836);
nand U5651 (N_5651,N_2715,N_2274);
and U5652 (N_5652,N_2727,N_2104);
nand U5653 (N_5653,N_1982,N_2790);
or U5654 (N_5654,N_584,N_3054);
and U5655 (N_5655,N_3884,N_3329);
and U5656 (N_5656,N_4901,N_222);
and U5657 (N_5657,N_1736,N_2687);
or U5658 (N_5658,N_546,N_4807);
nand U5659 (N_5659,N_2887,N_2510);
xnor U5660 (N_5660,N_459,N_4265);
nor U5661 (N_5661,N_2464,N_1511);
xnor U5662 (N_5662,N_920,N_714);
xnor U5663 (N_5663,N_18,N_146);
and U5664 (N_5664,N_2301,N_2838);
xnor U5665 (N_5665,N_4598,N_1213);
xnor U5666 (N_5666,N_264,N_211);
nor U5667 (N_5667,N_3744,N_2353);
nor U5668 (N_5668,N_3475,N_841);
or U5669 (N_5669,N_1815,N_1279);
nor U5670 (N_5670,N_1037,N_2434);
nand U5671 (N_5671,N_3827,N_3989);
nor U5672 (N_5672,N_2435,N_2255);
xnor U5673 (N_5673,N_4267,N_1880);
nand U5674 (N_5674,N_3247,N_4480);
nor U5675 (N_5675,N_962,N_4524);
xnor U5676 (N_5676,N_4659,N_555);
or U5677 (N_5677,N_4748,N_3582);
and U5678 (N_5678,N_2095,N_1492);
and U5679 (N_5679,N_1552,N_1107);
and U5680 (N_5680,N_2545,N_4518);
or U5681 (N_5681,N_4171,N_2769);
and U5682 (N_5682,N_3272,N_861);
and U5683 (N_5683,N_823,N_982);
or U5684 (N_5684,N_1885,N_3050);
nor U5685 (N_5685,N_3408,N_2743);
xnor U5686 (N_5686,N_2487,N_385);
nand U5687 (N_5687,N_564,N_2039);
xor U5688 (N_5688,N_1335,N_2015);
nand U5689 (N_5689,N_1077,N_3899);
and U5690 (N_5690,N_2304,N_3821);
and U5691 (N_5691,N_1376,N_1862);
or U5692 (N_5692,N_3324,N_3361);
nand U5693 (N_5693,N_137,N_4666);
or U5694 (N_5694,N_13,N_4868);
and U5695 (N_5695,N_2055,N_2643);
nor U5696 (N_5696,N_942,N_600);
and U5697 (N_5697,N_1630,N_2357);
nand U5698 (N_5698,N_4148,N_3809);
nand U5699 (N_5699,N_3326,N_4095);
nand U5700 (N_5700,N_3441,N_16);
nand U5701 (N_5701,N_3723,N_3476);
or U5702 (N_5702,N_1088,N_3924);
nor U5703 (N_5703,N_350,N_3730);
xor U5704 (N_5704,N_4085,N_47);
nand U5705 (N_5705,N_4760,N_3431);
nor U5706 (N_5706,N_1985,N_1615);
or U5707 (N_5707,N_3383,N_2249);
nor U5708 (N_5708,N_4756,N_1473);
nand U5709 (N_5709,N_4079,N_61);
and U5710 (N_5710,N_4601,N_4988);
nand U5711 (N_5711,N_4285,N_866);
xnor U5712 (N_5712,N_4195,N_4862);
and U5713 (N_5713,N_1760,N_1565);
and U5714 (N_5714,N_2475,N_598);
and U5715 (N_5715,N_859,N_1482);
nor U5716 (N_5716,N_4344,N_1735);
nand U5717 (N_5717,N_78,N_4440);
nand U5718 (N_5718,N_149,N_3192);
or U5719 (N_5719,N_2108,N_4602);
nand U5720 (N_5720,N_4512,N_1403);
nor U5721 (N_5721,N_3484,N_2154);
and U5722 (N_5722,N_4686,N_3555);
xnor U5723 (N_5723,N_2127,N_1720);
or U5724 (N_5724,N_2587,N_95);
or U5725 (N_5725,N_4236,N_2308);
and U5726 (N_5726,N_4432,N_699);
nor U5727 (N_5727,N_1442,N_1538);
xnor U5728 (N_5728,N_2092,N_3912);
nand U5729 (N_5729,N_4104,N_2000);
or U5730 (N_5730,N_1493,N_4466);
or U5731 (N_5731,N_709,N_470);
nand U5732 (N_5732,N_3813,N_1308);
and U5733 (N_5733,N_241,N_3133);
xor U5734 (N_5734,N_3089,N_390);
nor U5735 (N_5735,N_4533,N_3785);
or U5736 (N_5736,N_1637,N_3535);
nor U5737 (N_5737,N_2780,N_4361);
xnor U5738 (N_5738,N_1070,N_3269);
nand U5739 (N_5739,N_2508,N_4776);
xor U5740 (N_5740,N_2942,N_2855);
nand U5741 (N_5741,N_589,N_2128);
nand U5742 (N_5742,N_2812,N_3947);
or U5743 (N_5743,N_351,N_2857);
nor U5744 (N_5744,N_3267,N_320);
and U5745 (N_5745,N_1554,N_4515);
xor U5746 (N_5746,N_4619,N_2211);
xor U5747 (N_5747,N_3995,N_3694);
xnor U5748 (N_5748,N_3726,N_4715);
or U5749 (N_5749,N_4330,N_593);
nand U5750 (N_5750,N_2277,N_1437);
nor U5751 (N_5751,N_3149,N_3775);
or U5752 (N_5752,N_1048,N_100);
or U5753 (N_5753,N_1612,N_1507);
nor U5754 (N_5754,N_3156,N_3209);
or U5755 (N_5755,N_305,N_4102);
nor U5756 (N_5756,N_3734,N_229);
nand U5757 (N_5757,N_1681,N_1159);
nor U5758 (N_5758,N_2082,N_1834);
xnor U5759 (N_5759,N_1822,N_1201);
nor U5760 (N_5760,N_3304,N_3462);
or U5761 (N_5761,N_339,N_772);
nor U5762 (N_5762,N_3637,N_1794);
nand U5763 (N_5763,N_1941,N_1970);
nand U5764 (N_5764,N_973,N_2078);
xor U5765 (N_5765,N_4989,N_4105);
and U5766 (N_5766,N_3817,N_3282);
or U5767 (N_5767,N_174,N_1713);
nor U5768 (N_5768,N_2753,N_4347);
nand U5769 (N_5769,N_1100,N_967);
xnor U5770 (N_5770,N_4640,N_3323);
and U5771 (N_5771,N_3234,N_2501);
nor U5772 (N_5772,N_1766,N_4012);
xnor U5773 (N_5773,N_3465,N_195);
nor U5774 (N_5774,N_2831,N_3066);
and U5775 (N_5775,N_2399,N_4050);
or U5776 (N_5776,N_4706,N_1939);
xor U5777 (N_5777,N_2236,N_2086);
nand U5778 (N_5778,N_3240,N_3030);
or U5779 (N_5779,N_2358,N_1303);
and U5780 (N_5780,N_1638,N_2582);
nor U5781 (N_5781,N_3232,N_3752);
nor U5782 (N_5782,N_3202,N_1076);
and U5783 (N_5783,N_2986,N_4230);
and U5784 (N_5784,N_1154,N_4711);
and U5785 (N_5785,N_1243,N_4764);
xnor U5786 (N_5786,N_4568,N_4026);
or U5787 (N_5787,N_3102,N_2310);
nor U5788 (N_5788,N_2216,N_2307);
xnor U5789 (N_5789,N_3333,N_1842);
and U5790 (N_5790,N_1365,N_7);
or U5791 (N_5791,N_6,N_3229);
and U5792 (N_5792,N_4386,N_2426);
nor U5793 (N_5793,N_2945,N_416);
nand U5794 (N_5794,N_2217,N_2524);
and U5795 (N_5795,N_1451,N_2661);
or U5796 (N_5796,N_4443,N_4888);
xor U5797 (N_5797,N_1594,N_4936);
nor U5798 (N_5798,N_3891,N_3062);
and U5799 (N_5799,N_1930,N_1426);
xnor U5800 (N_5800,N_245,N_3018);
xor U5801 (N_5801,N_4877,N_3313);
nor U5802 (N_5802,N_4294,N_3650);
or U5803 (N_5803,N_3132,N_3065);
nand U5804 (N_5804,N_1518,N_2675);
nand U5805 (N_5805,N_3579,N_3766);
xor U5806 (N_5806,N_284,N_1764);
or U5807 (N_5807,N_392,N_656);
nor U5808 (N_5808,N_2290,N_4377);
nand U5809 (N_5809,N_3533,N_4444);
xnor U5810 (N_5810,N_2498,N_4564);
xnor U5811 (N_5811,N_3078,N_4650);
or U5812 (N_5812,N_3658,N_1953);
or U5813 (N_5813,N_45,N_2882);
or U5814 (N_5814,N_659,N_4098);
nor U5815 (N_5815,N_1468,N_4326);
xnor U5816 (N_5816,N_1130,N_4130);
and U5817 (N_5817,N_2639,N_3321);
nand U5818 (N_5818,N_3666,N_176);
or U5819 (N_5819,N_1350,N_4795);
and U5820 (N_5820,N_159,N_4593);
xnor U5821 (N_5821,N_3698,N_3352);
and U5822 (N_5822,N_109,N_3640);
nor U5823 (N_5823,N_491,N_2210);
nand U5824 (N_5824,N_3719,N_4712);
or U5825 (N_5825,N_4657,N_3194);
nand U5826 (N_5826,N_3980,N_2240);
and U5827 (N_5827,N_1520,N_1163);
nor U5828 (N_5828,N_3625,N_655);
and U5829 (N_5829,N_1046,N_2575);
or U5830 (N_5830,N_4371,N_2973);
nor U5831 (N_5831,N_4124,N_2458);
nand U5832 (N_5832,N_3592,N_3200);
nor U5833 (N_5833,N_36,N_987);
nor U5834 (N_5834,N_4832,N_558);
and U5835 (N_5835,N_1829,N_4334);
nand U5836 (N_5836,N_3617,N_4061);
nor U5837 (N_5837,N_4846,N_1900);
nor U5838 (N_5838,N_49,N_3088);
nand U5839 (N_5839,N_4031,N_1464);
or U5840 (N_5840,N_2635,N_198);
nor U5841 (N_5841,N_344,N_1363);
and U5842 (N_5842,N_4067,N_178);
nand U5843 (N_5843,N_774,N_4678);
or U5844 (N_5844,N_2705,N_4879);
and U5845 (N_5845,N_4156,N_2631);
nor U5846 (N_5846,N_3651,N_1725);
nand U5847 (N_5847,N_1639,N_2981);
nand U5848 (N_5848,N_482,N_4906);
nand U5849 (N_5849,N_2651,N_2117);
xor U5850 (N_5850,N_2559,N_1921);
nand U5851 (N_5851,N_55,N_4850);
or U5852 (N_5852,N_4177,N_2452);
xnor U5853 (N_5853,N_4221,N_4788);
or U5854 (N_5854,N_929,N_3036);
and U5855 (N_5855,N_3315,N_4616);
and U5856 (N_5856,N_4349,N_1606);
and U5857 (N_5857,N_279,N_2005);
xor U5858 (N_5858,N_3624,N_2077);
nand U5859 (N_5859,N_4379,N_4590);
xor U5860 (N_5860,N_3350,N_4537);
and U5861 (N_5861,N_1863,N_4165);
or U5862 (N_5862,N_1870,N_4903);
nand U5863 (N_5863,N_1745,N_3889);
xor U5864 (N_5864,N_3888,N_2819);
nor U5865 (N_5865,N_3742,N_3153);
nor U5866 (N_5866,N_571,N_4622);
nand U5867 (N_5867,N_2823,N_4971);
nor U5868 (N_5868,N_4867,N_2439);
or U5869 (N_5869,N_4946,N_4542);
nand U5870 (N_5870,N_4641,N_3957);
xor U5871 (N_5871,N_3648,N_662);
nand U5872 (N_5872,N_4099,N_1479);
or U5873 (N_5873,N_3250,N_4088);
or U5874 (N_5874,N_4905,N_3643);
nor U5875 (N_5875,N_3629,N_3653);
nor U5876 (N_5876,N_2828,N_2096);
and U5877 (N_5877,N_1908,N_1600);
and U5878 (N_5878,N_4917,N_293);
and U5879 (N_5879,N_3380,N_2205);
xnor U5880 (N_5880,N_900,N_2302);
or U5881 (N_5881,N_2449,N_1498);
xor U5882 (N_5882,N_363,N_4277);
or U5883 (N_5883,N_1922,N_3812);
or U5884 (N_5884,N_2161,N_1708);
nand U5885 (N_5885,N_3420,N_2541);
and U5886 (N_5886,N_2856,N_4147);
nor U5887 (N_5887,N_4032,N_30);
xnor U5888 (N_5888,N_918,N_4954);
and U5889 (N_5889,N_2554,N_4519);
xor U5890 (N_5890,N_4638,N_3057);
xor U5891 (N_5891,N_3770,N_3911);
nor U5892 (N_5892,N_2189,N_1641);
nor U5893 (N_5893,N_1718,N_3716);
nor U5894 (N_5894,N_1178,N_4474);
nor U5895 (N_5895,N_10,N_3283);
or U5896 (N_5896,N_1432,N_1608);
and U5897 (N_5897,N_3974,N_188);
nor U5898 (N_5898,N_1988,N_4346);
nor U5899 (N_5899,N_439,N_2503);
or U5900 (N_5900,N_1877,N_2622);
and U5901 (N_5901,N_283,N_3717);
nor U5902 (N_5902,N_544,N_2767);
nor U5903 (N_5903,N_2144,N_999);
or U5904 (N_5904,N_1546,N_2033);
and U5905 (N_5905,N_3094,N_115);
nand U5906 (N_5906,N_4375,N_2371);
and U5907 (N_5907,N_1959,N_690);
nand U5908 (N_5908,N_4964,N_2367);
xor U5909 (N_5909,N_3296,N_2282);
xnor U5910 (N_5910,N_3684,N_2774);
and U5911 (N_5911,N_797,N_1443);
nor U5912 (N_5912,N_412,N_1323);
and U5913 (N_5913,N_4881,N_3045);
nor U5914 (N_5914,N_1126,N_4983);
xor U5915 (N_5915,N_3603,N_249);
xor U5916 (N_5916,N_401,N_561);
and U5917 (N_5917,N_608,N_2561);
and U5918 (N_5918,N_3127,N_1917);
and U5919 (N_5919,N_960,N_373);
and U5920 (N_5920,N_1117,N_3340);
or U5921 (N_5921,N_1375,N_4431);
nor U5922 (N_5922,N_1542,N_1458);
and U5923 (N_5923,N_737,N_143);
and U5924 (N_5924,N_4308,N_3682);
nor U5925 (N_5925,N_4872,N_450);
nor U5926 (N_5926,N_4709,N_2678);
xor U5927 (N_5927,N_3765,N_2327);
nor U5928 (N_5928,N_3991,N_2018);
xor U5929 (N_5929,N_2873,N_85);
and U5930 (N_5930,N_2766,N_3397);
and U5931 (N_5931,N_4974,N_1322);
nand U5932 (N_5932,N_207,N_1741);
xor U5933 (N_5933,N_4818,N_3517);
xor U5934 (N_5934,N_4393,N_1906);
or U5935 (N_5935,N_1344,N_4114);
nand U5936 (N_5936,N_2995,N_3511);
or U5937 (N_5937,N_3895,N_1333);
xor U5938 (N_5938,N_2467,N_712);
nand U5939 (N_5939,N_1162,N_4778);
and U5940 (N_5940,N_2268,N_25);
nand U5941 (N_5941,N_1291,N_4237);
nand U5942 (N_5942,N_2553,N_2594);
nor U5943 (N_5943,N_4644,N_1689);
nand U5944 (N_5944,N_4609,N_60);
xnor U5945 (N_5945,N_4084,N_2021);
and U5946 (N_5946,N_2113,N_3227);
and U5947 (N_5947,N_4342,N_43);
nor U5948 (N_5948,N_2787,N_1390);
xor U5949 (N_5949,N_3107,N_847);
xor U5950 (N_5950,N_4694,N_3632);
xor U5951 (N_5951,N_2372,N_4970);
or U5952 (N_5952,N_725,N_4300);
xor U5953 (N_5953,N_1,N_4835);
and U5954 (N_5954,N_1371,N_4115);
or U5955 (N_5955,N_3958,N_2100);
or U5956 (N_5956,N_48,N_4549);
nand U5957 (N_5957,N_173,N_4794);
nand U5958 (N_5958,N_269,N_4965);
nand U5959 (N_5959,N_4193,N_753);
nor U5960 (N_5960,N_4845,N_4847);
nor U5961 (N_5961,N_2845,N_3949);
and U5962 (N_5962,N_2129,N_1765);
xnor U5963 (N_5963,N_1021,N_4476);
xor U5964 (N_5964,N_418,N_1358);
nand U5965 (N_5965,N_524,N_3866);
xor U5966 (N_5966,N_3831,N_3537);
nor U5967 (N_5967,N_2912,N_3138);
xnor U5968 (N_5968,N_4197,N_2595);
or U5969 (N_5969,N_1007,N_3865);
or U5970 (N_5970,N_3626,N_648);
nor U5971 (N_5971,N_4151,N_2065);
and U5972 (N_5972,N_4685,N_2007);
nor U5973 (N_5973,N_3600,N_3639);
nand U5974 (N_5974,N_4400,N_4087);
or U5975 (N_5975,N_4670,N_2829);
or U5976 (N_5976,N_2572,N_2657);
or U5977 (N_5977,N_365,N_4841);
or U5978 (N_5978,N_2962,N_3215);
or U5979 (N_5979,N_4509,N_1000);
nor U5980 (N_5980,N_265,N_1124);
nand U5981 (N_5981,N_3165,N_3986);
and U5982 (N_5982,N_1463,N_1932);
and U5983 (N_5983,N_4027,N_3279);
or U5984 (N_5984,N_4076,N_2752);
and U5985 (N_5985,N_1543,N_3370);
and U5986 (N_5986,N_4876,N_4500);
xor U5987 (N_5987,N_3979,N_1811);
xnor U5988 (N_5988,N_535,N_4690);
xor U5989 (N_5989,N_875,N_2135);
nor U5990 (N_5990,N_3369,N_128);
nand U5991 (N_5991,N_1971,N_3348);
nor U5992 (N_5992,N_1545,N_2751);
xor U5993 (N_5993,N_4608,N_1871);
xor U5994 (N_5994,N_560,N_607);
or U5995 (N_5995,N_3822,N_3972);
nor U5996 (N_5996,N_258,N_1915);
nor U5997 (N_5997,N_3051,N_2891);
or U5998 (N_5998,N_3549,N_3114);
xor U5999 (N_5999,N_1470,N_1184);
nor U6000 (N_6000,N_3574,N_1469);
or U6001 (N_6001,N_332,N_142);
nand U6002 (N_6002,N_3026,N_1675);
xor U6003 (N_6003,N_3520,N_1625);
or U6004 (N_6004,N_4737,N_147);
nand U6005 (N_6005,N_1429,N_2245);
and U6006 (N_6006,N_2459,N_4980);
nand U6007 (N_6007,N_1414,N_3175);
xor U6008 (N_6008,N_747,N_3594);
nor U6009 (N_6009,N_3155,N_4433);
xnor U6010 (N_6010,N_4672,N_3372);
nor U6011 (N_6011,N_66,N_4303);
nand U6012 (N_6012,N_1449,N_2448);
or U6013 (N_6013,N_3295,N_1113);
nor U6014 (N_6014,N_3907,N_710);
or U6015 (N_6015,N_3249,N_4020);
nor U6016 (N_6016,N_2447,N_3833);
xnor U6017 (N_6017,N_2782,N_2489);
nand U6018 (N_6018,N_1073,N_2048);
nand U6019 (N_6019,N_638,N_2827);
nor U6020 (N_6020,N_443,N_26);
nor U6021 (N_6021,N_4382,N_2621);
xor U6022 (N_6022,N_4961,N_4209);
nor U6023 (N_6023,N_2746,N_3930);
and U6024 (N_6024,N_1129,N_250);
or U6025 (N_6025,N_2160,N_1082);
xor U6026 (N_6026,N_354,N_705);
xor U6027 (N_6027,N_3032,N_171);
nor U6028 (N_6028,N_1433,N_2620);
xor U6029 (N_6029,N_4053,N_548);
nor U6030 (N_6030,N_1416,N_2030);
nor U6031 (N_6031,N_2865,N_2808);
nor U6032 (N_6032,N_4520,N_2340);
or U6033 (N_6033,N_1728,N_1972);
or U6034 (N_6034,N_3255,N_3031);
nor U6035 (N_6035,N_1032,N_210);
nor U6036 (N_6036,N_1207,N_4770);
nand U6037 (N_6037,N_4544,N_563);
xor U6038 (N_6038,N_956,N_565);
nand U6039 (N_6039,N_1678,N_1065);
xor U6040 (N_6040,N_799,N_3848);
nor U6041 (N_6041,N_4975,N_3028);
nand U6042 (N_6042,N_533,N_4525);
xor U6043 (N_6043,N_4028,N_1149);
or U6044 (N_6044,N_3125,N_4417);
nor U6045 (N_6045,N_2046,N_3566);
or U6046 (N_6046,N_3043,N_495);
and U6047 (N_6047,N_4231,N_2266);
or U6048 (N_6048,N_1685,N_706);
and U6049 (N_6049,N_3707,N_1890);
nand U6050 (N_6050,N_2300,N_1287);
nor U6051 (N_6051,N_986,N_3943);
xor U6052 (N_6052,N_3692,N_4135);
or U6053 (N_6053,N_4919,N_1040);
nand U6054 (N_6054,N_3703,N_2822);
nor U6055 (N_6055,N_3314,N_4991);
nand U6056 (N_6056,N_3837,N_4044);
and U6057 (N_6057,N_750,N_3767);
or U6058 (N_6058,N_719,N_1975);
xnor U6059 (N_6059,N_271,N_3506);
nand U6060 (N_6060,N_2576,N_2456);
nor U6061 (N_6061,N_2472,N_425);
and U6062 (N_6062,N_2366,N_17);
nor U6063 (N_6063,N_2002,N_1486);
or U6064 (N_6064,N_4293,N_3093);
and U6065 (N_6065,N_1029,N_3259);
and U6066 (N_6066,N_1066,N_2480);
xnor U6067 (N_6067,N_2646,N_2206);
nor U6068 (N_6068,N_1330,N_75);
nor U6069 (N_6069,N_1031,N_1683);
nor U6070 (N_6070,N_1099,N_4735);
nand U6071 (N_6071,N_4783,N_3404);
nor U6072 (N_6072,N_2571,N_1012);
or U6073 (N_6073,N_1956,N_2916);
xor U6074 (N_6074,N_4496,N_1072);
nor U6075 (N_6075,N_2259,N_937);
and U6076 (N_6076,N_4995,N_3117);
xor U6077 (N_6077,N_4610,N_3576);
nand U6078 (N_6078,N_4842,N_286);
or U6079 (N_6079,N_1937,N_4704);
nand U6080 (N_6080,N_679,N_4805);
nand U6081 (N_6081,N_4295,N_3774);
xnor U6082 (N_6082,N_3578,N_2341);
xnor U6083 (N_6083,N_92,N_2074);
or U6084 (N_6084,N_1205,N_2330);
or U6085 (N_6085,N_3802,N_2242);
or U6086 (N_6086,N_2215,N_1882);
xnor U6087 (N_6087,N_406,N_2773);
or U6088 (N_6088,N_2222,N_727);
or U6089 (N_6089,N_2241,N_298);
or U6090 (N_6090,N_3085,N_777);
xnor U6091 (N_6091,N_2276,N_3623);
or U6092 (N_6092,N_2858,N_3534);
and U6093 (N_6093,N_1051,N_4055);
or U6094 (N_6094,N_4721,N_2663);
or U6095 (N_6095,N_1283,N_4605);
xor U6096 (N_6096,N_120,N_4261);
nor U6097 (N_6097,N_1145,N_77);
and U6098 (N_6098,N_4116,N_3903);
nand U6099 (N_6099,N_4667,N_794);
or U6100 (N_6100,N_3409,N_3919);
or U6101 (N_6101,N_4460,N_4332);
nand U6102 (N_6102,N_522,N_667);
nand U6103 (N_6103,N_357,N_2786);
or U6104 (N_6104,N_588,N_4424);
or U6105 (N_6105,N_1998,N_1575);
nor U6106 (N_6106,N_322,N_2641);
nor U6107 (N_6107,N_1415,N_2234);
nor U6108 (N_6108,N_1034,N_4732);
nand U6109 (N_6109,N_1958,N_1412);
and U6110 (N_6110,N_3481,N_646);
xor U6111 (N_6111,N_3982,N_4145);
and U6112 (N_6112,N_4110,N_4069);
or U6113 (N_6113,N_405,N_1271);
xnor U6114 (N_6114,N_4861,N_4033);
and U6115 (N_6115,N_376,N_4373);
xor U6116 (N_6116,N_3798,N_1868);
and U6117 (N_6117,N_267,N_1512);
xor U6118 (N_6118,N_4998,N_1789);
nand U6119 (N_6119,N_4962,N_3160);
and U6120 (N_6120,N_951,N_3458);
and U6121 (N_6121,N_4278,N_3615);
nor U6122 (N_6122,N_2279,N_2137);
xor U6123 (N_6123,N_1487,N_375);
nor U6124 (N_6124,N_4719,N_1160);
and U6125 (N_6125,N_4495,N_421);
nand U6126 (N_6126,N_1298,N_3159);
or U6127 (N_6127,N_3001,N_2742);
nand U6128 (N_6128,N_3207,N_1395);
and U6129 (N_6129,N_4920,N_649);
xor U6130 (N_6130,N_353,N_2637);
and U6131 (N_6131,N_2717,N_1334);
or U6132 (N_6132,N_722,N_2321);
xor U6133 (N_6133,N_4652,N_4837);
or U6134 (N_6134,N_4508,N_1481);
nor U6135 (N_6135,N_2713,N_4937);
and U6136 (N_6136,N_429,N_616);
nor U6137 (N_6137,N_700,N_3396);
nand U6138 (N_6138,N_50,N_3407);
or U6139 (N_6139,N_2851,N_4489);
nor U6140 (N_6140,N_4728,N_745);
or U6141 (N_6141,N_3953,N_3733);
nand U6142 (N_6142,N_3245,N_4928);
nor U6143 (N_6143,N_2429,N_3647);
nand U6144 (N_6144,N_1043,N_3423);
nor U6145 (N_6145,N_3669,N_3213);
nand U6146 (N_6146,N_4306,N_204);
xor U6147 (N_6147,N_4753,N_1883);
or U6148 (N_6148,N_578,N_3778);
nand U6149 (N_6149,N_317,N_1155);
nand U6150 (N_6150,N_1467,N_2938);
and U6151 (N_6151,N_1832,N_2952);
nand U6152 (N_6152,N_3984,N_1150);
and U6153 (N_6153,N_1210,N_2339);
and U6154 (N_6154,N_3738,N_3112);
xnor U6155 (N_6155,N_4582,N_84);
and U6156 (N_6156,N_834,N_904);
xnor U6157 (N_6157,N_2284,N_4689);
and U6158 (N_6158,N_1292,N_1250);
or U6159 (N_6159,N_122,N_4080);
xnor U6160 (N_6160,N_610,N_995);
nand U6161 (N_6161,N_150,N_4968);
nand U6162 (N_6162,N_2722,N_3772);
or U6163 (N_6163,N_677,N_1527);
xor U6164 (N_6164,N_161,N_4126);
nand U6165 (N_6165,N_1485,N_4213);
or U6166 (N_6166,N_1445,N_1801);
xor U6167 (N_6167,N_2347,N_471);
or U6168 (N_6168,N_4477,N_3714);
nor U6169 (N_6169,N_2190,N_2450);
and U6170 (N_6170,N_1560,N_1419);
xor U6171 (N_6171,N_3387,N_4394);
or U6172 (N_6172,N_3331,N_4631);
nor U6173 (N_6173,N_4696,N_1267);
and U6174 (N_6174,N_151,N_1673);
nor U6175 (N_6175,N_4514,N_2612);
nand U6176 (N_6176,N_3786,N_3757);
or U6177 (N_6177,N_2788,N_888);
or U6178 (N_6178,N_1281,N_4297);
and U6179 (N_6179,N_4736,N_4266);
or U6180 (N_6180,N_1645,N_2591);
nor U6181 (N_6181,N_1296,N_102);
and U6182 (N_6182,N_411,N_3702);
nand U6183 (N_6183,N_4986,N_4503);
and U6184 (N_6184,N_83,N_911);
and U6185 (N_6185,N_3627,N_3335);
nor U6186 (N_6186,N_2083,N_1679);
nor U6187 (N_6187,N_1297,N_2172);
xor U6188 (N_6188,N_3187,N_4040);
nor U6189 (N_6189,N_3494,N_4383);
and U6190 (N_6190,N_2609,N_2671);
nand U6191 (N_6191,N_1574,N_3759);
nor U6192 (N_6192,N_1775,N_2906);
nor U6193 (N_6193,N_3019,N_1589);
or U6194 (N_6194,N_2931,N_4338);
nor U6195 (N_6195,N_1813,N_4123);
and U6196 (N_6196,N_4897,N_1895);
or U6197 (N_6197,N_1742,N_1698);
or U6198 (N_6198,N_685,N_4011);
and U6199 (N_6199,N_2585,N_769);
and U6200 (N_6200,N_1640,N_3589);
xnor U6201 (N_6201,N_1819,N_4389);
and U6202 (N_6202,N_3834,N_1476);
xnor U6203 (N_6203,N_498,N_4589);
nor U6204 (N_6204,N_1740,N_931);
or U6205 (N_6205,N_4227,N_1974);
xor U6206 (N_6206,N_945,N_4910);
or U6207 (N_6207,N_953,N_3236);
xnor U6208 (N_6208,N_474,N_4738);
nand U6209 (N_6209,N_1853,N_3988);
or U6210 (N_6210,N_4840,N_3934);
xor U6211 (N_6211,N_214,N_2719);
or U6212 (N_6212,N_2022,N_4572);
nor U6213 (N_6213,N_2654,N_3808);
or U6214 (N_6214,N_3206,N_3118);
or U6215 (N_6215,N_820,N_3436);
and U6216 (N_6216,N_1595,N_2862);
nand U6217 (N_6217,N_1509,N_4645);
xnor U6218 (N_6218,N_352,N_3302);
xnor U6219 (N_6219,N_4273,N_4113);
nand U6220 (N_6220,N_2151,N_3553);
xor U6221 (N_6221,N_2762,N_864);
or U6222 (N_6222,N_2164,N_4257);
nand U6223 (N_6223,N_3608,N_3437);
xor U6224 (N_6224,N_718,N_4022);
xor U6225 (N_6225,N_634,N_1023);
nand U6226 (N_6226,N_4107,N_2131);
xnor U6227 (N_6227,N_4136,N_3619);
nor U6228 (N_6228,N_2993,N_2305);
xnor U6229 (N_6229,N_1131,N_1614);
nand U6230 (N_6230,N_4716,N_3300);
nor U6231 (N_6231,N_552,N_3956);
and U6232 (N_6232,N_3067,N_2079);
nor U6233 (N_6233,N_3021,N_3925);
and U6234 (N_6234,N_2099,N_4772);
xnor U6235 (N_6235,N_4762,N_2648);
xor U6236 (N_6236,N_2626,N_4987);
and U6237 (N_6237,N_3522,N_1821);
xor U6238 (N_6238,N_3468,N_1239);
or U6239 (N_6239,N_952,N_3402);
or U6240 (N_6240,N_2984,N_316);
or U6241 (N_6241,N_1695,N_1796);
and U6242 (N_6242,N_247,N_179);
xnor U6243 (N_6243,N_506,N_559);
xor U6244 (N_6244,N_1733,N_1276);
xnor U6245 (N_6245,N_1300,N_1386);
xnor U6246 (N_6246,N_4318,N_1913);
nand U6247 (N_6247,N_4531,N_1629);
nor U6248 (N_6248,N_2085,N_2209);
xnor U6249 (N_6249,N_2379,N_1329);
nor U6250 (N_6250,N_99,N_101);
xor U6251 (N_6251,N_2320,N_2951);
nor U6252 (N_6252,N_2146,N_1997);
or U6253 (N_6253,N_1116,N_2854);
nand U6254 (N_6254,N_2198,N_1230);
or U6255 (N_6255,N_27,N_2546);
nor U6256 (N_6256,N_1784,N_4561);
nand U6257 (N_6257,N_2551,N_2888);
or U6258 (N_6258,N_3263,N_3630);
xor U6259 (N_6259,N_1274,N_1616);
and U6260 (N_6260,N_2978,N_3193);
nand U6261 (N_6261,N_1907,N_2431);
or U6262 (N_6262,N_890,N_3580);
nand U6263 (N_6263,N_2903,N_1876);
xor U6264 (N_6264,N_2650,N_4049);
xnor U6265 (N_6265,N_1653,N_4211);
nor U6266 (N_6266,N_2816,N_2967);
or U6267 (N_6267,N_278,N_3087);
xnor U6268 (N_6268,N_228,N_289);
nand U6269 (N_6269,N_1304,N_4830);
nand U6270 (N_6270,N_88,N_2755);
xnor U6271 (N_6271,N_1674,N_3131);
and U6272 (N_6272,N_630,N_2958);
nand U6273 (N_6273,N_2732,N_3058);
or U6274 (N_6274,N_2386,N_1172);
or U6275 (N_6275,N_3341,N_131);
or U6276 (N_6276,N_4320,N_2776);
nand U6277 (N_6277,N_4878,N_2204);
xnor U6278 (N_6278,N_4260,N_4959);
or U6279 (N_6279,N_2885,N_4337);
or U6280 (N_6280,N_2421,N_3881);
nand U6281 (N_6281,N_642,N_3524);
and U6282 (N_6282,N_505,N_1979);
nor U6283 (N_6283,N_683,N_2504);
and U6284 (N_6284,N_4090,N_1019);
nand U6285 (N_6285,N_224,N_2852);
nand U6286 (N_6286,N_2326,N_393);
nor U6287 (N_6287,N_3586,N_4584);
or U6288 (N_6288,N_1182,N_4545);
and U6289 (N_6289,N_1372,N_720);
and U6290 (N_6290,N_337,N_793);
nand U6291 (N_6291,N_4534,N_4773);
nor U6292 (N_6292,N_1188,N_3609);
xor U6293 (N_6293,N_2058,N_1366);
nor U6294 (N_6294,N_3338,N_2008);
and U6295 (N_6295,N_4204,N_2446);
or U6296 (N_6296,N_183,N_3832);
nand U6297 (N_6297,N_519,N_4857);
and U6298 (N_6298,N_666,N_4359);
or U6299 (N_6299,N_3900,N_2497);
or U6300 (N_6300,N_4839,N_917);
nand U6301 (N_6301,N_2814,N_1849);
and U6302 (N_6302,N_3025,N_3055);
nor U6303 (N_6303,N_3243,N_181);
nor U6304 (N_6304,N_1222,N_2684);
xnor U6305 (N_6305,N_1001,N_3910);
nor U6306 (N_6306,N_4219,N_3502);
and U6307 (N_6307,N_2260,N_4083);
and U6308 (N_6308,N_1806,N_4497);
and U6309 (N_6309,N_2881,N_73);
nand U6310 (N_6310,N_1233,N_3290);
nor U6311 (N_6311,N_2224,N_4385);
nor U6312 (N_6312,N_2907,N_905);
or U6313 (N_6313,N_818,N_3606);
or U6314 (N_6314,N_1943,N_1058);
nand U6315 (N_6315,N_2965,N_3406);
nor U6316 (N_6316,N_139,N_1513);
xnor U6317 (N_6317,N_1167,N_726);
and U6318 (N_6318,N_452,N_476);
nand U6319 (N_6319,N_2024,N_127);
nor U6320 (N_6320,N_1505,N_1633);
xor U6321 (N_6321,N_2522,N_3560);
nor U6322 (N_6322,N_1260,N_2598);
or U6323 (N_6323,N_1364,N_1892);
and U6324 (N_6324,N_2608,N_81);
and U6325 (N_6325,N_138,N_2724);
or U6326 (N_6326,N_1714,N_4391);
or U6327 (N_6327,N_1450,N_4916);
or U6328 (N_6328,N_594,N_1793);
xnor U6329 (N_6329,N_472,N_4216);
and U6330 (N_6330,N_3312,N_1132);
or U6331 (N_6331,N_3403,N_3357);
and U6332 (N_6332,N_3811,N_632);
nor U6333 (N_6333,N_1846,N_446);
nor U6334 (N_6334,N_467,N_1024);
nand U6335 (N_6335,N_124,N_3959);
and U6336 (N_6336,N_2688,N_2901);
xnor U6337 (N_6337,N_811,N_2655);
and U6338 (N_6338,N_1963,N_4471);
nand U6339 (N_6339,N_4201,N_3298);
and U6340 (N_6340,N_2558,N_4688);
and U6341 (N_6341,N_2401,N_4182);
or U6342 (N_6342,N_4513,N_1844);
xnor U6343 (N_6343,N_1047,N_3377);
or U6344 (N_6344,N_891,N_2049);
nor U6345 (N_6345,N_3424,N_4345);
and U6346 (N_6346,N_3697,N_520);
xor U6347 (N_6347,N_4671,N_3739);
or U6348 (N_6348,N_1218,N_1737);
or U6349 (N_6349,N_939,N_3796);
nor U6350 (N_6350,N_1867,N_517);
or U6351 (N_6351,N_627,N_3027);
and U6352 (N_6352,N_1079,N_947);
xnor U6353 (N_6353,N_1855,N_1701);
and U6354 (N_6354,N_4291,N_3011);
nor U6355 (N_6355,N_1254,N_2306);
or U6356 (N_6356,N_2272,N_1189);
and U6357 (N_6357,N_783,N_4323);
nand U6358 (N_6358,N_3342,N_4167);
or U6359 (N_6359,N_4769,N_2393);
nor U6360 (N_6360,N_1528,N_1715);
nor U6361 (N_6361,N_3795,N_4363);
nand U6362 (N_6362,N_4627,N_835);
and U6363 (N_6363,N_3503,N_2668);
or U6364 (N_6364,N_2573,N_2683);
nand U6365 (N_6365,N_3706,N_1564);
xor U6366 (N_6366,N_1823,N_958);
nand U6367 (N_6367,N_1568,N_2512);
nor U6368 (N_6368,N_3538,N_1462);
or U6369 (N_6369,N_4724,N_2257);
and U6370 (N_6370,N_155,N_2779);
and U6371 (N_6371,N_4315,N_4848);
xor U6372 (N_6372,N_4271,N_4999);
nor U6373 (N_6373,N_2175,N_927);
nand U6374 (N_6374,N_844,N_2485);
nor U6375 (N_6375,N_1547,N_654);
nand U6376 (N_6376,N_919,N_2396);
or U6377 (N_6377,N_2408,N_4210);
nor U6378 (N_6378,N_1388,N_3115);
nand U6379 (N_6379,N_3789,N_1774);
and U6380 (N_6380,N_313,N_3190);
and U6381 (N_6381,N_4411,N_3154);
and U6382 (N_6382,N_701,N_1050);
xnor U6383 (N_6383,N_3020,N_4454);
and U6384 (N_6384,N_4617,N_3135);
and U6385 (N_6385,N_4734,N_4153);
nand U6386 (N_6386,N_2318,N_2119);
nor U6387 (N_6387,N_2010,N_1305);
and U6388 (N_6388,N_2543,N_1156);
or U6389 (N_6389,N_2235,N_1888);
nand U6390 (N_6390,N_287,N_3562);
nand U6391 (N_6391,N_4312,N_2934);
and U6392 (N_6392,N_257,N_4409);
and U6393 (N_6393,N_2293,N_698);
nor U6394 (N_6394,N_2105,N_2054);
and U6395 (N_6395,N_1352,N_3758);
and U6396 (N_6396,N_4522,N_4352);
nand U6397 (N_6397,N_872,N_2700);
nand U6398 (N_6398,N_3141,N_3863);
and U6399 (N_6399,N_315,N_4569);
and U6400 (N_6400,N_2338,N_1247);
and U6401 (N_6401,N_4369,N_2747);
and U6402 (N_6402,N_330,N_3120);
nor U6403 (N_6403,N_4781,N_3654);
or U6404 (N_6404,N_673,N_3556);
and U6405 (N_6405,N_4676,N_1541);
or U6406 (N_6406,N_3737,N_631);
or U6407 (N_6407,N_4594,N_2390);
nand U6408 (N_6408,N_885,N_1659);
and U6409 (N_6409,N_1799,N_3090);
nor U6410 (N_6410,N_4969,N_3337);
or U6411 (N_6411,N_1055,N_4587);
xnor U6412 (N_6412,N_575,N_2623);
nand U6413 (N_6413,N_3166,N_1373);
xnor U6414 (N_6414,N_3668,N_3952);
and U6415 (N_6415,N_410,N_2676);
or U6416 (N_6416,N_3428,N_402);
xor U6417 (N_6417,N_4103,N_4045);
nand U6418 (N_6418,N_2644,N_2220);
or U6419 (N_6419,N_1488,N_2273);
nor U6420 (N_6420,N_1824,N_54);
xnor U6421 (N_6421,N_4588,N_4420);
nor U6422 (N_6422,N_438,N_387);
xor U6423 (N_6423,N_2032,N_998);
and U6424 (N_6424,N_1636,N_2493);
xnor U6425 (N_6425,N_2122,N_4718);
nand U6426 (N_6426,N_2805,N_881);
nor U6427 (N_6427,N_2990,N_2633);
and U6428 (N_6428,N_1875,N_1195);
and U6429 (N_6429,N_483,N_333);
and U6430 (N_6430,N_1175,N_1219);
or U6431 (N_6431,N_3628,N_200);
xnor U6432 (N_6432,N_2784,N_1181);
or U6433 (N_6433,N_2433,N_2323);
and U6434 (N_6434,N_2145,N_1121);
and U6435 (N_6435,N_403,N_2227);
or U6436 (N_6436,N_1743,N_33);
or U6437 (N_6437,N_1661,N_2328);
nor U6438 (N_6438,N_2619,N_2244);
nand U6439 (N_6439,N_2247,N_4674);
or U6440 (N_6440,N_3773,N_3878);
nor U6441 (N_6441,N_2478,N_3896);
nor U6442 (N_6442,N_1841,N_3618);
nor U6443 (N_6443,N_437,N_3756);
nor U6444 (N_6444,N_2170,N_3665);
nand U6445 (N_6445,N_208,N_424);
xnor U6446 (N_6446,N_3442,N_899);
or U6447 (N_6447,N_4560,N_3264);
nor U6448 (N_6448,N_3663,N_3042);
or U6449 (N_6449,N_2471,N_2407);
nor U6450 (N_6450,N_3478,N_2350);
or U6451 (N_6451,N_2089,N_1586);
nor U6452 (N_6452,N_3575,N_1649);
nand U6453 (N_6453,N_833,N_1474);
nor U6454 (N_6454,N_4239,N_4556);
nand U6455 (N_6455,N_4681,N_3542);
and U6456 (N_6456,N_3147,N_4246);
xnor U6457 (N_6457,N_70,N_2740);
nor U6458 (N_6458,N_4003,N_2384);
xnor U6459 (N_6459,N_2311,N_3843);
nor U6460 (N_6460,N_1501,N_4473);
nand U6461 (N_6461,N_1852,N_107);
or U6462 (N_6462,N_4396,N_3745);
nor U6463 (N_6463,N_2870,N_3753);
xnor U6464 (N_6464,N_3455,N_15);
or U6465 (N_6465,N_3599,N_3170);
and U6466 (N_6466,N_4557,N_4437);
nor U6467 (N_6467,N_2444,N_4526);
nor U6468 (N_6468,N_3079,N_4281);
or U6469 (N_6469,N_4698,N_2720);
xnor U6470 (N_6470,N_635,N_285);
and U6471 (N_6471,N_2789,N_2556);
and U6472 (N_6472,N_1387,N_4010);
or U6473 (N_6473,N_1306,N_887);
xnor U6474 (N_6474,N_2243,N_1623);
nor U6475 (N_6475,N_2948,N_2526);
or U6476 (N_6476,N_1724,N_1656);
or U6477 (N_6477,N_1805,N_2133);
or U6478 (N_6478,N_1626,N_1635);
nor U6479 (N_6479,N_4378,N_3219);
xnor U6480 (N_6480,N_3747,N_1526);
nor U6481 (N_6481,N_4573,N_2345);
xnor U6482 (N_6482,N_1302,N_1062);
and U6483 (N_6483,N_4206,N_1831);
xnor U6484 (N_6484,N_488,N_4319);
xnor U6485 (N_6485,N_3873,N_1865);
nor U6486 (N_6486,N_3690,N_2940);
and U6487 (N_6487,N_384,N_4527);
nor U6488 (N_6488,N_4418,N_3914);
and U6489 (N_6489,N_1759,N_4162);
and U6490 (N_6490,N_2966,N_4540);
nand U6491 (N_6491,N_4790,N_620);
or U6492 (N_6492,N_4516,N_235);
nand U6493 (N_6493,N_531,N_1074);
or U6494 (N_6494,N_4430,N_1459);
xor U6495 (N_6495,N_3681,N_4336);
or U6496 (N_6496,N_1986,N_3904);
nor U6497 (N_6497,N_1533,N_2972);
or U6498 (N_6498,N_466,N_2288);
and U6499 (N_6499,N_4710,N_3938);
or U6500 (N_6500,N_4854,N_3492);
and U6501 (N_6501,N_754,N_2894);
or U6502 (N_6502,N_1954,N_871);
nor U6503 (N_6503,N_3319,N_3709);
xnor U6504 (N_6504,N_3365,N_2846);
or U6505 (N_6505,N_2835,N_4001);
and U6506 (N_6506,N_31,N_3573);
and U6507 (N_6507,N_1164,N_695);
and U6508 (N_6508,N_1060,N_1704);
nor U6509 (N_6509,N_858,N_4996);
and U6510 (N_6510,N_2111,N_2652);
or U6511 (N_6511,N_444,N_12);
or U6512 (N_6512,N_838,N_4614);
and U6513 (N_6513,N_1585,N_2226);
or U6514 (N_6514,N_3140,N_1399);
and U6515 (N_6515,N_2035,N_1288);
nand U6516 (N_6516,N_325,N_276);
or U6517 (N_6517,N_4258,N_4743);
nor U6518 (N_6518,N_4427,N_4923);
or U6519 (N_6519,N_2336,N_2125);
nor U6520 (N_6520,N_2682,N_3926);
nand U6521 (N_6521,N_2890,N_1289);
nor U6522 (N_6522,N_4895,N_822);
or U6523 (N_6523,N_1671,N_226);
or U6524 (N_6524,N_2481,N_3923);
or U6525 (N_6525,N_2201,N_2525);
nor U6526 (N_6526,N_4254,N_132);
or U6527 (N_6527,N_1676,N_118);
nand U6528 (N_6528,N_3216,N_3330);
xor U6529 (N_6529,N_4161,N_4307);
or U6530 (N_6530,N_3012,N_1531);
nand U6531 (N_6531,N_3622,N_2694);
xnor U6532 (N_6532,N_1251,N_2840);
or U6533 (N_6533,N_1703,N_776);
nand U6534 (N_6534,N_1521,N_2153);
and U6535 (N_6535,N_3122,N_3515);
or U6536 (N_6536,N_4828,N_96);
nor U6537 (N_6537,N_2256,N_1918);
or U6538 (N_6538,N_300,N_3906);
xnor U6539 (N_6539,N_792,N_1221);
and U6540 (N_6540,N_2937,N_3096);
nor U6541 (N_6541,N_4152,N_4269);
nand U6542 (N_6542,N_4039,N_3495);
nor U6543 (N_6543,N_93,N_4452);
xor U6544 (N_6544,N_4803,N_1030);
nor U6545 (N_6545,N_874,N_825);
or U6546 (N_6546,N_2785,N_1549);
or U6547 (N_6547,N_3875,N_2383);
and U6548 (N_6548,N_455,N_3316);
and U6549 (N_6549,N_3992,N_4869);
xnor U6550 (N_6550,N_4665,N_407);
and U6551 (N_6551,N_2555,N_4621);
xnor U6552 (N_6552,N_1337,N_1069);
xnor U6553 (N_6553,N_515,N_4982);
nor U6554 (N_6554,N_134,N_3261);
nor U6555 (N_6555,N_2729,N_1327);
or U6556 (N_6556,N_4412,N_362);
nor U6557 (N_6557,N_3332,N_4904);
or U6558 (N_6558,N_2413,N_3426);
xor U6559 (N_6559,N_3505,N_3258);
xnor U6560 (N_6560,N_1807,N_3157);
xnor U6561 (N_6561,N_3939,N_349);
xor U6562 (N_6562,N_3595,N_2677);
or U6563 (N_6563,N_4190,N_72);
nand U6564 (N_6564,N_3238,N_3928);
xor U6565 (N_6565,N_3855,N_3993);
xnor U6566 (N_6566,N_3686,N_2970);
nor U6567 (N_6567,N_478,N_1763);
nor U6568 (N_6568,N_2754,N_1235);
or U6569 (N_6569,N_2542,N_2734);
xnor U6570 (N_6570,N_3847,N_1071);
or U6571 (N_6571,N_3996,N_579);
or U6572 (N_6572,N_4984,N_441);
nor U6573 (N_6573,N_1942,N_3109);
or U6574 (N_6574,N_449,N_893);
nor U6575 (N_6575,N_4600,N_1244);
nor U6576 (N_6576,N_3504,N_1110);
and U6577 (N_6577,N_1411,N_2613);
or U6578 (N_6578,N_537,N_2037);
nand U6579 (N_6579,N_1783,N_23);
xor U6580 (N_6580,N_629,N_3983);
nand U6581 (N_6581,N_2665,N_3405);
and U6582 (N_6582,N_3046,N_4506);
nand U6583 (N_6583,N_2315,N_4256);
and U6584 (N_6584,N_4006,N_3446);
nor U6585 (N_6585,N_2946,N_71);
nor U6586 (N_6586,N_602,N_2098);
and U6587 (N_6587,N_4408,N_2064);
and U6588 (N_6588,N_1422,N_4072);
or U6589 (N_6589,N_4343,N_3551);
and U6590 (N_6590,N_74,N_985);
nand U6591 (N_6591,N_3181,N_1301);
nand U6592 (N_6592,N_3169,N_4502);
or U6593 (N_6593,N_4047,N_4108);
and U6594 (N_6594,N_3781,N_4889);
nor U6595 (N_6595,N_1248,N_4255);
and U6596 (N_6596,N_1722,N_1142);
nor U6597 (N_6597,N_4056,N_817);
nor U6598 (N_6598,N_1534,N_2926);
xnor U6599 (N_6599,N_1710,N_2056);
or U6600 (N_6600,N_1240,N_766);
or U6601 (N_6601,N_4759,N_336);
nand U6602 (N_6602,N_2795,N_4112);
nand U6603 (N_6603,N_2979,N_925);
nor U6604 (N_6604,N_1135,N_329);
and U6605 (N_6605,N_1018,N_1648);
nor U6606 (N_6606,N_2252,N_1313);
xnor U6607 (N_6607,N_595,N_1699);
nor U6608 (N_6608,N_20,N_2659);
nand U6609 (N_6609,N_3400,N_4978);
nor U6610 (N_6610,N_2362,N_943);
xor U6611 (N_6611,N_815,N_2849);
or U6612 (N_6612,N_1946,N_4002);
xnor U6613 (N_6613,N_2492,N_1396);
nand U6614 (N_6614,N_2404,N_1086);
or U6615 (N_6615,N_2905,N_2586);
and U6616 (N_6616,N_4187,N_4708);
or U6617 (N_6617,N_4935,N_4532);
nor U6618 (N_6618,N_539,N_1711);
nor U6619 (N_6619,N_1802,N_3567);
or U6620 (N_6620,N_1196,N_3163);
xnor U6621 (N_6621,N_3385,N_1217);
nor U6622 (N_6622,N_3966,N_4882);
and U6623 (N_6623,N_1935,N_2983);
and U6624 (N_6624,N_69,N_803);
nor U6625 (N_6625,N_2728,N_503);
or U6626 (N_6626,N_814,N_2985);
nor U6627 (N_6627,N_2411,N_3188);
nor U6628 (N_6628,N_4654,N_67);
and U6629 (N_6629,N_4559,N_4146);
nor U6630 (N_6630,N_933,N_4403);
xnor U6631 (N_6631,N_4943,N_2801);
or U6632 (N_6632,N_1139,N_4450);
or U6633 (N_6633,N_3788,N_2052);
nand U6634 (N_6634,N_231,N_3123);
nor U6635 (N_6635,N_657,N_2692);
xor U6636 (N_6636,N_2880,N_3346);
nor U6637 (N_6637,N_2878,N_4899);
nand U6638 (N_6638,N_2441,N_2686);
nand U6639 (N_6639,N_4133,N_782);
nor U6640 (N_6640,N_4806,N_4853);
and U6641 (N_6641,N_723,N_3879);
xor U6642 (N_6642,N_4908,N_4566);
nor U6643 (N_6643,N_941,N_2476);
nor U6644 (N_6644,N_1894,N_4766);
or U6645 (N_6645,N_1569,N_1668);
xor U6646 (N_6646,N_788,N_4356);
or U6647 (N_6647,N_2730,N_1203);
xnor U6648 (N_6648,N_2094,N_3671);
nand U6649 (N_6649,N_2026,N_4967);
nand U6650 (N_6650,N_4166,N_3081);
or U6651 (N_6651,N_4911,N_2254);
or U6652 (N_6652,N_4100,N_3430);
nor U6653 (N_6653,N_4358,N_1202);
nor U6654 (N_6654,N_4768,N_3763);
or U6655 (N_6655,N_3731,N_1919);
xor U6656 (N_6656,N_4449,N_4360);
nand U6657 (N_6657,N_2126,N_1893);
xnor U6658 (N_6658,N_3929,N_2636);
nor U6659 (N_6659,N_1475,N_3791);
and U6660 (N_6660,N_2642,N_4037);
or U6661 (N_6661,N_3754,N_145);
xnor U6662 (N_6662,N_4313,N_3072);
and U6663 (N_6663,N_346,N_1664);
nor U6664 (N_6664,N_1677,N_1516);
xnor U6665 (N_6665,N_4535,N_2331);
nand U6666 (N_6666,N_1277,N_2348);
nor U6667 (N_6667,N_4159,N_1268);
or U6668 (N_6668,N_4930,N_1847);
xnor U6669 (N_6669,N_3443,N_4008);
or U6670 (N_6670,N_2861,N_2388);
nand U6671 (N_6671,N_3119,N_3680);
nor U6672 (N_6672,N_2600,N_2352);
and U6673 (N_6673,N_1826,N_708);
nand U6674 (N_6674,N_3183,N_3814);
nor U6675 (N_6675,N_112,N_1405);
xor U6676 (N_6676,N_1153,N_4483);
nor U6677 (N_6677,N_3284,N_1410);
or U6678 (N_6678,N_509,N_1576);
xor U6679 (N_6679,N_3645,N_557);
nand U6680 (N_6680,N_2382,N_4472);
and U6681 (N_6681,N_1294,N_2927);
nor U6682 (N_6682,N_3950,N_4577);
nand U6683 (N_6683,N_2953,N_1084);
xor U6684 (N_6684,N_3469,N_4567);
and U6685 (N_6685,N_611,N_1994);
and U6686 (N_6686,N_3004,N_63);
nand U6687 (N_6687,N_1646,N_4106);
and U6688 (N_6688,N_4081,N_3887);
nor U6689 (N_6689,N_3527,N_3704);
xnor U6690 (N_6690,N_1916,N_1326);
or U6691 (N_6691,N_3080,N_4228);
xor U6692 (N_6692,N_435,N_549);
nand U6693 (N_6693,N_1045,N_1496);
nand U6694 (N_6694,N_473,N_3199);
and U6695 (N_6695,N_1839,N_4422);
or U6696 (N_6696,N_3933,N_367);
nand U6697 (N_6697,N_1194,N_209);
and U6698 (N_6698,N_839,N_3417);
xnor U6699 (N_6699,N_3918,N_4725);
nor U6700 (N_6700,N_3872,N_2397);
xor U6701 (N_6701,N_697,N_3581);
and U6702 (N_6702,N_4801,N_3391);
or U6703 (N_6703,N_2212,N_4885);
and U6704 (N_6704,N_716,N_4249);
nor U6705 (N_6705,N_3226,N_3477);
or U6706 (N_6706,N_3212,N_2975);
or U6707 (N_6707,N_2173,N_2601);
xnor U6708 (N_6708,N_3121,N_4007);
and U6709 (N_6709,N_2625,N_2107);
xor U6710 (N_6710,N_3823,N_3356);
and U6711 (N_6711,N_3557,N_577);
xnor U6712 (N_6712,N_2772,N_299);
or U6713 (N_6713,N_3466,N_4073);
xor U6714 (N_6714,N_1989,N_2177);
nor U6715 (N_6715,N_304,N_3708);
and U6716 (N_6716,N_3008,N_1827);
nand U6717 (N_6717,N_116,N_2286);
nand U6718 (N_6718,N_169,N_399);
and U6719 (N_6719,N_2405,N_4633);
and U6720 (N_6720,N_1557,N_360);
and U6721 (N_6721,N_1495,N_1317);
or U6722 (N_6722,N_4948,N_3336);
nand U6723 (N_6723,N_4649,N_3677);
and U6724 (N_6724,N_3351,N_4000);
nand U6725 (N_6725,N_2440,N_2073);
and U6726 (N_6726,N_221,N_381);
or U6727 (N_6727,N_260,N_4155);
nor U6728 (N_6728,N_3824,N_167);
and U6729 (N_6729,N_2184,N_1500);
xnor U6730 (N_6730,N_1523,N_4702);
and U6731 (N_6731,N_3829,N_1967);
or U6732 (N_6732,N_4160,N_130);
nor U6733 (N_6733,N_1833,N_3710);
nor U6734 (N_6734,N_877,N_876);
or U6735 (N_6735,N_965,N_3362);
or U6736 (N_6736,N_1211,N_3675);
and U6737 (N_6737,N_2036,N_1454);
nor U6738 (N_6738,N_3718,N_4275);
xor U6739 (N_6739,N_3916,N_4934);
or U6740 (N_6740,N_2375,N_1619);
xnor U6741 (N_6741,N_4447,N_1256);
nand U6742 (N_6742,N_4655,N_1581);
and U6743 (N_6743,N_1122,N_1596);
and U6744 (N_6744,N_3486,N_3176);
nand U6745 (N_6745,N_1820,N_394);
xor U6746 (N_6746,N_4859,N_1529);
nand U6747 (N_6747,N_3349,N_4109);
nor U6748 (N_6748,N_4893,N_4914);
nor U6749 (N_6749,N_1914,N_4419);
and U6750 (N_6750,N_4731,N_711);
nor U6751 (N_6751,N_950,N_2799);
or U6752 (N_6752,N_2468,N_2333);
xnor U6753 (N_6753,N_4059,N_4912);
nor U6754 (N_6754,N_1185,N_1275);
or U6755 (N_6755,N_4208,N_4154);
nor U6756 (N_6756,N_2699,N_219);
nand U6757 (N_6757,N_694,N_3946);
and U6758 (N_6758,N_3281,N_2174);
or U6759 (N_6759,N_674,N_306);
and U6760 (N_6760,N_2470,N_1910);
and U6761 (N_6761,N_2183,N_4063);
nor U6762 (N_6762,N_2258,N_4630);
nand U6763 (N_6763,N_253,N_3293);
and U6764 (N_6764,N_3546,N_1817);
nor U6765 (N_6765,N_2701,N_4834);
nor U6766 (N_6766,N_1053,N_1319);
nor U6767 (N_6767,N_4335,N_592);
xor U6768 (N_6768,N_1991,N_3083);
nor U6769 (N_6769,N_4057,N_2777);
xor U6770 (N_6770,N_3877,N_4416);
nor U6771 (N_6771,N_2080,N_2171);
nor U6772 (N_6772,N_1192,N_4521);
xor U6773 (N_6773,N_4384,N_1654);
xnor U6774 (N_6774,N_4441,N_4445);
or U6775 (N_6775,N_4052,N_739);
nor U6776 (N_6776,N_1607,N_4238);
nor U6777 (N_6777,N_2269,N_165);
nand U6778 (N_6778,N_663,N_2319);
nor U6779 (N_6779,N_4703,N_4797);
or U6780 (N_6780,N_1896,N_2697);
nand U6781 (N_6781,N_932,N_2275);
or U6782 (N_6782,N_3061,N_4435);
nand U6783 (N_6783,N_4629,N_2569);
or U6784 (N_6784,N_480,N_850);
nand U6785 (N_6785,N_3655,N_2750);
nand U6786 (N_6786,N_3851,N_3470);
xnor U6787 (N_6787,N_244,N_3507);
or U6788 (N_6788,N_1886,N_3434);
nor U6789 (N_6789,N_3917,N_921);
and U6790 (N_6790,N_922,N_1761);
and U6791 (N_6791,N_3861,N_3815);
xnor U6792 (N_6792,N_1253,N_2351);
or U6793 (N_6793,N_4062,N_3584);
xnor U6794 (N_6794,N_2191,N_765);
or U6795 (N_6795,N_297,N_1394);
and U6796 (N_6796,N_4596,N_2749);
xnor U6797 (N_6797,N_2660,N_2714);
or U6798 (N_6798,N_4013,N_3500);
and U6799 (N_6799,N_4960,N_3970);
xnor U6800 (N_6800,N_2283,N_3898);
xnor U6801 (N_6801,N_693,N_2842);
nor U6802 (N_6802,N_4653,N_2602);
nand U6803 (N_6803,N_1191,N_2042);
and U6804 (N_6804,N_4241,N_2589);
or U6805 (N_6805,N_4578,N_2534);
nand U6806 (N_6806,N_2365,N_1960);
xnor U6807 (N_6807,N_3849,N_152);
nor U6808 (N_6808,N_4955,N_3002);
nand U6809 (N_6809,N_314,N_1510);
nor U6810 (N_6810,N_82,N_882);
nor U6811 (N_6811,N_2649,N_2298);
and U6812 (N_6812,N_3035,N_2672);
and U6813 (N_6813,N_3134,N_3457);
nor U6814 (N_6814,N_1613,N_3920);
or U6815 (N_6815,N_492,N_135);
nand U6816 (N_6816,N_2299,N_1762);
nand U6817 (N_6817,N_4591,N_4913);
and U6818 (N_6818,N_415,N_1339);
xnor U6819 (N_6819,N_2097,N_272);
and U6820 (N_6820,N_3039,N_3679);
and U6821 (N_6821,N_2578,N_1321);
xor U6822 (N_6822,N_2486,N_104);
nor U6823 (N_6823,N_4529,N_4994);
nand U6824 (N_6824,N_3178,N_3857);
nand U6825 (N_6825,N_1593,N_2193);
and U6826 (N_6826,N_4642,N_2817);
xnor U6827 (N_6827,N_21,N_4823);
or U6828 (N_6828,N_2783,N_606);
or U6829 (N_6829,N_1176,N_2596);
nor U6830 (N_6830,N_1848,N_1208);
nor U6831 (N_6831,N_3303,N_4463);
nand U6832 (N_6832,N_4701,N_3318);
nand U6833 (N_6833,N_3940,N_3271);
nand U6834 (N_6834,N_4976,N_4172);
and U6835 (N_6835,N_1952,N_4741);
or U6836 (N_6836,N_3539,N_639);
nand U6837 (N_6837,N_38,N_3310);
or U6838 (N_6838,N_3746,N_1461);
and U6839 (N_6839,N_3205,N_345);
and U6840 (N_6840,N_2999,N_4821);
or U6841 (N_6841,N_3086,N_4571);
nand U6842 (N_6842,N_4234,N_2599);
xnor U6843 (N_6843,N_3294,N_4207);
nor U6844 (N_6844,N_527,N_1400);
nand U6845 (N_6845,N_1539,N_4340);
xnor U6846 (N_6846,N_1299,N_2930);
and U6847 (N_6847,N_372,N_2103);
and U6848 (N_6848,N_220,N_669);
nor U6849 (N_6849,N_3631,N_4413);
or U6850 (N_6850,N_2843,N_3496);
xor U6851 (N_6851,N_434,N_1193);
and U6852 (N_6852,N_348,N_3254);
or U6853 (N_6853,N_3148,N_2900);
and U6854 (N_6854,N_3328,N_497);
xor U6855 (N_6855,N_187,N_2977);
nand U6856 (N_6856,N_3722,N_2935);
nor U6857 (N_6857,N_780,N_696);
or U6858 (N_6858,N_1686,N_2583);
xnor U6859 (N_6859,N_2563,N_2825);
and U6860 (N_6860,N_3179,N_1480);
nor U6861 (N_6861,N_832,N_4829);
nand U6862 (N_6862,N_3701,N_586);
nand U6863 (N_6863,N_3975,N_3104);
and U6864 (N_6864,N_4663,N_3779);
or U6865 (N_6865,N_4814,N_736);
xnor U6866 (N_6866,N_3531,N_233);
nand U6867 (N_6867,N_1436,N_1444);
or U6868 (N_6868,N_966,N_2537);
xor U6869 (N_6869,N_853,N_1466);
or U6870 (N_6870,N_417,N_2361);
or U6871 (N_6871,N_4775,N_603);
or U6872 (N_6872,N_1957,N_369);
and U6873 (N_6873,N_1125,N_4843);
or U6874 (N_6874,N_4815,N_4595);
or U6875 (N_6875,N_1756,N_2180);
nor U6876 (N_6876,N_3230,N_645);
nand U6877 (N_6877,N_489,N_661);
nand U6878 (N_6878,N_2239,N_296);
xor U6879 (N_6879,N_2342,N_1269);
or U6880 (N_6880,N_3649,N_1861);
nand U6881 (N_6881,N_514,N_1351);
nand U6882 (N_6882,N_1777,N_3945);
xor U6883 (N_6883,N_3755,N_4324);
nor U6884 (N_6884,N_680,N_2451);
nor U6885 (N_6885,N_309,N_4924);
and U6886 (N_6886,N_940,N_1452);
or U6887 (N_6887,N_3858,N_4058);
xor U6888 (N_6888,N_4883,N_3233);
or U6889 (N_6889,N_768,N_1166);
xor U6890 (N_6890,N_2208,N_2664);
or U6891 (N_6891,N_912,N_1360);
nand U6892 (N_6892,N_3068,N_1897);
xor U6893 (N_6893,N_2521,N_3512);
or U6894 (N_6894,N_3880,N_1859);
nor U6895 (N_6895,N_3260,N_1702);
nand U6896 (N_6896,N_1245,N_1804);
xor U6897 (N_6897,N_991,N_487);
or U6898 (N_6898,N_4700,N_1933);
nor U6899 (N_6899,N_1453,N_2118);
and U6900 (N_6900,N_4118,N_1729);
nand U6901 (N_6901,N_640,N_508);
nor U6902 (N_6902,N_4184,N_2038);
xor U6903 (N_6903,N_3728,N_42);
nor U6904 (N_6904,N_1726,N_189);
nand U6905 (N_6905,N_2614,N_1617);
nand U6906 (N_6906,N_2866,N_2815);
or U6907 (N_6907,N_199,N_1730);
and U6908 (N_6908,N_252,N_4224);
and U6909 (N_6909,N_2798,N_2590);
and U6910 (N_6910,N_4833,N_738);
xor U6911 (N_6911,N_2461,N_3964);
nor U6912 (N_6912,N_4620,N_1993);
nand U6913 (N_6913,N_4604,N_2369);
and U6914 (N_6914,N_1397,N_1393);
and U6915 (N_6915,N_1873,N_4933);
and U6916 (N_6916,N_1563,N_2519);
nor U6917 (N_6917,N_4782,N_3830);
nand U6918 (N_6918,N_978,N_1114);
or U6919 (N_6919,N_328,N_4078);
nand U6920 (N_6920,N_3670,N_290);
or U6921 (N_6921,N_1968,N_4041);
and U6922 (N_6922,N_4929,N_2950);
and U6923 (N_6923,N_2176,N_451);
or U6924 (N_6924,N_1440,N_1739);
nand U6925 (N_6925,N_4892,N_3604);
or U6926 (N_6926,N_4884,N_800);
nor U6927 (N_6927,N_1696,N_1965);
or U6928 (N_6928,N_3415,N_3676);
nor U6929 (N_6929,N_3460,N_37);
or U6930 (N_6930,N_3401,N_1025);
nor U6931 (N_6931,N_4851,N_3129);
and U6932 (N_6932,N_873,N_2316);
nand U6933 (N_6933,N_94,N_2028);
nand U6934 (N_6934,N_4015,N_4606);
nor U6935 (N_6935,N_98,N_2759);
and U6936 (N_6936,N_1771,N_212);
or U6937 (N_6937,N_2356,N_3270);
and U6938 (N_6938,N_4176,N_585);
nand U6939 (N_6939,N_2565,N_4235);
xor U6940 (N_6940,N_2531,N_3662);
and U6941 (N_6941,N_2084,N_3571);
xnor U6942 (N_6942,N_3860,N_1008);
and U6943 (N_6943,N_1962,N_295);
nor U6944 (N_6944,N_583,N_3760);
nor U6945 (N_6945,N_1767,N_2869);
xnor U6946 (N_6946,N_528,N_1104);
xor U6947 (N_6947,N_2061,N_485);
nor U6948 (N_6948,N_501,N_2020);
nand U6949 (N_6949,N_347,N_1263);
and U6950 (N_6950,N_4139,N_1061);
or U6951 (N_6951,N_4953,N_3084);
nor U6952 (N_6952,N_379,N_1361);
xnor U6953 (N_6953,N_4517,N_56);
and U6954 (N_6954,N_4046,N_1090);
or U6955 (N_6955,N_4370,N_1216);
nand U6956 (N_6956,N_1884,N_1969);
or U6957 (N_6957,N_3257,N_4217);
and U6958 (N_6958,N_2292,N_599);
nor U6959 (N_6959,N_3621,N_4481);
nand U6960 (N_6960,N_321,N_3422);
nand U6961 (N_6961,N_396,N_268);
nand U6962 (N_6962,N_4873,N_1223);
or U6963 (N_6963,N_177,N_2344);
and U6964 (N_6964,N_1092,N_2166);
or U6965 (N_6965,N_798,N_1955);
nor U6966 (N_6966,N_4029,N_1858);
nor U6967 (N_6967,N_4939,N_4844);
nand U6968 (N_6968,N_1354,N_493);
and U6969 (N_6969,N_2001,N_4305);
nor U6970 (N_6970,N_4547,N_3239);
xor U6971 (N_6971,N_1141,N_475);
or U6972 (N_6972,N_2403,N_3473);
nor U6973 (N_6973,N_3660,N_1259);
nor U6974 (N_6974,N_4510,N_622);
nand U6975 (N_6975,N_4932,N_3552);
nand U6976 (N_6976,N_326,N_1338);
or U6977 (N_6977,N_4179,N_1665);
nor U6978 (N_6978,N_4682,N_1085);
nand U6979 (N_6979,N_1435,N_4017);
xnor U6980 (N_6980,N_1905,N_4585);
and U6981 (N_6981,N_3037,N_206);
nor U6982 (N_6982,N_2987,N_728);
and U6983 (N_6983,N_4824,N_1901);
or U6984 (N_6984,N_675,N_4436);
or U6985 (N_6985,N_2886,N_4074);
and U6986 (N_6986,N_660,N_248);
nor U6987 (N_6987,N_2764,N_4940);
and U6988 (N_6988,N_3371,N_3908);
and U6989 (N_6989,N_202,N_2915);
nand U6990 (N_6990,N_3871,N_896);
xnor U6991 (N_6991,N_2506,N_2196);
or U6992 (N_6992,N_1731,N_3856);
or U6993 (N_6993,N_4244,N_3394);
and U6994 (N_6994,N_3355,N_4407);
or U6995 (N_6995,N_469,N_909);
nor U6996 (N_6996,N_2844,N_1374);
nor U6997 (N_6997,N_2289,N_2409);
xnor U6998 (N_6998,N_3360,N_1712);
nor U6999 (N_6999,N_3783,N_391);
nor U7000 (N_7000,N_4200,N_2287);
or U7001 (N_7001,N_809,N_4453);
xor U7002 (N_7002,N_2278,N_141);
or U7003 (N_7003,N_521,N_327);
xnor U7004 (N_7004,N_237,N_1382);
or U7005 (N_7005,N_52,N_4282);
and U7006 (N_7006,N_2627,N_218);
or U7007 (N_7007,N_3010,N_4491);
xor U7008 (N_7008,N_2792,N_4957);
nand U7009 (N_7009,N_2570,N_4479);
nand U7010 (N_7010,N_442,N_3513);
nor U7011 (N_7011,N_397,N_1753);
nor U7012 (N_7012,N_3418,N_2428);
nor U7013 (N_7013,N_4890,N_3354);
and U7014 (N_7014,N_2479,N_4150);
xor U7015 (N_7015,N_4274,N_3568);
or U7016 (N_7016,N_2415,N_3636);
and U7017 (N_7017,N_2883,N_1902);
xor U7018 (N_7018,N_3242,N_2530);
and U7019 (N_7019,N_3029,N_1610);
nor U7020 (N_7020,N_4196,N_1797);
or U7021 (N_7021,N_2374,N_5);
nor U7022 (N_7022,N_3596,N_2297);
nand U7023 (N_7023,N_633,N_2373);
or U7024 (N_7024,N_3840,N_3414);
or U7025 (N_7025,N_380,N_2989);
nor U7026 (N_7026,N_3167,N_4350);
nor U7027 (N_7027,N_3327,N_2368);
and U7028 (N_7028,N_3835,N_1644);
and U7029 (N_7029,N_948,N_4470);
nand U7030 (N_7030,N_2735,N_3806);
xor U7031 (N_7031,N_1845,N_8);
and U7032 (N_7032,N_944,N_1315);
nor U7033 (N_7033,N_828,N_3052);
and U7034 (N_7034,N_715,N_3071);
or U7035 (N_7035,N_1992,N_2527);
or U7036 (N_7036,N_3105,N_2346);
and U7037 (N_7037,N_86,N_2658);
xor U7038 (N_7038,N_2763,N_3749);
xor U7039 (N_7039,N_338,N_4684);
nor U7040 (N_7040,N_2593,N_2579);
nand U7041 (N_7041,N_1605,N_3014);
nor U7042 (N_7042,N_4339,N_4875);
or U7043 (N_7043,N_419,N_3461);
or U7044 (N_7044,N_2203,N_2443);
nand U7045 (N_7045,N_4977,N_1850);
nor U7046 (N_7046,N_936,N_90);
and U7047 (N_7047,N_1936,N_2387);
or U7048 (N_7048,N_1457,N_4562);
xnor U7049 (N_7049,N_1514,N_2902);
xnor U7050 (N_7050,N_4381,N_3736);
nor U7051 (N_7051,N_2031,N_3198);
or U7052 (N_7052,N_3016,N_496);
and U7053 (N_7053,N_4826,N_1666);
nor U7054 (N_7054,N_2516,N_1874);
xnor U7055 (N_7055,N_1647,N_3274);
or U7056 (N_7056,N_175,N_1377);
and U7057 (N_7057,N_4021,N_4950);
nor U7058 (N_7058,N_1006,N_2607);
nand U7059 (N_7059,N_3091,N_4902);
nor U7060 (N_7060,N_624,N_1409);
or U7061 (N_7061,N_3564,N_2148);
nand U7062 (N_7062,N_242,N_1406);
nor U7063 (N_7063,N_4802,N_408);
xnor U7064 (N_7064,N_1519,N_1026);
xor U7065 (N_7065,N_1020,N_3521);
and U7066 (N_7066,N_1669,N_3601);
or U7067 (N_7067,N_1120,N_4563);
and U7068 (N_7068,N_4963,N_3530);
and U7069 (N_7069,N_2460,N_1169);
nand U7070 (N_7070,N_2943,N_1923);
nor U7071 (N_7071,N_2427,N_802);
xor U7072 (N_7072,N_4140,N_2511);
nor U7073 (N_7073,N_713,N_464);
or U7074 (N_7074,N_1843,N_636);
and U7075 (N_7075,N_59,N_3184);
or U7076 (N_7076,N_981,N_2495);
and U7077 (N_7077,N_3922,N_3395);
xor U7078 (N_7078,N_1618,N_2850);
or U7079 (N_7079,N_4958,N_4351);
xnor U7080 (N_7080,N_2322,N_2744);
nand U7081 (N_7081,N_3204,N_2115);
xor U7082 (N_7082,N_3049,N_4639);
nand U7083 (N_7083,N_1798,N_2076);
nand U7084 (N_7084,N_1950,N_568);
or U7085 (N_7085,N_2969,N_2523);
nor U7086 (N_7086,N_540,N_785);
nand U7087 (N_7087,N_857,N_2378);
nand U7088 (N_7088,N_4259,N_2437);
nand U7089 (N_7089,N_2228,N_1978);
and U7090 (N_7090,N_2195,N_246);
nor U7091 (N_7091,N_4272,N_2548);
xor U7092 (N_7092,N_1265,N_1506);
or U7093 (N_7093,N_4750,N_3100);
nand U7094 (N_7094,N_4168,N_4907);
xnor U7095 (N_7095,N_1690,N_3588);
nand U7096 (N_7096,N_3130,N_430);
or U7097 (N_7097,N_4789,N_2884);
xnor U7098 (N_7098,N_1754,N_3550);
nor U7099 (N_7099,N_1588,N_2532);
nand U7100 (N_7100,N_216,N_1926);
nor U7101 (N_7101,N_414,N_2335);
and U7102 (N_7102,N_1524,N_370);
nand U7103 (N_7103,N_1684,N_2090);
nor U7104 (N_7104,N_2394,N_4767);
or U7105 (N_7105,N_4754,N_4651);
and U7106 (N_7106,N_463,N_4333);
or U7107 (N_7107,N_4612,N_2515);
nand U7108 (N_7108,N_3003,N_3359);
and U7109 (N_7109,N_193,N_1311);
nand U7110 (N_7110,N_3790,N_576);
nand U7111 (N_7111,N_3490,N_1785);
or U7112 (N_7112,N_481,N_468);
and U7113 (N_7113,N_1103,N_2053);
xor U7114 (N_7114,N_886,N_2014);
and U7115 (N_7115,N_4947,N_19);
xor U7116 (N_7116,N_821,N_3266);
nand U7117 (N_7117,N_4132,N_3960);
and U7118 (N_7118,N_3999,N_1056);
and U7119 (N_7119,N_2050,N_46);
xnor U7120 (N_7120,N_4699,N_3017);
or U7121 (N_7121,N_1769,N_2689);
xor U7122 (N_7122,N_389,N_4603);
nand U7123 (N_7123,N_166,N_2165);
nor U7124 (N_7124,N_1238,N_3038);
or U7125 (N_7125,N_2158,N_2976);
nor U7126 (N_7126,N_1112,N_4199);
xnor U7127 (N_7127,N_3339,N_1147);
and U7128 (N_7128,N_889,N_236);
xor U7129 (N_7129,N_3727,N_1295);
nor U7130 (N_7130,N_2009,N_240);
nor U7131 (N_7131,N_3309,N_1912);
nor U7132 (N_7132,N_1446,N_2959);
or U7133 (N_7133,N_732,N_4387);
xnor U7134 (N_7134,N_4648,N_3306);
xor U7135 (N_7135,N_3931,N_3776);
xnor U7136 (N_7136,N_2436,N_3544);
or U7137 (N_7137,N_916,N_1331);
or U7138 (N_7138,N_2027,N_2919);
nand U7139 (N_7139,N_1584,N_3203);
xnor U7140 (N_7140,N_254,N_840);
or U7141 (N_7141,N_4523,N_2535);
and U7142 (N_7142,N_2698,N_534);
nand U7143 (N_7143,N_3244,N_4185);
nand U7144 (N_7144,N_3593,N_3892);
and U7145 (N_7145,N_4886,N_1108);
nand U7146 (N_7146,N_870,N_217);
and U7147 (N_7147,N_1472,N_2149);
and U7148 (N_7148,N_1984,N_2968);
nand U7149 (N_7149,N_4623,N_1561);
or U7150 (N_7150,N_2072,N_465);
or U7151 (N_7151,N_3853,N_3793);
nand U7152 (N_7152,N_1096,N_2420);
and U7153 (N_7153,N_4101,N_2960);
xnor U7154 (N_7154,N_2332,N_1567);
xnor U7155 (N_7155,N_1747,N_1362);
or U7156 (N_7156,N_2956,N_2075);
xor U7157 (N_7157,N_1010,N_3015);
nand U7158 (N_7158,N_343,N_4091);
nand U7159 (N_7159,N_79,N_4175);
and U7160 (N_7160,N_263,N_1128);
or U7161 (N_7161,N_3110,N_4548);
and U7162 (N_7162,N_1611,N_3687);
nand U7163 (N_7163,N_764,N_2741);
or U7164 (N_7164,N_734,N_4511);
and U7165 (N_7165,N_4661,N_3101);
nand U7166 (N_7166,N_1199,N_590);
and U7167 (N_7167,N_4268,N_3523);
xnor U7168 (N_7168,N_4226,N_3803);
and U7169 (N_7169,N_1075,N_3435);
nand U7170 (N_7170,N_3948,N_2760);
xor U7171 (N_7171,N_3902,N_3985);
xnor U7172 (N_7172,N_763,N_3977);
or U7173 (N_7173,N_1097,N_3569);
or U7174 (N_7174,N_3305,N_4163);
nand U7175 (N_7175,N_225,N_4414);
or U7176 (N_7176,N_3536,N_4284);
xor U7177 (N_7177,N_2325,N_3638);
nand U7178 (N_7178,N_1682,N_500);
xnor U7179 (N_7179,N_3572,N_1200);
nand U7180 (N_7180,N_2718,N_767);
xor U7181 (N_7181,N_302,N_2309);
nand U7182 (N_7182,N_4972,N_837);
and U7183 (N_7183,N_2670,N_1455);
nand U7184 (N_7184,N_2045,N_4628);
and U7185 (N_7185,N_4341,N_3688);
nor U7186 (N_7186,N_1721,N_878);
or U7187 (N_7187,N_40,N_4765);
or U7188 (N_7188,N_1872,N_1052);
or U7189 (N_7189,N_4203,N_980);
xor U7190 (N_7190,N_1782,N_758);
or U7191 (N_7191,N_949,N_3724);
nor U7192 (N_7192,N_4816,N_3652);
or U7193 (N_7193,N_976,N_2693);
xor U7194 (N_7194,N_4966,N_3642);
and U7195 (N_7195,N_3048,N_4856);
or U7196 (N_7196,N_3713,N_1161);
or U7197 (N_7197,N_1133,N_22);
and U7198 (N_7198,N_992,N_4981);
nand U7199 (N_7199,N_1091,N_2876);
nand U7200 (N_7200,N_1687,N_3419);
nor U7201 (N_7201,N_935,N_4035);
nand U7202 (N_7202,N_129,N_3151);
xor U7203 (N_7203,N_3142,N_3480);
xnor U7204 (N_7204,N_4086,N_1709);
or U7205 (N_7205,N_4887,N_3124);
or U7206 (N_7206,N_3519,N_3367);
and U7207 (N_7207,N_621,N_2406);
and U7208 (N_7208,N_1336,N_2337);
nand U7209 (N_7209,N_3196,N_1036);
or U7210 (N_7210,N_2112,N_512);
nor U7211 (N_7211,N_4131,N_1407);
xor U7212 (N_7212,N_865,N_3384);
or U7213 (N_7213,N_3540,N_1650);
and U7214 (N_7214,N_4660,N_1456);
and U7215 (N_7215,N_4812,N_2044);
or U7216 (N_7216,N_4178,N_4173);
xnor U7217 (N_7217,N_1310,N_4283);
and U7218 (N_7218,N_550,N_1770);
or U7219 (N_7219,N_1838,N_3033);
xnor U7220 (N_7220,N_4354,N_4786);
xnor U7221 (N_7221,N_3410,N_2410);
or U7222 (N_7222,N_1934,N_448);
and U7223 (N_7223,N_4451,N_511);
nand U7224 (N_7224,N_721,N_4392);
nor U7225 (N_7225,N_619,N_2770);
nand U7226 (N_7226,N_1887,N_3006);
nand U7227 (N_7227,N_4325,N_3941);
nand U7228 (N_7228,N_4990,N_3041);
xor U7229 (N_7229,N_4607,N_4388);
nand U7230 (N_7230,N_4554,N_4276);
xnor U7231 (N_7231,N_494,N_3729);
or U7232 (N_7232,N_3547,N_1228);
or U7233 (N_7233,N_884,N_1347);
or U7234 (N_7234,N_4615,N_2859);
nand U7235 (N_7235,N_1039,N_1264);
or U7236 (N_7236,N_3897,N_1140);
and U7237 (N_7237,N_4279,N_1854);
and U7238 (N_7238,N_2469,N_2060);
nand U7239 (N_7239,N_2892,N_3868);
or U7240 (N_7240,N_3177,N_24);
xnor U7241 (N_7241,N_1165,N_62);
and U7242 (N_7242,N_4331,N_2933);
nor U7243 (N_7243,N_4687,N_2123);
nand U7244 (N_7244,N_2800,N_4122);
nand U7245 (N_7245,N_3792,N_2101);
and U7246 (N_7246,N_4288,N_3672);
xor U7247 (N_7247,N_1232,N_3748);
nand U7248 (N_7248,N_2577,N_1996);
nor U7249 (N_7249,N_2941,N_1342);
xnor U7250 (N_7250,N_2130,N_1869);
xor U7251 (N_7251,N_4785,N_3836);
nor U7252 (N_7252,N_4398,N_3445);
xor U7253 (N_7253,N_3805,N_1734);
nand U7254 (N_7254,N_1627,N_2088);
nand U7255 (N_7255,N_1417,N_1293);
and U7256 (N_7256,N_3695,N_1027);
nor U7257 (N_7257,N_1368,N_4499);
nand U7258 (N_7258,N_668,N_2538);
nand U7259 (N_7259,N_1494,N_1909);
nand U7260 (N_7260,N_2547,N_3467);
nand U7261 (N_7261,N_2136,N_3751);
or U7262 (N_7262,N_1808,N_3577);
xnor U7263 (N_7263,N_2231,N_1662);
xor U7264 (N_7264,N_3509,N_2771);
or U7265 (N_7265,N_4739,N_1663);
nand U7266 (N_7266,N_4921,N_4733);
xnor U7267 (N_7267,N_2832,N_729);
nor U7268 (N_7268,N_2618,N_1241);
and U7269 (N_7269,N_1749,N_3448);
nor U7270 (N_7270,N_4784,N_3095);
xnor U7271 (N_7271,N_1402,N_845);
xor U7272 (N_7272,N_1340,N_3846);
nor U7273 (N_7273,N_1925,N_1738);
or U7274 (N_7274,N_80,N_3620);
xnor U7275 (N_7275,N_1773,N_2913);
xor U7276 (N_7276,N_3150,N_0);
nand U7277 (N_7277,N_4488,N_1830);
xnor U7278 (N_7278,N_1080,N_4042);
and U7279 (N_7279,N_3951,N_972);
xor U7280 (N_7280,N_3563,N_4158);
xnor U7281 (N_7281,N_1005,N_3969);
and U7282 (N_7282,N_3489,N_3301);
nand U7283 (N_7283,N_1033,N_2280);
or U7284 (N_7284,N_3082,N_319);
xnor U7285 (N_7285,N_3459,N_846);
or U7286 (N_7286,N_3921,N_3113);
nor U7287 (N_7287,N_1148,N_4774);
xor U7288 (N_7288,N_201,N_2533);
xnor U7289 (N_7289,N_1212,N_2721);
or U7290 (N_7290,N_65,N_3570);
nand U7291 (N_7291,N_4442,N_140);
nand U7292 (N_7292,N_1864,N_3768);
xnor U7293 (N_7293,N_3363,N_3152);
or U7294 (N_7294,N_4880,N_4093);
or U7295 (N_7295,N_4457,N_1878);
nor U7296 (N_7296,N_318,N_1835);
nand U7297 (N_7297,N_2068,N_1717);
and U7298 (N_7298,N_1447,N_2802);
and U7299 (N_7299,N_1187,N_1127);
nor U7300 (N_7300,N_1903,N_2567);
xnor U7301 (N_7301,N_4310,N_382);
and U7302 (N_7302,N_4997,N_2818);
or U7303 (N_7303,N_9,N_1370);
xnor U7304 (N_7304,N_4493,N_1408);
and U7305 (N_7305,N_1706,N_2140);
xnor U7306 (N_7306,N_1553,N_2377);
nor U7307 (N_7307,N_2957,N_3915);
nor U7308 (N_7308,N_1719,N_4222);
nor U7309 (N_7309,N_2804,N_2453);
nor U7310 (N_7310,N_1651,N_2424);
and U7311 (N_7311,N_1535,N_830);
nor U7312 (N_7312,N_4635,N_2221);
nor U7313 (N_7313,N_2132,N_2864);
and U7314 (N_7314,N_751,N_4296);
or U7315 (N_7315,N_1692,N_4586);
nor U7316 (N_7316,N_1054,N_4024);
nand U7317 (N_7317,N_388,N_959);
nand U7318 (N_7318,N_2562,N_3825);
or U7319 (N_7319,N_1064,N_4191);
xnor U7320 (N_7320,N_4909,N_1134);
and U7321 (N_7321,N_3725,N_2143);
xnor U7322 (N_7322,N_1168,N_2251);
nand U7323 (N_7323,N_103,N_4117);
and U7324 (N_7324,N_3777,N_3413);
and U7325 (N_7325,N_4009,N_4583);
nor U7326 (N_7326,N_2768,N_2529);
xnor U7327 (N_7327,N_529,N_422);
or U7328 (N_7328,N_1004,N_1357);
nor U7329 (N_7329,N_2062,N_4311);
xor U7330 (N_7330,N_1899,N_3471);
nor U7331 (N_7331,N_1502,N_3211);
and U7332 (N_7332,N_51,N_1657);
nand U7333 (N_7333,N_930,N_4800);
nand U7334 (N_7334,N_1732,N_2756);
nor U7335 (N_7335,N_4729,N_3438);
and U7336 (N_7336,N_2949,N_807);
xnor U7337 (N_7337,N_1258,N_2666);
nand U7338 (N_7338,N_3937,N_3870);
xor U7339 (N_7339,N_2757,N_3667);
or U7340 (N_7340,N_2225,N_2192);
nand U7341 (N_7341,N_1578,N_3268);
nor U7342 (N_7342,N_359,N_2199);
xor U7343 (N_7343,N_262,N_1977);
nor U7344 (N_7344,N_867,N_3220);
xnor U7345 (N_7345,N_2640,N_1787);
nand U7346 (N_7346,N_3963,N_892);
and U7347 (N_7347,N_4555,N_4395);
nor U7348 (N_7348,N_516,N_1691);
xnor U7349 (N_7349,N_4944,N_4309);
and U7350 (N_7350,N_4779,N_2109);
nor U7351 (N_7351,N_3976,N_2738);
and U7352 (N_7352,N_2473,N_3659);
and U7353 (N_7353,N_4128,N_4693);
or U7354 (N_7354,N_1556,N_2380);
xnor U7355 (N_7355,N_3379,N_2412);
or U7356 (N_7356,N_4558,N_3616);
and U7357 (N_7357,N_3700,N_3499);
xor U7358 (N_7358,N_4289,N_2395);
and U7359 (N_7359,N_170,N_3472);
nor U7360 (N_7360,N_4134,N_2400);
and U7361 (N_7361,N_4149,N_3344);
nand U7362 (N_7362,N_1231,N_4270);
and U7363 (N_7363,N_530,N_4321);
or U7364 (N_7364,N_4751,N_4863);
nand U7365 (N_7365,N_158,N_3583);
and U7366 (N_7366,N_4242,N_192);
and U7367 (N_7367,N_801,N_4752);
nand U7368 (N_7368,N_1448,N_653);
nor U7369 (N_7369,N_4304,N_4212);
or U7370 (N_7370,N_3510,N_361);
xor U7371 (N_7371,N_1152,N_4);
and U7372 (N_7372,N_4543,N_1628);
nand U7373 (N_7373,N_4723,N_3280);
xnor U7374 (N_7374,N_4576,N_3721);
nor U7375 (N_7375,N_4329,N_3246);
nor U7376 (N_7376,N_2237,N_3276);
or U7377 (N_7377,N_928,N_3358);
and U7378 (N_7378,N_1700,N_1098);
or U7379 (N_7379,N_191,N_672);
xnor U7380 (N_7380,N_3942,N_294);
and U7381 (N_7381,N_3961,N_4581);
or U7382 (N_7382,N_1652,N_1522);
or U7383 (N_7383,N_2544,N_2606);
xnor U7384 (N_7384,N_4505,N_746);
nor U7385 (N_7385,N_28,N_4327);
or U7386 (N_7386,N_2071,N_2536);
nand U7387 (N_7387,N_4478,N_3098);
nand U7388 (N_7388,N_4415,N_1067);
and U7389 (N_7389,N_4927,N_4121);
xor U7390 (N_7390,N_4949,N_64);
and U7391 (N_7391,N_609,N_4181);
xor U7392 (N_7392,N_2928,N_2463);
nor U7393 (N_7393,N_1286,N_1170);
xnor U7394 (N_7394,N_2505,N_4243);
nand U7395 (N_7395,N_4727,N_4023);
nand U7396 (N_7396,N_1348,N_3699);
nor U7397 (N_7397,N_2317,N_4048);
xor U7398 (N_7398,N_3850,N_4871);
nor U7399 (N_7399,N_2877,N_310);
nand U7400 (N_7400,N_3073,N_547);
nand U7401 (N_7401,N_4780,N_4742);
or U7402 (N_7402,N_2707,N_3787);
or U7403 (N_7403,N_3195,N_926);
or U7404 (N_7404,N_282,N_730);
nand U7405 (N_7405,N_678,N_597);
nand U7406 (N_7406,N_1404,N_4634);
nand U7407 (N_7407,N_1115,N_2040);
and U7408 (N_7408,N_2185,N_168);
nor U7409 (N_7409,N_1465,N_3164);
nand U7410 (N_7410,N_2202,N_4348);
or U7411 (N_7411,N_1727,N_2218);
nand U7412 (N_7412,N_436,N_2034);
or U7413 (N_7413,N_2638,N_457);
and U7414 (N_7414,N_1011,N_2303);
and U7415 (N_7415,N_1755,N_2921);
or U7416 (N_7416,N_2425,N_4120);
and U7417 (N_7417,N_3559,N_1489);
nor U7418 (N_7418,N_1089,N_2716);
and U7419 (N_7419,N_2502,N_2496);
nand U7420 (N_7420,N_57,N_1723);
xor U7421 (N_7421,N_3936,N_4218);
and U7422 (N_7422,N_2483,N_97);
and U7423 (N_7423,N_3111,N_1226);
nor U7424 (N_7424,N_4611,N_3657);
nor U7425 (N_7425,N_4220,N_3299);
nor U7426 (N_7426,N_684,N_637);
nand U7427 (N_7427,N_946,N_4051);
or U7428 (N_7428,N_3780,N_4263);
nor U7429 (N_7429,N_117,N_4302);
nor U7430 (N_7430,N_4143,N_4082);
nand U7431 (N_7431,N_4198,N_3641);
xnor U7432 (N_7432,N_4697,N_1270);
or U7433 (N_7433,N_2250,N_4792);
nand U7434 (N_7434,N_3955,N_223);
or U7435 (N_7435,N_914,N_2120);
and U7436 (N_7436,N_4127,N_3990);
nand U7437 (N_7437,N_4138,N_775);
or U7438 (N_7438,N_1173,N_2457);
and U7439 (N_7439,N_162,N_3189);
or U7440 (N_7440,N_3040,N_2110);
xnor U7441 (N_7441,N_3334,N_4096);
and U7442 (N_7442,N_3252,N_3935);
or U7443 (N_7443,N_2630,N_4494);
and U7444 (N_7444,N_4019,N_3674);
nor U7445 (N_7445,N_2261,N_213);
or U7446 (N_7446,N_4714,N_4036);
and U7447 (N_7447,N_3210,N_2313);
and U7448 (N_7448,N_3185,N_3373);
and U7449 (N_7449,N_2588,N_3483);
nor U7450 (N_7450,N_2550,N_230);
nor U7451 (N_7451,N_1431,N_1081);
nor U7452 (N_7452,N_2811,N_4717);
nand U7453 (N_7453,N_4599,N_2168);
and U7454 (N_7454,N_4747,N_996);
nor U7455 (N_7455,N_1425,N_854);
xor U7456 (N_7456,N_1022,N_567);
nor U7457 (N_7457,N_4926,N_2679);
or U7458 (N_7458,N_3214,N_1418);
nand U7459 (N_7459,N_2634,N_1282);
nand U7460 (N_7460,N_1477,N_4299);
and U7461 (N_7461,N_1144,N_342);
xnor U7462 (N_7462,N_4498,N_2616);
nor U7463 (N_7463,N_1003,N_484);
nor U7464 (N_7464,N_2557,N_182);
nor U7465 (N_7465,N_458,N_2233);
nor U7466 (N_7466,N_1343,N_3452);
nor U7467 (N_7467,N_816,N_1225);
nand U7468 (N_7468,N_44,N_2758);
nor U7469 (N_7469,N_3291,N_1356);
xnor U7470 (N_7470,N_806,N_671);
nand U7471 (N_7471,N_4730,N_1517);
or U7472 (N_7472,N_554,N_1094);
xor U7473 (N_7473,N_1536,N_3376);
and U7474 (N_7474,N_1828,N_2863);
nand U7475 (N_7475,N_4475,N_910);
and U7476 (N_7476,N_2482,N_1158);
nor U7477 (N_7477,N_2285,N_114);
nor U7478 (N_7478,N_1778,N_1879);
nand U7479 (N_7479,N_3297,N_4726);
or U7480 (N_7480,N_1063,N_3064);
nand U7481 (N_7481,N_433,N_1525);
nor U7482 (N_7482,N_1602,N_3158);
nand U7483 (N_7483,N_3841,N_1812);
xor U7484 (N_7484,N_1632,N_4822);
or U7485 (N_7485,N_2454,N_2704);
nand U7486 (N_7486,N_2281,N_3678);
nand U7487 (N_7487,N_4043,N_1688);
or U7488 (N_7488,N_979,N_4632);
xor U7489 (N_7489,N_2029,N_2017);
or U7490 (N_7490,N_2156,N_2324);
nand U7491 (N_7491,N_848,N_3201);
nor U7492 (N_7492,N_988,N_126);
and U7493 (N_7493,N_504,N_2414);
nand U7494 (N_7494,N_3059,N_2004);
xnor U7495 (N_7495,N_4891,N_3289);
and U7496 (N_7496,N_3447,N_277);
xnor U7497 (N_7497,N_3056,N_125);
or U7498 (N_7498,N_3810,N_4870);
nand U7499 (N_7499,N_808,N_4819);
xnor U7500 (N_7500,N_4365,N_2144);
xnor U7501 (N_7501,N_634,N_1388);
nand U7502 (N_7502,N_4437,N_2844);
or U7503 (N_7503,N_992,N_473);
nand U7504 (N_7504,N_3860,N_4529);
or U7505 (N_7505,N_3046,N_1322);
or U7506 (N_7506,N_372,N_552);
xor U7507 (N_7507,N_4661,N_4602);
nand U7508 (N_7508,N_4191,N_2721);
or U7509 (N_7509,N_533,N_3889);
or U7510 (N_7510,N_1145,N_3608);
and U7511 (N_7511,N_1661,N_3359);
xor U7512 (N_7512,N_1922,N_1516);
nor U7513 (N_7513,N_3941,N_1636);
and U7514 (N_7514,N_16,N_1858);
and U7515 (N_7515,N_4363,N_3345);
xnor U7516 (N_7516,N_1267,N_4212);
nor U7517 (N_7517,N_3403,N_1888);
or U7518 (N_7518,N_3290,N_374);
or U7519 (N_7519,N_1511,N_4427);
and U7520 (N_7520,N_4381,N_741);
xor U7521 (N_7521,N_1441,N_2557);
nand U7522 (N_7522,N_3078,N_3243);
nor U7523 (N_7523,N_1302,N_3188);
nand U7524 (N_7524,N_3278,N_2731);
or U7525 (N_7525,N_550,N_4871);
or U7526 (N_7526,N_1603,N_390);
or U7527 (N_7527,N_2408,N_3045);
or U7528 (N_7528,N_4788,N_2826);
nor U7529 (N_7529,N_4570,N_2004);
nand U7530 (N_7530,N_1156,N_2673);
and U7531 (N_7531,N_2878,N_2660);
and U7532 (N_7532,N_4636,N_1527);
or U7533 (N_7533,N_2982,N_386);
or U7534 (N_7534,N_4335,N_2690);
or U7535 (N_7535,N_115,N_407);
nor U7536 (N_7536,N_4394,N_2308);
and U7537 (N_7537,N_166,N_2133);
nor U7538 (N_7538,N_3988,N_2410);
or U7539 (N_7539,N_3766,N_3490);
xnor U7540 (N_7540,N_3560,N_1522);
and U7541 (N_7541,N_2099,N_1455);
and U7542 (N_7542,N_4025,N_2132);
or U7543 (N_7543,N_1723,N_4875);
or U7544 (N_7544,N_815,N_3555);
xor U7545 (N_7545,N_3401,N_2165);
nor U7546 (N_7546,N_2099,N_3898);
nor U7547 (N_7547,N_759,N_4503);
or U7548 (N_7548,N_2332,N_2199);
nor U7549 (N_7549,N_1707,N_1006);
or U7550 (N_7550,N_1633,N_108);
xnor U7551 (N_7551,N_4438,N_4447);
nor U7552 (N_7552,N_779,N_2429);
and U7553 (N_7553,N_1230,N_1928);
nor U7554 (N_7554,N_853,N_1598);
nand U7555 (N_7555,N_233,N_2416);
nand U7556 (N_7556,N_2830,N_4035);
and U7557 (N_7557,N_3758,N_11);
or U7558 (N_7558,N_4459,N_753);
or U7559 (N_7559,N_3993,N_4351);
xor U7560 (N_7560,N_2751,N_2196);
nor U7561 (N_7561,N_560,N_4687);
xor U7562 (N_7562,N_3664,N_4115);
xnor U7563 (N_7563,N_297,N_2986);
nor U7564 (N_7564,N_350,N_2504);
xor U7565 (N_7565,N_1175,N_4200);
xor U7566 (N_7566,N_439,N_997);
xnor U7567 (N_7567,N_2488,N_178);
and U7568 (N_7568,N_2712,N_4638);
xor U7569 (N_7569,N_340,N_3094);
nor U7570 (N_7570,N_877,N_3396);
nor U7571 (N_7571,N_36,N_305);
nand U7572 (N_7572,N_3388,N_3142);
nand U7573 (N_7573,N_2536,N_3850);
nor U7574 (N_7574,N_701,N_1692);
xor U7575 (N_7575,N_2616,N_4111);
nor U7576 (N_7576,N_743,N_4489);
and U7577 (N_7577,N_590,N_3281);
xor U7578 (N_7578,N_266,N_2142);
and U7579 (N_7579,N_2094,N_2923);
xnor U7580 (N_7580,N_1347,N_4662);
or U7581 (N_7581,N_2129,N_3368);
and U7582 (N_7582,N_4485,N_2499);
and U7583 (N_7583,N_1836,N_2868);
nor U7584 (N_7584,N_1282,N_937);
xnor U7585 (N_7585,N_3465,N_3216);
xor U7586 (N_7586,N_4589,N_3301);
nor U7587 (N_7587,N_2033,N_1484);
xnor U7588 (N_7588,N_3823,N_4105);
xnor U7589 (N_7589,N_4777,N_53);
nand U7590 (N_7590,N_1610,N_3653);
and U7591 (N_7591,N_4407,N_551);
xnor U7592 (N_7592,N_3870,N_72);
nand U7593 (N_7593,N_2109,N_404);
nor U7594 (N_7594,N_3407,N_2155);
xnor U7595 (N_7595,N_4265,N_287);
nor U7596 (N_7596,N_4137,N_2404);
and U7597 (N_7597,N_1877,N_1192);
and U7598 (N_7598,N_4746,N_4381);
nor U7599 (N_7599,N_197,N_1967);
and U7600 (N_7600,N_1531,N_3053);
nor U7601 (N_7601,N_1011,N_181);
or U7602 (N_7602,N_2425,N_846);
or U7603 (N_7603,N_3320,N_3093);
or U7604 (N_7604,N_3026,N_2997);
xnor U7605 (N_7605,N_4855,N_2623);
and U7606 (N_7606,N_298,N_4807);
nand U7607 (N_7607,N_3553,N_1346);
nor U7608 (N_7608,N_14,N_808);
nand U7609 (N_7609,N_16,N_787);
and U7610 (N_7610,N_2481,N_294);
xnor U7611 (N_7611,N_1719,N_870);
xnor U7612 (N_7612,N_3374,N_505);
and U7613 (N_7613,N_2864,N_1278);
and U7614 (N_7614,N_2732,N_624);
xnor U7615 (N_7615,N_2677,N_3513);
and U7616 (N_7616,N_1582,N_570);
nor U7617 (N_7617,N_4948,N_427);
or U7618 (N_7618,N_1405,N_630);
nand U7619 (N_7619,N_443,N_1493);
nor U7620 (N_7620,N_2754,N_1038);
nand U7621 (N_7621,N_4972,N_2646);
or U7622 (N_7622,N_3253,N_4864);
xor U7623 (N_7623,N_41,N_4306);
nor U7624 (N_7624,N_4963,N_4054);
xor U7625 (N_7625,N_4353,N_3884);
nor U7626 (N_7626,N_2294,N_3396);
nor U7627 (N_7627,N_3649,N_3289);
nor U7628 (N_7628,N_3837,N_4448);
nand U7629 (N_7629,N_628,N_1336);
nor U7630 (N_7630,N_3607,N_2641);
nor U7631 (N_7631,N_803,N_167);
nand U7632 (N_7632,N_3333,N_3886);
xor U7633 (N_7633,N_2592,N_4196);
or U7634 (N_7634,N_522,N_2968);
nor U7635 (N_7635,N_4119,N_2385);
xnor U7636 (N_7636,N_3910,N_4552);
nor U7637 (N_7637,N_2487,N_576);
nor U7638 (N_7638,N_2057,N_2477);
nand U7639 (N_7639,N_3514,N_175);
nor U7640 (N_7640,N_353,N_27);
and U7641 (N_7641,N_4451,N_3086);
and U7642 (N_7642,N_4242,N_3791);
and U7643 (N_7643,N_1493,N_1913);
nand U7644 (N_7644,N_790,N_2095);
and U7645 (N_7645,N_2868,N_4213);
xnor U7646 (N_7646,N_1719,N_1880);
or U7647 (N_7647,N_4909,N_3120);
xor U7648 (N_7648,N_3708,N_919);
nand U7649 (N_7649,N_3221,N_1869);
nor U7650 (N_7650,N_2381,N_631);
nand U7651 (N_7651,N_3681,N_3483);
and U7652 (N_7652,N_124,N_3126);
xor U7653 (N_7653,N_3406,N_979);
nor U7654 (N_7654,N_1764,N_3187);
or U7655 (N_7655,N_2194,N_3802);
nand U7656 (N_7656,N_2434,N_2311);
xnor U7657 (N_7657,N_2708,N_43);
xnor U7658 (N_7658,N_3477,N_2472);
xor U7659 (N_7659,N_504,N_3674);
and U7660 (N_7660,N_775,N_4780);
or U7661 (N_7661,N_1908,N_389);
and U7662 (N_7662,N_3914,N_221);
nor U7663 (N_7663,N_3416,N_2955);
or U7664 (N_7664,N_1163,N_966);
xnor U7665 (N_7665,N_4630,N_2555);
nor U7666 (N_7666,N_1227,N_1882);
xnor U7667 (N_7667,N_541,N_1370);
and U7668 (N_7668,N_2506,N_4517);
xor U7669 (N_7669,N_693,N_2278);
or U7670 (N_7670,N_576,N_3855);
nor U7671 (N_7671,N_3304,N_4081);
and U7672 (N_7672,N_2998,N_3227);
xor U7673 (N_7673,N_2737,N_1607);
xnor U7674 (N_7674,N_2178,N_1925);
and U7675 (N_7675,N_2738,N_1060);
nand U7676 (N_7676,N_207,N_526);
and U7677 (N_7677,N_1618,N_4718);
nand U7678 (N_7678,N_2429,N_2207);
xnor U7679 (N_7679,N_194,N_233);
xnor U7680 (N_7680,N_3599,N_540);
nand U7681 (N_7681,N_196,N_689);
and U7682 (N_7682,N_1717,N_2883);
or U7683 (N_7683,N_2499,N_1190);
or U7684 (N_7684,N_1250,N_3314);
xnor U7685 (N_7685,N_2534,N_1174);
nor U7686 (N_7686,N_1286,N_2443);
and U7687 (N_7687,N_1577,N_3168);
and U7688 (N_7688,N_4367,N_4716);
or U7689 (N_7689,N_2971,N_3532);
nand U7690 (N_7690,N_3048,N_872);
nand U7691 (N_7691,N_2266,N_1588);
or U7692 (N_7692,N_232,N_4002);
or U7693 (N_7693,N_621,N_258);
xnor U7694 (N_7694,N_385,N_4953);
or U7695 (N_7695,N_3836,N_1428);
nor U7696 (N_7696,N_1302,N_938);
or U7697 (N_7697,N_4003,N_1870);
nand U7698 (N_7698,N_3913,N_3850);
nor U7699 (N_7699,N_4188,N_1353);
nor U7700 (N_7700,N_1892,N_4090);
xor U7701 (N_7701,N_3090,N_2601);
and U7702 (N_7702,N_1251,N_1938);
and U7703 (N_7703,N_2147,N_1840);
and U7704 (N_7704,N_3059,N_1906);
nor U7705 (N_7705,N_1190,N_1351);
and U7706 (N_7706,N_976,N_2601);
xor U7707 (N_7707,N_1010,N_562);
xor U7708 (N_7708,N_2394,N_1772);
nand U7709 (N_7709,N_4273,N_2327);
nor U7710 (N_7710,N_1499,N_4955);
xor U7711 (N_7711,N_1837,N_2372);
nand U7712 (N_7712,N_571,N_393);
xnor U7713 (N_7713,N_4741,N_1307);
nand U7714 (N_7714,N_2194,N_3562);
nor U7715 (N_7715,N_4001,N_3199);
nand U7716 (N_7716,N_2603,N_1423);
and U7717 (N_7717,N_1438,N_2757);
and U7718 (N_7718,N_3736,N_3204);
or U7719 (N_7719,N_3000,N_3610);
nor U7720 (N_7720,N_4427,N_1451);
or U7721 (N_7721,N_3105,N_2432);
nor U7722 (N_7722,N_2401,N_796);
nand U7723 (N_7723,N_3592,N_891);
nand U7724 (N_7724,N_4451,N_4564);
or U7725 (N_7725,N_3133,N_3179);
xnor U7726 (N_7726,N_408,N_612);
or U7727 (N_7727,N_1698,N_3553);
nand U7728 (N_7728,N_3476,N_675);
nor U7729 (N_7729,N_64,N_2284);
nand U7730 (N_7730,N_4945,N_3866);
and U7731 (N_7731,N_1698,N_2213);
xnor U7732 (N_7732,N_217,N_4225);
nor U7733 (N_7733,N_4336,N_3812);
xnor U7734 (N_7734,N_3855,N_1251);
or U7735 (N_7735,N_3354,N_3004);
nand U7736 (N_7736,N_2702,N_3618);
nor U7737 (N_7737,N_3347,N_2252);
nor U7738 (N_7738,N_3087,N_2880);
or U7739 (N_7739,N_3629,N_4330);
nor U7740 (N_7740,N_2227,N_3162);
xnor U7741 (N_7741,N_746,N_643);
nor U7742 (N_7742,N_4393,N_2782);
and U7743 (N_7743,N_704,N_1909);
or U7744 (N_7744,N_1505,N_2939);
or U7745 (N_7745,N_1893,N_1465);
nor U7746 (N_7746,N_3077,N_547);
or U7747 (N_7747,N_2785,N_1185);
and U7748 (N_7748,N_211,N_2926);
nor U7749 (N_7749,N_3289,N_2195);
and U7750 (N_7750,N_4953,N_4147);
xor U7751 (N_7751,N_3398,N_867);
nand U7752 (N_7752,N_4790,N_1138);
or U7753 (N_7753,N_4680,N_516);
xnor U7754 (N_7754,N_1757,N_3227);
or U7755 (N_7755,N_3108,N_4133);
or U7756 (N_7756,N_1238,N_610);
or U7757 (N_7757,N_802,N_1428);
and U7758 (N_7758,N_1276,N_3260);
xor U7759 (N_7759,N_1898,N_3144);
or U7760 (N_7760,N_4749,N_1099);
nand U7761 (N_7761,N_368,N_1960);
and U7762 (N_7762,N_2314,N_3754);
and U7763 (N_7763,N_2648,N_4974);
xor U7764 (N_7764,N_838,N_624);
or U7765 (N_7765,N_702,N_4924);
nand U7766 (N_7766,N_155,N_3659);
nand U7767 (N_7767,N_843,N_3775);
and U7768 (N_7768,N_3305,N_1297);
nand U7769 (N_7769,N_4798,N_4789);
nor U7770 (N_7770,N_1377,N_2955);
or U7771 (N_7771,N_1689,N_2275);
and U7772 (N_7772,N_2317,N_299);
nor U7773 (N_7773,N_1234,N_463);
xnor U7774 (N_7774,N_660,N_2359);
nor U7775 (N_7775,N_4280,N_3494);
nor U7776 (N_7776,N_4846,N_2679);
and U7777 (N_7777,N_1648,N_1874);
nand U7778 (N_7778,N_2266,N_4457);
xnor U7779 (N_7779,N_2074,N_1559);
and U7780 (N_7780,N_576,N_4990);
nand U7781 (N_7781,N_2025,N_1810);
xnor U7782 (N_7782,N_984,N_3079);
nor U7783 (N_7783,N_3446,N_352);
xor U7784 (N_7784,N_3294,N_1789);
xnor U7785 (N_7785,N_2549,N_4257);
or U7786 (N_7786,N_1563,N_4425);
xor U7787 (N_7787,N_801,N_964);
xor U7788 (N_7788,N_1197,N_4474);
xor U7789 (N_7789,N_452,N_859);
nor U7790 (N_7790,N_752,N_4524);
and U7791 (N_7791,N_909,N_846);
nand U7792 (N_7792,N_3418,N_3492);
xor U7793 (N_7793,N_3987,N_1253);
nor U7794 (N_7794,N_3015,N_637);
and U7795 (N_7795,N_1465,N_4302);
xnor U7796 (N_7796,N_3856,N_1882);
or U7797 (N_7797,N_1494,N_1502);
nor U7798 (N_7798,N_1280,N_4884);
nand U7799 (N_7799,N_179,N_4183);
nor U7800 (N_7800,N_889,N_3819);
or U7801 (N_7801,N_785,N_3562);
xor U7802 (N_7802,N_4521,N_3246);
nand U7803 (N_7803,N_3518,N_4500);
and U7804 (N_7804,N_4317,N_3753);
nand U7805 (N_7805,N_4252,N_877);
or U7806 (N_7806,N_147,N_1986);
nand U7807 (N_7807,N_2052,N_3147);
nor U7808 (N_7808,N_1329,N_99);
nand U7809 (N_7809,N_3881,N_2946);
xnor U7810 (N_7810,N_3777,N_525);
or U7811 (N_7811,N_4046,N_1022);
nand U7812 (N_7812,N_862,N_2246);
and U7813 (N_7813,N_3125,N_2214);
and U7814 (N_7814,N_2249,N_360);
or U7815 (N_7815,N_334,N_1157);
nor U7816 (N_7816,N_4549,N_3354);
nor U7817 (N_7817,N_4581,N_1529);
and U7818 (N_7818,N_1339,N_2949);
and U7819 (N_7819,N_4972,N_3045);
xnor U7820 (N_7820,N_1208,N_951);
xor U7821 (N_7821,N_4290,N_601);
or U7822 (N_7822,N_679,N_1465);
nor U7823 (N_7823,N_2754,N_2564);
nor U7824 (N_7824,N_3770,N_2634);
and U7825 (N_7825,N_764,N_3712);
nand U7826 (N_7826,N_1346,N_2842);
xnor U7827 (N_7827,N_3173,N_1998);
or U7828 (N_7828,N_4404,N_1551);
nor U7829 (N_7829,N_4546,N_207);
or U7830 (N_7830,N_1509,N_2070);
nor U7831 (N_7831,N_677,N_133);
or U7832 (N_7832,N_4142,N_2607);
and U7833 (N_7833,N_4832,N_1731);
nor U7834 (N_7834,N_2740,N_2587);
xor U7835 (N_7835,N_3693,N_4664);
nand U7836 (N_7836,N_3936,N_1037);
xor U7837 (N_7837,N_3623,N_3177);
nor U7838 (N_7838,N_1312,N_1065);
xor U7839 (N_7839,N_286,N_1736);
and U7840 (N_7840,N_854,N_4465);
or U7841 (N_7841,N_4170,N_3961);
nand U7842 (N_7842,N_963,N_4532);
and U7843 (N_7843,N_4685,N_389);
xnor U7844 (N_7844,N_3497,N_2910);
nand U7845 (N_7845,N_4622,N_2173);
and U7846 (N_7846,N_24,N_3753);
nand U7847 (N_7847,N_1037,N_2476);
nor U7848 (N_7848,N_2256,N_292);
nand U7849 (N_7849,N_4092,N_2542);
and U7850 (N_7850,N_4547,N_516);
nor U7851 (N_7851,N_811,N_3153);
and U7852 (N_7852,N_4315,N_2754);
nand U7853 (N_7853,N_3806,N_2295);
nor U7854 (N_7854,N_1974,N_3812);
and U7855 (N_7855,N_3934,N_1291);
nand U7856 (N_7856,N_4636,N_4179);
and U7857 (N_7857,N_2974,N_1116);
nor U7858 (N_7858,N_4843,N_3479);
or U7859 (N_7859,N_2094,N_2206);
and U7860 (N_7860,N_3329,N_3477);
nand U7861 (N_7861,N_4479,N_3791);
nand U7862 (N_7862,N_2326,N_3925);
nor U7863 (N_7863,N_4636,N_4176);
or U7864 (N_7864,N_1316,N_915);
nor U7865 (N_7865,N_405,N_4881);
and U7866 (N_7866,N_3606,N_674);
nor U7867 (N_7867,N_2032,N_2824);
or U7868 (N_7868,N_550,N_3255);
and U7869 (N_7869,N_2138,N_4412);
and U7870 (N_7870,N_1988,N_4167);
nand U7871 (N_7871,N_2501,N_2419);
or U7872 (N_7872,N_3121,N_2718);
or U7873 (N_7873,N_3223,N_1498);
xnor U7874 (N_7874,N_4964,N_606);
and U7875 (N_7875,N_1763,N_76);
or U7876 (N_7876,N_1780,N_2227);
and U7877 (N_7877,N_1939,N_1575);
nor U7878 (N_7878,N_3736,N_774);
and U7879 (N_7879,N_4255,N_4699);
or U7880 (N_7880,N_355,N_2686);
or U7881 (N_7881,N_4091,N_3992);
or U7882 (N_7882,N_3776,N_1350);
and U7883 (N_7883,N_3088,N_1261);
nor U7884 (N_7884,N_208,N_4250);
nand U7885 (N_7885,N_1793,N_1274);
nand U7886 (N_7886,N_4646,N_2123);
and U7887 (N_7887,N_4719,N_4627);
xor U7888 (N_7888,N_74,N_2119);
and U7889 (N_7889,N_153,N_3021);
and U7890 (N_7890,N_1497,N_2953);
or U7891 (N_7891,N_71,N_2730);
nor U7892 (N_7892,N_3937,N_2036);
xor U7893 (N_7893,N_111,N_2205);
or U7894 (N_7894,N_2624,N_4260);
xnor U7895 (N_7895,N_1442,N_4028);
or U7896 (N_7896,N_280,N_1030);
xnor U7897 (N_7897,N_1718,N_3954);
xnor U7898 (N_7898,N_1018,N_3864);
or U7899 (N_7899,N_713,N_3823);
nand U7900 (N_7900,N_3864,N_1079);
and U7901 (N_7901,N_2116,N_3058);
xnor U7902 (N_7902,N_2990,N_1716);
and U7903 (N_7903,N_4211,N_2443);
nor U7904 (N_7904,N_4710,N_1391);
nand U7905 (N_7905,N_2256,N_3671);
nor U7906 (N_7906,N_1630,N_1408);
and U7907 (N_7907,N_1647,N_4668);
and U7908 (N_7908,N_349,N_175);
or U7909 (N_7909,N_3777,N_1796);
nor U7910 (N_7910,N_2855,N_3896);
nand U7911 (N_7911,N_51,N_1328);
and U7912 (N_7912,N_3574,N_3443);
nor U7913 (N_7913,N_1152,N_3511);
nor U7914 (N_7914,N_4958,N_3955);
xor U7915 (N_7915,N_1507,N_3570);
nand U7916 (N_7916,N_1901,N_1189);
and U7917 (N_7917,N_3477,N_2931);
xor U7918 (N_7918,N_4984,N_806);
or U7919 (N_7919,N_2659,N_2596);
nor U7920 (N_7920,N_2062,N_291);
nand U7921 (N_7921,N_3520,N_3223);
xnor U7922 (N_7922,N_259,N_3726);
nor U7923 (N_7923,N_2579,N_751);
nor U7924 (N_7924,N_4103,N_4357);
xnor U7925 (N_7925,N_3364,N_1189);
xnor U7926 (N_7926,N_1043,N_420);
and U7927 (N_7927,N_2658,N_4850);
or U7928 (N_7928,N_65,N_3378);
nor U7929 (N_7929,N_3483,N_4246);
xnor U7930 (N_7930,N_1099,N_2460);
nand U7931 (N_7931,N_3807,N_751);
and U7932 (N_7932,N_1793,N_2587);
or U7933 (N_7933,N_3643,N_3807);
nand U7934 (N_7934,N_4547,N_1571);
nand U7935 (N_7935,N_530,N_4271);
nor U7936 (N_7936,N_2163,N_3018);
or U7937 (N_7937,N_3681,N_2786);
and U7938 (N_7938,N_534,N_2170);
nand U7939 (N_7939,N_969,N_1353);
nor U7940 (N_7940,N_3359,N_4679);
and U7941 (N_7941,N_3905,N_2248);
and U7942 (N_7942,N_1888,N_2475);
and U7943 (N_7943,N_3091,N_3875);
xnor U7944 (N_7944,N_1749,N_4583);
nand U7945 (N_7945,N_1666,N_31);
or U7946 (N_7946,N_2853,N_3915);
xnor U7947 (N_7947,N_4274,N_1251);
nand U7948 (N_7948,N_2777,N_2031);
and U7949 (N_7949,N_4578,N_2664);
nand U7950 (N_7950,N_2183,N_1060);
or U7951 (N_7951,N_4456,N_2678);
nor U7952 (N_7952,N_775,N_1085);
nand U7953 (N_7953,N_4538,N_1420);
or U7954 (N_7954,N_3345,N_4333);
xnor U7955 (N_7955,N_4873,N_485);
nor U7956 (N_7956,N_2482,N_353);
and U7957 (N_7957,N_573,N_3074);
nor U7958 (N_7958,N_3976,N_669);
or U7959 (N_7959,N_378,N_1284);
xor U7960 (N_7960,N_3496,N_3233);
and U7961 (N_7961,N_1760,N_4714);
and U7962 (N_7962,N_3989,N_94);
and U7963 (N_7963,N_2235,N_2076);
nand U7964 (N_7964,N_662,N_1298);
xnor U7965 (N_7965,N_203,N_4500);
nand U7966 (N_7966,N_4618,N_4791);
xor U7967 (N_7967,N_4620,N_1468);
and U7968 (N_7968,N_1742,N_103);
and U7969 (N_7969,N_577,N_4085);
nand U7970 (N_7970,N_3405,N_224);
nor U7971 (N_7971,N_2136,N_4679);
and U7972 (N_7972,N_4304,N_1775);
or U7973 (N_7973,N_416,N_4889);
nor U7974 (N_7974,N_1014,N_4960);
and U7975 (N_7975,N_1040,N_2812);
nand U7976 (N_7976,N_375,N_2919);
nor U7977 (N_7977,N_3133,N_1984);
and U7978 (N_7978,N_1134,N_1011);
xnor U7979 (N_7979,N_2941,N_4617);
or U7980 (N_7980,N_3929,N_432);
nor U7981 (N_7981,N_2081,N_595);
and U7982 (N_7982,N_3398,N_3586);
nor U7983 (N_7983,N_2925,N_3361);
and U7984 (N_7984,N_355,N_3260);
xnor U7985 (N_7985,N_3341,N_2444);
or U7986 (N_7986,N_396,N_2853);
and U7987 (N_7987,N_4688,N_2304);
nor U7988 (N_7988,N_148,N_3623);
nand U7989 (N_7989,N_4846,N_4529);
xor U7990 (N_7990,N_2686,N_2757);
nor U7991 (N_7991,N_4245,N_3105);
nor U7992 (N_7992,N_1764,N_906);
and U7993 (N_7993,N_849,N_3869);
or U7994 (N_7994,N_798,N_671);
and U7995 (N_7995,N_282,N_1126);
or U7996 (N_7996,N_2308,N_4602);
or U7997 (N_7997,N_2647,N_1038);
nand U7998 (N_7998,N_3463,N_4377);
nor U7999 (N_7999,N_2532,N_4006);
nand U8000 (N_8000,N_1974,N_1315);
nor U8001 (N_8001,N_776,N_156);
and U8002 (N_8002,N_1887,N_3494);
xnor U8003 (N_8003,N_321,N_755);
nor U8004 (N_8004,N_1153,N_4575);
and U8005 (N_8005,N_2434,N_2672);
or U8006 (N_8006,N_3292,N_441);
and U8007 (N_8007,N_4753,N_1306);
and U8008 (N_8008,N_1651,N_3988);
nor U8009 (N_8009,N_880,N_74);
or U8010 (N_8010,N_1360,N_2354);
and U8011 (N_8011,N_3659,N_266);
and U8012 (N_8012,N_4243,N_1824);
and U8013 (N_8013,N_4330,N_3636);
nor U8014 (N_8014,N_882,N_898);
and U8015 (N_8015,N_1655,N_737);
xor U8016 (N_8016,N_2885,N_1344);
xor U8017 (N_8017,N_3615,N_3386);
and U8018 (N_8018,N_4793,N_283);
nand U8019 (N_8019,N_3016,N_2148);
or U8020 (N_8020,N_1785,N_3866);
nor U8021 (N_8021,N_1584,N_1687);
nor U8022 (N_8022,N_3313,N_2428);
and U8023 (N_8023,N_1736,N_3902);
nor U8024 (N_8024,N_2720,N_4754);
or U8025 (N_8025,N_2804,N_2233);
or U8026 (N_8026,N_4043,N_1687);
nor U8027 (N_8027,N_2086,N_3642);
nor U8028 (N_8028,N_1733,N_3882);
or U8029 (N_8029,N_4197,N_642);
nor U8030 (N_8030,N_2336,N_256);
xnor U8031 (N_8031,N_4919,N_3494);
and U8032 (N_8032,N_495,N_3381);
xor U8033 (N_8033,N_2638,N_1334);
nor U8034 (N_8034,N_3231,N_2985);
nor U8035 (N_8035,N_535,N_2660);
and U8036 (N_8036,N_4039,N_838);
and U8037 (N_8037,N_3080,N_1893);
and U8038 (N_8038,N_2185,N_4826);
nand U8039 (N_8039,N_2349,N_1826);
nand U8040 (N_8040,N_1085,N_4936);
or U8041 (N_8041,N_4314,N_1298);
nor U8042 (N_8042,N_1062,N_3318);
and U8043 (N_8043,N_2721,N_4723);
or U8044 (N_8044,N_1333,N_1285);
or U8045 (N_8045,N_2562,N_3609);
and U8046 (N_8046,N_3392,N_495);
xor U8047 (N_8047,N_235,N_400);
xnor U8048 (N_8048,N_1362,N_1869);
nand U8049 (N_8049,N_4982,N_4349);
and U8050 (N_8050,N_3091,N_4376);
xnor U8051 (N_8051,N_4784,N_1518);
nor U8052 (N_8052,N_376,N_813);
nor U8053 (N_8053,N_1957,N_3172);
xor U8054 (N_8054,N_1875,N_592);
and U8055 (N_8055,N_2770,N_3257);
nor U8056 (N_8056,N_4567,N_1998);
nand U8057 (N_8057,N_1246,N_311);
nor U8058 (N_8058,N_4447,N_2463);
nor U8059 (N_8059,N_2027,N_3522);
nand U8060 (N_8060,N_3734,N_4726);
xor U8061 (N_8061,N_219,N_1817);
xor U8062 (N_8062,N_3298,N_2527);
xor U8063 (N_8063,N_3517,N_1429);
xor U8064 (N_8064,N_4735,N_3328);
nand U8065 (N_8065,N_1810,N_3321);
nor U8066 (N_8066,N_4477,N_395);
xnor U8067 (N_8067,N_1872,N_4543);
nor U8068 (N_8068,N_1265,N_4695);
or U8069 (N_8069,N_4465,N_2873);
and U8070 (N_8070,N_4982,N_4287);
xnor U8071 (N_8071,N_824,N_656);
nand U8072 (N_8072,N_1154,N_2774);
nor U8073 (N_8073,N_4847,N_184);
and U8074 (N_8074,N_371,N_3669);
xnor U8075 (N_8075,N_4019,N_1384);
nor U8076 (N_8076,N_3524,N_1456);
xor U8077 (N_8077,N_3553,N_3257);
nand U8078 (N_8078,N_1495,N_629);
nor U8079 (N_8079,N_589,N_658);
xor U8080 (N_8080,N_3908,N_87);
nand U8081 (N_8081,N_717,N_4729);
xor U8082 (N_8082,N_4038,N_3190);
nand U8083 (N_8083,N_1457,N_4580);
nor U8084 (N_8084,N_4316,N_1758);
and U8085 (N_8085,N_847,N_1478);
nand U8086 (N_8086,N_4225,N_1940);
nor U8087 (N_8087,N_743,N_3338);
and U8088 (N_8088,N_573,N_3155);
nand U8089 (N_8089,N_1721,N_1384);
and U8090 (N_8090,N_3657,N_831);
and U8091 (N_8091,N_2715,N_4392);
nand U8092 (N_8092,N_3219,N_2836);
nand U8093 (N_8093,N_301,N_4338);
xor U8094 (N_8094,N_617,N_3907);
nor U8095 (N_8095,N_1465,N_1572);
nor U8096 (N_8096,N_2930,N_509);
nor U8097 (N_8097,N_3090,N_3045);
or U8098 (N_8098,N_327,N_3804);
nand U8099 (N_8099,N_4591,N_894);
and U8100 (N_8100,N_3018,N_1550);
or U8101 (N_8101,N_3109,N_3737);
xnor U8102 (N_8102,N_2205,N_4303);
xnor U8103 (N_8103,N_2951,N_4106);
nor U8104 (N_8104,N_3667,N_1008);
xor U8105 (N_8105,N_1912,N_201);
nand U8106 (N_8106,N_4775,N_304);
or U8107 (N_8107,N_2786,N_4421);
nand U8108 (N_8108,N_279,N_2231);
and U8109 (N_8109,N_3304,N_4961);
or U8110 (N_8110,N_2111,N_240);
xnor U8111 (N_8111,N_588,N_787);
nand U8112 (N_8112,N_1091,N_2592);
nand U8113 (N_8113,N_2624,N_12);
nor U8114 (N_8114,N_4792,N_82);
nand U8115 (N_8115,N_3880,N_3661);
and U8116 (N_8116,N_4343,N_2853);
and U8117 (N_8117,N_2980,N_4334);
and U8118 (N_8118,N_2601,N_543);
and U8119 (N_8119,N_830,N_4116);
nor U8120 (N_8120,N_2526,N_4039);
nand U8121 (N_8121,N_4284,N_3231);
or U8122 (N_8122,N_3271,N_3552);
and U8123 (N_8123,N_4226,N_1406);
nand U8124 (N_8124,N_3579,N_4899);
xor U8125 (N_8125,N_1517,N_1350);
nor U8126 (N_8126,N_4657,N_4683);
and U8127 (N_8127,N_732,N_4938);
or U8128 (N_8128,N_3226,N_4765);
and U8129 (N_8129,N_192,N_834);
and U8130 (N_8130,N_3313,N_2655);
nand U8131 (N_8131,N_3771,N_1360);
and U8132 (N_8132,N_1547,N_754);
nor U8133 (N_8133,N_2543,N_1413);
and U8134 (N_8134,N_4543,N_4128);
xor U8135 (N_8135,N_2012,N_1724);
xor U8136 (N_8136,N_2195,N_4419);
and U8137 (N_8137,N_1609,N_82);
nor U8138 (N_8138,N_121,N_3783);
and U8139 (N_8139,N_3240,N_2296);
nor U8140 (N_8140,N_4497,N_2022);
nand U8141 (N_8141,N_1705,N_1489);
xor U8142 (N_8142,N_3726,N_4159);
nand U8143 (N_8143,N_1735,N_2350);
nand U8144 (N_8144,N_3144,N_559);
nor U8145 (N_8145,N_2053,N_1672);
or U8146 (N_8146,N_3084,N_1522);
nor U8147 (N_8147,N_57,N_1286);
and U8148 (N_8148,N_717,N_1318);
and U8149 (N_8149,N_1351,N_103);
or U8150 (N_8150,N_3409,N_2167);
xor U8151 (N_8151,N_3958,N_4847);
xnor U8152 (N_8152,N_4820,N_1584);
nand U8153 (N_8153,N_3251,N_4765);
xor U8154 (N_8154,N_1831,N_454);
and U8155 (N_8155,N_2624,N_523);
and U8156 (N_8156,N_1005,N_891);
nand U8157 (N_8157,N_2680,N_2681);
nand U8158 (N_8158,N_1388,N_2503);
xor U8159 (N_8159,N_4541,N_1006);
or U8160 (N_8160,N_797,N_4781);
nor U8161 (N_8161,N_4490,N_4651);
or U8162 (N_8162,N_2029,N_1621);
or U8163 (N_8163,N_4529,N_3325);
nor U8164 (N_8164,N_3374,N_1039);
xnor U8165 (N_8165,N_4917,N_1359);
or U8166 (N_8166,N_2852,N_879);
nand U8167 (N_8167,N_3221,N_2972);
and U8168 (N_8168,N_839,N_3242);
nor U8169 (N_8169,N_1533,N_678);
xnor U8170 (N_8170,N_1721,N_525);
nor U8171 (N_8171,N_2797,N_1946);
or U8172 (N_8172,N_2106,N_3623);
xnor U8173 (N_8173,N_4674,N_69);
nand U8174 (N_8174,N_3628,N_4873);
xnor U8175 (N_8175,N_2105,N_4585);
nor U8176 (N_8176,N_141,N_3603);
xor U8177 (N_8177,N_1990,N_4323);
nand U8178 (N_8178,N_4947,N_3707);
nand U8179 (N_8179,N_839,N_4990);
nand U8180 (N_8180,N_2908,N_1007);
or U8181 (N_8181,N_728,N_3794);
xnor U8182 (N_8182,N_4753,N_4255);
xnor U8183 (N_8183,N_1482,N_2673);
xor U8184 (N_8184,N_4361,N_1030);
xor U8185 (N_8185,N_3725,N_3715);
nor U8186 (N_8186,N_1716,N_2460);
nor U8187 (N_8187,N_3581,N_1263);
xnor U8188 (N_8188,N_4436,N_2110);
xnor U8189 (N_8189,N_3460,N_4787);
nor U8190 (N_8190,N_4100,N_2726);
or U8191 (N_8191,N_1046,N_731);
xnor U8192 (N_8192,N_4088,N_4014);
nor U8193 (N_8193,N_1846,N_4294);
nor U8194 (N_8194,N_669,N_2233);
or U8195 (N_8195,N_896,N_4828);
nand U8196 (N_8196,N_3733,N_110);
nand U8197 (N_8197,N_590,N_3704);
nor U8198 (N_8198,N_1596,N_4466);
nand U8199 (N_8199,N_1833,N_193);
nor U8200 (N_8200,N_3803,N_2966);
xnor U8201 (N_8201,N_1949,N_1392);
nor U8202 (N_8202,N_1417,N_2240);
nand U8203 (N_8203,N_1145,N_4494);
xnor U8204 (N_8204,N_3637,N_869);
nand U8205 (N_8205,N_3583,N_3659);
or U8206 (N_8206,N_2657,N_1609);
or U8207 (N_8207,N_1404,N_4400);
xnor U8208 (N_8208,N_4065,N_1493);
or U8209 (N_8209,N_3919,N_924);
nor U8210 (N_8210,N_2102,N_502);
and U8211 (N_8211,N_4163,N_3679);
nand U8212 (N_8212,N_1216,N_4824);
nand U8213 (N_8213,N_1058,N_1045);
or U8214 (N_8214,N_1916,N_4218);
nor U8215 (N_8215,N_2381,N_4669);
nor U8216 (N_8216,N_778,N_2304);
and U8217 (N_8217,N_2588,N_2359);
and U8218 (N_8218,N_789,N_4941);
nand U8219 (N_8219,N_3474,N_2306);
xnor U8220 (N_8220,N_4851,N_3327);
or U8221 (N_8221,N_4552,N_1465);
or U8222 (N_8222,N_4786,N_1113);
xor U8223 (N_8223,N_443,N_2198);
and U8224 (N_8224,N_4105,N_4869);
nand U8225 (N_8225,N_4728,N_2468);
nand U8226 (N_8226,N_4171,N_3009);
or U8227 (N_8227,N_2318,N_2189);
or U8228 (N_8228,N_1633,N_51);
or U8229 (N_8229,N_681,N_1606);
or U8230 (N_8230,N_1577,N_3683);
or U8231 (N_8231,N_59,N_2210);
nand U8232 (N_8232,N_2877,N_3825);
or U8233 (N_8233,N_2351,N_3610);
or U8234 (N_8234,N_3248,N_3886);
nor U8235 (N_8235,N_3981,N_2254);
nor U8236 (N_8236,N_1258,N_2375);
and U8237 (N_8237,N_353,N_1198);
nand U8238 (N_8238,N_414,N_4097);
nand U8239 (N_8239,N_1792,N_84);
or U8240 (N_8240,N_558,N_1262);
and U8241 (N_8241,N_3523,N_996);
nand U8242 (N_8242,N_301,N_4929);
nand U8243 (N_8243,N_2242,N_3775);
nor U8244 (N_8244,N_1992,N_3330);
and U8245 (N_8245,N_4697,N_2967);
nand U8246 (N_8246,N_2972,N_39);
and U8247 (N_8247,N_2069,N_4868);
or U8248 (N_8248,N_4849,N_1374);
nand U8249 (N_8249,N_2747,N_2921);
xnor U8250 (N_8250,N_4205,N_2726);
xnor U8251 (N_8251,N_625,N_1154);
xnor U8252 (N_8252,N_1708,N_2786);
nand U8253 (N_8253,N_2221,N_4287);
nor U8254 (N_8254,N_4658,N_4418);
nand U8255 (N_8255,N_595,N_3848);
xnor U8256 (N_8256,N_1413,N_2977);
xor U8257 (N_8257,N_3091,N_2800);
and U8258 (N_8258,N_3733,N_4262);
nand U8259 (N_8259,N_1772,N_169);
xor U8260 (N_8260,N_385,N_1624);
nor U8261 (N_8261,N_3728,N_3518);
nor U8262 (N_8262,N_4065,N_872);
xor U8263 (N_8263,N_3726,N_2999);
nor U8264 (N_8264,N_600,N_973);
and U8265 (N_8265,N_223,N_4085);
and U8266 (N_8266,N_3961,N_1231);
nor U8267 (N_8267,N_3673,N_2702);
and U8268 (N_8268,N_240,N_1934);
xnor U8269 (N_8269,N_390,N_750);
nand U8270 (N_8270,N_420,N_327);
or U8271 (N_8271,N_2923,N_1706);
nor U8272 (N_8272,N_2601,N_4119);
or U8273 (N_8273,N_1878,N_2349);
and U8274 (N_8274,N_4118,N_966);
nand U8275 (N_8275,N_3223,N_883);
nand U8276 (N_8276,N_4315,N_3304);
and U8277 (N_8277,N_570,N_625);
nand U8278 (N_8278,N_225,N_4828);
or U8279 (N_8279,N_3524,N_782);
nand U8280 (N_8280,N_3645,N_2863);
nand U8281 (N_8281,N_2674,N_1854);
and U8282 (N_8282,N_2970,N_2100);
nor U8283 (N_8283,N_1706,N_1557);
xnor U8284 (N_8284,N_2083,N_1447);
nand U8285 (N_8285,N_2143,N_4128);
and U8286 (N_8286,N_4701,N_569);
xnor U8287 (N_8287,N_4229,N_432);
or U8288 (N_8288,N_4051,N_3961);
and U8289 (N_8289,N_4082,N_3591);
xnor U8290 (N_8290,N_4443,N_4321);
or U8291 (N_8291,N_4411,N_3987);
nand U8292 (N_8292,N_61,N_1782);
nand U8293 (N_8293,N_3009,N_4083);
and U8294 (N_8294,N_3824,N_2147);
and U8295 (N_8295,N_28,N_133);
xnor U8296 (N_8296,N_506,N_2674);
xor U8297 (N_8297,N_2617,N_4282);
nor U8298 (N_8298,N_3144,N_1770);
or U8299 (N_8299,N_2156,N_890);
or U8300 (N_8300,N_7,N_4022);
or U8301 (N_8301,N_2793,N_91);
or U8302 (N_8302,N_3041,N_2614);
or U8303 (N_8303,N_2302,N_390);
nand U8304 (N_8304,N_1743,N_2554);
nor U8305 (N_8305,N_819,N_1366);
or U8306 (N_8306,N_4702,N_299);
or U8307 (N_8307,N_4645,N_3734);
nor U8308 (N_8308,N_1846,N_3964);
and U8309 (N_8309,N_1786,N_3543);
and U8310 (N_8310,N_4424,N_1128);
nor U8311 (N_8311,N_223,N_2102);
xnor U8312 (N_8312,N_2559,N_2223);
and U8313 (N_8313,N_4075,N_3315);
xnor U8314 (N_8314,N_4280,N_409);
and U8315 (N_8315,N_1726,N_1108);
nand U8316 (N_8316,N_2724,N_1255);
xnor U8317 (N_8317,N_2869,N_516);
nor U8318 (N_8318,N_1320,N_2309);
xnor U8319 (N_8319,N_4922,N_973);
and U8320 (N_8320,N_894,N_2670);
nand U8321 (N_8321,N_3915,N_3769);
nor U8322 (N_8322,N_2541,N_972);
nand U8323 (N_8323,N_21,N_518);
and U8324 (N_8324,N_2085,N_2298);
or U8325 (N_8325,N_4134,N_3485);
and U8326 (N_8326,N_1219,N_3878);
and U8327 (N_8327,N_1025,N_2280);
or U8328 (N_8328,N_48,N_4782);
and U8329 (N_8329,N_1208,N_1303);
nor U8330 (N_8330,N_4468,N_705);
xnor U8331 (N_8331,N_3731,N_3182);
or U8332 (N_8332,N_2232,N_4609);
or U8333 (N_8333,N_4948,N_854);
and U8334 (N_8334,N_947,N_1097);
or U8335 (N_8335,N_1955,N_4172);
xnor U8336 (N_8336,N_4698,N_4420);
nand U8337 (N_8337,N_189,N_2959);
nor U8338 (N_8338,N_2517,N_4106);
and U8339 (N_8339,N_3420,N_4915);
or U8340 (N_8340,N_2886,N_1724);
nor U8341 (N_8341,N_463,N_1632);
xor U8342 (N_8342,N_4188,N_2293);
nand U8343 (N_8343,N_1986,N_1240);
and U8344 (N_8344,N_2280,N_28);
nor U8345 (N_8345,N_955,N_4384);
nand U8346 (N_8346,N_4057,N_1405);
xor U8347 (N_8347,N_3266,N_2655);
and U8348 (N_8348,N_2245,N_2778);
and U8349 (N_8349,N_4396,N_3231);
and U8350 (N_8350,N_4754,N_652);
nand U8351 (N_8351,N_206,N_2883);
xnor U8352 (N_8352,N_1418,N_718);
and U8353 (N_8353,N_2336,N_2345);
and U8354 (N_8354,N_1483,N_3889);
nor U8355 (N_8355,N_625,N_2904);
or U8356 (N_8356,N_2995,N_4744);
or U8357 (N_8357,N_1229,N_3786);
nor U8358 (N_8358,N_3380,N_3959);
or U8359 (N_8359,N_2280,N_4910);
or U8360 (N_8360,N_4441,N_4567);
or U8361 (N_8361,N_2551,N_4598);
nand U8362 (N_8362,N_3394,N_801);
or U8363 (N_8363,N_3257,N_1631);
xnor U8364 (N_8364,N_1821,N_411);
xnor U8365 (N_8365,N_497,N_2850);
nor U8366 (N_8366,N_548,N_252);
or U8367 (N_8367,N_3114,N_548);
xnor U8368 (N_8368,N_26,N_4478);
or U8369 (N_8369,N_3590,N_2383);
nand U8370 (N_8370,N_4469,N_3393);
nand U8371 (N_8371,N_1178,N_2004);
nor U8372 (N_8372,N_4297,N_442);
and U8373 (N_8373,N_1812,N_51);
nor U8374 (N_8374,N_3099,N_3658);
xnor U8375 (N_8375,N_4750,N_2784);
xnor U8376 (N_8376,N_240,N_2684);
nand U8377 (N_8377,N_187,N_1924);
or U8378 (N_8378,N_4613,N_2263);
xor U8379 (N_8379,N_4416,N_4622);
nor U8380 (N_8380,N_3737,N_968);
xnor U8381 (N_8381,N_2092,N_3385);
nand U8382 (N_8382,N_2264,N_1468);
nor U8383 (N_8383,N_130,N_1101);
nor U8384 (N_8384,N_3949,N_1644);
nor U8385 (N_8385,N_1864,N_2626);
nand U8386 (N_8386,N_1993,N_1647);
xnor U8387 (N_8387,N_3382,N_3350);
nand U8388 (N_8388,N_4214,N_81);
xor U8389 (N_8389,N_631,N_452);
xnor U8390 (N_8390,N_4568,N_3504);
nand U8391 (N_8391,N_4938,N_3902);
nor U8392 (N_8392,N_4511,N_918);
and U8393 (N_8393,N_1002,N_2525);
or U8394 (N_8394,N_4123,N_3877);
nor U8395 (N_8395,N_541,N_3863);
and U8396 (N_8396,N_3153,N_3185);
xnor U8397 (N_8397,N_3551,N_1146);
xor U8398 (N_8398,N_4214,N_4882);
nor U8399 (N_8399,N_3880,N_2700);
and U8400 (N_8400,N_496,N_3378);
or U8401 (N_8401,N_930,N_1570);
xor U8402 (N_8402,N_3404,N_2636);
xnor U8403 (N_8403,N_3576,N_4066);
or U8404 (N_8404,N_2273,N_1067);
nor U8405 (N_8405,N_4159,N_2006);
nor U8406 (N_8406,N_618,N_885);
xnor U8407 (N_8407,N_4003,N_2772);
xor U8408 (N_8408,N_4276,N_1955);
nor U8409 (N_8409,N_3578,N_1600);
and U8410 (N_8410,N_3344,N_2022);
nor U8411 (N_8411,N_87,N_4050);
nand U8412 (N_8412,N_1279,N_202);
xnor U8413 (N_8413,N_4850,N_2547);
xnor U8414 (N_8414,N_2224,N_1970);
xnor U8415 (N_8415,N_2413,N_3596);
nor U8416 (N_8416,N_881,N_4338);
or U8417 (N_8417,N_1810,N_4822);
xnor U8418 (N_8418,N_387,N_1880);
xor U8419 (N_8419,N_4067,N_3243);
or U8420 (N_8420,N_2599,N_4425);
or U8421 (N_8421,N_2907,N_216);
nor U8422 (N_8422,N_4880,N_1254);
and U8423 (N_8423,N_2254,N_2622);
or U8424 (N_8424,N_269,N_1169);
xnor U8425 (N_8425,N_2128,N_2491);
nand U8426 (N_8426,N_3489,N_557);
nor U8427 (N_8427,N_2803,N_468);
nor U8428 (N_8428,N_2969,N_1465);
and U8429 (N_8429,N_3421,N_2637);
nand U8430 (N_8430,N_3612,N_1416);
xor U8431 (N_8431,N_1577,N_2848);
nor U8432 (N_8432,N_35,N_3797);
xnor U8433 (N_8433,N_4632,N_3375);
and U8434 (N_8434,N_679,N_171);
and U8435 (N_8435,N_3850,N_948);
nor U8436 (N_8436,N_1694,N_952);
nor U8437 (N_8437,N_4429,N_1331);
and U8438 (N_8438,N_3844,N_4577);
nor U8439 (N_8439,N_2106,N_973);
and U8440 (N_8440,N_3090,N_3374);
nand U8441 (N_8441,N_2423,N_2265);
xor U8442 (N_8442,N_3679,N_1725);
nand U8443 (N_8443,N_4484,N_1347);
or U8444 (N_8444,N_1343,N_1398);
nor U8445 (N_8445,N_1598,N_2963);
or U8446 (N_8446,N_3226,N_46);
and U8447 (N_8447,N_4778,N_2908);
nor U8448 (N_8448,N_2190,N_2329);
nor U8449 (N_8449,N_3143,N_4219);
nor U8450 (N_8450,N_175,N_3088);
xnor U8451 (N_8451,N_3974,N_2912);
and U8452 (N_8452,N_695,N_1094);
xor U8453 (N_8453,N_3979,N_294);
or U8454 (N_8454,N_3557,N_1934);
or U8455 (N_8455,N_4460,N_4139);
or U8456 (N_8456,N_2230,N_1379);
nor U8457 (N_8457,N_3266,N_3592);
nor U8458 (N_8458,N_377,N_2356);
and U8459 (N_8459,N_4215,N_2916);
or U8460 (N_8460,N_4553,N_1771);
and U8461 (N_8461,N_2180,N_116);
and U8462 (N_8462,N_1894,N_4876);
xor U8463 (N_8463,N_247,N_1678);
nand U8464 (N_8464,N_985,N_2968);
nand U8465 (N_8465,N_4590,N_1507);
and U8466 (N_8466,N_1219,N_2228);
and U8467 (N_8467,N_1125,N_1963);
and U8468 (N_8468,N_1038,N_637);
and U8469 (N_8469,N_2440,N_2865);
and U8470 (N_8470,N_530,N_1683);
or U8471 (N_8471,N_2230,N_859);
and U8472 (N_8472,N_2553,N_3350);
nand U8473 (N_8473,N_3522,N_63);
xnor U8474 (N_8474,N_1470,N_4135);
nand U8475 (N_8475,N_2911,N_629);
nand U8476 (N_8476,N_222,N_4649);
and U8477 (N_8477,N_3301,N_1407);
and U8478 (N_8478,N_2215,N_1911);
xor U8479 (N_8479,N_2777,N_1258);
and U8480 (N_8480,N_3532,N_456);
nor U8481 (N_8481,N_4182,N_3921);
nor U8482 (N_8482,N_3366,N_2426);
and U8483 (N_8483,N_4982,N_3005);
nor U8484 (N_8484,N_4460,N_3748);
nor U8485 (N_8485,N_3490,N_3589);
nor U8486 (N_8486,N_1068,N_3720);
and U8487 (N_8487,N_2691,N_3477);
or U8488 (N_8488,N_4,N_3447);
nand U8489 (N_8489,N_1412,N_3122);
nor U8490 (N_8490,N_3354,N_2427);
xor U8491 (N_8491,N_3832,N_4199);
or U8492 (N_8492,N_4608,N_1516);
nand U8493 (N_8493,N_2451,N_3706);
nand U8494 (N_8494,N_4711,N_4420);
nand U8495 (N_8495,N_2300,N_2910);
xor U8496 (N_8496,N_1250,N_3219);
nor U8497 (N_8497,N_3702,N_452);
nor U8498 (N_8498,N_1095,N_2808);
or U8499 (N_8499,N_1441,N_4873);
or U8500 (N_8500,N_2470,N_711);
nand U8501 (N_8501,N_2384,N_3186);
nor U8502 (N_8502,N_839,N_4923);
nand U8503 (N_8503,N_4108,N_2761);
xnor U8504 (N_8504,N_192,N_3942);
nor U8505 (N_8505,N_3007,N_3930);
and U8506 (N_8506,N_4250,N_1306);
and U8507 (N_8507,N_3388,N_406);
nor U8508 (N_8508,N_4434,N_3082);
nor U8509 (N_8509,N_824,N_1925);
nor U8510 (N_8510,N_1306,N_4973);
or U8511 (N_8511,N_2486,N_4855);
xor U8512 (N_8512,N_3649,N_3137);
nor U8513 (N_8513,N_827,N_530);
and U8514 (N_8514,N_1826,N_4256);
nand U8515 (N_8515,N_2963,N_2390);
or U8516 (N_8516,N_1878,N_2687);
nor U8517 (N_8517,N_2099,N_600);
nor U8518 (N_8518,N_1151,N_1994);
xor U8519 (N_8519,N_3520,N_2260);
nand U8520 (N_8520,N_137,N_4716);
nand U8521 (N_8521,N_1223,N_2752);
xor U8522 (N_8522,N_1103,N_4871);
and U8523 (N_8523,N_2846,N_3740);
nand U8524 (N_8524,N_4295,N_1319);
and U8525 (N_8525,N_4864,N_1342);
xnor U8526 (N_8526,N_1107,N_2105);
xor U8527 (N_8527,N_3576,N_1514);
and U8528 (N_8528,N_1436,N_1034);
nand U8529 (N_8529,N_1490,N_1522);
nor U8530 (N_8530,N_1425,N_867);
nor U8531 (N_8531,N_2415,N_3954);
or U8532 (N_8532,N_3930,N_4023);
nand U8533 (N_8533,N_2638,N_4842);
and U8534 (N_8534,N_1077,N_1359);
xnor U8535 (N_8535,N_4692,N_3690);
and U8536 (N_8536,N_4550,N_3503);
and U8537 (N_8537,N_1467,N_2550);
nor U8538 (N_8538,N_1527,N_1155);
nor U8539 (N_8539,N_1133,N_3838);
nor U8540 (N_8540,N_3523,N_2016);
nor U8541 (N_8541,N_3271,N_2776);
nor U8542 (N_8542,N_619,N_3376);
nand U8543 (N_8543,N_4279,N_3071);
and U8544 (N_8544,N_2570,N_1334);
xnor U8545 (N_8545,N_122,N_2753);
and U8546 (N_8546,N_783,N_1185);
nand U8547 (N_8547,N_4396,N_2285);
and U8548 (N_8548,N_4112,N_2554);
or U8549 (N_8549,N_1511,N_3496);
xnor U8550 (N_8550,N_3450,N_3409);
and U8551 (N_8551,N_432,N_129);
xnor U8552 (N_8552,N_1678,N_3062);
and U8553 (N_8553,N_3019,N_546);
or U8554 (N_8554,N_4715,N_4926);
or U8555 (N_8555,N_4085,N_2714);
nand U8556 (N_8556,N_446,N_1401);
nand U8557 (N_8557,N_1089,N_339);
nand U8558 (N_8558,N_1754,N_3956);
nor U8559 (N_8559,N_4320,N_3722);
nand U8560 (N_8560,N_2028,N_2898);
nand U8561 (N_8561,N_199,N_4067);
xor U8562 (N_8562,N_2238,N_4800);
nor U8563 (N_8563,N_717,N_2147);
and U8564 (N_8564,N_1242,N_507);
nand U8565 (N_8565,N_2703,N_4904);
nor U8566 (N_8566,N_2294,N_3435);
nor U8567 (N_8567,N_3218,N_3174);
xnor U8568 (N_8568,N_3547,N_1012);
nor U8569 (N_8569,N_1096,N_4910);
nor U8570 (N_8570,N_1777,N_2336);
nor U8571 (N_8571,N_1146,N_4840);
nand U8572 (N_8572,N_3120,N_130);
nor U8573 (N_8573,N_15,N_3287);
xnor U8574 (N_8574,N_2139,N_4818);
nor U8575 (N_8575,N_2983,N_3798);
xnor U8576 (N_8576,N_3411,N_3384);
nand U8577 (N_8577,N_4923,N_4128);
and U8578 (N_8578,N_3917,N_2401);
xor U8579 (N_8579,N_1360,N_676);
and U8580 (N_8580,N_4819,N_888);
and U8581 (N_8581,N_1172,N_510);
and U8582 (N_8582,N_3915,N_1940);
or U8583 (N_8583,N_756,N_3354);
xor U8584 (N_8584,N_4268,N_2040);
nor U8585 (N_8585,N_1207,N_2191);
nand U8586 (N_8586,N_642,N_2895);
xnor U8587 (N_8587,N_2403,N_860);
xor U8588 (N_8588,N_1289,N_712);
and U8589 (N_8589,N_994,N_672);
nand U8590 (N_8590,N_3340,N_3520);
nor U8591 (N_8591,N_3001,N_3602);
nand U8592 (N_8592,N_1199,N_4188);
and U8593 (N_8593,N_3565,N_3332);
and U8594 (N_8594,N_2410,N_2484);
nand U8595 (N_8595,N_4663,N_1153);
xor U8596 (N_8596,N_1885,N_1287);
nor U8597 (N_8597,N_1369,N_1678);
nor U8598 (N_8598,N_1344,N_47);
xnor U8599 (N_8599,N_4044,N_3475);
xnor U8600 (N_8600,N_2746,N_3553);
nor U8601 (N_8601,N_3896,N_2438);
or U8602 (N_8602,N_157,N_2296);
and U8603 (N_8603,N_4450,N_202);
nand U8604 (N_8604,N_1802,N_35);
and U8605 (N_8605,N_1136,N_2201);
xor U8606 (N_8606,N_3210,N_3736);
and U8607 (N_8607,N_2506,N_2407);
nand U8608 (N_8608,N_4799,N_1225);
nand U8609 (N_8609,N_3360,N_3425);
nor U8610 (N_8610,N_2216,N_2168);
or U8611 (N_8611,N_2457,N_1967);
nor U8612 (N_8612,N_1613,N_804);
nor U8613 (N_8613,N_2473,N_804);
nor U8614 (N_8614,N_4999,N_4932);
and U8615 (N_8615,N_895,N_1939);
xnor U8616 (N_8616,N_480,N_422);
nor U8617 (N_8617,N_2189,N_2447);
and U8618 (N_8618,N_1323,N_2900);
and U8619 (N_8619,N_4906,N_3836);
or U8620 (N_8620,N_2801,N_3339);
nand U8621 (N_8621,N_4640,N_1126);
nand U8622 (N_8622,N_1356,N_1018);
xor U8623 (N_8623,N_3516,N_46);
and U8624 (N_8624,N_2500,N_3794);
and U8625 (N_8625,N_2370,N_4485);
or U8626 (N_8626,N_3470,N_2948);
nand U8627 (N_8627,N_2482,N_2914);
nand U8628 (N_8628,N_4473,N_3212);
nor U8629 (N_8629,N_2170,N_2952);
nor U8630 (N_8630,N_4959,N_3596);
or U8631 (N_8631,N_678,N_4558);
nor U8632 (N_8632,N_460,N_41);
nor U8633 (N_8633,N_738,N_3002);
or U8634 (N_8634,N_2516,N_4161);
nand U8635 (N_8635,N_2094,N_1851);
or U8636 (N_8636,N_4652,N_1475);
and U8637 (N_8637,N_2649,N_3805);
nor U8638 (N_8638,N_2104,N_4006);
nor U8639 (N_8639,N_4667,N_4077);
nand U8640 (N_8640,N_799,N_4532);
and U8641 (N_8641,N_474,N_868);
nor U8642 (N_8642,N_2039,N_3820);
or U8643 (N_8643,N_2740,N_4811);
nor U8644 (N_8644,N_926,N_4101);
nor U8645 (N_8645,N_1899,N_2575);
or U8646 (N_8646,N_3274,N_3398);
nand U8647 (N_8647,N_263,N_3890);
xor U8648 (N_8648,N_1019,N_2673);
or U8649 (N_8649,N_1908,N_335);
xor U8650 (N_8650,N_4674,N_3169);
and U8651 (N_8651,N_878,N_716);
and U8652 (N_8652,N_2568,N_2577);
and U8653 (N_8653,N_2506,N_2149);
nor U8654 (N_8654,N_155,N_2665);
nor U8655 (N_8655,N_1545,N_247);
nand U8656 (N_8656,N_736,N_4230);
nand U8657 (N_8657,N_362,N_2705);
and U8658 (N_8658,N_1088,N_603);
xnor U8659 (N_8659,N_3038,N_2584);
and U8660 (N_8660,N_760,N_2380);
nand U8661 (N_8661,N_2896,N_3559);
nor U8662 (N_8662,N_3359,N_148);
or U8663 (N_8663,N_1966,N_2382);
or U8664 (N_8664,N_2051,N_3829);
and U8665 (N_8665,N_3328,N_2107);
nor U8666 (N_8666,N_1235,N_372);
nor U8667 (N_8667,N_2069,N_2844);
nor U8668 (N_8668,N_1265,N_479);
xor U8669 (N_8669,N_2251,N_1713);
xor U8670 (N_8670,N_1492,N_2434);
and U8671 (N_8671,N_2146,N_3216);
xor U8672 (N_8672,N_1388,N_611);
or U8673 (N_8673,N_4968,N_306);
and U8674 (N_8674,N_4973,N_2521);
nor U8675 (N_8675,N_699,N_3755);
xnor U8676 (N_8676,N_4642,N_1279);
and U8677 (N_8677,N_1427,N_4971);
nand U8678 (N_8678,N_3990,N_3774);
nand U8679 (N_8679,N_320,N_114);
or U8680 (N_8680,N_2278,N_532);
nor U8681 (N_8681,N_1906,N_469);
and U8682 (N_8682,N_597,N_4533);
and U8683 (N_8683,N_44,N_4016);
or U8684 (N_8684,N_4014,N_1498);
and U8685 (N_8685,N_3898,N_2771);
nand U8686 (N_8686,N_759,N_4808);
nand U8687 (N_8687,N_3594,N_680);
xnor U8688 (N_8688,N_2648,N_3201);
xnor U8689 (N_8689,N_4525,N_4712);
or U8690 (N_8690,N_1968,N_3006);
xnor U8691 (N_8691,N_4402,N_2951);
or U8692 (N_8692,N_1411,N_1306);
nand U8693 (N_8693,N_4654,N_2922);
nand U8694 (N_8694,N_4919,N_178);
and U8695 (N_8695,N_4433,N_3226);
nand U8696 (N_8696,N_3640,N_1583);
or U8697 (N_8697,N_2240,N_1063);
nand U8698 (N_8698,N_169,N_1343);
nand U8699 (N_8699,N_2498,N_4160);
nor U8700 (N_8700,N_265,N_4282);
or U8701 (N_8701,N_1017,N_4794);
and U8702 (N_8702,N_2717,N_2761);
xnor U8703 (N_8703,N_1576,N_4214);
or U8704 (N_8704,N_1892,N_4860);
nand U8705 (N_8705,N_2730,N_4765);
nand U8706 (N_8706,N_1777,N_3060);
nor U8707 (N_8707,N_4703,N_2376);
or U8708 (N_8708,N_4861,N_446);
and U8709 (N_8709,N_4193,N_2430);
nor U8710 (N_8710,N_3560,N_453);
nand U8711 (N_8711,N_3994,N_416);
nor U8712 (N_8712,N_3514,N_2638);
and U8713 (N_8713,N_3028,N_854);
nor U8714 (N_8714,N_1324,N_1365);
nand U8715 (N_8715,N_4782,N_3798);
xnor U8716 (N_8716,N_2743,N_1944);
nand U8717 (N_8717,N_590,N_227);
and U8718 (N_8718,N_3659,N_1788);
and U8719 (N_8719,N_3807,N_2724);
or U8720 (N_8720,N_1786,N_260);
nand U8721 (N_8721,N_1509,N_1567);
xnor U8722 (N_8722,N_966,N_2546);
nor U8723 (N_8723,N_3514,N_3126);
or U8724 (N_8724,N_3802,N_2738);
or U8725 (N_8725,N_3639,N_2503);
and U8726 (N_8726,N_4681,N_1280);
and U8727 (N_8727,N_4757,N_3581);
xor U8728 (N_8728,N_3289,N_4977);
and U8729 (N_8729,N_1175,N_1098);
nand U8730 (N_8730,N_19,N_1159);
or U8731 (N_8731,N_459,N_4400);
nor U8732 (N_8732,N_1119,N_1830);
nor U8733 (N_8733,N_1082,N_2289);
and U8734 (N_8734,N_2787,N_3835);
nand U8735 (N_8735,N_2624,N_3384);
xor U8736 (N_8736,N_1414,N_1157);
nor U8737 (N_8737,N_21,N_3670);
or U8738 (N_8738,N_576,N_2388);
and U8739 (N_8739,N_3421,N_3732);
and U8740 (N_8740,N_1026,N_714);
nand U8741 (N_8741,N_2594,N_3127);
nor U8742 (N_8742,N_2962,N_1825);
or U8743 (N_8743,N_745,N_4627);
or U8744 (N_8744,N_1184,N_3499);
nand U8745 (N_8745,N_2009,N_4643);
nor U8746 (N_8746,N_4621,N_3406);
or U8747 (N_8747,N_279,N_2442);
and U8748 (N_8748,N_4175,N_701);
xor U8749 (N_8749,N_2966,N_3419);
nor U8750 (N_8750,N_3334,N_3456);
and U8751 (N_8751,N_224,N_1724);
xnor U8752 (N_8752,N_1973,N_3647);
or U8753 (N_8753,N_2683,N_1426);
or U8754 (N_8754,N_3500,N_2181);
and U8755 (N_8755,N_3891,N_3058);
and U8756 (N_8756,N_4011,N_310);
xor U8757 (N_8757,N_3155,N_1948);
nor U8758 (N_8758,N_490,N_471);
nand U8759 (N_8759,N_4239,N_4361);
xnor U8760 (N_8760,N_693,N_4235);
and U8761 (N_8761,N_3518,N_3231);
and U8762 (N_8762,N_1882,N_3640);
nand U8763 (N_8763,N_4647,N_552);
and U8764 (N_8764,N_653,N_2115);
nand U8765 (N_8765,N_4059,N_1420);
and U8766 (N_8766,N_1250,N_416);
xor U8767 (N_8767,N_1827,N_505);
and U8768 (N_8768,N_3496,N_2643);
nand U8769 (N_8769,N_959,N_4219);
xor U8770 (N_8770,N_324,N_2395);
xor U8771 (N_8771,N_4410,N_1253);
nor U8772 (N_8772,N_852,N_4191);
nand U8773 (N_8773,N_3234,N_1177);
and U8774 (N_8774,N_4069,N_996);
nor U8775 (N_8775,N_1676,N_2055);
nor U8776 (N_8776,N_1196,N_4749);
or U8777 (N_8777,N_3634,N_4727);
or U8778 (N_8778,N_2707,N_1301);
or U8779 (N_8779,N_4744,N_1821);
nand U8780 (N_8780,N_4153,N_2953);
xnor U8781 (N_8781,N_3111,N_2123);
xor U8782 (N_8782,N_3234,N_4696);
nand U8783 (N_8783,N_3503,N_620);
nor U8784 (N_8784,N_4645,N_4190);
and U8785 (N_8785,N_3565,N_4273);
and U8786 (N_8786,N_3828,N_4655);
nand U8787 (N_8787,N_3332,N_2115);
nand U8788 (N_8788,N_3319,N_4951);
and U8789 (N_8789,N_3702,N_1342);
xor U8790 (N_8790,N_4076,N_2038);
or U8791 (N_8791,N_714,N_1898);
nand U8792 (N_8792,N_3634,N_634);
and U8793 (N_8793,N_4318,N_1281);
nand U8794 (N_8794,N_1706,N_2401);
xnor U8795 (N_8795,N_555,N_4435);
or U8796 (N_8796,N_2943,N_2020);
or U8797 (N_8797,N_4684,N_2607);
xor U8798 (N_8798,N_4095,N_549);
or U8799 (N_8799,N_1961,N_3620);
and U8800 (N_8800,N_3616,N_1465);
or U8801 (N_8801,N_2137,N_4473);
or U8802 (N_8802,N_958,N_4709);
nor U8803 (N_8803,N_4827,N_1659);
nor U8804 (N_8804,N_987,N_4493);
nor U8805 (N_8805,N_3528,N_4698);
or U8806 (N_8806,N_2563,N_2939);
xor U8807 (N_8807,N_3997,N_3791);
xnor U8808 (N_8808,N_206,N_4841);
nor U8809 (N_8809,N_3029,N_4207);
nor U8810 (N_8810,N_1918,N_4253);
xnor U8811 (N_8811,N_2403,N_3200);
nand U8812 (N_8812,N_2763,N_2385);
xnor U8813 (N_8813,N_406,N_552);
or U8814 (N_8814,N_3741,N_2102);
or U8815 (N_8815,N_1908,N_4228);
nand U8816 (N_8816,N_3669,N_4343);
or U8817 (N_8817,N_3218,N_512);
xnor U8818 (N_8818,N_76,N_370);
and U8819 (N_8819,N_1836,N_653);
or U8820 (N_8820,N_3482,N_4507);
and U8821 (N_8821,N_3468,N_2703);
or U8822 (N_8822,N_4415,N_3000);
nor U8823 (N_8823,N_4673,N_4770);
nand U8824 (N_8824,N_1386,N_3700);
or U8825 (N_8825,N_3569,N_3242);
and U8826 (N_8826,N_734,N_112);
nand U8827 (N_8827,N_1227,N_1498);
xnor U8828 (N_8828,N_3980,N_4676);
nor U8829 (N_8829,N_3239,N_2776);
and U8830 (N_8830,N_3555,N_1541);
and U8831 (N_8831,N_4982,N_4456);
nor U8832 (N_8832,N_4430,N_4975);
and U8833 (N_8833,N_1705,N_671);
and U8834 (N_8834,N_2668,N_3573);
xor U8835 (N_8835,N_4269,N_3724);
nor U8836 (N_8836,N_4433,N_4642);
and U8837 (N_8837,N_2794,N_561);
xnor U8838 (N_8838,N_3781,N_1539);
or U8839 (N_8839,N_4972,N_247);
xor U8840 (N_8840,N_3347,N_3214);
nor U8841 (N_8841,N_2410,N_648);
nand U8842 (N_8842,N_4932,N_1235);
nand U8843 (N_8843,N_1869,N_3863);
and U8844 (N_8844,N_4720,N_1859);
nand U8845 (N_8845,N_4284,N_439);
nor U8846 (N_8846,N_154,N_1148);
xor U8847 (N_8847,N_2668,N_2272);
and U8848 (N_8848,N_4897,N_3637);
nor U8849 (N_8849,N_1751,N_3596);
nor U8850 (N_8850,N_2462,N_3238);
xnor U8851 (N_8851,N_1490,N_1998);
nor U8852 (N_8852,N_2418,N_4558);
or U8853 (N_8853,N_2115,N_3677);
nand U8854 (N_8854,N_858,N_1836);
or U8855 (N_8855,N_4551,N_1049);
xor U8856 (N_8856,N_4141,N_4458);
nand U8857 (N_8857,N_3846,N_732);
xor U8858 (N_8858,N_3883,N_1496);
nand U8859 (N_8859,N_2457,N_4978);
or U8860 (N_8860,N_3348,N_3691);
nand U8861 (N_8861,N_1577,N_1396);
nand U8862 (N_8862,N_2946,N_780);
and U8863 (N_8863,N_2569,N_3988);
xnor U8864 (N_8864,N_3473,N_4150);
and U8865 (N_8865,N_2090,N_1082);
nand U8866 (N_8866,N_4361,N_2192);
nor U8867 (N_8867,N_591,N_2497);
nor U8868 (N_8868,N_805,N_2656);
nor U8869 (N_8869,N_2741,N_828);
xor U8870 (N_8870,N_1191,N_1368);
nand U8871 (N_8871,N_1584,N_1421);
or U8872 (N_8872,N_679,N_151);
nor U8873 (N_8873,N_1150,N_2812);
and U8874 (N_8874,N_767,N_147);
or U8875 (N_8875,N_2425,N_1635);
xor U8876 (N_8876,N_388,N_1173);
and U8877 (N_8877,N_2524,N_2564);
or U8878 (N_8878,N_3010,N_3454);
and U8879 (N_8879,N_2073,N_1371);
or U8880 (N_8880,N_1687,N_820);
or U8881 (N_8881,N_3320,N_296);
or U8882 (N_8882,N_1941,N_3088);
nor U8883 (N_8883,N_504,N_1984);
nor U8884 (N_8884,N_1863,N_4814);
nand U8885 (N_8885,N_4875,N_2362);
or U8886 (N_8886,N_1837,N_2892);
and U8887 (N_8887,N_3596,N_1931);
nand U8888 (N_8888,N_3283,N_924);
and U8889 (N_8889,N_3095,N_407);
nor U8890 (N_8890,N_4444,N_3240);
or U8891 (N_8891,N_3553,N_2607);
xor U8892 (N_8892,N_330,N_3549);
and U8893 (N_8893,N_742,N_2704);
and U8894 (N_8894,N_1449,N_2700);
or U8895 (N_8895,N_2025,N_1103);
xor U8896 (N_8896,N_2622,N_2602);
and U8897 (N_8897,N_4133,N_1228);
nor U8898 (N_8898,N_36,N_3456);
and U8899 (N_8899,N_4087,N_386);
and U8900 (N_8900,N_1296,N_1899);
nand U8901 (N_8901,N_1597,N_985);
nor U8902 (N_8902,N_3312,N_296);
xnor U8903 (N_8903,N_3427,N_4855);
nand U8904 (N_8904,N_1282,N_4189);
or U8905 (N_8905,N_2859,N_775);
or U8906 (N_8906,N_3258,N_4600);
nor U8907 (N_8907,N_1609,N_4981);
xnor U8908 (N_8908,N_677,N_2298);
nor U8909 (N_8909,N_2523,N_2070);
and U8910 (N_8910,N_3093,N_2665);
and U8911 (N_8911,N_1044,N_113);
xor U8912 (N_8912,N_4709,N_3855);
xnor U8913 (N_8913,N_3584,N_209);
and U8914 (N_8914,N_4984,N_4235);
nand U8915 (N_8915,N_3845,N_2805);
nor U8916 (N_8916,N_2661,N_465);
xor U8917 (N_8917,N_585,N_309);
or U8918 (N_8918,N_4633,N_1241);
xnor U8919 (N_8919,N_3325,N_4353);
xor U8920 (N_8920,N_2793,N_1682);
and U8921 (N_8921,N_2474,N_336);
and U8922 (N_8922,N_2075,N_4173);
and U8923 (N_8923,N_4393,N_632);
and U8924 (N_8924,N_26,N_1026);
or U8925 (N_8925,N_635,N_914);
and U8926 (N_8926,N_3872,N_2402);
and U8927 (N_8927,N_1680,N_68);
xnor U8928 (N_8928,N_3852,N_863);
nand U8929 (N_8929,N_2093,N_1484);
or U8930 (N_8930,N_4328,N_1388);
nor U8931 (N_8931,N_2673,N_2787);
or U8932 (N_8932,N_1694,N_3533);
nand U8933 (N_8933,N_4684,N_2874);
or U8934 (N_8934,N_2878,N_3789);
or U8935 (N_8935,N_3000,N_1106);
or U8936 (N_8936,N_1258,N_3093);
and U8937 (N_8937,N_2721,N_2853);
nor U8938 (N_8938,N_4941,N_1774);
nor U8939 (N_8939,N_4822,N_4025);
and U8940 (N_8940,N_1917,N_4368);
nor U8941 (N_8941,N_3033,N_2700);
xnor U8942 (N_8942,N_221,N_4815);
nor U8943 (N_8943,N_4346,N_2791);
nand U8944 (N_8944,N_3969,N_4172);
nor U8945 (N_8945,N_2629,N_674);
or U8946 (N_8946,N_2535,N_294);
xnor U8947 (N_8947,N_1271,N_4571);
xor U8948 (N_8948,N_3471,N_3381);
xor U8949 (N_8949,N_2014,N_723);
and U8950 (N_8950,N_2202,N_795);
nand U8951 (N_8951,N_2539,N_4111);
nor U8952 (N_8952,N_2168,N_1517);
nor U8953 (N_8953,N_2909,N_4450);
or U8954 (N_8954,N_4138,N_261);
and U8955 (N_8955,N_3656,N_772);
or U8956 (N_8956,N_1080,N_856);
nand U8957 (N_8957,N_4891,N_56);
xnor U8958 (N_8958,N_3820,N_1165);
nand U8959 (N_8959,N_2346,N_1);
nor U8960 (N_8960,N_3212,N_4457);
xor U8961 (N_8961,N_4044,N_3690);
or U8962 (N_8962,N_1021,N_936);
and U8963 (N_8963,N_4505,N_2109);
xnor U8964 (N_8964,N_3758,N_3307);
xnor U8965 (N_8965,N_2001,N_2154);
nand U8966 (N_8966,N_4410,N_2419);
xnor U8967 (N_8967,N_4806,N_3888);
nor U8968 (N_8968,N_2361,N_2081);
and U8969 (N_8969,N_3705,N_3908);
or U8970 (N_8970,N_924,N_4933);
nand U8971 (N_8971,N_3910,N_423);
nand U8972 (N_8972,N_1929,N_1856);
nand U8973 (N_8973,N_1396,N_2572);
xor U8974 (N_8974,N_482,N_4948);
or U8975 (N_8975,N_3205,N_1494);
and U8976 (N_8976,N_4346,N_1847);
and U8977 (N_8977,N_3230,N_3695);
xnor U8978 (N_8978,N_951,N_3350);
and U8979 (N_8979,N_3396,N_1159);
nor U8980 (N_8980,N_935,N_2844);
xnor U8981 (N_8981,N_516,N_3184);
nor U8982 (N_8982,N_878,N_3866);
nand U8983 (N_8983,N_2991,N_72);
xor U8984 (N_8984,N_428,N_3929);
or U8985 (N_8985,N_1164,N_2148);
nor U8986 (N_8986,N_2682,N_45);
or U8987 (N_8987,N_4170,N_2111);
and U8988 (N_8988,N_3902,N_3679);
nor U8989 (N_8989,N_332,N_2799);
xnor U8990 (N_8990,N_962,N_2379);
and U8991 (N_8991,N_2021,N_1964);
xor U8992 (N_8992,N_2274,N_1043);
nand U8993 (N_8993,N_4112,N_1705);
xnor U8994 (N_8994,N_3862,N_2493);
and U8995 (N_8995,N_3616,N_2997);
nor U8996 (N_8996,N_1571,N_4793);
or U8997 (N_8997,N_1639,N_1262);
or U8998 (N_8998,N_195,N_3806);
or U8999 (N_8999,N_3274,N_587);
or U9000 (N_9000,N_658,N_4844);
or U9001 (N_9001,N_3142,N_3613);
and U9002 (N_9002,N_264,N_1229);
nor U9003 (N_9003,N_374,N_3215);
nor U9004 (N_9004,N_626,N_4715);
nor U9005 (N_9005,N_4920,N_13);
xnor U9006 (N_9006,N_3439,N_2766);
or U9007 (N_9007,N_4033,N_3466);
xnor U9008 (N_9008,N_3002,N_2987);
or U9009 (N_9009,N_4611,N_569);
nor U9010 (N_9010,N_845,N_4456);
and U9011 (N_9011,N_1486,N_3948);
xor U9012 (N_9012,N_874,N_1489);
nor U9013 (N_9013,N_4778,N_1282);
nor U9014 (N_9014,N_3377,N_4097);
and U9015 (N_9015,N_3873,N_1663);
and U9016 (N_9016,N_4673,N_3191);
or U9017 (N_9017,N_20,N_2392);
nor U9018 (N_9018,N_2317,N_3334);
nand U9019 (N_9019,N_4026,N_4131);
nor U9020 (N_9020,N_4926,N_2587);
xnor U9021 (N_9021,N_3425,N_4779);
nor U9022 (N_9022,N_1153,N_4741);
or U9023 (N_9023,N_527,N_1108);
nor U9024 (N_9024,N_1944,N_1372);
and U9025 (N_9025,N_3378,N_3098);
xnor U9026 (N_9026,N_2773,N_4760);
or U9027 (N_9027,N_4396,N_3431);
or U9028 (N_9028,N_1183,N_3339);
nand U9029 (N_9029,N_305,N_1808);
and U9030 (N_9030,N_1617,N_807);
nand U9031 (N_9031,N_3855,N_3377);
xnor U9032 (N_9032,N_505,N_1205);
nor U9033 (N_9033,N_2160,N_892);
xnor U9034 (N_9034,N_3302,N_1540);
nor U9035 (N_9035,N_4632,N_2270);
nand U9036 (N_9036,N_2216,N_2267);
nand U9037 (N_9037,N_25,N_3414);
nor U9038 (N_9038,N_1518,N_1093);
nand U9039 (N_9039,N_1988,N_1099);
nand U9040 (N_9040,N_70,N_598);
or U9041 (N_9041,N_1482,N_4779);
xnor U9042 (N_9042,N_1201,N_3698);
and U9043 (N_9043,N_3280,N_597);
nand U9044 (N_9044,N_3556,N_3097);
nor U9045 (N_9045,N_3006,N_2790);
xnor U9046 (N_9046,N_3967,N_3345);
nor U9047 (N_9047,N_1264,N_4888);
and U9048 (N_9048,N_1013,N_678);
nand U9049 (N_9049,N_4011,N_2461);
xnor U9050 (N_9050,N_2088,N_239);
nand U9051 (N_9051,N_3953,N_4190);
and U9052 (N_9052,N_4494,N_3998);
or U9053 (N_9053,N_3237,N_4597);
and U9054 (N_9054,N_2508,N_4191);
and U9055 (N_9055,N_1910,N_383);
or U9056 (N_9056,N_2151,N_979);
xor U9057 (N_9057,N_2612,N_2576);
xnor U9058 (N_9058,N_4426,N_4842);
nand U9059 (N_9059,N_2316,N_1641);
or U9060 (N_9060,N_3999,N_3368);
and U9061 (N_9061,N_4275,N_4462);
xor U9062 (N_9062,N_4428,N_2100);
xor U9063 (N_9063,N_1368,N_3310);
xor U9064 (N_9064,N_2878,N_3792);
and U9065 (N_9065,N_2875,N_3970);
or U9066 (N_9066,N_202,N_3931);
and U9067 (N_9067,N_317,N_1123);
xnor U9068 (N_9068,N_857,N_2103);
and U9069 (N_9069,N_3633,N_2779);
xnor U9070 (N_9070,N_313,N_1682);
xor U9071 (N_9071,N_2506,N_2677);
nand U9072 (N_9072,N_3952,N_1902);
and U9073 (N_9073,N_2600,N_2040);
and U9074 (N_9074,N_1198,N_2802);
xor U9075 (N_9075,N_3095,N_1116);
nand U9076 (N_9076,N_4323,N_1471);
nor U9077 (N_9077,N_2342,N_4984);
xor U9078 (N_9078,N_793,N_1774);
or U9079 (N_9079,N_1646,N_3774);
nand U9080 (N_9080,N_1993,N_4362);
nor U9081 (N_9081,N_969,N_2157);
xor U9082 (N_9082,N_3236,N_3878);
and U9083 (N_9083,N_3335,N_4802);
or U9084 (N_9084,N_3648,N_529);
nand U9085 (N_9085,N_2838,N_1766);
or U9086 (N_9086,N_2857,N_4722);
xnor U9087 (N_9087,N_2441,N_1378);
xor U9088 (N_9088,N_1635,N_4254);
and U9089 (N_9089,N_2776,N_3664);
or U9090 (N_9090,N_3359,N_922);
xnor U9091 (N_9091,N_2406,N_2960);
or U9092 (N_9092,N_744,N_427);
or U9093 (N_9093,N_4842,N_485);
xnor U9094 (N_9094,N_1304,N_1514);
or U9095 (N_9095,N_1431,N_736);
and U9096 (N_9096,N_4647,N_845);
xor U9097 (N_9097,N_514,N_4613);
nor U9098 (N_9098,N_1401,N_11);
nor U9099 (N_9099,N_2983,N_2979);
or U9100 (N_9100,N_2292,N_3535);
xnor U9101 (N_9101,N_4334,N_1620);
or U9102 (N_9102,N_2896,N_439);
or U9103 (N_9103,N_3335,N_3826);
nor U9104 (N_9104,N_1711,N_313);
nand U9105 (N_9105,N_3328,N_331);
nor U9106 (N_9106,N_633,N_1618);
nand U9107 (N_9107,N_4075,N_1375);
nand U9108 (N_9108,N_1551,N_1550);
nor U9109 (N_9109,N_1309,N_325);
nand U9110 (N_9110,N_1915,N_1718);
or U9111 (N_9111,N_4545,N_3607);
nand U9112 (N_9112,N_3509,N_2847);
nor U9113 (N_9113,N_2875,N_4216);
and U9114 (N_9114,N_1976,N_4908);
and U9115 (N_9115,N_3937,N_4170);
or U9116 (N_9116,N_2284,N_27);
and U9117 (N_9117,N_3700,N_3733);
xnor U9118 (N_9118,N_1331,N_2702);
nor U9119 (N_9119,N_669,N_1729);
nand U9120 (N_9120,N_4132,N_730);
nor U9121 (N_9121,N_1832,N_1124);
or U9122 (N_9122,N_3420,N_909);
xor U9123 (N_9123,N_1219,N_365);
or U9124 (N_9124,N_1306,N_2394);
xnor U9125 (N_9125,N_1301,N_1712);
nor U9126 (N_9126,N_2256,N_3212);
or U9127 (N_9127,N_1554,N_1289);
and U9128 (N_9128,N_3224,N_620);
and U9129 (N_9129,N_4659,N_2213);
or U9130 (N_9130,N_641,N_4238);
nor U9131 (N_9131,N_1658,N_3773);
or U9132 (N_9132,N_4104,N_1325);
and U9133 (N_9133,N_3004,N_283);
or U9134 (N_9134,N_406,N_4634);
xor U9135 (N_9135,N_1517,N_3290);
nand U9136 (N_9136,N_414,N_3127);
nand U9137 (N_9137,N_4849,N_581);
nand U9138 (N_9138,N_1828,N_68);
or U9139 (N_9139,N_2674,N_2284);
or U9140 (N_9140,N_3717,N_1648);
nand U9141 (N_9141,N_1829,N_3034);
nor U9142 (N_9142,N_800,N_1845);
nand U9143 (N_9143,N_2690,N_3811);
xnor U9144 (N_9144,N_1187,N_4886);
xor U9145 (N_9145,N_3620,N_2599);
nor U9146 (N_9146,N_773,N_3411);
and U9147 (N_9147,N_459,N_1461);
nor U9148 (N_9148,N_1952,N_3099);
xor U9149 (N_9149,N_1955,N_4207);
nand U9150 (N_9150,N_1346,N_4968);
nor U9151 (N_9151,N_4049,N_1653);
nor U9152 (N_9152,N_4068,N_2527);
nor U9153 (N_9153,N_759,N_2102);
xor U9154 (N_9154,N_3834,N_2709);
or U9155 (N_9155,N_4814,N_4274);
nor U9156 (N_9156,N_2952,N_2476);
and U9157 (N_9157,N_2919,N_3360);
nor U9158 (N_9158,N_2153,N_3606);
nand U9159 (N_9159,N_1133,N_350);
nor U9160 (N_9160,N_597,N_1191);
nand U9161 (N_9161,N_546,N_4163);
nand U9162 (N_9162,N_1425,N_3557);
or U9163 (N_9163,N_3819,N_4669);
or U9164 (N_9164,N_661,N_1633);
nor U9165 (N_9165,N_957,N_4985);
nand U9166 (N_9166,N_3348,N_3593);
nand U9167 (N_9167,N_4815,N_2071);
xor U9168 (N_9168,N_1427,N_4496);
nand U9169 (N_9169,N_4206,N_3659);
or U9170 (N_9170,N_3696,N_2073);
or U9171 (N_9171,N_4971,N_2396);
and U9172 (N_9172,N_1510,N_852);
and U9173 (N_9173,N_2642,N_293);
nor U9174 (N_9174,N_4577,N_1294);
and U9175 (N_9175,N_1526,N_875);
nor U9176 (N_9176,N_1074,N_2276);
xor U9177 (N_9177,N_3003,N_4550);
or U9178 (N_9178,N_315,N_2421);
xnor U9179 (N_9179,N_639,N_4550);
xor U9180 (N_9180,N_2130,N_54);
nand U9181 (N_9181,N_384,N_1286);
and U9182 (N_9182,N_3363,N_2475);
nor U9183 (N_9183,N_532,N_707);
or U9184 (N_9184,N_457,N_332);
or U9185 (N_9185,N_3336,N_1784);
and U9186 (N_9186,N_2186,N_4380);
and U9187 (N_9187,N_4878,N_3260);
nand U9188 (N_9188,N_3970,N_3098);
or U9189 (N_9189,N_2014,N_3037);
and U9190 (N_9190,N_4245,N_547);
xnor U9191 (N_9191,N_1547,N_2518);
xor U9192 (N_9192,N_2818,N_2991);
or U9193 (N_9193,N_3577,N_1543);
xnor U9194 (N_9194,N_2182,N_2435);
xor U9195 (N_9195,N_4702,N_4958);
and U9196 (N_9196,N_197,N_1491);
nand U9197 (N_9197,N_196,N_1265);
xnor U9198 (N_9198,N_601,N_1620);
nand U9199 (N_9199,N_606,N_3780);
and U9200 (N_9200,N_4424,N_2030);
nand U9201 (N_9201,N_2686,N_1611);
nand U9202 (N_9202,N_1646,N_4919);
xor U9203 (N_9203,N_1499,N_279);
nand U9204 (N_9204,N_2215,N_3346);
or U9205 (N_9205,N_2186,N_3878);
or U9206 (N_9206,N_2538,N_4483);
nor U9207 (N_9207,N_1436,N_79);
nand U9208 (N_9208,N_2209,N_2137);
xor U9209 (N_9209,N_1464,N_1514);
nor U9210 (N_9210,N_4110,N_3422);
nand U9211 (N_9211,N_3615,N_4161);
xnor U9212 (N_9212,N_3467,N_4325);
nand U9213 (N_9213,N_1954,N_3264);
or U9214 (N_9214,N_4353,N_3551);
nand U9215 (N_9215,N_428,N_3570);
or U9216 (N_9216,N_15,N_3586);
xor U9217 (N_9217,N_3868,N_597);
nand U9218 (N_9218,N_1447,N_2304);
nand U9219 (N_9219,N_3394,N_4666);
nand U9220 (N_9220,N_4355,N_3310);
nand U9221 (N_9221,N_3032,N_4873);
or U9222 (N_9222,N_3650,N_859);
and U9223 (N_9223,N_4344,N_2411);
xor U9224 (N_9224,N_4962,N_3439);
and U9225 (N_9225,N_566,N_4484);
nor U9226 (N_9226,N_3955,N_3069);
xnor U9227 (N_9227,N_3912,N_778);
or U9228 (N_9228,N_4036,N_3067);
and U9229 (N_9229,N_1032,N_1325);
or U9230 (N_9230,N_1800,N_3292);
xor U9231 (N_9231,N_1194,N_2071);
nor U9232 (N_9232,N_1349,N_2407);
nor U9233 (N_9233,N_4161,N_2657);
nand U9234 (N_9234,N_4593,N_4311);
and U9235 (N_9235,N_3762,N_4282);
and U9236 (N_9236,N_456,N_885);
and U9237 (N_9237,N_373,N_3440);
nand U9238 (N_9238,N_3274,N_4554);
nor U9239 (N_9239,N_419,N_3456);
or U9240 (N_9240,N_2703,N_4989);
or U9241 (N_9241,N_3238,N_4095);
or U9242 (N_9242,N_4208,N_4339);
and U9243 (N_9243,N_654,N_4985);
and U9244 (N_9244,N_916,N_619);
or U9245 (N_9245,N_4452,N_497);
and U9246 (N_9246,N_2242,N_4802);
nand U9247 (N_9247,N_62,N_1415);
and U9248 (N_9248,N_1170,N_1964);
and U9249 (N_9249,N_4892,N_1033);
nor U9250 (N_9250,N_3726,N_3848);
xnor U9251 (N_9251,N_331,N_105);
nand U9252 (N_9252,N_3811,N_218);
or U9253 (N_9253,N_3109,N_1887);
nand U9254 (N_9254,N_1496,N_2888);
nand U9255 (N_9255,N_3233,N_175);
nor U9256 (N_9256,N_795,N_584);
xor U9257 (N_9257,N_3165,N_4966);
nor U9258 (N_9258,N_4298,N_2896);
and U9259 (N_9259,N_504,N_3553);
nand U9260 (N_9260,N_4835,N_671);
nand U9261 (N_9261,N_2693,N_3528);
and U9262 (N_9262,N_2839,N_2520);
or U9263 (N_9263,N_1131,N_2711);
and U9264 (N_9264,N_3672,N_2167);
nand U9265 (N_9265,N_2343,N_777);
nand U9266 (N_9266,N_134,N_254);
nand U9267 (N_9267,N_2302,N_725);
xnor U9268 (N_9268,N_646,N_4268);
nand U9269 (N_9269,N_2966,N_541);
and U9270 (N_9270,N_4505,N_3285);
nor U9271 (N_9271,N_4719,N_464);
and U9272 (N_9272,N_604,N_916);
nand U9273 (N_9273,N_1464,N_4299);
nor U9274 (N_9274,N_4592,N_1961);
or U9275 (N_9275,N_3759,N_3269);
or U9276 (N_9276,N_2822,N_1083);
xnor U9277 (N_9277,N_395,N_2931);
xor U9278 (N_9278,N_1479,N_2960);
and U9279 (N_9279,N_2837,N_4684);
xnor U9280 (N_9280,N_1280,N_390);
or U9281 (N_9281,N_3272,N_87);
nand U9282 (N_9282,N_4206,N_2330);
and U9283 (N_9283,N_4111,N_4596);
xnor U9284 (N_9284,N_2235,N_2026);
xor U9285 (N_9285,N_3305,N_4417);
nor U9286 (N_9286,N_4669,N_3822);
and U9287 (N_9287,N_2008,N_831);
or U9288 (N_9288,N_2985,N_1988);
xnor U9289 (N_9289,N_4386,N_1743);
xnor U9290 (N_9290,N_920,N_2079);
nand U9291 (N_9291,N_45,N_3178);
or U9292 (N_9292,N_1264,N_4410);
xnor U9293 (N_9293,N_1717,N_82);
nor U9294 (N_9294,N_1508,N_1676);
and U9295 (N_9295,N_1374,N_68);
or U9296 (N_9296,N_900,N_2433);
and U9297 (N_9297,N_1978,N_32);
nand U9298 (N_9298,N_216,N_856);
nor U9299 (N_9299,N_664,N_4829);
or U9300 (N_9300,N_799,N_797);
nor U9301 (N_9301,N_3001,N_4490);
nand U9302 (N_9302,N_969,N_3400);
or U9303 (N_9303,N_98,N_997);
or U9304 (N_9304,N_4301,N_2788);
and U9305 (N_9305,N_2364,N_1549);
xnor U9306 (N_9306,N_937,N_1573);
or U9307 (N_9307,N_3156,N_2002);
and U9308 (N_9308,N_3079,N_4554);
nor U9309 (N_9309,N_1033,N_1712);
nor U9310 (N_9310,N_2333,N_4810);
nand U9311 (N_9311,N_2376,N_4427);
and U9312 (N_9312,N_1282,N_4791);
nor U9313 (N_9313,N_1803,N_2246);
xnor U9314 (N_9314,N_1650,N_3032);
xor U9315 (N_9315,N_2521,N_4277);
and U9316 (N_9316,N_1946,N_2549);
and U9317 (N_9317,N_4370,N_4878);
nand U9318 (N_9318,N_4781,N_4716);
xor U9319 (N_9319,N_1649,N_1760);
nand U9320 (N_9320,N_4733,N_601);
or U9321 (N_9321,N_3109,N_1361);
and U9322 (N_9322,N_4426,N_4380);
xnor U9323 (N_9323,N_4944,N_744);
xnor U9324 (N_9324,N_1697,N_4068);
and U9325 (N_9325,N_4872,N_2173);
nand U9326 (N_9326,N_233,N_1463);
or U9327 (N_9327,N_1800,N_2906);
nor U9328 (N_9328,N_177,N_2955);
xor U9329 (N_9329,N_4639,N_2439);
xor U9330 (N_9330,N_3185,N_1076);
nor U9331 (N_9331,N_3523,N_985);
nand U9332 (N_9332,N_415,N_3714);
and U9333 (N_9333,N_3266,N_1579);
and U9334 (N_9334,N_4186,N_4048);
or U9335 (N_9335,N_112,N_251);
nor U9336 (N_9336,N_537,N_1317);
xnor U9337 (N_9337,N_4428,N_1922);
nor U9338 (N_9338,N_878,N_30);
or U9339 (N_9339,N_827,N_398);
xnor U9340 (N_9340,N_4440,N_2719);
nand U9341 (N_9341,N_4776,N_3513);
xnor U9342 (N_9342,N_4409,N_266);
nand U9343 (N_9343,N_2705,N_1144);
or U9344 (N_9344,N_1042,N_3530);
nor U9345 (N_9345,N_2603,N_1879);
nand U9346 (N_9346,N_525,N_4059);
and U9347 (N_9347,N_2631,N_3567);
or U9348 (N_9348,N_503,N_4665);
or U9349 (N_9349,N_2378,N_2599);
or U9350 (N_9350,N_305,N_4569);
and U9351 (N_9351,N_958,N_4564);
or U9352 (N_9352,N_1635,N_2965);
nor U9353 (N_9353,N_2515,N_509);
or U9354 (N_9354,N_2006,N_835);
or U9355 (N_9355,N_2134,N_152);
nand U9356 (N_9356,N_2704,N_1521);
xnor U9357 (N_9357,N_4918,N_533);
xnor U9358 (N_9358,N_3888,N_4889);
or U9359 (N_9359,N_2623,N_2643);
or U9360 (N_9360,N_3504,N_597);
or U9361 (N_9361,N_3037,N_4042);
and U9362 (N_9362,N_3848,N_3572);
nand U9363 (N_9363,N_4155,N_68);
xnor U9364 (N_9364,N_3281,N_3395);
or U9365 (N_9365,N_1284,N_1760);
nand U9366 (N_9366,N_2842,N_4308);
nor U9367 (N_9367,N_4804,N_3832);
or U9368 (N_9368,N_4932,N_2395);
nor U9369 (N_9369,N_4242,N_1672);
or U9370 (N_9370,N_4301,N_66);
nand U9371 (N_9371,N_4698,N_290);
and U9372 (N_9372,N_4774,N_577);
xnor U9373 (N_9373,N_1461,N_1839);
nand U9374 (N_9374,N_3384,N_4574);
and U9375 (N_9375,N_4116,N_1425);
and U9376 (N_9376,N_495,N_4553);
nor U9377 (N_9377,N_2775,N_4120);
nor U9378 (N_9378,N_4583,N_2053);
xnor U9379 (N_9379,N_1035,N_2710);
xnor U9380 (N_9380,N_4225,N_4981);
nand U9381 (N_9381,N_3233,N_922);
nand U9382 (N_9382,N_3741,N_3004);
xnor U9383 (N_9383,N_1763,N_4733);
or U9384 (N_9384,N_2427,N_1925);
nand U9385 (N_9385,N_479,N_4166);
xnor U9386 (N_9386,N_3000,N_1938);
nor U9387 (N_9387,N_2924,N_937);
or U9388 (N_9388,N_101,N_1508);
nand U9389 (N_9389,N_3051,N_1209);
or U9390 (N_9390,N_2994,N_2481);
and U9391 (N_9391,N_2713,N_4129);
nor U9392 (N_9392,N_1580,N_1667);
xnor U9393 (N_9393,N_3583,N_4014);
nand U9394 (N_9394,N_4240,N_2810);
nand U9395 (N_9395,N_4208,N_3496);
nand U9396 (N_9396,N_4378,N_3535);
and U9397 (N_9397,N_4087,N_4781);
or U9398 (N_9398,N_2913,N_1277);
and U9399 (N_9399,N_804,N_3204);
and U9400 (N_9400,N_537,N_3989);
nor U9401 (N_9401,N_845,N_4419);
nand U9402 (N_9402,N_3659,N_1967);
xor U9403 (N_9403,N_996,N_1363);
and U9404 (N_9404,N_1981,N_1192);
or U9405 (N_9405,N_1315,N_4292);
xor U9406 (N_9406,N_1372,N_3906);
nand U9407 (N_9407,N_157,N_2592);
nor U9408 (N_9408,N_3529,N_538);
xnor U9409 (N_9409,N_1270,N_1178);
xor U9410 (N_9410,N_3979,N_1486);
nor U9411 (N_9411,N_4444,N_3012);
and U9412 (N_9412,N_1837,N_2943);
nand U9413 (N_9413,N_4100,N_3147);
or U9414 (N_9414,N_1528,N_2147);
nor U9415 (N_9415,N_4773,N_4718);
xnor U9416 (N_9416,N_4142,N_1201);
or U9417 (N_9417,N_441,N_3258);
nor U9418 (N_9418,N_1948,N_3605);
xor U9419 (N_9419,N_4556,N_1485);
nand U9420 (N_9420,N_1573,N_705);
nor U9421 (N_9421,N_3141,N_4573);
nor U9422 (N_9422,N_1088,N_1362);
or U9423 (N_9423,N_1181,N_1299);
or U9424 (N_9424,N_240,N_4290);
nor U9425 (N_9425,N_2521,N_2007);
nand U9426 (N_9426,N_3417,N_3885);
or U9427 (N_9427,N_3477,N_4982);
xor U9428 (N_9428,N_4911,N_160);
nand U9429 (N_9429,N_3661,N_1722);
and U9430 (N_9430,N_4944,N_1968);
and U9431 (N_9431,N_521,N_245);
nand U9432 (N_9432,N_3644,N_4825);
and U9433 (N_9433,N_4753,N_176);
nor U9434 (N_9434,N_3695,N_4357);
nor U9435 (N_9435,N_781,N_3047);
and U9436 (N_9436,N_3213,N_498);
and U9437 (N_9437,N_3845,N_4719);
nand U9438 (N_9438,N_1979,N_3066);
nor U9439 (N_9439,N_4576,N_1983);
and U9440 (N_9440,N_4267,N_554);
nor U9441 (N_9441,N_3195,N_3108);
or U9442 (N_9442,N_4039,N_3490);
nor U9443 (N_9443,N_1174,N_728);
or U9444 (N_9444,N_4074,N_1735);
or U9445 (N_9445,N_4354,N_187);
xnor U9446 (N_9446,N_1571,N_3160);
or U9447 (N_9447,N_107,N_1228);
nand U9448 (N_9448,N_4050,N_4356);
xnor U9449 (N_9449,N_321,N_4500);
and U9450 (N_9450,N_713,N_2417);
nor U9451 (N_9451,N_3517,N_1907);
nor U9452 (N_9452,N_1401,N_4823);
nor U9453 (N_9453,N_4409,N_3618);
xnor U9454 (N_9454,N_605,N_2600);
nor U9455 (N_9455,N_1002,N_3707);
nand U9456 (N_9456,N_1304,N_691);
or U9457 (N_9457,N_2669,N_3964);
nor U9458 (N_9458,N_892,N_684);
xor U9459 (N_9459,N_2675,N_2126);
nand U9460 (N_9460,N_2525,N_4339);
nor U9461 (N_9461,N_2734,N_2252);
or U9462 (N_9462,N_729,N_4019);
nor U9463 (N_9463,N_2516,N_1951);
xor U9464 (N_9464,N_3943,N_388);
or U9465 (N_9465,N_3354,N_1841);
nand U9466 (N_9466,N_3840,N_3105);
and U9467 (N_9467,N_1934,N_413);
nand U9468 (N_9468,N_698,N_4624);
nand U9469 (N_9469,N_2958,N_117);
nor U9470 (N_9470,N_4452,N_4610);
xnor U9471 (N_9471,N_3029,N_4384);
or U9472 (N_9472,N_1800,N_4802);
and U9473 (N_9473,N_3591,N_4353);
and U9474 (N_9474,N_2884,N_4837);
xor U9475 (N_9475,N_4751,N_2594);
nand U9476 (N_9476,N_1438,N_4002);
and U9477 (N_9477,N_141,N_4999);
or U9478 (N_9478,N_2457,N_4197);
and U9479 (N_9479,N_2822,N_3597);
nor U9480 (N_9480,N_877,N_2197);
and U9481 (N_9481,N_260,N_3283);
xor U9482 (N_9482,N_3904,N_4126);
nor U9483 (N_9483,N_4992,N_3987);
nor U9484 (N_9484,N_4278,N_1953);
or U9485 (N_9485,N_4499,N_4120);
xnor U9486 (N_9486,N_1082,N_336);
or U9487 (N_9487,N_492,N_2778);
nor U9488 (N_9488,N_816,N_3565);
or U9489 (N_9489,N_4128,N_1036);
and U9490 (N_9490,N_1774,N_780);
nand U9491 (N_9491,N_3104,N_3548);
nor U9492 (N_9492,N_1017,N_3013);
or U9493 (N_9493,N_3525,N_3437);
and U9494 (N_9494,N_3772,N_407);
nand U9495 (N_9495,N_1084,N_2991);
and U9496 (N_9496,N_4721,N_4921);
and U9497 (N_9497,N_1493,N_4130);
xnor U9498 (N_9498,N_3923,N_1091);
or U9499 (N_9499,N_4441,N_2075);
and U9500 (N_9500,N_33,N_891);
xnor U9501 (N_9501,N_3220,N_168);
and U9502 (N_9502,N_2721,N_1534);
nor U9503 (N_9503,N_2212,N_1075);
nor U9504 (N_9504,N_600,N_4056);
xor U9505 (N_9505,N_1699,N_4250);
nand U9506 (N_9506,N_4904,N_2719);
or U9507 (N_9507,N_1078,N_841);
xor U9508 (N_9508,N_2621,N_1176);
nand U9509 (N_9509,N_4259,N_637);
nand U9510 (N_9510,N_4045,N_1908);
xnor U9511 (N_9511,N_3470,N_3944);
and U9512 (N_9512,N_1614,N_697);
xor U9513 (N_9513,N_4638,N_3064);
xor U9514 (N_9514,N_4139,N_2830);
xnor U9515 (N_9515,N_1096,N_4230);
and U9516 (N_9516,N_1812,N_1799);
and U9517 (N_9517,N_3393,N_1246);
and U9518 (N_9518,N_3801,N_3211);
or U9519 (N_9519,N_1418,N_4223);
or U9520 (N_9520,N_456,N_3841);
or U9521 (N_9521,N_3772,N_3124);
nor U9522 (N_9522,N_393,N_2466);
or U9523 (N_9523,N_4583,N_4634);
and U9524 (N_9524,N_873,N_3001);
nand U9525 (N_9525,N_3325,N_395);
and U9526 (N_9526,N_4720,N_3337);
xor U9527 (N_9527,N_906,N_557);
nand U9528 (N_9528,N_2830,N_940);
or U9529 (N_9529,N_0,N_71);
xor U9530 (N_9530,N_588,N_249);
nand U9531 (N_9531,N_4872,N_2804);
and U9532 (N_9532,N_25,N_4695);
or U9533 (N_9533,N_3598,N_2319);
nand U9534 (N_9534,N_4513,N_4688);
nor U9535 (N_9535,N_4947,N_43);
xor U9536 (N_9536,N_1525,N_3922);
or U9537 (N_9537,N_1207,N_394);
nor U9538 (N_9538,N_558,N_537);
or U9539 (N_9539,N_4276,N_4981);
nor U9540 (N_9540,N_4861,N_3312);
nand U9541 (N_9541,N_525,N_3647);
nand U9542 (N_9542,N_4009,N_2782);
xnor U9543 (N_9543,N_2798,N_784);
xnor U9544 (N_9544,N_4864,N_672);
nor U9545 (N_9545,N_2710,N_1197);
or U9546 (N_9546,N_2635,N_4235);
or U9547 (N_9547,N_846,N_714);
and U9548 (N_9548,N_3913,N_497);
and U9549 (N_9549,N_4330,N_1648);
nor U9550 (N_9550,N_1430,N_963);
xor U9551 (N_9551,N_3791,N_2740);
xnor U9552 (N_9552,N_179,N_2928);
and U9553 (N_9553,N_3592,N_829);
or U9554 (N_9554,N_1528,N_2615);
nand U9555 (N_9555,N_1654,N_1880);
xnor U9556 (N_9556,N_4435,N_20);
xnor U9557 (N_9557,N_4932,N_2892);
nand U9558 (N_9558,N_2829,N_2013);
nor U9559 (N_9559,N_3153,N_3274);
nor U9560 (N_9560,N_3489,N_4775);
and U9561 (N_9561,N_4813,N_1412);
and U9562 (N_9562,N_2017,N_1280);
nand U9563 (N_9563,N_2365,N_4519);
and U9564 (N_9564,N_2292,N_2560);
nand U9565 (N_9565,N_870,N_4915);
nand U9566 (N_9566,N_1151,N_601);
nand U9567 (N_9567,N_4505,N_3304);
and U9568 (N_9568,N_3555,N_1355);
or U9569 (N_9569,N_1878,N_4272);
nor U9570 (N_9570,N_4396,N_614);
nand U9571 (N_9571,N_396,N_2561);
xor U9572 (N_9572,N_3905,N_4792);
and U9573 (N_9573,N_4024,N_20);
nor U9574 (N_9574,N_433,N_1038);
nor U9575 (N_9575,N_868,N_1507);
or U9576 (N_9576,N_2010,N_281);
or U9577 (N_9577,N_1700,N_3734);
nor U9578 (N_9578,N_400,N_3085);
or U9579 (N_9579,N_2892,N_1338);
nand U9580 (N_9580,N_3906,N_3389);
nor U9581 (N_9581,N_3778,N_4923);
or U9582 (N_9582,N_1426,N_4317);
nand U9583 (N_9583,N_279,N_707);
and U9584 (N_9584,N_1807,N_473);
nand U9585 (N_9585,N_2464,N_606);
nand U9586 (N_9586,N_39,N_4217);
nand U9587 (N_9587,N_3334,N_2403);
nor U9588 (N_9588,N_1040,N_2465);
xor U9589 (N_9589,N_4215,N_3088);
nand U9590 (N_9590,N_4790,N_235);
nand U9591 (N_9591,N_3387,N_953);
nor U9592 (N_9592,N_47,N_1175);
or U9593 (N_9593,N_1123,N_1085);
or U9594 (N_9594,N_1799,N_3025);
nand U9595 (N_9595,N_638,N_589);
nor U9596 (N_9596,N_4818,N_682);
nor U9597 (N_9597,N_4599,N_763);
or U9598 (N_9598,N_3221,N_967);
nand U9599 (N_9599,N_2209,N_2746);
nor U9600 (N_9600,N_2044,N_545);
and U9601 (N_9601,N_2002,N_3970);
xor U9602 (N_9602,N_2306,N_1041);
and U9603 (N_9603,N_19,N_739);
and U9604 (N_9604,N_2235,N_3959);
nor U9605 (N_9605,N_468,N_2509);
xor U9606 (N_9606,N_2727,N_608);
and U9607 (N_9607,N_4445,N_3740);
or U9608 (N_9608,N_1176,N_2501);
and U9609 (N_9609,N_4792,N_1640);
xor U9610 (N_9610,N_4217,N_4629);
or U9611 (N_9611,N_6,N_4953);
nor U9612 (N_9612,N_2086,N_2906);
nor U9613 (N_9613,N_1574,N_3052);
and U9614 (N_9614,N_1468,N_362);
nor U9615 (N_9615,N_1780,N_3621);
nand U9616 (N_9616,N_3021,N_3098);
or U9617 (N_9617,N_68,N_445);
nor U9618 (N_9618,N_3751,N_4800);
nor U9619 (N_9619,N_1744,N_4107);
or U9620 (N_9620,N_3609,N_2775);
nand U9621 (N_9621,N_395,N_93);
or U9622 (N_9622,N_3159,N_1520);
nor U9623 (N_9623,N_181,N_4624);
or U9624 (N_9624,N_1023,N_1782);
and U9625 (N_9625,N_2748,N_4816);
nand U9626 (N_9626,N_1836,N_2168);
xnor U9627 (N_9627,N_591,N_2488);
or U9628 (N_9628,N_4947,N_105);
or U9629 (N_9629,N_4624,N_3360);
nand U9630 (N_9630,N_4378,N_1939);
xnor U9631 (N_9631,N_3030,N_3354);
xnor U9632 (N_9632,N_3254,N_2395);
nand U9633 (N_9633,N_2426,N_15);
nand U9634 (N_9634,N_380,N_4557);
nand U9635 (N_9635,N_3087,N_463);
nand U9636 (N_9636,N_4490,N_2108);
nor U9637 (N_9637,N_3451,N_558);
or U9638 (N_9638,N_4147,N_1369);
or U9639 (N_9639,N_703,N_4811);
nor U9640 (N_9640,N_1402,N_3455);
or U9641 (N_9641,N_4353,N_2524);
xnor U9642 (N_9642,N_1873,N_2717);
xnor U9643 (N_9643,N_2788,N_1341);
and U9644 (N_9644,N_2250,N_2040);
and U9645 (N_9645,N_383,N_1099);
nand U9646 (N_9646,N_4623,N_1086);
xor U9647 (N_9647,N_1103,N_4422);
nor U9648 (N_9648,N_2318,N_4278);
xor U9649 (N_9649,N_3960,N_3407);
and U9650 (N_9650,N_2912,N_1202);
nor U9651 (N_9651,N_3472,N_1851);
and U9652 (N_9652,N_2610,N_1964);
or U9653 (N_9653,N_1172,N_3199);
nor U9654 (N_9654,N_3654,N_3961);
nor U9655 (N_9655,N_4040,N_1507);
xor U9656 (N_9656,N_2503,N_3194);
or U9657 (N_9657,N_3815,N_2431);
xnor U9658 (N_9658,N_3799,N_1174);
xnor U9659 (N_9659,N_1395,N_4031);
or U9660 (N_9660,N_2583,N_735);
or U9661 (N_9661,N_173,N_1639);
nor U9662 (N_9662,N_1999,N_2055);
and U9663 (N_9663,N_4217,N_4936);
xor U9664 (N_9664,N_201,N_2911);
xnor U9665 (N_9665,N_1600,N_2310);
or U9666 (N_9666,N_1564,N_4492);
nor U9667 (N_9667,N_4680,N_4030);
or U9668 (N_9668,N_1813,N_859);
xor U9669 (N_9669,N_1255,N_190);
and U9670 (N_9670,N_2843,N_2314);
nor U9671 (N_9671,N_1526,N_3377);
or U9672 (N_9672,N_2214,N_2228);
or U9673 (N_9673,N_1700,N_1658);
and U9674 (N_9674,N_4700,N_2262);
nor U9675 (N_9675,N_2205,N_2255);
nor U9676 (N_9676,N_3324,N_4274);
nor U9677 (N_9677,N_1384,N_2283);
and U9678 (N_9678,N_4127,N_2318);
nand U9679 (N_9679,N_481,N_1801);
and U9680 (N_9680,N_4480,N_4632);
and U9681 (N_9681,N_842,N_676);
or U9682 (N_9682,N_2057,N_4615);
and U9683 (N_9683,N_68,N_4924);
nor U9684 (N_9684,N_2261,N_4824);
or U9685 (N_9685,N_3,N_3580);
nor U9686 (N_9686,N_780,N_4426);
nor U9687 (N_9687,N_3968,N_1809);
and U9688 (N_9688,N_67,N_3410);
or U9689 (N_9689,N_3099,N_2380);
and U9690 (N_9690,N_3582,N_3015);
and U9691 (N_9691,N_4062,N_1102);
nand U9692 (N_9692,N_1729,N_154);
nor U9693 (N_9693,N_4430,N_3941);
nand U9694 (N_9694,N_3919,N_3523);
or U9695 (N_9695,N_3406,N_4037);
nor U9696 (N_9696,N_1249,N_3262);
nand U9697 (N_9697,N_2095,N_2044);
and U9698 (N_9698,N_4990,N_3584);
nand U9699 (N_9699,N_4181,N_4223);
or U9700 (N_9700,N_1933,N_1299);
xor U9701 (N_9701,N_3523,N_767);
xor U9702 (N_9702,N_3791,N_2785);
nor U9703 (N_9703,N_2750,N_757);
nor U9704 (N_9704,N_2427,N_1477);
nor U9705 (N_9705,N_2741,N_4879);
nor U9706 (N_9706,N_3847,N_4622);
xor U9707 (N_9707,N_1529,N_1682);
or U9708 (N_9708,N_290,N_1765);
nor U9709 (N_9709,N_2319,N_2986);
nor U9710 (N_9710,N_369,N_88);
and U9711 (N_9711,N_940,N_1220);
xor U9712 (N_9712,N_1375,N_618);
nor U9713 (N_9713,N_340,N_4727);
and U9714 (N_9714,N_228,N_1792);
nand U9715 (N_9715,N_1921,N_948);
or U9716 (N_9716,N_2760,N_1135);
nand U9717 (N_9717,N_1752,N_857);
nand U9718 (N_9718,N_4528,N_884);
nor U9719 (N_9719,N_2929,N_442);
nor U9720 (N_9720,N_1688,N_1507);
xnor U9721 (N_9721,N_1035,N_4059);
nor U9722 (N_9722,N_4743,N_51);
nand U9723 (N_9723,N_3455,N_4284);
nor U9724 (N_9724,N_4391,N_1057);
xor U9725 (N_9725,N_777,N_3050);
xor U9726 (N_9726,N_3422,N_4609);
xor U9727 (N_9727,N_4498,N_4461);
or U9728 (N_9728,N_1908,N_4108);
nor U9729 (N_9729,N_3951,N_783);
xor U9730 (N_9730,N_2484,N_161);
nor U9731 (N_9731,N_4675,N_1211);
xor U9732 (N_9732,N_3709,N_2563);
nand U9733 (N_9733,N_323,N_3612);
and U9734 (N_9734,N_2975,N_2799);
xnor U9735 (N_9735,N_880,N_1424);
nand U9736 (N_9736,N_472,N_2776);
or U9737 (N_9737,N_3189,N_837);
and U9738 (N_9738,N_2120,N_736);
nor U9739 (N_9739,N_2793,N_1159);
xnor U9740 (N_9740,N_3985,N_4632);
nand U9741 (N_9741,N_1881,N_3459);
or U9742 (N_9742,N_1409,N_2046);
xnor U9743 (N_9743,N_4444,N_1129);
nor U9744 (N_9744,N_1744,N_3904);
nor U9745 (N_9745,N_4311,N_3345);
nand U9746 (N_9746,N_2243,N_4969);
and U9747 (N_9747,N_269,N_3);
nand U9748 (N_9748,N_2465,N_4010);
nand U9749 (N_9749,N_3572,N_4069);
and U9750 (N_9750,N_2735,N_1067);
nor U9751 (N_9751,N_2105,N_4964);
xor U9752 (N_9752,N_4050,N_167);
xor U9753 (N_9753,N_729,N_4204);
or U9754 (N_9754,N_857,N_2386);
xor U9755 (N_9755,N_3480,N_1726);
nor U9756 (N_9756,N_2298,N_2417);
nand U9757 (N_9757,N_4632,N_4658);
nor U9758 (N_9758,N_2604,N_86);
nor U9759 (N_9759,N_3692,N_4901);
or U9760 (N_9760,N_3959,N_3887);
and U9761 (N_9761,N_1623,N_4262);
xnor U9762 (N_9762,N_4207,N_3228);
xor U9763 (N_9763,N_1843,N_597);
nand U9764 (N_9764,N_561,N_2186);
or U9765 (N_9765,N_4404,N_635);
and U9766 (N_9766,N_727,N_76);
and U9767 (N_9767,N_2327,N_1245);
or U9768 (N_9768,N_2979,N_3225);
nand U9769 (N_9769,N_3367,N_1308);
xor U9770 (N_9770,N_3666,N_1650);
and U9771 (N_9771,N_1918,N_3255);
xor U9772 (N_9772,N_448,N_3953);
nand U9773 (N_9773,N_3570,N_4971);
or U9774 (N_9774,N_1250,N_3680);
and U9775 (N_9775,N_1,N_533);
nor U9776 (N_9776,N_1130,N_3907);
xnor U9777 (N_9777,N_457,N_3210);
nand U9778 (N_9778,N_3579,N_2957);
and U9779 (N_9779,N_117,N_3939);
nor U9780 (N_9780,N_1150,N_3001);
or U9781 (N_9781,N_3375,N_123);
nor U9782 (N_9782,N_638,N_1888);
or U9783 (N_9783,N_4446,N_300);
or U9784 (N_9784,N_917,N_3954);
or U9785 (N_9785,N_2065,N_2327);
or U9786 (N_9786,N_2414,N_3384);
xor U9787 (N_9787,N_3336,N_514);
nor U9788 (N_9788,N_3952,N_2300);
nand U9789 (N_9789,N_4423,N_133);
and U9790 (N_9790,N_1424,N_1429);
xnor U9791 (N_9791,N_3357,N_4035);
nand U9792 (N_9792,N_466,N_490);
nor U9793 (N_9793,N_429,N_2883);
nor U9794 (N_9794,N_649,N_2328);
and U9795 (N_9795,N_3031,N_2812);
or U9796 (N_9796,N_4712,N_1393);
or U9797 (N_9797,N_3763,N_97);
nor U9798 (N_9798,N_2859,N_216);
nand U9799 (N_9799,N_1621,N_2197);
and U9800 (N_9800,N_1102,N_106);
or U9801 (N_9801,N_1367,N_3212);
and U9802 (N_9802,N_4681,N_2888);
and U9803 (N_9803,N_1272,N_2616);
nor U9804 (N_9804,N_3885,N_3978);
and U9805 (N_9805,N_2649,N_2582);
and U9806 (N_9806,N_3169,N_251);
xnor U9807 (N_9807,N_829,N_360);
xor U9808 (N_9808,N_2553,N_4882);
nor U9809 (N_9809,N_4359,N_3811);
nor U9810 (N_9810,N_2757,N_3811);
nor U9811 (N_9811,N_2133,N_3445);
xor U9812 (N_9812,N_4595,N_3400);
nand U9813 (N_9813,N_1225,N_979);
nand U9814 (N_9814,N_2012,N_3765);
and U9815 (N_9815,N_926,N_1795);
and U9816 (N_9816,N_4316,N_469);
nand U9817 (N_9817,N_4015,N_732);
nor U9818 (N_9818,N_1131,N_749);
nor U9819 (N_9819,N_1369,N_4461);
and U9820 (N_9820,N_3459,N_1439);
xnor U9821 (N_9821,N_1746,N_3429);
xnor U9822 (N_9822,N_610,N_4619);
or U9823 (N_9823,N_1190,N_1939);
xnor U9824 (N_9824,N_1145,N_4952);
and U9825 (N_9825,N_1145,N_3452);
nand U9826 (N_9826,N_1380,N_3123);
or U9827 (N_9827,N_642,N_2745);
nand U9828 (N_9828,N_3232,N_2224);
nor U9829 (N_9829,N_1270,N_4667);
nand U9830 (N_9830,N_3117,N_553);
and U9831 (N_9831,N_4196,N_2003);
nand U9832 (N_9832,N_1361,N_1766);
and U9833 (N_9833,N_2169,N_2894);
and U9834 (N_9834,N_142,N_513);
or U9835 (N_9835,N_3328,N_4166);
or U9836 (N_9836,N_3632,N_482);
nor U9837 (N_9837,N_473,N_776);
xor U9838 (N_9838,N_1340,N_3031);
nor U9839 (N_9839,N_2109,N_217);
nor U9840 (N_9840,N_3632,N_1665);
and U9841 (N_9841,N_58,N_2948);
nand U9842 (N_9842,N_1595,N_803);
and U9843 (N_9843,N_3276,N_1478);
nand U9844 (N_9844,N_3395,N_1452);
nor U9845 (N_9845,N_2162,N_2844);
or U9846 (N_9846,N_1566,N_2986);
nand U9847 (N_9847,N_1628,N_3126);
or U9848 (N_9848,N_2576,N_4265);
nand U9849 (N_9849,N_386,N_4177);
xor U9850 (N_9850,N_40,N_3584);
and U9851 (N_9851,N_263,N_213);
nand U9852 (N_9852,N_2457,N_4757);
or U9853 (N_9853,N_2744,N_1591);
nor U9854 (N_9854,N_1639,N_451);
and U9855 (N_9855,N_4181,N_1953);
xor U9856 (N_9856,N_3693,N_804);
and U9857 (N_9857,N_2384,N_3309);
nor U9858 (N_9858,N_3664,N_3088);
nor U9859 (N_9859,N_27,N_3283);
or U9860 (N_9860,N_3542,N_2297);
nor U9861 (N_9861,N_2264,N_2009);
and U9862 (N_9862,N_973,N_248);
nor U9863 (N_9863,N_2528,N_790);
and U9864 (N_9864,N_2916,N_2457);
nand U9865 (N_9865,N_1251,N_2434);
nor U9866 (N_9866,N_1184,N_3524);
and U9867 (N_9867,N_3497,N_519);
or U9868 (N_9868,N_3393,N_4809);
and U9869 (N_9869,N_4685,N_3838);
and U9870 (N_9870,N_2706,N_3349);
xor U9871 (N_9871,N_3951,N_2608);
nand U9872 (N_9872,N_474,N_2235);
xor U9873 (N_9873,N_333,N_3428);
nand U9874 (N_9874,N_873,N_1864);
and U9875 (N_9875,N_1844,N_60);
or U9876 (N_9876,N_1916,N_32);
xor U9877 (N_9877,N_655,N_2703);
nand U9878 (N_9878,N_4998,N_4226);
xnor U9879 (N_9879,N_3718,N_2687);
nand U9880 (N_9880,N_3157,N_1039);
and U9881 (N_9881,N_237,N_4225);
and U9882 (N_9882,N_3395,N_3526);
nor U9883 (N_9883,N_2172,N_803);
xnor U9884 (N_9884,N_1766,N_4550);
or U9885 (N_9885,N_4277,N_1332);
and U9886 (N_9886,N_3124,N_3987);
nor U9887 (N_9887,N_554,N_1187);
or U9888 (N_9888,N_2903,N_513);
nor U9889 (N_9889,N_4540,N_804);
xor U9890 (N_9890,N_3151,N_3114);
nand U9891 (N_9891,N_2742,N_1481);
nand U9892 (N_9892,N_3322,N_2834);
nand U9893 (N_9893,N_4271,N_1809);
or U9894 (N_9894,N_662,N_2016);
or U9895 (N_9895,N_2019,N_3246);
or U9896 (N_9896,N_4102,N_3158);
xor U9897 (N_9897,N_3408,N_3104);
or U9898 (N_9898,N_3631,N_3252);
nor U9899 (N_9899,N_1788,N_3032);
xor U9900 (N_9900,N_3297,N_3188);
and U9901 (N_9901,N_2768,N_46);
nand U9902 (N_9902,N_3119,N_4574);
and U9903 (N_9903,N_959,N_4308);
and U9904 (N_9904,N_4639,N_4271);
nand U9905 (N_9905,N_4053,N_3142);
nand U9906 (N_9906,N_3188,N_1255);
nor U9907 (N_9907,N_2971,N_4664);
nor U9908 (N_9908,N_3820,N_2572);
xor U9909 (N_9909,N_982,N_523);
or U9910 (N_9910,N_2101,N_2978);
nor U9911 (N_9911,N_3699,N_4693);
nor U9912 (N_9912,N_4533,N_4068);
nand U9913 (N_9913,N_4887,N_4488);
nor U9914 (N_9914,N_461,N_268);
xnor U9915 (N_9915,N_2365,N_3636);
and U9916 (N_9916,N_4581,N_3143);
nor U9917 (N_9917,N_438,N_4413);
nor U9918 (N_9918,N_2227,N_2092);
nand U9919 (N_9919,N_3925,N_3246);
and U9920 (N_9920,N_4065,N_2018);
nand U9921 (N_9921,N_3777,N_1391);
xnor U9922 (N_9922,N_2123,N_2748);
or U9923 (N_9923,N_3396,N_1016);
xnor U9924 (N_9924,N_2910,N_4880);
nor U9925 (N_9925,N_4882,N_121);
and U9926 (N_9926,N_1047,N_1205);
xnor U9927 (N_9927,N_2969,N_1874);
nand U9928 (N_9928,N_4314,N_2666);
xor U9929 (N_9929,N_1188,N_854);
or U9930 (N_9930,N_684,N_497);
nor U9931 (N_9931,N_887,N_4642);
xnor U9932 (N_9932,N_4132,N_479);
and U9933 (N_9933,N_2261,N_4358);
nand U9934 (N_9934,N_3842,N_4218);
nand U9935 (N_9935,N_1106,N_3007);
xnor U9936 (N_9936,N_1566,N_1138);
xnor U9937 (N_9937,N_2693,N_3398);
or U9938 (N_9938,N_1103,N_2306);
nand U9939 (N_9939,N_857,N_1208);
and U9940 (N_9940,N_2523,N_2619);
and U9941 (N_9941,N_1751,N_3223);
and U9942 (N_9942,N_4696,N_4961);
xnor U9943 (N_9943,N_1036,N_3022);
nor U9944 (N_9944,N_1083,N_1450);
or U9945 (N_9945,N_3787,N_114);
nand U9946 (N_9946,N_1466,N_3678);
nor U9947 (N_9947,N_1017,N_2676);
nand U9948 (N_9948,N_1537,N_4724);
nor U9949 (N_9949,N_4145,N_1180);
nor U9950 (N_9950,N_2510,N_1706);
or U9951 (N_9951,N_1220,N_182);
or U9952 (N_9952,N_1286,N_3370);
xor U9953 (N_9953,N_3589,N_2069);
or U9954 (N_9954,N_292,N_4937);
or U9955 (N_9955,N_4128,N_2118);
and U9956 (N_9956,N_4070,N_798);
xnor U9957 (N_9957,N_3524,N_3384);
xor U9958 (N_9958,N_2550,N_4422);
and U9959 (N_9959,N_2791,N_2893);
or U9960 (N_9960,N_2848,N_1522);
and U9961 (N_9961,N_4400,N_1665);
xor U9962 (N_9962,N_3071,N_4223);
or U9963 (N_9963,N_580,N_891);
and U9964 (N_9964,N_1243,N_169);
and U9965 (N_9965,N_883,N_3141);
xnor U9966 (N_9966,N_1588,N_4029);
nor U9967 (N_9967,N_717,N_1486);
xor U9968 (N_9968,N_4177,N_4365);
or U9969 (N_9969,N_1137,N_4458);
xnor U9970 (N_9970,N_4542,N_3915);
xor U9971 (N_9971,N_655,N_546);
and U9972 (N_9972,N_2425,N_691);
xnor U9973 (N_9973,N_1125,N_3743);
xor U9974 (N_9974,N_2049,N_1534);
and U9975 (N_9975,N_401,N_4937);
or U9976 (N_9976,N_4382,N_3103);
nand U9977 (N_9977,N_2656,N_2987);
and U9978 (N_9978,N_2940,N_2560);
nand U9979 (N_9979,N_1214,N_328);
xnor U9980 (N_9980,N_679,N_3098);
nor U9981 (N_9981,N_4687,N_2007);
nor U9982 (N_9982,N_4569,N_217);
nor U9983 (N_9983,N_2100,N_3769);
or U9984 (N_9984,N_634,N_175);
xor U9985 (N_9985,N_1484,N_1817);
xnor U9986 (N_9986,N_1626,N_793);
nor U9987 (N_9987,N_2519,N_1347);
nor U9988 (N_9988,N_2336,N_1952);
nand U9989 (N_9989,N_1803,N_3016);
nand U9990 (N_9990,N_574,N_2902);
nor U9991 (N_9991,N_1571,N_3532);
nor U9992 (N_9992,N_2755,N_2980);
nand U9993 (N_9993,N_4723,N_3806);
or U9994 (N_9994,N_1894,N_438);
and U9995 (N_9995,N_395,N_2759);
and U9996 (N_9996,N_4891,N_3034);
or U9997 (N_9997,N_4462,N_3428);
xnor U9998 (N_9998,N_4109,N_2782);
and U9999 (N_9999,N_1197,N_4152);
nand U10000 (N_10000,N_7930,N_8399);
or U10001 (N_10001,N_9992,N_5725);
nor U10002 (N_10002,N_5420,N_5871);
or U10003 (N_10003,N_5796,N_6670);
or U10004 (N_10004,N_7707,N_8384);
nand U10005 (N_10005,N_5132,N_5357);
xnor U10006 (N_10006,N_8876,N_7058);
or U10007 (N_10007,N_7284,N_5947);
or U10008 (N_10008,N_8636,N_5605);
nor U10009 (N_10009,N_9211,N_6154);
xor U10010 (N_10010,N_7195,N_5957);
or U10011 (N_10011,N_8363,N_8905);
xnor U10012 (N_10012,N_5027,N_8612);
nor U10013 (N_10013,N_5421,N_7562);
and U10014 (N_10014,N_5496,N_8179);
nor U10015 (N_10015,N_6287,N_7504);
and U10016 (N_10016,N_7053,N_9934);
nand U10017 (N_10017,N_5094,N_8855);
nor U10018 (N_10018,N_7498,N_8209);
or U10019 (N_10019,N_8134,N_9837);
nor U10020 (N_10020,N_9898,N_9144);
nand U10021 (N_10021,N_8624,N_9330);
nor U10022 (N_10022,N_5278,N_8843);
nand U10023 (N_10023,N_7290,N_6948);
nor U10024 (N_10024,N_5855,N_6821);
and U10025 (N_10025,N_9410,N_8727);
nor U10026 (N_10026,N_8037,N_8819);
or U10027 (N_10027,N_6686,N_5151);
or U10028 (N_10028,N_9959,N_5021);
xor U10029 (N_10029,N_8758,N_9700);
nand U10030 (N_10030,N_6945,N_9301);
xor U10031 (N_10031,N_6045,N_5713);
xnor U10032 (N_10032,N_9504,N_5237);
nor U10033 (N_10033,N_7600,N_6743);
and U10034 (N_10034,N_9522,N_9253);
nand U10035 (N_10035,N_5490,N_8341);
nor U10036 (N_10036,N_5958,N_9053);
nand U10037 (N_10037,N_8487,N_9220);
or U10038 (N_10038,N_7673,N_8967);
or U10039 (N_10039,N_9237,N_7703);
or U10040 (N_10040,N_7887,N_9668);
nand U10041 (N_10041,N_8452,N_5146);
and U10042 (N_10042,N_6611,N_6121);
xnor U10043 (N_10043,N_5747,N_7704);
xor U10044 (N_10044,N_9641,N_5083);
nand U10045 (N_10045,N_6549,N_5281);
nand U10046 (N_10046,N_9938,N_8733);
and U10047 (N_10047,N_7386,N_8842);
and U10048 (N_10048,N_6851,N_9126);
nor U10049 (N_10049,N_7784,N_9247);
xnor U10050 (N_10050,N_9267,N_8949);
or U10051 (N_10051,N_9776,N_6243);
and U10052 (N_10052,N_5939,N_9475);
and U10053 (N_10053,N_7796,N_9532);
nand U10054 (N_10054,N_9678,N_6270);
nor U10055 (N_10055,N_5750,N_7370);
nor U10056 (N_10056,N_6685,N_5202);
and U10057 (N_10057,N_7235,N_7805);
nor U10058 (N_10058,N_7964,N_6845);
xnor U10059 (N_10059,N_8262,N_5693);
xor U10060 (N_10060,N_9850,N_5509);
xor U10061 (N_10061,N_9270,N_6667);
nand U10062 (N_10062,N_8306,N_9203);
and U10063 (N_10063,N_9390,N_9361);
or U10064 (N_10064,N_5308,N_8307);
nor U10065 (N_10065,N_7924,N_7438);
nand U10066 (N_10066,N_6252,N_8464);
xor U10067 (N_10067,N_5609,N_6759);
nor U10068 (N_10068,N_9179,N_5158);
nand U10069 (N_10069,N_9396,N_9230);
xnor U10070 (N_10070,N_7179,N_9561);
nor U10071 (N_10071,N_6340,N_5786);
and U10072 (N_10072,N_8995,N_7900);
xor U10073 (N_10073,N_9474,N_5676);
and U10074 (N_10074,N_6646,N_7789);
nor U10075 (N_10075,N_8635,N_9737);
and U10076 (N_10076,N_8069,N_9427);
xor U10077 (N_10077,N_8570,N_5839);
and U10078 (N_10078,N_6324,N_6242);
nand U10079 (N_10079,N_6001,N_5730);
nand U10080 (N_10080,N_9356,N_9659);
nand U10081 (N_10081,N_6145,N_6099);
nand U10082 (N_10082,N_6582,N_5238);
and U10083 (N_10083,N_6942,N_7208);
or U10084 (N_10084,N_5209,N_5296);
or U10085 (N_10085,N_8008,N_6820);
nor U10086 (N_10086,N_9242,N_9785);
and U10087 (N_10087,N_8327,N_7330);
and U10088 (N_10088,N_7361,N_6379);
and U10089 (N_10089,N_6296,N_7050);
and U10090 (N_10090,N_7170,N_9176);
or U10091 (N_10091,N_6216,N_9452);
and U10092 (N_10092,N_9285,N_5440);
and U10093 (N_10093,N_5683,N_6407);
nand U10094 (N_10094,N_9338,N_5689);
nand U10095 (N_10095,N_9064,N_5803);
nand U10096 (N_10096,N_6568,N_9949);
and U10097 (N_10097,N_7795,N_7176);
or U10098 (N_10098,N_7452,N_8868);
and U10099 (N_10099,N_7077,N_9988);
xor U10100 (N_10100,N_9600,N_7610);
and U10101 (N_10101,N_5459,N_9088);
and U10102 (N_10102,N_9863,N_8766);
xnor U10103 (N_10103,N_6372,N_8551);
xor U10104 (N_10104,N_6450,N_7635);
or U10105 (N_10105,N_6536,N_5731);
nand U10106 (N_10106,N_7872,N_6992);
or U10107 (N_10107,N_9403,N_9734);
or U10108 (N_10108,N_9888,N_6912);
nand U10109 (N_10109,N_5040,N_8197);
xnor U10110 (N_10110,N_9735,N_6239);
xor U10111 (N_10111,N_6694,N_5156);
xor U10112 (N_10112,N_5716,N_5612);
nor U10113 (N_10113,N_8161,N_7861);
nor U10114 (N_10114,N_9298,N_5611);
and U10115 (N_10115,N_7751,N_8491);
or U10116 (N_10116,N_7448,N_7993);
nor U10117 (N_10117,N_7803,N_7634);
nor U10118 (N_10118,N_8779,N_8050);
and U10119 (N_10119,N_8128,N_5243);
or U10120 (N_10120,N_9823,N_5899);
nor U10121 (N_10121,N_6342,N_7305);
xnor U10122 (N_10122,N_5236,N_8309);
and U10123 (N_10123,N_7519,N_5629);
or U10124 (N_10124,N_7379,N_7340);
nand U10125 (N_10125,N_7479,N_7173);
xor U10126 (N_10126,N_9508,N_9261);
or U10127 (N_10127,N_6018,N_9548);
and U10128 (N_10128,N_5301,N_9494);
nor U10129 (N_10129,N_6838,N_9894);
nand U10130 (N_10130,N_6853,N_7891);
and U10131 (N_10131,N_9759,N_7264);
and U10132 (N_10132,N_5869,N_9484);
and U10133 (N_10133,N_6292,N_5379);
nor U10134 (N_10134,N_5170,N_9831);
and U10135 (N_10135,N_7163,N_6002);
or U10136 (N_10136,N_6237,N_6614);
and U10137 (N_10137,N_5632,N_6333);
nor U10138 (N_10138,N_5257,N_5251);
xor U10139 (N_10139,N_6155,N_8597);
nand U10140 (N_10140,N_5789,N_9931);
and U10141 (N_10141,N_9792,N_7916);
and U10142 (N_10142,N_9882,N_5726);
or U10143 (N_10143,N_9841,N_9987);
nor U10144 (N_10144,N_8874,N_8291);
nand U10145 (N_10145,N_7197,N_8129);
and U10146 (N_10146,N_5322,N_8342);
nor U10147 (N_10147,N_7856,N_5906);
and U10148 (N_10148,N_7490,N_8567);
nor U10149 (N_10149,N_8418,N_7758);
nand U10150 (N_10150,N_6166,N_8755);
or U10151 (N_10151,N_6585,N_8155);
nor U10152 (N_10152,N_6390,N_7503);
and U10153 (N_10153,N_8783,N_7183);
xor U10154 (N_10154,N_8976,N_7339);
nor U10155 (N_10155,N_8709,N_5453);
and U10156 (N_10156,N_8998,N_5902);
nor U10157 (N_10157,N_6057,N_6870);
xnor U10158 (N_10158,N_8912,N_6225);
nand U10159 (N_10159,N_6291,N_8360);
xor U10160 (N_10160,N_8102,N_8238);
nand U10161 (N_10161,N_5804,N_8365);
nand U10162 (N_10162,N_7478,N_9736);
nand U10163 (N_10163,N_5401,N_7540);
xnor U10164 (N_10164,N_5633,N_5074);
xor U10165 (N_10165,N_7699,N_6055);
and U10166 (N_10166,N_7010,N_5386);
nand U10167 (N_10167,N_6832,N_6565);
or U10168 (N_10168,N_9535,N_9513);
xnor U10169 (N_10169,N_8939,N_7168);
nand U10170 (N_10170,N_8756,N_9180);
nand U10171 (N_10171,N_8115,N_7701);
and U10172 (N_10172,N_7022,N_6940);
nand U10173 (N_10173,N_9701,N_9777);
nand U10174 (N_10174,N_5193,N_6765);
nor U10175 (N_10175,N_7463,N_9000);
and U10176 (N_10176,N_8642,N_6541);
nor U10177 (N_10177,N_7845,N_5821);
xor U10178 (N_10178,N_5982,N_8334);
nor U10179 (N_10179,N_6959,N_8076);
and U10180 (N_10180,N_7988,N_7282);
nand U10181 (N_10181,N_8798,N_7632);
and U10182 (N_10182,N_8094,N_9957);
nor U10183 (N_10183,N_6530,N_6095);
nor U10184 (N_10184,N_6348,N_5186);
nor U10185 (N_10185,N_6844,N_5177);
or U10186 (N_10186,N_7491,N_9331);
and U10187 (N_10187,N_6757,N_8255);
and U10188 (N_10188,N_9703,N_7897);
nand U10189 (N_10189,N_6518,N_6344);
nor U10190 (N_10190,N_7210,N_7684);
nand U10191 (N_10191,N_9556,N_9101);
nand U10192 (N_10192,N_9585,N_5724);
or U10193 (N_10193,N_8547,N_8282);
nand U10194 (N_10194,N_8204,N_7437);
nor U10195 (N_10195,N_5858,N_5661);
xnor U10196 (N_10196,N_8663,N_8865);
or U10197 (N_10197,N_5521,N_8828);
xor U10198 (N_10198,N_5087,N_6039);
or U10199 (N_10199,N_9541,N_5823);
or U10200 (N_10200,N_7770,N_6978);
and U10201 (N_10201,N_6926,N_7351);
xor U10202 (N_10202,N_6627,N_7298);
and U10203 (N_10203,N_7487,N_6006);
nor U10204 (N_10204,N_9316,N_5447);
nand U10205 (N_10205,N_5403,N_8348);
or U10206 (N_10206,N_8029,N_9621);
or U10207 (N_10207,N_7613,N_6492);
nand U10208 (N_10208,N_7776,N_7692);
xor U10209 (N_10209,N_7798,N_8787);
or U10210 (N_10210,N_9821,N_5540);
xnor U10211 (N_10211,N_9836,N_7651);
nor U10212 (N_10212,N_7569,N_6801);
nor U10213 (N_10213,N_5338,N_5616);
nand U10214 (N_10214,N_9526,N_9334);
and U10215 (N_10215,N_7716,N_9813);
nor U10216 (N_10216,N_8110,N_6590);
and U10217 (N_10217,N_7908,N_6264);
and U10218 (N_10218,N_6920,N_9004);
and U10219 (N_10219,N_7574,N_6502);
or U10220 (N_10220,N_8431,N_8884);
nand U10221 (N_10221,N_7085,N_9090);
xor U10222 (N_10222,N_9583,N_9433);
xnor U10223 (N_10223,N_5976,N_5810);
or U10224 (N_10224,N_5875,N_5212);
and U10225 (N_10225,N_7743,N_9914);
and U10226 (N_10226,N_8379,N_9495);
xnor U10227 (N_10227,N_9842,N_5295);
nor U10228 (N_10228,N_5358,N_7767);
or U10229 (N_10229,N_8894,N_6423);
nor U10230 (N_10230,N_8084,N_7646);
and U10231 (N_10231,N_9281,N_9115);
nand U10232 (N_10232,N_6093,N_6393);
nand U10233 (N_10233,N_5738,N_5783);
and U10234 (N_10234,N_5856,N_5897);
nor U10235 (N_10235,N_6381,N_5797);
nand U10236 (N_10236,N_5334,N_5672);
and U10237 (N_10237,N_5117,N_5526);
xnor U10238 (N_10238,N_8652,N_8757);
nor U10239 (N_10239,N_5828,N_7943);
xnor U10240 (N_10240,N_9861,N_5610);
or U10241 (N_10241,N_8602,N_8982);
or U10242 (N_10242,N_7662,N_8596);
or U10243 (N_10243,N_5964,N_5697);
nor U10244 (N_10244,N_9212,N_7049);
nor U10245 (N_10245,N_5089,N_9069);
or U10246 (N_10246,N_6472,N_7782);
nand U10247 (N_10247,N_6365,N_6513);
and U10248 (N_10248,N_5501,N_8750);
nand U10249 (N_10249,N_6789,N_5949);
and U10250 (N_10250,N_7918,N_6835);
and U10251 (N_10251,N_5511,N_5734);
or U10252 (N_10252,N_9245,N_9071);
or U10253 (N_10253,N_5740,N_8538);
and U10254 (N_10254,N_5977,N_5013);
or U10255 (N_10255,N_5482,N_6418);
xor U10256 (N_10256,N_6280,N_5854);
and U10257 (N_10257,N_6501,N_8732);
or U10258 (N_10258,N_6671,N_7281);
xnor U10259 (N_10259,N_7056,N_6168);
nand U10260 (N_10260,N_9463,N_8614);
or U10261 (N_10261,N_6738,N_7299);
nor U10262 (N_10262,N_5993,N_8346);
nand U10263 (N_10263,N_8562,N_9870);
nand U10264 (N_10264,N_6719,N_8793);
and U10265 (N_10265,N_8242,N_8247);
nand U10266 (N_10266,N_9181,N_7871);
nand U10267 (N_10267,N_8304,N_5688);
nor U10268 (N_10268,N_7094,N_8368);
xnor U10269 (N_10269,N_5116,N_5100);
and U10270 (N_10270,N_7061,N_8677);
nand U10271 (N_10271,N_7655,N_9284);
nand U10272 (N_10272,N_6540,N_8034);
nor U10273 (N_10273,N_5945,N_7799);
or U10274 (N_10274,N_9102,N_8250);
xor U10275 (N_10275,N_9038,N_8981);
nor U10276 (N_10276,N_9848,N_6371);
or U10277 (N_10277,N_9711,N_8469);
or U10278 (N_10278,N_5478,N_7969);
or U10279 (N_10279,N_8513,N_8364);
xor U10280 (N_10280,N_8010,N_9733);
nand U10281 (N_10281,N_5455,N_7753);
or U10282 (N_10282,N_9726,N_8317);
xor U10283 (N_10283,N_6904,N_7890);
nor U10284 (N_10284,N_7260,N_9704);
or U10285 (N_10285,N_5385,N_9928);
or U10286 (N_10286,N_8303,N_9449);
nand U10287 (N_10287,N_6867,N_7862);
nand U10288 (N_10288,N_7737,N_9280);
xor U10289 (N_10289,N_9968,N_5345);
or U10290 (N_10290,N_9956,N_7729);
nor U10291 (N_10291,N_6865,N_9546);
and U10292 (N_10292,N_5306,N_9653);
xnor U10293 (N_10293,N_6566,N_8033);
and U10294 (N_10294,N_5001,N_7189);
nand U10295 (N_10295,N_9650,N_9969);
and U10296 (N_10296,N_5516,N_7378);
nand U10297 (N_10297,N_7267,N_8849);
nand U10298 (N_10298,N_6343,N_9388);
nand U10299 (N_10299,N_9887,N_8668);
and U10300 (N_10300,N_7353,N_8356);
nor U10301 (N_10301,N_9308,N_8457);
nand U10302 (N_10302,N_5293,N_5341);
nor U10303 (N_10303,N_5029,N_6804);
or U10304 (N_10304,N_7879,N_6717);
nor U10305 (N_10305,N_6941,N_6259);
or U10306 (N_10306,N_5229,N_6256);
and U10307 (N_10307,N_8575,N_7786);
xor U10308 (N_10308,N_9033,N_6446);
xor U10309 (N_10309,N_7015,N_8594);
and U10310 (N_10310,N_8739,N_8947);
or U10311 (N_10311,N_9393,N_8227);
or U10312 (N_10312,N_8603,N_9562);
nor U10313 (N_10313,N_5488,N_9244);
and U10314 (N_10314,N_7771,N_6402);
nand U10315 (N_10315,N_9829,N_6636);
and U10316 (N_10316,N_9802,N_7259);
nor U10317 (N_10317,N_8676,N_8377);
or U10318 (N_10318,N_8000,N_9906);
nor U10319 (N_10319,N_6519,N_6183);
or U10320 (N_10320,N_6297,N_7162);
xnor U10321 (N_10321,N_7146,N_7075);
nand U10322 (N_10322,N_5772,N_6211);
and U10323 (N_10323,N_8987,N_9877);
and U10324 (N_10324,N_9438,N_5025);
and U10325 (N_10325,N_6873,N_6293);
nand U10326 (N_10326,N_8460,N_5414);
or U10327 (N_10327,N_7016,N_7395);
xor U10328 (N_10328,N_9807,N_9875);
nand U10329 (N_10329,N_8283,N_5794);
and U10330 (N_10330,N_7164,N_6556);
xor U10331 (N_10331,N_8278,N_8933);
nand U10332 (N_10332,N_9110,N_9275);
and U10333 (N_10333,N_7702,N_5758);
or U10334 (N_10334,N_8999,N_7167);
xor U10335 (N_10335,N_5133,N_7874);
xor U10336 (N_10336,N_6439,N_5220);
xnor U10337 (N_10337,N_6029,N_6315);
xnor U10338 (N_10338,N_6861,N_6983);
nor U10339 (N_10339,N_5072,N_7691);
or U10340 (N_10340,N_5889,N_8300);
and U10341 (N_10341,N_7697,N_7660);
nand U10342 (N_10342,N_8759,N_7265);
xor U10343 (N_10343,N_6080,N_6204);
and U10344 (N_10344,N_8831,N_5573);
nor U10345 (N_10345,N_7787,N_6984);
or U10346 (N_10346,N_5196,N_8274);
nand U10347 (N_10347,N_8133,N_8498);
nand U10348 (N_10348,N_9209,N_8715);
or U10349 (N_10349,N_5266,N_6391);
xor U10350 (N_10350,N_7229,N_8644);
xnor U10351 (N_10351,N_8797,N_7190);
xnor U10352 (N_10352,N_7875,N_5062);
nand U10353 (N_10353,N_7652,N_8272);
nor U10354 (N_10354,N_8634,N_7810);
xnor U10355 (N_10355,N_5272,N_7772);
nor U10356 (N_10356,N_9998,N_8857);
and U10357 (N_10357,N_9922,N_8483);
or U10358 (N_10358,N_5848,N_9415);
nor U10359 (N_10359,N_5290,N_6486);
or U10360 (N_10360,N_5922,N_6149);
nand U10361 (N_10361,N_7790,N_5105);
or U10362 (N_10362,N_6535,N_9116);
and U10363 (N_10363,N_5475,N_5336);
xor U10364 (N_10364,N_7547,N_8295);
nor U10365 (N_10365,N_8434,N_8826);
or U10366 (N_10366,N_9972,N_6895);
nor U10367 (N_10367,N_6633,N_8022);
or U10368 (N_10368,N_6601,N_8692);
xnor U10369 (N_10369,N_7459,N_6461);
xor U10370 (N_10370,N_9442,N_5028);
and U10371 (N_10371,N_5102,N_6950);
nor U10372 (N_10372,N_7937,N_9867);
xnor U10373 (N_10373,N_6755,N_8914);
xnor U10374 (N_10374,N_6629,N_7791);
xor U10375 (N_10375,N_7637,N_7572);
nor U10376 (N_10376,N_5273,N_9486);
and U10377 (N_10377,N_8630,N_8007);
xnor U10378 (N_10378,N_5637,N_6284);
nand U10379 (N_10379,N_6321,N_6298);
or U10380 (N_10380,N_9854,N_7327);
nor U10381 (N_10381,N_6453,N_6786);
xor U10382 (N_10382,N_8293,N_8650);
and U10383 (N_10383,N_9994,N_8904);
nand U10384 (N_10384,N_9414,N_8256);
nor U10385 (N_10385,N_9304,N_5377);
xnor U10386 (N_10386,N_5152,N_5892);
and U10387 (N_10387,N_7069,N_7626);
or U10388 (N_10388,N_7440,N_5477);
nor U10389 (N_10389,N_5168,N_8132);
or U10390 (N_10390,N_5043,N_7566);
nand U10391 (N_10391,N_5349,N_7947);
nor U10392 (N_10392,N_7808,N_7272);
and U10393 (N_10393,N_6330,N_9707);
nor U10394 (N_10394,N_8131,N_6762);
nand U10395 (N_10395,N_8287,N_9691);
nand U10396 (N_10396,N_5569,N_7573);
xor U10397 (N_10397,N_7185,N_6064);
nand U10398 (N_10398,N_5944,N_7466);
and U10399 (N_10399,N_8028,N_9891);
nand U10400 (N_10400,N_7755,N_9603);
nor U10401 (N_10401,N_5571,N_6752);
and U10402 (N_10402,N_6610,N_8073);
or U10403 (N_10403,N_7923,N_8581);
nand U10404 (N_10404,N_6417,N_5798);
and U10405 (N_10405,N_6973,N_5228);
and U10406 (N_10406,N_8527,N_6299);
and U10407 (N_10407,N_9872,N_7232);
xor U10408 (N_10408,N_5389,N_9487);
nor U10409 (N_10409,N_6761,N_7241);
and U10410 (N_10410,N_7246,N_9536);
and U10411 (N_10411,N_8616,N_6131);
and U10412 (N_10412,N_9206,N_6993);
xnor U10413 (N_10413,N_5905,N_5143);
nand U10414 (N_10414,N_6648,N_8396);
or U10415 (N_10415,N_9341,N_9593);
or U10416 (N_10416,N_8956,N_6326);
and U10417 (N_10417,N_8821,N_5805);
and U10418 (N_10418,N_6213,N_8004);
or U10419 (N_10419,N_6124,N_6524);
nand U10420 (N_10420,N_8526,N_8684);
nor U10421 (N_10421,N_5502,N_7922);
nor U10422 (N_10422,N_8977,N_9423);
nand U10423 (N_10423,N_7506,N_7292);
or U10424 (N_10424,N_7268,N_8175);
xnor U10425 (N_10425,N_9811,N_7785);
xnor U10426 (N_10426,N_6400,N_5617);
nand U10427 (N_10427,N_6947,N_5224);
xor U10428 (N_10428,N_9873,N_5064);
and U10429 (N_10429,N_9571,N_9213);
xnor U10430 (N_10430,N_6014,N_6958);
nand U10431 (N_10431,N_6936,N_6431);
nor U10432 (N_10432,N_8560,N_8862);
and U10433 (N_10433,N_7417,N_5739);
nand U10434 (N_10434,N_6864,N_5325);
and U10435 (N_10435,N_8276,N_8711);
or U10436 (N_10436,N_6327,N_9772);
and U10437 (N_10437,N_5621,N_5352);
or U10438 (N_10438,N_9860,N_8164);
and U10439 (N_10439,N_6117,N_8349);
or U10440 (N_10440,N_9421,N_9710);
nand U10441 (N_10441,N_7827,N_9394);
nor U10442 (N_10442,N_7885,N_8366);
nand U10443 (N_10443,N_9576,N_8775);
nand U10444 (N_10444,N_9152,N_8322);
nor U10445 (N_10445,N_9890,N_5233);
or U10446 (N_10446,N_6012,N_7032);
nand U10447 (N_10447,N_6487,N_7431);
nand U10448 (N_10448,N_5390,N_9846);
nor U10449 (N_10449,N_5941,N_7468);
and U10450 (N_10450,N_7709,N_5240);
or U10451 (N_10451,N_8269,N_5709);
nand U10452 (N_10452,N_5678,N_9840);
and U10453 (N_10453,N_6703,N_6341);
nand U10454 (N_10454,N_9595,N_8494);
or U10455 (N_10455,N_6880,N_6787);
nor U10456 (N_10456,N_7853,N_6584);
and U10457 (N_10457,N_8350,N_7424);
xnor U10458 (N_10458,N_9313,N_9627);
or U10459 (N_10459,N_7888,N_9899);
and U10460 (N_10460,N_8052,N_6890);
xor U10461 (N_10461,N_8203,N_9944);
nor U10462 (N_10462,N_9544,N_5528);
and U10463 (N_10463,N_5407,N_6163);
nand U10464 (N_10464,N_6848,N_6054);
xnor U10465 (N_10465,N_7325,N_9510);
nor U10466 (N_10466,N_6999,N_8523);
nor U10467 (N_10467,N_8929,N_8601);
xnor U10468 (N_10468,N_5125,N_6778);
xnor U10469 (N_10469,N_9426,N_8508);
nor U10470 (N_10470,N_5047,N_9584);
or U10471 (N_10471,N_6058,N_5473);
nand U10472 (N_10472,N_9542,N_7182);
and U10473 (N_10473,N_6062,N_8973);
xnor U10474 (N_10474,N_9908,N_7215);
and U10475 (N_10475,N_8474,N_6422);
or U10476 (N_10476,N_9226,N_6139);
or U10477 (N_10477,N_6339,N_8576);
nor U10478 (N_10478,N_6798,N_8909);
and U10479 (N_10479,N_8503,N_5144);
xnor U10480 (N_10480,N_9793,N_5150);
nor U10481 (N_10481,N_5867,N_7470);
xnor U10482 (N_10482,N_8555,N_6359);
xor U10483 (N_10483,N_6153,N_8333);
or U10484 (N_10484,N_8109,N_5055);
xnor U10485 (N_10485,N_5597,N_8688);
nor U10486 (N_10486,N_5771,N_6282);
xnor U10487 (N_10487,N_6447,N_8323);
or U10488 (N_10488,N_8191,N_9514);
or U10489 (N_10489,N_9246,N_9465);
nor U10490 (N_10490,N_6653,N_7619);
xor U10491 (N_10491,N_5123,N_9200);
xnor U10492 (N_10492,N_6223,N_6129);
xor U10493 (N_10493,N_5818,N_9965);
and U10494 (N_10494,N_8328,N_7375);
xor U10495 (N_10495,N_8660,N_9493);
nand U10496 (N_10496,N_7368,N_8354);
xnor U10497 (N_10497,N_9596,N_6441);
nor U10498 (N_10498,N_8499,N_8902);
nand U10499 (N_10499,N_6693,N_8595);
nor U10500 (N_10500,N_5383,N_9391);
and U10501 (N_10501,N_7099,N_5067);
xor U10502 (N_10502,N_6806,N_5061);
nor U10503 (N_10503,N_7271,N_6911);
nand U10504 (N_10504,N_8608,N_9839);
xnor U10505 (N_10505,N_6678,N_5275);
xnor U10506 (N_10506,N_5148,N_7670);
nand U10507 (N_10507,N_8895,N_8806);
xor U10508 (N_10508,N_7402,N_5476);
nor U10509 (N_10509,N_7234,N_5835);
or U10510 (N_10510,N_6470,N_5780);
xnor U10511 (N_10511,N_9141,N_8609);
and U10512 (N_10512,N_8152,N_6421);
or U10513 (N_10513,N_9136,N_7680);
and U10514 (N_10514,N_9791,N_8850);
or U10515 (N_10515,N_9198,N_9859);
nand U10516 (N_10516,N_9309,N_6202);
nor U10517 (N_10517,N_7161,N_6953);
nand U10518 (N_10518,N_8736,N_7192);
and U10519 (N_10519,N_7344,N_9862);
nand U10520 (N_10520,N_9413,N_9236);
and U10521 (N_10521,N_8950,N_9238);
xor U10522 (N_10522,N_9815,N_7253);
nand U10523 (N_10523,N_7383,N_8728);
xor U10524 (N_10524,N_7693,N_8057);
nor U10525 (N_10525,N_9878,N_8626);
and U10526 (N_10526,N_7773,N_5594);
nand U10527 (N_10527,N_6825,N_8475);
and U10528 (N_10528,N_6723,N_6512);
nand U10529 (N_10529,N_6266,N_7096);
or U10530 (N_10530,N_6363,N_6369);
nand U10531 (N_10531,N_6304,N_8445);
or U10532 (N_10532,N_7659,N_7036);
and U10533 (N_10533,N_8722,N_8145);
nand U10534 (N_10534,N_6770,N_8921);
nand U10535 (N_10535,N_9095,N_8173);
nand U10536 (N_10536,N_9787,N_6278);
nor U10537 (N_10537,N_5698,N_8112);
nand U10538 (N_10538,N_6859,N_6069);
or U10539 (N_10539,N_6497,N_7008);
nor U10540 (N_10540,N_9800,N_7797);
xor U10541 (N_10541,N_5769,N_9507);
or U10542 (N_10542,N_5299,N_7242);
nand U10543 (N_10543,N_7846,N_7254);
xnor U10544 (N_10544,N_6060,N_9476);
xnor U10545 (N_10545,N_8748,N_8218);
nand U10546 (N_10546,N_7760,N_9408);
xor U10547 (N_10547,N_7133,N_9448);
nor U10548 (N_10548,N_8454,N_9827);
nand U10549 (N_10549,N_6273,N_7648);
nor U10550 (N_10550,N_6384,N_5631);
or U10551 (N_10551,N_5816,N_5645);
or U10552 (N_10552,N_5962,N_7471);
or U10553 (N_10553,N_8989,N_6526);
nor U10554 (N_10554,N_5995,N_6249);
and U10555 (N_10555,N_8092,N_5244);
xor U10556 (N_10556,N_7465,N_8081);
xor U10557 (N_10557,N_5464,N_5878);
or U10558 (N_10558,N_8448,N_6576);
or U10559 (N_10559,N_5392,N_8885);
xnor U10560 (N_10560,N_6736,N_8515);
and U10561 (N_10561,N_6797,N_8805);
and U10562 (N_10562,N_6668,N_8163);
or U10563 (N_10563,N_9639,N_9794);
and U10564 (N_10564,N_6882,N_8158);
xor U10565 (N_10565,N_8918,N_9739);
or U10566 (N_10566,N_6559,N_5520);
nor U10567 (N_10567,N_7997,N_9740);
or U10568 (N_10568,N_6573,N_5303);
nor U10569 (N_10569,N_8809,N_9254);
nand U10570 (N_10570,N_8358,N_5888);
or U10571 (N_10571,N_7996,N_9531);
xor U10572 (N_10572,N_9457,N_8625);
and U10573 (N_10573,N_6491,N_5362);
nor U10574 (N_10574,N_5111,N_6580);
xor U10575 (N_10575,N_6780,N_8180);
nand U10576 (N_10576,N_7389,N_6894);
xnor U10577 (N_10577,N_7859,N_8463);
nor U10578 (N_10578,N_6244,N_5784);
or U10579 (N_10579,N_5583,N_8889);
or U10580 (N_10580,N_9363,N_8693);
and U10581 (N_10581,N_6161,N_7076);
xor U10582 (N_10582,N_9816,N_5185);
nand U10583 (N_10583,N_8661,N_5653);
xor U10584 (N_10584,N_8281,N_5090);
xor U10585 (N_10585,N_7314,N_5007);
nor U10586 (N_10586,N_9521,N_7249);
and U10587 (N_10587,N_8955,N_8380);
or U10588 (N_10588,N_9266,N_5011);
and U10589 (N_10589,N_5756,N_7329);
or U10590 (N_10590,N_5530,N_9215);
xor U10591 (N_10591,N_9961,N_8063);
nor U10592 (N_10592,N_8439,N_5883);
and U10593 (N_10593,N_6428,N_5252);
nor U10594 (N_10594,N_8402,N_5051);
xnor U10595 (N_10595,N_6440,N_7523);
nor U10596 (N_10596,N_9057,N_9745);
xor U10597 (N_10597,N_9473,N_8689);
nor U10598 (N_10598,N_8923,N_6032);
or U10599 (N_10599,N_7994,N_8519);
nand U10600 (N_10600,N_8657,N_8335);
xor U10601 (N_10601,N_5615,N_6035);
nor U10602 (N_10602,N_7363,N_5312);
or U10603 (N_10603,N_6889,N_7322);
or U10604 (N_10604,N_5712,N_8564);
and U10605 (N_10605,N_5952,N_8373);
xnor U10606 (N_10606,N_7965,N_5012);
nand U10607 (N_10607,N_8301,N_9755);
nor U10608 (N_10608,N_9658,N_7457);
nand U10609 (N_10609,N_8936,N_6205);
or U10610 (N_10610,N_9626,N_9843);
nand U10611 (N_10611,N_6843,N_9321);
nand U10612 (N_10612,N_6969,N_6389);
and U10613 (N_10613,N_8591,N_8450);
nor U10614 (N_10614,N_7829,N_7426);
nand U10615 (N_10615,N_5483,N_8941);
nor U10616 (N_10616,N_7262,N_8592);
and U10617 (N_10617,N_5715,N_7833);
nor U10618 (N_10618,N_7397,N_8822);
xnor U10619 (N_10619,N_8796,N_8413);
xnor U10620 (N_10620,N_5608,N_5830);
nand U10621 (N_10621,N_9199,N_7263);
nand U10622 (N_10622,N_6427,N_5620);
xor U10623 (N_10623,N_7843,N_5710);
nand U10624 (N_10624,N_7738,N_9773);
or U10625 (N_10625,N_6241,N_7308);
nor U10626 (N_10626,N_5164,N_7920);
nand U10627 (N_10627,N_6961,N_5066);
xor U10628 (N_10628,N_5898,N_6933);
xor U10629 (N_10629,N_9059,N_5472);
or U10630 (N_10630,N_5396,N_7654);
or U10631 (N_10631,N_5582,N_6596);
and U10632 (N_10632,N_9397,N_6753);
or U10633 (N_10633,N_6442,N_6011);
xor U10634 (N_10634,N_8554,N_8896);
nand U10635 (N_10635,N_9738,N_5556);
nand U10636 (N_10636,N_8611,N_9241);
xnor U10637 (N_10637,N_9157,N_8853);
xnor U10638 (N_10638,N_9257,N_7238);
or U10639 (N_10639,N_5232,N_5287);
nor U10640 (N_10640,N_5927,N_5190);
nand U10641 (N_10641,N_9401,N_6935);
xnor U10642 (N_10642,N_9708,N_9684);
xor U10643 (N_10643,N_5280,N_7842);
nand U10644 (N_10644,N_8286,N_8093);
nor U10645 (N_10645,N_9979,N_9758);
and U10646 (N_10646,N_5247,N_8867);
or U10647 (N_10647,N_8339,N_6303);
nor U10648 (N_10648,N_8696,N_9657);
nand U10649 (N_10649,N_7726,N_7367);
nand U10650 (N_10650,N_9183,N_7992);
or U10651 (N_10651,N_7643,N_9079);
nand U10652 (N_10652,N_7449,N_8470);
and U10653 (N_10653,N_5536,N_5691);
xor U10654 (N_10654,N_9272,N_8529);
nor U10655 (N_10655,N_5541,N_6635);
xor U10656 (N_10656,N_8355,N_7712);
xnor U10657 (N_10657,N_9139,N_7629);
nor U10658 (N_10658,N_7201,N_6842);
nand U10659 (N_10659,N_8897,N_6238);
nor U10660 (N_10660,N_7226,N_8878);
nand U10661 (N_10661,N_5354,N_7777);
nand U10662 (N_10662,N_8325,N_7230);
and U10663 (N_10663,N_8667,N_5284);
nor U10664 (N_10664,N_8593,N_6688);
xor U10665 (N_10665,N_8014,N_8473);
nor U10666 (N_10666,N_5099,N_6645);
or U10667 (N_10667,N_6589,N_6621);
xor U10668 (N_10668,N_9328,N_6680);
nand U10669 (N_10669,N_8930,N_5974);
and U10670 (N_10670,N_5347,N_9468);
or U10671 (N_10671,N_7318,N_6017);
or U10672 (N_10672,N_7137,N_7472);
nor U10673 (N_10673,N_5986,N_8122);
and U10674 (N_10674,N_9697,N_8497);
xnor U10675 (N_10675,N_9904,N_5849);
or U10676 (N_10676,N_9995,N_6875);
xnor U10677 (N_10677,N_8845,N_8984);
nand U10678 (N_10678,N_5302,N_9900);
or U10679 (N_10679,N_9315,N_6963);
nand U10680 (N_10680,N_5149,N_5480);
nor U10681 (N_10681,N_8170,N_5961);
and U10682 (N_10682,N_7821,N_8623);
nor U10683 (N_10683,N_6550,N_7759);
nor U10684 (N_10684,N_9020,N_9092);
and U10685 (N_10685,N_5474,N_6721);
xnor U10686 (N_10686,N_7529,N_8540);
xnor U10687 (N_10687,N_9207,N_7730);
xor U10688 (N_10688,N_7101,N_5371);
xnor U10689 (N_10689,N_7690,N_8447);
nand U10690 (N_10690,N_6334,N_6622);
nor U10691 (N_10691,N_9025,N_8231);
xor U10692 (N_10692,N_9008,N_8101);
nor U10693 (N_10693,N_8343,N_6308);
xor U10694 (N_10694,N_8206,N_6997);
nor U10695 (N_10695,N_6790,N_7255);
xnor U10696 (N_10696,N_5417,N_6918);
xnor U10697 (N_10697,N_7388,N_9409);
or U10698 (N_10698,N_8861,N_7067);
xor U10699 (N_10699,N_6884,N_5097);
xnor U10700 (N_10700,N_5868,N_5122);
xnor U10701 (N_10701,N_6314,N_8680);
nand U10702 (N_10702,N_7461,N_7502);
or U10703 (N_10703,N_5191,N_7561);
or U10704 (N_10704,N_9817,N_9191);
or U10705 (N_10705,N_8517,N_7501);
xnor U10706 (N_10706,N_5807,N_7718);
nand U10707 (N_10707,N_5652,N_7906);
and U10708 (N_10708,N_7390,N_8928);
and U10709 (N_10709,N_8966,N_6871);
xnor U10710 (N_10710,N_9518,N_7027);
nand U10711 (N_10711,N_5776,N_9489);
or U10712 (N_10712,N_9349,N_7270);
or U10713 (N_10713,N_9530,N_6128);
nor U10714 (N_10714,N_6620,N_9225);
nor U10715 (N_10715,N_5866,N_7530);
xor U10716 (N_10716,N_6741,N_9122);
or U10717 (N_10717,N_7425,N_7051);
xnor U10718 (N_10718,N_8926,N_6415);
nor U10719 (N_10719,N_5655,N_9853);
or U10720 (N_10720,N_5005,N_5380);
and U10721 (N_10721,N_7765,N_7398);
xnor U10722 (N_10722,N_5570,N_9145);
and U10723 (N_10723,N_5262,N_9134);
xnor U10724 (N_10724,N_9167,N_7358);
and U10725 (N_10725,N_5084,N_8694);
nand U10726 (N_10726,N_6367,N_6877);
nor U10727 (N_10727,N_7636,N_6901);
nand U10728 (N_10728,N_5853,N_9712);
nor U10729 (N_10729,N_7645,N_5058);
or U10730 (N_10730,N_8111,N_6665);
or U10731 (N_10731,N_6137,N_8149);
and U10732 (N_10732,N_5861,N_7717);
nor U10733 (N_10733,N_7990,N_7858);
nor U10734 (N_10734,N_6126,N_6773);
and U10735 (N_10735,N_7552,N_8859);
or U10736 (N_10736,N_6016,N_6408);
or U10737 (N_10737,N_7590,N_9607);
xnor U10738 (N_10738,N_9400,N_6141);
and U10739 (N_10739,N_9306,N_6543);
or U10740 (N_10740,N_7860,N_6640);
or U10741 (N_10741,N_9077,N_9911);
xor U10742 (N_10742,N_5687,N_9278);
nor U10743 (N_10743,N_7435,N_5911);
and U10744 (N_10744,N_9999,N_7671);
xnor U10745 (N_10745,N_7919,N_7334);
or U10746 (N_10746,N_7960,N_7780);
nand U10747 (N_10747,N_7153,N_5529);
nor U10748 (N_10748,N_9366,N_7865);
and U10749 (N_10749,N_8792,N_5641);
or U10750 (N_10750,N_8318,N_5493);
or U10751 (N_10751,N_9178,N_7556);
nor U10752 (N_10752,N_6598,N_8182);
nand U10753 (N_10753,N_5165,N_5382);
nand U10754 (N_10754,N_7500,N_5259);
nand U10755 (N_10755,N_6104,N_7606);
and U10756 (N_10756,N_9830,N_5108);
xor U10757 (N_10757,N_6106,N_9512);
or U10758 (N_10758,N_6325,N_6910);
nor U10759 (N_10759,N_6522,N_8305);
nor U10760 (N_10760,N_7678,N_8708);
nand U10761 (N_10761,N_8193,N_5846);
nand U10762 (N_10762,N_6466,N_9456);
or U10763 (N_10763,N_7578,N_8275);
nor U10764 (N_10764,N_9194,N_9289);
or U10765 (N_10765,N_6727,N_6982);
nor U10766 (N_10766,N_8374,N_5258);
and U10767 (N_10767,N_6951,N_5624);
and U10768 (N_10768,N_5874,N_6283);
nand U10769 (N_10769,N_5800,N_5781);
xor U10770 (N_10770,N_6897,N_8598);
xnor U10771 (N_10771,N_6356,N_8372);
or U10772 (N_10772,N_8391,N_8901);
or U10773 (N_10773,N_5031,N_6398);
and U10774 (N_10774,N_7125,N_7532);
xor U10775 (N_10775,N_5218,N_9049);
xor U10776 (N_10776,N_5419,N_9833);
xnor U10777 (N_10777,N_9229,N_5923);
or U10778 (N_10778,N_8201,N_6854);
and U10779 (N_10779,N_9056,N_5204);
or U10780 (N_10780,N_6361,N_6575);
nor U10781 (N_10781,N_6994,N_5626);
and U10782 (N_10782,N_9419,N_5434);
nor U10783 (N_10783,N_6850,N_7026);
and U10784 (N_10784,N_6484,N_7217);
or U10785 (N_10785,N_9014,N_6548);
nand U10786 (N_10786,N_8451,N_9517);
nand U10787 (N_10787,N_6690,N_9326);
nor U10788 (N_10788,N_8455,N_7596);
and U10789 (N_10789,N_5175,N_9580);
xnor U10790 (N_10790,N_9293,N_9912);
and U10791 (N_10791,N_8428,N_6443);
nand U10792 (N_10792,N_8584,N_6506);
or U10793 (N_10793,N_6068,N_5216);
nor U10794 (N_10794,N_8395,N_7148);
nor U10795 (N_10795,N_9538,N_8243);
and U10796 (N_10796,N_6240,N_8534);
xor U10797 (N_10797,N_6038,N_7304);
nand U10798 (N_10798,N_7127,N_5817);
nor U10799 (N_10799,N_9451,N_8916);
or U10800 (N_10800,N_7555,N_9633);
nand U10801 (N_10801,N_6758,N_7819);
nor U10802 (N_10802,N_8162,N_5004);
nor U10803 (N_10803,N_9605,N_8118);
nand U10804 (N_10804,N_6800,N_7514);
nor U10805 (N_10805,N_5053,N_9174);
and U10806 (N_10806,N_7976,N_9825);
or U10807 (N_10807,N_8839,N_6027);
nor U10808 (N_10808,N_7451,N_5663);
or U10809 (N_10809,N_8500,N_8804);
xor U10810 (N_10810,N_6760,N_6781);
or U10811 (N_10811,N_9805,N_5348);
or U10812 (N_10812,N_7711,N_8810);
and U10813 (N_10813,N_7901,N_8085);
and U10814 (N_10814,N_7442,N_7086);
nand U10815 (N_10815,N_7068,N_8860);
xnor U10816 (N_10816,N_6525,N_7024);
nor U10817 (N_10817,N_5277,N_8714);
or U10818 (N_10818,N_7679,N_6534);
or U10819 (N_10819,N_9082,N_6679);
and U10820 (N_10820,N_9730,N_8730);
nand U10821 (N_10821,N_6785,N_6186);
nor U10822 (N_10822,N_5427,N_8412);
or U10823 (N_10823,N_6193,N_9041);
nor U10824 (N_10824,N_7126,N_7975);
or U10825 (N_10825,N_6836,N_5353);
nand U10826 (N_10826,N_5880,N_5760);
nand U10827 (N_10827,N_6764,N_8277);
and U10828 (N_10828,N_7244,N_7003);
xnor U10829 (N_10829,N_8665,N_9579);
or U10830 (N_10830,N_8233,N_5402);
or U10831 (N_10831,N_7039,N_5393);
or U10832 (N_10832,N_9147,N_6459);
nor U10833 (N_10833,N_5981,N_6542);
xor U10834 (N_10834,N_6210,N_7650);
xnor U10835 (N_10835,N_9378,N_8492);
nand U10836 (N_10836,N_6876,N_6040);
nor U10837 (N_10837,N_8716,N_6383);
xor U10838 (N_10838,N_9909,N_7319);
or U10839 (N_10839,N_5586,N_7293);
nor U10840 (N_10840,N_5285,N_9933);
or U10841 (N_10841,N_9170,N_5222);
or U10842 (N_10842,N_7278,N_8932);
nand U10843 (N_10843,N_6909,N_8313);
xnor U10844 (N_10844,N_7045,N_6111);
xnor U10845 (N_10845,N_9925,N_5991);
or U10846 (N_10846,N_6569,N_8749);
nor U10847 (N_10847,N_8710,N_5394);
xnor U10848 (N_10848,N_6405,N_9903);
or U10849 (N_10849,N_5773,N_9551);
or U10850 (N_10850,N_7204,N_7160);
or U10851 (N_10851,N_6477,N_8686);
nor U10852 (N_10852,N_8504,N_6514);
and U10853 (N_10853,N_8230,N_7295);
nand U10854 (N_10854,N_5877,N_7715);
and U10855 (N_10855,N_8443,N_7347);
xor U10856 (N_10856,N_8252,N_8521);
xor U10857 (N_10857,N_7144,N_6208);
nor U10858 (N_10858,N_6756,N_6015);
xnor U10859 (N_10859,N_5339,N_9695);
or U10860 (N_10860,N_6410,N_7725);
nand U10861 (N_10861,N_5929,N_8553);
nand U10862 (N_10862,N_9574,N_5696);
xnor U10863 (N_10863,N_7233,N_8606);
nor U10864 (N_10864,N_9417,N_8257);
xnor U10865 (N_10865,N_9406,N_7830);
xnor U10866 (N_10866,N_9460,N_9775);
or U10867 (N_10867,N_6426,N_5968);
nand U10868 (N_10868,N_5761,N_9483);
nand U10869 (N_10869,N_9804,N_9989);
nand U10870 (N_10870,N_8169,N_7736);
and U10871 (N_10871,N_6370,N_9670);
and U10872 (N_10872,N_9714,N_8186);
nand U10873 (N_10873,N_5033,N_9469);
and U10874 (N_10874,N_6647,N_6013);
nand U10875 (N_10875,N_8253,N_7496);
and U10876 (N_10876,N_9265,N_7410);
nand U10877 (N_10877,N_7907,N_9784);
and U10878 (N_10878,N_6499,N_8051);
nor U10879 (N_10879,N_8785,N_8009);
nand U10880 (N_10880,N_8142,N_8552);
xnor U10881 (N_10881,N_6323,N_9983);
and U10882 (N_10882,N_5433,N_5015);
xor U10883 (N_10883,N_9385,N_6980);
nor U10884 (N_10884,N_6063,N_8292);
nand U10885 (N_10885,N_7223,N_5042);
nor U10886 (N_10886,N_9303,N_6662);
and U10887 (N_10887,N_8123,N_5831);
nand U10888 (N_10888,N_7512,N_7222);
nand U10889 (N_10889,N_9905,N_6215);
or U10890 (N_10890,N_6811,N_6092);
and U10891 (N_10891,N_8021,N_8442);
nor U10892 (N_10892,N_6822,N_5411);
and U10893 (N_10893,N_5978,N_7557);
xor U10894 (N_10894,N_7605,N_8546);
or U10895 (N_10895,N_8319,N_6034);
xor U10896 (N_10896,N_8631,N_8615);
or U10897 (N_10897,N_6090,N_8167);
nor U10898 (N_10898,N_6148,N_8802);
xor U10899 (N_10899,N_6972,N_8471);
or U10900 (N_10900,N_5046,N_9335);
nor U10901 (N_10901,N_8747,N_9865);
xnor U10902 (N_10902,N_5890,N_7941);
and U10903 (N_10903,N_5956,N_7245);
xnor U10904 (N_10904,N_8062,N_5820);
and U10905 (N_10905,N_5872,N_5387);
xor U10906 (N_10906,N_5350,N_5391);
nor U10907 (N_10907,N_9523,N_7511);
nor U10908 (N_10908,N_5071,N_9052);
and U10909 (N_10909,N_5263,N_6366);
xnor U10910 (N_10910,N_6634,N_7653);
nor U10911 (N_10911,N_9838,N_5505);
nor U10912 (N_10912,N_6176,N_5600);
nand U10913 (N_10913,N_7042,N_8764);
and U10914 (N_10914,N_6539,N_8261);
xnor U10915 (N_10915,N_7762,N_5627);
or U10916 (N_10916,N_5704,N_7059);
or U10917 (N_10917,N_6891,N_9271);
and U10918 (N_10918,N_6116,N_9148);
or U10919 (N_10919,N_9031,N_7029);
and U10920 (N_10920,N_5162,N_7335);
or U10921 (N_10921,N_9017,N_7048);
xor U10922 (N_10922,N_5332,N_9011);
xnor U10923 (N_10923,N_5733,N_7571);
and U10924 (N_10924,N_7216,N_6538);
xor U10925 (N_10925,N_5885,N_6347);
nor U10926 (N_10926,N_9637,N_5468);
and U10927 (N_10927,N_9171,N_7849);
nand U10928 (N_10928,N_9617,N_9620);
xnor U10929 (N_10929,N_8137,N_7958);
nor U10930 (N_10930,N_9377,N_7899);
nand U10931 (N_10931,N_9425,N_5717);
nand U10932 (N_10932,N_8724,N_6810);
or U10933 (N_10933,N_7681,N_8633);
xnor U10934 (N_10934,N_9640,N_7418);
and U10935 (N_10935,N_6234,N_7741);
nand U10936 (N_10936,N_7213,N_5436);
and U10937 (N_10937,N_8096,N_5174);
or U10938 (N_10938,N_6500,N_7840);
nor U10939 (N_10939,N_9883,N_7483);
nand U10940 (N_10940,N_8703,N_8157);
nand U10941 (N_10941,N_8044,N_8707);
and U10942 (N_10942,N_8489,N_6046);
and U10943 (N_10943,N_5081,N_9674);
and U10944 (N_10944,N_9947,N_6630);
and U10945 (N_10945,N_8761,N_6118);
or U10946 (N_10946,N_8017,N_5095);
xnor U10947 (N_10947,N_7422,N_6373);
or U10948 (N_10948,N_5269,N_8429);
and U10949 (N_10949,N_6537,N_9874);
nand U10950 (N_10950,N_7649,N_6134);
nor U10951 (N_10951,N_6674,N_6042);
and U10952 (N_10952,N_7309,N_7687);
and U10953 (N_10953,N_6119,N_6140);
xor U10954 (N_10954,N_7674,N_7102);
nand U10955 (N_10955,N_6831,N_7129);
nor U10956 (N_10956,N_9010,N_6551);
and U10957 (N_10957,N_9428,N_7071);
nor U10958 (N_10958,N_6618,N_7275);
nor U10959 (N_10959,N_6311,N_8586);
or U10960 (N_10960,N_5599,N_8421);
or U10961 (N_10961,N_8963,N_8556);
or U10962 (N_10962,N_5658,N_6430);
and U10963 (N_10963,N_6623,N_6561);
xor U10964 (N_10964,N_5542,N_5121);
xnor U10965 (N_10965,N_5134,N_6476);
and U10966 (N_10966,N_6698,N_6588);
nand U10967 (N_10967,N_7060,N_7826);
and U10968 (N_10968,N_9322,N_6420);
nand U10969 (N_10969,N_6452,N_7825);
and U10970 (N_10970,N_6277,N_6914);
and U10971 (N_10971,N_7141,N_5328);
and U10972 (N_10972,N_6374,N_8388);
nand U10973 (N_10973,N_6082,N_6612);
and U10974 (N_10974,N_7630,N_7447);
nand U10975 (N_10975,N_8417,N_7439);
nor U10976 (N_10976,N_8039,N_8975);
nand U10977 (N_10977,N_5924,N_6127);
nor U10978 (N_10978,N_9832,N_7927);
or U10979 (N_10979,N_9948,N_5636);
nand U10980 (N_10980,N_8362,N_6482);
or U10981 (N_10981,N_5124,N_8908);
nor U10982 (N_10982,N_8254,N_5671);
and U10983 (N_10983,N_7847,N_8880);
and U10984 (N_10984,N_9075,N_6114);
or U10985 (N_10985,N_9680,N_7400);
nand U10986 (N_10986,N_8020,N_8852);
nand U10987 (N_10987,N_8035,N_6437);
nand U10988 (N_10988,N_6744,N_8403);
and U10989 (N_10989,N_6602,N_6110);
or U10990 (N_10990,N_8345,N_8524);
xnor U10991 (N_10991,N_9243,N_9138);
or U10992 (N_10992,N_7106,N_7978);
xnor U10993 (N_10993,N_9611,N_7893);
or U10994 (N_10994,N_7747,N_7647);
nand U10995 (N_10995,N_8210,N_8655);
or U10996 (N_10996,N_5585,N_6817);
nor U10997 (N_10997,N_8829,N_8531);
xor U10998 (N_10998,N_6837,N_8394);
or U10999 (N_10999,N_8385,N_7258);
nor U11000 (N_11000,N_7174,N_5666);
nor U11001 (N_11001,N_9648,N_7525);
nand U11002 (N_11002,N_9018,N_8064);
and U11003 (N_11003,N_7421,N_7999);
or U11004 (N_11004,N_8574,N_9371);
xor U11005 (N_11005,N_7535,N_6949);
and U11006 (N_11006,N_7946,N_5039);
or U11007 (N_11007,N_7291,N_8461);
nand U11008 (N_11008,N_8965,N_6767);
nand U11009 (N_11009,N_9376,N_8871);
and U11010 (N_11010,N_5841,N_7962);
nor U11011 (N_11011,N_9277,N_9622);
nor U11012 (N_11012,N_6527,N_7001);
or U11013 (N_11013,N_8701,N_8054);
or U11014 (N_11014,N_7474,N_9233);
nand U11015 (N_11015,N_5368,N_6350);
xor U11016 (N_11016,N_8468,N_7366);
and U11017 (N_11017,N_8430,N_5737);
or U11018 (N_11018,N_7385,N_5591);
and U11019 (N_11019,N_9656,N_6319);
nor U11020 (N_11020,N_9392,N_6180);
or U11021 (N_11021,N_9201,N_6246);
xnor U11022 (N_11022,N_8361,N_9193);
or U11023 (N_11023,N_8573,N_5565);
nor U11024 (N_11024,N_8639,N_8189);
nand U11025 (N_11025,N_8969,N_9009);
xor U11026 (N_11026,N_8847,N_7432);
and U11027 (N_11027,N_9029,N_8426);
nand U11028 (N_11028,N_8788,N_9849);
nor U11029 (N_11029,N_6489,N_5719);
nor U11030 (N_11030,N_6783,N_6261);
and U11031 (N_11031,N_5948,N_8026);
xnor U11032 (N_11032,N_8888,N_9725);
nor U11033 (N_11033,N_8682,N_8053);
nand U11034 (N_11034,N_7550,N_8205);
nand U11035 (N_11035,N_5320,N_9123);
nor U11036 (N_11036,N_9655,N_7266);
nand U11037 (N_11037,N_8619,N_9250);
or U11038 (N_11038,N_5754,N_8590);
xnor U11039 (N_11039,N_7769,N_7105);
nand U11040 (N_11040,N_7055,N_7537);
nor U11041 (N_11041,N_8883,N_7939);
nor U11042 (N_11042,N_7220,N_8208);
or U11043 (N_11043,N_9154,N_6766);
nor U11044 (N_11044,N_7159,N_6986);
nand U11045 (N_11045,N_7218,N_7228);
xor U11046 (N_11046,N_5943,N_6307);
nor U11047 (N_11047,N_9573,N_9572);
nand U11048 (N_11048,N_6077,N_7093);
xnor U11049 (N_11049,N_9150,N_8177);
nand U11050 (N_11050,N_9519,N_9205);
nor U11051 (N_11051,N_5907,N_9673);
nand U11052 (N_11052,N_7527,N_6254);
nor U11053 (N_11053,N_8479,N_7661);
or U11054 (N_11054,N_7114,N_8198);
nand U11055 (N_11055,N_9719,N_7531);
and U11056 (N_11056,N_8866,N_6964);
nand U11057 (N_11057,N_6651,N_9480);
nor U11058 (N_11058,N_9779,N_9107);
or U11059 (N_11059,N_6908,N_8266);
or U11060 (N_11060,N_9252,N_8925);
nand U11061 (N_11061,N_8297,N_8127);
nor U11062 (N_11062,N_7823,N_5925);
nor U11063 (N_11063,N_7300,N_7030);
and U11064 (N_11064,N_7303,N_6819);
xor U11065 (N_11065,N_5690,N_7337);
and U11066 (N_11066,N_6816,N_9902);
nor U11067 (N_11067,N_9525,N_8507);
nor U11068 (N_11068,N_7959,N_5500);
and U11069 (N_11069,N_5893,N_6714);
nor U11070 (N_11070,N_9789,N_6135);
nor U11071 (N_11071,N_6617,N_9430);
nand U11072 (N_11072,N_7507,N_6676);
and U11073 (N_11073,N_8838,N_5990);
nor U11074 (N_11074,N_9269,N_5160);
nand U11075 (N_11075,N_5806,N_7136);
nor U11076 (N_11076,N_8637,N_5171);
nand U11077 (N_11077,N_9771,N_6088);
or U11078 (N_11078,N_7130,N_7639);
xnor U11079 (N_11079,N_9629,N_6098);
nor U11080 (N_11080,N_9892,N_5928);
xor U11081 (N_11081,N_5469,N_9806);
xnor U11082 (N_11082,N_9689,N_5265);
nand U11083 (N_11083,N_8095,N_7884);
nor U11084 (N_11084,N_8067,N_8549);
or U11085 (N_11085,N_8216,N_5088);
nor U11086 (N_11086,N_6481,N_5708);
xnor U11087 (N_11087,N_5581,N_7766);
and U11088 (N_11088,N_6917,N_9694);
and U11089 (N_11089,N_9073,N_8097);
or U11090 (N_11090,N_8887,N_5602);
nor U11091 (N_11091,N_5270,N_6313);
nand U11092 (N_11092,N_7915,N_7034);
and U11093 (N_11093,N_5751,N_5510);
nor U11094 (N_11094,N_7430,N_9502);
and U11095 (N_11095,N_5418,N_5410);
nand U11096 (N_11096,N_8436,N_9990);
or U11097 (N_11097,N_7822,N_8340);
or U11098 (N_11098,N_7301,N_5009);
or U11099 (N_11099,N_8416,N_6751);
or U11100 (N_11100,N_9606,N_5462);
nand U11101 (N_11101,N_6943,N_7269);
and U11102 (N_11102,N_8482,N_7553);
nor U11103 (N_11103,N_6862,N_7898);
nand U11104 (N_11104,N_5546,N_9120);
nor U11105 (N_11105,N_8964,N_6067);
nand U11106 (N_11106,N_5532,N_5129);
nor U11107 (N_11107,N_9382,N_7250);
nor U11108 (N_11108,N_6631,N_5840);
xnor U11109 (N_11109,N_8196,N_8383);
and U11110 (N_11110,N_9628,N_5141);
and U11111 (N_11111,N_7793,N_9951);
or U11112 (N_11112,N_6414,N_6531);
nand U11113 (N_11113,N_5378,N_9782);
or U11114 (N_11114,N_5913,N_8913);
xnor U11115 (N_11115,N_8869,N_7276);
nand U11116 (N_11116,N_7694,N_6079);
and U11117 (N_11117,N_7012,N_8765);
nand U11118 (N_11118,N_8419,N_7427);
xor U11119 (N_11119,N_6085,N_8807);
nand U11120 (N_11120,N_6847,N_9255);
xnor U11121 (N_11121,N_9885,N_7544);
or U11122 (N_11122,N_8891,N_5648);
xnor U11123 (N_11123,N_8221,N_9422);
and U11124 (N_11124,N_8229,N_9781);
nand U11125 (N_11125,N_6929,N_6434);
or U11126 (N_11126,N_6998,N_7641);
xnor U11127 (N_11127,N_9558,N_7073);
or U11128 (N_11128,N_5596,N_8223);
and U11129 (N_11129,N_8458,N_5182);
xor U11130 (N_11130,N_5589,N_8882);
or U11131 (N_11131,N_5030,N_5606);
nand U11132 (N_11132,N_5137,N_6458);
and U11133 (N_11133,N_6445,N_8786);
nand U11134 (N_11134,N_6177,N_5613);
and U11135 (N_11135,N_8185,N_7565);
xor U11136 (N_11136,N_6707,N_9537);
xor U11137 (N_11137,N_6100,N_5588);
nor U11138 (N_11138,N_8214,N_5891);
xnor U11139 (N_11139,N_9155,N_9724);
or U11140 (N_11140,N_6289,N_7889);
xor U11141 (N_11141,N_5130,N_5579);
xor U11142 (N_11142,N_9963,N_8971);
xnor U11143 (N_11143,N_5745,N_9054);
or U11144 (N_11144,N_7019,N_5454);
nand U11145 (N_11145,N_9346,N_5194);
nand U11146 (N_11146,N_9188,N_9046);
or U11147 (N_11147,N_9750,N_8649);
or U11148 (N_11148,N_7870,N_5248);
nor U11149 (N_11149,N_9819,N_9169);
nor U11150 (N_11150,N_5300,N_8245);
and U11151 (N_11151,N_7848,N_9923);
or U11152 (N_11152,N_9012,N_7837);
nand U11153 (N_11153,N_7869,N_8600);
nor U11154 (N_11154,N_8533,N_6706);
nor U11155 (N_11155,N_5250,N_9380);
and U11156 (N_11156,N_7371,N_5525);
nand U11157 (N_11157,N_5908,N_5173);
and U11158 (N_11158,N_9654,N_7288);
or U11159 (N_11159,N_7231,N_5192);
and U11160 (N_11160,N_9826,N_5485);
xor U11161 (N_11161,N_5274,N_8326);
nand U11162 (N_11162,N_6232,N_6952);
or U11163 (N_11163,N_9039,N_9516);
nor U11164 (N_11164,N_5775,N_6830);
nor U11165 (N_11165,N_5860,N_6856);
nand U11166 (N_11166,N_6052,N_7166);
nand U11167 (N_11167,N_6779,N_6224);
xor U11168 (N_11168,N_7115,N_7481);
xor U11169 (N_11169,N_5707,N_9067);
or U11170 (N_11170,N_9260,N_5210);
nor U11171 (N_11171,N_7633,N_7564);
nand U11172 (N_11172,N_9880,N_9085);
nand U11173 (N_11173,N_9256,N_8993);
xor U11174 (N_11174,N_5372,N_6956);
xnor U11175 (N_11175,N_6144,N_7977);
or U11176 (N_11176,N_9752,N_7044);
xnor U11177 (N_11177,N_7723,N_6503);
nor U11178 (N_11178,N_6030,N_7445);
nor U11179 (N_11179,N_9550,N_7942);
nor U11180 (N_11180,N_9432,N_7180);
xor U11181 (N_11181,N_6478,N_9796);
and U11182 (N_11182,N_8763,N_9702);
nor U11183 (N_11183,N_8617,N_6863);
or U11184 (N_11184,N_6839,N_6174);
and U11185 (N_11185,N_7408,N_9117);
nor U11186 (N_11186,N_8353,N_8249);
nor U11187 (N_11187,N_9506,N_6188);
xor U11188 (N_11188,N_8446,N_8375);
xor U11189 (N_11189,N_7622,N_9986);
or U11190 (N_11190,N_7415,N_9910);
and U11191 (N_11191,N_9373,N_5862);
nand U11192 (N_11192,N_8338,N_7151);
and U11193 (N_11193,N_9884,N_7404);
or U11194 (N_11194,N_6606,N_8232);
xnor U11195 (N_11195,N_7065,N_6763);
or U11196 (N_11196,N_8146,N_5743);
or U11197 (N_11197,N_8087,N_5450);
or U11198 (N_11198,N_8958,N_6560);
nand U11199 (N_11199,N_7509,N_5324);
nor U11200 (N_11200,N_9093,N_6547);
nand U11201 (N_11201,N_9124,N_9375);
nand U11202 (N_11202,N_5076,N_5018);
nor U11203 (N_11203,N_7804,N_8687);
and U11204 (N_11204,N_6954,N_9021);
and U11205 (N_11205,N_5399,N_8139);
or U11206 (N_11206,N_7485,N_5288);
nor U11207 (N_11207,N_7000,N_8962);
or U11208 (N_11208,N_5759,N_8833);
xor U11209 (N_11209,N_6968,N_5344);
nand U11210 (N_11210,N_8740,N_9778);
xor U11211 (N_11211,N_8228,N_8289);
nand U11212 (N_11212,N_7113,N_5984);
nand U11213 (N_11213,N_8957,N_9223);
xor U11214 (N_11214,N_9240,N_6603);
xnor U11215 (N_11215,N_5471,N_5060);
xnor U11216 (N_11216,N_9754,N_6485);
xor U11217 (N_11217,N_9444,N_5439);
nand U11218 (N_11218,N_8924,N_9268);
nand U11219 (N_11219,N_8437,N_7948);
and U11220 (N_11220,N_9568,N_9458);
and U11221 (N_11221,N_8239,N_9159);
and U11222 (N_11222,N_6072,N_6990);
or U11223 (N_11223,N_5342,N_7735);
and U11224 (N_11224,N_8018,N_7328);
or U11225 (N_11225,N_9219,N_6985);
nand U11226 (N_11226,N_8780,N_5931);
or U11227 (N_11227,N_7618,N_5227);
xnor U11228 (N_11228,N_6834,N_8638);
and U11229 (N_11229,N_7046,N_9631);
nand U11230 (N_11230,N_7510,N_9632);
nand U11231 (N_11231,N_6591,N_9389);
or U11232 (N_11232,N_8036,N_7243);
xnor U11233 (N_11233,N_6625,N_6352);
xnor U11234 (N_11234,N_5523,N_6905);
xnor U11235 (N_11235,N_8835,N_9756);
nand U11236 (N_11236,N_6065,N_7446);
nand U11237 (N_11237,N_8263,N_8825);
nand U11238 (N_11238,N_9635,N_9044);
xnor U11239 (N_11239,N_8150,N_7877);
nor U11240 (N_11240,N_6654,N_9560);
or U11241 (N_11241,N_6613,N_7251);
or U11242 (N_11242,N_6300,N_9809);
and U11243 (N_11243,N_8268,N_8662);
nor U11244 (N_11244,N_6808,N_6849);
nor U11245 (N_11245,N_8820,N_9696);
nor U11246 (N_11246,N_7614,N_5309);
nand U11247 (N_11247,N_5801,N_5494);
xor U11248 (N_11248,N_7700,N_6209);
and U11249 (N_11249,N_8108,N_5140);
nor U11250 (N_11250,N_9946,N_7952);
nand U11251 (N_11251,N_9915,N_9103);
nand U11252 (N_11252,N_5538,N_6078);
xor U11253 (N_11253,N_9901,N_5446);
nor U11254 (N_11254,N_8522,N_5895);
or U11255 (N_11255,N_8422,N_8700);
and U11256 (N_11256,N_5049,N_6051);
and U11257 (N_11257,N_6269,N_9264);
nor U11258 (N_11258,N_9613,N_9612);
nor U11259 (N_11259,N_7955,N_5647);
nand U11260 (N_11260,N_9355,N_7814);
or U11261 (N_11261,N_6689,N_6987);
and U11262 (N_11262,N_7428,N_8959);
nor U11263 (N_11263,N_5879,N_6896);
nand U11264 (N_11264,N_9660,N_5980);
xnor U11265 (N_11265,N_7090,N_5331);
or U11266 (N_11266,N_7542,N_7956);
or U11267 (N_11267,N_9005,N_8726);
xor U11268 (N_11268,N_6558,N_7007);
or U11269 (N_11269,N_8005,N_9760);
or U11270 (N_11270,N_6607,N_5424);
xnor U11271 (N_11271,N_8016,N_6175);
xor U11272 (N_11272,N_8675,N_5207);
or U11273 (N_11273,N_7728,N_5370);
xnor U11274 (N_11274,N_7184,N_8284);
xor U11275 (N_11275,N_7200,N_9365);
xnor U11276 (N_11276,N_5901,N_9455);
and U11277 (N_11277,N_5481,N_6024);
and U11278 (N_11278,N_5595,N_8049);
nand U11279 (N_11279,N_5023,N_9524);
or U11280 (N_11280,N_7412,N_7841);
or U11281 (N_11281,N_8983,N_5988);
nand U11282 (N_11282,N_5008,N_6624);
nor U11283 (N_11283,N_5180,N_7454);
and U11284 (N_11284,N_6436,N_6720);
xor U11285 (N_11285,N_8390,N_8032);
or U11286 (N_11286,N_9960,N_9644);
nor U11287 (N_11287,N_6587,N_7310);
nand U11288 (N_11288,N_9940,N_6005);
and U11289 (N_11289,N_9360,N_6776);
nor U11290 (N_11290,N_7411,N_9491);
or U11291 (N_11291,N_8410,N_7928);
or U11292 (N_11292,N_7910,N_6498);
or U11293 (N_11293,N_7731,N_7714);
or U11294 (N_11294,N_9210,N_9672);
nor U11295 (N_11295,N_9685,N_7974);
nand U11296 (N_11296,N_6792,N_8119);
and U11297 (N_11297,N_9601,N_7638);
nor U11298 (N_11298,N_9564,N_6517);
or U11299 (N_11299,N_8120,N_6360);
and U11300 (N_11300,N_5514,N_5460);
and U11301 (N_11301,N_9453,N_8745);
nor U11302 (N_11302,N_5503,N_9112);
or U11303 (N_11303,N_9666,N_8219);
xor U11304 (N_11304,N_9582,N_7722);
xnor U11305 (N_11305,N_9855,N_5404);
xor U11306 (N_11306,N_7098,N_7313);
and U11307 (N_11307,N_6915,N_9973);
nand U11308 (N_11308,N_6151,N_9175);
xor U11309 (N_11309,N_5533,N_6302);
xnor U11310 (N_11310,N_7124,N_7103);
and U11311 (N_11311,N_8920,N_9786);
xnor U11312 (N_11312,N_8542,N_8992);
and U11313 (N_11313,N_8321,N_8927);
nand U11314 (N_11314,N_7111,N_7603);
nor U11315 (N_11315,N_9913,N_9790);
nand U11316 (N_11316,N_9643,N_7664);
xor U11317 (N_11317,N_9262,N_7631);
and U11318 (N_11318,N_9353,N_5063);
xnor U11319 (N_11319,N_7601,N_9395);
or U11320 (N_11320,N_6515,N_8324);
and U11321 (N_11321,N_7237,N_9450);
nor U11322 (N_11322,N_6974,N_6739);
nand U11323 (N_11323,N_9661,N_9345);
nor U11324 (N_11324,N_5515,N_8683);
or U11325 (N_11325,N_6649,N_6003);
and U11326 (N_11326,N_7720,N_6267);
or U11327 (N_11327,N_7855,N_9917);
nor U11328 (N_11328,N_8794,N_6883);
or U11329 (N_11329,N_7256,N_8389);
and U11330 (N_11330,N_7866,N_5085);
or U11331 (N_11331,N_8400,N_5953);
xnor U11332 (N_11332,N_8972,N_9570);
or U11333 (N_11333,N_5413,N_6795);
xor U11334 (N_11334,N_9383,N_6023);
and U11335 (N_11335,N_7156,N_5838);
nor U11336 (N_11336,N_5802,N_8104);
or U11337 (N_11337,N_9501,N_6194);
and U11338 (N_11338,N_7326,N_5767);
nand U11339 (N_11339,N_6906,N_5443);
nand U11340 (N_11340,N_5742,N_9481);
xnor U11341 (N_11341,N_8622,N_5271);
or U11342 (N_11342,N_6152,N_5307);
and U11343 (N_11343,N_6562,N_6494);
nand U11344 (N_11344,N_8991,N_7149);
xnor U11345 (N_11345,N_6386,N_8154);
nand U11346 (N_11346,N_8212,N_6637);
and U11347 (N_11347,N_9013,N_8100);
nand U11348 (N_11348,N_6730,N_6195);
or U11349 (N_11349,N_5578,N_7091);
nand U11350 (N_11350,N_5694,N_6784);
or U11351 (N_11351,N_5699,N_5634);
nand U11352 (N_11352,N_6619,N_9047);
xnor U11353 (N_11353,N_5077,N_5987);
and U11354 (N_11354,N_7221,N_6089);
xnor U11355 (N_11355,N_7041,N_7539);
and U11356 (N_11356,N_9216,N_5449);
xnor U11357 (N_11357,N_7343,N_5145);
xor U11358 (N_11358,N_9153,N_9368);
nor U11359 (N_11359,N_7929,N_5422);
and U11360 (N_11360,N_9224,N_9114);
xnor U11361 (N_11361,N_7399,N_8408);
nand U11362 (N_11362,N_6349,N_6146);
nand U11363 (N_11363,N_8045,N_9618);
and U11364 (N_11364,N_7534,N_8113);
nand U11365 (N_11365,N_9386,N_6938);
xor U11366 (N_11366,N_9985,N_5812);
or U11367 (N_11367,N_6782,N_8414);
xor U11368 (N_11368,N_9498,N_9937);
or U11369 (N_11369,N_9324,N_8188);
nor U11370 (N_11370,N_6201,N_5118);
nand U11371 (N_11371,N_6203,N_7627);
nor U11372 (N_11372,N_6236,N_7311);
nand U11373 (N_11373,N_8260,N_7211);
nand U11374 (N_11374,N_8486,N_8870);
or U11375 (N_11375,N_9467,N_7224);
nor U11376 (N_11376,N_7064,N_9381);
nor U11377 (N_11377,N_9587,N_8945);
and U11378 (N_11378,N_5549,N_7128);
nor U11379 (N_11379,N_7494,N_7548);
nor U11380 (N_11380,N_8378,N_8425);
or U11381 (N_11381,N_8900,N_6355);
nor U11382 (N_11382,N_5850,N_6022);
nand U11383 (N_11383,N_6488,N_6578);
nand U11384 (N_11384,N_5479,N_8501);
or U11385 (N_11385,N_8251,N_7536);
nor U11386 (N_11386,N_8194,N_6708);
nand U11387 (N_11387,N_6115,N_9332);
nor U11388 (N_11388,N_7802,N_9024);
nand U11389 (N_11389,N_8940,N_8099);
or U11390 (N_11390,N_6301,N_5768);
xnor U11391 (N_11391,N_7279,N_8502);
and U11392 (N_11392,N_7441,N_5711);
nand U11393 (N_11393,N_5261,N_7864);
nor U11394 (N_11394,N_6976,N_5184);
nand U11395 (N_11395,N_6840,N_5249);
and U11396 (N_11396,N_6290,N_6672);
and U11397 (N_11397,N_9630,N_6796);
nand U11398 (N_11398,N_7336,N_5881);
and U11399 (N_11399,N_5966,N_5106);
or U11400 (N_11400,N_7513,N_5279);
xor U11401 (N_11401,N_5491,N_6735);
or U11402 (N_11402,N_8509,N_6860);
or U11403 (N_11403,N_9509,N_8264);
nor U11404 (N_11404,N_8893,N_5813);
xnor U11405 (N_11405,N_7181,N_9096);
or U11406 (N_11406,N_7171,N_6212);
nand U11407 (N_11407,N_6406,N_6509);
or U11408 (N_11408,N_5593,N_6157);
nand U11409 (N_11409,N_5003,N_5409);
xnor U11410 (N_11410,N_8558,N_8041);
nor U11411 (N_11411,N_6404,N_8215);
xor U11412 (N_11412,N_8059,N_9137);
and U11413 (N_11413,N_6799,N_5700);
nor U11414 (N_11414,N_6310,N_5166);
nand U11415 (N_11415,N_6317,N_7354);
xor U11416 (N_11416,N_7345,N_7261);
nor U11417 (N_11417,N_8510,N_6167);
nand U11418 (N_11418,N_7925,N_7570);
or U11419 (N_11419,N_7986,N_6669);
nand U11420 (N_11420,N_6505,N_6869);
nand U11421 (N_11421,N_8587,N_5363);
and U11422 (N_11422,N_7214,N_8525);
nor U11423 (N_11423,N_9333,N_9416);
and U11424 (N_11424,N_9358,N_9930);
and U11425 (N_11425,N_7594,N_7807);
or U11426 (N_11426,N_9705,N_7863);
nor U11427 (N_11427,N_9731,N_8476);
xor U11428 (N_11428,N_5092,N_8176);
nor U11429 (N_11429,N_9173,N_9312);
nand U11430 (N_11430,N_6231,N_8308);
nand U11431 (N_11431,N_6247,N_9006);
and U11432 (N_11432,N_5305,N_8466);
nor U11433 (N_11433,N_9975,N_6087);
or U11434 (N_11434,N_9036,N_6378);
and U11435 (N_11435,N_8848,N_5260);
xor U11436 (N_11436,N_6818,N_7377);
or U11437 (N_11437,N_8259,N_7850);
nand U11438 (N_11438,N_5048,N_8381);
or U11439 (N_11439,N_8367,N_9350);
nand U11440 (N_11440,N_8645,N_5623);
nor U11441 (N_11441,N_8440,N_7813);
or U11442 (N_11442,N_5656,N_5429);
and U11443 (N_11443,N_8012,N_7052);
nor U11444 (N_11444,N_5456,N_5919);
xor U11445 (N_11445,N_6733,N_9539);
nor U11446 (N_11446,N_6608,N_9197);
nor U11447 (N_11447,N_6682,N_8271);
and U11448 (N_11448,N_9364,N_8279);
and U11449 (N_11449,N_5900,N_6966);
nand U11450 (N_11450,N_8427,N_6932);
xnor U11451 (N_11451,N_9251,N_5749);
nand U11452 (N_11452,N_8774,N_7092);
and U11453 (N_11453,N_8571,N_6364);
and U11454 (N_11454,N_6142,N_5314);
xnor U11455 (N_11455,N_7198,N_9828);
nand U11456 (N_11456,N_7721,N_9935);
xor U11457 (N_11457,N_8559,N_9834);
xor U11458 (N_11458,N_7005,N_7781);
xor U11459 (N_11459,N_8240,N_9981);
xor U11460 (N_11460,N_8217,N_8771);
or U11461 (N_11461,N_8808,N_5159);
or U11462 (N_11462,N_8702,N_6746);
nand U11463 (N_11463,N_5142,N_9671);
nor U11464 (N_11464,N_6841,N_9942);
and U11465 (N_11465,N_5096,N_9955);
and U11466 (N_11466,N_9747,N_9045);
xor U11467 (N_11467,N_5381,N_6388);
or U11468 (N_11468,N_9893,N_5685);
and U11469 (N_11469,N_5590,N_9847);
and U11470 (N_11470,N_5845,N_6105);
and U11471 (N_11471,N_9156,N_5431);
or U11472 (N_11472,N_9638,N_6874);
xnor U11473 (N_11473,N_8518,N_9586);
or U11474 (N_11474,N_9464,N_8298);
xnor U11475 (N_11475,N_7581,N_8086);
xnor U11476 (N_11476,N_7834,N_7131);
xor U11477 (N_11477,N_9761,N_6345);
or U11478 (N_11478,N_6156,N_7150);
xnor U11479 (N_11479,N_6444,N_9856);
nand U11480 (N_11480,N_5408,N_7257);
nor U11481 (N_11481,N_5361,N_6214);
xor U11482 (N_11482,N_6557,N_8207);
xnor U11483 (N_11483,N_7082,N_9926);
nor U11484 (N_11484,N_9625,N_8712);
nand U11485 (N_11485,N_5673,N_8979);
and U11486 (N_11486,N_7567,N_7881);
nor U11487 (N_11487,N_6309,N_6471);
nor U11488 (N_11488,N_7604,N_6335);
nor U11489 (N_11489,N_9814,N_7225);
and U11490 (N_11490,N_5499,N_6138);
nor U11491 (N_11491,N_8818,N_6677);
nand U11492 (N_11492,N_5376,N_5561);
or U11493 (N_11493,N_6354,N_7812);
nor U11494 (N_11494,N_5604,N_9763);
and U11495 (N_11495,N_8906,N_8784);
nor U11496 (N_11496,N_9026,N_5213);
or U11497 (N_11497,N_8664,N_5014);
nor U11498 (N_11498,N_5187,N_5465);
nor U11499 (N_11499,N_8423,N_8824);
nor U11500 (N_11500,N_9037,N_8988);
and U11501 (N_11501,N_7868,N_8211);
nand U11502 (N_11502,N_5512,N_6930);
xnor U11503 (N_11503,N_6409,N_5375);
nor U11504 (N_11504,N_9160,N_5829);
and U11505 (N_11505,N_6191,N_5346);
nand U11506 (N_11506,N_7037,N_5574);
or U11507 (N_11507,N_7533,N_9533);
xor U11508 (N_11508,N_5799,N_9070);
xor U11509 (N_11509,N_9976,N_6641);
and U11510 (N_11510,N_7982,N_9563);
xnor U11511 (N_11511,N_7521,N_7312);
nand U11512 (N_11512,N_9094,N_9259);
nand U11513 (N_11513,N_9097,N_9706);
nand U11514 (N_11514,N_8456,N_9325);
xor U11515 (N_11515,N_6657,N_7109);
nor U11516 (N_11516,N_9943,N_9447);
nor U11517 (N_11517,N_6658,N_6495);
nor U11518 (N_11518,N_8370,N_9446);
or U11519 (N_11519,N_5774,N_6265);
and U11520 (N_11520,N_6403,N_5365);
or U11521 (N_11521,N_5552,N_7436);
and U11522 (N_11522,N_6483,N_6346);
or U11523 (N_11523,N_9939,N_6887);
nor U11524 (N_11524,N_7683,N_9500);
nand U11525 (N_11525,N_7302,N_9398);
nor U11526 (N_11526,N_9540,N_8237);
nor U11527 (N_11527,N_6965,N_5153);
nor U11528 (N_11528,N_6338,N_8270);
xor U11529 (N_11529,N_9022,N_8296);
xor U11530 (N_11530,N_9142,N_5827);
nor U11531 (N_11531,N_6903,N_5065);
xor U11532 (N_11532,N_9042,N_8656);
nand U11533 (N_11533,N_7289,N_6170);
xor U11534 (N_11534,N_6049,N_9651);
or U11535 (N_11535,N_9048,N_6108);
nor U11536 (N_11536,N_6097,N_7944);
or U11537 (N_11537,N_8863,N_9227);
and U11538 (N_11538,N_7800,N_7880);
or U11539 (N_11539,N_9440,N_8974);
or U11540 (N_11540,N_9127,N_5335);
and U11541 (N_11541,N_8369,N_9399);
or U11542 (N_11542,N_6508,N_5837);
nor U11543 (N_11543,N_9125,N_9299);
and U11544 (N_11544,N_8061,N_7273);
nor U11545 (N_11545,N_6147,N_6171);
xnor U11546 (N_11546,N_9187,N_6581);
xor U11547 (N_11547,N_5234,N_6432);
nand U11548 (N_11548,N_9721,N_7392);
xor U11549 (N_11549,N_7489,N_7121);
and U11550 (N_11550,N_6775,N_9374);
or U11551 (N_11551,N_5545,N_8151);
xor U11552 (N_11552,N_9764,N_7497);
xnor U11553 (N_11553,N_7593,N_7450);
xor U11554 (N_11554,N_9868,N_5155);
and U11555 (N_11555,N_5555,N_7844);
xor U11556 (N_11556,N_6788,N_8856);
xor U11557 (N_11557,N_8997,N_7011);
nor U11558 (N_11558,N_5914,N_9876);
or U11559 (N_11559,N_7945,N_5179);
nor U11560 (N_11560,N_5200,N_9429);
xnor U11561 (N_11561,N_6083,N_8919);
nor U11562 (N_11562,N_9681,N_9741);
nor U11563 (N_11563,N_6433,N_5136);
and U11564 (N_11564,N_7545,N_5231);
and U11565 (N_11565,N_8544,N_5484);
xnor U11566 (N_11566,N_7817,N_6754);
nand U11567 (N_11567,N_5366,N_7320);
and U11568 (N_11568,N_6251,N_5553);
nor U11569 (N_11569,N_7508,N_7505);
xor U11570 (N_11570,N_5675,N_6724);
xnor U11571 (N_11571,N_5343,N_9609);
nor U11572 (N_11572,N_8585,N_8723);
nand U11573 (N_11573,N_9547,N_5297);
nand U11574 (N_11574,N_7006,N_6803);
and U11575 (N_11575,N_7820,N_7549);
or U11576 (N_11576,N_5732,N_5292);
and U11577 (N_11577,N_7615,N_8435);
nor U11578 (N_11578,N_7931,N_7985);
or U11579 (N_11579,N_6000,N_6136);
or U11580 (N_11580,N_7066,N_6886);
and U11581 (N_11581,N_9302,N_9810);
and U11582 (N_11582,N_5933,N_7349);
and U11583 (N_11583,N_6520,N_7352);
or U11584 (N_11584,N_8681,N_9445);
and U11585 (N_11585,N_8872,N_6260);
nand U11586 (N_11586,N_6197,N_5938);
nand U11587 (N_11587,N_5255,N_9528);
or U11588 (N_11588,N_6357,N_9723);
nor U11589 (N_11589,N_7719,N_8244);
nor U11590 (N_11590,N_6793,N_7420);
nor U11591 (N_11591,N_7088,N_7831);
or U11592 (N_11592,N_9118,N_7147);
or U11593 (N_11593,N_6970,N_6597);
nand U11594 (N_11594,N_5506,N_8678);
or U11595 (N_11595,N_6996,N_8090);
xor U11596 (N_11596,N_8387,N_7682);
xnor U11597 (N_11597,N_6934,N_5873);
and U11598 (N_11598,N_5668,N_5432);
xor U11599 (N_11599,N_8006,N_5435);
nand U11600 (N_11600,N_9557,N_6791);
xor U11601 (N_11601,N_5544,N_8124);
nor U11602 (N_11602,N_8729,N_5940);
nor U11603 (N_11603,N_8648,N_5614);
and U11604 (N_11604,N_7838,N_8738);
or U11605 (N_11605,N_9575,N_8532);
xor U11606 (N_11606,N_8183,N_9340);
nor U11607 (N_11607,N_5283,N_6169);
and U11608 (N_11608,N_6467,N_9294);
nor U11609 (N_11609,N_5495,N_5457);
nor U11610 (N_11610,N_7384,N_6294);
xnor U11611 (N_11611,N_8886,N_5844);
nand U11612 (N_11612,N_5833,N_6745);
nand U11613 (N_11613,N_6159,N_8548);
or U11614 (N_11614,N_5674,N_9287);
nor U11615 (N_11615,N_6713,N_5082);
nor U11616 (N_11616,N_6101,N_9844);
or U11617 (N_11617,N_8495,N_8098);
or U11618 (N_11618,N_5662,N_5628);
or U11619 (N_11619,N_6329,N_9477);
and U11620 (N_11620,N_8881,N_6563);
xor U11621 (N_11621,N_8520,N_9492);
and U11622 (N_11622,N_6061,N_8844);
nor U11623 (N_11623,N_9276,N_8875);
xor U11624 (N_11624,N_5826,N_5809);
nor U11625 (N_11625,N_8620,N_6892);
nand U11626 (N_11626,N_6749,N_7896);
or U11627 (N_11627,N_7792,N_8156);
or U11628 (N_11628,N_7403,N_9597);
nand U11629 (N_11629,N_8613,N_8800);
nand U11630 (N_11630,N_5795,N_7713);
nand U11631 (N_11631,N_8535,N_8672);
and U11632 (N_11632,N_5127,N_5998);
or U11633 (N_11633,N_9608,N_5785);
xor U11634 (N_11634,N_6826,N_7219);
or U11635 (N_11635,N_5497,N_8267);
xnor U11636 (N_11636,N_5226,N_7520);
nand U11637 (N_11637,N_9479,N_9554);
or U11638 (N_11638,N_8934,N_5139);
nand U11639 (N_11639,N_8068,N_6988);
or U11640 (N_11640,N_5351,N_9857);
nand U11641 (N_11641,N_7912,N_8148);
nor U11642 (N_11642,N_7733,N_5646);
and U11643 (N_11643,N_6715,N_8903);
xor U11644 (N_11644,N_6235,N_8481);
or U11645 (N_11645,N_9866,N_8827);
and U11646 (N_11646,N_5466,N_7142);
and U11647 (N_11647,N_5695,N_6710);
nor U11648 (N_11648,N_8153,N_8537);
nand U11649 (N_11649,N_5748,N_7333);
nor U11650 (N_11650,N_7953,N_5580);
xnor U11651 (N_11651,N_7346,N_8015);
nor U11652 (N_11652,N_7839,N_5920);
nor U11653 (N_11653,N_5753,N_6394);
or U11654 (N_11654,N_7391,N_7355);
and U11655 (N_11655,N_8116,N_9768);
xnor U11656 (N_11656,N_5963,N_5766);
and U11657 (N_11657,N_9128,N_9677);
nand U11658 (N_11658,N_9143,N_6026);
or U11659 (N_11659,N_5757,N_5310);
nand U11660 (N_11660,N_5323,N_7079);
nand U11661 (N_11661,N_5714,N_6967);
and U11662 (N_11662,N_6893,N_9945);
xor U11663 (N_11663,N_6946,N_6868);
xnor U11664 (N_11664,N_5254,N_6577);
and U11665 (N_11665,N_8165,N_6991);
nand U11666 (N_11666,N_6429,N_6268);
and U11667 (N_11667,N_9751,N_8651);
nand U11668 (N_11668,N_9675,N_5865);
nor U11669 (N_11669,N_5079,N_5183);
xor U11670 (N_11670,N_6019,N_5918);
xnor U11671 (N_11671,N_6979,N_8812);
or U11672 (N_11672,N_8143,N_8336);
or U11673 (N_11673,N_7369,N_7935);
or U11674 (N_11674,N_6944,N_5161);
xor U11675 (N_11675,N_6382,N_7588);
nand U11676 (N_11676,N_9722,N_5114);
nand U11677 (N_11677,N_5560,N_8222);
nor U11678 (N_11678,N_8003,N_9920);
and U11679 (N_11679,N_7818,N_9106);
or U11680 (N_11680,N_6878,N_5670);
nor U11681 (N_11681,N_8836,N_7014);
xor U11682 (N_11682,N_7433,N_6043);
or U11683 (N_11683,N_7824,N_6456);
or U11684 (N_11684,N_8299,N_8566);
nor U11685 (N_11685,N_7775,N_8172);
or U11686 (N_11686,N_5692,N_5554);
nand U11687 (N_11687,N_6033,N_6705);
xnor U11688 (N_11688,N_8106,N_5539);
xor U11689 (N_11689,N_7998,N_7287);
nand U11690 (N_11690,N_6207,N_5721);
nand U11691 (N_11691,N_7140,N_7984);
or U11692 (N_11692,N_6150,N_8140);
nand U11693 (N_11693,N_9434,N_7186);
and U11694 (N_11694,N_9202,N_5638);
nand U11695 (N_11695,N_9466,N_5172);
nor U11696 (N_11696,N_9133,N_9718);
xnor U11697 (N_11697,N_7518,N_8258);
xor U11698 (N_11698,N_7017,N_7132);
nand U11699 (N_11699,N_6457,N_9351);
nand U11700 (N_11700,N_7744,N_9034);
nand U11701 (N_11701,N_5534,N_5951);
or U11702 (N_11702,N_5112,N_7202);
nor U11703 (N_11703,N_7476,N_9757);
or U11704 (N_11704,N_5010,N_8776);
nor U11705 (N_11705,N_9520,N_5650);
nand U11706 (N_11706,N_9015,N_8746);
or U11707 (N_11707,N_9919,N_6995);
nand U11708 (N_11708,N_6226,N_5163);
and U11709 (N_11709,N_8001,N_8666);
or U11710 (N_11710,N_8773,N_7667);
or U11711 (N_11711,N_9598,N_5954);
xnor U11712 (N_11712,N_8405,N_8397);
xor U11713 (N_11713,N_8938,N_6464);
nand U11714 (N_11714,N_6742,N_9411);
and U11715 (N_11715,N_7493,N_6675);
xnor U11716 (N_11716,N_9623,N_8768);
nand U11717 (N_11717,N_7911,N_7108);
xor U11718 (N_11718,N_6178,N_8753);
xnor U11719 (N_11719,N_7934,N_7477);
nand U11720 (N_11720,N_5972,N_8138);
xnor U11721 (N_11721,N_9709,N_9439);
xnor U11722 (N_11722,N_8899,N_7867);
xnor U11723 (N_11723,N_9089,N_9932);
nor U11724 (N_11724,N_7196,N_8858);
or U11725 (N_11725,N_6412,N_5256);
and U11726 (N_11726,N_7732,N_7209);
or U11727 (N_11727,N_9616,N_6233);
nand U11728 (N_11728,N_9515,N_9030);
xor U11729 (N_11729,N_6455,N_5437);
xnor U11730 (N_11730,N_8790,N_5016);
xor U11731 (N_11731,N_9619,N_8125);
and U11732 (N_11732,N_9283,N_7028);
and U11733 (N_11733,N_9743,N_5701);
and U11734 (N_11734,N_8236,N_5188);
or U11735 (N_11735,N_7031,N_5397);
or U11736 (N_11736,N_9292,N_8089);
and U11737 (N_11737,N_7393,N_6218);
nor U11738 (N_11738,N_9649,N_7407);
nor U11739 (N_11739,N_5788,N_7640);
and U11740 (N_11740,N_5886,N_5559);
and U11741 (N_11741,N_5198,N_5568);
or U11742 (N_11742,N_8200,N_6306);
xnor U11743 (N_11743,N_9971,N_7306);
xor U11744 (N_11744,N_5782,N_9818);
nor U11745 (N_11745,N_7429,N_5444);
or U11746 (N_11746,N_6362,N_9405);
nand U11747 (N_11747,N_7515,N_9970);
or U11748 (N_11748,N_6041,N_7584);
or U11749 (N_11749,N_8031,N_8027);
xor U11750 (N_11750,N_8060,N_8719);
nor U11751 (N_11751,N_5566,N_7595);
or U11752 (N_11752,N_6768,N_7372);
xnor U11753 (N_11753,N_6336,N_8582);
xor U11754 (N_11754,N_6729,N_9370);
nand U11755 (N_11755,N_6425,N_9190);
nand U11756 (N_11756,N_7350,N_9505);
nand U11757 (N_11757,N_7467,N_5253);
or U11758 (N_11758,N_6748,N_9953);
nand U11759 (N_11759,N_7806,N_9319);
and U11760 (N_11760,N_5508,N_7966);
or U11761 (N_11761,N_7080,N_6650);
xnor U11762 (N_11762,N_5412,N_5640);
and U11763 (N_11763,N_5045,N_5316);
or U11764 (N_11764,N_7175,N_8970);
xor U11765 (N_11765,N_7423,N_8890);
xnor U11766 (N_11766,N_5131,N_5022);
nor U11767 (N_11767,N_6570,N_6605);
or U11768 (N_11768,N_6179,N_6616);
nand U11769 (N_11769,N_9443,N_9788);
nand U11770 (N_11770,N_7285,N_8734);
or U11771 (N_11771,N_9797,N_6716);
nand U11772 (N_11772,N_9614,N_9459);
or U11773 (N_11773,N_6411,N_7360);
xnor U11774 (N_11774,N_5311,N_8105);
or U11775 (N_11775,N_7710,N_9599);
xor U11776 (N_11776,N_5487,N_9001);
or U11777 (N_11777,N_5355,N_9511);
nor U11778 (N_11778,N_6143,N_6059);
and U11779 (N_11779,N_7575,N_6172);
xor U11780 (N_11780,N_7968,N_9166);
or U11781 (N_11781,N_8996,N_7621);
or U11782 (N_11782,N_9196,N_6109);
nor U11783 (N_11783,N_7227,N_6696);
nor U11784 (N_11784,N_7676,N_7206);
and U11785 (N_11785,N_8202,N_8653);
xor U11786 (N_11786,N_5930,N_8130);
nand U11787 (N_11787,N_9822,N_9019);
or U11788 (N_11788,N_9163,N_7921);
or U11789 (N_11789,N_5093,N_9602);
and U11790 (N_11790,N_5024,N_9565);
nand U11791 (N_11791,N_6385,N_9016);
nand U11792 (N_11792,N_6771,N_7434);
and U11793 (N_11793,N_8744,N_8737);
nand U11794 (N_11794,N_8042,N_9424);
or U11795 (N_11795,N_7905,N_9337);
nand U11796 (N_11796,N_6199,N_8072);
nor U11797 (N_11797,N_9766,N_8234);
xnor U11798 (N_11798,N_9699,N_9192);
xnor U11799 (N_11799,N_5822,N_8911);
nor U11800 (N_11800,N_6331,N_8411);
and U11801 (N_11801,N_9074,N_6532);
xor U11802 (N_11802,N_5438,N_5294);
and U11803 (N_11803,N_7991,N_5374);
or U11804 (N_11804,N_9688,N_8536);
nor U11805 (N_11805,N_6913,N_6902);
and U11806 (N_11806,N_7873,N_9727);
xnor U11807 (N_11807,N_5217,N_5887);
nor U11808 (N_11808,N_6274,N_6823);
nand U11809 (N_11809,N_5592,N_8199);
and U11810 (N_11810,N_6809,N_5843);
nand U11811 (N_11811,N_7475,N_7951);
xnor U11812 (N_11812,N_6091,N_9471);
or U11813 (N_11813,N_9470,N_6020);
and U11814 (N_11814,N_9993,N_7708);
or U11815 (N_11815,N_5406,N_7018);
nor U11816 (N_11816,N_7143,N_9168);
xor U11817 (N_11817,N_7074,N_8490);
and U11818 (N_11818,N_6687,N_6182);
and U11819 (N_11819,N_5318,N_6160);
xor U11820 (N_11820,N_7122,N_6960);
and U11821 (N_11821,N_6320,N_7373);
or U11822 (N_11822,N_9647,N_8985);
nand U11823 (N_11823,N_8632,N_7062);
xor U11824 (N_11824,N_7579,N_5109);
or U11825 (N_11825,N_6132,N_5967);
nor U11826 (N_11826,N_6460,N_5002);
or U11827 (N_11827,N_5104,N_9305);
or U11828 (N_11828,N_9369,N_7107);
xor U11829 (N_11829,N_6469,N_8898);
nor U11830 (N_11830,N_6262,N_8506);
and U11831 (N_11831,N_9679,N_5138);
nand U11832 (N_11832,N_5557,N_7835);
and U11833 (N_11833,N_5762,N_6815);
nand U11834 (N_11834,N_7376,N_7932);
nand U11835 (N_11835,N_5069,N_5622);
xor U11836 (N_11836,N_5932,N_7152);
or U11837 (N_11837,N_5706,N_5445);
nand U11838 (N_11838,N_5225,N_5630);
nor U11839 (N_11839,N_8485,N_5317);
xor U11840 (N_11840,N_9184,N_7212);
and U11841 (N_11841,N_7894,N_8978);
and U11842 (N_11842,N_8480,N_5398);
nor U11843 (N_11843,N_6493,N_9161);
nand U11844 (N_11844,N_8135,N_5815);
or U11845 (N_11845,N_6162,N_6219);
nor U11846 (N_11846,N_7961,N_8311);
nor U11847 (N_11847,N_5619,N_5517);
nand U11848 (N_11848,N_6829,N_9217);
nand U11849 (N_11849,N_8907,N_6594);
or U11850 (N_11850,N_9496,N_9742);
nor U11851 (N_11851,N_7809,N_9108);
xnor U11852 (N_11852,N_8472,N_9559);
and U11853 (N_11853,N_5654,N_9437);
xor U11854 (N_11854,N_9297,N_7973);
nor U11855 (N_11855,N_7576,N_7779);
and U11856 (N_11856,N_9146,N_6691);
xnor U11857 (N_11857,N_9062,N_6008);
nor U11858 (N_11858,N_9646,N_6924);
xnor U11859 (N_11859,N_6377,N_6583);
or U11860 (N_11860,N_6096,N_5857);
nor U11861 (N_11861,N_8647,N_8762);
nand U11862 (N_11862,N_5452,N_5916);
nor U11863 (N_11863,N_7558,N_9359);
xor U11864 (N_11864,N_7656,N_8799);
and U11865 (N_11865,N_8659,N_6731);
or U11866 (N_11866,N_8332,N_7677);
nor U11867 (N_11867,N_8310,N_7462);
or U11868 (N_11868,N_7665,N_7364);
and U11869 (N_11869,N_7642,N_9604);
nor U11870 (N_11870,N_6900,N_6666);
xor U11871 (N_11871,N_7455,N_9767);
nor U11872 (N_11872,N_8690,N_7495);
and U11873 (N_11873,N_6187,N_9231);
or U11874 (N_11874,N_8751,N_7989);
nor U11875 (N_11875,N_5598,N_5367);
and U11876 (N_11876,N_9352,N_5664);
and U11877 (N_11877,N_8530,N_7672);
and U11878 (N_11878,N_6813,N_9420);
xor U11879 (N_11879,N_6504,N_9072);
nor U11880 (N_11880,N_9927,N_6888);
nor U11881 (N_11881,N_8834,N_7486);
and U11882 (N_11882,N_5507,N_7035);
nor U11883 (N_11883,N_6009,N_6401);
xor U11884 (N_11884,N_8376,N_6712);
and U11885 (N_11885,N_7087,N_7033);
nor U11886 (N_11886,N_8393,N_6375);
xor U11887 (N_11887,N_8055,N_7488);
xnor U11888 (N_11888,N_9795,N_9897);
nand U11889 (N_11889,N_8493,N_7794);
nor U11890 (N_11890,N_6700,N_8285);
and U11891 (N_11891,N_9762,N_9545);
and U11892 (N_11892,N_5915,N_7374);
nor U11893 (N_11893,N_7611,N_8329);
xnor U11894 (N_11894,N_5770,N_9864);
nand U11895 (N_11895,N_5201,N_6732);
and U11896 (N_11896,N_9984,N_7815);
and U11897 (N_11897,N_6604,N_6567);
or U11898 (N_11898,N_8569,N_8777);
or U11899 (N_11899,N_6419,N_6435);
xnor U11900 (N_11900,N_6692,N_8330);
nor U11901 (N_11901,N_7696,N_5268);
nor U11902 (N_11902,N_5763,N_8743);
nor U11903 (N_11903,N_8910,N_9182);
xnor U11904 (N_11904,N_8599,N_7698);
xor U11905 (N_11905,N_8058,N_9111);
or U11906 (N_11906,N_5463,N_9686);
nand U11907 (N_11907,N_7883,N_7405);
nand U11908 (N_11908,N_8195,N_6396);
nor U11909 (N_11909,N_9966,N_6702);
or U11910 (N_11910,N_7100,N_9105);
or U11911 (N_11911,N_8066,N_7754);
xor U11912 (N_11912,N_5642,N_9407);
nand U11913 (N_11913,N_8181,N_6975);
and U11914 (N_11914,N_5686,N_6931);
or U11915 (N_11915,N_8561,N_9028);
nor U11916 (N_11916,N_7123,N_6276);
nor U11917 (N_11917,N_9098,N_7394);
and U11918 (N_11918,N_5037,N_5601);
nor U11919 (N_11919,N_5384,N_5221);
nand U11920 (N_11920,N_9820,N_6250);
and U11921 (N_11921,N_9258,N_6802);
nor U11922 (N_11922,N_9372,N_6263);
xor U11923 (N_11923,N_7987,N_7381);
or U11924 (N_11924,N_8543,N_7072);
and U11925 (N_11925,N_9490,N_8725);
xnor U11926 (N_11926,N_7277,N_6185);
xor U11927 (N_11927,N_5442,N_5955);
nand U11928 (N_11928,N_9228,N_9066);
and U11929 (N_11929,N_5859,N_7591);
xor U11930 (N_11930,N_6368,N_5531);
and U11931 (N_11931,N_6228,N_9078);
or U11932 (N_11932,N_9007,N_8628);
or U11933 (N_11933,N_7551,N_8038);
xor U11934 (N_11934,N_5098,N_5677);
nor U11935 (N_11935,N_5787,N_6102);
nand U11936 (N_11936,N_5513,N_6684);
or U11937 (N_11937,N_5052,N_6725);
nand U11938 (N_11938,N_6122,N_8449);
nand U11939 (N_11939,N_5537,N_5836);
and U11940 (N_11940,N_9958,N_7236);
or U11941 (N_11941,N_6709,N_9929);
and U11942 (N_11942,N_5038,N_7187);
and U11943 (N_11943,N_7705,N_9590);
nand U11944 (N_11944,N_9040,N_5832);
or U11945 (N_11945,N_7995,N_8704);
nor U11946 (N_11946,N_9109,N_7854);
xor U11947 (N_11947,N_6681,N_6774);
or U11948 (N_11948,N_8187,N_8147);
and U11949 (N_11949,N_6572,N_9924);
or U11950 (N_11950,N_6734,N_7745);
or U11951 (N_11951,N_5416,N_9063);
nor U11952 (N_11952,N_9964,N_8302);
or U11953 (N_11953,N_7409,N_8795);
xor U11954 (N_11954,N_5245,N_8401);
or U11955 (N_11955,N_5791,N_7543);
nor U11956 (N_11956,N_9248,N_8477);
xnor U11957 (N_11957,N_7191,N_7933);
nor U11958 (N_11958,N_5718,N_5178);
nor U11959 (N_11959,N_6047,N_8752);
nand U11960 (N_11960,N_6899,N_7443);
or U11961 (N_11961,N_6586,N_8917);
nor U11962 (N_11962,N_8512,N_8351);
xor U11963 (N_11963,N_8312,N_7612);
nor U11964 (N_11964,N_7895,N_6805);
and U11965 (N_11965,N_9936,N_7727);
nor U11966 (N_11966,N_5189,N_8441);
nand U11967 (N_11967,N_5808,N_6222);
and U11968 (N_11968,N_7783,N_6927);
and U11969 (N_11969,N_5997,N_9950);
and U11970 (N_11970,N_8347,N_5291);
xnor U11971 (N_11971,N_6683,N_5564);
and U11972 (N_11972,N_9907,N_7695);
xor U11973 (N_11973,N_9886,N_9131);
nand U11974 (N_11974,N_5230,N_6546);
xnor U11975 (N_11975,N_5882,N_7926);
xor U11976 (N_11976,N_5999,N_7473);
nand U11977 (N_11977,N_8079,N_9991);
nor U11978 (N_11978,N_8814,N_8126);
nand U11979 (N_11979,N_7460,N_8811);
nor U11980 (N_11980,N_7740,N_8670);
nor U11981 (N_11981,N_8873,N_9527);
xor U11982 (N_11982,N_5563,N_7110);
and U11983 (N_11983,N_7324,N_8691);
xor U11984 (N_11984,N_9068,N_8078);
or U11985 (N_11985,N_5649,N_6824);
or U11986 (N_11986,N_8462,N_9974);
and U11987 (N_11987,N_5852,N_8922);
or U11988 (N_11988,N_9130,N_5000);
nand U11989 (N_11989,N_7589,N_8371);
or U11990 (N_11990,N_9357,N_5973);
or U11991 (N_11991,N_7983,N_9295);
nor U11992 (N_11992,N_6094,N_7095);
nor U11993 (N_11993,N_5667,N_9667);
nand U11994 (N_11994,N_7517,N_6196);
and U11995 (N_11995,N_8698,N_8294);
or U11996 (N_11996,N_5057,N_5169);
or U11997 (N_11997,N_8224,N_5208);
and U11998 (N_11998,N_9221,N_5934);
nand U11999 (N_11999,N_9592,N_8951);
nand U12000 (N_12000,N_7980,N_7568);
or U12001 (N_12001,N_5790,N_6632);
and U12002 (N_12002,N_9503,N_7286);
nor U12003 (N_12003,N_9852,N_7582);
or U12004 (N_12004,N_6885,N_7541);
nor U12005 (N_12005,N_8589,N_5903);
and U12006 (N_12006,N_5489,N_9770);
or U12007 (N_12007,N_9310,N_9218);
nand U12008 (N_12008,N_9172,N_6086);
or U12009 (N_12009,N_7387,N_6523);
and U12010 (N_12010,N_9543,N_9317);
nor U12011 (N_12011,N_7669,N_9060);
xnor U12012 (N_12012,N_9645,N_6380);
nor U12013 (N_12013,N_8851,N_9812);
or U12014 (N_12014,N_7832,N_9412);
nor U12015 (N_12015,N_5577,N_8705);
xnor U12016 (N_12016,N_7836,N_6704);
nor U12017 (N_12017,N_8174,N_7178);
nand U12018 (N_12018,N_8550,N_8019);
or U12019 (N_12019,N_5405,N_8013);
or U12020 (N_12020,N_5777,N_5080);
nor U12021 (N_12021,N_9534,N_6777);
or U12022 (N_12022,N_5896,N_9803);
or U12023 (N_12023,N_7396,N_5971);
and U12024 (N_12024,N_8159,N_7464);
xor U12025 (N_12025,N_8953,N_7598);
or U12026 (N_12026,N_9589,N_7274);
and U12027 (N_12027,N_9858,N_7524);
and U12028 (N_12028,N_9663,N_5326);
and U12029 (N_12029,N_5682,N_9549);
and U12030 (N_12030,N_5498,N_5985);
and U12031 (N_12031,N_8438,N_7586);
xor U12032 (N_12032,N_9977,N_9871);
nand U12033 (N_12033,N_7240,N_6424);
and U12034 (N_12034,N_8960,N_6490);
xnor U12035 (N_12035,N_9104,N_7970);
nor U12036 (N_12036,N_9307,N_9478);
and U12037 (N_12037,N_5603,N_9652);
or U12038 (N_12038,N_6130,N_5223);
and U12039 (N_12039,N_9692,N_9482);
and U12040 (N_12040,N_6025,N_8273);
or U12041 (N_12041,N_8699,N_7563);
and U12042 (N_12042,N_9164,N_6056);
or U12043 (N_12043,N_6399,N_9099);
nand U12044 (N_12044,N_9642,N_6028);
nand U12045 (N_12045,N_9462,N_8915);
nor U12046 (N_12046,N_5847,N_7903);
and U12047 (N_12047,N_5625,N_6031);
nor U12048 (N_12048,N_5547,N_9896);
nand U12049 (N_12049,N_7484,N_8386);
xor U12050 (N_12050,N_7239,N_7620);
xor U12051 (N_12051,N_5458,N_8103);
and U12052 (N_12052,N_7453,N_7752);
nand U12053 (N_12053,N_8171,N_7546);
and U12054 (N_12054,N_8514,N_8107);
and U12055 (N_12055,N_8320,N_7307);
xnor U12056 (N_12056,N_7021,N_7559);
xor U12057 (N_12057,N_9799,N_7580);
nand U12058 (N_12058,N_6628,N_7583);
xor U12059 (N_12059,N_5373,N_7139);
nor U12060 (N_12060,N_8674,N_9918);
or U12061 (N_12061,N_8720,N_5824);
nand U12062 (N_12062,N_9798,N_8980);
xor U12063 (N_12063,N_7675,N_5975);
or U12064 (N_12064,N_7177,N_6279);
nand U12065 (N_12065,N_8516,N_8823);
or U12066 (N_12066,N_8994,N_9472);
or U12067 (N_12067,N_7587,N_8565);
or U12068 (N_12068,N_5304,N_6919);
and U12069 (N_12069,N_7764,N_6286);
or U12070 (N_12070,N_8767,N_9997);
and U12071 (N_12071,N_9744,N_8505);
nand U12072 (N_12072,N_6010,N_6852);
or U12073 (N_12073,N_6473,N_9748);
nand U12074 (N_12074,N_6184,N_7169);
nand U12075 (N_12075,N_5736,N_9314);
nor U12076 (N_12076,N_5779,N_6638);
and U12077 (N_12077,N_6021,N_7774);
xor U12078 (N_12078,N_6164,N_7043);
nor U12079 (N_12079,N_9404,N_8954);
xnor U12080 (N_12080,N_7616,N_5415);
nor U12081 (N_12081,N_9296,N_8024);
nor U12082 (N_12082,N_8136,N_8801);
xnor U12083 (N_12083,N_7348,N_6722);
nor U12084 (N_12084,N_5942,N_5470);
and U12085 (N_12085,N_9485,N_8961);
nand U12086 (N_12086,N_6827,N_5728);
nand U12087 (N_12087,N_6075,N_6376);
xor U12088 (N_12088,N_6074,N_7104);
or U12089 (N_12089,N_5239,N_8168);
nand U12090 (N_12090,N_5091,N_5103);
and U12091 (N_12091,N_6939,N_7857);
nand U12092 (N_12092,N_5147,N_8241);
nor U12093 (N_12093,N_5910,N_5120);
xnor U12094 (N_12094,N_7365,N_6449);
nand U12095 (N_12095,N_5235,N_7112);
or U12096 (N_12096,N_6165,N_8640);
and U12097 (N_12097,N_7750,N_7023);
nor U12098 (N_12098,N_8226,N_5154);
nor U12099 (N_12099,N_6173,N_7734);
nor U12100 (N_12100,N_7356,N_8070);
nor U12101 (N_12101,N_8314,N_8496);
and U12102 (N_12102,N_7341,N_5086);
or U12103 (N_12103,N_6496,N_5720);
or U12104 (N_12104,N_5205,N_8091);
nand U12105 (N_12105,N_6846,N_6462);
nor U12106 (N_12106,N_6528,N_5651);
nand U12107 (N_12107,N_8986,N_9282);
xor U12108 (N_12108,N_7247,N_9982);
xor U12109 (N_12109,N_5282,N_5126);
nor U12110 (N_12110,N_9693,N_6468);
nor U12111 (N_12111,N_8718,N_6663);
nor U12112 (N_12112,N_8465,N_5267);
nand U12113 (N_12113,N_5793,N_9687);
and U12114 (N_12114,N_7083,N_8568);
nand U12115 (N_12115,N_7538,N_7135);
nand U12116 (N_12116,N_5215,N_8280);
xor U12117 (N_12117,N_5056,N_7297);
nand U12118 (N_12118,N_8791,N_6571);
and U12119 (N_12119,N_8643,N_7742);
and U12120 (N_12120,N_9594,N_5965);
or U12121 (N_12121,N_9662,N_7057);
nand U12122 (N_12122,N_6395,N_7406);
nand U12123 (N_12123,N_5811,N_8056);
nor U12124 (N_12124,N_5876,N_5070);
xnor U12125 (N_12125,N_7748,N_9239);
or U12126 (N_12126,N_7499,N_6639);
xnor U12127 (N_12127,N_5135,N_9354);
nor U12128 (N_12128,N_7097,N_9339);
and U12129 (N_12129,N_8948,N_8742);
nor U12130 (N_12130,N_7644,N_9055);
nand U12131 (N_12131,N_6655,N_7081);
or U12132 (N_12132,N_6044,N_6479);
xnor U12133 (N_12133,N_7689,N_8265);
and U12134 (N_12134,N_9149,N_8641);
nor U12135 (N_12135,N_7739,N_5996);
and U12136 (N_12136,N_5657,N_8840);
or U12137 (N_12137,N_7316,N_7157);
nand U12138 (N_12138,N_8697,N_8478);
and U12139 (N_12139,N_7193,N_5548);
xor U12140 (N_12140,N_5912,N_7482);
nor U12141 (N_12141,N_7624,N_5989);
xnor U12142 (N_12142,N_6855,N_9567);
nor U12143 (N_12143,N_9080,N_7668);
or U12144 (N_12144,N_5050,N_5684);
nand U12145 (N_12145,N_9204,N_8935);
xnor U12146 (N_12146,N_8220,N_8944);
nor U12147 (N_12147,N_6037,N_8607);
and U12148 (N_12148,N_8420,N_8432);
xor U12149 (N_12149,N_5206,N_7009);
and U12150 (N_12150,N_5870,N_8488);
nor U12151 (N_12151,N_5926,N_5195);
xnor U12152 (N_12152,N_9436,N_9165);
nand U12153 (N_12153,N_8579,N_5550);
xor U12154 (N_12154,N_8741,N_5246);
and U12155 (N_12155,N_9669,N_5884);
or U12156 (N_12156,N_8075,N_9753);
nand U12157 (N_12157,N_9569,N_7761);
or U12158 (N_12158,N_8316,N_5073);
xor U12159 (N_12159,N_6351,N_7763);
and U12160 (N_12160,N_6451,N_7118);
and U12161 (N_12161,N_9441,N_8023);
and U12162 (N_12162,N_9952,N_6253);
nor U12163 (N_12163,N_9808,N_6053);
xor U12164 (N_12164,N_9320,N_5970);
nand U12165 (N_12165,N_5059,N_5395);
and U12166 (N_12166,N_9189,N_5765);
xnor U12167 (N_12167,N_8789,N_5735);
nand U12168 (N_12168,N_9488,N_6574);
nor U12169 (N_12169,N_8679,N_9774);
and U12170 (N_12170,N_7979,N_7469);
and U12171 (N_12171,N_5041,N_6747);
nor U12172 (N_12172,N_6070,N_5333);
and U12173 (N_12173,N_8065,N_7294);
and U12174 (N_12174,N_7002,N_6989);
and U12175 (N_12175,N_8359,N_5983);
or U12176 (N_12176,N_8160,N_6318);
nand U12177 (N_12177,N_8816,N_5792);
nor U12178 (N_12178,N_9384,N_7063);
xor U12179 (N_12179,N_5176,N_6728);
and U12180 (N_12180,N_9610,N_5203);
and U12181 (N_12181,N_7444,N_8846);
nor U12182 (N_12182,N_6353,N_7577);
or U12183 (N_12183,N_6463,N_9780);
xnor U12184 (N_12184,N_5115,N_5960);
nor U12185 (N_12185,N_7936,N_6872);
nand U12186 (N_12186,N_8046,N_9135);
xor U12187 (N_12187,N_6881,N_9288);
nor U12188 (N_12188,N_8837,N_5181);
and U12189 (N_12189,N_6076,N_9086);
or U12190 (N_12190,N_8671,N_6656);
nor U12191 (N_12191,N_5969,N_6600);
nand U12192 (N_12192,N_5329,N_6516);
and U12193 (N_12193,N_9327,N_8990);
nor U12194 (N_12194,N_7516,N_5959);
nand U12195 (N_12195,N_8382,N_9634);
nor U12196 (N_12196,N_5441,N_8453);
xor U12197 (N_12197,N_6181,N_7357);
and U12198 (N_12198,N_7597,N_8706);
and U12199 (N_12199,N_5388,N_9050);
xnor U12200 (N_12200,N_8629,N_5486);
or U12201 (N_12201,N_9061,N_8673);
nor U12202 (N_12202,N_8047,N_5639);
or U12203 (N_12203,N_8610,N_6358);
or U12204 (N_12204,N_7971,N_7070);
or U12205 (N_12205,N_5936,N_6626);
nand U12206 (N_12206,N_5337,N_5825);
nor U12207 (N_12207,N_5814,N_5722);
xnor U12208 (N_12208,N_8658,N_6328);
or U12209 (N_12209,N_6592,N_7456);
xor U12210 (N_12210,N_5994,N_8817);
nand U12211 (N_12211,N_6595,N_5110);
nor U12212 (N_12212,N_7362,N_8511);
xor U12213 (N_12213,N_9132,N_6272);
and U12214 (N_12214,N_8071,N_7686);
xnor U12215 (N_12215,N_9185,N_6922);
xnor U12216 (N_12216,N_6480,N_6217);
nor U12217 (N_12217,N_5618,N_6081);
and U12218 (N_12218,N_6507,N_6112);
nor U12219 (N_12219,N_5680,N_7886);
and U12220 (N_12220,N_6322,N_7757);
nand U12221 (N_12221,N_8654,N_6814);
or U12222 (N_12222,N_9235,N_9716);
nand U12223 (N_12223,N_6615,N_9311);
or U12224 (N_12224,N_6206,N_5006);
nand U12225 (N_12225,N_7323,N_6332);
nand U12226 (N_12226,N_6230,N_9978);
or U12227 (N_12227,N_7321,N_7778);
xor U12228 (N_12228,N_6120,N_8695);
xor U12229 (N_12229,N_5197,N_8088);
and U12230 (N_12230,N_6125,N_5313);
nand U12231 (N_12231,N_6198,N_7188);
and U12232 (N_12232,N_5119,N_7359);
or U12233 (N_12233,N_5921,N_9318);
or U12234 (N_12234,N_9002,N_5744);
nor U12235 (N_12235,N_9729,N_8114);
and U12236 (N_12236,N_6593,N_6275);
nand U12237 (N_12237,N_6879,N_9290);
and U12238 (N_12238,N_7158,N_7280);
and U12239 (N_12239,N_6281,N_5669);
or U12240 (N_12240,N_8528,N_5107);
or U12241 (N_12241,N_7592,N_8627);
and U12242 (N_12242,N_9552,N_5321);
nand U12243 (N_12243,N_9717,N_6113);
and U12244 (N_12244,N_5575,N_9529);
nand U12245 (N_12245,N_6643,N_5681);
or U12246 (N_12246,N_7205,N_7788);
nand U12247 (N_12247,N_8539,N_9027);
nor U12248 (N_12248,N_7940,N_6544);
and U12249 (N_12249,N_9879,N_7609);
or U12250 (N_12250,N_5764,N_7878);
nand U12251 (N_12251,N_7657,N_7909);
xor U12252 (N_12252,N_9083,N_6898);
or U12253 (N_12253,N_9058,N_6664);
and U12254 (N_12254,N_9336,N_5157);
nand U12255 (N_12255,N_6255,N_8879);
and U12256 (N_12256,N_6857,N_9845);
or U12257 (N_12257,N_9081,N_9435);
nand U12258 (N_12258,N_8467,N_6772);
and U12259 (N_12259,N_9121,N_6337);
or U12260 (N_12260,N_6071,N_7688);
xnor U12261 (N_12261,N_7914,N_6474);
and U12262 (N_12262,N_6438,N_8605);
nand U12263 (N_12263,N_7342,N_7331);
nor U12264 (N_12264,N_9151,N_8877);
nor U12265 (N_12265,N_6828,N_7458);
nand U12266 (N_12266,N_6529,N_6133);
nand U12267 (N_12267,N_8246,N_7117);
and U12268 (N_12268,N_6642,N_7047);
or U12269 (N_12269,N_7963,N_6288);
xor U12270 (N_12270,N_6794,N_9749);
nand U12271 (N_12271,N_8618,N_8604);
xor U12272 (N_12272,N_5834,N_9418);
nor U12273 (N_12273,N_7972,N_8077);
or U12274 (N_12274,N_9100,N_6257);
nand U12275 (N_12275,N_5979,N_7252);
or U12276 (N_12276,N_7528,N_9698);
nor U12277 (N_12277,N_6305,N_5426);
nand U12278 (N_12278,N_6697,N_8769);
and U12279 (N_12279,N_5644,N_5527);
nand U12280 (N_12280,N_7419,N_5423);
or U12281 (N_12281,N_6564,N_7904);
nor U12282 (N_12282,N_9869,N_5950);
or U12283 (N_12283,N_6220,N_7317);
and U12284 (N_12284,N_8685,N_6962);
or U12285 (N_12285,N_6554,N_7628);
and U12286 (N_12286,N_9555,N_5101);
and U12287 (N_12287,N_8892,N_9588);
nand U12288 (N_12288,N_8541,N_9431);
nand U12289 (N_12289,N_7967,N_8557);
nand U12290 (N_12290,N_6312,N_7025);
nor U12291 (N_12291,N_7756,N_5572);
nand U12292 (N_12292,N_8563,N_9566);
and U12293 (N_12293,N_6158,N_8184);
nor U12294 (N_12294,N_5551,N_7089);
or U12295 (N_12295,N_9954,N_9851);
xor U12296 (N_12296,N_6454,N_9263);
or U12297 (N_12297,N_8484,N_9996);
and U12298 (N_12298,N_6660,N_7199);
nand U12299 (N_12299,N_7957,N_6007);
or U12300 (N_12300,N_7401,N_6726);
or U12301 (N_12301,N_8830,N_7882);
or U12302 (N_12302,N_7416,N_8074);
nor U12303 (N_12303,N_8721,N_6103);
nor U12304 (N_12304,N_9624,N_5752);
xor U12305 (N_12305,N_9715,N_8415);
xor U12306 (N_12306,N_7768,N_8048);
nor U12307 (N_12307,N_8002,N_6977);
or U12308 (N_12308,N_5635,N_5746);
nor U12309 (N_12309,N_9084,N_8407);
and U12310 (N_12310,N_5576,N_9962);
or U12311 (N_12311,N_8043,N_7746);
nand U12312 (N_12312,N_8178,N_5167);
or U12313 (N_12313,N_8782,N_5584);
xor U12314 (N_12314,N_7013,N_7801);
and U12315 (N_12315,N_6609,N_5492);
xnor U12316 (N_12316,N_6579,N_8578);
and U12317 (N_12317,N_6190,N_7607);
and U12318 (N_12318,N_7876,N_7413);
and U12319 (N_12319,N_8192,N_5727);
xor U12320 (N_12320,N_5340,N_6229);
nand U12321 (N_12321,N_9323,N_8931);
or U12322 (N_12322,N_9274,N_5504);
nor U12323 (N_12323,N_8781,N_9087);
nor U12324 (N_12324,N_7949,N_6699);
nand U12325 (N_12325,N_7078,N_9286);
nand U12326 (N_12326,N_7414,N_9732);
nor U12327 (N_12327,N_7981,N_7666);
and U12328 (N_12328,N_5448,N_7116);
nor U12329 (N_12329,N_6545,N_6189);
xnor U12330 (N_12330,N_5755,N_7954);
nand U12331 (N_12331,N_5535,N_6316);
and U12332 (N_12332,N_7120,N_7480);
xnor U12333 (N_12333,N_8433,N_6511);
nor U12334 (N_12334,N_8952,N_6955);
and U12335 (N_12335,N_9720,N_9682);
xnor U12336 (N_12336,N_6807,N_9091);
xor U12337 (N_12337,N_8444,N_5937);
and U12338 (N_12338,N_9916,N_9461);
nor U12339 (N_12339,N_9676,N_8580);
nand U12340 (N_12340,N_5607,N_6036);
and U12341 (N_12341,N_8770,N_8772);
nor U12342 (N_12342,N_5741,N_8803);
and U12343 (N_12343,N_8646,N_8735);
nor U12344 (N_12344,N_5819,N_9195);
or U12345 (N_12345,N_9746,N_5075);
nand U12346 (N_12346,N_6652,N_7892);
or U12347 (N_12347,N_7145,N_8577);
xor U12348 (N_12348,N_9035,N_7194);
xor U12349 (N_12349,N_5241,N_6248);
nor U12350 (N_12350,N_6192,N_6413);
nand U12351 (N_12351,N_8166,N_9553);
nand U12352 (N_12352,N_7296,N_9881);
nand U12353 (N_12353,N_9387,N_6200);
or U12354 (N_12354,N_5032,N_5289);
nor U12355 (N_12355,N_6916,N_9273);
or U12356 (N_12356,N_6066,N_8404);
nand U12357 (N_12357,N_7203,N_6387);
xnor U12358 (N_12358,N_6907,N_6397);
and U12359 (N_12359,N_9578,N_6465);
and U12360 (N_12360,N_6695,N_5020);
and U12361 (N_12361,N_5904,N_9824);
and U12362 (N_12362,N_8942,N_7950);
and U12363 (N_12363,N_6599,N_5298);
or U12364 (N_12364,N_6833,N_5034);
xnor U12365 (N_12365,N_8813,N_5036);
and U12366 (N_12366,N_9234,N_7617);
nand U12367 (N_12367,N_5128,N_9636);
nand U12368 (N_12368,N_5729,N_5562);
or U12369 (N_12369,N_5286,N_5894);
nor U12370 (N_12370,N_5567,N_6521);
nor U12371 (N_12371,N_5264,N_6750);
or U12372 (N_12372,N_5078,N_9362);
or U12373 (N_12373,N_6123,N_5035);
and U12374 (N_12374,N_6553,N_5451);
xor U12375 (N_12375,N_6416,N_5946);
xnor U12376 (N_12376,N_7172,N_8190);
nor U12377 (N_12377,N_5524,N_5851);
and U12378 (N_12378,N_7554,N_6701);
nand U12379 (N_12379,N_5019,N_6448);
xor U12380 (N_12380,N_9158,N_6004);
xor U12381 (N_12381,N_6737,N_8083);
nor U12382 (N_12382,N_5017,N_8459);
or U12383 (N_12383,N_6923,N_5315);
or U12384 (N_12384,N_5327,N_9342);
nor U12385 (N_12385,N_7054,N_9454);
and U12386 (N_12386,N_8352,N_7913);
nor U12387 (N_12387,N_5863,N_9615);
or U12388 (N_12388,N_9232,N_9683);
or U12389 (N_12389,N_7599,N_8841);
xnor U12390 (N_12390,N_5113,N_8121);
xnor U12391 (N_12391,N_6971,N_9402);
xnor U12392 (N_12392,N_9113,N_5219);
xor U12393 (N_12393,N_8713,N_7332);
nor U12394 (N_12394,N_8025,N_9665);
or U12395 (N_12395,N_5909,N_5364);
xnor U12396 (N_12396,N_8344,N_5703);
and U12397 (N_12397,N_6084,N_9713);
nand U12398 (N_12398,N_7608,N_5242);
nor U12399 (N_12399,N_9591,N_9348);
nand U12400 (N_12400,N_6221,N_5467);
and U12401 (N_12401,N_6866,N_9783);
nand U12402 (N_12402,N_6769,N_9032);
nand U12403 (N_12403,N_6073,N_8717);
or U12404 (N_12404,N_7685,N_7040);
nor U12405 (N_12405,N_6812,N_9300);
and U12406 (N_12406,N_7625,N_9769);
and U12407 (N_12407,N_5026,N_5214);
nand U12408 (N_12408,N_6925,N_6858);
or U12409 (N_12409,N_9051,N_8331);
or U12410 (N_12410,N_8946,N_7134);
or U12411 (N_12411,N_8117,N_7749);
xor U12412 (N_12412,N_7492,N_7851);
xnor U12413 (N_12413,N_9664,N_9177);
nor U12414 (N_12414,N_8588,N_7207);
nand U12415 (N_12415,N_9801,N_9367);
and U12416 (N_12416,N_7816,N_6659);
xnor U12417 (N_12417,N_7585,N_9581);
nand U12418 (N_12418,N_7852,N_5461);
and U12419 (N_12419,N_8290,N_7154);
nand U12420 (N_12420,N_9921,N_9765);
nor U12421 (N_12421,N_8669,N_6981);
xor U12422 (N_12422,N_9980,N_8583);
nand U12423 (N_12423,N_9329,N_8011);
nand U12424 (N_12424,N_7119,N_7522);
and U12425 (N_12425,N_8141,N_5400);
nor U12426 (N_12426,N_9023,N_5679);
xnor U12427 (N_12427,N_8854,N_6245);
nor U12428 (N_12428,N_9065,N_8337);
and U12429 (N_12429,N_7248,N_7315);
and U12430 (N_12430,N_8409,N_9967);
or U12431 (N_12431,N_7155,N_5356);
and U12432 (N_12432,N_7724,N_6285);
xor U12433 (N_12433,N_8424,N_6048);
and U12434 (N_12434,N_9577,N_5864);
xor U12435 (N_12435,N_9728,N_9222);
and U12436 (N_12436,N_5425,N_9895);
nor U12437 (N_12437,N_7938,N_9347);
or U12438 (N_12438,N_7165,N_8815);
xnor U12439 (N_12439,N_5702,N_5330);
nor U12440 (N_12440,N_5660,N_7380);
nor U12441 (N_12441,N_5068,N_9379);
xor U12442 (N_12442,N_8778,N_9162);
and U12443 (N_12443,N_8082,N_5054);
nor U12444 (N_12444,N_6475,N_8621);
and U12445 (N_12445,N_5276,N_7004);
nand U12446 (N_12446,N_6644,N_6928);
or U12447 (N_12447,N_6937,N_8040);
and U12448 (N_12448,N_9003,N_5430);
xnor U12449 (N_12449,N_6740,N_8235);
nand U12450 (N_12450,N_5522,N_6107);
nand U12451 (N_12451,N_6271,N_5558);
nor U12452 (N_12452,N_5199,N_6718);
or U12453 (N_12453,N_6392,N_7138);
or U12454 (N_12454,N_9043,N_8968);
and U12455 (N_12455,N_5723,N_7602);
or U12456 (N_12456,N_9941,N_7526);
nor U12457 (N_12457,N_9129,N_5369);
or U12458 (N_12458,N_7283,N_8225);
xor U12459 (N_12459,N_9889,N_6050);
nor U12460 (N_12460,N_8357,N_8248);
or U12461 (N_12461,N_5360,N_7623);
and U12462 (N_12462,N_9344,N_6510);
xnor U12463 (N_12463,N_9499,N_8144);
xor U12464 (N_12464,N_7084,N_6711);
nor U12465 (N_12465,N_9279,N_9119);
or U12466 (N_12466,N_8943,N_6661);
nand U12467 (N_12467,N_6552,N_5992);
and U12468 (N_12468,N_8937,N_5211);
nor U12469 (N_12469,N_8760,N_7658);
xnor U12470 (N_12470,N_8864,N_6533);
nand U12471 (N_12471,N_8731,N_5044);
nand U12472 (N_12472,N_5518,N_9249);
nor U12473 (N_12473,N_6295,N_9214);
nor U12474 (N_12474,N_9140,N_9835);
or U12475 (N_12475,N_5917,N_7020);
and U12476 (N_12476,N_6227,N_9208);
nor U12477 (N_12477,N_8406,N_7382);
or U12478 (N_12478,N_8392,N_9076);
or U12479 (N_12479,N_6258,N_9497);
xor U12480 (N_12480,N_7706,N_5543);
or U12481 (N_12481,N_8754,N_8213);
xnor U12482 (N_12482,N_7828,N_5842);
nand U12483 (N_12483,N_7560,N_7917);
or U12484 (N_12484,N_6957,N_6555);
nand U12485 (N_12485,N_5659,N_8288);
nand U12486 (N_12486,N_8315,N_5665);
xor U12487 (N_12487,N_8080,N_5319);
nand U12488 (N_12488,N_6673,N_7811);
and U12489 (N_12489,N_5519,N_5705);
nor U12490 (N_12490,N_5587,N_5428);
and U12491 (N_12491,N_5643,N_8398);
xor U12492 (N_12492,N_9291,N_5778);
nand U12493 (N_12493,N_8545,N_6921);
or U12494 (N_12494,N_7663,N_8832);
nor U12495 (N_12495,N_7902,N_9186);
nor U12496 (N_12496,N_9343,N_5935);
or U12497 (N_12497,N_8572,N_8030);
and U12498 (N_12498,N_9690,N_7338);
nor U12499 (N_12499,N_7038,N_5359);
xor U12500 (N_12500,N_8034,N_7214);
and U12501 (N_12501,N_8629,N_9072);
and U12502 (N_12502,N_5140,N_5237);
and U12503 (N_12503,N_8310,N_5007);
nand U12504 (N_12504,N_9421,N_6250);
xor U12505 (N_12505,N_6601,N_8202);
nand U12506 (N_12506,N_7059,N_5995);
and U12507 (N_12507,N_9665,N_9637);
and U12508 (N_12508,N_7930,N_6655);
nor U12509 (N_12509,N_5490,N_7254);
and U12510 (N_12510,N_6745,N_9576);
xor U12511 (N_12511,N_7276,N_7278);
nor U12512 (N_12512,N_6888,N_6239);
nand U12513 (N_12513,N_7276,N_6383);
and U12514 (N_12514,N_5376,N_7822);
or U12515 (N_12515,N_9559,N_6522);
and U12516 (N_12516,N_8450,N_8981);
nor U12517 (N_12517,N_5846,N_6223);
and U12518 (N_12518,N_6690,N_8263);
nor U12519 (N_12519,N_6664,N_7452);
or U12520 (N_12520,N_6555,N_7675);
nor U12521 (N_12521,N_6548,N_7126);
nor U12522 (N_12522,N_9884,N_8740);
nor U12523 (N_12523,N_5216,N_8759);
nand U12524 (N_12524,N_7948,N_8925);
and U12525 (N_12525,N_6986,N_5243);
xnor U12526 (N_12526,N_6337,N_5683);
nand U12527 (N_12527,N_8923,N_6129);
xor U12528 (N_12528,N_9881,N_5649);
nor U12529 (N_12529,N_6142,N_8086);
xnor U12530 (N_12530,N_9035,N_9266);
nor U12531 (N_12531,N_6073,N_7608);
nor U12532 (N_12532,N_9519,N_6836);
xnor U12533 (N_12533,N_8529,N_7765);
nand U12534 (N_12534,N_5121,N_5703);
nand U12535 (N_12535,N_9219,N_6298);
and U12536 (N_12536,N_7459,N_8359);
xnor U12537 (N_12537,N_6412,N_5657);
nor U12538 (N_12538,N_9097,N_7638);
xor U12539 (N_12539,N_5977,N_5501);
or U12540 (N_12540,N_8519,N_6923);
nor U12541 (N_12541,N_7754,N_8664);
xnor U12542 (N_12542,N_7692,N_8986);
or U12543 (N_12543,N_6053,N_9531);
nand U12544 (N_12544,N_6441,N_5384);
and U12545 (N_12545,N_9226,N_9869);
or U12546 (N_12546,N_9246,N_9024);
or U12547 (N_12547,N_9710,N_5994);
and U12548 (N_12548,N_9602,N_6664);
nor U12549 (N_12549,N_9340,N_7016);
or U12550 (N_12550,N_5941,N_8890);
xnor U12551 (N_12551,N_7374,N_9147);
or U12552 (N_12552,N_5974,N_6977);
and U12553 (N_12553,N_8180,N_9019);
nand U12554 (N_12554,N_8327,N_8307);
and U12555 (N_12555,N_9030,N_6528);
or U12556 (N_12556,N_5185,N_5721);
or U12557 (N_12557,N_9507,N_6322);
xnor U12558 (N_12558,N_8631,N_9882);
or U12559 (N_12559,N_5471,N_5753);
and U12560 (N_12560,N_5477,N_5701);
and U12561 (N_12561,N_8652,N_7199);
nor U12562 (N_12562,N_8319,N_5057);
and U12563 (N_12563,N_7731,N_9072);
nor U12564 (N_12564,N_7158,N_9990);
xnor U12565 (N_12565,N_8593,N_5844);
and U12566 (N_12566,N_6275,N_5639);
nand U12567 (N_12567,N_7336,N_6881);
nor U12568 (N_12568,N_6085,N_6131);
or U12569 (N_12569,N_9162,N_8116);
and U12570 (N_12570,N_9732,N_6406);
and U12571 (N_12571,N_7318,N_7933);
xor U12572 (N_12572,N_5663,N_8901);
nand U12573 (N_12573,N_6107,N_6637);
and U12574 (N_12574,N_6796,N_6364);
and U12575 (N_12575,N_7993,N_6099);
nand U12576 (N_12576,N_5788,N_7015);
nand U12577 (N_12577,N_7634,N_9928);
xnor U12578 (N_12578,N_8299,N_8967);
or U12579 (N_12579,N_6891,N_9088);
nor U12580 (N_12580,N_7968,N_6230);
and U12581 (N_12581,N_7781,N_9486);
xor U12582 (N_12582,N_7229,N_8392);
or U12583 (N_12583,N_9804,N_7233);
nor U12584 (N_12584,N_9324,N_5769);
nor U12585 (N_12585,N_9215,N_7158);
nor U12586 (N_12586,N_9220,N_9410);
or U12587 (N_12587,N_6438,N_7043);
and U12588 (N_12588,N_8000,N_5807);
or U12589 (N_12589,N_7914,N_8313);
nand U12590 (N_12590,N_6004,N_6046);
or U12591 (N_12591,N_9826,N_5176);
xor U12592 (N_12592,N_6647,N_9363);
nand U12593 (N_12593,N_6611,N_5107);
or U12594 (N_12594,N_8363,N_9564);
xor U12595 (N_12595,N_5333,N_9014);
xnor U12596 (N_12596,N_5938,N_8399);
and U12597 (N_12597,N_9283,N_6593);
xor U12598 (N_12598,N_5106,N_7526);
nor U12599 (N_12599,N_5545,N_7097);
or U12600 (N_12600,N_8840,N_7040);
nand U12601 (N_12601,N_5843,N_8303);
nor U12602 (N_12602,N_6596,N_7717);
nand U12603 (N_12603,N_5701,N_6813);
nand U12604 (N_12604,N_6004,N_8070);
nor U12605 (N_12605,N_7937,N_5274);
nor U12606 (N_12606,N_7831,N_7420);
and U12607 (N_12607,N_9351,N_6013);
and U12608 (N_12608,N_9651,N_6499);
and U12609 (N_12609,N_8667,N_9541);
nand U12610 (N_12610,N_6304,N_9726);
nor U12611 (N_12611,N_8933,N_7140);
nand U12612 (N_12612,N_6582,N_9406);
nor U12613 (N_12613,N_6205,N_6124);
or U12614 (N_12614,N_8647,N_6597);
xnor U12615 (N_12615,N_7637,N_7589);
and U12616 (N_12616,N_6746,N_8861);
and U12617 (N_12617,N_9585,N_8095);
xnor U12618 (N_12618,N_8529,N_7441);
and U12619 (N_12619,N_5966,N_5320);
and U12620 (N_12620,N_8820,N_5641);
and U12621 (N_12621,N_6788,N_7322);
nand U12622 (N_12622,N_5852,N_7368);
nand U12623 (N_12623,N_5061,N_6409);
or U12624 (N_12624,N_6664,N_9690);
nor U12625 (N_12625,N_9708,N_8563);
and U12626 (N_12626,N_9643,N_6589);
nand U12627 (N_12627,N_6684,N_8324);
or U12628 (N_12628,N_5789,N_5766);
xor U12629 (N_12629,N_7152,N_8348);
xnor U12630 (N_12630,N_5521,N_8854);
and U12631 (N_12631,N_5323,N_8286);
and U12632 (N_12632,N_5917,N_8730);
or U12633 (N_12633,N_8445,N_6562);
or U12634 (N_12634,N_5179,N_9130);
and U12635 (N_12635,N_7504,N_7644);
nand U12636 (N_12636,N_6572,N_8280);
xnor U12637 (N_12637,N_8573,N_5095);
nor U12638 (N_12638,N_9842,N_9796);
and U12639 (N_12639,N_7925,N_7513);
nor U12640 (N_12640,N_7274,N_9535);
nand U12641 (N_12641,N_6592,N_5537);
or U12642 (N_12642,N_7876,N_7475);
nand U12643 (N_12643,N_5430,N_7026);
and U12644 (N_12644,N_9166,N_9293);
nor U12645 (N_12645,N_6083,N_5490);
or U12646 (N_12646,N_6134,N_9872);
xor U12647 (N_12647,N_9515,N_5326);
nand U12648 (N_12648,N_8305,N_8824);
nand U12649 (N_12649,N_5552,N_9106);
or U12650 (N_12650,N_8344,N_8079);
nor U12651 (N_12651,N_6373,N_5105);
xnor U12652 (N_12652,N_5469,N_6935);
or U12653 (N_12653,N_5359,N_8230);
nor U12654 (N_12654,N_9694,N_9863);
or U12655 (N_12655,N_5597,N_8799);
nor U12656 (N_12656,N_7997,N_5193);
nand U12657 (N_12657,N_5305,N_8478);
or U12658 (N_12658,N_8108,N_7565);
or U12659 (N_12659,N_5508,N_7503);
and U12660 (N_12660,N_5383,N_6392);
and U12661 (N_12661,N_8422,N_7783);
and U12662 (N_12662,N_5693,N_6239);
nand U12663 (N_12663,N_8503,N_5803);
nor U12664 (N_12664,N_6039,N_9110);
or U12665 (N_12665,N_8289,N_8339);
nand U12666 (N_12666,N_7509,N_5005);
nor U12667 (N_12667,N_6763,N_5470);
nand U12668 (N_12668,N_7507,N_7797);
nand U12669 (N_12669,N_6082,N_8484);
xnor U12670 (N_12670,N_9203,N_9445);
nand U12671 (N_12671,N_9524,N_8294);
nor U12672 (N_12672,N_6289,N_7360);
nand U12673 (N_12673,N_8172,N_7252);
nor U12674 (N_12674,N_8423,N_7935);
or U12675 (N_12675,N_7894,N_9986);
and U12676 (N_12676,N_7890,N_6413);
and U12677 (N_12677,N_9446,N_5362);
nand U12678 (N_12678,N_8415,N_9970);
or U12679 (N_12679,N_9319,N_6986);
and U12680 (N_12680,N_8086,N_7163);
or U12681 (N_12681,N_9314,N_9532);
nand U12682 (N_12682,N_5910,N_9858);
or U12683 (N_12683,N_7026,N_9245);
or U12684 (N_12684,N_8439,N_7591);
or U12685 (N_12685,N_8908,N_7131);
or U12686 (N_12686,N_8977,N_6022);
nor U12687 (N_12687,N_9647,N_9432);
xnor U12688 (N_12688,N_8779,N_8848);
or U12689 (N_12689,N_8371,N_7312);
nand U12690 (N_12690,N_7366,N_9773);
and U12691 (N_12691,N_9537,N_6393);
or U12692 (N_12692,N_5421,N_6312);
or U12693 (N_12693,N_8609,N_8255);
xor U12694 (N_12694,N_5284,N_5636);
xnor U12695 (N_12695,N_8933,N_6561);
or U12696 (N_12696,N_6310,N_7291);
and U12697 (N_12697,N_9327,N_6369);
and U12698 (N_12698,N_5323,N_5527);
nand U12699 (N_12699,N_7239,N_9321);
and U12700 (N_12700,N_8219,N_8979);
nor U12701 (N_12701,N_8996,N_9813);
xor U12702 (N_12702,N_5718,N_6348);
nand U12703 (N_12703,N_6649,N_5396);
and U12704 (N_12704,N_9573,N_5102);
nand U12705 (N_12705,N_5597,N_5808);
nor U12706 (N_12706,N_8654,N_7663);
nor U12707 (N_12707,N_8157,N_6714);
nor U12708 (N_12708,N_9881,N_7107);
xnor U12709 (N_12709,N_9253,N_8420);
and U12710 (N_12710,N_8831,N_5985);
nand U12711 (N_12711,N_9649,N_7415);
xnor U12712 (N_12712,N_6762,N_8721);
nor U12713 (N_12713,N_6798,N_5876);
nor U12714 (N_12714,N_5277,N_9204);
or U12715 (N_12715,N_9544,N_5816);
or U12716 (N_12716,N_5104,N_8342);
xor U12717 (N_12717,N_6342,N_5008);
nor U12718 (N_12718,N_6106,N_5043);
xnor U12719 (N_12719,N_9575,N_7833);
and U12720 (N_12720,N_5642,N_7812);
nor U12721 (N_12721,N_6503,N_8516);
nand U12722 (N_12722,N_8872,N_8250);
or U12723 (N_12723,N_6510,N_6418);
and U12724 (N_12724,N_5156,N_9876);
xor U12725 (N_12725,N_5380,N_6284);
nor U12726 (N_12726,N_9931,N_5767);
nand U12727 (N_12727,N_6820,N_6342);
nor U12728 (N_12728,N_6267,N_6814);
and U12729 (N_12729,N_6674,N_6425);
and U12730 (N_12730,N_5533,N_5572);
and U12731 (N_12731,N_6674,N_5883);
and U12732 (N_12732,N_5734,N_5599);
and U12733 (N_12733,N_7597,N_6875);
or U12734 (N_12734,N_7110,N_9973);
or U12735 (N_12735,N_7808,N_9557);
nand U12736 (N_12736,N_6447,N_6118);
and U12737 (N_12737,N_5797,N_7655);
and U12738 (N_12738,N_5233,N_7539);
or U12739 (N_12739,N_7894,N_8741);
and U12740 (N_12740,N_5865,N_7954);
and U12741 (N_12741,N_8596,N_7488);
nand U12742 (N_12742,N_6351,N_7894);
or U12743 (N_12743,N_8263,N_8910);
and U12744 (N_12744,N_9902,N_8099);
or U12745 (N_12745,N_8410,N_7586);
nand U12746 (N_12746,N_9387,N_6925);
xor U12747 (N_12747,N_9088,N_5128);
or U12748 (N_12748,N_6329,N_7758);
and U12749 (N_12749,N_8768,N_8218);
and U12750 (N_12750,N_9496,N_8942);
xnor U12751 (N_12751,N_7883,N_6350);
xnor U12752 (N_12752,N_5262,N_8461);
nand U12753 (N_12753,N_8439,N_7824);
xor U12754 (N_12754,N_9914,N_7931);
nor U12755 (N_12755,N_8485,N_5659);
and U12756 (N_12756,N_9732,N_5076);
or U12757 (N_12757,N_6702,N_9820);
nor U12758 (N_12758,N_7110,N_7317);
nor U12759 (N_12759,N_5063,N_8704);
xor U12760 (N_12760,N_7414,N_5174);
or U12761 (N_12761,N_5356,N_8963);
or U12762 (N_12762,N_6372,N_7516);
xor U12763 (N_12763,N_7769,N_9382);
nor U12764 (N_12764,N_9834,N_9163);
and U12765 (N_12765,N_7950,N_5419);
or U12766 (N_12766,N_7300,N_6592);
nor U12767 (N_12767,N_6422,N_8906);
xnor U12768 (N_12768,N_5501,N_7603);
nor U12769 (N_12769,N_7455,N_6067);
nor U12770 (N_12770,N_9484,N_5268);
or U12771 (N_12771,N_7811,N_6664);
or U12772 (N_12772,N_8758,N_6795);
nand U12773 (N_12773,N_9123,N_5176);
xnor U12774 (N_12774,N_9389,N_8519);
xor U12775 (N_12775,N_7691,N_9692);
xnor U12776 (N_12776,N_6889,N_7956);
nor U12777 (N_12777,N_6842,N_6105);
xor U12778 (N_12778,N_6690,N_5987);
xor U12779 (N_12779,N_7058,N_6096);
nor U12780 (N_12780,N_9536,N_7634);
or U12781 (N_12781,N_7879,N_9352);
nor U12782 (N_12782,N_7130,N_5748);
xor U12783 (N_12783,N_5244,N_7808);
nor U12784 (N_12784,N_9680,N_6991);
xor U12785 (N_12785,N_8888,N_6538);
or U12786 (N_12786,N_5795,N_5018);
and U12787 (N_12787,N_6113,N_9760);
nor U12788 (N_12788,N_7173,N_7353);
nand U12789 (N_12789,N_5728,N_5695);
nand U12790 (N_12790,N_6147,N_6430);
or U12791 (N_12791,N_6096,N_8765);
nor U12792 (N_12792,N_5417,N_9755);
and U12793 (N_12793,N_9488,N_7654);
and U12794 (N_12794,N_8724,N_9991);
nor U12795 (N_12795,N_6479,N_9090);
or U12796 (N_12796,N_6359,N_5362);
nand U12797 (N_12797,N_9695,N_8340);
and U12798 (N_12798,N_9227,N_6602);
and U12799 (N_12799,N_9197,N_5643);
and U12800 (N_12800,N_9964,N_7349);
nor U12801 (N_12801,N_5625,N_7577);
or U12802 (N_12802,N_6836,N_8044);
or U12803 (N_12803,N_7864,N_6887);
xnor U12804 (N_12804,N_5285,N_9934);
xor U12805 (N_12805,N_6725,N_5480);
or U12806 (N_12806,N_6864,N_8542);
nor U12807 (N_12807,N_7205,N_7104);
or U12808 (N_12808,N_5897,N_7979);
nand U12809 (N_12809,N_8186,N_8572);
nor U12810 (N_12810,N_7549,N_9601);
nor U12811 (N_12811,N_5048,N_5633);
and U12812 (N_12812,N_6437,N_7938);
and U12813 (N_12813,N_9146,N_9224);
xor U12814 (N_12814,N_9491,N_7597);
xnor U12815 (N_12815,N_9412,N_9968);
nor U12816 (N_12816,N_9101,N_6273);
nor U12817 (N_12817,N_6162,N_8817);
xor U12818 (N_12818,N_5152,N_6750);
xnor U12819 (N_12819,N_8415,N_6432);
nand U12820 (N_12820,N_5361,N_8932);
or U12821 (N_12821,N_6000,N_5437);
nor U12822 (N_12822,N_6052,N_9839);
and U12823 (N_12823,N_7692,N_7762);
or U12824 (N_12824,N_8386,N_7522);
xor U12825 (N_12825,N_7644,N_8371);
or U12826 (N_12826,N_7926,N_8806);
nand U12827 (N_12827,N_6655,N_5399);
nand U12828 (N_12828,N_5315,N_6742);
or U12829 (N_12829,N_5927,N_7351);
and U12830 (N_12830,N_7899,N_7284);
nand U12831 (N_12831,N_7519,N_9666);
or U12832 (N_12832,N_7169,N_8914);
nand U12833 (N_12833,N_7876,N_5190);
xor U12834 (N_12834,N_8516,N_6817);
xor U12835 (N_12835,N_8029,N_6318);
and U12836 (N_12836,N_5541,N_5035);
nand U12837 (N_12837,N_5906,N_9041);
or U12838 (N_12838,N_9440,N_6043);
or U12839 (N_12839,N_7603,N_7392);
or U12840 (N_12840,N_5319,N_8957);
nand U12841 (N_12841,N_6067,N_8809);
nand U12842 (N_12842,N_5276,N_9252);
and U12843 (N_12843,N_6119,N_5411);
or U12844 (N_12844,N_6636,N_5676);
nand U12845 (N_12845,N_6764,N_6901);
nand U12846 (N_12846,N_5220,N_6940);
or U12847 (N_12847,N_8166,N_8460);
nor U12848 (N_12848,N_6680,N_6388);
or U12849 (N_12849,N_5075,N_7669);
xor U12850 (N_12850,N_8076,N_9305);
xor U12851 (N_12851,N_7951,N_7304);
or U12852 (N_12852,N_8697,N_9599);
nor U12853 (N_12853,N_9760,N_5185);
or U12854 (N_12854,N_5814,N_8191);
and U12855 (N_12855,N_9908,N_8141);
or U12856 (N_12856,N_8313,N_9570);
nand U12857 (N_12857,N_8854,N_8517);
nand U12858 (N_12858,N_8408,N_5841);
xor U12859 (N_12859,N_6704,N_8187);
nand U12860 (N_12860,N_5581,N_5132);
and U12861 (N_12861,N_9903,N_8940);
nor U12862 (N_12862,N_5815,N_5125);
nor U12863 (N_12863,N_7792,N_9862);
nor U12864 (N_12864,N_6687,N_5041);
and U12865 (N_12865,N_8882,N_9294);
nand U12866 (N_12866,N_9374,N_7630);
xor U12867 (N_12867,N_7970,N_7333);
and U12868 (N_12868,N_8026,N_8443);
xnor U12869 (N_12869,N_8992,N_6079);
nor U12870 (N_12870,N_6561,N_8450);
nor U12871 (N_12871,N_8148,N_7803);
nand U12872 (N_12872,N_6163,N_6293);
or U12873 (N_12873,N_8867,N_5453);
and U12874 (N_12874,N_6100,N_5258);
xnor U12875 (N_12875,N_7341,N_6765);
nor U12876 (N_12876,N_5633,N_9340);
nand U12877 (N_12877,N_8749,N_8486);
nand U12878 (N_12878,N_6637,N_7597);
xnor U12879 (N_12879,N_7409,N_8603);
and U12880 (N_12880,N_8134,N_6754);
xnor U12881 (N_12881,N_9792,N_5711);
or U12882 (N_12882,N_8995,N_6824);
nand U12883 (N_12883,N_9010,N_9699);
or U12884 (N_12884,N_7349,N_6938);
xor U12885 (N_12885,N_8861,N_7633);
nand U12886 (N_12886,N_8220,N_9804);
nand U12887 (N_12887,N_8727,N_6760);
nor U12888 (N_12888,N_8124,N_5052);
nand U12889 (N_12889,N_7184,N_8137);
and U12890 (N_12890,N_6991,N_6083);
and U12891 (N_12891,N_6885,N_9139);
nand U12892 (N_12892,N_8402,N_6143);
nor U12893 (N_12893,N_6817,N_5233);
or U12894 (N_12894,N_9970,N_8034);
or U12895 (N_12895,N_5407,N_7731);
nand U12896 (N_12896,N_6644,N_9465);
xnor U12897 (N_12897,N_6035,N_6911);
xor U12898 (N_12898,N_6417,N_5684);
nand U12899 (N_12899,N_9274,N_6488);
nand U12900 (N_12900,N_5388,N_7720);
or U12901 (N_12901,N_8142,N_5154);
nand U12902 (N_12902,N_5257,N_8819);
and U12903 (N_12903,N_7072,N_7937);
nor U12904 (N_12904,N_6210,N_6971);
xnor U12905 (N_12905,N_9124,N_5723);
xor U12906 (N_12906,N_9780,N_5223);
or U12907 (N_12907,N_8317,N_5512);
xnor U12908 (N_12908,N_8235,N_6644);
xor U12909 (N_12909,N_7452,N_7848);
nor U12910 (N_12910,N_9370,N_6112);
and U12911 (N_12911,N_8705,N_6574);
nor U12912 (N_12912,N_8994,N_5813);
and U12913 (N_12913,N_9332,N_8919);
nor U12914 (N_12914,N_8399,N_9808);
or U12915 (N_12915,N_7169,N_9322);
and U12916 (N_12916,N_7743,N_5727);
nand U12917 (N_12917,N_7207,N_5136);
nor U12918 (N_12918,N_9974,N_9654);
and U12919 (N_12919,N_5093,N_9648);
xnor U12920 (N_12920,N_6311,N_8719);
and U12921 (N_12921,N_5627,N_6917);
nand U12922 (N_12922,N_5441,N_8123);
xor U12923 (N_12923,N_6181,N_5514);
and U12924 (N_12924,N_5704,N_6159);
nand U12925 (N_12925,N_8393,N_7236);
or U12926 (N_12926,N_8301,N_6298);
and U12927 (N_12927,N_6543,N_6768);
or U12928 (N_12928,N_5414,N_9852);
or U12929 (N_12929,N_5382,N_7968);
xor U12930 (N_12930,N_7283,N_7944);
nor U12931 (N_12931,N_7984,N_5030);
nand U12932 (N_12932,N_8133,N_7375);
and U12933 (N_12933,N_7862,N_6273);
nand U12934 (N_12934,N_5704,N_7686);
nor U12935 (N_12935,N_9200,N_6601);
xnor U12936 (N_12936,N_7509,N_6836);
nand U12937 (N_12937,N_9836,N_6984);
xnor U12938 (N_12938,N_9994,N_7142);
or U12939 (N_12939,N_8036,N_7047);
nand U12940 (N_12940,N_6387,N_6799);
or U12941 (N_12941,N_8991,N_6679);
nor U12942 (N_12942,N_9138,N_9495);
nor U12943 (N_12943,N_6309,N_9446);
xnor U12944 (N_12944,N_9087,N_8016);
xor U12945 (N_12945,N_6012,N_9675);
and U12946 (N_12946,N_9538,N_6801);
nor U12947 (N_12947,N_6406,N_6908);
xor U12948 (N_12948,N_6763,N_8231);
nand U12949 (N_12949,N_9864,N_6073);
xor U12950 (N_12950,N_5578,N_8515);
and U12951 (N_12951,N_6802,N_6562);
and U12952 (N_12952,N_7089,N_6708);
nor U12953 (N_12953,N_6480,N_8315);
or U12954 (N_12954,N_7568,N_7864);
nor U12955 (N_12955,N_5101,N_8249);
and U12956 (N_12956,N_9158,N_8192);
nand U12957 (N_12957,N_7255,N_7366);
nand U12958 (N_12958,N_8444,N_8165);
xor U12959 (N_12959,N_9680,N_7485);
xor U12960 (N_12960,N_9356,N_8732);
nor U12961 (N_12961,N_7154,N_7119);
and U12962 (N_12962,N_9123,N_9290);
nand U12963 (N_12963,N_8255,N_5991);
nor U12964 (N_12964,N_7589,N_5368);
or U12965 (N_12965,N_5628,N_9194);
nand U12966 (N_12966,N_7615,N_7702);
and U12967 (N_12967,N_8403,N_6215);
nor U12968 (N_12968,N_8710,N_9712);
nand U12969 (N_12969,N_7111,N_7791);
and U12970 (N_12970,N_8474,N_9728);
or U12971 (N_12971,N_6703,N_8906);
nand U12972 (N_12972,N_7269,N_6972);
nand U12973 (N_12973,N_9278,N_9059);
nor U12974 (N_12974,N_7516,N_8876);
nand U12975 (N_12975,N_9054,N_6768);
nor U12976 (N_12976,N_5957,N_8874);
and U12977 (N_12977,N_9069,N_6833);
nor U12978 (N_12978,N_5572,N_8272);
nand U12979 (N_12979,N_8475,N_9756);
xor U12980 (N_12980,N_6017,N_9588);
or U12981 (N_12981,N_5540,N_9062);
and U12982 (N_12982,N_9870,N_6164);
xnor U12983 (N_12983,N_8428,N_9437);
or U12984 (N_12984,N_9169,N_6127);
xnor U12985 (N_12985,N_8469,N_6852);
and U12986 (N_12986,N_9881,N_9364);
xnor U12987 (N_12987,N_5212,N_8835);
nand U12988 (N_12988,N_5904,N_6865);
and U12989 (N_12989,N_8657,N_5356);
nand U12990 (N_12990,N_9300,N_7789);
nand U12991 (N_12991,N_6258,N_5458);
nand U12992 (N_12992,N_9170,N_8358);
and U12993 (N_12993,N_7234,N_6714);
xor U12994 (N_12994,N_6223,N_8319);
or U12995 (N_12995,N_6823,N_5931);
nand U12996 (N_12996,N_8059,N_6768);
or U12997 (N_12997,N_8021,N_8449);
xor U12998 (N_12998,N_8351,N_8142);
nor U12999 (N_12999,N_6622,N_7428);
nor U13000 (N_13000,N_8959,N_5980);
or U13001 (N_13001,N_8690,N_5394);
xor U13002 (N_13002,N_6440,N_5361);
nand U13003 (N_13003,N_9017,N_6851);
and U13004 (N_13004,N_8231,N_6197);
and U13005 (N_13005,N_5620,N_7262);
xnor U13006 (N_13006,N_5030,N_6737);
nor U13007 (N_13007,N_9916,N_6123);
nor U13008 (N_13008,N_6868,N_5128);
xnor U13009 (N_13009,N_9734,N_9852);
or U13010 (N_13010,N_5310,N_9809);
nor U13011 (N_13011,N_8212,N_8148);
or U13012 (N_13012,N_5048,N_8149);
and U13013 (N_13013,N_9081,N_9898);
nor U13014 (N_13014,N_9883,N_7970);
nand U13015 (N_13015,N_9463,N_8174);
xor U13016 (N_13016,N_5715,N_6203);
nand U13017 (N_13017,N_7215,N_6423);
xnor U13018 (N_13018,N_7051,N_6878);
xnor U13019 (N_13019,N_7224,N_6920);
and U13020 (N_13020,N_6513,N_8988);
nor U13021 (N_13021,N_7953,N_9739);
or U13022 (N_13022,N_6689,N_7168);
xnor U13023 (N_13023,N_7525,N_6691);
nand U13024 (N_13024,N_8029,N_7062);
xor U13025 (N_13025,N_7081,N_9849);
nand U13026 (N_13026,N_8406,N_9541);
xor U13027 (N_13027,N_8550,N_9142);
nor U13028 (N_13028,N_7167,N_9978);
and U13029 (N_13029,N_9311,N_9951);
xor U13030 (N_13030,N_8462,N_9576);
or U13031 (N_13031,N_7717,N_8759);
xor U13032 (N_13032,N_6363,N_7005);
xnor U13033 (N_13033,N_6181,N_6120);
and U13034 (N_13034,N_5035,N_5034);
nor U13035 (N_13035,N_9591,N_8382);
or U13036 (N_13036,N_9523,N_6694);
nand U13037 (N_13037,N_8402,N_8034);
and U13038 (N_13038,N_8419,N_8534);
nor U13039 (N_13039,N_6630,N_7604);
nor U13040 (N_13040,N_6738,N_7417);
or U13041 (N_13041,N_7232,N_7221);
or U13042 (N_13042,N_9308,N_9981);
nor U13043 (N_13043,N_9911,N_5755);
or U13044 (N_13044,N_9473,N_8201);
nand U13045 (N_13045,N_7880,N_5665);
or U13046 (N_13046,N_7977,N_6423);
or U13047 (N_13047,N_7649,N_5809);
and U13048 (N_13048,N_6402,N_6588);
xnor U13049 (N_13049,N_9783,N_5899);
nand U13050 (N_13050,N_8991,N_8156);
or U13051 (N_13051,N_7339,N_5958);
and U13052 (N_13052,N_5898,N_8131);
or U13053 (N_13053,N_8573,N_5157);
xnor U13054 (N_13054,N_5768,N_7375);
and U13055 (N_13055,N_5243,N_5173);
or U13056 (N_13056,N_5088,N_7671);
or U13057 (N_13057,N_9392,N_8505);
and U13058 (N_13058,N_5882,N_7284);
nor U13059 (N_13059,N_8647,N_8138);
xnor U13060 (N_13060,N_6124,N_7548);
nand U13061 (N_13061,N_8727,N_8577);
nand U13062 (N_13062,N_5722,N_5616);
nor U13063 (N_13063,N_8832,N_7505);
xor U13064 (N_13064,N_8137,N_7327);
nor U13065 (N_13065,N_8166,N_8626);
nand U13066 (N_13066,N_8050,N_6430);
xor U13067 (N_13067,N_9040,N_8650);
xnor U13068 (N_13068,N_5300,N_7951);
xnor U13069 (N_13069,N_6850,N_7659);
nand U13070 (N_13070,N_7492,N_6070);
nor U13071 (N_13071,N_7568,N_5246);
xor U13072 (N_13072,N_8985,N_7983);
xor U13073 (N_13073,N_6890,N_7381);
or U13074 (N_13074,N_5599,N_7268);
xnor U13075 (N_13075,N_6294,N_5391);
nand U13076 (N_13076,N_8224,N_9199);
nand U13077 (N_13077,N_6371,N_5145);
nor U13078 (N_13078,N_6051,N_7005);
and U13079 (N_13079,N_7131,N_7680);
and U13080 (N_13080,N_8750,N_5899);
xor U13081 (N_13081,N_9004,N_9697);
nor U13082 (N_13082,N_7563,N_8700);
nand U13083 (N_13083,N_9231,N_5296);
or U13084 (N_13084,N_7866,N_7451);
nand U13085 (N_13085,N_9213,N_8434);
nor U13086 (N_13086,N_9609,N_7621);
nor U13087 (N_13087,N_8303,N_8715);
nand U13088 (N_13088,N_8006,N_8157);
and U13089 (N_13089,N_7122,N_7881);
or U13090 (N_13090,N_8511,N_6699);
and U13091 (N_13091,N_5052,N_9402);
and U13092 (N_13092,N_6931,N_8808);
nor U13093 (N_13093,N_8431,N_5715);
xnor U13094 (N_13094,N_6678,N_7470);
or U13095 (N_13095,N_5032,N_5727);
nor U13096 (N_13096,N_6058,N_9218);
or U13097 (N_13097,N_5729,N_6311);
or U13098 (N_13098,N_9078,N_7335);
or U13099 (N_13099,N_8197,N_8792);
and U13100 (N_13100,N_5325,N_9162);
and U13101 (N_13101,N_5411,N_8009);
or U13102 (N_13102,N_9500,N_9417);
nor U13103 (N_13103,N_6785,N_6470);
nor U13104 (N_13104,N_5018,N_9650);
nor U13105 (N_13105,N_6718,N_5328);
nor U13106 (N_13106,N_8485,N_8080);
xnor U13107 (N_13107,N_6461,N_9152);
nand U13108 (N_13108,N_5582,N_6514);
nor U13109 (N_13109,N_7654,N_7923);
xnor U13110 (N_13110,N_8162,N_5185);
and U13111 (N_13111,N_5616,N_8888);
and U13112 (N_13112,N_5738,N_5656);
nor U13113 (N_13113,N_5417,N_9521);
or U13114 (N_13114,N_7754,N_6922);
xor U13115 (N_13115,N_9204,N_7952);
and U13116 (N_13116,N_9084,N_6670);
or U13117 (N_13117,N_6109,N_5798);
and U13118 (N_13118,N_8156,N_7283);
or U13119 (N_13119,N_7942,N_7679);
and U13120 (N_13120,N_7802,N_9053);
or U13121 (N_13121,N_7391,N_6312);
xnor U13122 (N_13122,N_7477,N_6757);
nor U13123 (N_13123,N_9353,N_8979);
and U13124 (N_13124,N_7749,N_7720);
nand U13125 (N_13125,N_8916,N_8660);
nand U13126 (N_13126,N_7672,N_8988);
nand U13127 (N_13127,N_8184,N_8316);
nor U13128 (N_13128,N_6303,N_5113);
xor U13129 (N_13129,N_9916,N_7538);
and U13130 (N_13130,N_8972,N_9773);
xor U13131 (N_13131,N_8069,N_6743);
nand U13132 (N_13132,N_8603,N_8027);
nand U13133 (N_13133,N_9280,N_7860);
and U13134 (N_13134,N_7216,N_8531);
or U13135 (N_13135,N_7804,N_6695);
and U13136 (N_13136,N_8454,N_5785);
xnor U13137 (N_13137,N_9517,N_6381);
xnor U13138 (N_13138,N_6485,N_8794);
nor U13139 (N_13139,N_9188,N_8112);
nand U13140 (N_13140,N_5801,N_7246);
xnor U13141 (N_13141,N_9812,N_7863);
and U13142 (N_13142,N_9753,N_9124);
and U13143 (N_13143,N_6178,N_5683);
nand U13144 (N_13144,N_7843,N_5544);
and U13145 (N_13145,N_8315,N_9703);
nor U13146 (N_13146,N_5485,N_6378);
or U13147 (N_13147,N_5036,N_5895);
nor U13148 (N_13148,N_5902,N_5869);
nor U13149 (N_13149,N_9475,N_8630);
xnor U13150 (N_13150,N_9924,N_7866);
nor U13151 (N_13151,N_6274,N_6530);
xor U13152 (N_13152,N_9646,N_5864);
or U13153 (N_13153,N_5577,N_5792);
nand U13154 (N_13154,N_6322,N_6107);
nand U13155 (N_13155,N_8738,N_9177);
and U13156 (N_13156,N_7980,N_8073);
nand U13157 (N_13157,N_8447,N_7772);
nand U13158 (N_13158,N_7250,N_9756);
nor U13159 (N_13159,N_9872,N_9643);
xor U13160 (N_13160,N_7313,N_6737);
nor U13161 (N_13161,N_5198,N_6554);
nand U13162 (N_13162,N_5724,N_8669);
and U13163 (N_13163,N_6614,N_5650);
or U13164 (N_13164,N_6433,N_7968);
nor U13165 (N_13165,N_9297,N_6352);
nand U13166 (N_13166,N_6672,N_7758);
or U13167 (N_13167,N_8980,N_7181);
or U13168 (N_13168,N_8760,N_6134);
nor U13169 (N_13169,N_5732,N_6162);
or U13170 (N_13170,N_9540,N_8233);
xor U13171 (N_13171,N_6852,N_7460);
and U13172 (N_13172,N_5523,N_8371);
and U13173 (N_13173,N_6883,N_9477);
and U13174 (N_13174,N_6833,N_5976);
nand U13175 (N_13175,N_6642,N_5207);
nor U13176 (N_13176,N_5090,N_7853);
nor U13177 (N_13177,N_9052,N_9143);
nand U13178 (N_13178,N_8855,N_9222);
and U13179 (N_13179,N_9500,N_5528);
nand U13180 (N_13180,N_8930,N_5795);
nand U13181 (N_13181,N_7157,N_8614);
xnor U13182 (N_13182,N_7859,N_6507);
or U13183 (N_13183,N_8596,N_7231);
or U13184 (N_13184,N_7082,N_5815);
and U13185 (N_13185,N_6100,N_5965);
and U13186 (N_13186,N_9091,N_5140);
and U13187 (N_13187,N_5153,N_8580);
nand U13188 (N_13188,N_8579,N_6327);
nor U13189 (N_13189,N_9363,N_7102);
or U13190 (N_13190,N_6718,N_6276);
or U13191 (N_13191,N_7321,N_6966);
nand U13192 (N_13192,N_9160,N_5981);
nor U13193 (N_13193,N_6988,N_6849);
and U13194 (N_13194,N_7759,N_6143);
xor U13195 (N_13195,N_8400,N_5080);
or U13196 (N_13196,N_9699,N_9501);
nor U13197 (N_13197,N_6849,N_7113);
nor U13198 (N_13198,N_5473,N_5451);
or U13199 (N_13199,N_6222,N_9191);
nand U13200 (N_13200,N_7882,N_9945);
nand U13201 (N_13201,N_9836,N_8894);
nor U13202 (N_13202,N_8982,N_6527);
nor U13203 (N_13203,N_5899,N_8706);
nor U13204 (N_13204,N_5159,N_9203);
xnor U13205 (N_13205,N_6827,N_5227);
xor U13206 (N_13206,N_8578,N_8121);
nor U13207 (N_13207,N_8454,N_8998);
nor U13208 (N_13208,N_8023,N_6467);
xnor U13209 (N_13209,N_8288,N_6280);
nor U13210 (N_13210,N_6744,N_8441);
xnor U13211 (N_13211,N_8703,N_5703);
xor U13212 (N_13212,N_5736,N_7651);
nor U13213 (N_13213,N_8889,N_9568);
or U13214 (N_13214,N_7907,N_9886);
or U13215 (N_13215,N_7797,N_5865);
xor U13216 (N_13216,N_7464,N_7764);
nand U13217 (N_13217,N_7325,N_9149);
xnor U13218 (N_13218,N_8227,N_9889);
nand U13219 (N_13219,N_6955,N_7634);
nand U13220 (N_13220,N_6036,N_7577);
and U13221 (N_13221,N_7165,N_6568);
or U13222 (N_13222,N_6285,N_5837);
and U13223 (N_13223,N_6351,N_9272);
and U13224 (N_13224,N_9973,N_8501);
nor U13225 (N_13225,N_7781,N_6045);
nand U13226 (N_13226,N_9985,N_6337);
nand U13227 (N_13227,N_5330,N_9305);
nand U13228 (N_13228,N_5123,N_9520);
xnor U13229 (N_13229,N_5644,N_9001);
xnor U13230 (N_13230,N_5973,N_7718);
nor U13231 (N_13231,N_8041,N_5440);
and U13232 (N_13232,N_6384,N_6445);
nand U13233 (N_13233,N_6308,N_6651);
and U13234 (N_13234,N_5116,N_6715);
nand U13235 (N_13235,N_6221,N_5067);
and U13236 (N_13236,N_9096,N_9385);
nand U13237 (N_13237,N_8078,N_7614);
xnor U13238 (N_13238,N_6861,N_6474);
xnor U13239 (N_13239,N_5979,N_6130);
xor U13240 (N_13240,N_8021,N_7128);
xnor U13241 (N_13241,N_5586,N_9457);
xor U13242 (N_13242,N_7655,N_6241);
and U13243 (N_13243,N_7000,N_7071);
xnor U13244 (N_13244,N_5576,N_6238);
and U13245 (N_13245,N_7948,N_7153);
nand U13246 (N_13246,N_8444,N_8520);
nor U13247 (N_13247,N_9214,N_5471);
or U13248 (N_13248,N_5278,N_9483);
nor U13249 (N_13249,N_6835,N_5929);
nor U13250 (N_13250,N_8588,N_6837);
and U13251 (N_13251,N_9945,N_5802);
or U13252 (N_13252,N_7161,N_5751);
nand U13253 (N_13253,N_9103,N_8357);
xor U13254 (N_13254,N_8617,N_9781);
xnor U13255 (N_13255,N_6627,N_6112);
and U13256 (N_13256,N_7431,N_6598);
and U13257 (N_13257,N_6289,N_5882);
or U13258 (N_13258,N_9617,N_7901);
nor U13259 (N_13259,N_8740,N_9986);
and U13260 (N_13260,N_6853,N_5314);
nor U13261 (N_13261,N_6940,N_6747);
and U13262 (N_13262,N_6137,N_6735);
xor U13263 (N_13263,N_6573,N_6047);
nor U13264 (N_13264,N_6350,N_7606);
nand U13265 (N_13265,N_8356,N_8615);
and U13266 (N_13266,N_9111,N_9656);
or U13267 (N_13267,N_8420,N_5307);
and U13268 (N_13268,N_5075,N_6786);
nand U13269 (N_13269,N_5698,N_7840);
or U13270 (N_13270,N_7817,N_9300);
or U13271 (N_13271,N_6647,N_6033);
or U13272 (N_13272,N_9593,N_7008);
or U13273 (N_13273,N_5942,N_6651);
or U13274 (N_13274,N_8777,N_6212);
nand U13275 (N_13275,N_7883,N_8923);
xor U13276 (N_13276,N_5374,N_9327);
or U13277 (N_13277,N_7554,N_8155);
nand U13278 (N_13278,N_7298,N_8122);
xnor U13279 (N_13279,N_6142,N_8339);
xnor U13280 (N_13280,N_9765,N_5500);
nand U13281 (N_13281,N_7869,N_8834);
xor U13282 (N_13282,N_5911,N_6663);
or U13283 (N_13283,N_8488,N_9833);
xor U13284 (N_13284,N_6433,N_5403);
or U13285 (N_13285,N_7738,N_9880);
nand U13286 (N_13286,N_5718,N_5102);
and U13287 (N_13287,N_5593,N_9264);
or U13288 (N_13288,N_8525,N_9307);
nand U13289 (N_13289,N_5166,N_6911);
or U13290 (N_13290,N_6582,N_7311);
nand U13291 (N_13291,N_6519,N_9139);
nand U13292 (N_13292,N_9246,N_6081);
xnor U13293 (N_13293,N_8335,N_6961);
xor U13294 (N_13294,N_8786,N_9026);
or U13295 (N_13295,N_7220,N_7775);
and U13296 (N_13296,N_7149,N_7049);
xnor U13297 (N_13297,N_6056,N_8285);
nand U13298 (N_13298,N_8361,N_5772);
or U13299 (N_13299,N_6250,N_9411);
nor U13300 (N_13300,N_5456,N_5345);
nor U13301 (N_13301,N_9317,N_7649);
and U13302 (N_13302,N_7702,N_5513);
nand U13303 (N_13303,N_6514,N_9615);
and U13304 (N_13304,N_5634,N_5224);
and U13305 (N_13305,N_9424,N_5363);
nor U13306 (N_13306,N_9724,N_7204);
nor U13307 (N_13307,N_8718,N_5140);
xnor U13308 (N_13308,N_9417,N_6725);
xnor U13309 (N_13309,N_8480,N_8353);
xnor U13310 (N_13310,N_7847,N_9612);
nor U13311 (N_13311,N_9638,N_7049);
nand U13312 (N_13312,N_7276,N_5421);
or U13313 (N_13313,N_9951,N_8738);
nor U13314 (N_13314,N_9904,N_5721);
and U13315 (N_13315,N_6732,N_8024);
and U13316 (N_13316,N_7778,N_8640);
nand U13317 (N_13317,N_9810,N_8930);
and U13318 (N_13318,N_6938,N_9034);
and U13319 (N_13319,N_8462,N_5799);
or U13320 (N_13320,N_5994,N_5009);
and U13321 (N_13321,N_7862,N_8663);
and U13322 (N_13322,N_6091,N_9686);
nand U13323 (N_13323,N_7932,N_7761);
nand U13324 (N_13324,N_5588,N_8122);
nor U13325 (N_13325,N_5778,N_6995);
and U13326 (N_13326,N_7298,N_9849);
and U13327 (N_13327,N_5800,N_8217);
nand U13328 (N_13328,N_7475,N_8650);
and U13329 (N_13329,N_6642,N_6823);
nor U13330 (N_13330,N_8690,N_7053);
nand U13331 (N_13331,N_9128,N_6014);
or U13332 (N_13332,N_7925,N_9600);
nand U13333 (N_13333,N_5062,N_5497);
or U13334 (N_13334,N_7120,N_8967);
nand U13335 (N_13335,N_7519,N_7701);
or U13336 (N_13336,N_7489,N_5349);
nand U13337 (N_13337,N_5985,N_9542);
nor U13338 (N_13338,N_6782,N_6282);
nor U13339 (N_13339,N_9184,N_6810);
or U13340 (N_13340,N_6845,N_6864);
xnor U13341 (N_13341,N_7709,N_8314);
and U13342 (N_13342,N_5112,N_6237);
xor U13343 (N_13343,N_7786,N_9389);
nor U13344 (N_13344,N_8935,N_8776);
nand U13345 (N_13345,N_5879,N_6226);
or U13346 (N_13346,N_9743,N_5547);
nor U13347 (N_13347,N_9501,N_9308);
nor U13348 (N_13348,N_6206,N_5044);
nand U13349 (N_13349,N_6600,N_5914);
or U13350 (N_13350,N_5173,N_9714);
xnor U13351 (N_13351,N_8006,N_7469);
or U13352 (N_13352,N_5591,N_7911);
nand U13353 (N_13353,N_9765,N_9262);
xnor U13354 (N_13354,N_8218,N_9613);
or U13355 (N_13355,N_7304,N_6933);
or U13356 (N_13356,N_9261,N_5866);
nor U13357 (N_13357,N_6258,N_8611);
or U13358 (N_13358,N_8359,N_8699);
and U13359 (N_13359,N_9919,N_6203);
nor U13360 (N_13360,N_7864,N_8854);
nor U13361 (N_13361,N_9949,N_7261);
nor U13362 (N_13362,N_8888,N_5675);
nand U13363 (N_13363,N_5499,N_8266);
or U13364 (N_13364,N_7515,N_6286);
and U13365 (N_13365,N_9130,N_7895);
nand U13366 (N_13366,N_6329,N_8300);
xor U13367 (N_13367,N_8906,N_9454);
and U13368 (N_13368,N_8709,N_7037);
and U13369 (N_13369,N_8313,N_8208);
xnor U13370 (N_13370,N_7252,N_8449);
xor U13371 (N_13371,N_8768,N_7278);
nor U13372 (N_13372,N_5916,N_5097);
nor U13373 (N_13373,N_6522,N_5473);
xor U13374 (N_13374,N_8541,N_8623);
nand U13375 (N_13375,N_8213,N_9519);
and U13376 (N_13376,N_6655,N_9387);
and U13377 (N_13377,N_8348,N_8609);
nand U13378 (N_13378,N_8672,N_5083);
nor U13379 (N_13379,N_6366,N_6611);
nand U13380 (N_13380,N_9086,N_9779);
or U13381 (N_13381,N_7031,N_8808);
nand U13382 (N_13382,N_7735,N_5313);
xor U13383 (N_13383,N_9274,N_7845);
nor U13384 (N_13384,N_7040,N_8927);
xnor U13385 (N_13385,N_5052,N_7349);
and U13386 (N_13386,N_6331,N_5404);
nand U13387 (N_13387,N_8606,N_9814);
and U13388 (N_13388,N_9638,N_7909);
nand U13389 (N_13389,N_9081,N_5719);
nor U13390 (N_13390,N_9408,N_8964);
or U13391 (N_13391,N_7329,N_9231);
nand U13392 (N_13392,N_9285,N_9635);
nand U13393 (N_13393,N_5694,N_5125);
nor U13394 (N_13394,N_8684,N_6241);
and U13395 (N_13395,N_8275,N_8174);
nand U13396 (N_13396,N_8789,N_8480);
nor U13397 (N_13397,N_8830,N_8469);
nand U13398 (N_13398,N_6239,N_6644);
nand U13399 (N_13399,N_9252,N_5412);
and U13400 (N_13400,N_9573,N_9929);
and U13401 (N_13401,N_8264,N_5859);
or U13402 (N_13402,N_9151,N_9753);
nand U13403 (N_13403,N_5600,N_8692);
nand U13404 (N_13404,N_9103,N_5954);
nor U13405 (N_13405,N_6637,N_9310);
and U13406 (N_13406,N_9026,N_6109);
and U13407 (N_13407,N_6901,N_8041);
nor U13408 (N_13408,N_6209,N_8817);
xnor U13409 (N_13409,N_8198,N_7629);
nor U13410 (N_13410,N_7581,N_8577);
and U13411 (N_13411,N_6434,N_7346);
or U13412 (N_13412,N_7919,N_6703);
nor U13413 (N_13413,N_5482,N_5478);
or U13414 (N_13414,N_9062,N_8043);
xnor U13415 (N_13415,N_6169,N_9110);
nand U13416 (N_13416,N_8346,N_6488);
xor U13417 (N_13417,N_5535,N_8427);
nand U13418 (N_13418,N_7387,N_5697);
nand U13419 (N_13419,N_6870,N_5071);
xor U13420 (N_13420,N_8470,N_7859);
nand U13421 (N_13421,N_8707,N_8593);
nor U13422 (N_13422,N_9858,N_5232);
nor U13423 (N_13423,N_6307,N_8037);
nand U13424 (N_13424,N_9482,N_9430);
xnor U13425 (N_13425,N_5753,N_6427);
or U13426 (N_13426,N_8508,N_8628);
and U13427 (N_13427,N_5186,N_8595);
xnor U13428 (N_13428,N_5176,N_7072);
nand U13429 (N_13429,N_5103,N_5963);
xor U13430 (N_13430,N_8463,N_7839);
nand U13431 (N_13431,N_7855,N_6509);
and U13432 (N_13432,N_6296,N_6114);
xnor U13433 (N_13433,N_8874,N_6961);
nor U13434 (N_13434,N_7524,N_9184);
nor U13435 (N_13435,N_5033,N_9586);
xnor U13436 (N_13436,N_9073,N_9812);
nor U13437 (N_13437,N_8871,N_8358);
or U13438 (N_13438,N_5462,N_7848);
nand U13439 (N_13439,N_7091,N_8236);
nand U13440 (N_13440,N_8038,N_5173);
nor U13441 (N_13441,N_8530,N_8984);
and U13442 (N_13442,N_7286,N_7933);
or U13443 (N_13443,N_9967,N_9383);
nand U13444 (N_13444,N_9659,N_8232);
xor U13445 (N_13445,N_5981,N_8532);
nor U13446 (N_13446,N_8269,N_7243);
and U13447 (N_13447,N_6752,N_7682);
or U13448 (N_13448,N_5988,N_5208);
or U13449 (N_13449,N_7529,N_8353);
xor U13450 (N_13450,N_7105,N_5983);
and U13451 (N_13451,N_5241,N_6074);
or U13452 (N_13452,N_7667,N_7250);
xnor U13453 (N_13453,N_8226,N_5162);
nor U13454 (N_13454,N_8820,N_8200);
xor U13455 (N_13455,N_7084,N_7844);
xor U13456 (N_13456,N_8045,N_8497);
and U13457 (N_13457,N_9999,N_5511);
nand U13458 (N_13458,N_7261,N_5359);
nor U13459 (N_13459,N_6716,N_5223);
and U13460 (N_13460,N_7957,N_7231);
xnor U13461 (N_13461,N_9145,N_6575);
nand U13462 (N_13462,N_7783,N_9499);
xnor U13463 (N_13463,N_5900,N_8164);
or U13464 (N_13464,N_9648,N_5580);
or U13465 (N_13465,N_6125,N_5712);
nand U13466 (N_13466,N_6892,N_9548);
nor U13467 (N_13467,N_5076,N_7295);
nor U13468 (N_13468,N_8981,N_7014);
and U13469 (N_13469,N_8009,N_9637);
nand U13470 (N_13470,N_9146,N_9277);
and U13471 (N_13471,N_7855,N_9124);
nor U13472 (N_13472,N_9037,N_9216);
nor U13473 (N_13473,N_9463,N_5502);
nand U13474 (N_13474,N_6541,N_6373);
or U13475 (N_13475,N_8976,N_6206);
xnor U13476 (N_13476,N_5179,N_8577);
xnor U13477 (N_13477,N_9589,N_8026);
nor U13478 (N_13478,N_5117,N_6803);
and U13479 (N_13479,N_5598,N_7264);
nor U13480 (N_13480,N_8720,N_7254);
xor U13481 (N_13481,N_7588,N_9991);
and U13482 (N_13482,N_6510,N_6604);
xnor U13483 (N_13483,N_9875,N_8914);
and U13484 (N_13484,N_5010,N_5348);
nand U13485 (N_13485,N_5107,N_6380);
nand U13486 (N_13486,N_5569,N_5078);
nor U13487 (N_13487,N_7483,N_7366);
and U13488 (N_13488,N_7211,N_5765);
nand U13489 (N_13489,N_8799,N_6674);
and U13490 (N_13490,N_9481,N_6960);
nand U13491 (N_13491,N_6109,N_5257);
and U13492 (N_13492,N_7195,N_7731);
and U13493 (N_13493,N_8408,N_7539);
xnor U13494 (N_13494,N_8758,N_9313);
and U13495 (N_13495,N_8382,N_9401);
nor U13496 (N_13496,N_8530,N_9197);
xnor U13497 (N_13497,N_5459,N_8025);
or U13498 (N_13498,N_7295,N_6359);
nor U13499 (N_13499,N_7622,N_5093);
and U13500 (N_13500,N_8859,N_7157);
and U13501 (N_13501,N_6187,N_5223);
and U13502 (N_13502,N_5856,N_7531);
and U13503 (N_13503,N_7176,N_8448);
or U13504 (N_13504,N_6971,N_8505);
xor U13505 (N_13505,N_9007,N_6949);
nor U13506 (N_13506,N_7541,N_6108);
nand U13507 (N_13507,N_9687,N_7780);
nor U13508 (N_13508,N_8158,N_7867);
and U13509 (N_13509,N_8196,N_5588);
or U13510 (N_13510,N_6251,N_7858);
nand U13511 (N_13511,N_9174,N_5371);
or U13512 (N_13512,N_7450,N_9833);
xor U13513 (N_13513,N_8247,N_7650);
and U13514 (N_13514,N_9663,N_8360);
and U13515 (N_13515,N_7761,N_5940);
or U13516 (N_13516,N_6595,N_9984);
nor U13517 (N_13517,N_5202,N_8556);
nand U13518 (N_13518,N_9246,N_7795);
xor U13519 (N_13519,N_9821,N_6236);
nand U13520 (N_13520,N_7850,N_7863);
and U13521 (N_13521,N_6285,N_5192);
or U13522 (N_13522,N_8697,N_5723);
or U13523 (N_13523,N_8301,N_8186);
and U13524 (N_13524,N_5335,N_5640);
or U13525 (N_13525,N_8558,N_8368);
xor U13526 (N_13526,N_8335,N_9000);
xnor U13527 (N_13527,N_9339,N_9668);
or U13528 (N_13528,N_6570,N_5654);
and U13529 (N_13529,N_8947,N_9709);
and U13530 (N_13530,N_9615,N_8462);
xnor U13531 (N_13531,N_6299,N_5438);
nor U13532 (N_13532,N_7992,N_9218);
xnor U13533 (N_13533,N_8270,N_7456);
and U13534 (N_13534,N_5941,N_5224);
nor U13535 (N_13535,N_9630,N_9289);
and U13536 (N_13536,N_5173,N_9861);
xor U13537 (N_13537,N_7795,N_7775);
xor U13538 (N_13538,N_7139,N_6752);
and U13539 (N_13539,N_7435,N_6805);
or U13540 (N_13540,N_5220,N_8039);
xor U13541 (N_13541,N_8354,N_7890);
xor U13542 (N_13542,N_9062,N_7656);
nand U13543 (N_13543,N_7545,N_5453);
nor U13544 (N_13544,N_9750,N_9002);
and U13545 (N_13545,N_9055,N_9292);
and U13546 (N_13546,N_6255,N_5173);
nand U13547 (N_13547,N_8574,N_5902);
nor U13548 (N_13548,N_5349,N_6450);
xor U13549 (N_13549,N_5889,N_8713);
nor U13550 (N_13550,N_6180,N_5542);
xor U13551 (N_13551,N_5775,N_5370);
nor U13552 (N_13552,N_6917,N_7769);
and U13553 (N_13553,N_5422,N_9876);
nand U13554 (N_13554,N_7920,N_9097);
nor U13555 (N_13555,N_5898,N_6021);
nor U13556 (N_13556,N_8132,N_6149);
and U13557 (N_13557,N_7460,N_5440);
xor U13558 (N_13558,N_8356,N_7972);
nor U13559 (N_13559,N_7341,N_7051);
and U13560 (N_13560,N_5840,N_7911);
and U13561 (N_13561,N_5075,N_7882);
xnor U13562 (N_13562,N_6769,N_7166);
or U13563 (N_13563,N_8606,N_5647);
xnor U13564 (N_13564,N_6699,N_9641);
or U13565 (N_13565,N_9606,N_5935);
nand U13566 (N_13566,N_6591,N_6721);
xor U13567 (N_13567,N_8453,N_9033);
nand U13568 (N_13568,N_5095,N_8933);
or U13569 (N_13569,N_5552,N_6524);
xor U13570 (N_13570,N_5382,N_5668);
or U13571 (N_13571,N_7414,N_8763);
nand U13572 (N_13572,N_9865,N_5321);
nor U13573 (N_13573,N_6073,N_5172);
nor U13574 (N_13574,N_6413,N_6085);
nand U13575 (N_13575,N_6922,N_6770);
nor U13576 (N_13576,N_6422,N_8982);
or U13577 (N_13577,N_9344,N_6578);
and U13578 (N_13578,N_6132,N_7588);
nor U13579 (N_13579,N_8524,N_9824);
nor U13580 (N_13580,N_9660,N_8834);
xor U13581 (N_13581,N_8793,N_7619);
nor U13582 (N_13582,N_5191,N_7840);
or U13583 (N_13583,N_6982,N_6699);
or U13584 (N_13584,N_7760,N_7936);
nand U13585 (N_13585,N_8649,N_8961);
nand U13586 (N_13586,N_5349,N_6668);
nor U13587 (N_13587,N_9132,N_6333);
nand U13588 (N_13588,N_8576,N_5639);
or U13589 (N_13589,N_7835,N_6023);
and U13590 (N_13590,N_9425,N_8411);
nand U13591 (N_13591,N_6795,N_9363);
nand U13592 (N_13592,N_6079,N_8499);
or U13593 (N_13593,N_5090,N_6981);
nand U13594 (N_13594,N_6305,N_8814);
xnor U13595 (N_13595,N_7393,N_6424);
and U13596 (N_13596,N_6187,N_5835);
or U13597 (N_13597,N_5737,N_9953);
nand U13598 (N_13598,N_7850,N_8784);
xor U13599 (N_13599,N_5440,N_7347);
nor U13600 (N_13600,N_6083,N_9427);
and U13601 (N_13601,N_9041,N_9951);
or U13602 (N_13602,N_9550,N_6140);
nand U13603 (N_13603,N_8116,N_9534);
nand U13604 (N_13604,N_8207,N_7339);
xor U13605 (N_13605,N_5803,N_7853);
and U13606 (N_13606,N_9652,N_7804);
nor U13607 (N_13607,N_7661,N_7560);
nor U13608 (N_13608,N_9673,N_6493);
nor U13609 (N_13609,N_7040,N_8009);
or U13610 (N_13610,N_9609,N_8376);
xor U13611 (N_13611,N_9694,N_9596);
nand U13612 (N_13612,N_9539,N_7188);
and U13613 (N_13613,N_7245,N_9569);
nor U13614 (N_13614,N_5226,N_8190);
nor U13615 (N_13615,N_7140,N_9382);
nand U13616 (N_13616,N_9009,N_9633);
or U13617 (N_13617,N_9103,N_9305);
xor U13618 (N_13618,N_8598,N_6919);
nand U13619 (N_13619,N_8923,N_7902);
nand U13620 (N_13620,N_8176,N_5649);
and U13621 (N_13621,N_9421,N_6252);
xor U13622 (N_13622,N_6332,N_7875);
or U13623 (N_13623,N_7121,N_6236);
nor U13624 (N_13624,N_5022,N_8734);
or U13625 (N_13625,N_9710,N_9581);
or U13626 (N_13626,N_5223,N_6009);
or U13627 (N_13627,N_8638,N_9089);
xor U13628 (N_13628,N_9988,N_8262);
and U13629 (N_13629,N_9361,N_6550);
nand U13630 (N_13630,N_8783,N_7223);
nor U13631 (N_13631,N_8760,N_8174);
or U13632 (N_13632,N_7360,N_9264);
nand U13633 (N_13633,N_6846,N_9306);
or U13634 (N_13634,N_7643,N_9587);
or U13635 (N_13635,N_9551,N_9941);
nand U13636 (N_13636,N_5680,N_7271);
and U13637 (N_13637,N_6948,N_8870);
or U13638 (N_13638,N_6807,N_8697);
nand U13639 (N_13639,N_7857,N_8531);
xnor U13640 (N_13640,N_5093,N_7386);
and U13641 (N_13641,N_8314,N_5722);
or U13642 (N_13642,N_6569,N_7029);
or U13643 (N_13643,N_5946,N_7483);
and U13644 (N_13644,N_8745,N_6702);
xor U13645 (N_13645,N_9226,N_5350);
nand U13646 (N_13646,N_6546,N_5126);
or U13647 (N_13647,N_7404,N_7250);
nand U13648 (N_13648,N_5132,N_9901);
nand U13649 (N_13649,N_9522,N_6191);
nand U13650 (N_13650,N_5789,N_9908);
and U13651 (N_13651,N_5648,N_6297);
xnor U13652 (N_13652,N_5585,N_7353);
and U13653 (N_13653,N_7587,N_7736);
and U13654 (N_13654,N_7279,N_9413);
or U13655 (N_13655,N_8373,N_5048);
and U13656 (N_13656,N_9268,N_5573);
xor U13657 (N_13657,N_5314,N_8723);
or U13658 (N_13658,N_6732,N_8410);
nor U13659 (N_13659,N_9325,N_8997);
nor U13660 (N_13660,N_6119,N_7504);
or U13661 (N_13661,N_5675,N_9005);
nand U13662 (N_13662,N_7492,N_7810);
and U13663 (N_13663,N_9495,N_9393);
nand U13664 (N_13664,N_8251,N_7644);
nor U13665 (N_13665,N_6018,N_9360);
nor U13666 (N_13666,N_8964,N_8746);
and U13667 (N_13667,N_9580,N_5522);
or U13668 (N_13668,N_8127,N_6982);
nand U13669 (N_13669,N_5920,N_8076);
nor U13670 (N_13670,N_6420,N_9384);
nor U13671 (N_13671,N_5957,N_7518);
and U13672 (N_13672,N_5803,N_9939);
nand U13673 (N_13673,N_6830,N_5574);
and U13674 (N_13674,N_8697,N_9191);
nand U13675 (N_13675,N_9526,N_9202);
or U13676 (N_13676,N_9131,N_8643);
or U13677 (N_13677,N_7767,N_9645);
nand U13678 (N_13678,N_9968,N_5216);
xnor U13679 (N_13679,N_7121,N_5979);
nor U13680 (N_13680,N_9175,N_5674);
xnor U13681 (N_13681,N_7167,N_9246);
xnor U13682 (N_13682,N_6544,N_7347);
nand U13683 (N_13683,N_8831,N_9559);
or U13684 (N_13684,N_6076,N_5708);
and U13685 (N_13685,N_7011,N_8344);
xor U13686 (N_13686,N_9800,N_7484);
xnor U13687 (N_13687,N_8667,N_9629);
xor U13688 (N_13688,N_6875,N_6197);
nor U13689 (N_13689,N_6739,N_5839);
and U13690 (N_13690,N_9772,N_8708);
nand U13691 (N_13691,N_7067,N_7187);
or U13692 (N_13692,N_6462,N_6594);
nor U13693 (N_13693,N_6744,N_7633);
nor U13694 (N_13694,N_6270,N_7518);
nand U13695 (N_13695,N_9523,N_7295);
or U13696 (N_13696,N_7269,N_8260);
and U13697 (N_13697,N_6621,N_5048);
and U13698 (N_13698,N_7542,N_9738);
or U13699 (N_13699,N_9201,N_5879);
and U13700 (N_13700,N_9094,N_9582);
and U13701 (N_13701,N_5561,N_6360);
or U13702 (N_13702,N_8694,N_6224);
or U13703 (N_13703,N_9802,N_6375);
or U13704 (N_13704,N_6421,N_7112);
xor U13705 (N_13705,N_9631,N_8246);
and U13706 (N_13706,N_9536,N_5375);
or U13707 (N_13707,N_6272,N_6838);
nand U13708 (N_13708,N_7321,N_6821);
and U13709 (N_13709,N_5112,N_5731);
nand U13710 (N_13710,N_6344,N_7739);
xor U13711 (N_13711,N_5650,N_5514);
nand U13712 (N_13712,N_8358,N_9324);
and U13713 (N_13713,N_6786,N_9331);
nand U13714 (N_13714,N_9030,N_6182);
nor U13715 (N_13715,N_6867,N_7893);
xor U13716 (N_13716,N_5628,N_9766);
nor U13717 (N_13717,N_9961,N_8839);
or U13718 (N_13718,N_5433,N_9795);
or U13719 (N_13719,N_6889,N_9751);
nor U13720 (N_13720,N_6012,N_7027);
or U13721 (N_13721,N_6300,N_8978);
or U13722 (N_13722,N_5101,N_5666);
nor U13723 (N_13723,N_9237,N_5013);
nand U13724 (N_13724,N_8887,N_8471);
xnor U13725 (N_13725,N_8518,N_7086);
or U13726 (N_13726,N_7578,N_5816);
nand U13727 (N_13727,N_6429,N_6018);
nand U13728 (N_13728,N_8417,N_9349);
nor U13729 (N_13729,N_7626,N_8719);
xor U13730 (N_13730,N_5332,N_6004);
xnor U13731 (N_13731,N_9909,N_7645);
nand U13732 (N_13732,N_9392,N_7752);
nor U13733 (N_13733,N_7297,N_8891);
or U13734 (N_13734,N_9522,N_7617);
or U13735 (N_13735,N_8060,N_8552);
and U13736 (N_13736,N_8819,N_6448);
and U13737 (N_13737,N_9030,N_8698);
or U13738 (N_13738,N_8418,N_5650);
xnor U13739 (N_13739,N_8112,N_8446);
nand U13740 (N_13740,N_8500,N_5556);
and U13741 (N_13741,N_6492,N_7003);
nand U13742 (N_13742,N_9123,N_8012);
nand U13743 (N_13743,N_9425,N_8863);
nand U13744 (N_13744,N_5881,N_6189);
or U13745 (N_13745,N_7562,N_6347);
and U13746 (N_13746,N_6247,N_9651);
nor U13747 (N_13747,N_5808,N_9614);
xnor U13748 (N_13748,N_9359,N_5358);
xor U13749 (N_13749,N_6461,N_7298);
nor U13750 (N_13750,N_8003,N_7749);
and U13751 (N_13751,N_8062,N_8471);
xnor U13752 (N_13752,N_9229,N_9251);
and U13753 (N_13753,N_6544,N_8736);
xor U13754 (N_13754,N_8003,N_5345);
nand U13755 (N_13755,N_9731,N_6179);
and U13756 (N_13756,N_5793,N_9651);
or U13757 (N_13757,N_5163,N_7126);
xor U13758 (N_13758,N_9564,N_7630);
and U13759 (N_13759,N_8948,N_6471);
and U13760 (N_13760,N_9577,N_7810);
nor U13761 (N_13761,N_9837,N_5867);
nand U13762 (N_13762,N_8475,N_8367);
nor U13763 (N_13763,N_8457,N_8262);
or U13764 (N_13764,N_5042,N_6175);
and U13765 (N_13765,N_8480,N_5483);
xor U13766 (N_13766,N_6676,N_8116);
nor U13767 (N_13767,N_8125,N_5474);
nand U13768 (N_13768,N_9629,N_5157);
nor U13769 (N_13769,N_9315,N_9592);
or U13770 (N_13770,N_5829,N_7493);
and U13771 (N_13771,N_5024,N_6515);
and U13772 (N_13772,N_9892,N_8290);
and U13773 (N_13773,N_6433,N_8402);
or U13774 (N_13774,N_5245,N_8017);
xor U13775 (N_13775,N_7683,N_5102);
and U13776 (N_13776,N_6516,N_7246);
nor U13777 (N_13777,N_8134,N_8082);
or U13778 (N_13778,N_7925,N_9554);
or U13779 (N_13779,N_8582,N_9064);
nor U13780 (N_13780,N_6868,N_6472);
nor U13781 (N_13781,N_7129,N_6276);
nor U13782 (N_13782,N_6804,N_8105);
or U13783 (N_13783,N_9228,N_5870);
nand U13784 (N_13784,N_7129,N_6884);
or U13785 (N_13785,N_8330,N_9796);
xnor U13786 (N_13786,N_7830,N_9953);
or U13787 (N_13787,N_7420,N_7696);
nor U13788 (N_13788,N_8684,N_7273);
or U13789 (N_13789,N_5832,N_6869);
or U13790 (N_13790,N_8672,N_9340);
or U13791 (N_13791,N_6159,N_5124);
nand U13792 (N_13792,N_8571,N_7597);
or U13793 (N_13793,N_7923,N_7075);
xnor U13794 (N_13794,N_9398,N_8440);
nand U13795 (N_13795,N_5249,N_6624);
or U13796 (N_13796,N_7804,N_5874);
and U13797 (N_13797,N_7120,N_5364);
nor U13798 (N_13798,N_8927,N_7858);
nand U13799 (N_13799,N_5833,N_7727);
xnor U13800 (N_13800,N_5112,N_6450);
nand U13801 (N_13801,N_6903,N_6777);
nor U13802 (N_13802,N_5582,N_7209);
and U13803 (N_13803,N_6875,N_8250);
and U13804 (N_13804,N_9532,N_8347);
and U13805 (N_13805,N_6282,N_6467);
nor U13806 (N_13806,N_8105,N_7396);
and U13807 (N_13807,N_8120,N_7557);
and U13808 (N_13808,N_7726,N_7932);
xor U13809 (N_13809,N_9690,N_8107);
and U13810 (N_13810,N_6102,N_9897);
nand U13811 (N_13811,N_5049,N_6875);
and U13812 (N_13812,N_6591,N_5218);
nor U13813 (N_13813,N_7953,N_7615);
and U13814 (N_13814,N_8308,N_7869);
nor U13815 (N_13815,N_7119,N_8683);
and U13816 (N_13816,N_7878,N_6610);
or U13817 (N_13817,N_9698,N_8678);
or U13818 (N_13818,N_8878,N_7283);
or U13819 (N_13819,N_6482,N_5827);
or U13820 (N_13820,N_7774,N_7192);
nand U13821 (N_13821,N_5643,N_8135);
nand U13822 (N_13822,N_5867,N_6263);
xnor U13823 (N_13823,N_7165,N_5841);
or U13824 (N_13824,N_8298,N_8402);
nor U13825 (N_13825,N_6142,N_7765);
nand U13826 (N_13826,N_6737,N_8620);
nand U13827 (N_13827,N_5100,N_7307);
nor U13828 (N_13828,N_6388,N_5499);
nor U13829 (N_13829,N_9173,N_6244);
and U13830 (N_13830,N_6562,N_7968);
or U13831 (N_13831,N_9165,N_5925);
and U13832 (N_13832,N_6501,N_9297);
and U13833 (N_13833,N_6165,N_9155);
nor U13834 (N_13834,N_9682,N_7518);
nand U13835 (N_13835,N_7287,N_9860);
nor U13836 (N_13836,N_5471,N_8350);
and U13837 (N_13837,N_6317,N_8812);
nand U13838 (N_13838,N_5410,N_5442);
nand U13839 (N_13839,N_8716,N_9276);
nand U13840 (N_13840,N_7298,N_7767);
nor U13841 (N_13841,N_6223,N_6028);
or U13842 (N_13842,N_8449,N_5390);
nor U13843 (N_13843,N_7597,N_9190);
and U13844 (N_13844,N_8521,N_7856);
nor U13845 (N_13845,N_5897,N_9631);
and U13846 (N_13846,N_9905,N_9442);
xnor U13847 (N_13847,N_7848,N_8041);
and U13848 (N_13848,N_5807,N_9373);
xnor U13849 (N_13849,N_7518,N_5218);
xnor U13850 (N_13850,N_5375,N_5953);
nand U13851 (N_13851,N_5524,N_8797);
or U13852 (N_13852,N_6497,N_5092);
nand U13853 (N_13853,N_5411,N_6327);
and U13854 (N_13854,N_5716,N_5953);
nand U13855 (N_13855,N_5898,N_9004);
xor U13856 (N_13856,N_7988,N_8482);
and U13857 (N_13857,N_9632,N_8327);
or U13858 (N_13858,N_7977,N_8525);
nand U13859 (N_13859,N_9455,N_7238);
or U13860 (N_13860,N_5103,N_5846);
or U13861 (N_13861,N_6416,N_9854);
nor U13862 (N_13862,N_5628,N_7458);
nor U13863 (N_13863,N_5160,N_9541);
xor U13864 (N_13864,N_6060,N_7805);
nand U13865 (N_13865,N_7885,N_8869);
xnor U13866 (N_13866,N_9912,N_5587);
and U13867 (N_13867,N_5568,N_9146);
nor U13868 (N_13868,N_6867,N_7745);
nand U13869 (N_13869,N_7750,N_8113);
nor U13870 (N_13870,N_8962,N_6776);
nor U13871 (N_13871,N_9452,N_7523);
nand U13872 (N_13872,N_8247,N_5109);
nand U13873 (N_13873,N_8906,N_5744);
or U13874 (N_13874,N_7702,N_8990);
or U13875 (N_13875,N_5202,N_8170);
and U13876 (N_13876,N_9074,N_9517);
and U13877 (N_13877,N_5067,N_6918);
and U13878 (N_13878,N_6775,N_6795);
nand U13879 (N_13879,N_6195,N_5828);
xnor U13880 (N_13880,N_9876,N_9278);
xnor U13881 (N_13881,N_9173,N_9680);
nand U13882 (N_13882,N_9600,N_7180);
nand U13883 (N_13883,N_8923,N_8084);
and U13884 (N_13884,N_5019,N_7384);
xor U13885 (N_13885,N_9116,N_5655);
nand U13886 (N_13886,N_6980,N_7204);
nand U13887 (N_13887,N_8164,N_9900);
nor U13888 (N_13888,N_6598,N_6215);
and U13889 (N_13889,N_9349,N_6392);
nand U13890 (N_13890,N_9425,N_9429);
or U13891 (N_13891,N_6439,N_9070);
and U13892 (N_13892,N_7651,N_7407);
xor U13893 (N_13893,N_9246,N_5302);
nor U13894 (N_13894,N_5281,N_7044);
nand U13895 (N_13895,N_8234,N_9429);
nand U13896 (N_13896,N_8008,N_6426);
nor U13897 (N_13897,N_9004,N_6039);
or U13898 (N_13898,N_7767,N_7492);
or U13899 (N_13899,N_8527,N_5228);
nor U13900 (N_13900,N_8048,N_6310);
xnor U13901 (N_13901,N_6207,N_5744);
or U13902 (N_13902,N_8501,N_6786);
nand U13903 (N_13903,N_5651,N_8871);
and U13904 (N_13904,N_8651,N_8143);
nor U13905 (N_13905,N_7186,N_7174);
or U13906 (N_13906,N_5568,N_6920);
or U13907 (N_13907,N_5440,N_8154);
or U13908 (N_13908,N_9038,N_9483);
nand U13909 (N_13909,N_7497,N_9030);
or U13910 (N_13910,N_9787,N_6923);
or U13911 (N_13911,N_9331,N_9424);
or U13912 (N_13912,N_8199,N_6001);
and U13913 (N_13913,N_9461,N_7658);
and U13914 (N_13914,N_9570,N_5869);
nor U13915 (N_13915,N_9679,N_5657);
or U13916 (N_13916,N_5410,N_6168);
nor U13917 (N_13917,N_8805,N_6811);
nand U13918 (N_13918,N_9248,N_6971);
and U13919 (N_13919,N_6279,N_8916);
and U13920 (N_13920,N_6780,N_5831);
and U13921 (N_13921,N_7490,N_9455);
and U13922 (N_13922,N_6487,N_9964);
and U13923 (N_13923,N_9401,N_6286);
or U13924 (N_13924,N_6602,N_7668);
and U13925 (N_13925,N_8956,N_6379);
xnor U13926 (N_13926,N_7918,N_8859);
and U13927 (N_13927,N_9219,N_5920);
or U13928 (N_13928,N_8070,N_7456);
and U13929 (N_13929,N_6313,N_5190);
nand U13930 (N_13930,N_6681,N_8423);
and U13931 (N_13931,N_7297,N_6343);
nand U13932 (N_13932,N_7229,N_6373);
nor U13933 (N_13933,N_6679,N_8895);
and U13934 (N_13934,N_9259,N_8143);
and U13935 (N_13935,N_8834,N_7123);
xor U13936 (N_13936,N_5331,N_9643);
xnor U13937 (N_13937,N_9036,N_7998);
nand U13938 (N_13938,N_5497,N_6588);
nor U13939 (N_13939,N_7440,N_8145);
nor U13940 (N_13940,N_6634,N_8686);
nand U13941 (N_13941,N_8045,N_5055);
xnor U13942 (N_13942,N_7139,N_9816);
xnor U13943 (N_13943,N_6077,N_9955);
nand U13944 (N_13944,N_6133,N_8595);
or U13945 (N_13945,N_8437,N_9764);
xor U13946 (N_13946,N_5926,N_7566);
and U13947 (N_13947,N_7934,N_7807);
nand U13948 (N_13948,N_9769,N_8769);
nand U13949 (N_13949,N_5666,N_8456);
and U13950 (N_13950,N_7985,N_9332);
nand U13951 (N_13951,N_9673,N_5062);
or U13952 (N_13952,N_6804,N_8129);
xnor U13953 (N_13953,N_6652,N_7245);
nand U13954 (N_13954,N_6916,N_9286);
nand U13955 (N_13955,N_7180,N_8187);
xnor U13956 (N_13956,N_7712,N_9083);
and U13957 (N_13957,N_5840,N_9284);
and U13958 (N_13958,N_7530,N_9996);
nand U13959 (N_13959,N_8174,N_8582);
nand U13960 (N_13960,N_5880,N_9929);
and U13961 (N_13961,N_7731,N_6068);
or U13962 (N_13962,N_8728,N_6692);
xnor U13963 (N_13963,N_5840,N_6374);
nand U13964 (N_13964,N_6564,N_7636);
and U13965 (N_13965,N_6734,N_7633);
nand U13966 (N_13966,N_7086,N_6698);
and U13967 (N_13967,N_6147,N_7106);
nor U13968 (N_13968,N_7153,N_7822);
or U13969 (N_13969,N_5081,N_7306);
nor U13970 (N_13970,N_8019,N_5586);
and U13971 (N_13971,N_5767,N_5186);
nand U13972 (N_13972,N_9756,N_8452);
or U13973 (N_13973,N_9833,N_5637);
and U13974 (N_13974,N_5719,N_8841);
and U13975 (N_13975,N_5714,N_8983);
and U13976 (N_13976,N_7880,N_8880);
xnor U13977 (N_13977,N_9787,N_6932);
nand U13978 (N_13978,N_7833,N_8643);
and U13979 (N_13979,N_7346,N_6313);
and U13980 (N_13980,N_5238,N_9056);
and U13981 (N_13981,N_9985,N_9942);
nand U13982 (N_13982,N_7618,N_6757);
or U13983 (N_13983,N_8656,N_7834);
nor U13984 (N_13984,N_8033,N_8071);
nor U13985 (N_13985,N_9964,N_6898);
or U13986 (N_13986,N_7840,N_9902);
and U13987 (N_13987,N_5081,N_8729);
xor U13988 (N_13988,N_8535,N_5433);
nand U13989 (N_13989,N_5600,N_7948);
or U13990 (N_13990,N_5247,N_7799);
xor U13991 (N_13991,N_5154,N_9347);
or U13992 (N_13992,N_5084,N_5708);
and U13993 (N_13993,N_8643,N_5576);
nand U13994 (N_13994,N_9086,N_6083);
and U13995 (N_13995,N_9494,N_5225);
nand U13996 (N_13996,N_6284,N_7440);
xor U13997 (N_13997,N_7167,N_6807);
or U13998 (N_13998,N_5173,N_5005);
nor U13999 (N_13999,N_5373,N_6764);
and U14000 (N_14000,N_8600,N_9900);
xor U14001 (N_14001,N_8172,N_6554);
or U14002 (N_14002,N_9556,N_9959);
nand U14003 (N_14003,N_6535,N_9491);
xor U14004 (N_14004,N_9918,N_5712);
and U14005 (N_14005,N_5289,N_7772);
and U14006 (N_14006,N_8973,N_6907);
nand U14007 (N_14007,N_5780,N_6888);
nor U14008 (N_14008,N_9578,N_9231);
xor U14009 (N_14009,N_8975,N_8282);
nand U14010 (N_14010,N_9392,N_5090);
nor U14011 (N_14011,N_5778,N_8967);
nor U14012 (N_14012,N_6877,N_5083);
nor U14013 (N_14013,N_8261,N_7817);
and U14014 (N_14014,N_5125,N_6404);
or U14015 (N_14015,N_5230,N_5675);
nor U14016 (N_14016,N_7281,N_7748);
xnor U14017 (N_14017,N_8499,N_5059);
nand U14018 (N_14018,N_8173,N_8223);
and U14019 (N_14019,N_9763,N_5480);
or U14020 (N_14020,N_8238,N_5146);
and U14021 (N_14021,N_9212,N_8882);
and U14022 (N_14022,N_9171,N_5510);
or U14023 (N_14023,N_5248,N_5044);
xnor U14024 (N_14024,N_7333,N_7409);
nand U14025 (N_14025,N_8381,N_8600);
and U14026 (N_14026,N_9400,N_8738);
nand U14027 (N_14027,N_5010,N_6811);
nand U14028 (N_14028,N_8270,N_5764);
nand U14029 (N_14029,N_8346,N_7003);
and U14030 (N_14030,N_8068,N_5626);
and U14031 (N_14031,N_9413,N_9254);
nand U14032 (N_14032,N_5398,N_9105);
nor U14033 (N_14033,N_7693,N_9759);
or U14034 (N_14034,N_5985,N_9482);
xnor U14035 (N_14035,N_5252,N_6426);
xor U14036 (N_14036,N_5169,N_6277);
nor U14037 (N_14037,N_6687,N_7635);
nand U14038 (N_14038,N_9541,N_5670);
nand U14039 (N_14039,N_9074,N_5278);
and U14040 (N_14040,N_5431,N_6007);
nand U14041 (N_14041,N_6572,N_6672);
nor U14042 (N_14042,N_6822,N_6088);
nand U14043 (N_14043,N_5496,N_9377);
or U14044 (N_14044,N_9991,N_6880);
and U14045 (N_14045,N_9059,N_6606);
or U14046 (N_14046,N_7584,N_5685);
or U14047 (N_14047,N_9759,N_8487);
nand U14048 (N_14048,N_6603,N_5567);
nand U14049 (N_14049,N_5910,N_5819);
xnor U14050 (N_14050,N_8461,N_6411);
nand U14051 (N_14051,N_8857,N_8580);
and U14052 (N_14052,N_8043,N_9614);
nor U14053 (N_14053,N_8242,N_9588);
xnor U14054 (N_14054,N_9015,N_6112);
nor U14055 (N_14055,N_9499,N_6520);
and U14056 (N_14056,N_8772,N_8912);
nand U14057 (N_14057,N_6575,N_8424);
nand U14058 (N_14058,N_5603,N_9668);
xor U14059 (N_14059,N_6616,N_5444);
nand U14060 (N_14060,N_7108,N_9159);
xor U14061 (N_14061,N_7782,N_7706);
and U14062 (N_14062,N_5281,N_7085);
or U14063 (N_14063,N_9148,N_5804);
and U14064 (N_14064,N_8173,N_9617);
or U14065 (N_14065,N_8971,N_5498);
xnor U14066 (N_14066,N_5718,N_8273);
nor U14067 (N_14067,N_6389,N_6877);
nand U14068 (N_14068,N_6366,N_8082);
or U14069 (N_14069,N_5152,N_7760);
and U14070 (N_14070,N_6090,N_5338);
xor U14071 (N_14071,N_5190,N_7752);
or U14072 (N_14072,N_8560,N_5835);
and U14073 (N_14073,N_5951,N_5290);
nand U14074 (N_14074,N_8275,N_8615);
or U14075 (N_14075,N_9375,N_6059);
nor U14076 (N_14076,N_5557,N_6021);
or U14077 (N_14077,N_8594,N_6780);
xnor U14078 (N_14078,N_7422,N_8441);
and U14079 (N_14079,N_6667,N_9169);
nor U14080 (N_14080,N_9089,N_7083);
or U14081 (N_14081,N_8077,N_5138);
nand U14082 (N_14082,N_6358,N_5243);
nor U14083 (N_14083,N_6654,N_5314);
nor U14084 (N_14084,N_6125,N_6793);
or U14085 (N_14085,N_6885,N_9453);
or U14086 (N_14086,N_5713,N_5675);
nand U14087 (N_14087,N_6757,N_9810);
and U14088 (N_14088,N_5775,N_9185);
xnor U14089 (N_14089,N_9822,N_9076);
nand U14090 (N_14090,N_7070,N_9656);
nor U14091 (N_14091,N_5828,N_8071);
or U14092 (N_14092,N_8412,N_5156);
and U14093 (N_14093,N_5513,N_5141);
nor U14094 (N_14094,N_9836,N_8313);
xor U14095 (N_14095,N_9313,N_8919);
nor U14096 (N_14096,N_5002,N_9430);
or U14097 (N_14097,N_6866,N_6539);
nand U14098 (N_14098,N_7316,N_7227);
xnor U14099 (N_14099,N_7473,N_8434);
nand U14100 (N_14100,N_9690,N_5321);
nor U14101 (N_14101,N_7602,N_7506);
and U14102 (N_14102,N_5164,N_7876);
nor U14103 (N_14103,N_9969,N_7423);
xor U14104 (N_14104,N_5041,N_7825);
nor U14105 (N_14105,N_8839,N_6939);
xor U14106 (N_14106,N_9771,N_7709);
nand U14107 (N_14107,N_5760,N_5481);
nand U14108 (N_14108,N_9424,N_8813);
and U14109 (N_14109,N_6349,N_5437);
and U14110 (N_14110,N_6948,N_9128);
xnor U14111 (N_14111,N_9900,N_6433);
and U14112 (N_14112,N_8742,N_7351);
xnor U14113 (N_14113,N_5531,N_9230);
nand U14114 (N_14114,N_8925,N_5148);
nand U14115 (N_14115,N_6025,N_5731);
nand U14116 (N_14116,N_6885,N_7435);
xnor U14117 (N_14117,N_7413,N_6977);
and U14118 (N_14118,N_8122,N_5625);
and U14119 (N_14119,N_5978,N_9892);
nand U14120 (N_14120,N_5098,N_9690);
nand U14121 (N_14121,N_8803,N_8305);
nand U14122 (N_14122,N_6203,N_8745);
and U14123 (N_14123,N_7297,N_6801);
nor U14124 (N_14124,N_7529,N_6368);
xnor U14125 (N_14125,N_9193,N_5905);
xor U14126 (N_14126,N_7992,N_6595);
or U14127 (N_14127,N_5826,N_7358);
nor U14128 (N_14128,N_8808,N_6374);
nand U14129 (N_14129,N_8474,N_9048);
and U14130 (N_14130,N_7952,N_6668);
xnor U14131 (N_14131,N_8596,N_6150);
xor U14132 (N_14132,N_7445,N_8746);
or U14133 (N_14133,N_8879,N_6157);
nor U14134 (N_14134,N_6028,N_5227);
xnor U14135 (N_14135,N_6906,N_6845);
or U14136 (N_14136,N_8369,N_6721);
and U14137 (N_14137,N_5312,N_8396);
or U14138 (N_14138,N_6331,N_9983);
xnor U14139 (N_14139,N_6856,N_6028);
and U14140 (N_14140,N_8982,N_6631);
nor U14141 (N_14141,N_8629,N_5379);
xnor U14142 (N_14142,N_6030,N_9529);
nand U14143 (N_14143,N_7182,N_7672);
or U14144 (N_14144,N_5384,N_5996);
nor U14145 (N_14145,N_5117,N_7454);
nand U14146 (N_14146,N_7794,N_7019);
xnor U14147 (N_14147,N_7890,N_6278);
nand U14148 (N_14148,N_8241,N_9413);
nor U14149 (N_14149,N_6408,N_8381);
nor U14150 (N_14150,N_8075,N_6029);
or U14151 (N_14151,N_6006,N_8464);
xnor U14152 (N_14152,N_7541,N_6861);
nor U14153 (N_14153,N_7048,N_7637);
or U14154 (N_14154,N_7407,N_8331);
nand U14155 (N_14155,N_7017,N_7663);
xnor U14156 (N_14156,N_6387,N_7305);
and U14157 (N_14157,N_6993,N_5403);
nor U14158 (N_14158,N_7981,N_8337);
or U14159 (N_14159,N_8952,N_8041);
nor U14160 (N_14160,N_9595,N_5690);
nand U14161 (N_14161,N_6973,N_6993);
nand U14162 (N_14162,N_8186,N_5104);
nand U14163 (N_14163,N_7935,N_8428);
xor U14164 (N_14164,N_6581,N_6818);
and U14165 (N_14165,N_8197,N_8238);
and U14166 (N_14166,N_8538,N_6634);
nand U14167 (N_14167,N_6304,N_6685);
nor U14168 (N_14168,N_9669,N_9968);
nor U14169 (N_14169,N_8120,N_8939);
or U14170 (N_14170,N_6574,N_9194);
or U14171 (N_14171,N_5631,N_6099);
or U14172 (N_14172,N_6432,N_8448);
nor U14173 (N_14173,N_5724,N_8149);
xnor U14174 (N_14174,N_5411,N_7123);
xnor U14175 (N_14175,N_5504,N_5798);
and U14176 (N_14176,N_6010,N_7114);
xnor U14177 (N_14177,N_8242,N_6727);
xnor U14178 (N_14178,N_9226,N_7320);
and U14179 (N_14179,N_8485,N_7907);
nor U14180 (N_14180,N_7952,N_9044);
or U14181 (N_14181,N_5943,N_8129);
and U14182 (N_14182,N_7723,N_9029);
and U14183 (N_14183,N_7055,N_7314);
and U14184 (N_14184,N_6789,N_8865);
xor U14185 (N_14185,N_8584,N_9129);
or U14186 (N_14186,N_8936,N_7555);
nand U14187 (N_14187,N_9526,N_7513);
or U14188 (N_14188,N_7151,N_6978);
nor U14189 (N_14189,N_6657,N_6492);
nor U14190 (N_14190,N_7932,N_6672);
nor U14191 (N_14191,N_5726,N_7192);
nor U14192 (N_14192,N_6324,N_6209);
nor U14193 (N_14193,N_8600,N_6341);
or U14194 (N_14194,N_9433,N_6952);
nand U14195 (N_14195,N_9830,N_9548);
nor U14196 (N_14196,N_9597,N_6080);
or U14197 (N_14197,N_9891,N_8604);
nand U14198 (N_14198,N_7613,N_6143);
and U14199 (N_14199,N_8309,N_7268);
nor U14200 (N_14200,N_7871,N_7643);
or U14201 (N_14201,N_7314,N_9042);
nor U14202 (N_14202,N_8945,N_5255);
and U14203 (N_14203,N_7358,N_6770);
or U14204 (N_14204,N_8648,N_6157);
and U14205 (N_14205,N_6049,N_6520);
nand U14206 (N_14206,N_7717,N_8432);
and U14207 (N_14207,N_6352,N_9136);
nand U14208 (N_14208,N_5107,N_9049);
nand U14209 (N_14209,N_8570,N_8427);
nor U14210 (N_14210,N_8526,N_7992);
xor U14211 (N_14211,N_9765,N_8992);
xnor U14212 (N_14212,N_6187,N_8307);
and U14213 (N_14213,N_8619,N_5322);
xor U14214 (N_14214,N_5134,N_8436);
or U14215 (N_14215,N_9411,N_5536);
nor U14216 (N_14216,N_9634,N_6977);
and U14217 (N_14217,N_6903,N_9980);
xnor U14218 (N_14218,N_9134,N_9620);
and U14219 (N_14219,N_7361,N_8918);
nand U14220 (N_14220,N_9922,N_9569);
nor U14221 (N_14221,N_6691,N_7129);
or U14222 (N_14222,N_8658,N_6853);
or U14223 (N_14223,N_6029,N_5552);
xor U14224 (N_14224,N_7551,N_8797);
xor U14225 (N_14225,N_6964,N_9689);
xnor U14226 (N_14226,N_7990,N_5825);
and U14227 (N_14227,N_8586,N_5005);
or U14228 (N_14228,N_6825,N_9118);
nand U14229 (N_14229,N_5079,N_8127);
and U14230 (N_14230,N_5232,N_7089);
nor U14231 (N_14231,N_8323,N_9002);
xnor U14232 (N_14232,N_9554,N_5245);
nand U14233 (N_14233,N_6536,N_9891);
nor U14234 (N_14234,N_6339,N_7878);
nand U14235 (N_14235,N_5114,N_7947);
or U14236 (N_14236,N_7171,N_7438);
and U14237 (N_14237,N_9791,N_6216);
nor U14238 (N_14238,N_6643,N_6623);
or U14239 (N_14239,N_9632,N_6682);
xor U14240 (N_14240,N_6708,N_6473);
and U14241 (N_14241,N_5574,N_9977);
nor U14242 (N_14242,N_8013,N_6357);
nor U14243 (N_14243,N_9826,N_6604);
or U14244 (N_14244,N_7230,N_6571);
and U14245 (N_14245,N_5196,N_5442);
nand U14246 (N_14246,N_5102,N_5741);
and U14247 (N_14247,N_8199,N_6490);
xnor U14248 (N_14248,N_6132,N_6780);
xnor U14249 (N_14249,N_7498,N_9385);
nor U14250 (N_14250,N_6733,N_7281);
nand U14251 (N_14251,N_8930,N_5902);
nand U14252 (N_14252,N_5445,N_8963);
and U14253 (N_14253,N_9473,N_7675);
nand U14254 (N_14254,N_9368,N_9966);
nor U14255 (N_14255,N_6047,N_9142);
nand U14256 (N_14256,N_5587,N_7272);
and U14257 (N_14257,N_5086,N_8321);
and U14258 (N_14258,N_5153,N_7689);
nor U14259 (N_14259,N_8207,N_5713);
xnor U14260 (N_14260,N_8376,N_6408);
or U14261 (N_14261,N_9441,N_7705);
and U14262 (N_14262,N_5179,N_6725);
nor U14263 (N_14263,N_6464,N_6050);
nand U14264 (N_14264,N_6335,N_7239);
or U14265 (N_14265,N_6569,N_8811);
xnor U14266 (N_14266,N_8891,N_5639);
and U14267 (N_14267,N_6722,N_5579);
nand U14268 (N_14268,N_6353,N_5887);
nor U14269 (N_14269,N_8492,N_6897);
xor U14270 (N_14270,N_6957,N_5117);
and U14271 (N_14271,N_7452,N_7852);
and U14272 (N_14272,N_8962,N_7519);
and U14273 (N_14273,N_6753,N_8532);
nor U14274 (N_14274,N_8541,N_6632);
nand U14275 (N_14275,N_8453,N_7615);
xor U14276 (N_14276,N_5820,N_8487);
nand U14277 (N_14277,N_7933,N_5047);
nand U14278 (N_14278,N_5083,N_6399);
xnor U14279 (N_14279,N_6734,N_5946);
nand U14280 (N_14280,N_8669,N_7188);
nor U14281 (N_14281,N_7363,N_6647);
nand U14282 (N_14282,N_9317,N_8424);
and U14283 (N_14283,N_9417,N_9245);
nand U14284 (N_14284,N_7445,N_5344);
nand U14285 (N_14285,N_9533,N_5213);
or U14286 (N_14286,N_5022,N_7411);
or U14287 (N_14287,N_5378,N_8477);
or U14288 (N_14288,N_5189,N_6661);
nor U14289 (N_14289,N_9542,N_8752);
nor U14290 (N_14290,N_9115,N_9396);
or U14291 (N_14291,N_9601,N_6671);
and U14292 (N_14292,N_5691,N_8912);
nor U14293 (N_14293,N_7590,N_6304);
xnor U14294 (N_14294,N_9197,N_9245);
xnor U14295 (N_14295,N_9786,N_9333);
xor U14296 (N_14296,N_9458,N_5648);
nand U14297 (N_14297,N_9731,N_6496);
nand U14298 (N_14298,N_8266,N_5152);
xor U14299 (N_14299,N_7323,N_6287);
nor U14300 (N_14300,N_9819,N_7723);
xor U14301 (N_14301,N_7771,N_6453);
and U14302 (N_14302,N_5236,N_8587);
nor U14303 (N_14303,N_9002,N_7327);
nand U14304 (N_14304,N_7848,N_5153);
or U14305 (N_14305,N_5516,N_9519);
xnor U14306 (N_14306,N_6225,N_5852);
xor U14307 (N_14307,N_5703,N_9552);
nor U14308 (N_14308,N_9407,N_9040);
and U14309 (N_14309,N_8531,N_8113);
and U14310 (N_14310,N_6288,N_7329);
and U14311 (N_14311,N_6623,N_8847);
and U14312 (N_14312,N_5790,N_9986);
nor U14313 (N_14313,N_8237,N_7368);
xor U14314 (N_14314,N_6099,N_5861);
nand U14315 (N_14315,N_9411,N_9737);
nand U14316 (N_14316,N_5047,N_7530);
or U14317 (N_14317,N_7939,N_8123);
and U14318 (N_14318,N_7791,N_6778);
and U14319 (N_14319,N_5210,N_6743);
xor U14320 (N_14320,N_9470,N_7829);
xnor U14321 (N_14321,N_6318,N_6316);
nand U14322 (N_14322,N_5344,N_9665);
or U14323 (N_14323,N_8140,N_8210);
or U14324 (N_14324,N_5647,N_6458);
xnor U14325 (N_14325,N_6940,N_5979);
nor U14326 (N_14326,N_5674,N_8158);
nand U14327 (N_14327,N_6907,N_6260);
nor U14328 (N_14328,N_9763,N_8455);
or U14329 (N_14329,N_6386,N_5146);
nand U14330 (N_14330,N_7452,N_9642);
nand U14331 (N_14331,N_7992,N_9529);
xor U14332 (N_14332,N_9779,N_9238);
nand U14333 (N_14333,N_8766,N_6723);
nand U14334 (N_14334,N_5095,N_6733);
xnor U14335 (N_14335,N_7141,N_6345);
or U14336 (N_14336,N_9596,N_5742);
nor U14337 (N_14337,N_6370,N_6827);
nand U14338 (N_14338,N_8185,N_5756);
and U14339 (N_14339,N_9804,N_9748);
or U14340 (N_14340,N_6250,N_8474);
xnor U14341 (N_14341,N_8684,N_9399);
and U14342 (N_14342,N_8016,N_8116);
xnor U14343 (N_14343,N_5083,N_6347);
nand U14344 (N_14344,N_6378,N_9714);
nor U14345 (N_14345,N_7113,N_8937);
nor U14346 (N_14346,N_7761,N_5782);
or U14347 (N_14347,N_6328,N_8561);
nor U14348 (N_14348,N_7550,N_9412);
and U14349 (N_14349,N_5125,N_9392);
nor U14350 (N_14350,N_5734,N_6069);
or U14351 (N_14351,N_8601,N_9366);
or U14352 (N_14352,N_7237,N_8831);
or U14353 (N_14353,N_7566,N_7594);
and U14354 (N_14354,N_5054,N_7451);
or U14355 (N_14355,N_7740,N_5565);
and U14356 (N_14356,N_8327,N_9226);
xnor U14357 (N_14357,N_8816,N_6748);
and U14358 (N_14358,N_8659,N_7881);
nor U14359 (N_14359,N_7833,N_8972);
nor U14360 (N_14360,N_5641,N_6058);
nor U14361 (N_14361,N_6807,N_7361);
xor U14362 (N_14362,N_8483,N_6859);
or U14363 (N_14363,N_7737,N_5510);
or U14364 (N_14364,N_7345,N_5794);
xor U14365 (N_14365,N_5448,N_6985);
or U14366 (N_14366,N_9061,N_8478);
nand U14367 (N_14367,N_9996,N_9593);
nor U14368 (N_14368,N_5751,N_9942);
nor U14369 (N_14369,N_6655,N_8098);
and U14370 (N_14370,N_8634,N_9219);
xnor U14371 (N_14371,N_7408,N_7851);
and U14372 (N_14372,N_7059,N_6031);
or U14373 (N_14373,N_9916,N_9614);
and U14374 (N_14374,N_5633,N_6004);
or U14375 (N_14375,N_7111,N_9911);
or U14376 (N_14376,N_5896,N_8598);
xor U14377 (N_14377,N_8516,N_5683);
nand U14378 (N_14378,N_9723,N_8215);
xnor U14379 (N_14379,N_9479,N_5851);
xnor U14380 (N_14380,N_9053,N_7523);
and U14381 (N_14381,N_6608,N_8561);
or U14382 (N_14382,N_8270,N_8844);
nand U14383 (N_14383,N_6387,N_7236);
xor U14384 (N_14384,N_8577,N_5235);
nor U14385 (N_14385,N_5829,N_8050);
nand U14386 (N_14386,N_7728,N_6098);
xor U14387 (N_14387,N_8950,N_7373);
nor U14388 (N_14388,N_9330,N_7906);
or U14389 (N_14389,N_5051,N_5594);
xor U14390 (N_14390,N_6989,N_8416);
nor U14391 (N_14391,N_5765,N_8496);
and U14392 (N_14392,N_9258,N_9818);
and U14393 (N_14393,N_6719,N_5725);
xor U14394 (N_14394,N_9468,N_5259);
or U14395 (N_14395,N_6080,N_6177);
or U14396 (N_14396,N_7074,N_8081);
xnor U14397 (N_14397,N_8607,N_9826);
and U14398 (N_14398,N_7461,N_6112);
xnor U14399 (N_14399,N_8648,N_9951);
nand U14400 (N_14400,N_9618,N_6496);
xor U14401 (N_14401,N_9746,N_9929);
or U14402 (N_14402,N_5480,N_9247);
or U14403 (N_14403,N_5274,N_8048);
or U14404 (N_14404,N_6356,N_5499);
nor U14405 (N_14405,N_7650,N_7417);
xor U14406 (N_14406,N_7156,N_9537);
nor U14407 (N_14407,N_8394,N_9102);
nor U14408 (N_14408,N_7499,N_7669);
or U14409 (N_14409,N_8339,N_7495);
or U14410 (N_14410,N_8648,N_9719);
or U14411 (N_14411,N_6215,N_8504);
and U14412 (N_14412,N_9238,N_8268);
xor U14413 (N_14413,N_5762,N_5060);
nor U14414 (N_14414,N_8904,N_7357);
or U14415 (N_14415,N_8624,N_9005);
and U14416 (N_14416,N_8061,N_6256);
nor U14417 (N_14417,N_8655,N_6168);
nand U14418 (N_14418,N_5879,N_9843);
nand U14419 (N_14419,N_8513,N_7432);
xnor U14420 (N_14420,N_5045,N_7254);
xnor U14421 (N_14421,N_7637,N_7049);
or U14422 (N_14422,N_5558,N_6201);
nor U14423 (N_14423,N_5400,N_7384);
xnor U14424 (N_14424,N_6807,N_5904);
and U14425 (N_14425,N_5386,N_5376);
xor U14426 (N_14426,N_9605,N_7223);
nand U14427 (N_14427,N_6424,N_6502);
nand U14428 (N_14428,N_6594,N_9377);
xnor U14429 (N_14429,N_7003,N_6273);
and U14430 (N_14430,N_7932,N_7687);
or U14431 (N_14431,N_6666,N_9187);
xnor U14432 (N_14432,N_5886,N_5234);
nor U14433 (N_14433,N_9884,N_5184);
nor U14434 (N_14434,N_6394,N_9448);
nor U14435 (N_14435,N_5601,N_7379);
and U14436 (N_14436,N_5130,N_6075);
nor U14437 (N_14437,N_8036,N_9630);
xor U14438 (N_14438,N_7730,N_6958);
and U14439 (N_14439,N_5823,N_8589);
xnor U14440 (N_14440,N_7971,N_7368);
xor U14441 (N_14441,N_9742,N_5586);
or U14442 (N_14442,N_6340,N_8401);
xnor U14443 (N_14443,N_7768,N_9886);
nor U14444 (N_14444,N_7919,N_9535);
nor U14445 (N_14445,N_8086,N_7780);
or U14446 (N_14446,N_5094,N_6391);
and U14447 (N_14447,N_8813,N_9716);
nand U14448 (N_14448,N_7427,N_8994);
nand U14449 (N_14449,N_8549,N_5726);
xnor U14450 (N_14450,N_8394,N_9613);
or U14451 (N_14451,N_9979,N_7528);
nor U14452 (N_14452,N_6132,N_6229);
and U14453 (N_14453,N_9730,N_8896);
and U14454 (N_14454,N_8740,N_9303);
or U14455 (N_14455,N_7362,N_6885);
xnor U14456 (N_14456,N_7937,N_8830);
nand U14457 (N_14457,N_6975,N_8072);
or U14458 (N_14458,N_7028,N_6219);
xor U14459 (N_14459,N_9293,N_7256);
nor U14460 (N_14460,N_8988,N_9921);
and U14461 (N_14461,N_7765,N_5738);
xnor U14462 (N_14462,N_6937,N_6226);
nor U14463 (N_14463,N_6465,N_5668);
xnor U14464 (N_14464,N_9279,N_5988);
nand U14465 (N_14465,N_5216,N_8195);
xor U14466 (N_14466,N_6979,N_7636);
nor U14467 (N_14467,N_9675,N_5200);
or U14468 (N_14468,N_5187,N_6334);
and U14469 (N_14469,N_5592,N_6631);
or U14470 (N_14470,N_9717,N_8482);
and U14471 (N_14471,N_7599,N_6538);
or U14472 (N_14472,N_8433,N_5056);
nor U14473 (N_14473,N_7390,N_7341);
and U14474 (N_14474,N_5378,N_6308);
nor U14475 (N_14475,N_7872,N_6411);
and U14476 (N_14476,N_5833,N_9674);
nand U14477 (N_14477,N_9480,N_6962);
xor U14478 (N_14478,N_8841,N_5314);
nand U14479 (N_14479,N_5131,N_8875);
and U14480 (N_14480,N_9295,N_9614);
nand U14481 (N_14481,N_8679,N_5838);
or U14482 (N_14482,N_7659,N_6540);
nand U14483 (N_14483,N_8189,N_7155);
xnor U14484 (N_14484,N_9512,N_8556);
xnor U14485 (N_14485,N_9662,N_5146);
nand U14486 (N_14486,N_5291,N_6737);
xor U14487 (N_14487,N_5921,N_9474);
and U14488 (N_14488,N_6092,N_8701);
or U14489 (N_14489,N_8390,N_5028);
and U14490 (N_14490,N_7346,N_6765);
and U14491 (N_14491,N_9793,N_9585);
and U14492 (N_14492,N_8931,N_6929);
xor U14493 (N_14493,N_7547,N_8546);
nand U14494 (N_14494,N_6010,N_7484);
nor U14495 (N_14495,N_9011,N_8955);
nand U14496 (N_14496,N_9954,N_6332);
nand U14497 (N_14497,N_8186,N_9559);
nand U14498 (N_14498,N_6404,N_5993);
xnor U14499 (N_14499,N_7326,N_7817);
or U14500 (N_14500,N_6637,N_9176);
nor U14501 (N_14501,N_7972,N_8377);
nand U14502 (N_14502,N_5297,N_7550);
xor U14503 (N_14503,N_9791,N_6504);
and U14504 (N_14504,N_9776,N_9811);
and U14505 (N_14505,N_9133,N_7689);
nor U14506 (N_14506,N_7459,N_9529);
xnor U14507 (N_14507,N_8650,N_9275);
xnor U14508 (N_14508,N_7002,N_7110);
or U14509 (N_14509,N_5803,N_6626);
or U14510 (N_14510,N_8424,N_6370);
nor U14511 (N_14511,N_5721,N_7635);
and U14512 (N_14512,N_8705,N_7749);
and U14513 (N_14513,N_6499,N_8521);
xnor U14514 (N_14514,N_7363,N_6371);
or U14515 (N_14515,N_8754,N_5629);
and U14516 (N_14516,N_9750,N_6653);
or U14517 (N_14517,N_5173,N_8111);
nand U14518 (N_14518,N_9051,N_5557);
nor U14519 (N_14519,N_9842,N_7451);
nand U14520 (N_14520,N_5809,N_9442);
nand U14521 (N_14521,N_5091,N_9927);
or U14522 (N_14522,N_6585,N_9314);
xor U14523 (N_14523,N_9258,N_6851);
or U14524 (N_14524,N_8352,N_9522);
xor U14525 (N_14525,N_6971,N_8585);
or U14526 (N_14526,N_5292,N_5530);
nand U14527 (N_14527,N_9604,N_9460);
nor U14528 (N_14528,N_5021,N_8030);
xor U14529 (N_14529,N_8866,N_9089);
or U14530 (N_14530,N_6343,N_6857);
nand U14531 (N_14531,N_5776,N_9686);
xnor U14532 (N_14532,N_9726,N_8354);
nand U14533 (N_14533,N_7653,N_7261);
xor U14534 (N_14534,N_8814,N_6751);
or U14535 (N_14535,N_7526,N_9598);
nand U14536 (N_14536,N_8587,N_7930);
nor U14537 (N_14537,N_9745,N_5951);
xor U14538 (N_14538,N_9957,N_5018);
nand U14539 (N_14539,N_7162,N_8836);
or U14540 (N_14540,N_8955,N_5656);
xor U14541 (N_14541,N_7268,N_8142);
xnor U14542 (N_14542,N_8597,N_7492);
xor U14543 (N_14543,N_7238,N_5864);
nand U14544 (N_14544,N_7263,N_7260);
nor U14545 (N_14545,N_9620,N_6363);
nand U14546 (N_14546,N_7764,N_6502);
nor U14547 (N_14547,N_7628,N_6701);
nand U14548 (N_14548,N_8735,N_9038);
and U14549 (N_14549,N_8118,N_6194);
nor U14550 (N_14550,N_7226,N_5638);
or U14551 (N_14551,N_7662,N_5394);
xnor U14552 (N_14552,N_5819,N_8461);
and U14553 (N_14553,N_5634,N_6988);
nor U14554 (N_14554,N_5085,N_5579);
xor U14555 (N_14555,N_8199,N_5620);
nor U14556 (N_14556,N_9544,N_5313);
nor U14557 (N_14557,N_5023,N_7694);
nand U14558 (N_14558,N_6589,N_9579);
or U14559 (N_14559,N_5866,N_9214);
nand U14560 (N_14560,N_7972,N_9288);
nor U14561 (N_14561,N_8600,N_8704);
or U14562 (N_14562,N_7938,N_7378);
xor U14563 (N_14563,N_5708,N_6681);
nand U14564 (N_14564,N_5026,N_5806);
or U14565 (N_14565,N_7533,N_7484);
and U14566 (N_14566,N_7671,N_5528);
or U14567 (N_14567,N_5125,N_6882);
xnor U14568 (N_14568,N_6644,N_9109);
nand U14569 (N_14569,N_6927,N_8591);
and U14570 (N_14570,N_6895,N_6921);
and U14571 (N_14571,N_5560,N_7272);
nor U14572 (N_14572,N_7394,N_6052);
or U14573 (N_14573,N_6435,N_5147);
nor U14574 (N_14574,N_8517,N_6873);
and U14575 (N_14575,N_9227,N_7592);
nand U14576 (N_14576,N_9004,N_8952);
nor U14577 (N_14577,N_7437,N_6060);
nand U14578 (N_14578,N_9922,N_9309);
nand U14579 (N_14579,N_9593,N_5255);
xor U14580 (N_14580,N_9103,N_6383);
or U14581 (N_14581,N_8632,N_6378);
xor U14582 (N_14582,N_6606,N_8443);
xnor U14583 (N_14583,N_6579,N_9634);
and U14584 (N_14584,N_8755,N_5014);
xnor U14585 (N_14585,N_8262,N_6441);
xnor U14586 (N_14586,N_6675,N_8986);
and U14587 (N_14587,N_5244,N_6764);
or U14588 (N_14588,N_7762,N_7517);
and U14589 (N_14589,N_6523,N_6970);
and U14590 (N_14590,N_9557,N_7792);
nor U14591 (N_14591,N_7227,N_5451);
and U14592 (N_14592,N_7051,N_6692);
nor U14593 (N_14593,N_6681,N_8521);
nand U14594 (N_14594,N_9108,N_7667);
or U14595 (N_14595,N_9464,N_8217);
nor U14596 (N_14596,N_7192,N_6042);
and U14597 (N_14597,N_5360,N_9765);
nand U14598 (N_14598,N_6143,N_9378);
xor U14599 (N_14599,N_7525,N_6117);
or U14600 (N_14600,N_5569,N_5915);
xor U14601 (N_14601,N_6786,N_8005);
xnor U14602 (N_14602,N_8756,N_6907);
and U14603 (N_14603,N_8380,N_7565);
nand U14604 (N_14604,N_5801,N_6876);
xnor U14605 (N_14605,N_9576,N_9712);
or U14606 (N_14606,N_7124,N_9405);
xor U14607 (N_14607,N_5276,N_5949);
and U14608 (N_14608,N_7137,N_8942);
and U14609 (N_14609,N_9107,N_8808);
or U14610 (N_14610,N_6962,N_8885);
nand U14611 (N_14611,N_8007,N_6014);
and U14612 (N_14612,N_9489,N_6850);
nand U14613 (N_14613,N_6202,N_5660);
and U14614 (N_14614,N_8876,N_7692);
and U14615 (N_14615,N_7914,N_6020);
xor U14616 (N_14616,N_6161,N_7361);
nand U14617 (N_14617,N_8934,N_6153);
nand U14618 (N_14618,N_7686,N_6887);
xnor U14619 (N_14619,N_9504,N_9980);
nand U14620 (N_14620,N_7422,N_7525);
nor U14621 (N_14621,N_6671,N_9180);
or U14622 (N_14622,N_7881,N_5150);
and U14623 (N_14623,N_7518,N_6246);
nand U14624 (N_14624,N_7472,N_9173);
and U14625 (N_14625,N_8288,N_7295);
and U14626 (N_14626,N_8817,N_9342);
xnor U14627 (N_14627,N_5147,N_8689);
nand U14628 (N_14628,N_8095,N_8323);
xor U14629 (N_14629,N_7484,N_8995);
or U14630 (N_14630,N_7216,N_6249);
nor U14631 (N_14631,N_9316,N_5001);
xnor U14632 (N_14632,N_9452,N_6570);
and U14633 (N_14633,N_5982,N_7467);
nor U14634 (N_14634,N_7298,N_8431);
or U14635 (N_14635,N_7950,N_5357);
xor U14636 (N_14636,N_6001,N_7694);
or U14637 (N_14637,N_6318,N_8706);
xor U14638 (N_14638,N_8698,N_9752);
or U14639 (N_14639,N_5068,N_9784);
xnor U14640 (N_14640,N_5988,N_9013);
or U14641 (N_14641,N_5793,N_9614);
nand U14642 (N_14642,N_6172,N_9651);
and U14643 (N_14643,N_8390,N_5902);
nor U14644 (N_14644,N_9884,N_5521);
or U14645 (N_14645,N_6153,N_9673);
and U14646 (N_14646,N_7180,N_7473);
or U14647 (N_14647,N_9702,N_9073);
nand U14648 (N_14648,N_6054,N_9417);
xor U14649 (N_14649,N_9358,N_7644);
nor U14650 (N_14650,N_6444,N_7797);
nor U14651 (N_14651,N_9815,N_7100);
nor U14652 (N_14652,N_9614,N_5973);
nand U14653 (N_14653,N_6963,N_6428);
nand U14654 (N_14654,N_8029,N_9300);
or U14655 (N_14655,N_6816,N_8355);
or U14656 (N_14656,N_9218,N_7335);
nand U14657 (N_14657,N_5066,N_8098);
nor U14658 (N_14658,N_7846,N_8327);
or U14659 (N_14659,N_9039,N_6807);
nor U14660 (N_14660,N_8440,N_5888);
nor U14661 (N_14661,N_6415,N_5841);
xor U14662 (N_14662,N_9294,N_5825);
nand U14663 (N_14663,N_7008,N_5268);
nand U14664 (N_14664,N_5850,N_6207);
or U14665 (N_14665,N_5250,N_9995);
nand U14666 (N_14666,N_6949,N_8717);
and U14667 (N_14667,N_6802,N_6719);
or U14668 (N_14668,N_8837,N_7148);
and U14669 (N_14669,N_7968,N_6040);
or U14670 (N_14670,N_9726,N_6176);
nand U14671 (N_14671,N_5417,N_9298);
xor U14672 (N_14672,N_5227,N_8268);
and U14673 (N_14673,N_7513,N_9460);
or U14674 (N_14674,N_5615,N_5202);
nor U14675 (N_14675,N_7605,N_5331);
xor U14676 (N_14676,N_8045,N_6124);
xnor U14677 (N_14677,N_7418,N_6670);
or U14678 (N_14678,N_8846,N_5455);
and U14679 (N_14679,N_6002,N_6718);
xnor U14680 (N_14680,N_8306,N_5349);
nor U14681 (N_14681,N_6827,N_6430);
nand U14682 (N_14682,N_7799,N_7676);
nor U14683 (N_14683,N_8110,N_8781);
nand U14684 (N_14684,N_8084,N_9868);
and U14685 (N_14685,N_8994,N_7214);
nand U14686 (N_14686,N_6422,N_7533);
nand U14687 (N_14687,N_5161,N_5037);
nor U14688 (N_14688,N_6959,N_7635);
nand U14689 (N_14689,N_9770,N_7175);
nand U14690 (N_14690,N_8185,N_5537);
nor U14691 (N_14691,N_7423,N_6438);
nor U14692 (N_14692,N_8341,N_8315);
or U14693 (N_14693,N_7886,N_8446);
xor U14694 (N_14694,N_5136,N_9084);
nor U14695 (N_14695,N_9536,N_7400);
or U14696 (N_14696,N_6505,N_5912);
nor U14697 (N_14697,N_5199,N_7783);
xor U14698 (N_14698,N_7715,N_7668);
nor U14699 (N_14699,N_7985,N_9552);
nand U14700 (N_14700,N_9669,N_9530);
or U14701 (N_14701,N_7080,N_6808);
and U14702 (N_14702,N_8229,N_8031);
or U14703 (N_14703,N_6025,N_8171);
xor U14704 (N_14704,N_8863,N_9196);
and U14705 (N_14705,N_5019,N_8661);
nor U14706 (N_14706,N_8517,N_8070);
nand U14707 (N_14707,N_6651,N_9230);
nor U14708 (N_14708,N_6254,N_9834);
nand U14709 (N_14709,N_7899,N_7563);
xor U14710 (N_14710,N_5894,N_7853);
nand U14711 (N_14711,N_8162,N_6471);
or U14712 (N_14712,N_6539,N_7893);
nand U14713 (N_14713,N_6537,N_8475);
and U14714 (N_14714,N_7520,N_9679);
and U14715 (N_14715,N_8995,N_8756);
nor U14716 (N_14716,N_6802,N_6098);
and U14717 (N_14717,N_6578,N_7024);
nor U14718 (N_14718,N_9559,N_6637);
nor U14719 (N_14719,N_6289,N_7849);
nor U14720 (N_14720,N_7611,N_7583);
nand U14721 (N_14721,N_5628,N_7644);
xor U14722 (N_14722,N_9066,N_6981);
xor U14723 (N_14723,N_7654,N_8839);
nor U14724 (N_14724,N_7134,N_8807);
nand U14725 (N_14725,N_9462,N_8624);
or U14726 (N_14726,N_9721,N_8821);
nand U14727 (N_14727,N_9961,N_6562);
nand U14728 (N_14728,N_7359,N_8857);
xnor U14729 (N_14729,N_9763,N_5314);
nor U14730 (N_14730,N_6563,N_7171);
nor U14731 (N_14731,N_6274,N_9570);
or U14732 (N_14732,N_8535,N_6629);
and U14733 (N_14733,N_5423,N_8190);
or U14734 (N_14734,N_9866,N_5215);
and U14735 (N_14735,N_9680,N_9247);
or U14736 (N_14736,N_9365,N_8954);
or U14737 (N_14737,N_5483,N_5718);
nand U14738 (N_14738,N_5084,N_9487);
nor U14739 (N_14739,N_6853,N_9788);
nor U14740 (N_14740,N_6617,N_7065);
xnor U14741 (N_14741,N_8192,N_7093);
nand U14742 (N_14742,N_8795,N_9108);
or U14743 (N_14743,N_5337,N_6980);
nor U14744 (N_14744,N_8240,N_8134);
nand U14745 (N_14745,N_9367,N_8832);
and U14746 (N_14746,N_7402,N_8213);
and U14747 (N_14747,N_7342,N_7997);
or U14748 (N_14748,N_6957,N_9593);
nand U14749 (N_14749,N_7105,N_6194);
and U14750 (N_14750,N_8401,N_5944);
nand U14751 (N_14751,N_7016,N_8747);
or U14752 (N_14752,N_7691,N_6287);
nor U14753 (N_14753,N_8235,N_9774);
nor U14754 (N_14754,N_6475,N_9660);
xnor U14755 (N_14755,N_8988,N_5223);
and U14756 (N_14756,N_9806,N_9824);
xnor U14757 (N_14757,N_8292,N_9207);
and U14758 (N_14758,N_7763,N_6405);
or U14759 (N_14759,N_7547,N_6032);
nand U14760 (N_14760,N_6065,N_6792);
xnor U14761 (N_14761,N_8682,N_5923);
or U14762 (N_14762,N_9133,N_7641);
and U14763 (N_14763,N_8632,N_9019);
nor U14764 (N_14764,N_6136,N_6240);
nand U14765 (N_14765,N_6111,N_8678);
or U14766 (N_14766,N_8356,N_7281);
nand U14767 (N_14767,N_6070,N_9525);
xnor U14768 (N_14768,N_6979,N_7561);
and U14769 (N_14769,N_5559,N_6595);
or U14770 (N_14770,N_9617,N_6365);
or U14771 (N_14771,N_6673,N_8786);
xor U14772 (N_14772,N_6207,N_7120);
and U14773 (N_14773,N_8455,N_7217);
and U14774 (N_14774,N_7333,N_7254);
nand U14775 (N_14775,N_6431,N_6125);
nand U14776 (N_14776,N_8160,N_6859);
or U14777 (N_14777,N_5937,N_5371);
and U14778 (N_14778,N_6904,N_6434);
xnor U14779 (N_14779,N_6314,N_7213);
nor U14780 (N_14780,N_6188,N_5881);
or U14781 (N_14781,N_9153,N_6557);
xnor U14782 (N_14782,N_6260,N_8104);
xor U14783 (N_14783,N_7065,N_5292);
and U14784 (N_14784,N_9856,N_8638);
nand U14785 (N_14785,N_5108,N_7134);
xor U14786 (N_14786,N_5747,N_8241);
or U14787 (N_14787,N_6870,N_9705);
nor U14788 (N_14788,N_9565,N_5029);
nor U14789 (N_14789,N_8192,N_6554);
or U14790 (N_14790,N_6893,N_5571);
or U14791 (N_14791,N_8485,N_6202);
and U14792 (N_14792,N_5529,N_8571);
nand U14793 (N_14793,N_8148,N_6820);
nor U14794 (N_14794,N_7048,N_6123);
nor U14795 (N_14795,N_7514,N_9053);
or U14796 (N_14796,N_6536,N_8712);
nand U14797 (N_14797,N_8238,N_5514);
or U14798 (N_14798,N_8703,N_9457);
nand U14799 (N_14799,N_7690,N_7972);
nand U14800 (N_14800,N_8413,N_8373);
nand U14801 (N_14801,N_8833,N_9174);
and U14802 (N_14802,N_9377,N_9517);
xnor U14803 (N_14803,N_7412,N_6426);
xor U14804 (N_14804,N_6902,N_8902);
xor U14805 (N_14805,N_7990,N_9429);
and U14806 (N_14806,N_5799,N_5620);
nand U14807 (N_14807,N_9091,N_8587);
nand U14808 (N_14808,N_6074,N_8399);
nand U14809 (N_14809,N_5396,N_6012);
or U14810 (N_14810,N_5245,N_7132);
nor U14811 (N_14811,N_8297,N_7613);
or U14812 (N_14812,N_6967,N_6985);
or U14813 (N_14813,N_7605,N_7410);
nor U14814 (N_14814,N_8508,N_6811);
and U14815 (N_14815,N_8137,N_8834);
or U14816 (N_14816,N_7751,N_6920);
nand U14817 (N_14817,N_9189,N_9540);
nor U14818 (N_14818,N_5006,N_9736);
nand U14819 (N_14819,N_5011,N_6977);
xor U14820 (N_14820,N_9596,N_6846);
xor U14821 (N_14821,N_8148,N_5806);
nand U14822 (N_14822,N_6611,N_7349);
nand U14823 (N_14823,N_5143,N_8287);
xor U14824 (N_14824,N_8457,N_7996);
xor U14825 (N_14825,N_5267,N_7180);
and U14826 (N_14826,N_9338,N_5587);
and U14827 (N_14827,N_6851,N_9045);
nor U14828 (N_14828,N_7372,N_9228);
or U14829 (N_14829,N_6794,N_9067);
or U14830 (N_14830,N_6189,N_7714);
xnor U14831 (N_14831,N_7136,N_7836);
nor U14832 (N_14832,N_5611,N_6370);
xor U14833 (N_14833,N_6312,N_8541);
and U14834 (N_14834,N_9019,N_7907);
xnor U14835 (N_14835,N_5409,N_5728);
nand U14836 (N_14836,N_9286,N_6535);
xnor U14837 (N_14837,N_5357,N_9712);
nand U14838 (N_14838,N_5186,N_9410);
or U14839 (N_14839,N_8722,N_7163);
xor U14840 (N_14840,N_7794,N_8896);
xor U14841 (N_14841,N_5885,N_6456);
nand U14842 (N_14842,N_9836,N_9980);
nor U14843 (N_14843,N_5315,N_5715);
nand U14844 (N_14844,N_9530,N_5897);
and U14845 (N_14845,N_7965,N_6308);
nand U14846 (N_14846,N_5562,N_5998);
xor U14847 (N_14847,N_8499,N_6217);
or U14848 (N_14848,N_6200,N_7401);
xnor U14849 (N_14849,N_8115,N_5262);
nor U14850 (N_14850,N_7498,N_8501);
nor U14851 (N_14851,N_5136,N_6743);
nand U14852 (N_14852,N_6373,N_9077);
and U14853 (N_14853,N_8626,N_5918);
and U14854 (N_14854,N_7568,N_5432);
and U14855 (N_14855,N_7014,N_6975);
and U14856 (N_14856,N_7852,N_8794);
nor U14857 (N_14857,N_5444,N_7035);
xnor U14858 (N_14858,N_9014,N_8604);
nor U14859 (N_14859,N_5649,N_6154);
xor U14860 (N_14860,N_6646,N_6234);
nor U14861 (N_14861,N_6763,N_9248);
xor U14862 (N_14862,N_8468,N_6246);
xor U14863 (N_14863,N_7874,N_5020);
nor U14864 (N_14864,N_8986,N_7352);
or U14865 (N_14865,N_6273,N_7115);
xnor U14866 (N_14866,N_5575,N_6491);
nor U14867 (N_14867,N_9344,N_8034);
nor U14868 (N_14868,N_6683,N_7549);
nor U14869 (N_14869,N_9411,N_9339);
and U14870 (N_14870,N_7811,N_9689);
nor U14871 (N_14871,N_7241,N_5075);
nand U14872 (N_14872,N_8345,N_5677);
or U14873 (N_14873,N_6425,N_7867);
xnor U14874 (N_14874,N_7615,N_5511);
nand U14875 (N_14875,N_5828,N_6912);
nor U14876 (N_14876,N_8325,N_7154);
xnor U14877 (N_14877,N_5344,N_6808);
nor U14878 (N_14878,N_7200,N_7818);
or U14879 (N_14879,N_6908,N_5673);
nor U14880 (N_14880,N_6248,N_9351);
and U14881 (N_14881,N_5798,N_9853);
or U14882 (N_14882,N_8985,N_5844);
or U14883 (N_14883,N_9161,N_7576);
nand U14884 (N_14884,N_8271,N_9562);
or U14885 (N_14885,N_5683,N_7597);
or U14886 (N_14886,N_8432,N_7549);
or U14887 (N_14887,N_6314,N_9588);
and U14888 (N_14888,N_7332,N_8243);
xnor U14889 (N_14889,N_7059,N_8083);
or U14890 (N_14890,N_5710,N_6426);
and U14891 (N_14891,N_5158,N_6004);
nor U14892 (N_14892,N_8540,N_5170);
nand U14893 (N_14893,N_6426,N_5962);
xnor U14894 (N_14894,N_6400,N_8167);
or U14895 (N_14895,N_6714,N_9332);
nand U14896 (N_14896,N_9242,N_9631);
xor U14897 (N_14897,N_5412,N_9270);
or U14898 (N_14898,N_7955,N_6869);
nand U14899 (N_14899,N_5646,N_6797);
nor U14900 (N_14900,N_5598,N_7981);
nor U14901 (N_14901,N_7885,N_7075);
nand U14902 (N_14902,N_7138,N_6316);
xor U14903 (N_14903,N_6446,N_6782);
nor U14904 (N_14904,N_5324,N_9779);
xnor U14905 (N_14905,N_9078,N_6879);
xor U14906 (N_14906,N_9568,N_8032);
nand U14907 (N_14907,N_6782,N_7952);
or U14908 (N_14908,N_7091,N_8056);
and U14909 (N_14909,N_9182,N_6445);
nor U14910 (N_14910,N_5857,N_9929);
nor U14911 (N_14911,N_6221,N_9114);
and U14912 (N_14912,N_6437,N_7350);
nand U14913 (N_14913,N_7510,N_7988);
or U14914 (N_14914,N_7758,N_9069);
xor U14915 (N_14915,N_7110,N_8298);
and U14916 (N_14916,N_8428,N_7077);
or U14917 (N_14917,N_9424,N_6664);
or U14918 (N_14918,N_6282,N_6279);
nor U14919 (N_14919,N_9056,N_9431);
xor U14920 (N_14920,N_9530,N_8588);
nand U14921 (N_14921,N_5446,N_9689);
xor U14922 (N_14922,N_6622,N_5979);
and U14923 (N_14923,N_7911,N_5087);
xnor U14924 (N_14924,N_9030,N_6642);
xnor U14925 (N_14925,N_7317,N_7223);
and U14926 (N_14926,N_7625,N_9505);
and U14927 (N_14927,N_9478,N_9606);
nor U14928 (N_14928,N_7698,N_9343);
nor U14929 (N_14929,N_5778,N_9059);
xnor U14930 (N_14930,N_9668,N_7186);
and U14931 (N_14931,N_7159,N_6168);
nand U14932 (N_14932,N_6306,N_8299);
or U14933 (N_14933,N_9315,N_7039);
or U14934 (N_14934,N_6555,N_6559);
xnor U14935 (N_14935,N_9898,N_6971);
nor U14936 (N_14936,N_5975,N_8724);
nor U14937 (N_14937,N_8414,N_8526);
and U14938 (N_14938,N_7671,N_8565);
or U14939 (N_14939,N_8050,N_9689);
or U14940 (N_14940,N_6537,N_7446);
nand U14941 (N_14941,N_7333,N_7656);
nor U14942 (N_14942,N_7116,N_9631);
nor U14943 (N_14943,N_8051,N_5514);
xnor U14944 (N_14944,N_7054,N_9994);
or U14945 (N_14945,N_7022,N_6069);
nor U14946 (N_14946,N_8249,N_7674);
nand U14947 (N_14947,N_5659,N_8871);
or U14948 (N_14948,N_8636,N_7196);
and U14949 (N_14949,N_5284,N_8812);
nand U14950 (N_14950,N_9959,N_9724);
or U14951 (N_14951,N_8805,N_7976);
and U14952 (N_14952,N_5736,N_9755);
or U14953 (N_14953,N_9079,N_8234);
or U14954 (N_14954,N_7573,N_7545);
xnor U14955 (N_14955,N_6101,N_8341);
nor U14956 (N_14956,N_7041,N_7774);
nand U14957 (N_14957,N_7706,N_7438);
xor U14958 (N_14958,N_9520,N_9524);
and U14959 (N_14959,N_7861,N_6201);
and U14960 (N_14960,N_6274,N_6455);
nand U14961 (N_14961,N_5502,N_9596);
and U14962 (N_14962,N_5415,N_6378);
and U14963 (N_14963,N_9704,N_7243);
or U14964 (N_14964,N_7696,N_8106);
nor U14965 (N_14965,N_6098,N_6245);
nor U14966 (N_14966,N_9719,N_8574);
xor U14967 (N_14967,N_6989,N_8537);
nor U14968 (N_14968,N_9653,N_6437);
or U14969 (N_14969,N_8887,N_6224);
xnor U14970 (N_14970,N_7857,N_9778);
nor U14971 (N_14971,N_5265,N_8607);
xor U14972 (N_14972,N_7539,N_6017);
xor U14973 (N_14973,N_9357,N_5453);
xor U14974 (N_14974,N_7385,N_6854);
nor U14975 (N_14975,N_8432,N_9992);
or U14976 (N_14976,N_5759,N_6960);
and U14977 (N_14977,N_7468,N_5699);
and U14978 (N_14978,N_8721,N_6766);
nand U14979 (N_14979,N_7935,N_9695);
or U14980 (N_14980,N_8770,N_6037);
nand U14981 (N_14981,N_7063,N_8331);
xor U14982 (N_14982,N_6391,N_6233);
or U14983 (N_14983,N_6448,N_6390);
nand U14984 (N_14984,N_9318,N_7794);
nand U14985 (N_14985,N_8912,N_9049);
nand U14986 (N_14986,N_8617,N_8006);
xnor U14987 (N_14987,N_9635,N_6207);
nand U14988 (N_14988,N_6207,N_9049);
nand U14989 (N_14989,N_7135,N_7053);
or U14990 (N_14990,N_5510,N_9381);
nor U14991 (N_14991,N_8273,N_6486);
xor U14992 (N_14992,N_7077,N_9678);
nand U14993 (N_14993,N_9400,N_8586);
xnor U14994 (N_14994,N_6925,N_9195);
and U14995 (N_14995,N_8125,N_9066);
and U14996 (N_14996,N_7304,N_8707);
and U14997 (N_14997,N_7110,N_8032);
nand U14998 (N_14998,N_6258,N_5420);
nand U14999 (N_14999,N_8422,N_5174);
or U15000 (N_15000,N_11392,N_10798);
nand U15001 (N_15001,N_12196,N_11375);
nor U15002 (N_15002,N_14476,N_12626);
or U15003 (N_15003,N_13837,N_11386);
xor U15004 (N_15004,N_10773,N_14390);
and U15005 (N_15005,N_12120,N_12886);
nor U15006 (N_15006,N_14058,N_13708);
xnor U15007 (N_15007,N_13523,N_10235);
nand U15008 (N_15008,N_13423,N_12484);
nor U15009 (N_15009,N_10608,N_12706);
nor U15010 (N_15010,N_13511,N_11132);
or U15011 (N_15011,N_12372,N_14013);
and U15012 (N_15012,N_11697,N_10119);
xor U15013 (N_15013,N_14195,N_11018);
nor U15014 (N_15014,N_10888,N_11026);
nor U15015 (N_15015,N_11755,N_13202);
or U15016 (N_15016,N_11297,N_12302);
nand U15017 (N_15017,N_12423,N_10917);
and U15018 (N_15018,N_13994,N_11658);
nor U15019 (N_15019,N_10405,N_11876);
and U15020 (N_15020,N_12123,N_11007);
and U15021 (N_15021,N_12308,N_11129);
nor U15022 (N_15022,N_14338,N_11332);
or U15023 (N_15023,N_10480,N_14630);
nand U15024 (N_15024,N_14523,N_10421);
or U15025 (N_15025,N_11793,N_13271);
and U15026 (N_15026,N_13684,N_11499);
or U15027 (N_15027,N_11929,N_11896);
nor U15028 (N_15028,N_12777,N_13910);
nand U15029 (N_15029,N_11789,N_11081);
and U15030 (N_15030,N_14499,N_12292);
or U15031 (N_15031,N_14371,N_10072);
or U15032 (N_15032,N_10971,N_11585);
or U15033 (N_15033,N_13111,N_12782);
or U15034 (N_15034,N_14242,N_12742);
nor U15035 (N_15035,N_10040,N_11781);
nand U15036 (N_15036,N_10374,N_10567);
or U15037 (N_15037,N_10981,N_10687);
nor U15038 (N_15038,N_12448,N_13235);
nor U15039 (N_15039,N_11293,N_12903);
and U15040 (N_15040,N_14652,N_14840);
or U15041 (N_15041,N_13510,N_12958);
nand U15042 (N_15042,N_12344,N_10786);
and U15043 (N_15043,N_10822,N_11477);
nor U15044 (N_15044,N_13718,N_14947);
or U15045 (N_15045,N_11150,N_11468);
xor U15046 (N_15046,N_11742,N_11837);
or U15047 (N_15047,N_11356,N_13443);
and U15048 (N_15048,N_14654,N_11899);
or U15049 (N_15049,N_13299,N_11681);
xor U15050 (N_15050,N_10781,N_10661);
xnor U15051 (N_15051,N_11811,N_10574);
nor U15052 (N_15052,N_10482,N_12208);
or U15053 (N_15053,N_13195,N_11607);
xor U15054 (N_15054,N_12470,N_10655);
xor U15055 (N_15055,N_14509,N_14387);
nand U15056 (N_15056,N_13875,N_11131);
xor U15057 (N_15057,N_13629,N_13360);
or U15058 (N_15058,N_12189,N_14177);
nand U15059 (N_15059,N_13306,N_13618);
and U15060 (N_15060,N_10027,N_11688);
xor U15061 (N_15061,N_11219,N_13258);
and U15062 (N_15062,N_12238,N_12451);
or U15063 (N_15063,N_14742,N_13373);
nor U15064 (N_15064,N_13182,N_13126);
and U15065 (N_15065,N_10400,N_12396);
nor U15066 (N_15066,N_11657,N_12354);
nand U15067 (N_15067,N_10429,N_12294);
xor U15068 (N_15068,N_14039,N_14651);
nor U15069 (N_15069,N_14196,N_11398);
or U15070 (N_15070,N_11826,N_12227);
and U15071 (N_15071,N_13642,N_14370);
xor U15072 (N_15072,N_14901,N_14855);
or U15073 (N_15073,N_12728,N_11986);
or U15074 (N_15074,N_13637,N_13246);
xnor U15075 (N_15075,N_12422,N_13931);
or U15076 (N_15076,N_14324,N_11331);
nor U15077 (N_15077,N_10023,N_14398);
and U15078 (N_15078,N_10006,N_13660);
nor U15079 (N_15079,N_10444,N_12951);
xor U15080 (N_15080,N_12299,N_13915);
and U15081 (N_15081,N_13901,N_13193);
or U15082 (N_15082,N_11539,N_11413);
xor U15083 (N_15083,N_13025,N_12268);
or U15084 (N_15084,N_10930,N_10869);
or U15085 (N_15085,N_11732,N_10675);
or U15086 (N_15086,N_14050,N_10637);
nor U15087 (N_15087,N_13526,N_12065);
or U15088 (N_15088,N_13686,N_13919);
and U15089 (N_15089,N_12289,N_10606);
or U15090 (N_15090,N_12513,N_13638);
or U15091 (N_15091,N_12855,N_12838);
nand U15092 (N_15092,N_12609,N_12824);
nor U15093 (N_15093,N_12535,N_13644);
xnor U15094 (N_15094,N_14780,N_14256);
xnor U15095 (N_15095,N_12566,N_12881);
xor U15096 (N_15096,N_12987,N_11222);
xor U15097 (N_15097,N_14986,N_13079);
nor U15098 (N_15098,N_12485,N_10752);
and U15099 (N_15099,N_13008,N_13216);
nor U15100 (N_15100,N_11576,N_11393);
nor U15101 (N_15101,N_10513,N_10819);
or U15102 (N_15102,N_10902,N_11164);
nand U15103 (N_15103,N_11261,N_14702);
and U15104 (N_15104,N_10633,N_10406);
nand U15105 (N_15105,N_12282,N_14047);
nor U15106 (N_15106,N_13154,N_11547);
or U15107 (N_15107,N_11556,N_14666);
xor U15108 (N_15108,N_10247,N_12009);
or U15109 (N_15109,N_12873,N_13856);
or U15110 (N_15110,N_12032,N_11889);
xnor U15111 (N_15111,N_11472,N_10207);
or U15112 (N_15112,N_13930,N_12935);
and U15113 (N_15113,N_13515,N_14545);
xor U15114 (N_15114,N_13279,N_13949);
or U15115 (N_15115,N_14072,N_12187);
and U15116 (N_15116,N_10468,N_14428);
nor U15117 (N_15117,N_12226,N_12370);
or U15118 (N_15118,N_13859,N_10762);
xnor U15119 (N_15119,N_12468,N_13338);
nand U15120 (N_15120,N_13018,N_11751);
nor U15121 (N_15121,N_10999,N_10282);
nand U15122 (N_15122,N_10539,N_13825);
nand U15123 (N_15123,N_10139,N_14667);
or U15124 (N_15124,N_13680,N_10208);
or U15125 (N_15125,N_10621,N_13779);
xnor U15126 (N_15126,N_10309,N_10266);
nand U15127 (N_15127,N_12870,N_11453);
or U15128 (N_15128,N_13453,N_13074);
or U15129 (N_15129,N_12042,N_14537);
nand U15130 (N_15130,N_12731,N_14410);
or U15131 (N_15131,N_13112,N_14424);
nand U15132 (N_15132,N_10760,N_13976);
and U15133 (N_15133,N_13539,N_13251);
nand U15134 (N_15134,N_13761,N_14136);
and U15135 (N_15135,N_11877,N_10367);
or U15136 (N_15136,N_12165,N_12981);
and U15137 (N_15137,N_14110,N_11652);
nor U15138 (N_15138,N_13694,N_13148);
xor U15139 (N_15139,N_11913,N_12510);
nand U15140 (N_15140,N_10018,N_13054);
nand U15141 (N_15141,N_10958,N_10636);
xnor U15142 (N_15142,N_12989,N_11725);
nor U15143 (N_15143,N_14157,N_13822);
nor U15144 (N_15144,N_12826,N_11613);
or U15145 (N_15145,N_13156,N_13816);
nor U15146 (N_15146,N_12582,N_11636);
nand U15147 (N_15147,N_14237,N_10544);
xor U15148 (N_15148,N_11945,N_10071);
xor U15149 (N_15149,N_13575,N_13044);
nor U15150 (N_15150,N_10627,N_12150);
nor U15151 (N_15151,N_11285,N_14987);
and U15152 (N_15152,N_13744,N_10431);
nor U15153 (N_15153,N_13060,N_14930);
or U15154 (N_15154,N_12457,N_12539);
nand U15155 (N_15155,N_12141,N_12964);
nand U15156 (N_15156,N_13614,N_14349);
and U15157 (N_15157,N_14734,N_12880);
nor U15158 (N_15158,N_10263,N_14323);
nor U15159 (N_15159,N_11606,N_13566);
xnor U15160 (N_15160,N_12286,N_10586);
nand U15161 (N_15161,N_14182,N_14127);
xnor U15162 (N_15162,N_10547,N_11210);
xnor U15163 (N_15163,N_14887,N_10488);
and U15164 (N_15164,N_13952,N_14123);
nand U15165 (N_15165,N_12615,N_11473);
or U15166 (N_15166,N_11241,N_12979);
or U15167 (N_15167,N_10402,N_13574);
nand U15168 (N_15168,N_12952,N_10111);
or U15169 (N_15169,N_11374,N_12041);
and U15170 (N_15170,N_10699,N_13780);
nand U15171 (N_15171,N_12489,N_13345);
nand U15172 (N_15172,N_14698,N_14151);
nor U15173 (N_15173,N_12211,N_12505);
xnor U15174 (N_15174,N_13220,N_13398);
and U15175 (N_15175,N_14041,N_12047);
nand U15176 (N_15176,N_14009,N_10115);
xnor U15177 (N_15177,N_12638,N_14315);
nand U15178 (N_15178,N_13912,N_10200);
or U15179 (N_15179,N_11816,N_12511);
nand U15180 (N_15180,N_12810,N_10164);
xnor U15181 (N_15181,N_12406,N_10479);
xor U15182 (N_15182,N_14845,N_13124);
and U15183 (N_15183,N_14462,N_14459);
nor U15184 (N_15184,N_12195,N_13966);
xnor U15185 (N_15185,N_10691,N_14191);
nand U15186 (N_15186,N_12433,N_14624);
nand U15187 (N_15187,N_12221,N_12117);
or U15188 (N_15188,N_14198,N_14068);
and U15189 (N_15189,N_13091,N_11822);
xor U15190 (N_15190,N_14895,N_10083);
and U15191 (N_15191,N_13550,N_10747);
nand U15192 (N_15192,N_14866,N_14900);
nand U15193 (N_15193,N_11451,N_13722);
xor U15194 (N_15194,N_10784,N_11237);
nand U15195 (N_15195,N_11305,N_14310);
xnor U15196 (N_15196,N_12478,N_13376);
nor U15197 (N_15197,N_13675,N_13935);
nand U15198 (N_15198,N_12658,N_11033);
or U15199 (N_15199,N_13992,N_10022);
nand U15200 (N_15200,N_10149,N_11156);
nand U15201 (N_15201,N_14430,N_10991);
xnor U15202 (N_15202,N_10649,N_13346);
or U15203 (N_15203,N_14801,N_11310);
nor U15204 (N_15204,N_13237,N_10680);
nor U15205 (N_15205,N_12254,N_14382);
nand U15206 (N_15206,N_14452,N_12711);
nor U15207 (N_15207,N_14583,N_13864);
xor U15208 (N_15208,N_10946,N_12602);
and U15209 (N_15209,N_11009,N_10327);
nand U15210 (N_15210,N_11010,N_11872);
nor U15211 (N_15211,N_11171,N_10088);
xor U15212 (N_15212,N_12106,N_14994);
and U15213 (N_15213,N_12859,N_14492);
xor U15214 (N_15214,N_14621,N_14946);
nor U15215 (N_15215,N_14373,N_12531);
xnor U15216 (N_15216,N_11296,N_10458);
or U15217 (N_15217,N_10223,N_11491);
nand U15218 (N_15218,N_11922,N_10318);
nor U15219 (N_15219,N_14273,N_13303);
xnor U15220 (N_15220,N_12960,N_10857);
nor U15221 (N_15221,N_11315,N_14915);
xnor U15222 (N_15222,N_12383,N_14216);
xnor U15223 (N_15223,N_12064,N_12417);
and U15224 (N_15224,N_13493,N_14388);
and U15225 (N_15225,N_10188,N_13666);
and U15226 (N_15226,N_12203,N_10926);
nand U15227 (N_15227,N_11013,N_13040);
nor U15228 (N_15228,N_10689,N_14000);
xnor U15229 (N_15229,N_12022,N_12143);
and U15230 (N_15230,N_10162,N_12850);
nor U15231 (N_15231,N_14961,N_11863);
xnor U15232 (N_15232,N_10683,N_12095);
or U15233 (N_15233,N_13503,N_11741);
nor U15234 (N_15234,N_14470,N_12339);
or U15235 (N_15235,N_12229,N_11645);
nand U15236 (N_15236,N_10685,N_14951);
or U15237 (N_15237,N_10166,N_11988);
and U15238 (N_15238,N_13563,N_13134);
nand U15239 (N_15239,N_10470,N_14688);
or U15240 (N_15240,N_11367,N_10171);
and U15241 (N_15241,N_13723,N_13657);
xnor U15242 (N_15242,N_14612,N_14941);
nor U15243 (N_15243,N_14079,N_13845);
xor U15244 (N_15244,N_10907,N_11181);
xnor U15245 (N_15245,N_12382,N_14678);
or U15246 (N_15246,N_11493,N_10933);
nand U15247 (N_15247,N_12581,N_13768);
xnor U15248 (N_15248,N_14362,N_13261);
nor U15249 (N_15249,N_10044,N_12699);
xnor U15250 (N_15250,N_10684,N_10693);
nor U15251 (N_15251,N_10635,N_11841);
nor U15252 (N_15252,N_14354,N_13364);
nor U15253 (N_15253,N_12893,N_10777);
nor U15254 (N_15254,N_12912,N_13399);
xnor U15255 (N_15255,N_10383,N_10451);
or U15256 (N_15256,N_14640,N_11648);
or U15257 (N_15257,N_12916,N_11707);
nor U15258 (N_15258,N_12193,N_10439);
nor U15259 (N_15259,N_10799,N_12937);
or U15260 (N_15260,N_12716,N_13129);
xnor U15261 (N_15261,N_12757,N_13142);
nor U15262 (N_15262,N_11311,N_10074);
or U15263 (N_15263,N_12201,N_13959);
nand U15264 (N_15264,N_11133,N_10825);
and U15265 (N_15265,N_11059,N_11105);
or U15266 (N_15266,N_11247,N_14687);
nor U15267 (N_15267,N_10565,N_12703);
nand U15268 (N_15268,N_13923,N_12083);
and U15269 (N_15269,N_12999,N_11731);
or U15270 (N_15270,N_11765,N_13424);
xor U15271 (N_15271,N_13161,N_12391);
xnor U15272 (N_15272,N_14201,N_10177);
or U15273 (N_15273,N_10756,N_12906);
nor U15274 (N_15274,N_10624,N_12991);
xnor U15275 (N_15275,N_14168,N_13438);
nor U15276 (N_15276,N_12385,N_14632);
nor U15277 (N_15277,N_11855,N_10913);
xor U15278 (N_15278,N_10806,N_14730);
or U15279 (N_15279,N_10733,N_10754);
or U15280 (N_15280,N_12154,N_14577);
xor U15281 (N_15281,N_13269,N_12928);
and U15282 (N_15282,N_11430,N_13710);
or U15283 (N_15283,N_14910,N_12860);
xnor U15284 (N_15284,N_13643,N_11488);
and U15285 (N_15285,N_14814,N_10920);
xor U15286 (N_15286,N_11750,N_14313);
and U15287 (N_15287,N_12016,N_12390);
or U15288 (N_15288,N_13858,N_10277);
xnor U15289 (N_15289,N_13862,N_11037);
and U15290 (N_15290,N_12879,N_11828);
or U15291 (N_15291,N_10304,N_11061);
nand U15292 (N_15292,N_12732,N_12657);
and U15293 (N_15293,N_12823,N_14350);
nor U15294 (N_15294,N_14141,N_12246);
and U15295 (N_15295,N_13445,N_13766);
xor U15296 (N_15296,N_14303,N_12670);
and U15297 (N_15297,N_12033,N_10441);
and U15298 (N_15298,N_13500,N_10978);
nor U15299 (N_15299,N_13953,N_14137);
nand U15300 (N_15300,N_11093,N_11489);
and U15301 (N_15301,N_10715,N_13184);
nor U15302 (N_15302,N_13649,N_10213);
or U15303 (N_15303,N_13712,N_11107);
nor U15304 (N_15304,N_10082,N_12895);
xor U15305 (N_15305,N_12532,N_10815);
nor U15306 (N_15306,N_11716,N_12572);
nand U15307 (N_15307,N_13247,N_14144);
nand U15308 (N_15308,N_12491,N_10990);
nor U15309 (N_15309,N_13255,N_10051);
or U15310 (N_15310,N_12147,N_11853);
xnor U15311 (N_15311,N_10548,N_14084);
nand U15312 (N_15312,N_10601,N_13372);
and U15313 (N_15313,N_14448,N_10230);
or U15314 (N_15314,N_10026,N_10343);
or U15315 (N_15315,N_10276,N_12314);
and U15316 (N_15316,N_10280,N_10738);
and U15317 (N_15317,N_10258,N_11337);
nand U15318 (N_15318,N_12082,N_10927);
nor U15319 (N_15319,N_13045,N_13808);
or U15320 (N_15320,N_10214,N_14701);
nor U15321 (N_15321,N_11938,N_13576);
and U15322 (N_15322,N_12520,N_10057);
xnor U15323 (N_15323,N_10523,N_13835);
or U15324 (N_15324,N_10005,N_12324);
xor U15325 (N_15325,N_11667,N_12668);
and U15326 (N_15326,N_10271,N_14658);
nand U15327 (N_15327,N_13565,N_11207);
nor U15328 (N_15328,N_11575,N_13022);
nor U15329 (N_15329,N_12788,N_10404);
nor U15330 (N_15330,N_10438,N_11909);
nor U15331 (N_15331,N_11683,N_14451);
or U15332 (N_15332,N_10906,N_12684);
and U15333 (N_15333,N_14083,N_13662);
nor U15334 (N_15334,N_11847,N_13996);
nor U15335 (N_15335,N_13774,N_12791);
xnor U15336 (N_15336,N_11792,N_12553);
and U15337 (N_15337,N_13149,N_14408);
nor U15338 (N_15338,N_13521,N_10724);
and U15339 (N_15339,N_11975,N_11982);
nor U15340 (N_15340,N_13738,N_10062);
nand U15341 (N_15341,N_11329,N_12522);
nand U15342 (N_15342,N_13038,N_11824);
or U15343 (N_15343,N_12963,N_10344);
or U15344 (N_15344,N_11004,N_14322);
xor U15345 (N_15345,N_12034,N_12005);
and U15346 (N_15346,N_11062,N_14538);
xor U15347 (N_15347,N_13902,N_13739);
nand U15348 (N_15348,N_14560,N_12050);
nor U15349 (N_15349,N_10135,N_11701);
nand U15350 (N_15350,N_10007,N_13650);
nand U15351 (N_15351,N_12361,N_12639);
nor U15352 (N_15352,N_10775,N_12063);
xnor U15353 (N_15353,N_14588,N_11827);
and U15354 (N_15354,N_12772,N_13089);
and U15355 (N_15355,N_11109,N_11802);
or U15356 (N_15356,N_12381,N_14858);
nand U15357 (N_15357,N_13878,N_10395);
xor U15358 (N_15358,N_10519,N_14655);
and U15359 (N_15359,N_14711,N_11362);
xnor U15360 (N_15360,N_14593,N_13681);
nand U15361 (N_15361,N_13573,N_11144);
and U15362 (N_15362,N_14106,N_14844);
xnor U15363 (N_15363,N_13366,N_10239);
and U15364 (N_15364,N_12770,N_10910);
xnor U15365 (N_15365,N_11940,N_10914);
and U15366 (N_15366,N_11000,N_14097);
nand U15367 (N_15367,N_14581,N_13733);
nand U15368 (N_15368,N_14359,N_11264);
or U15369 (N_15369,N_10332,N_14145);
or U15370 (N_15370,N_13365,N_10889);
nor U15371 (N_15371,N_10667,N_10126);
xor U15372 (N_15372,N_11813,N_11268);
nand U15373 (N_15373,N_13970,N_11608);
nor U15374 (N_15374,N_13706,N_10351);
nand U15375 (N_15375,N_11366,N_12965);
or U15376 (N_15376,N_12759,N_14914);
nand U15377 (N_15377,N_10143,N_11342);
xor U15378 (N_15378,N_13987,N_11201);
xor U15379 (N_15379,N_13551,N_10873);
and U15380 (N_15380,N_13475,N_11592);
or U15381 (N_15381,N_10851,N_11942);
and U15382 (N_15382,N_11160,N_11966);
or U15383 (N_15383,N_14890,N_12035);
nor U15384 (N_15384,N_14376,N_10833);
and U15385 (N_15385,N_11715,N_13892);
nand U15386 (N_15386,N_12142,N_11357);
xor U15387 (N_15387,N_12801,N_10887);
nor U15388 (N_15388,N_13672,N_14043);
xor U15389 (N_15389,N_12799,N_13831);
xor U15390 (N_15390,N_12377,N_13327);
nor U15391 (N_15391,N_10844,N_13478);
nand U15392 (N_15392,N_14880,N_13536);
and U15393 (N_15393,N_11275,N_11842);
or U15394 (N_15394,N_13944,N_11204);
and U15395 (N_15395,N_10363,N_12523);
or U15396 (N_15396,N_10264,N_11086);
nor U15397 (N_15397,N_10033,N_10161);
and U15398 (N_15398,N_12435,N_11687);
and U15399 (N_15399,N_12936,N_12309);
nand U15400 (N_15400,N_14319,N_12449);
or U15401 (N_15401,N_13474,N_10501);
nor U15402 (N_15402,N_13014,N_10285);
nand U15403 (N_15403,N_10493,N_11330);
xor U15404 (N_15404,N_11183,N_14609);
or U15405 (N_15405,N_14437,N_13098);
and U15406 (N_15406,N_13896,N_14515);
or U15407 (N_15407,N_10987,N_11794);
nand U15408 (N_15408,N_13685,N_14825);
and U15409 (N_15409,N_11787,N_11085);
xor U15410 (N_15410,N_13585,N_12662);
xnor U15411 (N_15411,N_10440,N_11796);
and U15412 (N_15412,N_11353,N_12183);
nor U15413 (N_15413,N_11581,N_11690);
and U15414 (N_15414,N_11005,N_14817);
xor U15415 (N_15415,N_13941,N_14815);
nor U15416 (N_15416,N_14740,N_13762);
nor U15417 (N_15417,N_14233,N_11968);
nand U15418 (N_15418,N_14007,N_11312);
and U15419 (N_15419,N_11435,N_14569);
and U15420 (N_15420,N_13753,N_13707);
and U15421 (N_15421,N_13888,N_13340);
nand U15422 (N_15422,N_14042,N_12326);
nand U15423 (N_15423,N_14952,N_10729);
or U15424 (N_15424,N_11864,N_14173);
or U15425 (N_15425,N_11269,N_13415);
xnor U15426 (N_15426,N_11996,N_13270);
nor U15427 (N_15427,N_10619,N_11812);
nand U15428 (N_15428,N_14343,N_10291);
and U15429 (N_15429,N_10995,N_11180);
xnor U15430 (N_15430,N_11424,N_12653);
nand U15431 (N_15431,N_14826,N_11051);
or U15432 (N_15432,N_10397,N_11936);
or U15433 (N_15433,N_13064,N_12817);
nand U15434 (N_15434,N_11744,N_10076);
xnor U15435 (N_15435,N_12179,N_12144);
xor U15436 (N_15436,N_12643,N_12062);
or U15437 (N_15437,N_14235,N_13209);
xor U15438 (N_15438,N_10707,N_13117);
or U15439 (N_15439,N_13505,N_13654);
xnor U15440 (N_15440,N_14415,N_12258);
or U15441 (N_15441,N_13297,N_10789);
nor U15442 (N_15442,N_12547,N_14636);
nand U15443 (N_15443,N_14119,N_11278);
or U15444 (N_15444,N_11536,N_14409);
or U15445 (N_15445,N_11932,N_13807);
or U15446 (N_15446,N_10965,N_13215);
and U15447 (N_15447,N_10384,N_10909);
nand U15448 (N_15448,N_13464,N_14602);
and U15449 (N_15449,N_13337,N_13777);
nor U15450 (N_15450,N_14328,N_12571);
nor U15451 (N_15451,N_10466,N_13602);
or U15452 (N_15452,N_14589,N_10219);
nand U15453 (N_15453,N_12669,N_12429);
nor U15454 (N_15454,N_10764,N_10357);
nand U15455 (N_15455,N_10948,N_14750);
xor U15456 (N_15456,N_10701,N_13608);
xor U15457 (N_15457,N_12729,N_10757);
nor U15458 (N_15458,N_12894,N_12833);
nor U15459 (N_15459,N_13012,N_11038);
or U15460 (N_15460,N_11660,N_10178);
nand U15461 (N_15461,N_11927,N_12461);
nand U15462 (N_15462,N_13653,N_12512);
nand U15463 (N_15463,N_10287,N_12495);
or U15464 (N_15464,N_13052,N_10763);
xnor U15465 (N_15465,N_14896,N_12934);
xnor U15466 (N_15466,N_13205,N_14715);
nand U15467 (N_15467,N_14756,N_10576);
and U15468 (N_15468,N_11773,N_13813);
and U15469 (N_15469,N_14438,N_13834);
nor U15470 (N_15470,N_11217,N_13799);
xor U15471 (N_15471,N_13242,N_12704);
nand U15472 (N_15472,N_10003,N_10510);
nor U15473 (N_15473,N_12456,N_13313);
nand U15474 (N_15474,N_10145,N_14277);
nor U15475 (N_15475,N_14197,N_13371);
nand U15476 (N_15476,N_14990,N_12092);
or U15477 (N_15477,N_13725,N_14638);
xnor U15478 (N_15478,N_14317,N_12414);
xor U15479 (N_15479,N_13924,N_12586);
and U15480 (N_15480,N_14575,N_10896);
nand U15481 (N_15481,N_12910,N_14207);
or U15482 (N_15482,N_11244,N_11779);
or U15483 (N_15483,N_13903,N_10950);
and U15484 (N_15484,N_14999,N_13479);
nand U15485 (N_15485,N_12310,N_11380);
xor U15486 (N_15486,N_14361,N_13559);
or U15487 (N_15487,N_10108,N_14967);
and U15488 (N_15488,N_12774,N_12868);
xnor U15489 (N_15489,N_11412,N_13754);
xnor U15490 (N_15490,N_11860,N_12629);
xnor U15491 (N_15491,N_14754,N_14278);
and U15492 (N_15492,N_14641,N_12116);
and U15493 (N_15493,N_14653,N_13080);
xnor U15494 (N_15494,N_11239,N_12940);
xor U15495 (N_15495,N_11120,N_12020);
xor U15496 (N_15496,N_13818,N_11523);
xor U15497 (N_15497,N_12184,N_10472);
and U15498 (N_15498,N_11630,N_14501);
xnor U15499 (N_15499,N_10564,N_10362);
nand U15500 (N_15500,N_11558,N_11320);
xnor U15501 (N_15501,N_14179,N_12335);
nand U15502 (N_15502,N_12052,N_11843);
nand U15503 (N_15503,N_13354,N_11602);
nor U15504 (N_15504,N_12548,N_11739);
xor U15505 (N_15505,N_14767,N_14553);
and U15506 (N_15506,N_14070,N_13958);
xor U15507 (N_15507,N_14040,N_11321);
nand U15508 (N_15508,N_11987,N_10788);
nor U15509 (N_15509,N_10463,N_12129);
xor U15510 (N_15510,N_10864,N_11561);
and U15511 (N_15511,N_13490,N_10538);
nand U15512 (N_15512,N_14253,N_10521);
and U15513 (N_15513,N_12597,N_13395);
xnor U15514 (N_15514,N_14795,N_14379);
nor U15515 (N_15515,N_13636,N_14019);
nand U15516 (N_15516,N_12399,N_10376);
nor U15517 (N_15517,N_12714,N_10078);
or U15518 (N_15518,N_11359,N_13311);
nand U15519 (N_15519,N_12200,N_13187);
xnor U15520 (N_15520,N_14080,N_10678);
xnor U15521 (N_15521,N_14768,N_12792);
nand U15522 (N_15522,N_11341,N_10568);
and U15523 (N_15523,N_11090,N_13316);
nand U15524 (N_15524,N_10550,N_13452);
nor U15525 (N_15525,N_10616,N_14676);
and U15526 (N_15526,N_10620,N_14209);
xor U15527 (N_15527,N_11168,N_13887);
nor U15528 (N_15528,N_14561,N_13449);
or U15529 (N_15529,N_14166,N_11821);
nor U15530 (N_15530,N_10996,N_14366);
xnor U15531 (N_15531,N_10163,N_11372);
and U15532 (N_15532,N_10956,N_10960);
xor U15533 (N_15533,N_12002,N_11963);
xor U15534 (N_15534,N_12966,N_10221);
and U15535 (N_15535,N_10634,N_11229);
nor U15536 (N_15536,N_11888,N_13448);
or U15537 (N_15537,N_14629,N_13989);
nand U15538 (N_15538,N_11050,N_14685);
nand U15539 (N_15539,N_14506,N_14504);
or U15540 (N_15540,N_11277,N_14220);
or U15541 (N_15541,N_12865,N_13757);
nor U15542 (N_15542,N_12984,N_11919);
nand U15543 (N_15543,N_14773,N_12672);
or U15544 (N_15544,N_14139,N_11322);
xnor U15545 (N_15545,N_11256,N_12504);
nor U15546 (N_15546,N_12579,N_10793);
nor U15547 (N_15547,N_11475,N_10516);
and U15548 (N_15548,N_13389,N_13665);
nor U15549 (N_15549,N_13609,N_14126);
xor U15550 (N_15550,N_14149,N_11740);
nor U15551 (N_15551,N_13099,N_12554);
nor U15552 (N_15552,N_14018,N_12306);
or U15553 (N_15553,N_12848,N_11351);
nand U15554 (N_15554,N_12917,N_14949);
xor U15555 (N_15555,N_13592,N_10012);
xnor U15556 (N_15556,N_13732,N_13146);
and U15557 (N_15557,N_13552,N_11333);
nand U15558 (N_15558,N_14567,N_11417);
or U15559 (N_15559,N_13582,N_14114);
nand U15560 (N_15560,N_12152,N_10986);
nand U15561 (N_15561,N_10622,N_14045);
and U15562 (N_15562,N_12135,N_13874);
and U15563 (N_15563,N_11125,N_12724);
nand U15564 (N_15564,N_10443,N_10494);
xnor U15565 (N_15565,N_14697,N_13264);
nor U15566 (N_15566,N_11343,N_11231);
nor U15567 (N_15567,N_12166,N_10250);
nand U15568 (N_15568,N_12596,N_10838);
or U15569 (N_15569,N_10805,N_11846);
xnor U15570 (N_15570,N_11941,N_10205);
xnor U15571 (N_15571,N_13635,N_11578);
nand U15572 (N_15572,N_12459,N_11775);
nand U15573 (N_15573,N_13691,N_12105);
nor U15574 (N_15574,N_11483,N_12321);
nand U15575 (N_15575,N_11505,N_11067);
nor U15576 (N_15576,N_11911,N_11825);
nand U15577 (N_15577,N_11777,N_11737);
and U15578 (N_15578,N_14977,N_11918);
or U15579 (N_15579,N_14439,N_13867);
or U15580 (N_15580,N_11980,N_12705);
or U15581 (N_15581,N_10359,N_14614);
nand U15582 (N_15582,N_11895,N_11456);
nand U15583 (N_15583,N_14808,N_11024);
nand U15584 (N_15584,N_11484,N_12160);
nor U15585 (N_15585,N_12098,N_13428);
and U15586 (N_15586,N_12046,N_14998);
nand U15587 (N_15587,N_14848,N_14975);
or U15588 (N_15588,N_14378,N_12127);
or U15589 (N_15589,N_11629,N_14976);
or U15590 (N_15590,N_11957,N_10337);
and U15591 (N_15591,N_11890,N_14170);
nand U15592 (N_15592,N_14238,N_11083);
xnor U15593 (N_15593,N_10060,N_11914);
or U15594 (N_15594,N_11385,N_12194);
xor U15595 (N_15595,N_12413,N_13107);
and U15596 (N_15596,N_13606,N_14229);
nor U15597 (N_15597,N_11112,N_11962);
or U15598 (N_15598,N_13230,N_10849);
and U15599 (N_15599,N_14546,N_13849);
nor U15600 (N_15600,N_11702,N_14464);
nand U15601 (N_15601,N_11901,N_11161);
or U15602 (N_15602,N_12632,N_14076);
nand U15603 (N_15603,N_12055,N_12186);
nand U15604 (N_15604,N_13198,N_13975);
nand U15605 (N_15605,N_13743,N_12760);
and U15606 (N_15606,N_11465,N_13283);
nor U15607 (N_15607,N_13175,N_11440);
nor U15608 (N_15608,N_14029,N_13711);
xor U15609 (N_15609,N_10180,N_10647);
nor U15610 (N_15610,N_13988,N_11723);
or U15611 (N_15611,N_14781,N_11496);
nand U15612 (N_15612,N_10240,N_12175);
xor U15613 (N_15613,N_11555,N_12350);
nor U15614 (N_15614,N_13361,N_11983);
xnor U15615 (N_15615,N_13820,N_14983);
xor U15616 (N_15616,N_12618,N_10010);
nand U15617 (N_15617,N_11016,N_10238);
nand U15618 (N_15618,N_11622,N_11350);
xnor U15619 (N_15619,N_10575,N_13088);
nand U15620 (N_15620,N_13317,N_13437);
xor U15621 (N_15621,N_12407,N_11881);
or U15622 (N_15622,N_10144,N_12994);
nand U15623 (N_15623,N_11950,N_10242);
nor U15624 (N_15624,N_10209,N_14518);
and U15625 (N_15625,N_10515,N_12255);
xnor U15626 (N_15626,N_12901,N_10569);
and U15627 (N_15627,N_13023,N_11504);
or U15628 (N_15628,N_12630,N_10642);
or U15629 (N_15629,N_10054,N_14101);
nor U15630 (N_15630,N_14416,N_10121);
and U15631 (N_15631,N_13096,N_10134);
and U15632 (N_15632,N_13347,N_11509);
xnor U15633 (N_15633,N_12167,N_11313);
nand U15634 (N_15634,N_13236,N_14153);
nor U15635 (N_15635,N_12453,N_11384);
or U15636 (N_15636,N_12825,N_13153);
xor U15637 (N_15637,N_14783,N_10089);
or U15638 (N_15638,N_13262,N_10537);
nor U15639 (N_15639,N_12573,N_14514);
and U15640 (N_15640,N_13513,N_10973);
or U15641 (N_15641,N_10881,N_13291);
nand U15642 (N_15642,N_13403,N_10695);
xor U15643 (N_15643,N_11002,N_11589);
nor U15644 (N_15644,N_14790,N_12830);
or U15645 (N_15645,N_14929,N_13851);
nor U15646 (N_15646,N_13633,N_11528);
or U15647 (N_15647,N_13226,N_13554);
xor U15648 (N_15648,N_12017,N_13487);
and U15649 (N_15649,N_13778,N_12325);
xor U15650 (N_15650,N_11034,N_12739);
or U15651 (N_15651,N_11628,N_12562);
nor U15652 (N_15652,N_13720,N_14348);
nor U15653 (N_15653,N_13323,N_11830);
xor U15654 (N_15654,N_13103,N_10941);
xor U15655 (N_15655,N_10810,N_12405);
xnor U15656 (N_15656,N_11596,N_12080);
or U15657 (N_15657,N_11522,N_14854);
and U15658 (N_15658,N_11517,N_12526);
xor U15659 (N_15659,N_10029,N_12272);
xnor U15660 (N_15660,N_14661,N_12516);
and U15661 (N_15661,N_11772,N_14147);
nor U15662 (N_15662,N_13883,N_11949);
nor U15663 (N_15663,N_13804,N_11266);
xor U15664 (N_15664,N_10323,N_10049);
nand U15665 (N_15665,N_13601,N_10492);
nand U15666 (N_15666,N_11173,N_11178);
xnor U15667 (N_15667,N_12701,N_12463);
and U15668 (N_15668,N_10227,N_12988);
xor U15669 (N_15669,N_11415,N_13561);
xor U15670 (N_15670,N_12450,N_12748);
xnor U15671 (N_15671,N_12455,N_10711);
nor U15672 (N_15672,N_10787,N_13514);
nand U15673 (N_15673,N_13508,N_10929);
nand U15674 (N_15674,N_13301,N_14879);
xor U15675 (N_15675,N_12717,N_13751);
and U15676 (N_15676,N_12460,N_14098);
or U15677 (N_15677,N_11309,N_12775);
or U15678 (N_15678,N_11035,N_11800);
nor U15679 (N_15679,N_11762,N_13728);
and U15680 (N_15680,N_11437,N_10453);
and U15681 (N_15681,N_13884,N_13674);
nand U15682 (N_15682,N_14307,N_13027);
nand U15683 (N_15683,N_12931,N_11867);
and U15684 (N_15684,N_14406,N_12733);
nor U15685 (N_15685,N_14978,N_11151);
nand U15686 (N_15686,N_12389,N_14884);
and U15687 (N_15687,N_12054,N_10722);
and U15688 (N_15688,N_13932,N_11993);
xnor U15689 (N_15689,N_12665,N_10561);
xor U15690 (N_15690,N_13979,N_12056);
nor U15691 (N_15691,N_10670,N_12275);
or U15692 (N_15692,N_11703,N_11916);
and U15693 (N_15693,N_14600,N_11623);
nor U15694 (N_15694,N_13290,N_14759);
xnor U15695 (N_15695,N_11926,N_10630);
nand U15696 (N_15696,N_12343,N_10278);
and U15697 (N_15697,N_11075,N_13793);
nand U15698 (N_15698,N_11603,N_11527);
or U15699 (N_15699,N_14036,N_10413);
xnor U15700 (N_15700,N_14766,N_11220);
nand U15701 (N_15701,N_14226,N_12869);
or U15702 (N_15702,N_14477,N_14700);
or U15703 (N_15703,N_14924,N_11325);
nand U15704 (N_15704,N_10915,N_12920);
or U15705 (N_15705,N_14557,N_14245);
and U15706 (N_15706,N_14611,N_14919);
or U15707 (N_15707,N_10605,N_12752);
nand U15708 (N_15708,N_11790,N_11080);
xnor U15709 (N_15709,N_10419,N_14747);
or U15710 (N_15710,N_11196,N_12358);
nor U15711 (N_15711,N_13035,N_11840);
xor U15712 (N_15712,N_10460,N_14091);
or U15713 (N_15713,N_14936,N_10094);
nand U15714 (N_15714,N_14064,N_14731);
and U15715 (N_15715,N_11422,N_13263);
and U15716 (N_15716,N_13073,N_10713);
and U15717 (N_15717,N_13420,N_10690);
and U15718 (N_15718,N_13906,N_14507);
nor U15719 (N_15719,N_13152,N_14104);
or U15720 (N_15720,N_13197,N_13447);
nor U15721 (N_15721,N_12075,N_14931);
nor U15722 (N_15722,N_14512,N_10916);
and U15723 (N_15723,N_12472,N_11140);
or U15724 (N_15724,N_12827,N_10355);
nor U15725 (N_15725,N_10597,N_10901);
or U15726 (N_15726,N_14917,N_12436);
or U15727 (N_15727,N_14933,N_11439);
and U15728 (N_15728,N_10750,N_12871);
nand U15729 (N_15729,N_10843,N_12718);
or U15730 (N_15730,N_11521,N_12114);
nor U15731 (N_15731,N_10554,N_14035);
xnor U15732 (N_15732,N_14836,N_12188);
or U15733 (N_15733,N_14205,N_11759);
and U15734 (N_15734,N_12137,N_14057);
and U15735 (N_15735,N_12734,N_13043);
nor U15736 (N_15736,N_11545,N_10422);
and U15737 (N_15737,N_12260,N_13519);
xnor U15738 (N_15738,N_10369,N_10983);
xnor U15739 (N_15739,N_11533,N_10710);
nor U15740 (N_15740,N_12636,N_13679);
nor U15741 (N_15741,N_13570,N_10897);
nor U15742 (N_15742,N_13199,N_14832);
xor U15743 (N_15743,N_14802,N_11421);
xnor U15744 (N_15744,N_11810,N_12322);
nand U15745 (N_15745,N_14120,N_12276);
nand U15746 (N_15746,N_10095,N_11191);
nor U15747 (N_15747,N_13036,N_13544);
xor U15748 (N_15748,N_10912,N_12971);
xor U15749 (N_15749,N_11947,N_14860);
and U15750 (N_15750,N_12329,N_12228);
nor U15751 (N_15751,N_11912,N_13705);
xor U15752 (N_15752,N_12939,N_14939);
xnor U15753 (N_15753,N_10963,N_11166);
and U15754 (N_15754,N_13033,N_10342);
and U15755 (N_15755,N_10511,N_13538);
nand U15756 (N_15756,N_14922,N_10490);
nor U15757 (N_15757,N_14761,N_11236);
or U15758 (N_15758,N_13714,N_12696);
nor U15759 (N_15759,N_14033,N_11965);
and U15760 (N_15760,N_10031,N_14244);
and U15761 (N_15761,N_14082,N_10452);
and U15762 (N_15762,N_10530,N_14265);
or U15763 (N_15763,N_13410,N_10871);
nand U15764 (N_15764,N_11640,N_11363);
and U15765 (N_15765,N_11101,N_11195);
and U15766 (N_15766,N_14351,N_10640);
nor U15767 (N_15767,N_10385,N_10603);
and U15768 (N_15768,N_13309,N_13769);
nor U15769 (N_15769,N_13239,N_13071);
and U15770 (N_15770,N_11544,N_11396);
xnor U15771 (N_15771,N_10234,N_13329);
or U15772 (N_15772,N_12036,N_10955);
or U15773 (N_15773,N_11134,N_13108);
nand U15774 (N_15774,N_13477,N_14336);
nor U15775 (N_15775,N_12012,N_14794);
and U15776 (N_15776,N_12592,N_14942);
xnor U15777 (N_15777,N_10270,N_10546);
nand U15778 (N_15778,N_12296,N_10382);
nand U15779 (N_15779,N_14837,N_10317);
nor U15780 (N_15780,N_13321,N_11600);
or U15781 (N_15781,N_10281,N_12749);
nor U15782 (N_15782,N_12437,N_10542);
or U15783 (N_15783,N_12647,N_14591);
nor U15784 (N_15784,N_14703,N_14958);
and U15785 (N_15785,N_12493,N_14527);
or U15786 (N_15786,N_14656,N_13541);
xnor U15787 (N_15787,N_12404,N_12909);
or U15788 (N_15788,N_14269,N_10954);
nand U15789 (N_15789,N_12969,N_11143);
or U15790 (N_15790,N_10845,N_13363);
nor U15791 (N_15791,N_13367,N_12598);
or U15792 (N_15792,N_12536,N_12765);
and U15793 (N_15793,N_14178,N_11579);
nor U15794 (N_15794,N_14727,N_14834);
or U15795 (N_15795,N_13077,N_13426);
or U15796 (N_15796,N_13085,N_12546);
nand U15797 (N_15797,N_14142,N_14935);
nand U15798 (N_15798,N_10248,N_11757);
nor U15799 (N_15799,N_14094,N_12755);
nand U15800 (N_15800,N_13531,N_11295);
nand U15801 (N_15801,N_14012,N_11267);
nor U15802 (N_15802,N_11593,N_14525);
nor U15803 (N_15803,N_14647,N_10654);
nor U15804 (N_15804,N_14736,N_13758);
and U15805 (N_15805,N_11803,N_10063);
or U15806 (N_15806,N_10409,N_13560);
or U15807 (N_15807,N_14889,N_13225);
or U15808 (N_15808,N_14878,N_12431);
and U15809 (N_15809,N_12247,N_11611);
and U15810 (N_15810,N_10672,N_10084);
nand U15811 (N_15811,N_10096,N_12073);
and U15812 (N_15812,N_14391,N_12086);
xnor U15813 (N_15813,N_11187,N_10809);
xnor U15814 (N_15814,N_11709,N_12664);
nand U15815 (N_15815,N_13991,N_11552);
nor U15816 (N_15816,N_14934,N_11956);
nand U15817 (N_15817,N_12215,N_12069);
xor U15818 (N_15818,N_10828,N_10442);
nand U15819 (N_15819,N_14241,N_14270);
xnor U15820 (N_15820,N_13196,N_11515);
nand U15821 (N_15821,N_13177,N_14429);
nor U15822 (N_15822,N_14115,N_11141);
nand U15823 (N_15823,N_10069,N_11429);
nand U15824 (N_15824,N_14096,N_12756);
or U15825 (N_15825,N_14240,N_10222);
nand U15826 (N_15826,N_14456,N_11203);
and U15827 (N_15827,N_14552,N_12819);
or U15828 (N_15828,N_10854,N_14871);
and U15829 (N_15829,N_11402,N_12274);
nor U15830 (N_15830,N_14472,N_13121);
and U15831 (N_15831,N_12071,N_14920);
xor U15832 (N_15832,N_14375,N_14160);
nor U15833 (N_15833,N_14729,N_14713);
nand U15834 (N_15834,N_10522,N_14670);
xnor U15835 (N_15835,N_11695,N_14916);
or U15836 (N_15836,N_10922,N_10184);
xor U15837 (N_15837,N_14927,N_14564);
nand U15838 (N_15838,N_11526,N_14176);
nor U15839 (N_15839,N_11336,N_11252);
nand U15840 (N_15840,N_11469,N_12967);
and U15841 (N_15841,N_13105,N_10604);
nand U15842 (N_15842,N_13588,N_12975);
xor U15843 (N_15843,N_12222,N_12371);
nor U15844 (N_15844,N_12060,N_14034);
nand U15845 (N_15845,N_12441,N_12171);
nand U15846 (N_15846,N_12411,N_12259);
nand U15847 (N_15847,N_11619,N_12778);
xnor U15848 (N_15848,N_11055,N_10292);
nand U15849 (N_15849,N_13530,N_14298);
nor U15850 (N_15850,N_10345,N_12692);
nand U15851 (N_15851,N_14526,N_10628);
nand U15852 (N_15852,N_14210,N_14980);
and U15853 (N_15853,N_11023,N_12605);
xor U15854 (N_15854,N_13441,N_10712);
or U15855 (N_15855,N_11272,N_14870);
nor U15856 (N_15856,N_14485,N_12678);
xor U15857 (N_15857,N_12675,N_10830);
and U15858 (N_15858,N_13512,N_10943);
nand U15859 (N_15859,N_11167,N_11177);
xor U15860 (N_15860,N_14052,N_10424);
nor U15861 (N_15861,N_12497,N_11511);
and U15862 (N_15862,N_10064,N_13009);
nand U15863 (N_15863,N_12319,N_11419);
nand U15864 (N_15864,N_13458,N_13058);
xor U15865 (N_15865,N_13048,N_11795);
or U15866 (N_15866,N_10467,N_12442);
and U15867 (N_15867,N_11653,N_12947);
or U15868 (N_15868,N_13248,N_14014);
and U15869 (N_15869,N_10185,N_13425);
or U15870 (N_15870,N_11728,N_12133);
and U15871 (N_15871,N_10949,N_11441);
or U15872 (N_15872,N_14318,N_13580);
nor U15873 (N_15873,N_12925,N_13860);
nand U15874 (N_15874,N_10590,N_11569);
and U15875 (N_15875,N_14113,N_10646);
and U15876 (N_15876,N_13159,N_10925);
and U15877 (N_15877,N_12304,N_12241);
nor U15878 (N_15878,N_11128,N_13249);
nor U15879 (N_15879,N_13136,N_13461);
nor U15880 (N_15880,N_14494,N_14116);
or U15881 (N_15881,N_10253,N_14744);
or U15882 (N_15882,N_10106,N_13529);
nand U15883 (N_15883,N_12281,N_13375);
and U15884 (N_15884,N_13100,N_11257);
nand U15885 (N_15885,N_14519,N_11327);
nand U15886 (N_15886,N_13164,N_13432);
xor U15887 (N_15887,N_12483,N_13362);
or U15888 (N_15888,N_13534,N_14227);
or U15889 (N_15889,N_10761,N_14056);
and U15890 (N_15890,N_12543,N_12003);
and U15891 (N_15891,N_13929,N_12872);
xnor U15892 (N_15892,N_11891,N_14888);
nor U15893 (N_15893,N_14957,N_10485);
and U15894 (N_15894,N_10335,N_12445);
or U15895 (N_15895,N_11130,N_13776);
or U15896 (N_15896,N_12191,N_11292);
xnor U15897 (N_15897,N_11232,N_11369);
xor U15898 (N_15898,N_14665,N_14066);
and U15899 (N_15899,N_12233,N_12156);
xnor U15900 (N_15900,N_14230,N_10137);
nand U15901 (N_15901,N_11099,N_11524);
or U15902 (N_15902,N_11011,N_12168);
nand U15903 (N_15903,N_12576,N_14522);
xnor U15904 (N_15904,N_10150,N_10610);
and U15905 (N_15905,N_10032,N_11079);
xor U15906 (N_15906,N_14516,N_13188);
and U15907 (N_15907,N_11717,N_12307);
or U15908 (N_15908,N_13557,N_11387);
nand U15909 (N_15909,N_12763,N_11635);
or U15910 (N_15910,N_14105,N_11019);
or U15911 (N_15911,N_10462,N_13517);
or U15912 (N_15912,N_12138,N_10269);
nand U15913 (N_15913,N_14148,N_14635);
or U15914 (N_15914,N_14363,N_13599);
and U15915 (N_15915,N_13781,N_11442);
xor U15916 (N_15916,N_14484,N_12575);
xor U15917 (N_15917,N_13522,N_14962);
or U15918 (N_15918,N_14469,N_14260);
or U15919 (N_15919,N_13046,N_11908);
and U15920 (N_15920,N_13083,N_13465);
nor U15921 (N_15921,N_11193,N_10483);
nand U15922 (N_15922,N_12420,N_12533);
nor U15923 (N_15923,N_14749,N_10540);
xor U15924 (N_15924,N_13459,N_13020);
nor U15925 (N_15925,N_10218,N_14357);
nand U15926 (N_15926,N_14407,N_10093);
nand U15927 (N_15927,N_10349,N_14211);
and U15928 (N_15928,N_13870,N_14221);
nor U15929 (N_15929,N_14586,N_13502);
xnor U15930 (N_15930,N_13972,N_14547);
or U15931 (N_15931,N_12205,N_12887);
nand U15932 (N_15932,N_11818,N_13130);
xnor U15933 (N_15933,N_13854,N_11985);
nand U15934 (N_15934,N_11878,N_12239);
xnor U15935 (N_15935,N_14473,N_13222);
and U15936 (N_15936,N_11289,N_13203);
or U15937 (N_15937,N_14811,N_10246);
or U15938 (N_15938,N_14948,N_10525);
or U15939 (N_15939,N_14460,N_13413);
xnor U15940 (N_15940,N_14886,N_14249);
and U15941 (N_15941,N_13748,N_13259);
nor U15942 (N_15942,N_11948,N_11307);
or U15943 (N_15943,N_14053,N_13368);
nor U15944 (N_15944,N_10127,N_13179);
xnor U15945 (N_15945,N_10587,N_12798);
nand U15946 (N_15946,N_11072,N_11154);
nor U15947 (N_15947,N_13756,N_14503);
nand U15948 (N_15948,N_11786,N_10879);
or U15949 (N_15949,N_12333,N_10275);
xor U15950 (N_15950,N_14596,N_12145);
nor U15951 (N_15951,N_11303,N_14997);
xor U15952 (N_15952,N_10988,N_13170);
or U15953 (N_15953,N_13165,N_13954);
nand U15954 (N_15954,N_12182,N_10599);
xor U15955 (N_15955,N_10692,N_12612);
and U15956 (N_15956,N_11286,N_10097);
nand U15957 (N_15957,N_12642,N_10566);
nand U15958 (N_15958,N_14705,N_14722);
xnor U15959 (N_15959,N_10358,N_11774);
nor U15960 (N_15960,N_13701,N_12722);
nor U15961 (N_15961,N_13980,N_13167);
and U15962 (N_15962,N_11226,N_11567);
nor U15963 (N_15963,N_13488,N_11006);
and U15964 (N_15964,N_11928,N_11584);
xor U15965 (N_15965,N_10745,N_11260);
nor U15966 (N_15966,N_14598,N_14074);
nand U15967 (N_15967,N_11328,N_11959);
nand U15968 (N_15968,N_12067,N_14925);
xor U15969 (N_15969,N_11214,N_14130);
xor U15970 (N_15970,N_12883,N_14274);
xnor U15971 (N_15971,N_10398,N_13784);
and U15972 (N_15972,N_13349,N_11283);
nor U15973 (N_15973,N_10194,N_10609);
xor U15974 (N_15974,N_13607,N_14721);
xnor U15975 (N_15975,N_13330,N_13676);
and U15976 (N_15976,N_11411,N_14449);
or U15977 (N_15977,N_14285,N_13210);
xor U15978 (N_15978,N_10884,N_10147);
or U15979 (N_15979,N_14185,N_10340);
nor U15980 (N_15980,N_14289,N_14183);
or U15981 (N_15981,N_13305,N_14342);
nand U15982 (N_15982,N_10079,N_13624);
and U15983 (N_15983,N_11202,N_11871);
nor U15984 (N_15984,N_13352,N_14234);
and U15985 (N_15985,N_10721,N_12836);
and U15986 (N_15986,N_11532,N_11745);
nor U15987 (N_15987,N_11216,N_14255);
nor U15988 (N_15988,N_11153,N_10290);
and U15989 (N_15989,N_11175,N_10972);
and U15990 (N_15990,N_13162,N_12181);
nor U15991 (N_15991,N_10940,N_14521);
nand U15992 (N_15992,N_12613,N_11651);
nand U15993 (N_15993,N_14165,N_14427);
nor U15994 (N_15994,N_12001,N_13127);
and U15995 (N_15995,N_10120,N_11447);
or U15996 (N_15996,N_13617,N_14520);
nor U15997 (N_15997,N_12583,N_12723);
or U15998 (N_15998,N_14312,N_10296);
or U15999 (N_15999,N_13377,N_10414);
and U16000 (N_16000,N_13422,N_12128);
xor U16001 (N_16001,N_12337,N_10308);
and U16002 (N_16002,N_13387,N_13639);
or U16003 (N_16003,N_12527,N_14446);
nor U16004 (N_16004,N_13116,N_14026);
nor U16005 (N_16005,N_13911,N_14161);
nor U16006 (N_16006,N_13984,N_12768);
xor U16007 (N_16007,N_14762,N_13603);
or U16008 (N_16008,N_12161,N_10878);
nor U16009 (N_16009,N_14247,N_13457);
xor U16010 (N_16010,N_10346,N_12659);
and U16011 (N_16011,N_10151,N_11814);
nand U16012 (N_16012,N_13034,N_13968);
or U16013 (N_16013,N_12248,N_14551);
and U16014 (N_16014,N_14789,N_12781);
or U16015 (N_16015,N_10716,N_11691);
and U16016 (N_16016,N_12709,N_11348);
xor U16017 (N_16017,N_12927,N_14341);
nor U16018 (N_16018,N_10759,N_11225);
or U16019 (N_16019,N_12037,N_12563);
and U16020 (N_16020,N_12375,N_12224);
nor U16021 (N_16021,N_13234,N_10976);
nand U16022 (N_16022,N_10418,N_12885);
and U16023 (N_16023,N_10997,N_11068);
and U16024 (N_16024,N_10053,N_13335);
and U16025 (N_16025,N_10212,N_10708);
nor U16026 (N_16026,N_13589,N_13041);
or U16027 (N_16027,N_12323,N_13843);
nand U16028 (N_16028,N_11454,N_12366);
nor U16029 (N_16029,N_14276,N_13749);
and U16030 (N_16030,N_13336,N_12849);
nor U16031 (N_16031,N_13274,N_10645);
xnor U16032 (N_16032,N_11124,N_14086);
and U16033 (N_16033,N_14095,N_12637);
or U16034 (N_16034,N_12185,N_14292);
or U16035 (N_16035,N_10299,N_10653);
nor U16036 (N_16036,N_10322,N_12359);
nor U16037 (N_16037,N_10411,N_11506);
nand U16038 (N_16038,N_13794,N_14291);
or U16039 (N_16039,N_14309,N_13207);
or U16040 (N_16040,N_10272,N_10176);
xnor U16041 (N_16041,N_14006,N_11710);
or U16042 (N_16042,N_14981,N_12680);
nand U16043 (N_16043,N_13946,N_10837);
nor U16044 (N_16044,N_11672,N_12068);
xor U16045 (N_16045,N_13591,N_11049);
and U16046 (N_16046,N_10663,N_14777);
and U16047 (N_16047,N_13451,N_13118);
and U16048 (N_16048,N_13855,N_10210);
or U16049 (N_16049,N_10228,N_10450);
xnor U16050 (N_16050,N_14748,N_11060);
xor U16051 (N_16051,N_10136,N_14765);
and U16052 (N_16052,N_12506,N_10232);
and U16053 (N_16053,N_13324,N_12574);
and U16054 (N_16054,N_13548,N_12891);
or U16055 (N_16055,N_12387,N_10593);
xnor U16056 (N_16056,N_12301,N_14544);
nand U16057 (N_16057,N_14965,N_14380);
xnor U16058 (N_16058,N_10004,N_10551);
nand U16059 (N_16059,N_10428,N_11678);
nor U16060 (N_16060,N_14490,N_14737);
nor U16061 (N_16061,N_12283,N_13087);
or U16062 (N_16062,N_12393,N_12689);
nor U16063 (N_16063,N_13905,N_12856);
or U16064 (N_16064,N_13891,N_13584);
or U16065 (N_16065,N_11563,N_14436);
or U16066 (N_16066,N_13257,N_14660);
xnor U16067 (N_16067,N_11146,N_11460);
or U16068 (N_16068,N_10391,N_11599);
and U16069 (N_16069,N_14372,N_11228);
xnor U16070 (N_16070,N_11729,N_13682);
xor U16071 (N_16071,N_11615,N_12822);
nand U16072 (N_16072,N_14392,N_14955);
nand U16073 (N_16073,N_13240,N_10899);
and U16074 (N_16074,N_13914,N_10961);
nand U16075 (N_16075,N_13898,N_10900);
nand U16076 (N_16076,N_14798,N_11215);
xnor U16077 (N_16077,N_13282,N_13070);
xor U16078 (N_16078,N_10736,N_13620);
or U16079 (N_16079,N_14625,N_11092);
or U16080 (N_16080,N_13651,N_12986);
nand U16081 (N_16081,N_12726,N_10375);
nor U16082 (N_16082,N_10244,N_14550);
nand U16083 (N_16083,N_13119,N_14356);
nor U16084 (N_16084,N_11066,N_10455);
and U16085 (N_16085,N_10998,N_13933);
and U16086 (N_16086,N_14266,N_13455);
and U16087 (N_16087,N_13567,N_14818);
and U16088 (N_16088,N_14943,N_11408);
xnor U16089 (N_16089,N_14002,N_12110);
and U16090 (N_16090,N_11298,N_11063);
or U16091 (N_16091,N_12784,N_14708);
or U16092 (N_16092,N_11553,N_14467);
nand U16093 (N_16093,N_11643,N_12108);
and U16094 (N_16094,N_11832,N_11549);
and U16095 (N_16095,N_10725,N_13532);
and U16096 (N_16096,N_11764,N_10138);
or U16097 (N_16097,N_12905,N_10254);
or U16098 (N_16098,N_11617,N_13186);
nand U16099 (N_16099,N_11960,N_12266);
and U16100 (N_16100,N_10582,N_10588);
or U16101 (N_16101,N_13973,N_11137);
or U16102 (N_16102,N_12544,N_13397);
xor U16103 (N_16103,N_12614,N_14689);
nor U16104 (N_16104,N_10436,N_11582);
nand U16105 (N_16105,N_10100,N_11700);
xnor U16106 (N_16106,N_12261,N_14723);
or U16107 (N_16107,N_11588,N_11121);
nor U16108 (N_16108,N_12236,N_11094);
and U16109 (N_16109,N_13571,N_10812);
and U16110 (N_16110,N_12595,N_14623);
nor U16111 (N_16111,N_11763,N_10034);
nor U16112 (N_16112,N_14769,N_14993);
nor U16113 (N_16113,N_10334,N_12089);
and U16114 (N_16114,N_10652,N_14724);
or U16115 (N_16115,N_10489,N_12503);
and U16116 (N_16116,N_14985,N_14495);
xnor U16117 (N_16117,N_13414,N_14180);
and U16118 (N_16118,N_14434,N_10437);
and U16119 (N_16119,N_11915,N_13590);
nor U16120 (N_16120,N_14192,N_14824);
and U16121 (N_16121,N_13059,N_12834);
or U16122 (N_16122,N_14297,N_12346);
or U16123 (N_16123,N_13265,N_14782);
or U16124 (N_16124,N_11903,N_10648);
nor U16125 (N_16125,N_11087,N_12367);
nand U16126 (N_16126,N_13664,N_11807);
nand U16127 (N_16127,N_14953,N_13577);
or U16128 (N_16128,N_14710,N_13407);
and U16129 (N_16129,N_10779,N_12434);
and U16130 (N_16130,N_10356,N_11017);
nand U16131 (N_16131,N_11179,N_14530);
and U16132 (N_16132,N_10774,N_13764);
xnor U16133 (N_16133,N_10928,N_10937);
xor U16134 (N_16134,N_11609,N_11438);
nand U16135 (N_16135,N_10688,N_11481);
and U16136 (N_16136,N_14597,N_12832);
and U16137 (N_16137,N_10016,N_13429);
nand U16138 (N_16138,N_10874,N_11753);
or U16139 (N_16139,N_10201,N_11371);
xnor U16140 (N_16140,N_14664,N_14709);
xor U16141 (N_16141,N_11866,N_12348);
and U16142 (N_16142,N_11937,N_14619);
or U16143 (N_16143,N_13871,N_14534);
nor U16144 (N_16144,N_12474,N_10796);
nor U16145 (N_16145,N_14048,N_12443);
and U16146 (N_16146,N_12029,N_12776);
and U16147 (N_16147,N_12681,N_13024);
and U16148 (N_16148,N_11809,N_14496);
nand U16149 (N_16149,N_12623,N_10297);
and U16150 (N_16150,N_14374,N_10107);
xor U16151 (N_16151,N_12746,N_13621);
xnor U16152 (N_16152,N_13470,N_12519);
or U16153 (N_16153,N_10643,N_14212);
or U16154 (N_16154,N_13595,N_13547);
nor U16155 (N_16155,N_13320,N_12290);
and U16156 (N_16156,N_14992,N_12685);
xor U16157 (N_16157,N_14944,N_12844);
nor U16158 (N_16158,N_10251,N_13863);
xor U16159 (N_16159,N_14764,N_13102);
xor U16160 (N_16160,N_12192,N_13504);
and U16161 (N_16161,N_11147,N_14268);
or U16162 (N_16162,N_12458,N_12839);
nand U16163 (N_16163,N_14046,N_13402);
nand U16164 (N_16164,N_10694,N_12898);
nor U16165 (N_16165,N_12769,N_12197);
nand U16166 (N_16166,N_12218,N_11471);
nand U16167 (N_16167,N_14251,N_12753);
xnor U16168 (N_16168,N_10841,N_12688);
nor U16169 (N_16169,N_10245,N_12993);
xor U16170 (N_16170,N_11339,N_10333);
xor U16171 (N_16171,N_12923,N_10481);
or U16172 (N_16172,N_10305,N_13208);
xnor U16173 (N_16173,N_14617,N_11944);
and U16174 (N_16174,N_10430,N_14038);
nor U16175 (N_16175,N_10331,N_11730);
and U16176 (N_16176,N_10737,N_13628);
nand U16177 (N_16177,N_10050,N_12245);
nand U16178 (N_16178,N_11907,N_11665);
nor U16179 (N_16179,N_14991,N_14457);
nor U16180 (N_16180,N_14087,N_11967);
xnor U16181 (N_16181,N_13409,N_10967);
and U16182 (N_16182,N_14846,N_12518);
or U16183 (N_16183,N_13907,N_10705);
and U16184 (N_16184,N_10703,N_10199);
nor U16185 (N_16185,N_14584,N_11254);
nand U16186 (N_16186,N_12252,N_11302);
xnor U16187 (N_16187,N_12297,N_10935);
and U16188 (N_16188,N_10908,N_10128);
and U16189 (N_16189,N_11610,N_13605);
xor U16190 (N_16190,N_11512,N_14109);
or U16191 (N_16191,N_10478,N_13527);
and U16192 (N_16192,N_11030,N_12976);
nand U16193 (N_16193,N_14395,N_13341);
xnor U16194 (N_16194,N_11245,N_12015);
nor U16195 (N_16195,N_12401,N_14063);
or U16196 (N_16196,N_10433,N_14851);
or U16197 (N_16197,N_11208,N_14804);
nor U16198 (N_16198,N_12112,N_13238);
and U16199 (N_16199,N_10019,N_10109);
nor U16200 (N_16200,N_14184,N_12567);
nand U16201 (N_16201,N_10260,N_13833);
nor U16202 (N_16202,N_11693,N_14140);
nand U16203 (N_16203,N_12004,N_10921);
and U16204 (N_16204,N_10066,N_12924);
and U16205 (N_16205,N_14299,N_12364);
or U16206 (N_16206,N_14563,N_12590);
nand U16207 (N_16207,N_12126,N_12795);
nand U16208 (N_16208,N_11849,N_10206);
xor U16209 (N_16209,N_12486,N_10170);
or U16210 (N_16210,N_14150,N_11383);
or U16211 (N_16211,N_13713,N_14259);
and U16212 (N_16212,N_13067,N_14912);
nor U16213 (N_16213,N_11423,N_12369);
xnor U16214 (N_16214,N_13788,N_14807);
and U16215 (N_16215,N_10686,N_13667);
xnor U16216 (N_16216,N_12076,N_11485);
xor U16217 (N_16217,N_11542,N_13063);
nor U16218 (N_16218,N_14337,N_12214);
or U16219 (N_16219,N_14011,N_11649);
and U16220 (N_16220,N_13745,N_12622);
and U16221 (N_16221,N_12627,N_13292);
and U16222 (N_16222,N_13285,N_14894);
nand U16223 (N_16223,N_14421,N_12682);
xor U16224 (N_16224,N_10030,N_13293);
or U16225 (N_16225,N_11211,N_13061);
nor U16226 (N_16226,N_10425,N_11601);
nor U16227 (N_16227,N_14686,N_14483);
xnor U16228 (N_16228,N_12040,N_12151);
and U16229 (N_16229,N_10893,N_12648);
or U16230 (N_16230,N_10744,N_13194);
nand U16231 (N_16231,N_11642,N_13796);
nor U16232 (N_16232,N_11969,N_10098);
nand U16233 (N_16233,N_12550,N_11186);
xnor U16234 (N_16234,N_10816,N_13302);
nand U16235 (N_16235,N_13838,N_14417);
nand U16236 (N_16236,N_11192,N_13110);
xnor U16237 (N_16237,N_13689,N_14345);
xor U16238 (N_16238,N_12502,N_13031);
and U16239 (N_16239,N_13823,N_12537);
and U16240 (N_16240,N_10461,N_13715);
and U16241 (N_16241,N_13936,N_11212);
and U16242 (N_16242,N_12217,N_10831);
nor U16243 (N_16243,N_13431,N_11082);
nand U16244 (N_16244,N_10541,N_13655);
nor U16245 (N_16245,N_12787,N_11184);
xor U16246 (N_16246,N_13704,N_12852);
nor U16247 (N_16247,N_10361,N_11288);
nand U16248 (N_16248,N_10600,N_12962);
nor U16249 (N_16249,N_12634,N_10080);
or U16250 (N_16250,N_10225,N_14683);
nor U16251 (N_16251,N_14017,N_14725);
and U16252 (N_16252,N_10168,N_12588);
or U16253 (N_16253,N_12340,N_13047);
and U16254 (N_16254,N_11754,N_12889);
xor U16255 (N_16255,N_12243,N_12313);
xor U16256 (N_16256,N_10840,N_10310);
xor U16257 (N_16257,N_12911,N_11271);
xnor U16258 (N_16258,N_10339,N_11284);
nand U16259 (N_16259,N_14628,N_10497);
and U16260 (N_16260,N_12424,N_10380);
and U16261 (N_16261,N_11098,N_11897);
or U16262 (N_16262,N_13019,N_10193);
nor U16263 (N_16263,N_14284,N_10289);
or U16264 (N_16264,N_13692,N_14394);
nand U16265 (N_16265,N_11364,N_11259);
and U16266 (N_16266,N_11381,N_10778);
xor U16267 (N_16267,N_10038,N_12589);
xnor U16268 (N_16268,N_11498,N_14704);
xor U16269 (N_16269,N_13760,N_13339);
nand U16270 (N_16270,N_12426,N_12534);
or U16271 (N_16271,N_11494,N_12101);
or U16272 (N_16272,N_12521,N_10969);
nor U16273 (N_16273,N_14488,N_14797);
xor U16274 (N_16274,N_10632,N_11282);
nor U16275 (N_16275,N_11159,N_11486);
nor U16276 (N_16276,N_14536,N_10379);
nor U16277 (N_16277,N_12300,N_12454);
nor U16278 (N_16278,N_12694,N_14236);
nor U16279 (N_16279,N_10826,N_11537);
nor U16280 (N_16280,N_10252,N_13999);
xor U16281 (N_16281,N_13233,N_10353);
or U16282 (N_16282,N_14022,N_11427);
xnor U16283 (N_16283,N_14796,N_12113);
nor U16284 (N_16284,N_13801,N_13206);
xnor U16285 (N_16285,N_10449,N_13333);
or U16286 (N_16286,N_10052,N_13746);
xnor U16287 (N_16287,N_10832,N_14208);
nor U16288 (N_16288,N_13383,N_13056);
or U16289 (N_16289,N_13934,N_10782);
or U16290 (N_16290,N_11377,N_14326);
nand U16291 (N_16291,N_11894,N_12061);
nand U16292 (N_16292,N_10563,N_11198);
and U16293 (N_16293,N_12180,N_11463);
xor U16294 (N_16294,N_11508,N_13955);
or U16295 (N_16295,N_13440,N_13583);
and U16296 (N_16296,N_13357,N_14695);
nor U16297 (N_16297,N_14314,N_10571);
nor U16298 (N_16298,N_12481,N_12416);
xor U16299 (N_16299,N_12149,N_14639);
or U16300 (N_16300,N_11152,N_13600);
and U16301 (N_16301,N_10427,N_11249);
and U16302 (N_16302,N_11587,N_11979);
nand U16303 (N_16303,N_11559,N_14960);
xnor U16304 (N_16304,N_13696,N_14906);
and U16305 (N_16305,N_11981,N_12851);
or U16306 (N_16306,N_11573,N_12710);
nor U16307 (N_16307,N_14707,N_11668);
nand U16308 (N_16308,N_11248,N_11931);
nand U16309 (N_16309,N_10202,N_13497);
nand U16310 (N_16310,N_10035,N_14169);
nand U16311 (N_16311,N_13374,N_12978);
or U16312 (N_16312,N_11084,N_14092);
and U16313 (N_16313,N_11586,N_10502);
nor U16314 (N_16314,N_11597,N_10804);
nand U16315 (N_16315,N_13631,N_14330);
or U16316 (N_16316,N_13937,N_14732);
or U16317 (N_16317,N_13332,N_13861);
and U16318 (N_16318,N_11713,N_12861);
xor U16319 (N_16319,N_14893,N_14202);
xor U16320 (N_16320,N_10865,N_13252);
nand U16321 (N_16321,N_12480,N_12628);
or U16322 (N_16322,N_10811,N_11263);
or U16323 (N_16323,N_13412,N_11174);
nand U16324 (N_16324,N_12479,N_13581);
nand U16325 (N_16325,N_11352,N_13553);
and U16326 (N_16326,N_14248,N_11654);
or U16327 (N_16327,N_12330,N_14979);
nand U16328 (N_16328,N_11457,N_13886);
xor U16329 (N_16329,N_11319,N_12608);
nand U16330 (N_16330,N_10231,N_10148);
xnor U16331 (N_16331,N_13267,N_13123);
xor U16332 (N_16332,N_10723,N_12890);
nor U16333 (N_16333,N_13709,N_13005);
nor U16334 (N_16334,N_12365,N_10099);
nor U16335 (N_16335,N_14214,N_13113);
nor U16336 (N_16336,N_13765,N_12624);
and U16337 (N_16337,N_10953,N_12279);
nor U16338 (N_16338,N_12528,N_14690);
nand U16339 (N_16339,N_10167,N_12896);
or U16340 (N_16340,N_10860,N_11314);
or U16341 (N_16341,N_14839,N_10390);
xor U16342 (N_16342,N_12469,N_10673);
nor U16343 (N_16343,N_12649,N_14305);
nor U16344 (N_16344,N_13850,N_13865);
or U16345 (N_16345,N_12835,N_14869);
or U16346 (N_16346,N_13670,N_12477);
and U16347 (N_16347,N_13115,N_12741);
xor U16348 (N_16348,N_12432,N_12794);
xor U16349 (N_16349,N_12857,N_10146);
nand U16350 (N_16350,N_11756,N_14254);
and U16351 (N_16351,N_11379,N_11999);
or U16352 (N_16352,N_10717,N_11388);
nor U16353 (N_16353,N_12345,N_14060);
xnor U16354 (N_16354,N_12673,N_13880);
and U16355 (N_16355,N_10169,N_14133);
nor U16356 (N_16356,N_12332,N_14051);
or U16357 (N_16357,N_14607,N_11605);
xnor U16358 (N_16358,N_10945,N_11104);
xnor U16359 (N_16359,N_10267,N_14938);
nand U16360 (N_16360,N_12267,N_13401);
xor U16361 (N_16361,N_11743,N_11028);
xor U16362 (N_16362,N_13817,N_10536);
nor U16363 (N_16363,N_11974,N_14859);
nor U16364 (N_16364,N_12049,N_13729);
nand U16365 (N_16365,N_12633,N_10882);
nand U16366 (N_16366,N_12646,N_11831);
xor U16367 (N_16367,N_13671,N_12109);
and U16368 (N_16368,N_12545,N_12900);
and U16369 (N_16369,N_11784,N_14358);
xor U16370 (N_16370,N_10500,N_11414);
nor U16371 (N_16371,N_13922,N_12652);
or U16372 (N_16372,N_13382,N_10257);
xor U16373 (N_16373,N_13543,N_11780);
nor U16374 (N_16374,N_10249,N_13229);
and U16375 (N_16375,N_14847,N_14720);
and U16376 (N_16376,N_11834,N_11326);
xnor U16377 (N_16377,N_14044,N_13520);
or U16378 (N_16378,N_11058,N_11022);
or U16379 (N_16379,N_11924,N_11925);
xnor U16380 (N_16380,N_14078,N_14918);
and U16381 (N_16381,N_14644,N_13775);
xnor U16382 (N_16382,N_14121,N_13759);
xor U16383 (N_16383,N_14015,N_14604);
and U16384 (N_16384,N_14419,N_12148);
nand U16385 (N_16385,N_11291,N_11923);
xnor U16386 (N_16386,N_12542,N_11998);
nor U16387 (N_16387,N_14118,N_11012);
xor U16388 (N_16388,N_10298,N_13138);
and U16389 (N_16389,N_11835,N_11360);
and U16390 (N_16390,N_13829,N_13169);
xor U16391 (N_16391,N_11036,N_12140);
nand U16392 (N_16392,N_10664,N_10217);
or U16393 (N_16393,N_14805,N_10780);
and U16394 (N_16394,N_11875,N_12285);
nor U16395 (N_16395,N_11276,N_10730);
and U16396 (N_16396,N_11952,N_12078);
nand U16397 (N_16397,N_13558,N_12780);
xnor U16398 (N_16398,N_14486,N_12708);
and U16399 (N_16399,N_10158,N_11815);
and U16400 (N_16400,N_10839,N_10102);
or U16401 (N_16401,N_13030,N_11238);
xor U16402 (N_16402,N_13663,N_13180);
and U16403 (N_16403,N_12244,N_13750);
xnor U16404 (N_16404,N_10677,N_10765);
xor U16405 (N_16405,N_13010,N_11870);
or U16406 (N_16406,N_12269,N_14365);
and U16407 (N_16407,N_12957,N_10347);
and U16408 (N_16408,N_12515,N_11224);
or U16409 (N_16409,N_11290,N_13528);
nand U16410 (N_16410,N_12230,N_10682);
nand U16411 (N_16411,N_14543,N_10306);
or U16412 (N_16412,N_12000,N_14673);
and U16413 (N_16413,N_14443,N_13647);
and U16414 (N_16414,N_13542,N_11287);
or U16415 (N_16415,N_13882,N_12271);
nor U16416 (N_16416,N_12316,N_12496);
xor U16417 (N_16417,N_13741,N_12525);
or U16418 (N_16418,N_13231,N_12730);
and U16419 (N_16419,N_12607,N_10434);
and U16420 (N_16420,N_10518,N_13114);
xor U16421 (N_16421,N_13218,N_12096);
and U16422 (N_16422,N_10014,N_14649);
nand U16423 (N_16423,N_10446,N_12341);
xor U16424 (N_16424,N_11088,N_13795);
xnor U16425 (N_16425,N_14691,N_12882);
xor U16426 (N_16426,N_13957,N_14932);
nand U16427 (N_16427,N_14090,N_14841);
nor U16428 (N_16428,N_13369,N_13844);
nand U16429 (N_16429,N_11616,N_13806);
xnor U16430 (N_16430,N_14134,N_14065);
xor U16431 (N_16431,N_11091,N_13125);
or U16432 (N_16432,N_10553,N_13384);
nand U16433 (N_16433,N_14921,N_10191);
xor U16434 (N_16434,N_10898,N_13518);
and U16435 (N_16435,N_11699,N_12691);
xor U16436 (N_16436,N_14505,N_13462);
nand U16437 (N_16437,N_11158,N_10024);
nand U16438 (N_16438,N_12280,N_13325);
xnor U16439 (N_16439,N_11614,N_13176);
xor U16440 (N_16440,N_13466,N_13982);
xor U16441 (N_16441,N_13192,N_11738);
nor U16442 (N_16442,N_11661,N_11823);
and U16443 (N_16443,N_12921,N_13960);
and U16444 (N_16444,N_12177,N_14739);
or U16445 (N_16445,N_13260,N_11185);
or U16446 (N_16446,N_14799,N_13857);
xor U16447 (N_16447,N_12996,N_13963);
and U16448 (N_16448,N_14601,N_10265);
xnor U16449 (N_16449,N_10328,N_14217);
nand U16450 (N_16450,N_10435,N_11548);
nor U16451 (N_16451,N_14891,N_12044);
nand U16452 (N_16452,N_10204,N_13962);
nand U16453 (N_16453,N_11612,N_14788);
nor U16454 (N_16454,N_13698,N_13797);
xnor U16455 (N_16455,N_12006,N_13658);
nand U16456 (N_16456,N_10932,N_12977);
xor U16457 (N_16457,N_11748,N_10307);
xnor U16458 (N_16458,N_13158,N_12311);
nand U16459 (N_16459,N_11108,N_10122);
or U16460 (N_16460,N_14696,N_12225);
and U16461 (N_16461,N_12210,N_14028);
nor U16462 (N_16462,N_10399,N_12570);
or U16463 (N_16463,N_12464,N_11747);
or U16464 (N_16464,N_11844,N_12164);
xnor U16465 (N_16465,N_13028,N_10445);
or U16466 (N_16466,N_10658,N_13824);
xnor U16467 (N_16467,N_11014,N_13496);
nor U16468 (N_16468,N_11274,N_13082);
or U16469 (N_16469,N_11324,N_11852);
nor U16470 (N_16470,N_10613,N_13244);
or U16471 (N_16471,N_14037,N_10966);
or U16472 (N_16472,N_11455,N_10676);
nand U16473 (N_16473,N_14719,N_14215);
and U16474 (N_16474,N_14290,N_12577);
nand U16475 (N_16475,N_14637,N_13151);
xnor U16476 (N_16476,N_11705,N_14124);
nor U16477 (N_16477,N_10484,N_14386);
nand U16478 (N_16478,N_14758,N_12030);
xnor U16479 (N_16479,N_12111,N_11664);
or U16480 (N_16480,N_10962,N_12264);
or U16481 (N_16481,N_14355,N_13057);
and U16482 (N_16482,N_11106,N_13610);
nand U16483 (N_16483,N_10741,N_14088);
xor U16484 (N_16484,N_14966,N_14189);
xnor U16485 (N_16485,N_11659,N_14831);
nand U16486 (N_16486,N_13997,N_14774);
or U16487 (N_16487,N_12057,N_14699);
nand U16488 (N_16488,N_13683,N_10312);
xnor U16489 (N_16489,N_14027,N_12874);
nor U16490 (N_16490,N_13050,N_14779);
or U16491 (N_16491,N_14904,N_11136);
and U16492 (N_16492,N_10918,N_14302);
and U16493 (N_16493,N_10847,N_11639);
xor U16494 (N_16494,N_14020,N_12645);
nor U16495 (N_16495,N_10656,N_12352);
nand U16496 (N_16496,N_12351,N_13467);
nor U16497 (N_16497,N_14030,N_13348);
and U16498 (N_16498,N_14743,N_14680);
nor U16499 (N_16499,N_11804,N_13540);
nor U16500 (N_16500,N_14928,N_10036);
or U16501 (N_16501,N_12059,N_12476);
xnor U16502 (N_16502,N_12088,N_12631);
nor U16503 (N_16503,N_10477,N_12955);
nand U16504 (N_16504,N_12591,N_10140);
nand U16505 (N_16505,N_10157,N_11543);
nand U16506 (N_16506,N_10092,N_10133);
nor U16507 (N_16507,N_13981,N_10229);
xor U16508 (N_16508,N_13827,N_11206);
xor U16509 (N_16509,N_14393,N_14250);
nand U16510 (N_16510,N_14281,N_10572);
and U16511 (N_16511,N_10728,N_14555);
or U16512 (N_16512,N_14385,N_11676);
or U16513 (N_16513,N_10842,N_10589);
nand U16514 (N_16514,N_14347,N_13611);
nor U16515 (N_16515,N_14810,N_10284);
nor U16516 (N_16516,N_12494,N_14352);
or U16517 (N_16517,N_14875,N_12438);
or U16518 (N_16518,N_14684,N_13740);
and U16519 (N_16519,N_11436,N_14471);
nand U16520 (N_16520,N_13562,N_12419);
nand U16521 (N_16521,N_14970,N_13343);
or U16522 (N_16522,N_14411,N_12802);
or U16523 (N_16523,N_10262,N_11450);
xor U16524 (N_16524,N_11397,N_13893);
or U16525 (N_16525,N_14404,N_13545);
and U16526 (N_16526,N_13081,N_10381);
and U16527 (N_16527,N_14257,N_12124);
nor U16528 (N_16528,N_10591,N_13578);
or U16529 (N_16529,N_12619,N_12256);
nand U16530 (N_16530,N_14571,N_13172);
nor U16531 (N_16531,N_11917,N_13076);
or U16532 (N_16532,N_11304,N_10617);
or U16533 (N_16533,N_12773,N_11487);
and U16534 (N_16534,N_11502,N_13331);
and U16535 (N_16535,N_14458,N_11520);
xnor U16536 (N_16536,N_13418,N_13140);
nand U16537 (N_16537,N_12943,N_11935);
nand U16538 (N_16538,N_12336,N_13417);
and U16539 (N_16539,N_10393,N_14279);
or U16540 (N_16540,N_11122,N_13471);
xor U16541 (N_16541,N_14535,N_13173);
or U16542 (N_16542,N_10131,N_12974);
nor U16543 (N_16543,N_10562,N_13181);
xnor U16544 (N_16544,N_13615,N_10364);
and U16545 (N_16545,N_14016,N_13104);
nor U16546 (N_16546,N_12051,N_11760);
nor U16547 (N_16547,N_13612,N_11626);
xnor U16548 (N_16548,N_14320,N_14275);
and U16549 (N_16549,N_14396,N_10320);
nor U16550 (N_16550,N_11808,N_11409);
xor U16551 (N_16551,N_12972,N_10215);
nor U16552 (N_16552,N_13144,N_10061);
and U16553 (N_16553,N_11076,N_14763);
xor U16554 (N_16554,N_10175,N_14827);
and U16555 (N_16555,N_11410,N_11577);
nor U16556 (N_16556,N_13546,N_10037);
or U16557 (N_16557,N_13967,N_11365);
nor U16558 (N_16558,N_13141,N_12444);
and U16559 (N_16559,N_14295,N_11769);
and U16560 (N_16560,N_14294,N_12198);
nor U16561 (N_16561,N_11991,N_14186);
xor U16562 (N_16562,N_11358,N_10982);
or U16563 (N_16563,N_11650,N_11934);
xor U16564 (N_16564,N_13983,N_13640);
nor U16565 (N_16565,N_11046,N_11669);
xnor U16566 (N_16566,N_12053,N_14397);
nor U16567 (N_16567,N_12702,N_12758);
nor U16568 (N_16568,N_11299,N_14972);
xor U16569 (N_16569,N_10159,N_10216);
xor U16570 (N_16570,N_13069,N_13281);
nor U16571 (N_16571,N_13042,N_11791);
or U16572 (N_16572,N_13224,N_13731);
or U16573 (N_16573,N_12843,N_10944);
and U16574 (N_16574,N_11656,N_11720);
nand U16575 (N_16575,N_11189,N_10476);
or U16576 (N_16576,N_14809,N_14267);
and U16577 (N_16577,N_10528,N_10890);
and U16578 (N_16578,N_10524,N_13810);
nand U16579 (N_16579,N_11065,N_12091);
nor U16580 (N_16580,N_10611,N_11692);
or U16581 (N_16581,N_13494,N_12783);
or U16582 (N_16582,N_11163,N_14959);
xor U16583 (N_16583,N_12837,N_10048);
xor U16584 (N_16584,N_10301,N_14493);
xnor U16585 (N_16585,N_12915,N_10526);
or U16586 (N_16586,N_12403,N_11677);
nor U16587 (N_16587,N_11258,N_14111);
and U16588 (N_16588,N_12698,N_14399);
xnor U16589 (N_16589,N_12785,N_10372);
xnor U16590 (N_16590,N_14422,N_11188);
xnor U16591 (N_16591,N_11262,N_12530);
xor U16592 (N_16592,N_12287,N_10612);
or U16593 (N_16593,N_10432,N_12097);
and U16594 (N_16594,N_12918,N_13985);
nor U16595 (N_16595,N_12206,N_13742);
nor U16596 (N_16596,N_14874,N_14646);
and U16597 (N_16597,N_11971,N_11213);
xor U16598 (N_16598,N_14187,N_14663);
nor U16599 (N_16599,N_11097,N_11025);
nor U16600 (N_16600,N_14204,N_12427);
nand U16601 (N_16601,N_13798,N_12743);
and U16602 (N_16602,N_10073,N_11631);
nand U16603 (N_16603,N_12507,N_10527);
nand U16604 (N_16604,N_13805,N_14633);
xor U16605 (N_16605,N_11718,N_13245);
or U16606 (N_16606,N_10938,N_10514);
nor U16607 (N_16607,N_14306,N_11115);
xor U16608 (N_16608,N_14580,N_13084);
nor U16609 (N_16609,N_13147,N_10758);
nand U16610 (N_16610,N_12908,N_12007);
xnor U16611 (N_16611,N_14194,N_12440);
and U16612 (N_16612,N_11801,N_11031);
and U16613 (N_16613,N_13241,N_10341);
xnor U16614 (N_16614,N_11859,N_10447);
and U16615 (N_16615,N_14077,N_13011);
xnor U16616 (N_16616,N_13436,N_11042);
or U16617 (N_16617,N_11119,N_14728);
or U16618 (N_16618,N_14500,N_11733);
and U16619 (N_16619,N_13627,N_11354);
and U16620 (N_16620,N_10067,N_14772);
nand U16621 (N_16621,N_12394,N_11673);
xor U16622 (N_16622,N_14672,N_14502);
or U16623 (N_16623,N_14786,N_14032);
xnor U16624 (N_16624,N_11984,N_11535);
or U16625 (N_16625,N_13097,N_10977);
xor U16626 (N_16626,N_10742,N_10503);
nor U16627 (N_16627,N_14480,N_12045);
or U16628 (N_16628,N_14175,N_12808);
xnor U16629 (N_16629,N_14129,N_14107);
xor U16630 (N_16630,N_14718,N_12913);
or U16631 (N_16631,N_11771,N_12490);
or U16632 (N_16632,N_14280,N_12942);
nand U16633 (N_16633,N_12829,N_11869);
and U16634 (N_16634,N_11711,N_11958);
and U16635 (N_16635,N_13659,N_14883);
xnor U16636 (N_16636,N_12800,N_10748);
or U16637 (N_16637,N_12786,N_11406);
xnor U16638 (N_16638,N_12816,N_10880);
nand U16639 (N_16639,N_11391,N_14634);
nor U16640 (N_16640,N_11480,N_12262);
nor U16641 (N_16641,N_12253,N_12320);
nor U16642 (N_16642,N_13948,N_11253);
and U16643 (N_16643,N_12278,N_12360);
xnor U16644 (N_16644,N_13278,N_13294);
nand U16645 (N_16645,N_14054,N_12818);
or U16646 (N_16646,N_10803,N_11503);
or U16647 (N_16647,N_12676,N_12099);
nand U16648 (N_16648,N_11420,N_14674);
nand U16649 (N_16649,N_14816,N_11641);
nand U16650 (N_16650,N_14005,N_13646);
or U16651 (N_16651,N_10583,N_11221);
nor U16652 (N_16652,N_13648,N_10508);
nand U16653 (N_16653,N_13993,N_12926);
xor U16654 (N_16654,N_14131,N_12611);
or U16655 (N_16655,N_12617,N_13388);
and U16656 (N_16656,N_13379,N_13408);
nor U16657 (N_16657,N_12026,N_10696);
or U16658 (N_16658,N_14610,N_13095);
and U16659 (N_16659,N_14574,N_12594);
nand U16660 (N_16660,N_10529,N_12207);
nor U16661 (N_16661,N_13454,N_14882);
nor U16662 (N_16662,N_10877,N_14842);
and U16663 (N_16663,N_12118,N_11170);
xnor U16664 (N_16664,N_14576,N_11459);
xnor U16665 (N_16665,N_13516,N_12651);
xnor U16666 (N_16666,N_12747,N_14679);
or U16667 (N_16667,N_12713,N_13013);
xnor U16668 (N_16668,N_12933,N_10734);
nor U16669 (N_16669,N_11838,N_13956);
and U16670 (N_16670,N_13163,N_12072);
xnor U16671 (N_16671,N_11308,N_14599);
or U16672 (N_16672,N_13853,N_12250);
nand U16673 (N_16673,N_12119,N_10183);
or U16674 (N_16674,N_11500,N_12712);
or U16675 (N_16675,N_12878,N_12293);
and U16676 (N_16676,N_12568,N_13212);
nand U16677 (N_16677,N_12565,N_12767);
and U16678 (N_16678,N_14511,N_11047);
and U16679 (N_16679,N_14243,N_10863);
or U16680 (N_16680,N_13885,N_13790);
nor U16681 (N_16681,N_14529,N_10718);
nand U16682 (N_16682,N_11100,N_10124);
nand U16683 (N_16683,N_11043,N_12039);
or U16684 (N_16684,N_12650,N_11997);
xor U16685 (N_16685,N_12018,N_14746);
or U16686 (N_16686,N_13342,N_11848);
xnor U16687 (N_16687,N_12467,N_10615);
xnor U16688 (N_16688,N_10474,N_12693);
nor U16689 (N_16689,N_11666,N_14021);
nand U16690 (N_16690,N_10268,N_10091);
xor U16691 (N_16691,N_10330,N_12327);
nor U16692 (N_16692,N_14833,N_13965);
or U16693 (N_16693,N_12961,N_11323);
nand U16694 (N_16694,N_14856,N_10814);
and U16695 (N_16695,N_11155,N_10979);
and U16696 (N_16696,N_14595,N_11675);
xnor U16697 (N_16697,N_11405,N_10172);
and U16698 (N_16698,N_14631,N_11734);
and U16699 (N_16699,N_13904,N_13697);
xor U16700 (N_16700,N_11233,N_10156);
xor U16701 (N_16701,N_11845,N_10895);
nand U16702 (N_16702,N_12487,N_11003);
or U16703 (N_16703,N_11978,N_12813);
xor U16704 (N_16704,N_11990,N_12397);
and U16705 (N_16705,N_12644,N_11052);
xnor U16706 (N_16706,N_11376,N_14100);
nand U16707 (N_16707,N_13139,N_10584);
nor U16708 (N_16708,N_12103,N_10070);
or U16709 (N_16709,N_13189,N_14262);
nand U16710 (N_16710,N_11646,N_14821);
nand U16711 (N_16711,N_13998,N_14867);
nor U16712 (N_16712,N_11338,N_13396);
nand U16713 (N_16713,N_14381,N_11474);
nor U16714 (N_16714,N_13909,N_10389);
nor U16715 (N_16715,N_10824,N_10552);
nor U16716 (N_16716,N_12697,N_10086);
and U16717 (N_16717,N_13695,N_12421);
and U16718 (N_16718,N_14822,N_10087);
xnor U16719 (N_16719,N_10520,N_13356);
nand U16720 (N_16720,N_14353,N_13632);
or U16721 (N_16721,N_12985,N_14585);
nand U16722 (N_16722,N_14620,N_13256);
nand U16723 (N_16723,N_14171,N_14335);
xor U16724 (N_16724,N_13677,N_14286);
and U16725 (N_16725,N_11316,N_12740);
nand U16726 (N_16726,N_11008,N_11476);
nand U16727 (N_16727,N_10187,N_14413);
xor U16728 (N_16728,N_14712,N_11482);
xnor U16729 (N_16729,N_13921,N_12158);
xor U16730 (N_16730,N_11378,N_12779);
nand U16731 (N_16731,N_12998,N_11467);
and U16732 (N_16732,N_13007,N_12944);
and U16733 (N_16733,N_10236,N_10802);
nand U16734 (N_16734,N_10801,N_10039);
xnor U16735 (N_16735,N_10706,N_11418);
and U16736 (N_16736,N_11218,N_11501);
xnor U16737 (N_16737,N_10058,N_13204);
xnor U16738 (N_16738,N_14717,N_10401);
xnor U16739 (N_16739,N_12353,N_13273);
xor U16740 (N_16740,N_11598,N_14565);
nand U16741 (N_16741,N_10771,N_11516);
or U16742 (N_16742,N_11403,N_10794);
or U16743 (N_16743,N_11149,N_11044);
xnor U16744 (N_16744,N_14650,N_13734);
xnor U16745 (N_16745,N_10198,N_10846);
nand U16746 (N_16746,N_10261,N_13463);
and U16747 (N_16747,N_11621,N_11538);
nor U16748 (N_16748,N_11724,N_13460);
nand U16749 (N_16749,N_14099,N_13476);
nand U16750 (N_16750,N_12863,N_12616);
and U16751 (N_16751,N_10464,N_10939);
or U16752 (N_16752,N_11904,N_14885);
xor U16753 (N_16753,N_10753,N_10465);
xor U16754 (N_16754,N_12517,N_11722);
xnor U16755 (N_16755,N_13391,N_10179);
nand U16756 (N_16756,N_10665,N_14261);
nor U16757 (N_16757,N_11390,N_13812);
nand U16758 (N_16758,N_13876,N_13003);
xor U16759 (N_16759,N_14463,N_11027);
or U16760 (N_16760,N_12159,N_14897);
nand U16761 (N_16761,N_13872,N_11345);
and U16762 (N_16762,N_11873,N_12725);
xnor U16763 (N_16763,N_13174,N_12600);
xor U16764 (N_16764,N_10657,N_13877);
nand U16765 (N_16765,N_14193,N_11041);
and U16766 (N_16766,N_14103,N_12471);
and U16767 (N_16767,N_10103,N_12875);
and U16768 (N_16768,N_10186,N_13016);
nand U16769 (N_16769,N_10316,N_13243);
or U16770 (N_16770,N_11551,N_12265);
nand U16771 (N_16771,N_12357,N_11973);
or U16772 (N_16772,N_11887,N_12687);
or U16773 (N_16773,N_11407,N_12866);
xnor U16774 (N_16774,N_11746,N_12010);
xor U16775 (N_16775,N_11698,N_12273);
nand U16776 (N_16776,N_10059,N_11445);
and U16777 (N_16777,N_12315,N_14913);
nor U16778 (N_16778,N_10795,N_12284);
nand U16779 (N_16779,N_13535,N_12805);
and U16780 (N_16780,N_11497,N_12745);
nor U16781 (N_16781,N_13619,N_10237);
nand U16782 (N_16782,N_13727,N_14971);
or U16783 (N_16783,N_10731,N_11490);
and U16784 (N_16784,N_13678,N_11200);
nand U16785 (N_16785,N_13157,N_11479);
xor U16786 (N_16786,N_14533,N_12331);
nor U16787 (N_16787,N_11280,N_14510);
or U16788 (N_16788,N_10867,N_12840);
nand U16789 (N_16789,N_11858,N_10302);
or U16790 (N_16790,N_12074,N_10951);
and U16791 (N_16791,N_13485,N_12402);
nand U16792 (N_16792,N_12263,N_12907);
xnor U16793 (N_16793,N_13484,N_11638);
xor U16794 (N_16794,N_14579,N_11633);
xnor U16795 (N_16795,N_10829,N_12277);
nor U16796 (N_16796,N_13062,N_11461);
or U16797 (N_16797,N_13752,N_10055);
and U16798 (N_16798,N_13763,N_13964);
or U16799 (N_16799,N_10154,N_13406);
xnor U16800 (N_16800,N_12021,N_13894);
nor U16801 (N_16801,N_12342,N_10852);
or U16802 (N_16802,N_14031,N_11534);
and U16803 (N_16803,N_13770,N_14426);
and U16804 (N_16804,N_12425,N_13787);
or U16805 (N_16805,N_10041,N_11382);
nor U16806 (N_16806,N_14154,N_12170);
xnor U16807 (N_16807,N_11550,N_11689);
nand U16808 (N_16808,N_13213,N_12750);
nand U16809 (N_16809,N_11223,N_10570);
xnor U16810 (N_16810,N_14745,N_11444);
or U16811 (N_16811,N_13555,N_14899);
and U16812 (N_16812,N_14508,N_10110);
nand U16813 (N_16813,N_10989,N_14272);
and U16814 (N_16814,N_11726,N_11583);
and U16815 (N_16815,N_12686,N_10473);
nand U16816 (N_16816,N_10423,N_12814);
nor U16817 (N_16817,N_13926,N_10578);
and U16818 (N_16818,N_12671,N_12131);
xor U16819 (N_16819,N_12240,N_10934);
nand U16820 (N_16820,N_11205,N_13122);
xor U16821 (N_16821,N_10295,N_14093);
xnor U16822 (N_16822,N_11954,N_11069);
and U16823 (N_16823,N_14549,N_12288);
nor U16824 (N_16824,N_13066,N_11053);
and U16825 (N_16825,N_11373,N_14877);
and U16826 (N_16826,N_13353,N_10668);
nand U16827 (N_16827,N_10160,N_14067);
nor U16828 (N_16828,N_13131,N_13392);
and U16829 (N_16829,N_14146,N_12555);
or U16830 (N_16830,N_11230,N_10797);
xor U16831 (N_16831,N_13128,N_13266);
or U16832 (N_16832,N_12347,N_12803);
or U16833 (N_16833,N_11355,N_12790);
nand U16834 (N_16834,N_12155,N_14475);
xnor U16835 (N_16835,N_14225,N_10117);
or U16836 (N_16836,N_11625,N_11644);
or U16837 (N_16837,N_11560,N_10607);
and U16838 (N_16838,N_11370,N_14974);
and U16839 (N_16839,N_14073,N_13661);
or U16840 (N_16840,N_12121,N_11712);
nand U16841 (N_16841,N_12409,N_11162);
nand U16842 (N_16842,N_13939,N_10618);
nor U16843 (N_16843,N_10767,N_11604);
nand U16844 (N_16844,N_11727,N_13492);
and U16845 (N_16845,N_14528,N_11394);
nor U16846 (N_16846,N_11056,N_11021);
xnor U16847 (N_16847,N_13800,N_11970);
nor U16848 (N_16848,N_13272,N_12845);
or U16849 (N_16849,N_12811,N_12892);
nand U16850 (N_16850,N_10123,N_10850);
nand U16851 (N_16851,N_10531,N_10985);
nor U16852 (N_16852,N_10274,N_13168);
and U16853 (N_16853,N_14450,N_14969);
nand U16854 (N_16854,N_10499,N_13001);
nand U16855 (N_16855,N_10727,N_11995);
xor U16856 (N_16856,N_12132,N_10129);
and U16857 (N_16857,N_12793,N_14956);
xor U16858 (N_16858,N_12695,N_12392);
nor U16859 (N_16859,N_11246,N_11001);
or U16860 (N_16860,N_13832,N_10905);
nor U16861 (N_16861,N_10669,N_10714);
nor U16862 (N_16862,N_12719,N_10704);
and U16863 (N_16863,N_13847,N_12362);
nor U16864 (N_16864,N_12945,N_13669);
nand U16865 (N_16865,N_12587,N_14122);
or U16866 (N_16866,N_14988,N_13699);
or U16867 (N_16867,N_10313,N_14062);
and U16868 (N_16868,N_11531,N_11361);
nand U16869 (N_16869,N_13928,N_10165);
xor U16870 (N_16870,N_11165,N_14940);
xor U16871 (N_16871,N_14819,N_11554);
xor U16872 (N_16872,N_12376,N_13310);
nand U16873 (N_16873,N_10625,N_10817);
xor U16874 (N_16874,N_12677,N_12368);
and U16875 (N_16875,N_10769,N_12556);
and U16876 (N_16876,N_14716,N_10293);
or U16877 (N_16877,N_11096,N_11806);
nand U16878 (N_16878,N_10768,N_11458);
xnor U16879 (N_16879,N_14852,N_14735);
and U16880 (N_16880,N_10836,N_14643);
or U16881 (N_16881,N_10203,N_12559);
xor U16882 (N_16882,N_14482,N_12488);
xnor U16883 (N_16883,N_11294,N_14864);
and U16884 (N_16884,N_11250,N_11431);
xor U16885 (N_16885,N_13586,N_12884);
nor U16886 (N_16886,N_13491,N_13026);
nand U16887 (N_16887,N_10321,N_10579);
or U16888 (N_16888,N_14222,N_11829);
nor U16889 (N_16889,N_12771,N_11114);
or U16890 (N_16890,N_14592,N_13879);
nor U16891 (N_16891,N_11157,N_13359);
or U16892 (N_16892,N_13501,N_12220);
nand U16893 (N_16893,N_11570,N_13866);
xor U16894 (N_16894,N_10025,N_12223);
or U16895 (N_16895,N_14368,N_12136);
nand U16896 (N_16896,N_13482,N_12430);
nand U16897 (N_16897,N_10626,N_14344);
and U16898 (N_16898,N_10862,N_14264);
nand U16899 (N_16899,N_14613,N_11404);
nand U16900 (N_16900,N_11953,N_10557);
nor U16901 (N_16901,N_14531,N_14923);
nand U16902 (N_16902,N_14263,N_12902);
or U16903 (N_16903,N_13385,N_11368);
and U16904 (N_16904,N_11850,N_12008);
or U16905 (N_16905,N_11240,N_13767);
and U16906 (N_16906,N_12914,N_14089);
or U16907 (N_16907,N_13703,N_12038);
nand U16908 (N_16908,N_11541,N_13444);
nand U16909 (N_16909,N_12178,N_12482);
xnor U16910 (N_16910,N_10792,N_12620);
and U16911 (N_16911,N_13370,N_12968);
and U16912 (N_16912,N_10104,N_14112);
or U16913 (N_16913,N_11251,N_12084);
and U16914 (N_16914,N_11138,N_13908);
and U16915 (N_16915,N_11778,N_13852);
nand U16916 (N_16916,N_11102,N_12661);
xnor U16917 (N_16917,N_12540,N_12919);
nand U16918 (N_16918,N_12237,N_12318);
or U16919 (N_16919,N_14071,N_14442);
xor U16920 (N_16920,N_14431,N_10336);
or U16921 (N_16921,N_13652,N_14849);
and U16922 (N_16922,N_10130,N_10651);
nand U16923 (N_16923,N_11113,N_10533);
or U16924 (N_16924,N_10504,N_13312);
and U16925 (N_16925,N_13090,N_10116);
nand U16926 (N_16926,N_11634,N_11749);
nor U16927 (N_16927,N_12831,N_14995);
nand U16928 (N_16928,N_11797,N_13319);
xnor U16929 (N_16929,N_11674,N_10827);
nand U16930 (N_16930,N_14857,N_13287);
nand U16931 (N_16931,N_13000,N_13439);
and U16932 (N_16932,N_12312,N_12093);
nor U16933 (N_16933,N_10614,N_12251);
or U16934 (N_16934,N_11880,N_13065);
xnor U16935 (N_16935,N_13525,N_13053);
nand U16936 (N_16936,N_11300,N_11194);
nand U16937 (N_16937,N_14455,N_14432);
or U16938 (N_16938,N_14296,N_14025);
xnor U16939 (N_16939,N_13253,N_13506);
and U16940 (N_16940,N_12374,N_10595);
nand U16941 (N_16941,N_13498,N_10360);
nor U16942 (N_16942,N_10952,N_12204);
xnor U16943 (N_16943,N_13307,N_14775);
nor U16944 (N_16944,N_13938,N_14675);
nor U16945 (N_16945,N_12561,N_10505);
xor U16946 (N_16946,N_12807,N_14714);
and U16947 (N_16947,N_12466,N_12992);
nor U16948 (N_16948,N_14706,N_10559);
nor U16949 (N_16949,N_13435,N_13773);
xnor U16950 (N_16950,N_10931,N_11054);
and U16951 (N_16951,N_11694,N_12821);
and U16952 (N_16952,N_13811,N_12603);
or U16953 (N_16953,N_10495,N_13072);
nand U16954 (N_16954,N_11955,N_11139);
and U16955 (N_16955,N_12538,N_13978);
nor U16956 (N_16956,N_10959,N_14132);
xor U16957 (N_16957,N_10674,N_14004);
nor U16958 (N_16958,N_13344,N_14252);
and U16959 (N_16959,N_13700,N_14143);
xor U16960 (N_16960,N_13950,N_14174);
nand U16961 (N_16961,N_13250,N_14075);
and U16962 (N_16962,N_10326,N_14367);
and U16963 (N_16963,N_13942,N_10823);
nor U16964 (N_16964,N_13598,N_14425);
xnor U16965 (N_16965,N_14162,N_13456);
or U16966 (N_16966,N_13916,N_10000);
xor U16967 (N_16967,N_13630,N_11566);
nand U16968 (N_16968,N_13890,N_14791);
and U16969 (N_16969,N_12549,N_14539);
and U16970 (N_16970,N_12305,N_10924);
xnor U16971 (N_16971,N_11243,N_12812);
nand U16972 (N_16972,N_12379,N_12761);
nand U16973 (N_16973,N_14283,N_12610);
nor U16974 (N_16974,N_11077,N_14853);
and U16975 (N_16975,N_12388,N_13378);
xnor U16976 (N_16976,N_14108,N_12115);
or U16977 (N_16977,N_14287,N_10662);
and U16978 (N_16978,N_12751,N_10872);
nand U16979 (N_16979,N_13183,N_13145);
or U16980 (N_16980,N_10923,N_12922);
and U16981 (N_16981,N_11833,N_13473);
or U16982 (N_16982,N_13995,N_13190);
nand U16983 (N_16983,N_13755,N_10417);
nor U16984 (N_16984,N_10013,N_10314);
xor U16985 (N_16985,N_11679,N_10720);
nor U16986 (N_16986,N_12234,N_11946);
nor U16987 (N_16987,N_14023,N_10543);
xnor U16988 (N_16988,N_11820,N_12948);
and U16989 (N_16989,N_14843,N_12104);
nor U16990 (N_16990,N_12809,N_13288);
and U16991 (N_16991,N_11117,N_12028);
xnor U16992 (N_16992,N_10994,N_13925);
nor U16993 (N_16993,N_10535,N_10751);
or U16994 (N_16994,N_11721,N_14954);
and U16995 (N_16995,N_11197,N_11318);
xnor U16996 (N_16996,N_12190,N_13143);
or U16997 (N_16997,N_14085,N_14199);
and U16998 (N_16998,N_14206,N_11564);
and U16999 (N_16999,N_12317,N_14152);
xor U17000 (N_17000,N_13489,N_14445);
nor U17001 (N_17001,N_14562,N_10173);
nor U17002 (N_17002,N_12270,N_12232);
xnor U17003 (N_17003,N_14751,N_10011);
xor U17004 (N_17004,N_10412,N_12085);
and U17005 (N_17005,N_12298,N_10197);
and U17006 (N_17006,N_14402,N_14453);
nand U17007 (N_17007,N_14223,N_13951);
xnor U17008 (N_17008,N_11839,N_14339);
xnor U17009 (N_17009,N_14377,N_14590);
or U17010 (N_17010,N_13390,N_10226);
and U17011 (N_17011,N_13300,N_12079);
nand U17012 (N_17012,N_11126,N_10388);
xnor U17013 (N_17013,N_10580,N_14907);
nand U17014 (N_17014,N_12560,N_10631);
xnor U17015 (N_17015,N_11964,N_12475);
nor U17016 (N_17016,N_14364,N_14325);
or U17017 (N_17017,N_12146,N_10629);
nor U17018 (N_17018,N_13427,N_14155);
xor U17019 (N_17019,N_11920,N_14213);
nand U17020 (N_17020,N_13524,N_13604);
or U17021 (N_17021,N_10300,N_11655);
xnor U17022 (N_17022,N_12212,N_10974);
xnor U17023 (N_17023,N_11618,N_10017);
nand U17024 (N_17024,N_13092,N_14414);
nor U17025 (N_17025,N_11478,N_14677);
or U17026 (N_17026,N_12163,N_14461);
nor U17027 (N_17027,N_13032,N_11270);
and U17028 (N_17028,N_13897,N_12384);
xor U17029 (N_17029,N_14622,N_13690);
nor U17030 (N_17030,N_10211,N_10118);
or U17031 (N_17031,N_11752,N_10020);
and U17032 (N_17032,N_11735,N_14102);
or U17033 (N_17033,N_13308,N_14489);
xnor U17034 (N_17034,N_10556,N_12500);
nand U17035 (N_17035,N_12956,N_10700);
xor U17036 (N_17036,N_14024,N_10919);
nor U17037 (N_17037,N_11647,N_10808);
nor U17038 (N_17038,N_10697,N_11452);
or U17039 (N_17039,N_13421,N_12418);
or U17040 (N_17040,N_11565,N_11719);
nor U17041 (N_17041,N_10870,N_10045);
nor U17042 (N_17042,N_13160,N_13275);
nand U17043 (N_17043,N_11470,N_10861);
or U17044 (N_17044,N_10602,N_10387);
nor U17045 (N_17045,N_14163,N_12139);
and U17046 (N_17046,N_12058,N_12011);
and U17047 (N_17047,N_11670,N_13039);
nand U17048 (N_17048,N_12514,N_11519);
nor U17049 (N_17049,N_10125,N_12363);
xor U17050 (N_17050,N_13771,N_12949);
nand U17051 (N_17051,N_11594,N_13687);
nor U17052 (N_17052,N_10132,N_13446);
xnor U17053 (N_17053,N_13135,N_11529);
xor U17054 (N_17054,N_14984,N_14776);
or U17055 (N_17055,N_12970,N_14369);
xor U17056 (N_17056,N_13480,N_14540);
or U17057 (N_17057,N_12938,N_12941);
and U17058 (N_17058,N_14973,N_10755);
xnor U17059 (N_17059,N_10021,N_12552);
or U17060 (N_17060,N_10980,N_13280);
or U17061 (N_17061,N_14117,N_14478);
and U17062 (N_17062,N_13839,N_13673);
nand U17063 (N_17063,N_12295,N_10876);
or U17064 (N_17064,N_12492,N_14603);
xnor U17065 (N_17065,N_10415,N_11029);
or U17066 (N_17066,N_10813,N_12599);
xnor U17067 (N_17067,N_11426,N_13623);
or U17068 (N_17068,N_13726,N_12031);
or U17069 (N_17069,N_11736,N_13093);
nor U17070 (N_17070,N_11344,N_13622);
xnor U17071 (N_17071,N_13315,N_11768);
xnor U17072 (N_17072,N_10487,N_10457);
and U17073 (N_17073,N_14181,N_13836);
nor U17074 (N_17074,N_12235,N_13556);
or U17075 (N_17075,N_10666,N_10152);
and U17076 (N_17076,N_12932,N_11865);
nand U17077 (N_17077,N_14785,N_10181);
nand U17078 (N_17078,N_10459,N_10220);
xor U17079 (N_17079,N_11989,N_10911);
or U17080 (N_17080,N_11070,N_13721);
nand U17081 (N_17081,N_10660,N_13889);
or U17082 (N_17082,N_14903,N_10875);
xnor U17083 (N_17083,N_10835,N_11346);
xnor U17084 (N_17084,N_13961,N_14669);
xnor U17085 (N_17085,N_10015,N_14850);
nor U17086 (N_17086,N_11399,N_14231);
nor U17087 (N_17087,N_12014,N_14778);
nand U17088 (N_17088,N_12174,N_12904);
nand U17089 (N_17089,N_11492,N_14905);
xnor U17090 (N_17090,N_13296,N_10456);
nor U17091 (N_17091,N_14008,N_10155);
nand U17092 (N_17092,N_14820,N_14465);
or U17093 (N_17093,N_10790,N_10848);
nor U17094 (N_17094,N_13450,N_11349);
or U17095 (N_17095,N_10746,N_13393);
xnor U17096 (N_17096,N_13782,N_13221);
xor U17097 (N_17097,N_12744,N_11591);
and U17098 (N_17098,N_14055,N_14334);
xnor U17099 (N_17099,N_14135,N_13037);
and U17100 (N_17100,N_12584,N_10975);
nor U17101 (N_17101,N_14945,N_10288);
nand U17102 (N_17102,N_11992,N_10370);
and U17103 (N_17103,N_14876,N_10558);
nor U17104 (N_17104,N_11874,N_12349);
xor U17105 (N_17105,N_14898,N_11568);
nor U17106 (N_17106,N_12656,N_11462);
and U17107 (N_17107,N_12395,N_13736);
xnor U17108 (N_17108,N_11449,N_14733);
and U17109 (N_17109,N_14308,N_10532);
or U17110 (N_17110,N_11518,N_14403);
nor U17111 (N_17111,N_10726,N_10732);
or U17112 (N_17112,N_12070,N_10448);
and U17113 (N_17113,N_10324,N_11443);
or U17114 (N_17114,N_10368,N_13789);
nand U17115 (N_17115,N_13211,N_13868);
nand U17116 (N_17116,N_13895,N_13404);
nor U17117 (N_17117,N_10396,N_13881);
and U17118 (N_17118,N_11227,N_10190);
or U17119 (N_17119,N_10420,N_11696);
nor U17120 (N_17120,N_12841,N_10189);
or U17121 (N_17121,N_10286,N_12219);
and U17122 (N_17122,N_13150,N_10373);
and U17123 (N_17123,N_14331,N_14787);
or U17124 (N_17124,N_10365,N_10001);
or U17125 (N_17125,N_10233,N_11680);
and U17126 (N_17126,N_10224,N_14156);
xnor U17127 (N_17127,N_10255,N_10856);
and U17128 (N_17128,N_12216,N_11073);
and U17129 (N_17129,N_14806,N_10112);
xor U17130 (N_17130,N_13977,N_12736);
xor U17131 (N_17131,N_14433,N_13286);
nand U17132 (N_17132,N_11884,N_12593);
and U17133 (N_17133,N_12990,N_13078);
and U17134 (N_17134,N_11868,N_10964);
and U17135 (N_17135,N_12806,N_12328);
nand U17136 (N_17136,N_11389,N_10885);
nor U17137 (N_17137,N_10142,N_11434);
xor U17138 (N_17138,N_11910,N_13634);
or U17139 (N_17139,N_13314,N_14556);
nand U17140 (N_17140,N_14311,N_13785);
nand U17141 (N_17141,N_10681,N_10740);
or U17142 (N_17142,N_14671,N_12509);
nand U17143 (N_17143,N_11057,N_14401);
or U17144 (N_17144,N_14594,N_14645);
and U17145 (N_17145,N_12663,N_11557);
or U17146 (N_17146,N_14167,N_14159);
nor U17147 (N_17147,N_12737,N_12738);
nand U17148 (N_17148,N_13015,N_12122);
and U17149 (N_17149,N_10377,N_14059);
nor U17150 (N_17150,N_11279,N_14682);
and U17151 (N_17151,N_13106,N_14190);
xnor U17152 (N_17152,N_12654,N_11900);
and U17153 (N_17153,N_11595,N_14542);
nand U17154 (N_17154,N_12660,N_13641);
or U17155 (N_17155,N_11921,N_10325);
and U17156 (N_17156,N_14333,N_11190);
and U17157 (N_17157,N_11799,N_14950);
and U17158 (N_17158,N_11466,N_12789);
xor U17159 (N_17159,N_12954,N_14524);
and U17160 (N_17160,N_14753,N_10749);
or U17161 (N_17161,N_12355,N_14568);
or U17162 (N_17162,N_11788,N_11851);
and U17163 (N_17163,N_12378,N_10315);
xor U17164 (N_17164,N_11856,N_10182);
and U17165 (N_17165,N_11015,N_13828);
nand U17166 (N_17166,N_10378,N_10894);
xor U17167 (N_17167,N_14937,N_14188);
nand U17168 (N_17168,N_11682,N_13483);
xor U17169 (N_17169,N_12157,N_10783);
xnor U17170 (N_17170,N_13486,N_13716);
nand U17171 (N_17171,N_13730,N_12700);
nand U17172 (N_17172,N_12578,N_10512);
xor U17173 (N_17173,N_14288,N_11317);
xnor U17174 (N_17174,N_14760,N_10192);
xnor U17175 (N_17175,N_14474,N_11879);
nand U17176 (N_17176,N_13569,N_14963);
xnor U17177 (N_17177,N_13656,N_12077);
nor U17178 (N_17178,N_14321,N_10283);
nand U17179 (N_17179,N_10141,N_12027);
xnor U17180 (N_17180,N_14479,N_11078);
nand U17181 (N_17181,N_12580,N_14813);
nand U17182 (N_17182,N_14346,N_14541);
or U17183 (N_17183,N_13334,N_12066);
nor U17184 (N_17184,N_11265,N_13625);
nand U17185 (N_17185,N_10047,N_11039);
or U17186 (N_17186,N_10471,N_11089);
or U17187 (N_17187,N_14293,N_11111);
nand U17188 (N_17188,N_10866,N_13101);
xnor U17189 (N_17189,N_13899,N_12973);
or U17190 (N_17190,N_14792,N_10338);
nand U17191 (N_17191,N_12023,N_14861);
or U17192 (N_17192,N_10090,N_14158);
nand U17193 (N_17193,N_14757,N_13094);
xnor U17194 (N_17194,N_14657,N_13869);
nor U17195 (N_17195,N_10486,N_14360);
and U17196 (N_17196,N_12134,N_12446);
or U17197 (N_17197,N_11433,N_13289);
nand U17198 (N_17198,N_11685,N_13017);
xnor U17199 (N_17199,N_13004,N_12452);
xnor U17200 (N_17200,N_13803,N_11273);
nor U17201 (N_17201,N_11590,N_10719);
nand U17202 (N_17202,N_14908,N_14608);
nand U17203 (N_17203,N_14989,N_10957);
nand U17204 (N_17204,N_11951,N_10868);
and U17205 (N_17205,N_11148,N_13326);
and U17206 (N_17206,N_11933,N_12100);
nand U17207 (N_17207,N_13841,N_11854);
xnor U17208 (N_17208,N_10992,N_14741);
or U17209 (N_17209,N_12959,N_10408);
and U17210 (N_17210,N_12410,N_11885);
xnor U17211 (N_17211,N_13783,N_14662);
nor U17212 (N_17212,N_12529,N_13411);
or U17213 (N_17213,N_13481,N_12946);
or U17214 (N_17214,N_13355,N_11446);
nand U17215 (N_17215,N_13772,N_10259);
xor U17216 (N_17216,N_12162,N_11572);
nor U17217 (N_17217,N_11883,N_11306);
nor U17218 (N_17218,N_11861,N_11395);
or U17219 (N_17219,N_12043,N_14873);
or U17220 (N_17220,N_12715,N_12173);
xnor U17221 (N_17221,N_14812,N_13842);
and U17222 (N_17222,N_11805,N_13171);
and U17223 (N_17223,N_14648,N_10903);
nor U17224 (N_17224,N_11671,N_10883);
nand U17225 (N_17225,N_13533,N_10855);
xor U17226 (N_17226,N_13613,N_10174);
xor U17227 (N_17227,N_14497,N_12558);
nand U17228 (N_17228,N_12408,N_10028);
nor U17229 (N_17229,N_12024,N_13021);
xnor U17230 (N_17230,N_14332,N_13049);
nor U17231 (N_17231,N_14926,N_13200);
nand U17232 (N_17232,N_13927,N_13920);
nand U17233 (N_17233,N_14559,N_10671);
nor U17234 (N_17234,N_11976,N_14627);
nand U17235 (N_17235,N_11714,N_12667);
xor U17236 (N_17236,N_12125,N_13568);
and U17237 (N_17237,N_10821,N_10820);
nand U17238 (N_17238,N_10042,N_11127);
nand U17239 (N_17239,N_10555,N_13468);
nor U17240 (N_17240,N_13549,N_11782);
nand U17241 (N_17241,N_10545,N_11172);
nand U17242 (N_17242,N_13155,N_13873);
and U17243 (N_17243,N_12107,N_12601);
nand U17244 (N_17244,N_12541,N_11819);
nor U17245 (N_17245,N_11562,N_12153);
and U17246 (N_17246,N_11116,N_13430);
or U17247 (N_17247,N_13120,N_11546);
xor U17248 (N_17248,N_11972,N_12982);
nor U17249 (N_17249,N_14405,N_10639);
or U17250 (N_17250,N_14770,N_14271);
or U17251 (N_17251,N_14340,N_14566);
nor U17252 (N_17252,N_10068,N_14081);
nor U17253 (N_17253,N_12762,N_13419);
xnor U17254 (N_17254,N_10776,N_13304);
nand U17255 (N_17255,N_14447,N_14582);
and U17256 (N_17256,N_12820,N_14829);
and U17257 (N_17257,N_14863,N_14693);
xnor U17258 (N_17258,N_13137,N_12524);
and U17259 (N_17259,N_10650,N_12102);
nand U17260 (N_17260,N_14554,N_12338);
and U17261 (N_17261,N_13507,N_11142);
and U17262 (N_17262,N_10772,N_13593);
nand U17263 (N_17263,N_10534,N_10577);
nor U17264 (N_17264,N_14435,N_10475);
xnor U17265 (N_17265,N_12815,N_14572);
xor U17266 (N_17266,N_13814,N_10592);
nand U17267 (N_17267,N_13055,N_10818);
and U17268 (N_17268,N_12447,N_10319);
and U17269 (N_17269,N_10936,N_11857);
and U17270 (N_17270,N_13940,N_13380);
nand U17271 (N_17271,N_14738,N_11182);
xor U17272 (N_17272,N_13394,N_11961);
xnor U17273 (N_17273,N_11335,N_14441);
nor U17274 (N_17274,N_10549,N_11906);
nor U17275 (N_17275,N_14892,N_14616);
xor U17276 (N_17276,N_12950,N_14400);
and U17277 (N_17277,N_10984,N_13228);
nand U17278 (N_17278,N_11281,N_14578);
nand U17279 (N_17279,N_14003,N_14771);
or U17280 (N_17280,N_13185,N_13002);
nor U17281 (N_17281,N_12766,N_11242);
nand U17282 (N_17282,N_14615,N_11893);
and U17283 (N_17283,N_10273,N_10294);
or U17284 (N_17284,N_10598,N_10426);
nand U17285 (N_17285,N_10105,N_10410);
nand U17286 (N_17286,N_11347,N_12635);
xnor U17287 (N_17287,N_14911,N_13693);
and U17288 (N_17288,N_13645,N_14383);
xnor U17289 (N_17289,N_14626,N_13668);
xor U17290 (N_17290,N_12877,N_14784);
xnor U17291 (N_17291,N_11209,N_11663);
or U17292 (N_17292,N_11525,N_13298);
nor U17293 (N_17293,N_13509,N_13223);
or U17294 (N_17294,N_12428,N_14909);
nand U17295 (N_17295,N_10311,N_13400);
xnor U17296 (N_17296,N_10506,N_10350);
xnor U17297 (N_17297,N_14803,N_11892);
nand U17298 (N_17298,N_14329,N_11045);
or U17299 (N_17299,N_12797,N_12213);
or U17300 (N_17300,N_10766,N_10454);
nor U17301 (N_17301,N_11428,N_14316);
nor U17302 (N_17302,N_13791,N_11334);
xnor U17303 (N_17303,N_12754,N_11662);
nand U17304 (N_17304,N_10386,N_13969);
xnor U17305 (N_17305,N_13846,N_11416);
nor U17306 (N_17306,N_12980,N_10496);
xor U17307 (N_17307,N_11902,N_12604);
nor U17308 (N_17308,N_13840,N_13596);
xnor U17309 (N_17309,N_10498,N_11767);
and U17310 (N_17310,N_10659,N_13971);
nand U17311 (N_17311,N_13499,N_12953);
nand U17312 (N_17312,N_10241,N_13068);
nand U17313 (N_17313,N_13351,N_12683);
or U17314 (N_17314,N_13109,N_12465);
xor U17315 (N_17315,N_11048,N_12462);
xor U17316 (N_17316,N_11145,N_10644);
and U17317 (N_17317,N_11176,N_13227);
and U17318 (N_17318,N_14232,N_14659);
nor U17319 (N_17319,N_10968,N_13434);
nor U17320 (N_17320,N_13830,N_12585);
xnor U17321 (N_17321,N_10904,N_11110);
and U17322 (N_17322,N_14570,N_10702);
or U17323 (N_17323,N_13719,N_14010);
or U17324 (N_17324,N_12025,N_14835);
xnor U17325 (N_17325,N_12231,N_14752);
and U17326 (N_17326,N_13295,N_14838);
and U17327 (N_17327,N_13214,N_12854);
or U17328 (N_17328,N_11301,N_12291);
xor U17329 (N_17329,N_10892,N_12897);
and U17330 (N_17330,N_11123,N_13802);
and U17331 (N_17331,N_13594,N_13688);
and U17332 (N_17332,N_12847,N_11169);
nand U17333 (N_17333,N_10623,N_12876);
xor U17334 (N_17334,N_14164,N_13219);
nand U17335 (N_17335,N_11020,N_12498);
nor U17336 (N_17336,N_13918,N_10113);
xor U17337 (N_17337,N_10256,N_12094);
nand U17338 (N_17338,N_13217,N_14203);
nand U17339 (N_17339,N_13572,N_13029);
and U17340 (N_17340,N_12796,N_12666);
xor U17341 (N_17341,N_14304,N_12842);
nand U17342 (N_17342,N_14498,N_14606);
xnor U17343 (N_17343,N_14532,N_10947);
nand U17344 (N_17344,N_10009,N_13086);
nor U17345 (N_17345,N_12828,N_14384);
nor U17346 (N_17346,N_14200,N_12508);
nor U17347 (N_17347,N_14605,N_14246);
nand U17348 (N_17348,N_10354,N_13191);
and U17349 (N_17349,N_11766,N_11637);
nor U17350 (N_17350,N_12853,N_11994);
or U17351 (N_17351,N_13277,N_10800);
nand U17352 (N_17352,N_13717,N_13974);
and U17353 (N_17353,N_12557,N_13201);
nor U17354 (N_17354,N_13986,N_10785);
or U17355 (N_17355,N_11032,N_11898);
nand U17356 (N_17356,N_14219,N_14258);
xor U17357 (N_17357,N_14793,N_12995);
xnor U17358 (N_17358,N_10791,N_11977);
or U17359 (N_17359,N_14301,N_10886);
nand U17360 (N_17360,N_13166,N_13826);
or U17361 (N_17361,N_10581,N_14668);
and U17362 (N_17362,N_13735,N_13232);
or U17363 (N_17363,N_12864,N_13917);
xor U17364 (N_17364,N_10056,N_12690);
xnor U17365 (N_17365,N_14282,N_12087);
nand U17366 (N_17366,N_13350,N_13616);
xnor U17367 (N_17367,N_11040,N_14513);
nor U17368 (N_17368,N_11930,N_13416);
nor U17369 (N_17369,N_11400,N_12130);
nand U17370 (N_17370,N_14642,N_13276);
and U17371 (N_17371,N_11507,N_14001);
nand U17372 (N_17372,N_10743,N_10008);
or U17373 (N_17373,N_13133,N_10585);
or U17374 (N_17374,N_13178,N_12564);
nor U17375 (N_17375,N_12398,N_11836);
and U17376 (N_17376,N_12735,N_10698);
xnor U17377 (N_17377,N_10858,N_11425);
and U17378 (N_17378,N_13442,N_11199);
nand U17379 (N_17379,N_14862,N_13990);
xnor U17380 (N_17380,N_10641,N_13579);
or U17381 (N_17381,N_10891,N_11905);
nor U17382 (N_17382,N_14228,N_11770);
nor U17383 (N_17383,N_12356,N_13702);
or U17384 (N_17384,N_12983,N_12867);
nand U17385 (N_17385,N_13564,N_14418);
nand U17386 (N_17386,N_11632,N_14420);
or U17387 (N_17387,N_11706,N_11513);
nor U17388 (N_17388,N_10407,N_10196);
nor U17389 (N_17389,N_11135,N_12930);
and U17390 (N_17390,N_14487,N_12081);
or U17391 (N_17391,N_13821,N_12640);
nor U17392 (N_17392,N_13472,N_11624);
nor U17393 (N_17393,N_13947,N_13737);
nor U17394 (N_17394,N_13433,N_11464);
or U17395 (N_17395,N_10807,N_14172);
nand U17396 (N_17396,N_11340,N_12249);
nand U17397 (N_17397,N_12707,N_14902);
and U17398 (N_17398,N_14558,N_12242);
and U17399 (N_17399,N_11255,N_11882);
xor U17400 (N_17400,N_10077,N_10081);
nand U17401 (N_17401,N_12846,N_13792);
xnor U17402 (N_17402,N_13626,N_12176);
xor U17403 (N_17403,N_11886,N_13913);
and U17404 (N_17404,N_11064,N_10416);
xor U17405 (N_17405,N_11758,N_14481);
xnor U17406 (N_17406,N_12997,N_14049);
nor U17407 (N_17407,N_10279,N_13943);
nor U17408 (N_17408,N_10046,N_10043);
nor U17409 (N_17409,N_13405,N_14681);
xor U17410 (N_17410,N_12569,N_12415);
nor U17411 (N_17411,N_12400,N_12202);
nand U17412 (N_17412,N_10573,N_13358);
nand U17413 (N_17413,N_12048,N_12090);
nor U17414 (N_17414,N_10491,N_12169);
or U17415 (N_17415,N_11776,N_12019);
and U17416 (N_17416,N_10075,N_10859);
and U17417 (N_17417,N_11686,N_10993);
nand U17418 (N_17418,N_12551,N_12172);
or U17419 (N_17419,N_13597,N_10392);
xor U17420 (N_17420,N_10371,N_14239);
or U17421 (N_17421,N_11540,N_14968);
and U17422 (N_17422,N_14454,N_10834);
nand U17423 (N_17423,N_12641,N_11103);
nand U17424 (N_17424,N_12727,N_11817);
nand U17425 (N_17425,N_12412,N_12386);
xor U17426 (N_17426,N_14823,N_14300);
xor U17427 (N_17427,N_13747,N_14573);
nor U17428 (N_17428,N_11574,N_14412);
or U17429 (N_17429,N_10970,N_14865);
nor U17430 (N_17430,N_10509,N_14694);
xnor U17431 (N_17431,N_12929,N_11939);
xor U17432 (N_17432,N_11118,N_11510);
and U17433 (N_17433,N_10085,N_11495);
or U17434 (N_17434,N_11234,N_12862);
nor U17435 (N_17435,N_12764,N_14444);
nand U17436 (N_17436,N_13495,N_10403);
nand U17437 (N_17437,N_11684,N_14830);
or U17438 (N_17438,N_10596,N_14726);
nand U17439 (N_17439,N_11785,N_10735);
or U17440 (N_17440,N_14061,N_13945);
nor U17441 (N_17441,N_13132,N_13318);
or U17442 (N_17442,N_11708,N_10507);
nor U17443 (N_17443,N_12380,N_12721);
xor U17444 (N_17444,N_14389,N_13254);
and U17445 (N_17445,N_10195,N_11448);
and U17446 (N_17446,N_13006,N_12804);
or U17447 (N_17447,N_14996,N_12334);
xor U17448 (N_17448,N_10594,N_13815);
xnor U17449 (N_17449,N_13284,N_10853);
xor U17450 (N_17450,N_12679,N_10679);
nor U17451 (N_17451,N_14964,N_11432);
nor U17452 (N_17452,N_10153,N_14128);
nand U17453 (N_17453,N_14548,N_11580);
and U17454 (N_17454,N_11235,N_10770);
and U17455 (N_17455,N_14069,N_14125);
nand U17456 (N_17456,N_10348,N_14224);
nand U17457 (N_17457,N_10942,N_11401);
xor U17458 (N_17458,N_14755,N_14800);
and U17459 (N_17459,N_13809,N_13469);
nand U17460 (N_17460,N_14218,N_13786);
or U17461 (N_17461,N_12373,N_14692);
xor U17462 (N_17462,N_13381,N_10394);
xor U17463 (N_17463,N_10065,N_11783);
xnor U17464 (N_17464,N_13587,N_12257);
and U17465 (N_17465,N_10243,N_12625);
xnor U17466 (N_17466,N_13724,N_12858);
nand U17467 (N_17467,N_13268,N_13848);
nor U17468 (N_17468,N_11095,N_12199);
xor U17469 (N_17469,N_10303,N_14587);
or U17470 (N_17470,N_12013,N_10709);
and U17471 (N_17471,N_13819,N_10739);
nand U17472 (N_17472,N_11514,N_11071);
and U17473 (N_17473,N_13537,N_12621);
or U17474 (N_17474,N_14491,N_12888);
nor U17475 (N_17475,N_14327,N_14466);
xor U17476 (N_17476,N_10114,N_10638);
xnor U17477 (N_17477,N_12473,N_12674);
and U17478 (N_17478,N_13900,N_14138);
nand U17479 (N_17479,N_11620,N_13386);
xor U17480 (N_17480,N_14618,N_13051);
nor U17481 (N_17481,N_10329,N_14468);
or U17482 (N_17482,N_13322,N_10366);
or U17483 (N_17483,N_11530,N_12606);
nor U17484 (N_17484,N_14868,N_10469);
and U17485 (N_17485,N_14872,N_12720);
and U17486 (N_17486,N_12439,N_11943);
nor U17487 (N_17487,N_11704,N_11862);
xor U17488 (N_17488,N_12303,N_14881);
and U17489 (N_17489,N_12499,N_10101);
nand U17490 (N_17490,N_11627,N_11074);
nand U17491 (N_17491,N_12899,N_14517);
or U17492 (N_17492,N_14423,N_11571);
xnor U17493 (N_17493,N_11798,N_14440);
xor U17494 (N_17494,N_14982,N_13328);
or U17495 (N_17495,N_12655,N_13075);
nand U17496 (N_17496,N_10560,N_10002);
nor U17497 (N_17497,N_10517,N_12501);
xnor U17498 (N_17498,N_14828,N_11761);
xnor U17499 (N_17499,N_12209,N_10352);
nor U17500 (N_17500,N_14608,N_12938);
nor U17501 (N_17501,N_10154,N_14439);
xnor U17502 (N_17502,N_13419,N_14966);
or U17503 (N_17503,N_13535,N_10070);
nor U17504 (N_17504,N_12339,N_11370);
or U17505 (N_17505,N_14340,N_10050);
nand U17506 (N_17506,N_11079,N_10882);
and U17507 (N_17507,N_11151,N_11750);
or U17508 (N_17508,N_12004,N_13961);
xor U17509 (N_17509,N_14093,N_14880);
and U17510 (N_17510,N_10787,N_13543);
or U17511 (N_17511,N_11561,N_12841);
and U17512 (N_17512,N_11137,N_11447);
nand U17513 (N_17513,N_10637,N_14509);
nand U17514 (N_17514,N_10118,N_11147);
nor U17515 (N_17515,N_10187,N_12995);
and U17516 (N_17516,N_13646,N_13626);
and U17517 (N_17517,N_10997,N_13840);
and U17518 (N_17518,N_11914,N_11249);
or U17519 (N_17519,N_13617,N_12966);
nor U17520 (N_17520,N_13020,N_12545);
or U17521 (N_17521,N_13653,N_11813);
nand U17522 (N_17522,N_13599,N_12884);
xor U17523 (N_17523,N_12592,N_14980);
or U17524 (N_17524,N_13595,N_14730);
or U17525 (N_17525,N_13770,N_12429);
and U17526 (N_17526,N_11700,N_14569);
xor U17527 (N_17527,N_14507,N_12390);
or U17528 (N_17528,N_14989,N_11484);
xnor U17529 (N_17529,N_11553,N_10683);
xnor U17530 (N_17530,N_14178,N_13447);
and U17531 (N_17531,N_14326,N_10346);
and U17532 (N_17532,N_12432,N_10642);
or U17533 (N_17533,N_11154,N_10778);
or U17534 (N_17534,N_13972,N_14021);
nand U17535 (N_17535,N_13428,N_11211);
nand U17536 (N_17536,N_13968,N_12334);
nand U17537 (N_17537,N_11696,N_12720);
nor U17538 (N_17538,N_10699,N_12229);
and U17539 (N_17539,N_11628,N_10707);
and U17540 (N_17540,N_13068,N_12818);
or U17541 (N_17541,N_12689,N_11290);
nand U17542 (N_17542,N_10171,N_14634);
nand U17543 (N_17543,N_14422,N_12960);
and U17544 (N_17544,N_11185,N_13513);
and U17545 (N_17545,N_12583,N_10306);
or U17546 (N_17546,N_11681,N_12477);
xor U17547 (N_17547,N_12208,N_11260);
and U17548 (N_17548,N_14854,N_12023);
nor U17549 (N_17549,N_12296,N_11310);
and U17550 (N_17550,N_13050,N_10154);
nor U17551 (N_17551,N_11401,N_10530);
or U17552 (N_17552,N_10842,N_12429);
or U17553 (N_17553,N_10777,N_10293);
or U17554 (N_17554,N_10701,N_12310);
nand U17555 (N_17555,N_10221,N_10310);
or U17556 (N_17556,N_13065,N_13180);
or U17557 (N_17557,N_13220,N_10534);
nor U17558 (N_17558,N_10225,N_10044);
nor U17559 (N_17559,N_13182,N_11297);
and U17560 (N_17560,N_14044,N_14635);
xnor U17561 (N_17561,N_10744,N_14007);
nand U17562 (N_17562,N_13543,N_13032);
or U17563 (N_17563,N_11537,N_13535);
xor U17564 (N_17564,N_10738,N_10540);
xnor U17565 (N_17565,N_12071,N_10462);
xnor U17566 (N_17566,N_14679,N_12168);
nor U17567 (N_17567,N_13024,N_13995);
nand U17568 (N_17568,N_12265,N_13135);
nor U17569 (N_17569,N_11633,N_14093);
or U17570 (N_17570,N_12530,N_13770);
or U17571 (N_17571,N_11866,N_12903);
xnor U17572 (N_17572,N_13023,N_13211);
and U17573 (N_17573,N_10152,N_12559);
nand U17574 (N_17574,N_14784,N_10382);
and U17575 (N_17575,N_11137,N_10389);
or U17576 (N_17576,N_12666,N_12527);
nor U17577 (N_17577,N_11481,N_10125);
nand U17578 (N_17578,N_13118,N_10267);
and U17579 (N_17579,N_14178,N_13719);
xor U17580 (N_17580,N_14058,N_14594);
or U17581 (N_17581,N_12537,N_11574);
and U17582 (N_17582,N_10852,N_12246);
or U17583 (N_17583,N_14361,N_11135);
xor U17584 (N_17584,N_11972,N_11998);
or U17585 (N_17585,N_12770,N_12940);
or U17586 (N_17586,N_11270,N_12698);
xnor U17587 (N_17587,N_13362,N_12670);
or U17588 (N_17588,N_11313,N_14800);
nor U17589 (N_17589,N_13185,N_12998);
nor U17590 (N_17590,N_11554,N_10000);
nand U17591 (N_17591,N_11522,N_14707);
and U17592 (N_17592,N_12587,N_13957);
nand U17593 (N_17593,N_12139,N_14359);
nand U17594 (N_17594,N_11996,N_13690);
nand U17595 (N_17595,N_12918,N_11315);
nand U17596 (N_17596,N_13542,N_10819);
and U17597 (N_17597,N_12848,N_13691);
or U17598 (N_17598,N_12950,N_13709);
xor U17599 (N_17599,N_14367,N_12718);
or U17600 (N_17600,N_14847,N_14559);
xor U17601 (N_17601,N_14349,N_11861);
or U17602 (N_17602,N_10364,N_11889);
or U17603 (N_17603,N_14392,N_11513);
or U17604 (N_17604,N_12577,N_11517);
and U17605 (N_17605,N_10636,N_10043);
or U17606 (N_17606,N_13409,N_13724);
and U17607 (N_17607,N_13592,N_10014);
nand U17608 (N_17608,N_10092,N_10065);
xor U17609 (N_17609,N_12260,N_14288);
xor U17610 (N_17610,N_13063,N_14288);
nor U17611 (N_17611,N_12361,N_13407);
xnor U17612 (N_17612,N_11977,N_10648);
or U17613 (N_17613,N_13214,N_14961);
or U17614 (N_17614,N_13173,N_11500);
or U17615 (N_17615,N_12012,N_14487);
or U17616 (N_17616,N_13346,N_10872);
or U17617 (N_17617,N_14201,N_14714);
and U17618 (N_17618,N_14921,N_13753);
nand U17619 (N_17619,N_11070,N_12054);
xor U17620 (N_17620,N_10589,N_14326);
nand U17621 (N_17621,N_13622,N_13775);
and U17622 (N_17622,N_14874,N_10109);
nand U17623 (N_17623,N_12309,N_12580);
or U17624 (N_17624,N_11763,N_14414);
and U17625 (N_17625,N_14751,N_10631);
or U17626 (N_17626,N_12486,N_10691);
or U17627 (N_17627,N_12682,N_14394);
and U17628 (N_17628,N_11685,N_12039);
or U17629 (N_17629,N_11635,N_12999);
or U17630 (N_17630,N_13154,N_10346);
xor U17631 (N_17631,N_13540,N_12640);
nand U17632 (N_17632,N_14414,N_13810);
nor U17633 (N_17633,N_14067,N_13305);
nor U17634 (N_17634,N_12960,N_12784);
nand U17635 (N_17635,N_11666,N_12675);
xor U17636 (N_17636,N_14771,N_13842);
nand U17637 (N_17637,N_13469,N_14889);
and U17638 (N_17638,N_10133,N_10136);
nand U17639 (N_17639,N_11041,N_14956);
nor U17640 (N_17640,N_13741,N_10414);
nand U17641 (N_17641,N_14389,N_10795);
nand U17642 (N_17642,N_12440,N_10856);
and U17643 (N_17643,N_14017,N_11584);
xnor U17644 (N_17644,N_12247,N_13655);
nor U17645 (N_17645,N_11321,N_12292);
and U17646 (N_17646,N_11101,N_11350);
nor U17647 (N_17647,N_13711,N_10998);
xor U17648 (N_17648,N_12451,N_12984);
xor U17649 (N_17649,N_11926,N_11442);
nand U17650 (N_17650,N_11964,N_10620);
nand U17651 (N_17651,N_13018,N_14928);
nand U17652 (N_17652,N_10394,N_14857);
nand U17653 (N_17653,N_12913,N_10190);
and U17654 (N_17654,N_10445,N_14883);
or U17655 (N_17655,N_11411,N_13095);
nand U17656 (N_17656,N_14803,N_10341);
or U17657 (N_17657,N_12905,N_10406);
nand U17658 (N_17658,N_14504,N_13069);
nand U17659 (N_17659,N_12602,N_10459);
or U17660 (N_17660,N_13649,N_13367);
xor U17661 (N_17661,N_14957,N_11497);
or U17662 (N_17662,N_13507,N_10510);
nor U17663 (N_17663,N_13272,N_12987);
nor U17664 (N_17664,N_12623,N_13188);
nand U17665 (N_17665,N_13800,N_11509);
or U17666 (N_17666,N_11491,N_10987);
nand U17667 (N_17667,N_12342,N_12704);
nor U17668 (N_17668,N_11327,N_13003);
or U17669 (N_17669,N_14173,N_13783);
and U17670 (N_17670,N_10414,N_10533);
and U17671 (N_17671,N_14027,N_14770);
nand U17672 (N_17672,N_12303,N_13451);
nand U17673 (N_17673,N_12626,N_10508);
or U17674 (N_17674,N_10964,N_11147);
nor U17675 (N_17675,N_14991,N_14481);
nor U17676 (N_17676,N_12123,N_12837);
nor U17677 (N_17677,N_14235,N_14767);
xnor U17678 (N_17678,N_12950,N_12408);
nand U17679 (N_17679,N_13436,N_13008);
nand U17680 (N_17680,N_14233,N_12370);
nor U17681 (N_17681,N_11080,N_11108);
nor U17682 (N_17682,N_13544,N_10539);
and U17683 (N_17683,N_10053,N_14678);
and U17684 (N_17684,N_10496,N_14872);
or U17685 (N_17685,N_12343,N_13307);
or U17686 (N_17686,N_10104,N_11693);
nand U17687 (N_17687,N_11562,N_10579);
nor U17688 (N_17688,N_11848,N_10770);
or U17689 (N_17689,N_13708,N_10222);
and U17690 (N_17690,N_12916,N_12314);
nand U17691 (N_17691,N_12678,N_11969);
nor U17692 (N_17692,N_10123,N_10563);
nor U17693 (N_17693,N_11992,N_14376);
nor U17694 (N_17694,N_14331,N_14981);
and U17695 (N_17695,N_13828,N_10921);
nand U17696 (N_17696,N_14350,N_12883);
or U17697 (N_17697,N_11980,N_12129);
and U17698 (N_17698,N_14807,N_11928);
nand U17699 (N_17699,N_13849,N_12340);
xor U17700 (N_17700,N_11660,N_12153);
nand U17701 (N_17701,N_11677,N_11984);
xnor U17702 (N_17702,N_12004,N_10478);
xnor U17703 (N_17703,N_10029,N_13374);
nor U17704 (N_17704,N_13852,N_12043);
nor U17705 (N_17705,N_12253,N_14636);
and U17706 (N_17706,N_11932,N_12832);
and U17707 (N_17707,N_11048,N_13799);
xnor U17708 (N_17708,N_12152,N_14663);
nand U17709 (N_17709,N_14893,N_14640);
or U17710 (N_17710,N_14023,N_14470);
nor U17711 (N_17711,N_13531,N_14538);
nand U17712 (N_17712,N_13325,N_10644);
and U17713 (N_17713,N_10855,N_10010);
and U17714 (N_17714,N_11387,N_12545);
or U17715 (N_17715,N_14365,N_11298);
and U17716 (N_17716,N_10244,N_11293);
or U17717 (N_17717,N_10473,N_14012);
or U17718 (N_17718,N_12252,N_12385);
nor U17719 (N_17719,N_12956,N_14131);
or U17720 (N_17720,N_11459,N_13347);
nand U17721 (N_17721,N_14893,N_13687);
xnor U17722 (N_17722,N_11302,N_12311);
or U17723 (N_17723,N_10212,N_11817);
xnor U17724 (N_17724,N_10484,N_12341);
and U17725 (N_17725,N_13098,N_14456);
or U17726 (N_17726,N_14804,N_13964);
and U17727 (N_17727,N_12911,N_12045);
xnor U17728 (N_17728,N_10845,N_12073);
or U17729 (N_17729,N_14438,N_14664);
xor U17730 (N_17730,N_13690,N_10142);
and U17731 (N_17731,N_13427,N_14757);
xnor U17732 (N_17732,N_10048,N_14296);
or U17733 (N_17733,N_13298,N_11560);
or U17734 (N_17734,N_13870,N_14254);
and U17735 (N_17735,N_14108,N_14714);
nor U17736 (N_17736,N_13930,N_10883);
xor U17737 (N_17737,N_13348,N_11261);
and U17738 (N_17738,N_13203,N_14687);
nor U17739 (N_17739,N_10195,N_12202);
xnor U17740 (N_17740,N_11493,N_14525);
and U17741 (N_17741,N_11582,N_11229);
nor U17742 (N_17742,N_13694,N_11682);
and U17743 (N_17743,N_12170,N_13119);
nor U17744 (N_17744,N_12431,N_13295);
nor U17745 (N_17745,N_12072,N_12985);
nor U17746 (N_17746,N_12901,N_11345);
nor U17747 (N_17747,N_14531,N_11683);
nor U17748 (N_17748,N_11924,N_13161);
nor U17749 (N_17749,N_12908,N_10720);
nand U17750 (N_17750,N_11919,N_13993);
xnor U17751 (N_17751,N_11145,N_14089);
nand U17752 (N_17752,N_12515,N_14809);
xnor U17753 (N_17753,N_10229,N_13565);
and U17754 (N_17754,N_13360,N_13488);
nand U17755 (N_17755,N_10304,N_13746);
nand U17756 (N_17756,N_10132,N_14477);
xnor U17757 (N_17757,N_13548,N_11229);
xnor U17758 (N_17758,N_14634,N_12285);
and U17759 (N_17759,N_12083,N_10493);
xor U17760 (N_17760,N_13118,N_11230);
nand U17761 (N_17761,N_11308,N_12075);
or U17762 (N_17762,N_10561,N_10086);
nor U17763 (N_17763,N_12076,N_13513);
nand U17764 (N_17764,N_12839,N_14745);
nand U17765 (N_17765,N_10826,N_10608);
and U17766 (N_17766,N_10996,N_13784);
nand U17767 (N_17767,N_10212,N_12325);
nor U17768 (N_17768,N_12571,N_11494);
and U17769 (N_17769,N_12912,N_14351);
xnor U17770 (N_17770,N_11196,N_13034);
and U17771 (N_17771,N_13422,N_11270);
nand U17772 (N_17772,N_11588,N_14252);
nand U17773 (N_17773,N_13222,N_14367);
xnor U17774 (N_17774,N_10512,N_10645);
nor U17775 (N_17775,N_14136,N_11953);
xnor U17776 (N_17776,N_11064,N_14072);
nor U17777 (N_17777,N_13625,N_11442);
or U17778 (N_17778,N_10162,N_11202);
nor U17779 (N_17779,N_13246,N_11457);
or U17780 (N_17780,N_12301,N_12275);
or U17781 (N_17781,N_14397,N_12833);
or U17782 (N_17782,N_13872,N_14602);
nor U17783 (N_17783,N_10778,N_12049);
or U17784 (N_17784,N_13961,N_10381);
xor U17785 (N_17785,N_12075,N_13041);
or U17786 (N_17786,N_11055,N_10293);
xnor U17787 (N_17787,N_10111,N_11181);
and U17788 (N_17788,N_10370,N_14540);
or U17789 (N_17789,N_13184,N_12387);
nor U17790 (N_17790,N_12104,N_11743);
xor U17791 (N_17791,N_14256,N_14803);
nand U17792 (N_17792,N_13430,N_12087);
nand U17793 (N_17793,N_11196,N_11487);
or U17794 (N_17794,N_13395,N_11642);
and U17795 (N_17795,N_12544,N_10221);
and U17796 (N_17796,N_11449,N_14891);
nor U17797 (N_17797,N_13883,N_12761);
nand U17798 (N_17798,N_14753,N_14470);
or U17799 (N_17799,N_12457,N_14230);
nor U17800 (N_17800,N_10465,N_14024);
xor U17801 (N_17801,N_13391,N_14074);
xor U17802 (N_17802,N_11713,N_10877);
xnor U17803 (N_17803,N_10120,N_14684);
nor U17804 (N_17804,N_11321,N_14588);
nand U17805 (N_17805,N_14578,N_12084);
xor U17806 (N_17806,N_10521,N_11675);
and U17807 (N_17807,N_13138,N_10389);
or U17808 (N_17808,N_12866,N_11145);
xor U17809 (N_17809,N_14216,N_10248);
and U17810 (N_17810,N_14092,N_14283);
or U17811 (N_17811,N_10138,N_14835);
and U17812 (N_17812,N_11445,N_11583);
and U17813 (N_17813,N_13223,N_11206);
or U17814 (N_17814,N_12087,N_10299);
and U17815 (N_17815,N_10731,N_12277);
xnor U17816 (N_17816,N_11117,N_12707);
nor U17817 (N_17817,N_11683,N_13349);
nand U17818 (N_17818,N_11778,N_11266);
or U17819 (N_17819,N_12761,N_11951);
nor U17820 (N_17820,N_10402,N_14172);
nor U17821 (N_17821,N_12070,N_14382);
nand U17822 (N_17822,N_10014,N_13035);
and U17823 (N_17823,N_10282,N_12114);
or U17824 (N_17824,N_13634,N_11962);
or U17825 (N_17825,N_13680,N_11759);
and U17826 (N_17826,N_13980,N_13553);
or U17827 (N_17827,N_11450,N_10744);
and U17828 (N_17828,N_10518,N_13855);
and U17829 (N_17829,N_13861,N_13639);
nor U17830 (N_17830,N_13787,N_10377);
nor U17831 (N_17831,N_12525,N_12891);
or U17832 (N_17832,N_11373,N_10379);
and U17833 (N_17833,N_11665,N_11976);
and U17834 (N_17834,N_10861,N_10391);
nand U17835 (N_17835,N_13867,N_12862);
and U17836 (N_17836,N_10694,N_11853);
or U17837 (N_17837,N_12852,N_12906);
and U17838 (N_17838,N_13473,N_12794);
and U17839 (N_17839,N_12021,N_11343);
or U17840 (N_17840,N_13369,N_12046);
or U17841 (N_17841,N_13632,N_10399);
nor U17842 (N_17842,N_12283,N_10982);
nand U17843 (N_17843,N_11493,N_11640);
xnor U17844 (N_17844,N_14540,N_14014);
and U17845 (N_17845,N_14752,N_10067);
nand U17846 (N_17846,N_10214,N_10552);
nor U17847 (N_17847,N_11699,N_13775);
nor U17848 (N_17848,N_12223,N_13881);
nand U17849 (N_17849,N_13048,N_11460);
nand U17850 (N_17850,N_14479,N_10182);
and U17851 (N_17851,N_14803,N_13264);
and U17852 (N_17852,N_10903,N_14586);
xnor U17853 (N_17853,N_13447,N_12989);
xnor U17854 (N_17854,N_12037,N_14609);
nand U17855 (N_17855,N_13274,N_14545);
nor U17856 (N_17856,N_12137,N_11308);
and U17857 (N_17857,N_14072,N_11660);
xor U17858 (N_17858,N_12836,N_14913);
and U17859 (N_17859,N_13010,N_12619);
nor U17860 (N_17860,N_12905,N_14582);
or U17861 (N_17861,N_14055,N_12849);
nand U17862 (N_17862,N_11693,N_12069);
xor U17863 (N_17863,N_12116,N_14985);
nand U17864 (N_17864,N_12754,N_12421);
xnor U17865 (N_17865,N_13850,N_13337);
and U17866 (N_17866,N_12326,N_13427);
and U17867 (N_17867,N_10367,N_14894);
or U17868 (N_17868,N_13080,N_14016);
xnor U17869 (N_17869,N_14036,N_12593);
nand U17870 (N_17870,N_12428,N_10670);
xor U17871 (N_17871,N_14465,N_10778);
or U17872 (N_17872,N_14450,N_11064);
and U17873 (N_17873,N_13542,N_14962);
and U17874 (N_17874,N_10184,N_10213);
nand U17875 (N_17875,N_11227,N_10608);
nor U17876 (N_17876,N_12057,N_11146);
or U17877 (N_17877,N_13211,N_14344);
xnor U17878 (N_17878,N_10511,N_10247);
xor U17879 (N_17879,N_10050,N_14634);
nand U17880 (N_17880,N_11804,N_10750);
nand U17881 (N_17881,N_11480,N_14599);
xnor U17882 (N_17882,N_12446,N_13070);
nand U17883 (N_17883,N_14265,N_12735);
nor U17884 (N_17884,N_11176,N_11419);
nand U17885 (N_17885,N_12205,N_10021);
nor U17886 (N_17886,N_11045,N_13629);
or U17887 (N_17887,N_12366,N_12261);
or U17888 (N_17888,N_14778,N_13307);
or U17889 (N_17889,N_14206,N_13797);
or U17890 (N_17890,N_13041,N_10331);
nand U17891 (N_17891,N_14565,N_13212);
or U17892 (N_17892,N_13790,N_10462);
nor U17893 (N_17893,N_11444,N_11409);
and U17894 (N_17894,N_10988,N_10809);
or U17895 (N_17895,N_11091,N_10949);
or U17896 (N_17896,N_12512,N_12012);
nand U17897 (N_17897,N_14579,N_12325);
nor U17898 (N_17898,N_14795,N_14438);
xor U17899 (N_17899,N_11988,N_14626);
xor U17900 (N_17900,N_10851,N_11887);
and U17901 (N_17901,N_14787,N_13685);
or U17902 (N_17902,N_11127,N_11508);
nor U17903 (N_17903,N_11361,N_10016);
and U17904 (N_17904,N_12842,N_11328);
nand U17905 (N_17905,N_10044,N_10821);
nor U17906 (N_17906,N_12650,N_11145);
nor U17907 (N_17907,N_13726,N_13151);
and U17908 (N_17908,N_14313,N_14259);
xor U17909 (N_17909,N_13837,N_11869);
xnor U17910 (N_17910,N_13386,N_14915);
and U17911 (N_17911,N_13652,N_14907);
or U17912 (N_17912,N_13945,N_12642);
or U17913 (N_17913,N_11474,N_12928);
and U17914 (N_17914,N_14147,N_11477);
nor U17915 (N_17915,N_12274,N_13829);
nor U17916 (N_17916,N_14720,N_13616);
xor U17917 (N_17917,N_13930,N_11376);
or U17918 (N_17918,N_13496,N_14517);
nand U17919 (N_17919,N_14242,N_14490);
xor U17920 (N_17920,N_14357,N_14876);
xor U17921 (N_17921,N_10839,N_10569);
or U17922 (N_17922,N_12185,N_12900);
xnor U17923 (N_17923,N_12968,N_13214);
and U17924 (N_17924,N_13693,N_13570);
nand U17925 (N_17925,N_10299,N_13214);
nand U17926 (N_17926,N_11007,N_13372);
xor U17927 (N_17927,N_11054,N_10409);
or U17928 (N_17928,N_12428,N_13308);
or U17929 (N_17929,N_14225,N_13219);
xor U17930 (N_17930,N_11632,N_13634);
nand U17931 (N_17931,N_13465,N_10844);
nand U17932 (N_17932,N_14471,N_11873);
nor U17933 (N_17933,N_12709,N_10230);
nor U17934 (N_17934,N_11852,N_12717);
xor U17935 (N_17935,N_11558,N_12984);
nor U17936 (N_17936,N_14032,N_14843);
xor U17937 (N_17937,N_14781,N_12887);
xnor U17938 (N_17938,N_13501,N_11259);
and U17939 (N_17939,N_13561,N_12764);
nand U17940 (N_17940,N_14380,N_14528);
or U17941 (N_17941,N_14257,N_14627);
xnor U17942 (N_17942,N_13686,N_13179);
xor U17943 (N_17943,N_12955,N_14416);
nand U17944 (N_17944,N_14631,N_12738);
nor U17945 (N_17945,N_14096,N_12286);
nand U17946 (N_17946,N_13327,N_13022);
nand U17947 (N_17947,N_10743,N_11282);
and U17948 (N_17948,N_14739,N_11281);
nor U17949 (N_17949,N_12668,N_13145);
and U17950 (N_17950,N_12918,N_10549);
nor U17951 (N_17951,N_11559,N_11801);
nor U17952 (N_17952,N_13925,N_11395);
and U17953 (N_17953,N_10200,N_11849);
nor U17954 (N_17954,N_11842,N_14678);
nor U17955 (N_17955,N_13023,N_13117);
nor U17956 (N_17956,N_13890,N_14881);
nor U17957 (N_17957,N_13627,N_14842);
nand U17958 (N_17958,N_10791,N_14406);
or U17959 (N_17959,N_11985,N_14086);
nor U17960 (N_17960,N_11560,N_10965);
or U17961 (N_17961,N_11515,N_10932);
nand U17962 (N_17962,N_14205,N_12508);
and U17963 (N_17963,N_14337,N_11218);
xor U17964 (N_17964,N_10677,N_10594);
and U17965 (N_17965,N_10391,N_14067);
or U17966 (N_17966,N_14116,N_13654);
and U17967 (N_17967,N_13787,N_10438);
nand U17968 (N_17968,N_13910,N_11650);
nand U17969 (N_17969,N_13550,N_14214);
nand U17970 (N_17970,N_12405,N_11963);
xor U17971 (N_17971,N_12612,N_11055);
xor U17972 (N_17972,N_13298,N_14283);
xnor U17973 (N_17973,N_12727,N_13281);
nor U17974 (N_17974,N_14879,N_11144);
nor U17975 (N_17975,N_12299,N_10239);
nand U17976 (N_17976,N_10448,N_13262);
xor U17977 (N_17977,N_14115,N_12528);
or U17978 (N_17978,N_10815,N_13192);
and U17979 (N_17979,N_12953,N_14147);
xnor U17980 (N_17980,N_13907,N_13899);
xnor U17981 (N_17981,N_12910,N_10430);
nor U17982 (N_17982,N_13893,N_10641);
or U17983 (N_17983,N_14479,N_12398);
nor U17984 (N_17984,N_13821,N_10639);
and U17985 (N_17985,N_10198,N_14301);
or U17986 (N_17986,N_12531,N_11134);
and U17987 (N_17987,N_14689,N_11710);
xnor U17988 (N_17988,N_11908,N_12799);
xor U17989 (N_17989,N_14788,N_14817);
nand U17990 (N_17990,N_11395,N_13416);
nor U17991 (N_17991,N_11488,N_11232);
or U17992 (N_17992,N_10101,N_13935);
and U17993 (N_17993,N_14708,N_10863);
xnor U17994 (N_17994,N_10403,N_14381);
and U17995 (N_17995,N_11318,N_10448);
and U17996 (N_17996,N_11925,N_10644);
nand U17997 (N_17997,N_10829,N_14832);
or U17998 (N_17998,N_14839,N_13813);
nor U17999 (N_17999,N_12691,N_14772);
and U18000 (N_18000,N_12148,N_13385);
xnor U18001 (N_18001,N_14817,N_14225);
and U18002 (N_18002,N_14056,N_11469);
nor U18003 (N_18003,N_14161,N_14092);
and U18004 (N_18004,N_14737,N_12169);
nand U18005 (N_18005,N_11316,N_11903);
xnor U18006 (N_18006,N_14089,N_11246);
nand U18007 (N_18007,N_14644,N_11073);
nor U18008 (N_18008,N_11535,N_12344);
nand U18009 (N_18009,N_12915,N_14403);
xnor U18010 (N_18010,N_13311,N_10194);
nor U18011 (N_18011,N_10399,N_12692);
xor U18012 (N_18012,N_10050,N_14996);
nand U18013 (N_18013,N_11765,N_14161);
and U18014 (N_18014,N_12697,N_12481);
xor U18015 (N_18015,N_11242,N_10245);
or U18016 (N_18016,N_11986,N_12081);
nor U18017 (N_18017,N_10725,N_11411);
xor U18018 (N_18018,N_14362,N_13928);
or U18019 (N_18019,N_14628,N_13675);
nand U18020 (N_18020,N_13954,N_13739);
or U18021 (N_18021,N_12445,N_10073);
nor U18022 (N_18022,N_10378,N_10793);
xor U18023 (N_18023,N_10109,N_13515);
nand U18024 (N_18024,N_14150,N_14268);
xnor U18025 (N_18025,N_12856,N_11308);
and U18026 (N_18026,N_14860,N_12254);
nor U18027 (N_18027,N_12671,N_13555);
xnor U18028 (N_18028,N_14545,N_12960);
xor U18029 (N_18029,N_13507,N_12470);
nor U18030 (N_18030,N_11692,N_10163);
nand U18031 (N_18031,N_14706,N_14063);
nand U18032 (N_18032,N_14489,N_11428);
or U18033 (N_18033,N_12006,N_10320);
or U18034 (N_18034,N_13252,N_11208);
nand U18035 (N_18035,N_14499,N_10164);
nand U18036 (N_18036,N_10322,N_14750);
xor U18037 (N_18037,N_11706,N_13004);
xor U18038 (N_18038,N_13496,N_12116);
and U18039 (N_18039,N_13536,N_10225);
xnor U18040 (N_18040,N_14173,N_13544);
nor U18041 (N_18041,N_11699,N_12587);
and U18042 (N_18042,N_11903,N_14631);
nand U18043 (N_18043,N_12353,N_14828);
or U18044 (N_18044,N_12739,N_14879);
or U18045 (N_18045,N_14919,N_13814);
and U18046 (N_18046,N_13698,N_12445);
nor U18047 (N_18047,N_13821,N_12467);
or U18048 (N_18048,N_14686,N_11272);
and U18049 (N_18049,N_14459,N_11673);
nor U18050 (N_18050,N_13386,N_11171);
xnor U18051 (N_18051,N_10084,N_13056);
nor U18052 (N_18052,N_11402,N_12506);
xor U18053 (N_18053,N_13481,N_10756);
xnor U18054 (N_18054,N_11674,N_12222);
xnor U18055 (N_18055,N_13926,N_10722);
nand U18056 (N_18056,N_14622,N_13509);
xor U18057 (N_18057,N_10096,N_14665);
xor U18058 (N_18058,N_13448,N_13551);
or U18059 (N_18059,N_13364,N_14561);
or U18060 (N_18060,N_12756,N_12617);
and U18061 (N_18061,N_11509,N_11900);
nor U18062 (N_18062,N_13660,N_13739);
or U18063 (N_18063,N_13755,N_11104);
nor U18064 (N_18064,N_10910,N_12268);
nor U18065 (N_18065,N_12594,N_11543);
nor U18066 (N_18066,N_14117,N_11839);
nor U18067 (N_18067,N_14699,N_10785);
nor U18068 (N_18068,N_10686,N_12709);
nor U18069 (N_18069,N_13746,N_11124);
and U18070 (N_18070,N_12701,N_13909);
and U18071 (N_18071,N_14292,N_12890);
xnor U18072 (N_18072,N_13692,N_14010);
or U18073 (N_18073,N_14875,N_12289);
xor U18074 (N_18074,N_13198,N_12410);
xor U18075 (N_18075,N_13534,N_13827);
xnor U18076 (N_18076,N_14735,N_11197);
nand U18077 (N_18077,N_12304,N_11943);
xnor U18078 (N_18078,N_14560,N_13220);
nor U18079 (N_18079,N_11767,N_10850);
xor U18080 (N_18080,N_12637,N_10733);
and U18081 (N_18081,N_10232,N_13133);
and U18082 (N_18082,N_11441,N_12415);
xnor U18083 (N_18083,N_13287,N_13190);
nand U18084 (N_18084,N_14903,N_13994);
and U18085 (N_18085,N_14869,N_10274);
nor U18086 (N_18086,N_11275,N_11411);
nand U18087 (N_18087,N_10335,N_10983);
nand U18088 (N_18088,N_10022,N_10864);
nand U18089 (N_18089,N_11010,N_13225);
nand U18090 (N_18090,N_12127,N_11716);
nor U18091 (N_18091,N_14551,N_12608);
xnor U18092 (N_18092,N_13513,N_12871);
nor U18093 (N_18093,N_12555,N_11783);
or U18094 (N_18094,N_14939,N_14443);
xor U18095 (N_18095,N_14302,N_12648);
or U18096 (N_18096,N_13728,N_12547);
xnor U18097 (N_18097,N_13408,N_10825);
and U18098 (N_18098,N_12186,N_12309);
nor U18099 (N_18099,N_12115,N_10705);
or U18100 (N_18100,N_14888,N_10184);
and U18101 (N_18101,N_13312,N_13243);
or U18102 (N_18102,N_10512,N_12975);
or U18103 (N_18103,N_12119,N_11415);
nand U18104 (N_18104,N_14063,N_14689);
xnor U18105 (N_18105,N_14896,N_14347);
and U18106 (N_18106,N_10035,N_12982);
or U18107 (N_18107,N_12175,N_14899);
and U18108 (N_18108,N_14763,N_10687);
nand U18109 (N_18109,N_14074,N_13386);
xnor U18110 (N_18110,N_14899,N_11083);
nor U18111 (N_18111,N_14168,N_14829);
or U18112 (N_18112,N_14214,N_11978);
or U18113 (N_18113,N_10578,N_13731);
nand U18114 (N_18114,N_10426,N_14471);
nor U18115 (N_18115,N_12226,N_11516);
and U18116 (N_18116,N_10358,N_11115);
and U18117 (N_18117,N_12417,N_10235);
nor U18118 (N_18118,N_14293,N_12378);
nand U18119 (N_18119,N_12120,N_10192);
nor U18120 (N_18120,N_11403,N_10680);
xnor U18121 (N_18121,N_14036,N_14223);
nand U18122 (N_18122,N_14908,N_11026);
and U18123 (N_18123,N_13239,N_13590);
xor U18124 (N_18124,N_12775,N_14615);
and U18125 (N_18125,N_13233,N_12345);
and U18126 (N_18126,N_11247,N_13780);
nor U18127 (N_18127,N_11644,N_13554);
xnor U18128 (N_18128,N_13720,N_14574);
xnor U18129 (N_18129,N_14251,N_11400);
nor U18130 (N_18130,N_14431,N_10998);
or U18131 (N_18131,N_13612,N_13189);
nand U18132 (N_18132,N_14878,N_14074);
nand U18133 (N_18133,N_14607,N_11141);
nor U18134 (N_18134,N_11171,N_13962);
xor U18135 (N_18135,N_11216,N_10994);
nor U18136 (N_18136,N_14403,N_12668);
nor U18137 (N_18137,N_12315,N_11958);
or U18138 (N_18138,N_14961,N_13444);
xor U18139 (N_18139,N_11126,N_10090);
nor U18140 (N_18140,N_14955,N_10293);
nand U18141 (N_18141,N_12246,N_13690);
and U18142 (N_18142,N_12316,N_11627);
xnor U18143 (N_18143,N_10175,N_14087);
nand U18144 (N_18144,N_10265,N_12344);
or U18145 (N_18145,N_13234,N_11562);
and U18146 (N_18146,N_10789,N_10096);
or U18147 (N_18147,N_12802,N_12099);
xor U18148 (N_18148,N_10378,N_12211);
and U18149 (N_18149,N_10006,N_10574);
or U18150 (N_18150,N_10158,N_12796);
xnor U18151 (N_18151,N_14425,N_10266);
or U18152 (N_18152,N_10789,N_11738);
nor U18153 (N_18153,N_12524,N_12778);
nor U18154 (N_18154,N_10112,N_10177);
nor U18155 (N_18155,N_11150,N_12145);
nor U18156 (N_18156,N_13891,N_14963);
or U18157 (N_18157,N_10033,N_11779);
or U18158 (N_18158,N_12837,N_10332);
xnor U18159 (N_18159,N_11054,N_10578);
xnor U18160 (N_18160,N_11739,N_10638);
and U18161 (N_18161,N_14085,N_11077);
xor U18162 (N_18162,N_10519,N_11076);
nor U18163 (N_18163,N_12503,N_10416);
xor U18164 (N_18164,N_11540,N_14285);
nor U18165 (N_18165,N_11221,N_12592);
and U18166 (N_18166,N_11328,N_14570);
or U18167 (N_18167,N_13260,N_12137);
xor U18168 (N_18168,N_10561,N_11800);
or U18169 (N_18169,N_11660,N_10970);
xor U18170 (N_18170,N_10216,N_10673);
or U18171 (N_18171,N_10661,N_11507);
and U18172 (N_18172,N_14808,N_14551);
xnor U18173 (N_18173,N_11512,N_12774);
nand U18174 (N_18174,N_12219,N_12118);
and U18175 (N_18175,N_12036,N_14496);
xor U18176 (N_18176,N_13402,N_11279);
nand U18177 (N_18177,N_12711,N_14806);
and U18178 (N_18178,N_12698,N_13677);
xnor U18179 (N_18179,N_14252,N_14386);
and U18180 (N_18180,N_13059,N_14556);
xor U18181 (N_18181,N_14308,N_12806);
nor U18182 (N_18182,N_14592,N_14405);
nand U18183 (N_18183,N_10729,N_13528);
nand U18184 (N_18184,N_10937,N_13254);
xor U18185 (N_18185,N_12281,N_12116);
and U18186 (N_18186,N_11333,N_14590);
xnor U18187 (N_18187,N_11307,N_14984);
xnor U18188 (N_18188,N_11510,N_13267);
or U18189 (N_18189,N_11739,N_13483);
xnor U18190 (N_18190,N_11809,N_13999);
or U18191 (N_18191,N_14848,N_13894);
nand U18192 (N_18192,N_11495,N_14168);
nor U18193 (N_18193,N_10082,N_13728);
and U18194 (N_18194,N_12303,N_13376);
and U18195 (N_18195,N_14689,N_11422);
or U18196 (N_18196,N_12021,N_12875);
or U18197 (N_18197,N_14351,N_10450);
nor U18198 (N_18198,N_13664,N_14378);
xor U18199 (N_18199,N_13647,N_14304);
and U18200 (N_18200,N_13974,N_14463);
nor U18201 (N_18201,N_12194,N_10292);
nor U18202 (N_18202,N_14238,N_10635);
and U18203 (N_18203,N_10112,N_11264);
xor U18204 (N_18204,N_11464,N_13692);
nor U18205 (N_18205,N_11926,N_10908);
nand U18206 (N_18206,N_10486,N_14487);
and U18207 (N_18207,N_10122,N_14767);
xnor U18208 (N_18208,N_12104,N_10558);
xor U18209 (N_18209,N_10403,N_14996);
nor U18210 (N_18210,N_10307,N_11481);
xnor U18211 (N_18211,N_14697,N_13544);
and U18212 (N_18212,N_12330,N_10199);
nor U18213 (N_18213,N_14602,N_11825);
nor U18214 (N_18214,N_13073,N_13993);
nor U18215 (N_18215,N_12983,N_13085);
nor U18216 (N_18216,N_13189,N_12616);
or U18217 (N_18217,N_10951,N_13192);
and U18218 (N_18218,N_14916,N_14079);
nor U18219 (N_18219,N_11918,N_14290);
nand U18220 (N_18220,N_13228,N_12747);
or U18221 (N_18221,N_11904,N_11672);
xor U18222 (N_18222,N_14419,N_11399);
nor U18223 (N_18223,N_10582,N_14370);
nor U18224 (N_18224,N_10148,N_14199);
nor U18225 (N_18225,N_11432,N_13022);
nor U18226 (N_18226,N_10757,N_12006);
and U18227 (N_18227,N_14501,N_12789);
nand U18228 (N_18228,N_13005,N_11389);
nor U18229 (N_18229,N_13561,N_14262);
nor U18230 (N_18230,N_13294,N_12789);
xnor U18231 (N_18231,N_12794,N_12502);
xnor U18232 (N_18232,N_13164,N_13412);
or U18233 (N_18233,N_10504,N_11804);
and U18234 (N_18234,N_11236,N_10758);
nand U18235 (N_18235,N_14628,N_11230);
and U18236 (N_18236,N_13237,N_11602);
xnor U18237 (N_18237,N_12896,N_11386);
and U18238 (N_18238,N_14858,N_12113);
nand U18239 (N_18239,N_10189,N_12542);
nand U18240 (N_18240,N_10486,N_12152);
xnor U18241 (N_18241,N_14384,N_14730);
xor U18242 (N_18242,N_10991,N_13011);
or U18243 (N_18243,N_12951,N_11204);
nor U18244 (N_18244,N_11874,N_12895);
nor U18245 (N_18245,N_12044,N_14627);
or U18246 (N_18246,N_11502,N_11509);
nand U18247 (N_18247,N_12319,N_13489);
and U18248 (N_18248,N_11691,N_10786);
nor U18249 (N_18249,N_11594,N_13816);
and U18250 (N_18250,N_12057,N_12393);
and U18251 (N_18251,N_12126,N_14114);
xor U18252 (N_18252,N_12328,N_13141);
or U18253 (N_18253,N_14747,N_14454);
xor U18254 (N_18254,N_12118,N_14175);
xor U18255 (N_18255,N_12729,N_11978);
or U18256 (N_18256,N_14604,N_14291);
xnor U18257 (N_18257,N_11083,N_10518);
xor U18258 (N_18258,N_13977,N_13559);
nand U18259 (N_18259,N_12857,N_11604);
and U18260 (N_18260,N_11051,N_12084);
and U18261 (N_18261,N_14158,N_12327);
nor U18262 (N_18262,N_14888,N_11981);
xor U18263 (N_18263,N_12976,N_13933);
nor U18264 (N_18264,N_12271,N_10801);
or U18265 (N_18265,N_14328,N_13185);
and U18266 (N_18266,N_14057,N_13046);
nand U18267 (N_18267,N_14348,N_12172);
and U18268 (N_18268,N_12122,N_14722);
nor U18269 (N_18269,N_12800,N_10929);
and U18270 (N_18270,N_12726,N_12665);
nor U18271 (N_18271,N_12387,N_13289);
nand U18272 (N_18272,N_12376,N_11456);
xnor U18273 (N_18273,N_13344,N_11282);
and U18274 (N_18274,N_12912,N_11324);
xnor U18275 (N_18275,N_13653,N_14413);
or U18276 (N_18276,N_12310,N_14834);
and U18277 (N_18277,N_14275,N_11097);
nand U18278 (N_18278,N_12327,N_10853);
nor U18279 (N_18279,N_12211,N_13892);
or U18280 (N_18280,N_11698,N_13677);
and U18281 (N_18281,N_10752,N_13836);
and U18282 (N_18282,N_10997,N_11268);
nand U18283 (N_18283,N_13162,N_10472);
nand U18284 (N_18284,N_12648,N_14176);
nand U18285 (N_18285,N_13049,N_12028);
xnor U18286 (N_18286,N_14645,N_13760);
nand U18287 (N_18287,N_13141,N_11483);
nor U18288 (N_18288,N_14699,N_13620);
nand U18289 (N_18289,N_12737,N_10287);
nor U18290 (N_18290,N_11571,N_12459);
and U18291 (N_18291,N_13187,N_12671);
and U18292 (N_18292,N_12218,N_14448);
and U18293 (N_18293,N_13074,N_13250);
or U18294 (N_18294,N_14867,N_11204);
nand U18295 (N_18295,N_10546,N_13596);
nor U18296 (N_18296,N_10956,N_14864);
xnor U18297 (N_18297,N_11639,N_10625);
nor U18298 (N_18298,N_14718,N_11342);
nor U18299 (N_18299,N_11316,N_13723);
xor U18300 (N_18300,N_13984,N_10693);
nand U18301 (N_18301,N_11243,N_11413);
or U18302 (N_18302,N_11199,N_14832);
or U18303 (N_18303,N_14700,N_11736);
xor U18304 (N_18304,N_12031,N_12138);
or U18305 (N_18305,N_14980,N_12548);
nand U18306 (N_18306,N_11294,N_10692);
and U18307 (N_18307,N_12591,N_11191);
and U18308 (N_18308,N_13036,N_10897);
nor U18309 (N_18309,N_10007,N_11542);
nor U18310 (N_18310,N_13490,N_13210);
or U18311 (N_18311,N_11043,N_11354);
or U18312 (N_18312,N_10536,N_12482);
xnor U18313 (N_18313,N_14169,N_10283);
xor U18314 (N_18314,N_11818,N_10542);
nor U18315 (N_18315,N_11695,N_12123);
nand U18316 (N_18316,N_14066,N_12460);
nor U18317 (N_18317,N_14870,N_12620);
nand U18318 (N_18318,N_11651,N_12981);
nor U18319 (N_18319,N_13093,N_12254);
nor U18320 (N_18320,N_12291,N_11379);
nor U18321 (N_18321,N_12509,N_11654);
and U18322 (N_18322,N_11289,N_13988);
nand U18323 (N_18323,N_14657,N_11320);
or U18324 (N_18324,N_13459,N_11432);
nor U18325 (N_18325,N_12233,N_11503);
or U18326 (N_18326,N_14551,N_10861);
nor U18327 (N_18327,N_12000,N_13044);
nor U18328 (N_18328,N_12436,N_11073);
or U18329 (N_18329,N_13612,N_12467);
nand U18330 (N_18330,N_12136,N_10621);
xor U18331 (N_18331,N_13451,N_11152);
nand U18332 (N_18332,N_10726,N_13624);
nor U18333 (N_18333,N_11890,N_12037);
nor U18334 (N_18334,N_10990,N_13747);
or U18335 (N_18335,N_14185,N_10940);
or U18336 (N_18336,N_12797,N_14988);
xnor U18337 (N_18337,N_10758,N_13262);
nand U18338 (N_18338,N_13807,N_12748);
or U18339 (N_18339,N_11421,N_14974);
or U18340 (N_18340,N_10756,N_10207);
nor U18341 (N_18341,N_10150,N_12141);
xnor U18342 (N_18342,N_11642,N_10119);
nand U18343 (N_18343,N_10661,N_14230);
and U18344 (N_18344,N_13310,N_12412);
and U18345 (N_18345,N_12259,N_12875);
or U18346 (N_18346,N_13136,N_12139);
nor U18347 (N_18347,N_11955,N_10094);
nor U18348 (N_18348,N_12673,N_14085);
nor U18349 (N_18349,N_14729,N_12188);
and U18350 (N_18350,N_10206,N_11975);
and U18351 (N_18351,N_12068,N_12519);
xor U18352 (N_18352,N_10513,N_14106);
or U18353 (N_18353,N_14917,N_10410);
nand U18354 (N_18354,N_11623,N_14410);
or U18355 (N_18355,N_12675,N_13332);
nand U18356 (N_18356,N_11899,N_10828);
and U18357 (N_18357,N_13867,N_14858);
or U18358 (N_18358,N_11443,N_14745);
nor U18359 (N_18359,N_11941,N_12590);
nand U18360 (N_18360,N_13522,N_12114);
or U18361 (N_18361,N_13666,N_13789);
or U18362 (N_18362,N_11891,N_10182);
xnor U18363 (N_18363,N_12842,N_13996);
xor U18364 (N_18364,N_11933,N_10469);
nor U18365 (N_18365,N_14173,N_13384);
nand U18366 (N_18366,N_10315,N_14324);
nor U18367 (N_18367,N_14190,N_13379);
or U18368 (N_18368,N_12805,N_12780);
and U18369 (N_18369,N_11201,N_12150);
nor U18370 (N_18370,N_13141,N_13727);
or U18371 (N_18371,N_10774,N_12204);
or U18372 (N_18372,N_10622,N_13843);
xnor U18373 (N_18373,N_10143,N_10294);
and U18374 (N_18374,N_12400,N_12385);
nor U18375 (N_18375,N_12749,N_11714);
or U18376 (N_18376,N_10030,N_14471);
and U18377 (N_18377,N_12238,N_12868);
or U18378 (N_18378,N_10453,N_12462);
nor U18379 (N_18379,N_12964,N_13985);
and U18380 (N_18380,N_11432,N_10728);
xor U18381 (N_18381,N_12911,N_10898);
and U18382 (N_18382,N_10407,N_13911);
and U18383 (N_18383,N_13437,N_11526);
and U18384 (N_18384,N_13835,N_10636);
and U18385 (N_18385,N_10816,N_12558);
xor U18386 (N_18386,N_11587,N_12368);
and U18387 (N_18387,N_12403,N_12781);
nand U18388 (N_18388,N_12560,N_11672);
xnor U18389 (N_18389,N_11636,N_13374);
xnor U18390 (N_18390,N_13682,N_11620);
or U18391 (N_18391,N_14033,N_10381);
and U18392 (N_18392,N_13741,N_10178);
nor U18393 (N_18393,N_10314,N_12440);
xnor U18394 (N_18394,N_10521,N_14735);
and U18395 (N_18395,N_12544,N_11381);
and U18396 (N_18396,N_13593,N_13123);
or U18397 (N_18397,N_14549,N_14821);
nor U18398 (N_18398,N_11019,N_10776);
nor U18399 (N_18399,N_13293,N_13927);
nor U18400 (N_18400,N_11566,N_10006);
nor U18401 (N_18401,N_12681,N_10088);
or U18402 (N_18402,N_10764,N_14133);
and U18403 (N_18403,N_11495,N_12057);
xnor U18404 (N_18404,N_13277,N_12003);
xor U18405 (N_18405,N_12156,N_14837);
nand U18406 (N_18406,N_11612,N_12666);
nand U18407 (N_18407,N_14486,N_14587);
or U18408 (N_18408,N_14491,N_11881);
nor U18409 (N_18409,N_11336,N_13432);
xnor U18410 (N_18410,N_14458,N_10291);
or U18411 (N_18411,N_13168,N_14278);
xnor U18412 (N_18412,N_13138,N_13881);
or U18413 (N_18413,N_11602,N_12480);
nand U18414 (N_18414,N_12716,N_14112);
nand U18415 (N_18415,N_11699,N_11395);
and U18416 (N_18416,N_11687,N_11192);
nor U18417 (N_18417,N_14248,N_12483);
or U18418 (N_18418,N_10904,N_10962);
nand U18419 (N_18419,N_12849,N_10214);
xnor U18420 (N_18420,N_11762,N_12831);
xor U18421 (N_18421,N_12404,N_13662);
and U18422 (N_18422,N_14014,N_10423);
xnor U18423 (N_18423,N_14634,N_14728);
xnor U18424 (N_18424,N_12247,N_14257);
or U18425 (N_18425,N_14967,N_14744);
xor U18426 (N_18426,N_13212,N_10373);
nor U18427 (N_18427,N_14903,N_12510);
nand U18428 (N_18428,N_14235,N_11635);
and U18429 (N_18429,N_11857,N_10373);
and U18430 (N_18430,N_12094,N_13415);
nor U18431 (N_18431,N_12329,N_14587);
nor U18432 (N_18432,N_10457,N_13567);
xnor U18433 (N_18433,N_13832,N_12209);
and U18434 (N_18434,N_11570,N_13266);
nor U18435 (N_18435,N_11782,N_11554);
and U18436 (N_18436,N_12802,N_10064);
nand U18437 (N_18437,N_12775,N_12411);
and U18438 (N_18438,N_11471,N_10547);
nand U18439 (N_18439,N_12153,N_11837);
xnor U18440 (N_18440,N_11214,N_11074);
nor U18441 (N_18441,N_13620,N_10696);
or U18442 (N_18442,N_12967,N_10941);
nor U18443 (N_18443,N_10122,N_12310);
nand U18444 (N_18444,N_14802,N_11313);
nand U18445 (N_18445,N_14146,N_13345);
nand U18446 (N_18446,N_14107,N_12851);
xor U18447 (N_18447,N_14578,N_11660);
and U18448 (N_18448,N_14371,N_13522);
nor U18449 (N_18449,N_12892,N_13105);
nand U18450 (N_18450,N_14874,N_13375);
nand U18451 (N_18451,N_13417,N_13437);
and U18452 (N_18452,N_11774,N_10270);
and U18453 (N_18453,N_14235,N_14517);
and U18454 (N_18454,N_11472,N_10050);
nor U18455 (N_18455,N_10500,N_12473);
nor U18456 (N_18456,N_12245,N_12969);
or U18457 (N_18457,N_10341,N_10096);
xor U18458 (N_18458,N_11627,N_11020);
and U18459 (N_18459,N_10386,N_12461);
xnor U18460 (N_18460,N_12485,N_10656);
nor U18461 (N_18461,N_13580,N_13511);
or U18462 (N_18462,N_10356,N_13815);
nor U18463 (N_18463,N_10902,N_10378);
and U18464 (N_18464,N_12415,N_14188);
nor U18465 (N_18465,N_13441,N_11440);
nor U18466 (N_18466,N_12445,N_11948);
or U18467 (N_18467,N_14887,N_13062);
and U18468 (N_18468,N_10440,N_11435);
nand U18469 (N_18469,N_10297,N_10832);
nand U18470 (N_18470,N_12103,N_11589);
nor U18471 (N_18471,N_10116,N_12425);
nand U18472 (N_18472,N_11325,N_13135);
and U18473 (N_18473,N_11169,N_13778);
xor U18474 (N_18474,N_11973,N_12807);
nand U18475 (N_18475,N_12847,N_10416);
xnor U18476 (N_18476,N_11253,N_10341);
xor U18477 (N_18477,N_10083,N_13568);
nor U18478 (N_18478,N_12812,N_14286);
and U18479 (N_18479,N_11377,N_11229);
xor U18480 (N_18480,N_11052,N_10625);
xor U18481 (N_18481,N_14996,N_13234);
nand U18482 (N_18482,N_14517,N_14299);
or U18483 (N_18483,N_12394,N_12430);
nor U18484 (N_18484,N_10808,N_12746);
or U18485 (N_18485,N_14455,N_10949);
xnor U18486 (N_18486,N_13842,N_12699);
and U18487 (N_18487,N_10043,N_12377);
or U18488 (N_18488,N_11069,N_13236);
or U18489 (N_18489,N_12609,N_14252);
nand U18490 (N_18490,N_14194,N_13197);
nand U18491 (N_18491,N_10938,N_14445);
and U18492 (N_18492,N_10685,N_10243);
or U18493 (N_18493,N_12358,N_10237);
nor U18494 (N_18494,N_10775,N_12348);
nand U18495 (N_18495,N_10056,N_11654);
nand U18496 (N_18496,N_12257,N_13898);
and U18497 (N_18497,N_14598,N_13060);
and U18498 (N_18498,N_13249,N_12051);
or U18499 (N_18499,N_12144,N_11479);
nand U18500 (N_18500,N_13622,N_10590);
nand U18501 (N_18501,N_10388,N_13834);
and U18502 (N_18502,N_10485,N_12275);
nor U18503 (N_18503,N_12444,N_10331);
nand U18504 (N_18504,N_10564,N_14574);
nand U18505 (N_18505,N_10723,N_12440);
nor U18506 (N_18506,N_12341,N_13731);
nor U18507 (N_18507,N_12655,N_12407);
nand U18508 (N_18508,N_12370,N_11188);
and U18509 (N_18509,N_13120,N_13302);
xor U18510 (N_18510,N_14126,N_13004);
nor U18511 (N_18511,N_12582,N_10909);
nand U18512 (N_18512,N_10080,N_14823);
and U18513 (N_18513,N_12927,N_14959);
nand U18514 (N_18514,N_11027,N_11226);
nor U18515 (N_18515,N_12109,N_10799);
nand U18516 (N_18516,N_11672,N_12015);
and U18517 (N_18517,N_12550,N_12160);
and U18518 (N_18518,N_10346,N_13316);
and U18519 (N_18519,N_12691,N_12856);
and U18520 (N_18520,N_12543,N_13362);
xor U18521 (N_18521,N_14216,N_13647);
and U18522 (N_18522,N_13662,N_13670);
nand U18523 (N_18523,N_13251,N_10419);
xnor U18524 (N_18524,N_14097,N_11336);
and U18525 (N_18525,N_13641,N_13342);
and U18526 (N_18526,N_13556,N_14407);
xnor U18527 (N_18527,N_10901,N_10821);
nor U18528 (N_18528,N_14872,N_13563);
nor U18529 (N_18529,N_10212,N_14140);
nor U18530 (N_18530,N_11900,N_12954);
nor U18531 (N_18531,N_11301,N_14418);
xnor U18532 (N_18532,N_12413,N_13689);
or U18533 (N_18533,N_12838,N_10331);
xnor U18534 (N_18534,N_11395,N_12225);
nor U18535 (N_18535,N_11271,N_13578);
xor U18536 (N_18536,N_11389,N_12831);
nor U18537 (N_18537,N_12606,N_12543);
xor U18538 (N_18538,N_10460,N_11337);
and U18539 (N_18539,N_11868,N_10721);
and U18540 (N_18540,N_12026,N_12220);
or U18541 (N_18541,N_11171,N_12701);
nand U18542 (N_18542,N_10520,N_14547);
and U18543 (N_18543,N_10469,N_13572);
nand U18544 (N_18544,N_14832,N_10485);
or U18545 (N_18545,N_12300,N_11589);
or U18546 (N_18546,N_10702,N_14050);
or U18547 (N_18547,N_13244,N_12315);
xor U18548 (N_18548,N_13526,N_12205);
xor U18549 (N_18549,N_10344,N_11456);
or U18550 (N_18550,N_14194,N_11281);
nand U18551 (N_18551,N_12372,N_13073);
and U18552 (N_18552,N_11960,N_14354);
and U18553 (N_18553,N_11440,N_12787);
or U18554 (N_18554,N_12612,N_14305);
nand U18555 (N_18555,N_14255,N_14414);
xor U18556 (N_18556,N_13086,N_10186);
nand U18557 (N_18557,N_14868,N_14520);
and U18558 (N_18558,N_14054,N_10427);
nor U18559 (N_18559,N_10974,N_11804);
or U18560 (N_18560,N_11941,N_13934);
or U18561 (N_18561,N_11092,N_14196);
and U18562 (N_18562,N_11142,N_11163);
or U18563 (N_18563,N_11465,N_11574);
xor U18564 (N_18564,N_10636,N_12129);
nor U18565 (N_18565,N_10011,N_10072);
or U18566 (N_18566,N_13130,N_12310);
nand U18567 (N_18567,N_12457,N_12219);
xor U18568 (N_18568,N_13103,N_14438);
xnor U18569 (N_18569,N_13389,N_11000);
nor U18570 (N_18570,N_14737,N_13235);
nand U18571 (N_18571,N_10383,N_11990);
or U18572 (N_18572,N_11615,N_10113);
or U18573 (N_18573,N_14477,N_13388);
nand U18574 (N_18574,N_12083,N_14878);
nand U18575 (N_18575,N_13731,N_10243);
nor U18576 (N_18576,N_11872,N_10398);
nor U18577 (N_18577,N_11011,N_14978);
or U18578 (N_18578,N_11409,N_10949);
nand U18579 (N_18579,N_13169,N_11191);
xnor U18580 (N_18580,N_12763,N_10228);
nand U18581 (N_18581,N_14170,N_11289);
or U18582 (N_18582,N_14349,N_12347);
xor U18583 (N_18583,N_13160,N_11043);
nor U18584 (N_18584,N_11885,N_13084);
and U18585 (N_18585,N_11984,N_14747);
xor U18586 (N_18586,N_13932,N_13491);
and U18587 (N_18587,N_12785,N_12095);
and U18588 (N_18588,N_11492,N_12114);
nand U18589 (N_18589,N_10628,N_13299);
nor U18590 (N_18590,N_14104,N_11271);
xnor U18591 (N_18591,N_13023,N_10812);
nor U18592 (N_18592,N_10852,N_12488);
and U18593 (N_18593,N_14859,N_11912);
nand U18594 (N_18594,N_12615,N_10872);
nand U18595 (N_18595,N_12196,N_12411);
and U18596 (N_18596,N_10139,N_13816);
nand U18597 (N_18597,N_10527,N_11552);
xnor U18598 (N_18598,N_13610,N_14194);
or U18599 (N_18599,N_10591,N_12923);
xnor U18600 (N_18600,N_10891,N_13100);
or U18601 (N_18601,N_14450,N_14504);
xor U18602 (N_18602,N_13544,N_12647);
or U18603 (N_18603,N_11234,N_11416);
xor U18604 (N_18604,N_13624,N_14162);
or U18605 (N_18605,N_11735,N_12115);
nand U18606 (N_18606,N_10754,N_14559);
or U18607 (N_18607,N_13865,N_13924);
or U18608 (N_18608,N_13570,N_14308);
nor U18609 (N_18609,N_13942,N_11388);
nor U18610 (N_18610,N_10163,N_10339);
nor U18611 (N_18611,N_12265,N_13927);
nand U18612 (N_18612,N_13942,N_14111);
nor U18613 (N_18613,N_13419,N_14036);
nor U18614 (N_18614,N_10845,N_14383);
xor U18615 (N_18615,N_10847,N_12117);
xor U18616 (N_18616,N_10517,N_12246);
nor U18617 (N_18617,N_14553,N_11593);
nand U18618 (N_18618,N_13581,N_10506);
nor U18619 (N_18619,N_13844,N_12891);
and U18620 (N_18620,N_13686,N_11037);
and U18621 (N_18621,N_13005,N_14036);
xor U18622 (N_18622,N_13931,N_10740);
or U18623 (N_18623,N_14240,N_10439);
nand U18624 (N_18624,N_10663,N_10588);
nand U18625 (N_18625,N_14498,N_11738);
and U18626 (N_18626,N_11245,N_12110);
nor U18627 (N_18627,N_10762,N_11555);
nand U18628 (N_18628,N_10739,N_13664);
xnor U18629 (N_18629,N_11297,N_10598);
xor U18630 (N_18630,N_14344,N_13308);
xor U18631 (N_18631,N_11819,N_14514);
nor U18632 (N_18632,N_11276,N_10731);
or U18633 (N_18633,N_13237,N_14900);
or U18634 (N_18634,N_14565,N_12437);
xor U18635 (N_18635,N_11723,N_11825);
or U18636 (N_18636,N_11488,N_10330);
and U18637 (N_18637,N_11451,N_10531);
and U18638 (N_18638,N_10847,N_11839);
or U18639 (N_18639,N_12533,N_12404);
nand U18640 (N_18640,N_11811,N_11252);
nor U18641 (N_18641,N_11559,N_14423);
and U18642 (N_18642,N_10792,N_13005);
xnor U18643 (N_18643,N_14269,N_12588);
nor U18644 (N_18644,N_10116,N_10713);
and U18645 (N_18645,N_13625,N_10586);
or U18646 (N_18646,N_10718,N_11991);
xor U18647 (N_18647,N_10752,N_14228);
and U18648 (N_18648,N_14323,N_11357);
or U18649 (N_18649,N_10635,N_11744);
nor U18650 (N_18650,N_13963,N_11773);
or U18651 (N_18651,N_13545,N_11084);
and U18652 (N_18652,N_11322,N_14538);
xor U18653 (N_18653,N_10861,N_10384);
nand U18654 (N_18654,N_10424,N_12899);
xor U18655 (N_18655,N_11932,N_10797);
nand U18656 (N_18656,N_10099,N_14037);
xor U18657 (N_18657,N_14517,N_14198);
xor U18658 (N_18658,N_10707,N_12816);
nor U18659 (N_18659,N_14078,N_13554);
nand U18660 (N_18660,N_14493,N_14468);
nand U18661 (N_18661,N_13968,N_14961);
nor U18662 (N_18662,N_11627,N_12816);
xor U18663 (N_18663,N_11670,N_10384);
and U18664 (N_18664,N_14029,N_14632);
nor U18665 (N_18665,N_13518,N_13348);
xnor U18666 (N_18666,N_11238,N_11557);
or U18667 (N_18667,N_11605,N_10855);
or U18668 (N_18668,N_12994,N_10285);
or U18669 (N_18669,N_14016,N_13425);
nand U18670 (N_18670,N_13028,N_13063);
or U18671 (N_18671,N_12019,N_10944);
nor U18672 (N_18672,N_12501,N_12449);
or U18673 (N_18673,N_12122,N_10280);
or U18674 (N_18674,N_12608,N_13647);
xnor U18675 (N_18675,N_13873,N_14691);
or U18676 (N_18676,N_12677,N_12946);
xnor U18677 (N_18677,N_14145,N_11066);
or U18678 (N_18678,N_12961,N_12401);
or U18679 (N_18679,N_14271,N_14121);
or U18680 (N_18680,N_11297,N_11525);
nor U18681 (N_18681,N_11663,N_14778);
nand U18682 (N_18682,N_10788,N_10974);
xor U18683 (N_18683,N_14286,N_11372);
nor U18684 (N_18684,N_10749,N_14967);
nand U18685 (N_18685,N_14040,N_10800);
nand U18686 (N_18686,N_11659,N_10927);
or U18687 (N_18687,N_13664,N_14371);
or U18688 (N_18688,N_11888,N_13113);
or U18689 (N_18689,N_14899,N_12530);
nor U18690 (N_18690,N_12199,N_11639);
or U18691 (N_18691,N_13364,N_11351);
xnor U18692 (N_18692,N_13264,N_14614);
xnor U18693 (N_18693,N_13417,N_12292);
xnor U18694 (N_18694,N_12572,N_12986);
xnor U18695 (N_18695,N_13151,N_11890);
nor U18696 (N_18696,N_11578,N_14624);
and U18697 (N_18697,N_10413,N_10590);
or U18698 (N_18698,N_12914,N_11766);
nand U18699 (N_18699,N_13567,N_13683);
or U18700 (N_18700,N_10728,N_10649);
or U18701 (N_18701,N_12977,N_14008);
xnor U18702 (N_18702,N_11130,N_12989);
and U18703 (N_18703,N_13127,N_12831);
and U18704 (N_18704,N_11811,N_11278);
nand U18705 (N_18705,N_12315,N_11807);
xor U18706 (N_18706,N_10459,N_14500);
nand U18707 (N_18707,N_14310,N_14749);
nand U18708 (N_18708,N_12364,N_13432);
xnor U18709 (N_18709,N_12657,N_10796);
xor U18710 (N_18710,N_14528,N_11556);
or U18711 (N_18711,N_14526,N_11372);
or U18712 (N_18712,N_11609,N_14016);
or U18713 (N_18713,N_14628,N_14984);
nor U18714 (N_18714,N_12836,N_10683);
and U18715 (N_18715,N_13207,N_10334);
and U18716 (N_18716,N_12342,N_12110);
nor U18717 (N_18717,N_11829,N_13191);
and U18718 (N_18718,N_11171,N_14115);
and U18719 (N_18719,N_14818,N_14104);
or U18720 (N_18720,N_10527,N_10815);
nand U18721 (N_18721,N_11736,N_14123);
xor U18722 (N_18722,N_10577,N_11839);
and U18723 (N_18723,N_13849,N_10948);
xnor U18724 (N_18724,N_12622,N_14108);
or U18725 (N_18725,N_14422,N_14792);
nor U18726 (N_18726,N_11968,N_10999);
and U18727 (N_18727,N_11475,N_12245);
and U18728 (N_18728,N_11874,N_14379);
nand U18729 (N_18729,N_12064,N_11293);
or U18730 (N_18730,N_12228,N_11157);
and U18731 (N_18731,N_10567,N_13466);
and U18732 (N_18732,N_10629,N_12891);
xnor U18733 (N_18733,N_14103,N_12399);
and U18734 (N_18734,N_12528,N_11825);
xor U18735 (N_18735,N_11438,N_13775);
or U18736 (N_18736,N_12060,N_10574);
or U18737 (N_18737,N_12281,N_13752);
and U18738 (N_18738,N_10424,N_10062);
nor U18739 (N_18739,N_14089,N_14442);
or U18740 (N_18740,N_11943,N_12583);
nor U18741 (N_18741,N_12065,N_14922);
and U18742 (N_18742,N_12135,N_10453);
xor U18743 (N_18743,N_10369,N_10744);
nor U18744 (N_18744,N_12733,N_13548);
or U18745 (N_18745,N_14266,N_11340);
nor U18746 (N_18746,N_13107,N_10406);
or U18747 (N_18747,N_14704,N_10980);
xor U18748 (N_18748,N_11543,N_13507);
or U18749 (N_18749,N_14154,N_13175);
and U18750 (N_18750,N_12251,N_12602);
nand U18751 (N_18751,N_12360,N_14197);
or U18752 (N_18752,N_12785,N_13295);
nand U18753 (N_18753,N_13670,N_13482);
nand U18754 (N_18754,N_10646,N_10656);
or U18755 (N_18755,N_14716,N_11532);
nand U18756 (N_18756,N_10469,N_10040);
or U18757 (N_18757,N_14055,N_13689);
or U18758 (N_18758,N_14288,N_12178);
or U18759 (N_18759,N_10882,N_10743);
nand U18760 (N_18760,N_13954,N_10912);
nand U18761 (N_18761,N_14452,N_14140);
nand U18762 (N_18762,N_10358,N_11078);
and U18763 (N_18763,N_10634,N_14828);
nand U18764 (N_18764,N_11003,N_14478);
nor U18765 (N_18765,N_12889,N_11461);
or U18766 (N_18766,N_10792,N_13496);
nand U18767 (N_18767,N_10973,N_14820);
and U18768 (N_18768,N_13674,N_12516);
and U18769 (N_18769,N_11958,N_14963);
nor U18770 (N_18770,N_10601,N_12452);
nand U18771 (N_18771,N_11665,N_12985);
or U18772 (N_18772,N_11643,N_14868);
or U18773 (N_18773,N_11423,N_14797);
xor U18774 (N_18774,N_11169,N_11794);
or U18775 (N_18775,N_13687,N_11929);
or U18776 (N_18776,N_12741,N_14801);
nor U18777 (N_18777,N_10691,N_10485);
xor U18778 (N_18778,N_14327,N_12099);
nor U18779 (N_18779,N_13359,N_14539);
or U18780 (N_18780,N_11868,N_10729);
nor U18781 (N_18781,N_13038,N_11605);
nor U18782 (N_18782,N_12134,N_10700);
nand U18783 (N_18783,N_14836,N_12008);
nor U18784 (N_18784,N_11987,N_12570);
or U18785 (N_18785,N_11058,N_11737);
nor U18786 (N_18786,N_13787,N_11472);
xor U18787 (N_18787,N_14053,N_13849);
nand U18788 (N_18788,N_13395,N_11893);
nor U18789 (N_18789,N_10696,N_11137);
or U18790 (N_18790,N_10365,N_13466);
nor U18791 (N_18791,N_13467,N_14092);
xor U18792 (N_18792,N_13348,N_10378);
nor U18793 (N_18793,N_13790,N_12633);
nand U18794 (N_18794,N_10083,N_11384);
nor U18795 (N_18795,N_10305,N_14800);
xnor U18796 (N_18796,N_11648,N_12546);
and U18797 (N_18797,N_12181,N_11389);
nand U18798 (N_18798,N_11058,N_13133);
and U18799 (N_18799,N_12095,N_11922);
nor U18800 (N_18800,N_12608,N_11788);
or U18801 (N_18801,N_11999,N_11888);
xor U18802 (N_18802,N_13919,N_12904);
and U18803 (N_18803,N_11246,N_14000);
nand U18804 (N_18804,N_13957,N_10384);
nand U18805 (N_18805,N_14689,N_11715);
nor U18806 (N_18806,N_12181,N_14221);
nor U18807 (N_18807,N_12955,N_10061);
nand U18808 (N_18808,N_14144,N_10220);
xor U18809 (N_18809,N_10541,N_13271);
and U18810 (N_18810,N_12575,N_14101);
nand U18811 (N_18811,N_11774,N_12028);
or U18812 (N_18812,N_12689,N_14734);
and U18813 (N_18813,N_10255,N_13595);
or U18814 (N_18814,N_14506,N_13930);
nor U18815 (N_18815,N_11828,N_11264);
nand U18816 (N_18816,N_13730,N_10283);
nor U18817 (N_18817,N_12910,N_10957);
xnor U18818 (N_18818,N_13203,N_12075);
or U18819 (N_18819,N_11257,N_10133);
nand U18820 (N_18820,N_14605,N_13949);
nand U18821 (N_18821,N_12170,N_14885);
or U18822 (N_18822,N_11742,N_11080);
or U18823 (N_18823,N_12088,N_12531);
nor U18824 (N_18824,N_11199,N_12157);
nor U18825 (N_18825,N_14147,N_10244);
nor U18826 (N_18826,N_13404,N_10458);
nand U18827 (N_18827,N_12878,N_12208);
and U18828 (N_18828,N_13784,N_10801);
or U18829 (N_18829,N_14468,N_10584);
and U18830 (N_18830,N_14114,N_13796);
nor U18831 (N_18831,N_10401,N_10322);
or U18832 (N_18832,N_11069,N_13126);
xnor U18833 (N_18833,N_12122,N_13939);
nor U18834 (N_18834,N_10534,N_10482);
xor U18835 (N_18835,N_10393,N_10914);
nor U18836 (N_18836,N_11463,N_14410);
and U18837 (N_18837,N_12333,N_12265);
xnor U18838 (N_18838,N_14637,N_12275);
and U18839 (N_18839,N_14256,N_14765);
xor U18840 (N_18840,N_10925,N_10530);
or U18841 (N_18841,N_12676,N_13446);
or U18842 (N_18842,N_14486,N_10294);
nor U18843 (N_18843,N_14594,N_14214);
and U18844 (N_18844,N_12167,N_14316);
or U18845 (N_18845,N_13428,N_11684);
or U18846 (N_18846,N_13281,N_13975);
or U18847 (N_18847,N_10105,N_12085);
or U18848 (N_18848,N_11712,N_12703);
and U18849 (N_18849,N_11117,N_10887);
or U18850 (N_18850,N_12708,N_13650);
or U18851 (N_18851,N_11831,N_14315);
nand U18852 (N_18852,N_12701,N_13975);
xor U18853 (N_18853,N_10939,N_12966);
nand U18854 (N_18854,N_14578,N_10874);
nand U18855 (N_18855,N_14517,N_11155);
nand U18856 (N_18856,N_11240,N_10291);
nor U18857 (N_18857,N_13451,N_13077);
xor U18858 (N_18858,N_10818,N_13284);
or U18859 (N_18859,N_10059,N_10429);
or U18860 (N_18860,N_12471,N_14895);
nand U18861 (N_18861,N_12698,N_12330);
xnor U18862 (N_18862,N_14181,N_11488);
or U18863 (N_18863,N_10672,N_14551);
or U18864 (N_18864,N_12000,N_13135);
nor U18865 (N_18865,N_10872,N_14606);
and U18866 (N_18866,N_10219,N_12291);
nand U18867 (N_18867,N_10721,N_12652);
xor U18868 (N_18868,N_11184,N_10849);
or U18869 (N_18869,N_12378,N_13286);
and U18870 (N_18870,N_11222,N_13584);
nor U18871 (N_18871,N_12432,N_10176);
nor U18872 (N_18872,N_10739,N_11660);
nand U18873 (N_18873,N_14827,N_11376);
or U18874 (N_18874,N_12570,N_14226);
or U18875 (N_18875,N_14392,N_10263);
or U18876 (N_18876,N_11577,N_11056);
or U18877 (N_18877,N_13010,N_12790);
xor U18878 (N_18878,N_11654,N_10006);
and U18879 (N_18879,N_13850,N_14302);
or U18880 (N_18880,N_12306,N_13968);
xor U18881 (N_18881,N_11818,N_12292);
nor U18882 (N_18882,N_12787,N_14667);
nor U18883 (N_18883,N_13479,N_11898);
and U18884 (N_18884,N_12797,N_13999);
xnor U18885 (N_18885,N_13488,N_14584);
and U18886 (N_18886,N_12582,N_12833);
and U18887 (N_18887,N_11219,N_12304);
or U18888 (N_18888,N_12756,N_10745);
nor U18889 (N_18889,N_10064,N_14520);
xor U18890 (N_18890,N_11159,N_13519);
and U18891 (N_18891,N_14051,N_11915);
xnor U18892 (N_18892,N_12633,N_10083);
xor U18893 (N_18893,N_11837,N_11913);
xnor U18894 (N_18894,N_10716,N_13601);
and U18895 (N_18895,N_13408,N_14389);
xnor U18896 (N_18896,N_14785,N_11246);
nand U18897 (N_18897,N_12956,N_12717);
nor U18898 (N_18898,N_12025,N_13926);
or U18899 (N_18899,N_10574,N_14920);
and U18900 (N_18900,N_11798,N_11144);
nand U18901 (N_18901,N_14595,N_10488);
and U18902 (N_18902,N_13783,N_13896);
nor U18903 (N_18903,N_11162,N_13488);
or U18904 (N_18904,N_11115,N_10154);
nand U18905 (N_18905,N_14350,N_12763);
and U18906 (N_18906,N_10371,N_12275);
xor U18907 (N_18907,N_10036,N_10360);
xnor U18908 (N_18908,N_11003,N_12575);
and U18909 (N_18909,N_13689,N_10555);
xor U18910 (N_18910,N_13169,N_12326);
nand U18911 (N_18911,N_12937,N_12419);
nand U18912 (N_18912,N_11969,N_11779);
and U18913 (N_18913,N_14650,N_13784);
xnor U18914 (N_18914,N_13321,N_12998);
xor U18915 (N_18915,N_11603,N_10978);
or U18916 (N_18916,N_11777,N_11240);
and U18917 (N_18917,N_11155,N_10667);
xnor U18918 (N_18918,N_12623,N_10667);
nand U18919 (N_18919,N_14687,N_12934);
or U18920 (N_18920,N_12908,N_11431);
xnor U18921 (N_18921,N_10298,N_14494);
xor U18922 (N_18922,N_12640,N_14251);
and U18923 (N_18923,N_13723,N_11750);
or U18924 (N_18924,N_14492,N_13401);
nor U18925 (N_18925,N_13236,N_13846);
or U18926 (N_18926,N_12030,N_11910);
nor U18927 (N_18927,N_11638,N_11204);
and U18928 (N_18928,N_11692,N_12074);
nand U18929 (N_18929,N_10728,N_14584);
or U18930 (N_18930,N_13269,N_14379);
and U18931 (N_18931,N_13368,N_13063);
and U18932 (N_18932,N_14152,N_12018);
or U18933 (N_18933,N_13313,N_13368);
xor U18934 (N_18934,N_12508,N_11092);
nor U18935 (N_18935,N_10751,N_13916);
nand U18936 (N_18936,N_13209,N_12797);
or U18937 (N_18937,N_10598,N_12898);
or U18938 (N_18938,N_10949,N_11548);
xor U18939 (N_18939,N_13704,N_11896);
nand U18940 (N_18940,N_12230,N_12841);
nand U18941 (N_18941,N_14914,N_13931);
or U18942 (N_18942,N_11324,N_12057);
and U18943 (N_18943,N_11795,N_11346);
nand U18944 (N_18944,N_10272,N_10106);
xnor U18945 (N_18945,N_12064,N_13091);
or U18946 (N_18946,N_14682,N_14961);
or U18947 (N_18947,N_13535,N_11015);
and U18948 (N_18948,N_13031,N_14989);
nor U18949 (N_18949,N_14923,N_10178);
and U18950 (N_18950,N_11980,N_14369);
xor U18951 (N_18951,N_11498,N_11312);
or U18952 (N_18952,N_12525,N_12619);
and U18953 (N_18953,N_13911,N_13414);
nor U18954 (N_18954,N_14815,N_10856);
nor U18955 (N_18955,N_10694,N_14718);
nand U18956 (N_18956,N_11713,N_14856);
xor U18957 (N_18957,N_13841,N_13772);
nand U18958 (N_18958,N_10193,N_10434);
or U18959 (N_18959,N_12354,N_13108);
nand U18960 (N_18960,N_10252,N_12072);
xnor U18961 (N_18961,N_14030,N_14864);
or U18962 (N_18962,N_11571,N_12244);
nand U18963 (N_18963,N_13958,N_14695);
xnor U18964 (N_18964,N_13701,N_13219);
nor U18965 (N_18965,N_10481,N_11730);
or U18966 (N_18966,N_11066,N_12117);
and U18967 (N_18967,N_10286,N_12292);
and U18968 (N_18968,N_11785,N_13164);
and U18969 (N_18969,N_14157,N_11133);
and U18970 (N_18970,N_10819,N_11119);
nor U18971 (N_18971,N_11192,N_11205);
and U18972 (N_18972,N_10922,N_10673);
nand U18973 (N_18973,N_13131,N_11031);
or U18974 (N_18974,N_13023,N_12786);
and U18975 (N_18975,N_11910,N_12475);
xnor U18976 (N_18976,N_13784,N_14546);
xor U18977 (N_18977,N_13221,N_12043);
xnor U18978 (N_18978,N_13851,N_13998);
xor U18979 (N_18979,N_14208,N_12293);
nand U18980 (N_18980,N_14923,N_14306);
xor U18981 (N_18981,N_11642,N_14361);
nand U18982 (N_18982,N_12785,N_12469);
xor U18983 (N_18983,N_13141,N_12204);
xnor U18984 (N_18984,N_13148,N_12909);
or U18985 (N_18985,N_12054,N_11427);
or U18986 (N_18986,N_10199,N_14217);
and U18987 (N_18987,N_10242,N_10325);
or U18988 (N_18988,N_12106,N_11151);
nor U18989 (N_18989,N_11021,N_10720);
or U18990 (N_18990,N_13029,N_14130);
or U18991 (N_18991,N_14587,N_14470);
and U18992 (N_18992,N_14088,N_14067);
xnor U18993 (N_18993,N_11191,N_13338);
xor U18994 (N_18994,N_11430,N_11528);
nor U18995 (N_18995,N_11014,N_14145);
or U18996 (N_18996,N_14579,N_14977);
xnor U18997 (N_18997,N_13477,N_14235);
nor U18998 (N_18998,N_10396,N_10487);
or U18999 (N_18999,N_13931,N_11071);
nor U19000 (N_19000,N_11537,N_13619);
xnor U19001 (N_19001,N_12159,N_14068);
and U19002 (N_19002,N_10196,N_14394);
nor U19003 (N_19003,N_14222,N_13024);
and U19004 (N_19004,N_14794,N_12851);
xor U19005 (N_19005,N_10643,N_13142);
xnor U19006 (N_19006,N_14355,N_10778);
nor U19007 (N_19007,N_12193,N_11905);
nand U19008 (N_19008,N_11343,N_11451);
or U19009 (N_19009,N_10169,N_14068);
xor U19010 (N_19010,N_14367,N_13675);
nor U19011 (N_19011,N_14359,N_12998);
and U19012 (N_19012,N_10921,N_13491);
or U19013 (N_19013,N_14458,N_11858);
xor U19014 (N_19014,N_10602,N_11755);
xor U19015 (N_19015,N_12460,N_14074);
nand U19016 (N_19016,N_13642,N_13758);
and U19017 (N_19017,N_14719,N_10094);
xor U19018 (N_19018,N_10838,N_11248);
or U19019 (N_19019,N_10191,N_12537);
nand U19020 (N_19020,N_10264,N_10122);
nand U19021 (N_19021,N_11293,N_14997);
nand U19022 (N_19022,N_11809,N_10915);
nand U19023 (N_19023,N_14934,N_14297);
nor U19024 (N_19024,N_12748,N_11490);
or U19025 (N_19025,N_11009,N_13438);
nor U19026 (N_19026,N_12219,N_12692);
xnor U19027 (N_19027,N_10143,N_12692);
nand U19028 (N_19028,N_12433,N_11943);
nand U19029 (N_19029,N_13686,N_10105);
xnor U19030 (N_19030,N_10991,N_12099);
nand U19031 (N_19031,N_14725,N_14241);
nor U19032 (N_19032,N_13200,N_10246);
nand U19033 (N_19033,N_12458,N_14195);
nor U19034 (N_19034,N_14068,N_12592);
or U19035 (N_19035,N_14868,N_12774);
xnor U19036 (N_19036,N_13425,N_10657);
nor U19037 (N_19037,N_10056,N_10654);
nor U19038 (N_19038,N_13397,N_12540);
xnor U19039 (N_19039,N_11554,N_12236);
or U19040 (N_19040,N_10230,N_10191);
nand U19041 (N_19041,N_13538,N_13540);
or U19042 (N_19042,N_12858,N_14643);
and U19043 (N_19043,N_12567,N_12750);
or U19044 (N_19044,N_10132,N_11307);
nor U19045 (N_19045,N_14153,N_12185);
or U19046 (N_19046,N_12611,N_11260);
xor U19047 (N_19047,N_13907,N_14192);
and U19048 (N_19048,N_11248,N_12408);
and U19049 (N_19049,N_12865,N_12039);
or U19050 (N_19050,N_11138,N_13772);
and U19051 (N_19051,N_13031,N_10902);
or U19052 (N_19052,N_13607,N_14358);
nor U19053 (N_19053,N_11865,N_13813);
and U19054 (N_19054,N_12871,N_11260);
xor U19055 (N_19055,N_14219,N_13622);
xnor U19056 (N_19056,N_12780,N_13660);
nor U19057 (N_19057,N_11440,N_10437);
nor U19058 (N_19058,N_13930,N_14910);
nor U19059 (N_19059,N_14400,N_10929);
and U19060 (N_19060,N_13790,N_13106);
and U19061 (N_19061,N_14874,N_14934);
and U19062 (N_19062,N_11822,N_14068);
nand U19063 (N_19063,N_11037,N_11608);
xnor U19064 (N_19064,N_14233,N_13900);
nor U19065 (N_19065,N_12660,N_11876);
xor U19066 (N_19066,N_10612,N_12023);
nor U19067 (N_19067,N_11550,N_12985);
nand U19068 (N_19068,N_12227,N_14509);
nand U19069 (N_19069,N_14938,N_13161);
xor U19070 (N_19070,N_12088,N_10290);
xnor U19071 (N_19071,N_10675,N_10445);
nor U19072 (N_19072,N_11109,N_12678);
nand U19073 (N_19073,N_14679,N_14792);
nand U19074 (N_19074,N_14572,N_12817);
nand U19075 (N_19075,N_12873,N_11816);
nand U19076 (N_19076,N_12555,N_13118);
and U19077 (N_19077,N_14115,N_13667);
and U19078 (N_19078,N_14807,N_11102);
xor U19079 (N_19079,N_12866,N_11352);
xor U19080 (N_19080,N_11830,N_12949);
xor U19081 (N_19081,N_12686,N_14279);
xnor U19082 (N_19082,N_14313,N_10748);
nand U19083 (N_19083,N_13637,N_14953);
nor U19084 (N_19084,N_12053,N_12568);
nor U19085 (N_19085,N_13809,N_14400);
xor U19086 (N_19086,N_14230,N_13052);
or U19087 (N_19087,N_14296,N_12716);
nor U19088 (N_19088,N_13980,N_14720);
nor U19089 (N_19089,N_14853,N_10104);
nand U19090 (N_19090,N_10327,N_10632);
nand U19091 (N_19091,N_10742,N_11952);
nand U19092 (N_19092,N_10151,N_14611);
or U19093 (N_19093,N_10545,N_10702);
xnor U19094 (N_19094,N_13118,N_14230);
xor U19095 (N_19095,N_11559,N_10620);
xor U19096 (N_19096,N_10120,N_11354);
nand U19097 (N_19097,N_13777,N_12616);
nor U19098 (N_19098,N_14986,N_11032);
nor U19099 (N_19099,N_13822,N_10468);
or U19100 (N_19100,N_12728,N_12130);
nor U19101 (N_19101,N_13194,N_13990);
and U19102 (N_19102,N_14715,N_14698);
nor U19103 (N_19103,N_14531,N_11551);
and U19104 (N_19104,N_12413,N_12021);
nor U19105 (N_19105,N_10178,N_13444);
and U19106 (N_19106,N_12524,N_14401);
or U19107 (N_19107,N_10185,N_10217);
or U19108 (N_19108,N_10980,N_11356);
xnor U19109 (N_19109,N_11056,N_14474);
xnor U19110 (N_19110,N_13475,N_14398);
and U19111 (N_19111,N_10459,N_11923);
and U19112 (N_19112,N_11698,N_14534);
and U19113 (N_19113,N_10345,N_12336);
nand U19114 (N_19114,N_14793,N_14597);
nand U19115 (N_19115,N_14548,N_10504);
and U19116 (N_19116,N_10261,N_14295);
nand U19117 (N_19117,N_11128,N_10254);
and U19118 (N_19118,N_14210,N_10167);
or U19119 (N_19119,N_11648,N_11552);
nor U19120 (N_19120,N_14196,N_12755);
xor U19121 (N_19121,N_12005,N_14441);
or U19122 (N_19122,N_10866,N_14064);
and U19123 (N_19123,N_10849,N_10255);
xnor U19124 (N_19124,N_11300,N_11312);
or U19125 (N_19125,N_13231,N_12875);
xnor U19126 (N_19126,N_14599,N_14570);
xor U19127 (N_19127,N_13662,N_14632);
xor U19128 (N_19128,N_12096,N_14085);
or U19129 (N_19129,N_14801,N_10163);
xor U19130 (N_19130,N_14748,N_13928);
xnor U19131 (N_19131,N_11076,N_11168);
and U19132 (N_19132,N_11789,N_13805);
and U19133 (N_19133,N_14828,N_13174);
nor U19134 (N_19134,N_10097,N_11850);
or U19135 (N_19135,N_11958,N_10643);
nand U19136 (N_19136,N_13740,N_11887);
and U19137 (N_19137,N_13406,N_12691);
nand U19138 (N_19138,N_10021,N_10476);
and U19139 (N_19139,N_10350,N_12208);
xnor U19140 (N_19140,N_11135,N_14226);
nand U19141 (N_19141,N_13651,N_11951);
nand U19142 (N_19142,N_12508,N_10003);
and U19143 (N_19143,N_12599,N_11014);
and U19144 (N_19144,N_11820,N_13855);
and U19145 (N_19145,N_11226,N_11258);
or U19146 (N_19146,N_14208,N_11577);
and U19147 (N_19147,N_11935,N_10840);
nand U19148 (N_19148,N_11636,N_11954);
xnor U19149 (N_19149,N_10153,N_14183);
or U19150 (N_19150,N_13498,N_10722);
or U19151 (N_19151,N_13523,N_13654);
nand U19152 (N_19152,N_10938,N_11099);
or U19153 (N_19153,N_13237,N_13060);
nor U19154 (N_19154,N_11898,N_13439);
and U19155 (N_19155,N_12307,N_12944);
nand U19156 (N_19156,N_10894,N_10867);
nand U19157 (N_19157,N_11086,N_14842);
nor U19158 (N_19158,N_14234,N_14647);
or U19159 (N_19159,N_11251,N_10088);
nor U19160 (N_19160,N_11347,N_12959);
or U19161 (N_19161,N_12829,N_14026);
and U19162 (N_19162,N_12690,N_13153);
and U19163 (N_19163,N_10658,N_14647);
nor U19164 (N_19164,N_10059,N_12600);
and U19165 (N_19165,N_14503,N_12227);
nor U19166 (N_19166,N_14875,N_14817);
xor U19167 (N_19167,N_10640,N_11121);
xnor U19168 (N_19168,N_10578,N_11222);
nand U19169 (N_19169,N_13733,N_13307);
xnor U19170 (N_19170,N_10654,N_14853);
or U19171 (N_19171,N_14046,N_10236);
nor U19172 (N_19172,N_14752,N_11358);
xnor U19173 (N_19173,N_13736,N_14659);
nand U19174 (N_19174,N_12765,N_11853);
xnor U19175 (N_19175,N_11447,N_10458);
and U19176 (N_19176,N_12520,N_10165);
nor U19177 (N_19177,N_12695,N_11166);
xor U19178 (N_19178,N_10750,N_11056);
xor U19179 (N_19179,N_12859,N_14377);
xnor U19180 (N_19180,N_12367,N_13612);
nor U19181 (N_19181,N_12723,N_11894);
xnor U19182 (N_19182,N_10572,N_12243);
or U19183 (N_19183,N_12793,N_10717);
or U19184 (N_19184,N_12736,N_11400);
and U19185 (N_19185,N_14986,N_12925);
nand U19186 (N_19186,N_10146,N_13295);
xor U19187 (N_19187,N_11698,N_14789);
or U19188 (N_19188,N_13917,N_10079);
and U19189 (N_19189,N_11954,N_13325);
and U19190 (N_19190,N_11480,N_10679);
xor U19191 (N_19191,N_13226,N_10740);
xnor U19192 (N_19192,N_11116,N_10674);
nor U19193 (N_19193,N_10251,N_11836);
or U19194 (N_19194,N_11255,N_13920);
nor U19195 (N_19195,N_13565,N_13883);
and U19196 (N_19196,N_14535,N_13099);
xor U19197 (N_19197,N_13864,N_14217);
and U19198 (N_19198,N_12092,N_11880);
or U19199 (N_19199,N_11042,N_11962);
nand U19200 (N_19200,N_11215,N_11605);
nand U19201 (N_19201,N_12941,N_10089);
nand U19202 (N_19202,N_14819,N_10114);
xnor U19203 (N_19203,N_14696,N_12392);
nand U19204 (N_19204,N_10661,N_11214);
and U19205 (N_19205,N_12905,N_12767);
and U19206 (N_19206,N_14219,N_11021);
nand U19207 (N_19207,N_13080,N_10774);
or U19208 (N_19208,N_12377,N_12187);
or U19209 (N_19209,N_14723,N_11713);
and U19210 (N_19210,N_12175,N_12079);
nor U19211 (N_19211,N_14136,N_13170);
nor U19212 (N_19212,N_10697,N_10341);
nand U19213 (N_19213,N_11292,N_14308);
and U19214 (N_19214,N_13594,N_12967);
nand U19215 (N_19215,N_13338,N_11773);
xnor U19216 (N_19216,N_13423,N_12244);
xnor U19217 (N_19217,N_13425,N_14321);
nor U19218 (N_19218,N_10303,N_14524);
and U19219 (N_19219,N_14767,N_14453);
nand U19220 (N_19220,N_11553,N_12489);
or U19221 (N_19221,N_12926,N_14986);
or U19222 (N_19222,N_13969,N_13276);
xor U19223 (N_19223,N_14554,N_12679);
xnor U19224 (N_19224,N_12353,N_12749);
nand U19225 (N_19225,N_14453,N_13308);
or U19226 (N_19226,N_10992,N_13718);
or U19227 (N_19227,N_14223,N_14507);
nand U19228 (N_19228,N_11529,N_10869);
nor U19229 (N_19229,N_12950,N_12458);
xor U19230 (N_19230,N_10821,N_13245);
nor U19231 (N_19231,N_13627,N_10798);
nand U19232 (N_19232,N_12679,N_14598);
and U19233 (N_19233,N_12868,N_14268);
or U19234 (N_19234,N_14143,N_14040);
nor U19235 (N_19235,N_11464,N_10532);
xnor U19236 (N_19236,N_12813,N_11836);
nor U19237 (N_19237,N_10444,N_13399);
or U19238 (N_19238,N_13026,N_12769);
and U19239 (N_19239,N_14433,N_12627);
xnor U19240 (N_19240,N_13957,N_11825);
and U19241 (N_19241,N_14791,N_10944);
xnor U19242 (N_19242,N_14306,N_10628);
nand U19243 (N_19243,N_10337,N_10542);
or U19244 (N_19244,N_13562,N_10919);
nand U19245 (N_19245,N_10621,N_11365);
nand U19246 (N_19246,N_10799,N_10457);
nor U19247 (N_19247,N_11246,N_10038);
and U19248 (N_19248,N_10976,N_12269);
nor U19249 (N_19249,N_13847,N_12804);
nand U19250 (N_19250,N_13976,N_13475);
nand U19251 (N_19251,N_13350,N_13770);
xor U19252 (N_19252,N_14316,N_14521);
and U19253 (N_19253,N_11989,N_10371);
nor U19254 (N_19254,N_11975,N_14495);
and U19255 (N_19255,N_14913,N_11779);
nor U19256 (N_19256,N_14059,N_12396);
or U19257 (N_19257,N_11253,N_11164);
xnor U19258 (N_19258,N_11762,N_11692);
xnor U19259 (N_19259,N_10016,N_12272);
nor U19260 (N_19260,N_10952,N_11459);
xnor U19261 (N_19261,N_14248,N_14425);
nand U19262 (N_19262,N_10440,N_11100);
nand U19263 (N_19263,N_10966,N_10092);
or U19264 (N_19264,N_11573,N_14092);
nand U19265 (N_19265,N_10016,N_14743);
and U19266 (N_19266,N_13818,N_11345);
nand U19267 (N_19267,N_14149,N_11278);
nor U19268 (N_19268,N_12379,N_11757);
xor U19269 (N_19269,N_12794,N_12890);
and U19270 (N_19270,N_10932,N_10310);
nand U19271 (N_19271,N_11612,N_11041);
and U19272 (N_19272,N_13416,N_12754);
nor U19273 (N_19273,N_10153,N_14614);
and U19274 (N_19274,N_10775,N_11540);
and U19275 (N_19275,N_13739,N_12985);
or U19276 (N_19276,N_12081,N_14157);
and U19277 (N_19277,N_11832,N_14796);
xnor U19278 (N_19278,N_12111,N_13148);
nor U19279 (N_19279,N_10920,N_13062);
and U19280 (N_19280,N_12717,N_13055);
nand U19281 (N_19281,N_10804,N_12068);
xnor U19282 (N_19282,N_13193,N_13978);
and U19283 (N_19283,N_13764,N_12310);
nand U19284 (N_19284,N_14217,N_14148);
and U19285 (N_19285,N_10561,N_10535);
xor U19286 (N_19286,N_13841,N_10712);
nor U19287 (N_19287,N_10647,N_10127);
and U19288 (N_19288,N_12964,N_14947);
nand U19289 (N_19289,N_10323,N_11081);
nand U19290 (N_19290,N_11321,N_13607);
xnor U19291 (N_19291,N_14886,N_12270);
and U19292 (N_19292,N_10314,N_11365);
nand U19293 (N_19293,N_11642,N_10678);
xnor U19294 (N_19294,N_14231,N_14549);
and U19295 (N_19295,N_13097,N_14940);
and U19296 (N_19296,N_10511,N_14698);
nand U19297 (N_19297,N_12189,N_13164);
or U19298 (N_19298,N_12934,N_14100);
xnor U19299 (N_19299,N_14690,N_14320);
xor U19300 (N_19300,N_13096,N_14687);
nand U19301 (N_19301,N_13438,N_10433);
or U19302 (N_19302,N_11953,N_10051);
xnor U19303 (N_19303,N_11554,N_11656);
or U19304 (N_19304,N_11146,N_12372);
nand U19305 (N_19305,N_10505,N_13362);
nor U19306 (N_19306,N_11794,N_11291);
or U19307 (N_19307,N_12469,N_10247);
nor U19308 (N_19308,N_10194,N_14216);
or U19309 (N_19309,N_11315,N_13757);
xnor U19310 (N_19310,N_14817,N_11193);
xor U19311 (N_19311,N_14513,N_13370);
nand U19312 (N_19312,N_13703,N_11814);
nand U19313 (N_19313,N_10750,N_12387);
nand U19314 (N_19314,N_11788,N_10188);
and U19315 (N_19315,N_11334,N_13192);
or U19316 (N_19316,N_11075,N_12209);
or U19317 (N_19317,N_12424,N_14050);
nor U19318 (N_19318,N_14754,N_13089);
or U19319 (N_19319,N_14038,N_14011);
nor U19320 (N_19320,N_12864,N_13014);
and U19321 (N_19321,N_13882,N_10147);
nor U19322 (N_19322,N_12020,N_11003);
or U19323 (N_19323,N_14541,N_11014);
and U19324 (N_19324,N_11332,N_11823);
xnor U19325 (N_19325,N_14215,N_13675);
nor U19326 (N_19326,N_13059,N_11062);
and U19327 (N_19327,N_14555,N_11260);
and U19328 (N_19328,N_12160,N_13762);
or U19329 (N_19329,N_13398,N_12275);
nand U19330 (N_19330,N_10765,N_10771);
xnor U19331 (N_19331,N_12388,N_11586);
and U19332 (N_19332,N_11530,N_12015);
nand U19333 (N_19333,N_13066,N_13205);
or U19334 (N_19334,N_11487,N_14271);
nor U19335 (N_19335,N_14657,N_12459);
nand U19336 (N_19336,N_12348,N_10411);
xor U19337 (N_19337,N_11719,N_12090);
nand U19338 (N_19338,N_14430,N_11247);
nand U19339 (N_19339,N_10027,N_13986);
xnor U19340 (N_19340,N_11980,N_11189);
xnor U19341 (N_19341,N_13422,N_10624);
or U19342 (N_19342,N_12187,N_13887);
xor U19343 (N_19343,N_10062,N_13386);
nand U19344 (N_19344,N_13336,N_11607);
xor U19345 (N_19345,N_13756,N_12637);
or U19346 (N_19346,N_14603,N_10829);
and U19347 (N_19347,N_11405,N_13623);
xor U19348 (N_19348,N_10701,N_14397);
and U19349 (N_19349,N_11835,N_14341);
xnor U19350 (N_19350,N_13823,N_14960);
nor U19351 (N_19351,N_12181,N_11727);
or U19352 (N_19352,N_12766,N_14840);
nand U19353 (N_19353,N_13293,N_14062);
nor U19354 (N_19354,N_13970,N_13859);
xnor U19355 (N_19355,N_10968,N_11200);
and U19356 (N_19356,N_13506,N_13321);
or U19357 (N_19357,N_14342,N_11990);
nor U19358 (N_19358,N_11183,N_14026);
or U19359 (N_19359,N_13572,N_13229);
or U19360 (N_19360,N_11017,N_12918);
nand U19361 (N_19361,N_14687,N_10050);
or U19362 (N_19362,N_13765,N_11952);
nand U19363 (N_19363,N_14819,N_12305);
nor U19364 (N_19364,N_10408,N_10217);
nand U19365 (N_19365,N_12632,N_14808);
or U19366 (N_19366,N_14033,N_10235);
and U19367 (N_19367,N_12720,N_14911);
nor U19368 (N_19368,N_10436,N_12760);
nand U19369 (N_19369,N_14545,N_14217);
or U19370 (N_19370,N_14384,N_14237);
or U19371 (N_19371,N_13141,N_14646);
or U19372 (N_19372,N_11114,N_13525);
nand U19373 (N_19373,N_13227,N_14712);
xnor U19374 (N_19374,N_11092,N_12281);
nand U19375 (N_19375,N_11705,N_12438);
nand U19376 (N_19376,N_11410,N_12866);
and U19377 (N_19377,N_12174,N_14768);
or U19378 (N_19378,N_12006,N_11555);
nor U19379 (N_19379,N_10091,N_12270);
nor U19380 (N_19380,N_13656,N_11077);
and U19381 (N_19381,N_12157,N_10215);
and U19382 (N_19382,N_10344,N_14262);
nand U19383 (N_19383,N_13596,N_10081);
or U19384 (N_19384,N_14691,N_11887);
nor U19385 (N_19385,N_12694,N_10170);
and U19386 (N_19386,N_14353,N_13077);
or U19387 (N_19387,N_11358,N_13044);
xor U19388 (N_19388,N_13977,N_13366);
nor U19389 (N_19389,N_13471,N_13551);
nand U19390 (N_19390,N_14124,N_12563);
nand U19391 (N_19391,N_12461,N_14880);
nor U19392 (N_19392,N_10234,N_10863);
nor U19393 (N_19393,N_13262,N_10605);
nor U19394 (N_19394,N_10790,N_14326);
nand U19395 (N_19395,N_10231,N_12184);
nand U19396 (N_19396,N_11624,N_12427);
nand U19397 (N_19397,N_10579,N_10476);
nor U19398 (N_19398,N_11417,N_10768);
nor U19399 (N_19399,N_12821,N_14456);
or U19400 (N_19400,N_14512,N_14587);
nand U19401 (N_19401,N_14598,N_11692);
xor U19402 (N_19402,N_10623,N_10316);
nor U19403 (N_19403,N_13479,N_14928);
and U19404 (N_19404,N_10261,N_12053);
nor U19405 (N_19405,N_11128,N_14400);
or U19406 (N_19406,N_10040,N_13844);
nand U19407 (N_19407,N_11653,N_14764);
and U19408 (N_19408,N_13238,N_11717);
nand U19409 (N_19409,N_13491,N_13351);
and U19410 (N_19410,N_10564,N_13829);
xnor U19411 (N_19411,N_12662,N_14452);
and U19412 (N_19412,N_13411,N_12129);
nor U19413 (N_19413,N_13127,N_12184);
nor U19414 (N_19414,N_14279,N_14499);
nor U19415 (N_19415,N_10253,N_14600);
and U19416 (N_19416,N_11841,N_13167);
and U19417 (N_19417,N_14333,N_10940);
or U19418 (N_19418,N_12046,N_12199);
and U19419 (N_19419,N_11678,N_11967);
or U19420 (N_19420,N_10811,N_12694);
nand U19421 (N_19421,N_12469,N_10335);
nor U19422 (N_19422,N_13320,N_13803);
nor U19423 (N_19423,N_10853,N_12037);
and U19424 (N_19424,N_11736,N_12841);
xnor U19425 (N_19425,N_13718,N_13378);
nand U19426 (N_19426,N_11430,N_10291);
nand U19427 (N_19427,N_11331,N_10637);
nand U19428 (N_19428,N_10230,N_11812);
nand U19429 (N_19429,N_14140,N_13928);
and U19430 (N_19430,N_12388,N_13344);
nor U19431 (N_19431,N_13326,N_12203);
xor U19432 (N_19432,N_14442,N_13533);
or U19433 (N_19433,N_13440,N_13597);
nor U19434 (N_19434,N_10447,N_10051);
or U19435 (N_19435,N_13798,N_13416);
and U19436 (N_19436,N_13868,N_14852);
or U19437 (N_19437,N_11813,N_10362);
nand U19438 (N_19438,N_10555,N_11505);
nor U19439 (N_19439,N_11380,N_10326);
and U19440 (N_19440,N_12924,N_11194);
nand U19441 (N_19441,N_14686,N_12976);
and U19442 (N_19442,N_11449,N_14908);
nand U19443 (N_19443,N_14564,N_12339);
or U19444 (N_19444,N_13465,N_14604);
nand U19445 (N_19445,N_11263,N_12610);
and U19446 (N_19446,N_12397,N_13012);
xor U19447 (N_19447,N_10689,N_10369);
nand U19448 (N_19448,N_11344,N_14118);
nand U19449 (N_19449,N_13342,N_14558);
nor U19450 (N_19450,N_13323,N_11192);
or U19451 (N_19451,N_11312,N_11757);
and U19452 (N_19452,N_14099,N_14705);
nand U19453 (N_19453,N_13569,N_11018);
nor U19454 (N_19454,N_10970,N_14632);
or U19455 (N_19455,N_12053,N_14977);
nor U19456 (N_19456,N_14499,N_14650);
xnor U19457 (N_19457,N_13896,N_11146);
nor U19458 (N_19458,N_10982,N_11798);
nor U19459 (N_19459,N_11056,N_11537);
nand U19460 (N_19460,N_11740,N_14255);
nor U19461 (N_19461,N_10411,N_12711);
and U19462 (N_19462,N_11419,N_10367);
nand U19463 (N_19463,N_14742,N_12345);
and U19464 (N_19464,N_12463,N_13433);
or U19465 (N_19465,N_11186,N_10509);
nor U19466 (N_19466,N_14475,N_14417);
nand U19467 (N_19467,N_14625,N_14294);
or U19468 (N_19468,N_11932,N_10519);
xor U19469 (N_19469,N_12468,N_11082);
nor U19470 (N_19470,N_10140,N_12047);
xor U19471 (N_19471,N_12573,N_13395);
xnor U19472 (N_19472,N_14725,N_14887);
nor U19473 (N_19473,N_11004,N_12471);
and U19474 (N_19474,N_11727,N_10616);
or U19475 (N_19475,N_13465,N_12431);
nand U19476 (N_19476,N_14534,N_13101);
xor U19477 (N_19477,N_11255,N_11315);
nor U19478 (N_19478,N_10705,N_14614);
nand U19479 (N_19479,N_11650,N_14283);
and U19480 (N_19480,N_12817,N_14073);
or U19481 (N_19481,N_14548,N_14684);
xnor U19482 (N_19482,N_10343,N_12881);
nor U19483 (N_19483,N_12447,N_12658);
xnor U19484 (N_19484,N_11026,N_13956);
nand U19485 (N_19485,N_13472,N_12527);
nand U19486 (N_19486,N_12922,N_11319);
xor U19487 (N_19487,N_13085,N_14090);
or U19488 (N_19488,N_13695,N_10680);
xor U19489 (N_19489,N_10163,N_11574);
xor U19490 (N_19490,N_13868,N_13290);
xnor U19491 (N_19491,N_13661,N_10268);
nor U19492 (N_19492,N_14333,N_11710);
nor U19493 (N_19493,N_11609,N_10371);
or U19494 (N_19494,N_14055,N_10687);
xnor U19495 (N_19495,N_13009,N_10058);
nand U19496 (N_19496,N_12988,N_13946);
and U19497 (N_19497,N_12529,N_14393);
xnor U19498 (N_19498,N_11779,N_13703);
nand U19499 (N_19499,N_11121,N_14219);
and U19500 (N_19500,N_11538,N_14247);
xnor U19501 (N_19501,N_10603,N_13852);
xnor U19502 (N_19502,N_12039,N_10277);
or U19503 (N_19503,N_10357,N_10991);
nand U19504 (N_19504,N_12951,N_14323);
xor U19505 (N_19505,N_10420,N_14052);
nor U19506 (N_19506,N_14376,N_11713);
nand U19507 (N_19507,N_14491,N_13301);
nand U19508 (N_19508,N_14893,N_13302);
xor U19509 (N_19509,N_10723,N_14576);
or U19510 (N_19510,N_13233,N_10282);
xor U19511 (N_19511,N_11302,N_13154);
nor U19512 (N_19512,N_11935,N_12349);
xnor U19513 (N_19513,N_13015,N_14491);
xor U19514 (N_19514,N_13906,N_11071);
and U19515 (N_19515,N_11187,N_11169);
and U19516 (N_19516,N_11328,N_10788);
xnor U19517 (N_19517,N_14371,N_13647);
nor U19518 (N_19518,N_14371,N_13187);
or U19519 (N_19519,N_13941,N_11433);
nor U19520 (N_19520,N_14547,N_12308);
and U19521 (N_19521,N_14774,N_14547);
and U19522 (N_19522,N_12616,N_13115);
nand U19523 (N_19523,N_12039,N_13469);
or U19524 (N_19524,N_14952,N_14616);
and U19525 (N_19525,N_12480,N_10516);
or U19526 (N_19526,N_13118,N_13384);
nor U19527 (N_19527,N_13882,N_13228);
or U19528 (N_19528,N_12389,N_13881);
xor U19529 (N_19529,N_12511,N_10030);
or U19530 (N_19530,N_10511,N_13396);
nand U19531 (N_19531,N_12504,N_13694);
xor U19532 (N_19532,N_11014,N_14548);
or U19533 (N_19533,N_10977,N_11651);
nor U19534 (N_19534,N_14767,N_13268);
nand U19535 (N_19535,N_14749,N_14763);
xnor U19536 (N_19536,N_11480,N_11284);
nor U19537 (N_19537,N_13905,N_10127);
and U19538 (N_19538,N_10718,N_11472);
and U19539 (N_19539,N_14600,N_13663);
nor U19540 (N_19540,N_12835,N_10926);
and U19541 (N_19541,N_12473,N_10950);
nor U19542 (N_19542,N_13051,N_14357);
nand U19543 (N_19543,N_13075,N_13932);
xnor U19544 (N_19544,N_11028,N_12376);
and U19545 (N_19545,N_14587,N_14901);
nand U19546 (N_19546,N_14758,N_11752);
or U19547 (N_19547,N_14607,N_11452);
and U19548 (N_19548,N_13088,N_14833);
and U19549 (N_19549,N_10747,N_13769);
xor U19550 (N_19550,N_11653,N_13244);
nand U19551 (N_19551,N_12377,N_14437);
xor U19552 (N_19552,N_14207,N_10399);
and U19553 (N_19553,N_14257,N_14167);
nand U19554 (N_19554,N_11847,N_13772);
nor U19555 (N_19555,N_14176,N_11868);
nor U19556 (N_19556,N_14973,N_13188);
nor U19557 (N_19557,N_13327,N_13875);
or U19558 (N_19558,N_13343,N_14398);
nor U19559 (N_19559,N_11268,N_12303);
nand U19560 (N_19560,N_12735,N_11912);
xnor U19561 (N_19561,N_10764,N_13549);
and U19562 (N_19562,N_10535,N_13697);
xor U19563 (N_19563,N_12422,N_11380);
nor U19564 (N_19564,N_11674,N_10089);
nand U19565 (N_19565,N_13646,N_13480);
and U19566 (N_19566,N_10119,N_10386);
xnor U19567 (N_19567,N_10725,N_14139);
nor U19568 (N_19568,N_14379,N_11661);
and U19569 (N_19569,N_14033,N_11924);
nor U19570 (N_19570,N_12881,N_14543);
xor U19571 (N_19571,N_10421,N_14814);
nor U19572 (N_19572,N_12583,N_11851);
or U19573 (N_19573,N_11058,N_12127);
and U19574 (N_19574,N_13557,N_12042);
xor U19575 (N_19575,N_10334,N_13935);
and U19576 (N_19576,N_14401,N_12265);
nand U19577 (N_19577,N_11541,N_14775);
xor U19578 (N_19578,N_14944,N_14702);
nand U19579 (N_19579,N_13195,N_12432);
xnor U19580 (N_19580,N_13293,N_10750);
nor U19581 (N_19581,N_12431,N_11245);
xor U19582 (N_19582,N_11580,N_12963);
nor U19583 (N_19583,N_14742,N_10085);
xnor U19584 (N_19584,N_11437,N_12457);
and U19585 (N_19585,N_10818,N_13315);
and U19586 (N_19586,N_10145,N_14070);
and U19587 (N_19587,N_12860,N_12025);
nor U19588 (N_19588,N_14184,N_14739);
nand U19589 (N_19589,N_10763,N_14220);
or U19590 (N_19590,N_11217,N_14051);
or U19591 (N_19591,N_13000,N_14781);
xnor U19592 (N_19592,N_14162,N_13362);
or U19593 (N_19593,N_14076,N_12841);
nor U19594 (N_19594,N_14148,N_11578);
nor U19595 (N_19595,N_13360,N_12921);
and U19596 (N_19596,N_11532,N_14741);
and U19597 (N_19597,N_13398,N_11449);
or U19598 (N_19598,N_12088,N_10695);
and U19599 (N_19599,N_11978,N_13424);
or U19600 (N_19600,N_10636,N_13603);
nand U19601 (N_19601,N_13626,N_13085);
or U19602 (N_19602,N_10932,N_10568);
and U19603 (N_19603,N_11510,N_13026);
nor U19604 (N_19604,N_11311,N_14325);
nand U19605 (N_19605,N_11305,N_13210);
nand U19606 (N_19606,N_12529,N_13974);
nand U19607 (N_19607,N_10545,N_12801);
or U19608 (N_19608,N_12311,N_11574);
and U19609 (N_19609,N_13281,N_14555);
and U19610 (N_19610,N_12884,N_10271);
nand U19611 (N_19611,N_14365,N_13304);
xnor U19612 (N_19612,N_12397,N_12697);
nand U19613 (N_19613,N_14551,N_13680);
xor U19614 (N_19614,N_13065,N_11723);
xnor U19615 (N_19615,N_14228,N_10165);
nand U19616 (N_19616,N_10932,N_14046);
or U19617 (N_19617,N_12519,N_13761);
xnor U19618 (N_19618,N_11828,N_13943);
nand U19619 (N_19619,N_12148,N_13007);
xnor U19620 (N_19620,N_12368,N_14848);
or U19621 (N_19621,N_10675,N_12086);
xnor U19622 (N_19622,N_12742,N_11407);
xnor U19623 (N_19623,N_12336,N_11266);
nor U19624 (N_19624,N_10251,N_10469);
nand U19625 (N_19625,N_11693,N_12230);
and U19626 (N_19626,N_14024,N_14107);
and U19627 (N_19627,N_12222,N_10716);
nand U19628 (N_19628,N_12674,N_13272);
xor U19629 (N_19629,N_10876,N_12863);
xor U19630 (N_19630,N_13292,N_12945);
or U19631 (N_19631,N_14159,N_11019);
xor U19632 (N_19632,N_13487,N_14111);
nand U19633 (N_19633,N_11226,N_13062);
nor U19634 (N_19634,N_12822,N_14417);
nand U19635 (N_19635,N_13296,N_14937);
nor U19636 (N_19636,N_12406,N_12369);
nor U19637 (N_19637,N_10200,N_12591);
nor U19638 (N_19638,N_10856,N_12743);
nand U19639 (N_19639,N_13133,N_14182);
xor U19640 (N_19640,N_10828,N_13825);
nor U19641 (N_19641,N_14971,N_11940);
or U19642 (N_19642,N_11830,N_11493);
and U19643 (N_19643,N_13928,N_11943);
or U19644 (N_19644,N_14640,N_11070);
nor U19645 (N_19645,N_14450,N_12758);
and U19646 (N_19646,N_14147,N_10766);
and U19647 (N_19647,N_11956,N_10859);
and U19648 (N_19648,N_10547,N_12271);
nor U19649 (N_19649,N_14152,N_13752);
nor U19650 (N_19650,N_12771,N_12846);
nand U19651 (N_19651,N_12303,N_10443);
xnor U19652 (N_19652,N_14727,N_13708);
nand U19653 (N_19653,N_10413,N_14711);
nor U19654 (N_19654,N_10119,N_14088);
and U19655 (N_19655,N_10382,N_11427);
nor U19656 (N_19656,N_14936,N_13661);
or U19657 (N_19657,N_12669,N_10552);
nor U19658 (N_19658,N_11874,N_13586);
nor U19659 (N_19659,N_10075,N_12245);
nand U19660 (N_19660,N_14040,N_13466);
and U19661 (N_19661,N_10102,N_13093);
nor U19662 (N_19662,N_12634,N_13343);
and U19663 (N_19663,N_14804,N_10347);
xor U19664 (N_19664,N_10506,N_10793);
or U19665 (N_19665,N_14235,N_11619);
xnor U19666 (N_19666,N_11534,N_12531);
and U19667 (N_19667,N_12678,N_13214);
or U19668 (N_19668,N_13389,N_14332);
and U19669 (N_19669,N_14719,N_12976);
or U19670 (N_19670,N_12645,N_11099);
nand U19671 (N_19671,N_11022,N_10831);
nor U19672 (N_19672,N_10009,N_13227);
nand U19673 (N_19673,N_11769,N_11094);
nor U19674 (N_19674,N_12395,N_13745);
xor U19675 (N_19675,N_11575,N_13577);
and U19676 (N_19676,N_14732,N_10058);
nor U19677 (N_19677,N_14869,N_12477);
xor U19678 (N_19678,N_12617,N_13494);
nor U19679 (N_19679,N_14783,N_14581);
or U19680 (N_19680,N_13974,N_13694);
xnor U19681 (N_19681,N_10527,N_10366);
and U19682 (N_19682,N_10985,N_14507);
and U19683 (N_19683,N_12528,N_12211);
xnor U19684 (N_19684,N_11328,N_14225);
xor U19685 (N_19685,N_13870,N_11785);
nor U19686 (N_19686,N_13472,N_14551);
xnor U19687 (N_19687,N_12574,N_13176);
xor U19688 (N_19688,N_14202,N_11011);
nand U19689 (N_19689,N_11402,N_13450);
nand U19690 (N_19690,N_13112,N_10552);
or U19691 (N_19691,N_13324,N_14967);
nor U19692 (N_19692,N_13919,N_14180);
nand U19693 (N_19693,N_11168,N_11763);
or U19694 (N_19694,N_12808,N_10169);
xor U19695 (N_19695,N_13378,N_14038);
nand U19696 (N_19696,N_11556,N_11735);
and U19697 (N_19697,N_10149,N_12388);
xor U19698 (N_19698,N_12610,N_10883);
xor U19699 (N_19699,N_13197,N_11900);
nand U19700 (N_19700,N_14701,N_12506);
nor U19701 (N_19701,N_12807,N_14692);
nor U19702 (N_19702,N_13714,N_10300);
nand U19703 (N_19703,N_10950,N_12227);
or U19704 (N_19704,N_10024,N_12180);
or U19705 (N_19705,N_12158,N_10096);
or U19706 (N_19706,N_13363,N_13312);
xnor U19707 (N_19707,N_14793,N_14980);
nand U19708 (N_19708,N_13286,N_11679);
nand U19709 (N_19709,N_14919,N_12272);
xor U19710 (N_19710,N_11291,N_12092);
nor U19711 (N_19711,N_13873,N_11718);
nand U19712 (N_19712,N_11318,N_11160);
or U19713 (N_19713,N_12487,N_10536);
nand U19714 (N_19714,N_13138,N_12239);
or U19715 (N_19715,N_12041,N_11450);
xor U19716 (N_19716,N_11162,N_14815);
or U19717 (N_19717,N_10407,N_12263);
xor U19718 (N_19718,N_13337,N_11048);
nand U19719 (N_19719,N_11037,N_11469);
nand U19720 (N_19720,N_12141,N_14338);
xnor U19721 (N_19721,N_12609,N_14151);
nor U19722 (N_19722,N_10893,N_12889);
xor U19723 (N_19723,N_10464,N_13424);
nor U19724 (N_19724,N_13308,N_12240);
nor U19725 (N_19725,N_10375,N_13418);
and U19726 (N_19726,N_11585,N_14702);
and U19727 (N_19727,N_12514,N_10329);
nor U19728 (N_19728,N_12916,N_12499);
nand U19729 (N_19729,N_14742,N_12842);
nor U19730 (N_19730,N_12891,N_11730);
xor U19731 (N_19731,N_11615,N_14172);
or U19732 (N_19732,N_14918,N_13430);
nand U19733 (N_19733,N_14243,N_14832);
or U19734 (N_19734,N_14060,N_12206);
xor U19735 (N_19735,N_12013,N_13118);
xor U19736 (N_19736,N_14357,N_13851);
nand U19737 (N_19737,N_14241,N_10740);
and U19738 (N_19738,N_13722,N_10190);
nand U19739 (N_19739,N_14312,N_10902);
nand U19740 (N_19740,N_10117,N_14132);
or U19741 (N_19741,N_14021,N_14997);
or U19742 (N_19742,N_14948,N_14647);
xnor U19743 (N_19743,N_12183,N_10485);
or U19744 (N_19744,N_14804,N_11088);
or U19745 (N_19745,N_12347,N_13291);
and U19746 (N_19746,N_11302,N_12052);
xor U19747 (N_19747,N_13129,N_13677);
or U19748 (N_19748,N_11563,N_13058);
and U19749 (N_19749,N_11312,N_14147);
xor U19750 (N_19750,N_11305,N_14523);
and U19751 (N_19751,N_10579,N_13084);
nand U19752 (N_19752,N_11987,N_13473);
nor U19753 (N_19753,N_13242,N_14538);
and U19754 (N_19754,N_12541,N_12619);
or U19755 (N_19755,N_11354,N_11568);
nand U19756 (N_19756,N_11332,N_14902);
or U19757 (N_19757,N_11398,N_14532);
and U19758 (N_19758,N_11673,N_12308);
and U19759 (N_19759,N_13340,N_13455);
nand U19760 (N_19760,N_13244,N_13567);
or U19761 (N_19761,N_14055,N_13756);
xor U19762 (N_19762,N_11900,N_10405);
xor U19763 (N_19763,N_12898,N_11081);
nand U19764 (N_19764,N_14054,N_13844);
or U19765 (N_19765,N_10426,N_13815);
xor U19766 (N_19766,N_14227,N_14791);
xor U19767 (N_19767,N_10937,N_11989);
or U19768 (N_19768,N_14883,N_10775);
nand U19769 (N_19769,N_14647,N_11162);
nor U19770 (N_19770,N_12427,N_14080);
nor U19771 (N_19771,N_14968,N_11717);
and U19772 (N_19772,N_14108,N_13990);
nand U19773 (N_19773,N_14692,N_14611);
and U19774 (N_19774,N_12765,N_11666);
nor U19775 (N_19775,N_14448,N_14547);
nor U19776 (N_19776,N_12961,N_10223);
xor U19777 (N_19777,N_14855,N_10618);
xor U19778 (N_19778,N_10512,N_14230);
and U19779 (N_19779,N_12464,N_10914);
xnor U19780 (N_19780,N_11966,N_14243);
and U19781 (N_19781,N_13690,N_11788);
nor U19782 (N_19782,N_12776,N_12837);
and U19783 (N_19783,N_12813,N_10254);
nor U19784 (N_19784,N_12517,N_12943);
or U19785 (N_19785,N_11389,N_10789);
nor U19786 (N_19786,N_12290,N_12925);
nand U19787 (N_19787,N_12506,N_14494);
and U19788 (N_19788,N_14963,N_14708);
xor U19789 (N_19789,N_14477,N_10802);
or U19790 (N_19790,N_12446,N_10484);
and U19791 (N_19791,N_12517,N_10601);
nand U19792 (N_19792,N_10959,N_10567);
nand U19793 (N_19793,N_12090,N_11953);
xnor U19794 (N_19794,N_14729,N_13363);
nor U19795 (N_19795,N_11791,N_13243);
and U19796 (N_19796,N_13090,N_11948);
nand U19797 (N_19797,N_11754,N_13570);
nand U19798 (N_19798,N_12666,N_13893);
xnor U19799 (N_19799,N_11907,N_12111);
nand U19800 (N_19800,N_10207,N_10607);
nor U19801 (N_19801,N_11736,N_13281);
xor U19802 (N_19802,N_10664,N_11694);
nor U19803 (N_19803,N_14333,N_12928);
nor U19804 (N_19804,N_10512,N_12054);
and U19805 (N_19805,N_14834,N_12839);
or U19806 (N_19806,N_10231,N_13336);
nor U19807 (N_19807,N_10479,N_12696);
nand U19808 (N_19808,N_11115,N_14610);
nand U19809 (N_19809,N_14884,N_13608);
and U19810 (N_19810,N_11580,N_13595);
or U19811 (N_19811,N_13752,N_11412);
xor U19812 (N_19812,N_11313,N_14291);
nand U19813 (N_19813,N_11333,N_12862);
and U19814 (N_19814,N_12992,N_11043);
nand U19815 (N_19815,N_12305,N_14328);
nand U19816 (N_19816,N_13906,N_12733);
xor U19817 (N_19817,N_14220,N_12301);
xnor U19818 (N_19818,N_13807,N_13305);
and U19819 (N_19819,N_14630,N_12143);
xor U19820 (N_19820,N_14484,N_12265);
nor U19821 (N_19821,N_14644,N_10886);
nor U19822 (N_19822,N_10542,N_13917);
and U19823 (N_19823,N_14728,N_14290);
nand U19824 (N_19824,N_10294,N_10268);
nand U19825 (N_19825,N_14586,N_11802);
and U19826 (N_19826,N_12773,N_13990);
nor U19827 (N_19827,N_11696,N_11713);
and U19828 (N_19828,N_10864,N_11932);
xor U19829 (N_19829,N_14122,N_13231);
xnor U19830 (N_19830,N_12703,N_10301);
nand U19831 (N_19831,N_11563,N_14144);
xor U19832 (N_19832,N_12049,N_10602);
or U19833 (N_19833,N_11851,N_14287);
and U19834 (N_19834,N_14659,N_10957);
nor U19835 (N_19835,N_11013,N_11271);
and U19836 (N_19836,N_11053,N_14237);
or U19837 (N_19837,N_13902,N_14838);
nand U19838 (N_19838,N_10339,N_11927);
nand U19839 (N_19839,N_11560,N_10869);
or U19840 (N_19840,N_14687,N_14394);
nand U19841 (N_19841,N_14320,N_13022);
and U19842 (N_19842,N_14568,N_10625);
or U19843 (N_19843,N_12156,N_10201);
nor U19844 (N_19844,N_10776,N_13331);
or U19845 (N_19845,N_10629,N_14581);
xor U19846 (N_19846,N_11593,N_14443);
nor U19847 (N_19847,N_10381,N_13059);
nand U19848 (N_19848,N_12252,N_13138);
nor U19849 (N_19849,N_12336,N_13410);
nor U19850 (N_19850,N_10712,N_10476);
and U19851 (N_19851,N_13815,N_12034);
and U19852 (N_19852,N_12202,N_13973);
or U19853 (N_19853,N_12357,N_11707);
nand U19854 (N_19854,N_11833,N_11346);
nor U19855 (N_19855,N_13652,N_11898);
xor U19856 (N_19856,N_11894,N_12087);
xor U19857 (N_19857,N_10614,N_12436);
and U19858 (N_19858,N_13602,N_12463);
nor U19859 (N_19859,N_10592,N_12824);
nor U19860 (N_19860,N_12873,N_13591);
xor U19861 (N_19861,N_11779,N_11844);
and U19862 (N_19862,N_12710,N_13222);
and U19863 (N_19863,N_12850,N_11836);
xor U19864 (N_19864,N_13946,N_14282);
and U19865 (N_19865,N_11729,N_13285);
xor U19866 (N_19866,N_11143,N_12001);
nor U19867 (N_19867,N_10030,N_14971);
nor U19868 (N_19868,N_12536,N_10708);
nor U19869 (N_19869,N_11890,N_12171);
xnor U19870 (N_19870,N_13683,N_11296);
nand U19871 (N_19871,N_12396,N_10951);
and U19872 (N_19872,N_13361,N_10608);
nor U19873 (N_19873,N_14147,N_13671);
nor U19874 (N_19874,N_12404,N_13931);
and U19875 (N_19875,N_11273,N_11172);
nor U19876 (N_19876,N_11143,N_12386);
and U19877 (N_19877,N_14181,N_13215);
or U19878 (N_19878,N_14448,N_14836);
xor U19879 (N_19879,N_10011,N_13343);
nand U19880 (N_19880,N_12017,N_13782);
xnor U19881 (N_19881,N_10020,N_14329);
nand U19882 (N_19882,N_11392,N_14067);
nor U19883 (N_19883,N_14168,N_10895);
nand U19884 (N_19884,N_14391,N_13142);
nor U19885 (N_19885,N_11000,N_12584);
nor U19886 (N_19886,N_12047,N_14848);
xnor U19887 (N_19887,N_11854,N_12266);
and U19888 (N_19888,N_13213,N_13389);
nor U19889 (N_19889,N_11610,N_13352);
and U19890 (N_19890,N_13579,N_10839);
and U19891 (N_19891,N_10137,N_10355);
and U19892 (N_19892,N_11025,N_10854);
and U19893 (N_19893,N_10269,N_14663);
nand U19894 (N_19894,N_11740,N_13946);
xor U19895 (N_19895,N_11428,N_12101);
xnor U19896 (N_19896,N_12412,N_10024);
nor U19897 (N_19897,N_11347,N_14955);
and U19898 (N_19898,N_12758,N_13217);
or U19899 (N_19899,N_12760,N_10716);
nand U19900 (N_19900,N_12192,N_14027);
and U19901 (N_19901,N_11230,N_10904);
nand U19902 (N_19902,N_11762,N_13481);
nor U19903 (N_19903,N_11501,N_13990);
or U19904 (N_19904,N_14282,N_14443);
xnor U19905 (N_19905,N_13451,N_12055);
xnor U19906 (N_19906,N_11270,N_13645);
nor U19907 (N_19907,N_11925,N_11233);
and U19908 (N_19908,N_13470,N_11679);
and U19909 (N_19909,N_14338,N_11052);
nor U19910 (N_19910,N_10941,N_13478);
or U19911 (N_19911,N_10729,N_12179);
nand U19912 (N_19912,N_14970,N_13576);
nor U19913 (N_19913,N_12494,N_14385);
nor U19914 (N_19914,N_11907,N_11947);
nor U19915 (N_19915,N_11865,N_14704);
nand U19916 (N_19916,N_12063,N_13844);
and U19917 (N_19917,N_13403,N_10839);
nand U19918 (N_19918,N_11707,N_11291);
xor U19919 (N_19919,N_13475,N_10659);
nor U19920 (N_19920,N_11315,N_11942);
nor U19921 (N_19921,N_14568,N_10945);
nand U19922 (N_19922,N_13793,N_13323);
xor U19923 (N_19923,N_11094,N_10702);
nand U19924 (N_19924,N_14544,N_14416);
or U19925 (N_19925,N_11054,N_13208);
or U19926 (N_19926,N_14963,N_14224);
or U19927 (N_19927,N_14553,N_11914);
nand U19928 (N_19928,N_10255,N_13257);
xor U19929 (N_19929,N_10491,N_11965);
nor U19930 (N_19930,N_10985,N_10655);
xnor U19931 (N_19931,N_12234,N_10406);
and U19932 (N_19932,N_14067,N_12878);
and U19933 (N_19933,N_11487,N_10553);
nor U19934 (N_19934,N_14044,N_14897);
nor U19935 (N_19935,N_13852,N_11177);
and U19936 (N_19936,N_13719,N_10345);
nor U19937 (N_19937,N_13798,N_12045);
and U19938 (N_19938,N_13229,N_11413);
and U19939 (N_19939,N_10512,N_13258);
nand U19940 (N_19940,N_10442,N_11542);
nand U19941 (N_19941,N_14002,N_11489);
xnor U19942 (N_19942,N_10120,N_12969);
and U19943 (N_19943,N_11322,N_11829);
or U19944 (N_19944,N_14676,N_13798);
nand U19945 (N_19945,N_11496,N_10791);
nor U19946 (N_19946,N_13613,N_13483);
nand U19947 (N_19947,N_11059,N_14404);
nor U19948 (N_19948,N_11451,N_14467);
or U19949 (N_19949,N_10064,N_11015);
or U19950 (N_19950,N_12485,N_14622);
xor U19951 (N_19951,N_12415,N_13699);
and U19952 (N_19952,N_14324,N_13788);
xor U19953 (N_19953,N_14949,N_11473);
nand U19954 (N_19954,N_10318,N_10615);
nor U19955 (N_19955,N_13570,N_10575);
nor U19956 (N_19956,N_11656,N_13327);
or U19957 (N_19957,N_11103,N_13743);
nor U19958 (N_19958,N_10360,N_12088);
nand U19959 (N_19959,N_11730,N_13914);
xor U19960 (N_19960,N_11433,N_12342);
nor U19961 (N_19961,N_14040,N_12544);
and U19962 (N_19962,N_12970,N_10386);
xnor U19963 (N_19963,N_13465,N_10230);
nand U19964 (N_19964,N_12130,N_12870);
or U19965 (N_19965,N_12323,N_14729);
or U19966 (N_19966,N_11095,N_13280);
nor U19967 (N_19967,N_10739,N_11918);
or U19968 (N_19968,N_10413,N_10693);
nor U19969 (N_19969,N_12094,N_11230);
xnor U19970 (N_19970,N_14309,N_12617);
and U19971 (N_19971,N_14757,N_10102);
nand U19972 (N_19972,N_10572,N_14559);
nor U19973 (N_19973,N_13571,N_11536);
and U19974 (N_19974,N_13347,N_13936);
xor U19975 (N_19975,N_10439,N_11928);
or U19976 (N_19976,N_12316,N_14730);
xnor U19977 (N_19977,N_13301,N_10348);
nand U19978 (N_19978,N_11607,N_12455);
nand U19979 (N_19979,N_12586,N_14887);
xnor U19980 (N_19980,N_13017,N_13883);
or U19981 (N_19981,N_13726,N_13492);
nand U19982 (N_19982,N_11560,N_11112);
or U19983 (N_19983,N_14399,N_10163);
or U19984 (N_19984,N_13663,N_14493);
and U19985 (N_19985,N_14054,N_13895);
or U19986 (N_19986,N_10921,N_14547);
or U19987 (N_19987,N_13440,N_10404);
and U19988 (N_19988,N_11457,N_11586);
nor U19989 (N_19989,N_10883,N_14576);
xor U19990 (N_19990,N_13751,N_13254);
xnor U19991 (N_19991,N_14826,N_12865);
nor U19992 (N_19992,N_12125,N_12256);
nand U19993 (N_19993,N_14520,N_10391);
xnor U19994 (N_19994,N_13027,N_13983);
and U19995 (N_19995,N_12341,N_10180);
nor U19996 (N_19996,N_12680,N_11919);
xnor U19997 (N_19997,N_12686,N_11876);
xor U19998 (N_19998,N_13488,N_13718);
or U19999 (N_19999,N_12922,N_12122);
xnor U20000 (N_20000,N_15632,N_16709);
nor U20001 (N_20001,N_18615,N_15537);
nor U20002 (N_20002,N_19398,N_16794);
and U20003 (N_20003,N_16681,N_19750);
nor U20004 (N_20004,N_19678,N_19170);
and U20005 (N_20005,N_19448,N_17046);
nand U20006 (N_20006,N_18340,N_18589);
xor U20007 (N_20007,N_15225,N_16148);
or U20008 (N_20008,N_18606,N_17952);
xnor U20009 (N_20009,N_16616,N_15682);
nand U20010 (N_20010,N_16765,N_18778);
or U20011 (N_20011,N_19633,N_15931);
xor U20012 (N_20012,N_15589,N_18146);
xnor U20013 (N_20013,N_18953,N_16370);
nand U20014 (N_20014,N_15079,N_18038);
xor U20015 (N_20015,N_15509,N_18926);
nand U20016 (N_20016,N_18062,N_19708);
or U20017 (N_20017,N_18289,N_18434);
nor U20018 (N_20018,N_19126,N_16491);
and U20019 (N_20019,N_19489,N_17051);
and U20020 (N_20020,N_19308,N_16625);
xor U20021 (N_20021,N_16732,N_17944);
and U20022 (N_20022,N_18908,N_15268);
and U20023 (N_20023,N_16345,N_16246);
and U20024 (N_20024,N_16596,N_15446);
or U20025 (N_20025,N_19339,N_17583);
and U20026 (N_20026,N_19189,N_18624);
nor U20027 (N_20027,N_16831,N_18706);
nor U20028 (N_20028,N_18413,N_16319);
and U20029 (N_20029,N_19920,N_16744);
and U20030 (N_20030,N_17553,N_16091);
or U20031 (N_20031,N_15940,N_19981);
xor U20032 (N_20032,N_19233,N_15508);
and U20033 (N_20033,N_18870,N_16297);
xnor U20034 (N_20034,N_19322,N_16181);
nor U20035 (N_20035,N_15449,N_17276);
and U20036 (N_20036,N_18239,N_17642);
and U20037 (N_20037,N_19713,N_18861);
or U20038 (N_20038,N_17123,N_18035);
or U20039 (N_20039,N_16380,N_15377);
xor U20040 (N_20040,N_18659,N_16296);
xnor U20041 (N_20041,N_17181,N_18839);
and U20042 (N_20042,N_15310,N_16541);
nor U20043 (N_20043,N_19254,N_15739);
nand U20044 (N_20044,N_19897,N_18500);
or U20045 (N_20045,N_18002,N_15425);
and U20046 (N_20046,N_19621,N_18126);
xor U20047 (N_20047,N_16802,N_16511);
xor U20048 (N_20048,N_19315,N_17531);
nand U20049 (N_20049,N_19351,N_17846);
xnor U20050 (N_20050,N_19153,N_18172);
and U20051 (N_20051,N_18282,N_17066);
nand U20052 (N_20052,N_15922,N_19790);
and U20053 (N_20053,N_15021,N_18066);
or U20054 (N_20054,N_15878,N_17721);
xnor U20055 (N_20055,N_15477,N_18543);
nor U20056 (N_20056,N_19063,N_17275);
and U20057 (N_20057,N_15895,N_17355);
nor U20058 (N_20058,N_17119,N_15703);
nor U20059 (N_20059,N_16656,N_16562);
and U20060 (N_20060,N_15843,N_16067);
nor U20061 (N_20061,N_19843,N_16219);
nand U20062 (N_20062,N_18341,N_16904);
xnor U20063 (N_20063,N_18833,N_18810);
and U20064 (N_20064,N_17338,N_19648);
xor U20065 (N_20065,N_18705,N_19326);
or U20066 (N_20066,N_19813,N_16005);
nand U20067 (N_20067,N_15213,N_19471);
and U20068 (N_20068,N_18580,N_16305);
xnor U20069 (N_20069,N_17710,N_18812);
nand U20070 (N_20070,N_15686,N_16956);
or U20071 (N_20071,N_16875,N_17077);
or U20072 (N_20072,N_19327,N_19537);
nand U20073 (N_20073,N_17070,N_17759);
nand U20074 (N_20074,N_17218,N_15595);
nor U20075 (N_20075,N_15999,N_16584);
and U20076 (N_20076,N_18233,N_19477);
and U20077 (N_20077,N_15609,N_18387);
or U20078 (N_20078,N_18482,N_18645);
nor U20079 (N_20079,N_16789,N_17715);
or U20080 (N_20080,N_15665,N_19154);
nor U20081 (N_20081,N_19280,N_15381);
xor U20082 (N_20082,N_15012,N_17628);
nand U20083 (N_20083,N_18945,N_16226);
or U20084 (N_20084,N_15140,N_18583);
nand U20085 (N_20085,N_16530,N_19918);
nor U20086 (N_20086,N_17502,N_18797);
xnor U20087 (N_20087,N_16339,N_18018);
or U20088 (N_20088,N_18834,N_19038);
xor U20089 (N_20089,N_18904,N_16374);
and U20090 (N_20090,N_19355,N_17784);
nand U20091 (N_20091,N_19856,N_19418);
and U20092 (N_20092,N_17567,N_18318);
or U20093 (N_20093,N_18088,N_16605);
and U20094 (N_20094,N_18327,N_19396);
and U20095 (N_20095,N_15748,N_18127);
nor U20096 (N_20096,N_17454,N_19915);
xor U20097 (N_20097,N_19823,N_15771);
or U20098 (N_20098,N_15283,N_17742);
nor U20099 (N_20099,N_18489,N_17354);
xor U20100 (N_20100,N_19965,N_19048);
nor U20101 (N_20101,N_19746,N_16688);
or U20102 (N_20102,N_18649,N_15633);
or U20103 (N_20103,N_18915,N_19803);
nand U20104 (N_20104,N_16679,N_17898);
and U20105 (N_20105,N_17030,N_16347);
and U20106 (N_20106,N_16349,N_16400);
xnor U20107 (N_20107,N_19910,N_19580);
and U20108 (N_20108,N_19286,N_15976);
xnor U20109 (N_20109,N_15583,N_16902);
nand U20110 (N_20110,N_18895,N_18347);
xor U20111 (N_20111,N_19806,N_16220);
and U20112 (N_20112,N_17498,N_18253);
nand U20113 (N_20113,N_16918,N_19564);
and U20114 (N_20114,N_17970,N_15025);
nand U20115 (N_20115,N_16440,N_16986);
xor U20116 (N_20116,N_16798,N_17886);
nor U20117 (N_20117,N_16313,N_16730);
or U20118 (N_20118,N_16818,N_15904);
or U20119 (N_20119,N_18545,N_17778);
xnor U20120 (N_20120,N_17474,N_17258);
and U20121 (N_20121,N_17381,N_17505);
or U20122 (N_20122,N_16391,N_17932);
xor U20123 (N_20123,N_16830,N_16170);
nor U20124 (N_20124,N_18271,N_16809);
nor U20125 (N_20125,N_17521,N_15235);
nand U20126 (N_20126,N_17496,N_16773);
nor U20127 (N_20127,N_17373,N_18249);
or U20128 (N_20128,N_17653,N_18665);
nand U20129 (N_20129,N_17489,N_19523);
nand U20130 (N_20130,N_15276,N_16166);
or U20131 (N_20131,N_19963,N_17903);
or U20132 (N_20132,N_17314,N_17876);
xor U20133 (N_20133,N_18419,N_15844);
nand U20134 (N_20134,N_16238,N_15629);
xnor U20135 (N_20135,N_15037,N_15405);
or U20136 (N_20136,N_19776,N_18377);
nor U20137 (N_20137,N_17257,N_19367);
xnor U20138 (N_20138,N_15651,N_16423);
or U20139 (N_20139,N_15138,N_18941);
or U20140 (N_20140,N_19206,N_19120);
nor U20141 (N_20141,N_18558,N_19698);
nor U20142 (N_20142,N_18421,N_19866);
nor U20143 (N_20143,N_15286,N_17221);
and U20144 (N_20144,N_17093,N_17029);
nor U20145 (N_20145,N_16072,N_18905);
and U20146 (N_20146,N_17767,N_19936);
and U20147 (N_20147,N_18855,N_19954);
or U20148 (N_20148,N_17666,N_16415);
nor U20149 (N_20149,N_19437,N_18345);
or U20150 (N_20150,N_18224,N_17271);
nor U20151 (N_20151,N_15220,N_16320);
nand U20152 (N_20152,N_16650,N_19852);
and U20153 (N_20153,N_16668,N_15707);
xnor U20154 (N_20154,N_15673,N_17821);
xor U20155 (N_20155,N_19131,N_18256);
nor U20156 (N_20156,N_16707,N_18399);
or U20157 (N_20157,N_19271,N_16954);
nor U20158 (N_20158,N_15496,N_17985);
or U20159 (N_20159,N_16567,N_19588);
and U20160 (N_20160,N_17801,N_19508);
nand U20161 (N_20161,N_17728,N_17228);
and U20162 (N_20162,N_17601,N_15476);
nand U20163 (N_20163,N_19744,N_18620);
and U20164 (N_20164,N_15628,N_19433);
nor U20165 (N_20165,N_15302,N_16648);
nor U20166 (N_20166,N_15863,N_15663);
nand U20167 (N_20167,N_17399,N_15608);
or U20168 (N_20168,N_18053,N_18889);
or U20169 (N_20169,N_18965,N_18028);
nand U20170 (N_20170,N_19660,N_16204);
nor U20171 (N_20171,N_15824,N_15702);
nand U20172 (N_20172,N_18844,N_16436);
xnor U20173 (N_20173,N_18228,N_17648);
or U20174 (N_20174,N_16350,N_18843);
xnor U20175 (N_20175,N_19578,N_16791);
nand U20176 (N_20176,N_16711,N_17220);
or U20177 (N_20177,N_19362,N_19811);
nor U20178 (N_20178,N_17855,N_19664);
and U20179 (N_20179,N_17617,N_15781);
or U20180 (N_20180,N_18221,N_15104);
xor U20181 (N_20181,N_15888,N_15561);
nand U20182 (N_20182,N_19608,N_15164);
nor U20183 (N_20183,N_15577,N_17036);
nand U20184 (N_20184,N_15601,N_15814);
or U20185 (N_20185,N_19090,N_16360);
xor U20186 (N_20186,N_19095,N_18990);
xor U20187 (N_20187,N_18913,N_18763);
and U20188 (N_20188,N_16402,N_15669);
or U20189 (N_20189,N_15184,N_17391);
and U20190 (N_20190,N_15144,N_17164);
nand U20191 (N_20191,N_15203,N_15614);
nand U20192 (N_20192,N_16674,N_15178);
xor U20193 (N_20193,N_17991,N_18007);
and U20194 (N_20194,N_15334,N_16050);
and U20195 (N_20195,N_17914,N_15499);
nand U20196 (N_20196,N_17610,N_15558);
nand U20197 (N_20197,N_17114,N_15581);
and U20198 (N_20198,N_17349,N_17321);
or U20199 (N_20199,N_19614,N_18217);
nand U20200 (N_20200,N_19949,N_16086);
or U20201 (N_20201,N_18086,N_18732);
xor U20202 (N_20202,N_16793,N_16076);
or U20203 (N_20203,N_17544,N_19465);
nor U20204 (N_20204,N_18806,N_15366);
nand U20205 (N_20205,N_19876,N_17834);
and U20206 (N_20206,N_19613,N_18792);
or U20207 (N_20207,N_18004,N_15038);
nand U20208 (N_20208,N_17313,N_17635);
and U20209 (N_20209,N_18588,N_19216);
or U20210 (N_20210,N_18911,N_18738);
xor U20211 (N_20211,N_16309,N_15852);
and U20212 (N_20212,N_17669,N_19479);
xnor U20213 (N_20213,N_18368,N_18962);
nor U20214 (N_20214,N_15638,N_18655);
xor U20215 (N_20215,N_19328,N_18757);
and U20216 (N_20216,N_19911,N_15088);
nor U20217 (N_20217,N_18747,N_18090);
xnor U20218 (N_20218,N_18788,N_16102);
and U20219 (N_20219,N_17796,N_17266);
nor U20220 (N_20220,N_18200,N_19719);
and U20221 (N_20221,N_16083,N_16623);
xnor U20222 (N_20222,N_19478,N_17472);
or U20223 (N_20223,N_17217,N_15625);
and U20224 (N_20224,N_18385,N_17014);
nor U20225 (N_20225,N_19199,N_15403);
nor U20226 (N_20226,N_16587,N_16554);
xnor U20227 (N_20227,N_19848,N_19446);
nand U20228 (N_20228,N_19023,N_16641);
nand U20229 (N_20229,N_18652,N_18560);
nand U20230 (N_20230,N_16643,N_15556);
or U20231 (N_20231,N_17296,N_16367);
nand U20232 (N_20232,N_16578,N_17219);
nor U20233 (N_20233,N_15237,N_19006);
or U20234 (N_20234,N_16630,N_15315);
and U20235 (N_20235,N_18454,N_15946);
xnor U20236 (N_20236,N_18938,N_19325);
or U20237 (N_20237,N_18107,N_16343);
nor U20238 (N_20238,N_17435,N_17329);
xor U20239 (N_20239,N_18559,N_19042);
nand U20240 (N_20240,N_16093,N_18106);
nor U20241 (N_20241,N_18847,N_16441);
xnor U20242 (N_20242,N_18582,N_19575);
and U20243 (N_20243,N_17862,N_17517);
or U20244 (N_20244,N_15872,N_18936);
nor U20245 (N_20245,N_18414,N_15085);
and U20246 (N_20246,N_19935,N_15547);
nand U20247 (N_20247,N_16131,N_18484);
xor U20248 (N_20248,N_18912,N_17394);
nor U20249 (N_20249,N_19764,N_16368);
xnor U20250 (N_20250,N_19293,N_17144);
or U20251 (N_20251,N_16920,N_16257);
or U20252 (N_20252,N_19344,N_19980);
nor U20253 (N_20253,N_18978,N_15480);
nor U20254 (N_20254,N_19188,N_17245);
and U20255 (N_20255,N_18651,N_15098);
nand U20256 (N_20256,N_17363,N_17009);
or U20257 (N_20257,N_17649,N_17259);
and U20258 (N_20258,N_18835,N_18262);
nor U20259 (N_20259,N_18346,N_19198);
nor U20260 (N_20260,N_15465,N_17148);
nand U20261 (N_20261,N_18917,N_18805);
and U20262 (N_20262,N_17773,N_15199);
and U20263 (N_20263,N_18487,N_17339);
and U20264 (N_20264,N_17833,N_17933);
xnor U20265 (N_20265,N_18301,N_17169);
nor U20266 (N_20266,N_19807,N_15969);
nand U20267 (N_20267,N_19461,N_16949);
xnor U20268 (N_20268,N_15386,N_16048);
and U20269 (N_20269,N_15524,N_16375);
or U20270 (N_20270,N_15357,N_17269);
or U20271 (N_20271,N_15110,N_18512);
and U20272 (N_20272,N_16827,N_18435);
or U20273 (N_20273,N_18240,N_19140);
nor U20274 (N_20274,N_15719,N_19606);
nor U20275 (N_20275,N_19145,N_16645);
or U20276 (N_20276,N_18058,N_15009);
nor U20277 (N_20277,N_15239,N_15950);
or U20278 (N_20278,N_16095,N_18140);
or U20279 (N_20279,N_18077,N_18252);
nor U20280 (N_20280,N_19817,N_18799);
xnor U20281 (N_20281,N_15807,N_17350);
and U20282 (N_20282,N_16342,N_18231);
nor U20283 (N_20283,N_17462,N_16116);
nor U20284 (N_20284,N_19135,N_18569);
nor U20285 (N_20285,N_17265,N_16774);
nand U20286 (N_20286,N_18669,N_17019);
nor U20287 (N_20287,N_16951,N_18299);
and U20288 (N_20288,N_17912,N_15860);
nand U20289 (N_20289,N_17015,N_15964);
xor U20290 (N_20290,N_19905,N_16034);
nand U20291 (N_20291,N_18476,N_17662);
and U20292 (N_20292,N_17809,N_15920);
and U20293 (N_20293,N_18247,N_18483);
and U20294 (N_20294,N_19840,N_19321);
or U20295 (N_20295,N_18991,N_16447);
nor U20296 (N_20296,N_15913,N_16610);
nor U20297 (N_20297,N_19600,N_16200);
nand U20298 (N_20298,N_16886,N_19672);
or U20299 (N_20299,N_16040,N_16944);
nor U20300 (N_20300,N_18376,N_17779);
and U20301 (N_20301,N_15658,N_17063);
nand U20302 (N_20302,N_19710,N_17331);
xnor U20303 (N_20303,N_18869,N_17356);
nor U20304 (N_20304,N_15684,N_16743);
and U20305 (N_20305,N_19889,N_15796);
or U20306 (N_20306,N_18822,N_18405);
or U20307 (N_20307,N_17510,N_17684);
or U20308 (N_20308,N_15389,N_16130);
nor U20309 (N_20309,N_16253,N_15296);
xor U20310 (N_20310,N_15903,N_16272);
xor U20311 (N_20311,N_17732,N_16387);
nor U20312 (N_20312,N_17301,N_19881);
nand U20313 (N_20313,N_18470,N_19970);
and U20314 (N_20314,N_19128,N_16202);
xor U20315 (N_20315,N_19707,N_18122);
xnor U20316 (N_20316,N_16509,N_15955);
nor U20317 (N_20317,N_18308,N_19679);
nor U20318 (N_20318,N_16290,N_17017);
or U20319 (N_20319,N_17386,N_17040);
nand U20320 (N_20320,N_19360,N_15906);
nand U20321 (N_20321,N_16221,N_18030);
or U20322 (N_20322,N_15122,N_15223);
and U20323 (N_20323,N_19788,N_17982);
nor U20324 (N_20324,N_16482,N_16576);
nor U20325 (N_20325,N_17334,N_15986);
and U20326 (N_20326,N_18670,N_16751);
or U20327 (N_20327,N_17436,N_16039);
or U20328 (N_20328,N_16619,N_16042);
nand U20329 (N_20329,N_19838,N_15972);
or U20330 (N_20330,N_15031,N_19000);
and U20331 (N_20331,N_19507,N_17103);
nor U20332 (N_20332,N_16861,N_16850);
nor U20333 (N_20333,N_19442,N_19323);
and U20334 (N_20334,N_17121,N_16722);
nand U20335 (N_20335,N_15907,N_17563);
or U20336 (N_20336,N_15637,N_16031);
and U20337 (N_20337,N_15507,N_18397);
and U20338 (N_20338,N_17958,N_16685);
or U20339 (N_20339,N_15434,N_15528);
or U20340 (N_20340,N_16718,N_15724);
nor U20341 (N_20341,N_19445,N_19278);
xor U20342 (N_20342,N_17926,N_17290);
or U20343 (N_20343,N_17761,N_16432);
nand U20344 (N_20344,N_19341,N_16999);
nand U20345 (N_20345,N_16810,N_18339);
nor U20346 (N_20346,N_19775,N_17882);
and U20347 (N_20347,N_15754,N_16026);
xor U20348 (N_20348,N_18828,N_17626);
nand U20349 (N_20349,N_15497,N_16869);
or U20350 (N_20350,N_16377,N_16540);
or U20351 (N_20351,N_17828,N_18618);
xnor U20352 (N_20352,N_15960,N_19676);
nor U20353 (N_20353,N_15160,N_15887);
xnor U20354 (N_20354,N_18444,N_15078);
xnor U20355 (N_20355,N_19671,N_16165);
and U20356 (N_20356,N_15185,N_19574);
nor U20357 (N_20357,N_18459,N_15475);
or U20358 (N_20358,N_19825,N_19598);
nand U20359 (N_20359,N_17600,N_18691);
and U20360 (N_20360,N_18048,N_16976);
xor U20361 (N_20361,N_17414,N_19332);
nand U20362 (N_20362,N_18390,N_16728);
nand U20363 (N_20363,N_16962,N_17061);
or U20364 (N_20364,N_18450,N_15287);
nor U20365 (N_20365,N_17021,N_18143);
nor U20366 (N_20366,N_16358,N_19755);
nand U20367 (N_20367,N_16479,N_19522);
xnor U20368 (N_20368,N_17083,N_16465);
and U20369 (N_20369,N_19833,N_19570);
and U20370 (N_20370,N_15414,N_17942);
xnor U20371 (N_20371,N_17272,N_19995);
or U20372 (N_20372,N_16586,N_18125);
nor U20373 (N_20373,N_17412,N_18370);
nor U20374 (N_20374,N_17254,N_18621);
nand U20375 (N_20375,N_19822,N_15322);
and U20376 (N_20376,N_19392,N_18374);
and U20377 (N_20377,N_15693,N_18207);
and U20378 (N_20378,N_19432,N_16526);
nand U20379 (N_20379,N_16153,N_16662);
or U20380 (N_20380,N_19155,N_15847);
and U20381 (N_20381,N_18523,N_15309);
nor U20382 (N_20382,N_17528,N_17174);
and U20383 (N_20383,N_16263,N_19407);
nand U20384 (N_20384,N_15522,N_18557);
xor U20385 (N_20385,N_17185,N_17509);
or U20386 (N_20386,N_19898,N_15933);
and U20387 (N_20387,N_16515,N_16485);
xnor U20388 (N_20388,N_19184,N_15065);
or U20389 (N_20389,N_16860,N_16770);
and U20390 (N_20390,N_17380,N_15156);
nand U20391 (N_20391,N_17611,N_18296);
nand U20392 (N_20392,N_18758,N_17532);
xnor U20393 (N_20393,N_17387,N_18392);
and U20394 (N_20394,N_15474,N_15026);
nor U20395 (N_20395,N_15194,N_17237);
xnor U20396 (N_20396,N_19704,N_18456);
nor U20397 (N_20397,N_16488,N_17561);
or U20398 (N_20398,N_15889,N_16232);
nor U20399 (N_20399,N_19429,N_19193);
xnor U20400 (N_20400,N_19076,N_19207);
or U20401 (N_20401,N_16628,N_18883);
nand U20402 (N_20402,N_19747,N_19521);
or U20403 (N_20403,N_18932,N_19997);
xor U20404 (N_20404,N_15606,N_18786);
nor U20405 (N_20405,N_16484,N_16085);
xor U20406 (N_20406,N_18598,N_17018);
or U20407 (N_20407,N_15846,N_16973);
and U20408 (N_20408,N_16336,N_16283);
nor U20409 (N_20409,N_17515,N_17848);
nand U20410 (N_20410,N_19110,N_16328);
or U20411 (N_20411,N_19659,N_15421);
nor U20412 (N_20412,N_18553,N_17470);
and U20413 (N_20413,N_16492,N_15788);
nand U20414 (N_20414,N_16348,N_17364);
nand U20415 (N_20415,N_16197,N_15206);
nor U20416 (N_20416,N_15699,N_16982);
or U20417 (N_20417,N_19637,N_17790);
nand U20418 (N_20418,N_15598,N_16560);
nor U20419 (N_20419,N_18098,N_16943);
xnor U20420 (N_20420,N_18765,N_19349);
or U20421 (N_20421,N_16241,N_17538);
nand U20422 (N_20422,N_17636,N_17191);
nor U20423 (N_20423,N_16803,N_17889);
xnor U20424 (N_20424,N_16813,N_15112);
xor U20425 (N_20425,N_15909,N_15033);
and U20426 (N_20426,N_16405,N_18698);
nor U20427 (N_20427,N_19005,N_19594);
and U20428 (N_20428,N_16428,N_15557);
and U20429 (N_20429,N_16457,N_17695);
xor U20430 (N_20430,N_15265,N_18635);
nand U20431 (N_20431,N_18718,N_18064);
nor U20432 (N_20432,N_17755,N_18804);
xnor U20433 (N_20433,N_17211,N_16775);
xnor U20434 (N_20434,N_19767,N_18174);
nand U20435 (N_20435,N_16110,N_18964);
nand U20436 (N_20436,N_16250,N_17554);
or U20437 (N_20437,N_18488,N_19491);
nor U20438 (N_20438,N_18429,N_16989);
and U20439 (N_20439,N_17333,N_18037);
or U20440 (N_20440,N_16425,N_19087);
and U20441 (N_20441,N_15813,N_16010);
or U20442 (N_20442,N_17465,N_19861);
and U20443 (N_20443,N_18350,N_18235);
nor U20444 (N_20444,N_18416,N_18856);
nand U20445 (N_20445,N_15457,N_19681);
and U20446 (N_20446,N_16388,N_19015);
and U20447 (N_20447,N_16068,N_18216);
and U20448 (N_20448,N_15181,N_16088);
nand U20449 (N_20449,N_16114,N_18182);
and U20450 (N_20450,N_17894,N_18739);
xor U20451 (N_20451,N_19809,N_15828);
or U20452 (N_20452,N_17581,N_15498);
nor U20453 (N_20453,N_19439,N_16318);
or U20454 (N_20454,N_16672,N_17162);
nand U20455 (N_20455,N_16849,N_19894);
nor U20456 (N_20456,N_18531,N_16742);
or U20457 (N_20457,N_18940,N_15858);
nand U20458 (N_20458,N_15299,N_15029);
nor U20459 (N_20459,N_17327,N_16359);
nand U20460 (N_20460,N_19099,N_16703);
nand U20461 (N_20461,N_17859,N_17922);
nor U20462 (N_20462,N_19195,N_17943);
nand U20463 (N_20463,N_16559,N_16483);
nor U20464 (N_20464,N_16779,N_15196);
or U20465 (N_20465,N_16639,N_18285);
and U20466 (N_20466,N_15354,N_16531);
nand U20467 (N_20467,N_16527,N_17607);
xnor U20468 (N_20468,N_16105,N_18496);
or U20469 (N_20469,N_18295,N_19631);
and U20470 (N_20470,N_18178,N_16287);
xnor U20471 (N_20471,N_15330,N_16523);
or U20472 (N_20472,N_17246,N_19912);
and U20473 (N_20473,N_18193,N_15382);
xor U20474 (N_20474,N_17129,N_18430);
nor U20475 (N_20475,N_18284,N_18731);
and U20476 (N_20476,N_18830,N_16061);
xor U20477 (N_20477,N_16876,N_17945);
or U20478 (N_20478,N_17749,N_17788);
and U20479 (N_20479,N_18266,N_19831);
xor U20480 (N_20480,N_15761,N_18012);
nand U20481 (N_20481,N_16780,N_17974);
xnor U20482 (N_20482,N_19228,N_16635);
nand U20483 (N_20483,N_17667,N_16315);
or U20484 (N_20484,N_15444,N_18097);
or U20485 (N_20485,N_18727,N_16642);
nand U20486 (N_20486,N_17145,N_18762);
or U20487 (N_20487,N_17622,N_16490);
xnor U20488 (N_20488,N_19238,N_19307);
nor U20489 (N_20489,N_19390,N_17307);
nand U20490 (N_20490,N_16256,N_16424);
or U20491 (N_20491,N_17540,N_16749);
or U20492 (N_20492,N_16341,N_17722);
nand U20493 (N_20493,N_17877,N_19690);
xnor U20494 (N_20494,N_18729,N_16948);
nand U20495 (N_20495,N_16379,N_15704);
nand U20496 (N_20496,N_17905,N_18309);
nand U20497 (N_20497,N_17996,N_18068);
and U20498 (N_20498,N_16450,N_15427);
nor U20499 (N_20499,N_19040,N_18780);
xnor U20500 (N_20500,N_19868,N_18261);
nor U20501 (N_20501,N_18115,N_19799);
nand U20502 (N_20502,N_19640,N_19143);
nand U20503 (N_20503,N_18020,N_16208);
xor U20504 (N_20504,N_15631,N_17948);
and U20505 (N_20505,N_15770,N_17957);
nor U20506 (N_20506,N_16146,N_19159);
or U20507 (N_20507,N_17207,N_15097);
xnor U20508 (N_20508,N_18579,N_19655);
or U20509 (N_20509,N_18794,N_15179);
nand U20510 (N_20510,N_18505,N_18796);
nand U20511 (N_20511,N_17423,N_17753);
or U20512 (N_20512,N_16461,N_19787);
xnor U20513 (N_20513,N_19180,N_17810);
or U20514 (N_20514,N_15851,N_15827);
xor U20515 (N_20515,N_17183,N_16453);
and U20516 (N_20516,N_18208,N_18867);
nor U20517 (N_20517,N_16829,N_17639);
and U20518 (N_20518,N_17647,N_16198);
nor U20519 (N_20519,N_19104,N_17078);
and U20520 (N_20520,N_19256,N_16442);
and U20521 (N_20521,N_15169,N_19568);
or U20522 (N_20522,N_17418,N_17464);
nor U20523 (N_20523,N_16437,N_15512);
nand U20524 (N_20524,N_16251,N_19619);
and U20525 (N_20525,N_18333,N_18680);
nand U20526 (N_20526,N_17797,N_17085);
and U20527 (N_20527,N_16781,N_15981);
nand U20528 (N_20528,N_18710,N_17816);
nand U20529 (N_20529,N_18540,N_17518);
nand U20530 (N_20530,N_15068,N_16323);
xor U20531 (N_20531,N_17137,N_15494);
and U20532 (N_20532,N_16723,N_16476);
and U20533 (N_20533,N_19529,N_19654);
nand U20534 (N_20534,N_15672,N_19039);
or U20535 (N_20535,N_18325,N_18594);
or U20536 (N_20536,N_18360,N_15411);
nor U20537 (N_20537,N_18473,N_16879);
or U20538 (N_20538,N_15942,N_16938);
and U20539 (N_20539,N_15572,N_19409);
nor U20540 (N_20540,N_19336,N_15221);
nor U20541 (N_20541,N_15753,N_17672);
or U20542 (N_20542,N_19701,N_15594);
nand U20543 (N_20543,N_16945,N_18597);
nand U20544 (N_20544,N_17201,N_16613);
and U20545 (N_20545,N_15681,N_16868);
or U20546 (N_20546,N_18250,N_16937);
xor U20547 (N_20547,N_18236,N_15540);
nor U20548 (N_20548,N_18417,N_16733);
nand U20549 (N_20549,N_17150,N_16249);
xnor U20550 (N_20550,N_17865,N_19171);
nor U20551 (N_20551,N_15586,N_16652);
xor U20552 (N_20552,N_17965,N_15792);
and U20553 (N_20553,N_17693,N_15648);
and U20554 (N_20554,N_16929,N_18059);
nand U20555 (N_20555,N_18303,N_18190);
or U20556 (N_20556,N_16503,N_19132);
nor U20557 (N_20557,N_18882,N_16247);
xnor U20558 (N_20558,N_18631,N_19275);
or U20559 (N_20559,N_19372,N_18836);
xor U20560 (N_20560,N_18436,N_19319);
xor U20561 (N_20561,N_15013,N_16536);
nand U20562 (N_20562,N_17564,N_18168);
and U20563 (N_20563,N_15319,N_17817);
and U20564 (N_20564,N_19998,N_19075);
nor U20565 (N_20565,N_18845,N_17155);
nand U20566 (N_20566,N_15740,N_16907);
nand U20567 (N_20567,N_16702,N_17482);
nand U20568 (N_20568,N_19045,N_15766);
nor U20569 (N_20569,N_19052,N_17978);
xor U20570 (N_20570,N_19169,N_15339);
xnor U20571 (N_20571,N_19078,N_15035);
xnor U20572 (N_20572,N_15915,N_15615);
xnor U20573 (N_20573,N_17654,N_17997);
xor U20574 (N_20574,N_18201,N_19636);
and U20575 (N_20575,N_16079,N_19643);
or U20576 (N_20576,N_16990,N_19844);
nand U20577 (N_20577,N_19097,N_17478);
and U20578 (N_20578,N_19089,N_19878);
or U20579 (N_20579,N_16027,N_18664);
and U20580 (N_20580,N_18492,N_17632);
nor U20581 (N_20581,N_18603,N_17800);
nand U20582 (N_20582,N_19794,N_15874);
nand U20583 (N_20583,N_15613,N_17508);
and U20584 (N_20584,N_16155,N_17455);
and U20585 (N_20585,N_17747,N_18149);
xnor U20586 (N_20586,N_18943,N_17971);
nand U20587 (N_20587,N_18326,N_19452);
or U20588 (N_20588,N_17253,N_17679);
or U20589 (N_20589,N_18952,N_15391);
xor U20590 (N_20590,N_19670,N_17921);
nor U20591 (N_20591,N_16163,N_16021);
nor U20592 (N_20592,N_17336,N_15782);
xor U20593 (N_20593,N_18114,N_16444);
and U20594 (N_20594,N_18394,N_18966);
and U20595 (N_20595,N_18842,N_19134);
and U20596 (N_20596,N_18191,N_15621);
and U20597 (N_20597,N_15373,N_17694);
and U20598 (N_20598,N_16382,N_17681);
xor U20599 (N_20599,N_16538,N_18342);
and U20600 (N_20600,N_16699,N_19234);
xor U20601 (N_20601,N_18666,N_15757);
or U20602 (N_20602,N_17707,N_18396);
or U20603 (N_20603,N_18752,N_16329);
or U20604 (N_20604,N_15859,N_17775);
xnor U20605 (N_20605,N_16960,N_17383);
xnor U20606 (N_20606,N_17726,N_17741);
or U20607 (N_20607,N_19211,N_19692);
nor U20608 (N_20608,N_18654,N_16636);
nand U20609 (N_20609,N_15831,N_15876);
and U20610 (N_20610,N_17153,N_16271);
nand U20611 (N_20611,N_17372,N_19172);
or U20612 (N_20612,N_17634,N_18442);
or U20613 (N_20613,N_15376,N_15061);
or U20614 (N_20614,N_15819,N_19547);
nor U20615 (N_20615,N_17122,N_17225);
xnor U20616 (N_20616,N_16126,N_18741);
nor U20617 (N_20617,N_19700,N_19149);
or U20618 (N_20618,N_19284,N_16456);
nand U20619 (N_20619,N_15820,N_17442);
and U20620 (N_20620,N_18682,N_17916);
nor U20621 (N_20621,N_19842,N_19950);
nor U20622 (N_20622,N_19812,N_19514);
and U20623 (N_20623,N_15855,N_15593);
xnor U20624 (N_20624,N_18837,N_16236);
nand U20625 (N_20625,N_15324,N_17449);
nand U20626 (N_20626,N_17294,N_16658);
nor U20627 (N_20627,N_17353,N_18985);
and U20628 (N_20628,N_16510,N_15800);
nor U20629 (N_20629,N_15550,N_16577);
or U20630 (N_20630,N_18721,N_15186);
nor U20631 (N_20631,N_16690,N_17194);
nand U20632 (N_20632,N_15886,N_16915);
nor U20633 (N_20633,N_16724,N_15838);
nor U20634 (N_20634,N_17319,N_18320);
nor U20635 (N_20635,N_17309,N_16946);
or U20636 (N_20636,N_15930,N_15086);
xor U20637 (N_20637,N_16245,N_18013);
and U20638 (N_20638,N_19603,N_17738);
or U20639 (N_20639,N_15742,N_17227);
and U20640 (N_20640,N_18081,N_19955);
nor U20641 (N_20641,N_18798,N_19836);
nor U20642 (N_20642,N_15227,N_19506);
and U20643 (N_20643,N_19236,N_16255);
xor U20644 (N_20644,N_16609,N_16138);
xor U20645 (N_20645,N_17831,N_16549);
or U20646 (N_20646,N_17766,N_18614);
or U20647 (N_20647,N_17637,N_19966);
xor U20648 (N_20648,N_15934,N_18637);
nor U20649 (N_20649,N_18948,N_19988);
xnor U20650 (N_20650,N_17757,N_15388);
and U20651 (N_20651,N_19541,N_19309);
xnor U20652 (N_20652,N_19960,N_17335);
nand U20653 (N_20653,N_18298,N_18006);
xnor U20654 (N_20654,N_19368,N_19532);
or U20655 (N_20655,N_17913,N_19653);
nor U20656 (N_20656,N_19779,N_18034);
or U20657 (N_20657,N_15114,N_18046);
and U20658 (N_20658,N_15230,N_18000);
nor U20659 (N_20659,N_18584,N_16115);
xnor U20660 (N_20660,N_17870,N_19953);
or U20661 (N_20661,N_17404,N_15849);
xnor U20662 (N_20662,N_18970,N_16664);
and U20663 (N_20663,N_17573,N_15527);
and U20664 (N_20664,N_18117,N_17798);
or U20665 (N_20665,N_15470,N_16118);
or U20666 (N_20666,N_19819,N_16135);
nor U20667 (N_20667,N_18744,N_19650);
and U20668 (N_20668,N_16772,N_17663);
and U20669 (N_20669,N_16820,N_17032);
nor U20670 (N_20670,N_16841,N_16404);
or U20671 (N_20671,N_15728,N_16545);
nor U20672 (N_20672,N_15036,N_19517);
nor U20673 (N_20673,N_17752,N_19573);
or U20674 (N_20674,N_19101,N_17097);
nand U20675 (N_20675,N_16859,N_15927);
or U20676 (N_20676,N_17420,N_18619);
nand U20677 (N_20677,N_15549,N_18009);
and U20678 (N_20678,N_19330,N_17107);
xor U20679 (N_20679,N_16867,N_17138);
and U20680 (N_20680,N_18375,N_16332);
and U20681 (N_20681,N_15304,N_17631);
or U20682 (N_20682,N_18029,N_19926);
or U20683 (N_20683,N_18657,N_16337);
xor U20684 (N_20684,N_17534,N_16771);
or U20685 (N_20685,N_18297,N_15344);
or U20686 (N_20686,N_19387,N_16007);
xnor U20687 (N_20687,N_15706,N_18042);
and U20688 (N_20688,N_16495,N_15243);
xor U20689 (N_20689,N_16008,N_19577);
or U20690 (N_20690,N_16838,N_18388);
nand U20691 (N_20691,N_16932,N_17342);
and U20692 (N_20692,N_18973,N_17365);
xnor U20693 (N_20693,N_17249,N_16002);
or U20694 (N_20694,N_17007,N_18858);
nand U20695 (N_20695,N_19020,N_17836);
xnor U20696 (N_20696,N_18975,N_16203);
nand U20697 (N_20697,N_17909,N_16970);
nor U20698 (N_20698,N_18113,N_15147);
nor U20699 (N_20699,N_19657,N_16967);
and U20700 (N_20700,N_18181,N_17823);
nor U20701 (N_20701,N_15242,N_18723);
xor U20702 (N_20702,N_19941,N_18923);
nor U20703 (N_20703,N_19074,N_19420);
or U20704 (N_20704,N_15610,N_16143);
and U20705 (N_20705,N_19302,N_16211);
nand U20706 (N_20706,N_17463,N_18186);
and U20707 (N_20707,N_15195,N_17044);
nor U20708 (N_20708,N_16726,N_16145);
nor U20709 (N_20709,N_15316,N_18141);
xor U20710 (N_20710,N_15074,N_19250);
xor U20711 (N_20711,N_16745,N_18872);
and U20712 (N_20712,N_16043,N_18503);
or U20713 (N_20713,N_18363,N_16410);
nor U20714 (N_20714,N_19869,N_15275);
or U20715 (N_20715,N_19994,N_19549);
and U20716 (N_20716,N_19406,N_18769);
nor U20717 (N_20717,N_19595,N_18897);
xor U20718 (N_20718,N_18535,N_19638);
xnor U20719 (N_20719,N_19977,N_17937);
or U20720 (N_20720,N_19921,N_16262);
and U20721 (N_20721,N_15562,N_15918);
xor U20722 (N_20722,N_18715,N_16659);
or U20723 (N_20723,N_18518,N_18969);
nand U20724 (N_20724,N_15717,N_18562);
nor U20725 (N_20725,N_18021,N_16899);
xnor U20726 (N_20726,N_17366,N_19828);
nand U20727 (N_20727,N_15552,N_18565);
and U20728 (N_20728,N_18108,N_17664);
and U20729 (N_20729,N_18587,N_16958);
xor U20730 (N_20730,N_18552,N_15829);
nor U20731 (N_20731,N_19300,N_17530);
and U20732 (N_20732,N_19297,N_18623);
xnor U20733 (N_20733,N_15129,N_15657);
nor U20734 (N_20734,N_15236,N_18093);
xor U20735 (N_20735,N_19417,N_17557);
xor U20736 (N_20736,N_17128,N_16267);
nand U20737 (N_20737,N_17452,N_15866);
nand U20738 (N_20738,N_15518,N_17720);
or U20739 (N_20739,N_18676,N_17703);
and U20740 (N_20740,N_15202,N_16366);
or U20741 (N_20741,N_19683,N_17956);
and U20742 (N_20742,N_19551,N_18424);
nor U20743 (N_20743,N_19901,N_18490);
nor U20744 (N_20744,N_19348,N_19394);
xor U20745 (N_20745,N_17106,N_16851);
xnor U20746 (N_20746,N_19624,N_15865);
xor U20747 (N_20747,N_17906,N_18819);
nor U20748 (N_20748,N_18022,N_15124);
and U20749 (N_20749,N_17130,N_15102);
or U20750 (N_20750,N_16910,N_16666);
nand U20751 (N_20751,N_17511,N_15359);
or U20752 (N_20752,N_19985,N_19524);
or U20753 (N_20753,N_19246,N_19401);
or U20754 (N_20754,N_19203,N_16224);
nand U20755 (N_20755,N_19179,N_18668);
xnor U20756 (N_20756,N_19780,N_17579);
and U20757 (N_20757,N_19352,N_15209);
and U20758 (N_20758,N_17892,N_16354);
nor U20759 (N_20759,N_18199,N_17547);
nand U20760 (N_20760,N_16569,N_19770);
and U20761 (N_20761,N_16448,N_16676);
or U20762 (N_20762,N_17791,N_19556);
nand U20763 (N_20763,N_17160,N_18566);
or U20764 (N_20764,N_19877,N_17764);
and U20765 (N_20765,N_19093,N_18329);
nand U20766 (N_20766,N_16637,N_19051);
xor U20767 (N_20767,N_18486,N_18644);
or U20768 (N_20768,N_16183,N_16980);
nand U20769 (N_20769,N_16878,N_15240);
xor U20770 (N_20770,N_19992,N_17367);
nand U20771 (N_20771,N_16385,N_19884);
nand U20772 (N_20772,N_15952,N_19397);
and U20773 (N_20773,N_18403,N_19258);
xnor U20774 (N_20774,N_16696,N_16431);
nand U20775 (N_20775,N_17481,N_15718);
nor U20776 (N_20776,N_16925,N_15900);
xor U20777 (N_20777,N_15328,N_15912);
and U20778 (N_20778,N_18087,N_16419);
nand U20779 (N_20779,N_17993,N_18924);
or U20780 (N_20780,N_16383,N_16365);
nor U20781 (N_20781,N_19191,N_15826);
nor U20782 (N_20782,N_19425,N_19421);
nand U20783 (N_20783,N_17392,N_15341);
nand U20784 (N_20784,N_19847,N_19008);
xor U20785 (N_20785,N_15488,N_18104);
nor U20786 (N_20786,N_16308,N_15043);
or U20787 (N_20787,N_18226,N_15002);
nor U20788 (N_20788,N_17475,N_18920);
nor U20789 (N_20789,N_15654,N_16640);
xnor U20790 (N_20790,N_16978,N_16903);
xor U20791 (N_20791,N_15456,N_19928);
or U20792 (N_20792,N_15671,N_17680);
or U20793 (N_20793,N_16063,N_17777);
and U20794 (N_20794,N_19804,N_15337);
and U20795 (N_20795,N_18091,N_16158);
nand U20796 (N_20796,N_17024,N_16883);
xnor U20797 (N_20797,N_15292,N_19096);
xor U20798 (N_20798,N_15256,N_15966);
xor U20799 (N_20799,N_15599,N_17038);
nor U20800 (N_20800,N_17055,N_18139);
and U20801 (N_20801,N_19117,N_17189);
nor U20802 (N_20802,N_15925,N_16760);
xnor U20803 (N_20803,N_15580,N_16784);
nand U20804 (N_20804,N_16969,N_16633);
nor U20805 (N_20805,N_17638,N_17872);
nand U20806 (N_20806,N_15652,N_16409);
xor U20807 (N_20807,N_17090,N_16047);
or U20808 (N_20808,N_18520,N_18348);
and U20809 (N_20809,N_15332,N_17188);
or U20810 (N_20810,N_17289,N_16053);
xnor U20811 (N_20811,N_17947,N_17559);
and U20812 (N_20812,N_17504,N_16568);
xor U20813 (N_20813,N_17458,N_19972);
nor U20814 (N_20814,N_16109,N_18056);
or U20815 (N_20815,N_19832,N_18779);
xnor U20816 (N_20816,N_19338,N_15180);
xor U20817 (N_20817,N_17552,N_16129);
and U20818 (N_20818,N_19716,N_19263);
or U20819 (N_20819,N_19444,N_15331);
nor U20820 (N_20820,N_17057,N_17069);
and U20821 (N_20821,N_16394,N_18134);
or U20822 (N_20822,N_15662,N_19265);
nand U20823 (N_20823,N_17376,N_16139);
nand U20824 (N_20824,N_15034,N_19778);
xor U20825 (N_20825,N_16496,N_18313);
xnor U20826 (N_20826,N_17723,N_16865);
nand U20827 (N_20827,N_15216,N_17902);
or U20828 (N_20828,N_15516,N_16649);
xnor U20829 (N_20829,N_19497,N_19138);
xnor U20830 (N_20830,N_18465,N_17807);
or U20831 (N_20831,N_19160,N_15387);
and U20832 (N_20832,N_15117,N_17173);
nor U20833 (N_20833,N_18400,N_17507);
nand U20834 (N_20834,N_18891,N_18750);
xnor U20835 (N_20835,N_17255,N_15278);
xor U20836 (N_20836,N_15161,N_18572);
nand U20837 (N_20837,N_17597,N_18072);
and U20838 (N_20838,N_19296,N_19993);
xnor U20839 (N_20839,N_19539,N_18031);
and U20840 (N_20840,N_17964,N_18099);
xor U20841 (N_20841,N_17871,N_18754);
nand U20842 (N_20842,N_19244,N_17743);
and U20843 (N_20843,N_15176,N_19802);
and U20844 (N_20844,N_18876,N_19656);
nor U20845 (N_20845,N_17685,N_17494);
nand U20846 (N_20846,N_16125,N_17999);
xor U20847 (N_20847,N_17593,N_15326);
nor U20848 (N_20848,N_19167,N_16914);
nor U20849 (N_20849,N_18324,N_15362);
or U20850 (N_20850,N_15869,N_19520);
or U20851 (N_20851,N_18745,N_17966);
xor U20852 (N_20852,N_19702,N_18711);
nand U20853 (N_20853,N_15075,N_19224);
nor U20854 (N_20854,N_16279,N_18898);
nor U20855 (N_20855,N_17960,N_19290);
nor U20856 (N_20856,N_18384,N_17323);
nand U20857 (N_20857,N_19879,N_19187);
or U20858 (N_20858,N_15407,N_16884);
nor U20859 (N_20859,N_17197,N_16647);
and U20860 (N_20860,N_17954,N_15384);
xnor U20861 (N_20861,N_16895,N_19071);
nor U20862 (N_20862,N_15254,N_19333);
nor U20863 (N_20863,N_18092,N_19181);
xor U20864 (N_20864,N_16615,N_18462);
and U20865 (N_20865,N_19632,N_15297);
and U20866 (N_20866,N_18466,N_17113);
or U20867 (N_20867,N_17292,N_15090);
xor U20868 (N_20868,N_17071,N_18410);
and U20869 (N_20869,N_16243,N_15785);
and U20870 (N_20870,N_16225,N_17422);
nand U20871 (N_20871,N_16836,N_16963);
nor U20872 (N_20872,N_19058,N_18862);
xor U20873 (N_20873,N_17729,N_18025);
or U20874 (N_20874,N_19628,N_18120);
nor U20875 (N_20875,N_18156,N_18305);
nand U20876 (N_20876,N_17252,N_19939);
nor U20877 (N_20877,N_16874,N_16171);
and U20878 (N_20878,N_18420,N_18640);
xor U20879 (N_20879,N_16692,N_19304);
xnor U20880 (N_20880,N_15306,N_18269);
nand U20881 (N_20881,N_19798,N_18213);
nand U20882 (N_20882,N_19572,N_16128);
or U20883 (N_20883,N_15410,N_19400);
nor U20884 (N_20884,N_16762,N_17575);
nor U20885 (N_20885,N_19510,N_17989);
or U20886 (N_20886,N_17614,N_15574);
xor U20887 (N_20887,N_15491,N_15664);
xnor U20888 (N_20888,N_16843,N_16352);
nand U20889 (N_20889,N_16327,N_17895);
xnor U20890 (N_20890,N_16543,N_16124);
or U20891 (N_20891,N_16862,N_18188);
and U20892 (N_20892,N_18129,N_18277);
nand U20893 (N_20893,N_16856,N_15170);
nand U20894 (N_20894,N_16149,N_16304);
nor U20895 (N_20895,N_15442,N_15076);
nand U20896 (N_20896,N_19536,N_18427);
nand U20897 (N_20897,N_16059,N_16740);
or U20898 (N_20898,N_16154,N_15511);
nor U20899 (N_20899,N_15805,N_18770);
or U20900 (N_20900,N_19100,N_18032);
xor U20901 (N_20901,N_15471,N_18761);
or U20902 (N_20902,N_17286,N_17689);
nand U20903 (N_20903,N_17198,N_15690);
nand U20904 (N_20904,N_17439,N_18371);
xnor U20905 (N_20905,N_18043,N_18353);
nand U20906 (N_20906,N_17430,N_19611);
and U20907 (N_20907,N_16512,N_17250);
xor U20908 (N_20908,N_15500,N_15674);
or U20909 (N_20909,N_15776,N_19642);
nor U20910 (N_20910,N_17487,N_16766);
nor U20911 (N_20911,N_16016,N_16629);
and U20912 (N_20912,N_18827,N_17405);
xor U20913 (N_20913,N_19900,N_15259);
or U20914 (N_20914,N_17224,N_19667);
and U20915 (N_20915,N_17159,N_19973);
or U20916 (N_20916,N_19870,N_18958);
xor U20917 (N_20917,N_17901,N_19902);
and U20918 (N_20918,N_18218,N_15821);
nand U20919 (N_20919,N_15736,N_15726);
and U20920 (N_20920,N_16470,N_16824);
nand U20921 (N_20921,N_19711,N_19158);
nor U20922 (N_20922,N_17127,N_15121);
xor U20923 (N_20923,N_17533,N_17891);
and U20924 (N_20924,N_17303,N_19106);
xnor U20925 (N_20925,N_19438,N_19112);
nor U20926 (N_20926,N_16070,N_19105);
nor U20927 (N_20927,N_17180,N_16695);
nand U20928 (N_20928,N_19511,N_17787);
nor U20929 (N_20929,N_17963,N_17133);
or U20930 (N_20930,N_15692,N_16854);
nand U20931 (N_20931,N_17545,N_17116);
nand U20932 (N_20932,N_16912,N_16140);
nor U20933 (N_20933,N_16189,N_19035);
xnor U20934 (N_20934,N_16514,N_17318);
and U20935 (N_20935,N_16078,N_15945);
xnor U20936 (N_20936,N_18901,N_18073);
or U20937 (N_20937,N_17908,N_18590);
or U20938 (N_20938,N_19455,N_18626);
nor U20939 (N_20939,N_17026,N_17427);
or U20940 (N_20940,N_16396,N_17751);
or U20941 (N_20941,N_15485,N_19885);
and U20942 (N_20942,N_17825,N_16055);
and U20943 (N_20943,N_18161,N_19129);
nor U20944 (N_20944,N_17052,N_15956);
nand U20945 (N_20945,N_18463,N_17598);
or U20946 (N_20946,N_18052,N_16094);
nor U20947 (N_20947,N_15525,N_17629);
or U20948 (N_20948,N_17176,N_18461);
nand U20949 (N_20949,N_16179,N_15408);
nor U20950 (N_20950,N_18817,N_15760);
and U20951 (N_20951,N_18001,N_17934);
xnor U20952 (N_20952,N_17195,N_15573);
xnor U20953 (N_20953,N_17028,N_17857);
or U20954 (N_20954,N_15317,N_18524);
nor U20955 (N_20955,N_18981,N_15984);
nor U20956 (N_20956,N_18244,N_15649);
nor U20957 (N_20957,N_17984,N_16783);
nand U20958 (N_20958,N_15284,N_18438);
nor U20959 (N_20959,N_16757,N_19976);
and U20960 (N_20960,N_16218,N_18395);
xnor U20961 (N_20961,N_19651,N_16678);
nor U20962 (N_20962,N_16863,N_17497);
and U20963 (N_20963,N_19243,N_17034);
and U20964 (N_20964,N_17260,N_19944);
nand U20965 (N_20965,N_18748,N_18616);
xnor U20966 (N_20966,N_15113,N_15789);
nor U20967 (N_20967,N_18003,N_17105);
nand U20968 (N_20968,N_15746,N_15338);
and U20969 (N_20969,N_16481,N_16891);
nand U20970 (N_20970,N_16306,N_15368);
xnor U20971 (N_20971,N_18696,N_19085);
xor U20972 (N_20972,N_15459,N_19291);
xnor U20973 (N_20973,N_18265,N_17092);
nor U20974 (N_20974,N_18169,N_18783);
xnor U20975 (N_20975,N_18982,N_17223);
nand U20976 (N_20976,N_16727,N_18431);
nor U20977 (N_20977,N_18449,N_15249);
xor U20978 (N_20978,N_16472,N_17371);
or U20979 (N_20979,N_16322,N_16389);
xnor U20980 (N_20980,N_19065,N_15871);
nor U20981 (N_20981,N_17279,N_18890);
or U20982 (N_20982,N_18391,N_15385);
nand U20983 (N_20983,N_19176,N_19274);
nand U20984 (N_20984,N_18322,N_17035);
nand U20985 (N_20985,N_18036,N_16168);
nand U20986 (N_20986,N_16498,N_17591);
and U20987 (N_20987,N_17351,N_17031);
and U20988 (N_20988,N_15279,N_18795);
and U20989 (N_20989,N_15048,N_18079);
and U20990 (N_20990,N_17087,N_17199);
and U20991 (N_20991,N_18753,N_19846);
or U20992 (N_20992,N_19695,N_17758);
nand U20993 (N_20993,N_16776,N_18154);
or U20994 (N_20994,N_15157,N_16687);
or U20995 (N_20995,N_16324,N_19729);
or U20996 (N_20996,N_19055,N_19130);
xnor U20997 (N_20997,N_18076,N_16417);
xor U20998 (N_20998,N_16084,N_17337);
or U20999 (N_20999,N_17262,N_16719);
or U21000 (N_21000,N_17995,N_18793);
and U21001 (N_21001,N_17402,N_16266);
nor U21002 (N_21002,N_16556,N_19723);
and U21003 (N_21003,N_15810,N_19411);
and U21004 (N_21004,N_18386,N_15653);
xnor U21005 (N_21005,N_18534,N_16880);
and U21006 (N_21006,N_17242,N_16855);
nor U21007 (N_21007,N_16671,N_16430);
or U21008 (N_21008,N_19194,N_15543);
or U21009 (N_21009,N_15255,N_18633);
and U21010 (N_21010,N_19402,N_15729);
and U21011 (N_21011,N_18634,N_18777);
nor U21012 (N_21012,N_15914,N_19923);
and U21013 (N_21013,N_16111,N_18137);
nand U21014 (N_21014,N_15705,N_16866);
xnor U21015 (N_21015,N_16612,N_16667);
nor U21016 (N_21016,N_17754,N_15118);
nor U21017 (N_21017,N_16673,N_17981);
nand U21018 (N_21018,N_17516,N_18934);
xor U21019 (N_21019,N_19735,N_15017);
nor U21020 (N_21020,N_18274,N_18577);
xnor U21021 (N_21021,N_19816,N_15361);
and U21022 (N_21022,N_19509,N_15045);
xnor U21023 (N_21023,N_18067,N_19466);
nand U21024 (N_21024,N_16700,N_19255);
nand U21025 (N_21025,N_16756,N_19305);
nand U21026 (N_21026,N_19546,N_15011);
nand U21027 (N_21027,N_15634,N_16331);
nand U21028 (N_21028,N_15545,N_16215);
nor U21029 (N_21029,N_16940,N_18601);
and U21030 (N_21030,N_15908,N_16737);
nor U21031 (N_21031,N_16303,N_19553);
nor U21032 (N_21032,N_19982,N_17158);
or U21033 (N_21033,N_19230,N_16054);
and U21034 (N_21034,N_19017,N_19384);
and U21035 (N_21035,N_18096,N_17043);
nor U21036 (N_21036,N_18548,N_15655);
nand U21037 (N_21037,N_15794,N_15032);
or U21038 (N_21038,N_17804,N_16930);
nand U21039 (N_21039,N_19826,N_19472);
xnor U21040 (N_21040,N_19674,N_19314);
or U21041 (N_21041,N_15579,N_17683);
nor U21042 (N_21042,N_15398,N_19462);
nor U21043 (N_21043,N_18246,N_19620);
or U21044 (N_21044,N_17839,N_17830);
nand U21045 (N_21045,N_15938,N_18726);
or U21046 (N_21046,N_17012,N_16837);
or U21047 (N_21047,N_16858,N_16934);
or U21048 (N_21048,N_18415,N_18831);
or U21049 (N_21049,N_16477,N_15492);
xnor U21050 (N_21050,N_18865,N_18533);
or U21051 (N_21051,N_18238,N_18352);
xnor U21052 (N_21052,N_15926,N_18445);
and U21053 (N_21053,N_18846,N_19430);
nor U21054 (N_21054,N_16412,N_15815);
nor U21055 (N_21055,N_15643,N_16965);
xnor U21056 (N_21056,N_19694,N_17744);
nand U21057 (N_21057,N_19709,N_17045);
nor U21058 (N_21058,N_15919,N_18697);
and U21059 (N_21059,N_15688,N_16528);
or U21060 (N_21060,N_17630,N_15222);
nand U21061 (N_21061,N_16119,N_18254);
and U21062 (N_21062,N_17988,N_19929);
nor U21063 (N_21063,N_18443,N_17360);
and U21064 (N_21064,N_16746,N_19257);
or U21065 (N_21065,N_17082,N_17446);
nand U21066 (N_21066,N_16190,N_18848);
or U21067 (N_21067,N_17500,N_15082);
xor U21068 (N_21068,N_16454,N_18967);
nor U21069 (N_21069,N_16012,N_17657);
nor U21070 (N_21070,N_18935,N_17918);
xor U21071 (N_21071,N_18781,N_18927);
and U21072 (N_21072,N_16957,N_16782);
or U21073 (N_21073,N_16178,N_18205);
and U21074 (N_21074,N_15049,N_19987);
and U21075 (N_21075,N_18749,N_19909);
nor U21076 (N_21076,N_18954,N_16959);
nor U21077 (N_21077,N_17291,N_19358);
nor U21078 (N_21078,N_17101,N_16953);
nand U21079 (N_21079,N_18885,N_15103);
nand U21080 (N_21080,N_16062,N_19373);
xor U21081 (N_21081,N_19386,N_19582);
xnor U21082 (N_21082,N_19734,N_19122);
nand U21083 (N_21083,N_19649,N_16092);
xor U21084 (N_21084,N_15775,N_18684);
or U21085 (N_21085,N_17525,N_19617);
xor U21086 (N_21086,N_17856,N_15921);
and U21087 (N_21087,N_16689,N_16121);
nand U21088 (N_21088,N_15801,N_16585);
and U21089 (N_21089,N_16075,N_16468);
nand U21090 (N_21090,N_19531,N_15379);
nand U21091 (N_21091,N_17297,N_16191);
nor U21092 (N_21092,N_16571,N_17646);
and U21093 (N_21093,N_17730,N_15063);
xor U21094 (N_21094,N_15383,N_17020);
or U21095 (N_21095,N_17733,N_15780);
or U21096 (N_21096,N_18756,N_16502);
nor U21097 (N_21097,N_19760,N_16435);
nand U21098 (N_21098,N_15095,N_17536);
xnor U21099 (N_21099,N_17852,N_18922);
or U21100 (N_21100,N_18625,N_19753);
or U21101 (N_21101,N_18380,N_16787);
nand U21102 (N_21102,N_16254,N_17328);
or U21103 (N_21103,N_18679,N_19086);
nand U21104 (N_21104,N_19473,N_17979);
nor U21105 (N_21105,N_19590,N_18515);
nor U21106 (N_21106,N_15285,N_15183);
nor U21107 (N_21107,N_15340,N_16000);
nor U21108 (N_21108,N_18251,N_17039);
nand U21109 (N_21109,N_15694,N_19527);
or U21110 (N_21110,N_15730,N_18017);
or U21111 (N_21111,N_18728,N_17675);
xor U21112 (N_21112,N_17459,N_17930);
nor U21113 (N_21113,N_15797,N_16420);
and U21114 (N_21114,N_17467,N_19287);
nand U21115 (N_21115,N_19615,N_16142);
xnor U21116 (N_21116,N_17433,N_16030);
nand U21117 (N_21117,N_17962,N_17134);
nand U21118 (N_21118,N_15784,N_16564);
or U21119 (N_21119,N_15635,N_15404);
or U21120 (N_21120,N_19605,N_18439);
xnor U21121 (N_21121,N_19313,N_17210);
nor U21122 (N_21122,N_19303,N_18928);
and U21123 (N_21123,N_16195,N_16983);
and U21124 (N_21124,N_18661,N_15772);
and U21125 (N_21125,N_16548,N_19917);
nand U21126 (N_21126,N_19141,N_16292);
nand U21127 (N_21127,N_19264,N_15143);
and U21128 (N_21128,N_18095,N_19001);
xnor U21129 (N_21129,N_18994,N_18575);
xor U21130 (N_21130,N_15396,N_19370);
xor U21131 (N_21131,N_17311,N_18563);
xor U21132 (N_21132,N_19686,N_15008);
nor U21133 (N_21133,N_18135,N_17763);
xor U21134 (N_21134,N_19538,N_17893);
nor U21135 (N_21135,N_15311,N_19652);
nand U21136 (N_21136,N_18382,N_18145);
and U21137 (N_21137,N_18356,N_17927);
nand U21138 (N_21138,N_16845,N_15174);
xnor U21139 (N_21139,N_18050,N_18100);
nor U21140 (N_21140,N_19999,N_15248);
xor U21141 (N_21141,N_16565,N_15336);
and U21142 (N_21142,N_17840,N_17479);
nand U21143 (N_21143,N_18452,N_17236);
or U21144 (N_21144,N_17299,N_16408);
nand U21145 (N_21145,N_16748,N_15064);
xnor U21146 (N_21146,N_15261,N_17099);
nand U21147 (N_21147,N_19299,N_18671);
nand U21148 (N_21148,N_18782,N_16575);
nand U21149 (N_21149,N_15529,N_19567);
nor U21150 (N_21150,N_17771,N_18702);
and U21151 (N_21151,N_17549,N_18195);
xor U21152 (N_21152,N_17718,N_19292);
nand U21153 (N_21153,N_17650,N_15661);
nand U21154 (N_21154,N_15957,N_15062);
xnor U21155 (N_21155,N_17813,N_19453);
nor U21156 (N_21156,N_17154,N_19593);
and U21157 (N_21157,N_15817,N_18051);
or U21158 (N_21158,N_18121,N_18701);
nand U21159 (N_21159,N_15932,N_16011);
nor U21160 (N_21160,N_16908,N_17806);
nand U21161 (N_21161,N_17756,N_19925);
nand U21162 (N_21162,N_19518,N_16653);
or U21163 (N_21163,N_16955,N_15100);
or U21164 (N_21164,N_19226,N_15591);
nand U21165 (N_21165,N_17359,N_18060);
nor U21166 (N_21166,N_17278,N_18225);
and U21167 (N_21167,N_15660,N_19200);
nor U21168 (N_21168,N_17413,N_17596);
xor U21169 (N_21169,N_16141,N_16767);
nor U21170 (N_21170,N_16573,N_15534);
nor U21171 (N_21171,N_16018,N_19118);
xnor U21172 (N_21172,N_15501,N_15504);
xnor U21173 (N_21173,N_18642,N_18902);
nand U21174 (N_21174,N_18974,N_15327);
nor U21175 (N_21175,N_19948,N_18477);
nand U21176 (N_21176,N_18281,N_19859);
or U21177 (N_21177,N_15646,N_18818);
nand U21178 (N_21178,N_16182,N_17873);
nor U21179 (N_21179,N_18428,N_15171);
xnor U21180 (N_21180,N_19718,N_18537);
or U21181 (N_21181,N_18527,N_15148);
nor U21182 (N_21182,N_15346,N_16159);
nor U21183 (N_21183,N_15620,N_19476);
nor U21184 (N_21184,N_18344,N_19830);
nor U21185 (N_21185,N_19289,N_15093);
xnor U21186 (N_21186,N_17620,N_16796);
nand U21187 (N_21187,N_18825,N_19726);
and U21188 (N_21188,N_15928,N_15233);
nand U21189 (N_21189,N_17760,N_19459);
xnor U21190 (N_21190,N_16073,N_17203);
or U21191 (N_21191,N_19666,N_16516);
or U21192 (N_21192,N_15641,N_17702);
xnor U21193 (N_21193,N_18612,N_15146);
or U21194 (N_21194,N_17330,N_18546);
nand U21195 (N_21195,N_15042,N_16071);
xnor U21196 (N_21196,N_19498,N_17992);
and U21197 (N_21197,N_15046,N_16205);
and U21198 (N_21198,N_18131,N_15862);
nand U21199 (N_21199,N_17698,N_19212);
and U21200 (N_21200,N_15723,N_16680);
nor U21201 (N_21201,N_17200,N_15967);
xor U21202 (N_21202,N_18170,N_18230);
or U21203 (N_21203,N_16581,N_19810);
nand U21204 (N_21204,N_16614,N_18334);
xnor U21205 (N_21205,N_16001,N_19204);
nor U21206 (N_21206,N_17149,N_17789);
nor U21207 (N_21207,N_19136,N_19316);
and U21208 (N_21208,N_15198,N_15190);
nor U21209 (N_21209,N_17904,N_17973);
nand U21210 (N_21210,N_15260,N_17866);
or U21211 (N_21211,N_17987,N_19178);
and U21212 (N_21212,N_18774,N_16493);
nor U21213 (N_21213,N_17382,N_19782);
and U21214 (N_21214,N_17434,N_18875);
and U21215 (N_21215,N_19616,N_15390);
nand U21216 (N_21216,N_17868,N_18629);
and U21217 (N_21217,N_18514,N_15725);
or U21218 (N_21218,N_17668,N_16797);
or U21219 (N_21219,N_19014,N_15226);
xnor U21220 (N_21220,N_15172,N_18681);
nor U21221 (N_21221,N_17132,N_17523);
or U21222 (N_21222,N_15060,N_18933);
xor U21223 (N_21223,N_17177,N_16230);
and U21224 (N_21224,N_18422,N_17074);
nand U21225 (N_21225,N_16550,N_17736);
nor U21226 (N_21226,N_15553,N_18667);
and U21227 (N_21227,N_16233,N_16421);
xor U21228 (N_21228,N_15149,N_18210);
xor U21229 (N_21229,N_17022,N_19174);
xnor U21230 (N_21230,N_19451,N_18678);
nand U21231 (N_21231,N_16214,N_19589);
nor U21232 (N_21232,N_18283,N_18404);
or U21233 (N_21233,N_15258,N_17416);
or U21234 (N_21234,N_18838,N_18914);
nand U21235 (N_21235,N_19663,N_19913);
and U21236 (N_21236,N_17421,N_15791);
xnor U21237 (N_21237,N_18080,N_17375);
and U21238 (N_21238,N_18389,N_18198);
xnor U21239 (N_21239,N_18128,N_16669);
and U21240 (N_21240,N_16877,N_16873);
and U21241 (N_21241,N_18192,N_17951);
nor U21242 (N_21242,N_16852,N_16896);
nor U21243 (N_21243,N_19634,N_18693);
or U21244 (N_21244,N_17576,N_17938);
nand U21245 (N_21245,N_17261,N_19797);
xnor U21246 (N_21246,N_16731,N_19364);
and U21247 (N_21247,N_16777,N_16497);
or U21248 (N_21248,N_17118,N_19152);
xnor U21249 (N_21249,N_15530,N_15438);
and U21250 (N_21250,N_16261,N_19854);
or U21251 (N_21251,N_16582,N_18716);
and U21252 (N_21252,N_18894,N_16655);
xnor U21253 (N_21253,N_16307,N_18622);
xor U21254 (N_21254,N_16822,N_15487);
nor U21255 (N_21255,N_15349,N_16258);
xor U21256 (N_21256,N_18148,N_17135);
and U21257 (N_21257,N_19720,N_15510);
and U21258 (N_21258,N_19053,N_15563);
or U21259 (N_21259,N_19561,N_17900);
nor U21260 (N_21260,N_17048,N_19121);
nand U21261 (N_21261,N_18504,N_16936);
or U21262 (N_21262,N_19559,N_18700);
and U21263 (N_21263,N_19748,N_17503);
nand U21264 (N_21264,N_18879,N_17578);
nor U21265 (N_21265,N_16734,N_19119);
or U21266 (N_21266,N_15979,N_18315);
and U21267 (N_21267,N_17456,N_18237);
nand U21268 (N_21268,N_18730,N_19475);
nand U21269 (N_21269,N_17447,N_16363);
and U21270 (N_21270,N_17486,N_19310);
nor U21271 (N_21271,N_17287,N_18019);
xnor U21272 (N_21272,N_19064,N_15128);
nor U21273 (N_21273,N_18993,N_18860);
or U21274 (N_21274,N_19662,N_17824);
nand U21275 (N_21275,N_15899,N_15127);
and U21276 (N_21276,N_16291,N_18585);
xnor U21277 (N_21277,N_16277,N_18268);
nor U21278 (N_21278,N_15452,N_18275);
nor U21279 (N_21279,N_19763,N_15364);
nor U21280 (N_21280,N_19237,N_15004);
or U21281 (N_21281,N_18290,N_15054);
xor U21282 (N_21282,N_18866,N_17473);
or U21283 (N_21283,N_19454,N_17706);
nand U21284 (N_21284,N_18089,N_18498);
nand U21285 (N_21285,N_17621,N_15832);
nand U21286 (N_21286,N_17379,N_16992);
or U21287 (N_21287,N_17929,N_16196);
and U21288 (N_21288,N_19612,N_18245);
nor U21289 (N_21289,N_15071,N_16593);
xnor U21290 (N_21290,N_19163,N_18641);
or U21291 (N_21291,N_17161,N_15314);
nor U21292 (N_21292,N_18499,N_15192);
or U21293 (N_21293,N_15998,N_19789);
xnor U21294 (N_21294,N_16213,N_16761);
nand U21295 (N_21295,N_17765,N_18516);
nand U21296 (N_21296,N_17346,N_17986);
xor U21297 (N_21297,N_15901,N_18773);
nand U21298 (N_21298,N_18026,N_19888);
nand U21299 (N_21299,N_18508,N_19808);
xnor U21300 (N_21300,N_16505,N_16351);
nand U21301 (N_21301,N_15450,N_19591);
xor U21302 (N_21302,N_18925,N_15155);
xor U21303 (N_21303,N_16714,N_17179);
or U21304 (N_21304,N_17233,N_17950);
or U21305 (N_21305,N_17700,N_18455);
xor U21306 (N_21306,N_18673,N_16947);
nand U21307 (N_21307,N_16552,N_17854);
xnor U21308 (N_21308,N_16414,N_17762);
nand U21309 (N_21309,N_15989,N_15187);
and U21310 (N_21310,N_17899,N_19139);
nand U21311 (N_21311,N_19259,N_16570);
or U21312 (N_21312,N_19504,N_16041);
nand U21313 (N_21313,N_18144,N_17072);
nor U21314 (N_21314,N_16599,N_16294);
or U21315 (N_21315,N_16459,N_15245);
and U21316 (N_21316,N_19706,N_15028);
and U21317 (N_21317,N_16439,N_17424);
nand U21318 (N_21318,N_17058,N_19253);
nand U21319 (N_21319,N_15335,N_19385);
nor U21320 (N_21320,N_17527,N_15752);
and U21321 (N_21321,N_18992,N_15535);
and U21322 (N_21322,N_17772,N_19645);
or U21323 (N_21323,N_15473,N_17403);
xor U21324 (N_21324,N_18722,N_17170);
or U21325 (N_21325,N_19345,N_18939);
xnor U21326 (N_21326,N_17468,N_19192);
or U21327 (N_21327,N_16187,N_18328);
and U21328 (N_21328,N_15417,N_15970);
nor U21329 (N_21329,N_17660,N_18485);
or U21330 (N_21330,N_18229,N_19359);
nor U21331 (N_21331,N_16136,N_17506);
nor U21332 (N_21332,N_16286,N_17448);
xnor U21333 (N_21333,N_15083,N_17687);
nor U21334 (N_21334,N_19705,N_16480);
or U21335 (N_21335,N_15592,N_18433);
nor U21336 (N_21336,N_18255,N_18063);
nand U21337 (N_21337,N_19363,N_19088);
xor U21338 (N_21338,N_15214,N_18636);
nor U21339 (N_21339,N_15041,N_19533);
nor U21340 (N_21340,N_18863,N_19766);
nand U21341 (N_21341,N_18526,N_18132);
xnor U21342 (N_21342,N_15308,N_19738);
and U21343 (N_21343,N_17049,N_18646);
or U21344 (N_21344,N_19535,N_18823);
and U21345 (N_21345,N_15806,N_17524);
or U21346 (N_21346,N_19604,N_18852);
and U21347 (N_21347,N_17820,N_18074);
nor U21348 (N_21348,N_18854,N_16248);
xnor U21349 (N_21349,N_18118,N_15420);
and U21350 (N_21350,N_15839,N_18311);
or U21351 (N_21351,N_19783,N_19443);
and U21352 (N_21352,N_18085,N_16038);
nand U21353 (N_21353,N_15616,N_16192);
nand U21354 (N_21354,N_16317,N_15519);
and U21355 (N_21355,N_19635,N_19940);
nand U21356 (N_21356,N_15167,N_18820);
nand U21357 (N_21357,N_16013,N_18707);
and U21358 (N_21358,N_19412,N_17604);
nor U21359 (N_21359,N_17285,N_17925);
nand U21360 (N_21360,N_17053,N_19239);
and U21361 (N_21361,N_18258,N_15024);
and U21362 (N_21362,N_16631,N_17480);
nor U21363 (N_21363,N_19156,N_18024);
nor U21364 (N_21364,N_17229,N_15428);
nand U21365 (N_21365,N_19685,N_17212);
nand U21366 (N_21366,N_17477,N_17401);
and U21367 (N_21367,N_19665,N_15264);
nor U21368 (N_21368,N_17111,N_16799);
and U21369 (N_21369,N_19043,N_18942);
nand U21370 (N_21370,N_15218,N_18203);
and U21371 (N_21371,N_16222,N_19951);
xnor U21372 (N_21372,N_18379,N_17705);
and U21373 (N_21373,N_18539,N_19080);
nand U21374 (N_21374,N_18215,N_17878);
or U21375 (N_21375,N_19684,N_17389);
xnor U21376 (N_21376,N_16968,N_15582);
xor U21377 (N_21377,N_18658,N_18398);
nand U21378 (N_21378,N_17555,N_17645);
xnor U21379 (N_21379,N_19749,N_16758);
nand U21380 (N_21380,N_17143,N_17885);
xor U21381 (N_21381,N_15745,N_18692);
and U21382 (N_21382,N_18593,N_18302);
or U21383 (N_21383,N_16123,N_19743);
nor U21384 (N_21384,N_18023,N_19703);
nand U21385 (N_21385,N_18607,N_19011);
and U21386 (N_21386,N_19197,N_16014);
or U21387 (N_21387,N_17745,N_19784);
nand U21388 (N_21388,N_15689,N_18907);
xnor U21389 (N_21389,N_17589,N_16694);
xor U21390 (N_21390,N_18071,N_16897);
nor U21391 (N_21391,N_19301,N_19677);
nand U21392 (N_21392,N_19312,N_15342);
nand U21393 (N_21393,N_16759,N_16463);
nor U21394 (N_21394,N_18759,N_17658);
nand U21395 (N_21395,N_17923,N_15749);
nor U21396 (N_21396,N_16022,N_17443);
xor U21397 (N_21397,N_16020,N_15802);
and U21398 (N_21398,N_17915,N_15804);
and U21399 (N_21399,N_15056,N_19343);
xnor U21400 (N_21400,N_17659,N_16941);
and U21401 (N_21401,N_15734,N_17274);
nand U21402 (N_21402,N_17222,N_17117);
nor U21403 (N_21403,N_19010,N_18663);
or U21404 (N_21404,N_19161,N_17068);
or U21405 (N_21405,N_18719,N_15569);
and U21406 (N_21406,N_15619,N_18411);
or U21407 (N_21407,N_16098,N_17599);
nand U21408 (N_21408,N_16157,N_17104);
xor U21409 (N_21409,N_19252,N_18776);
or U21410 (N_21410,N_19835,N_15370);
or U21411 (N_21411,N_19469,N_18930);
and U21412 (N_21412,N_19447,N_16390);
or U21413 (N_21413,N_19404,N_17780);
xnor U21414 (N_21414,N_15656,N_15066);
nor U21415 (N_21415,N_19081,N_15313);
nor U21416 (N_21416,N_16411,N_16763);
nor U21417 (N_21417,N_18751,N_16994);
xor U21418 (N_21418,N_18660,N_17182);
and U21419 (N_21419,N_16721,N_15720);
nand U21420 (N_21420,N_15441,N_19699);
nand U21421 (N_21421,N_15318,N_18123);
nand U21422 (N_21422,N_16927,N_16864);
and U21423 (N_21423,N_19123,N_16590);
and U21424 (N_21424,N_15571,N_19487);
nand U21425 (N_21425,N_19873,N_18189);
or U21426 (N_21426,N_16933,N_18381);
or U21427 (N_21427,N_16755,N_18312);
and U21428 (N_21428,N_17949,N_18358);
and U21429 (N_21429,N_18292,N_19742);
xnor U21430 (N_21430,N_17247,N_19285);
xnor U21431 (N_21431,N_16344,N_15395);
and U21432 (N_21432,N_15917,N_15253);
nor U21433 (N_21433,N_19858,N_18929);
and U21434 (N_21434,N_15612,N_16993);
xnor U21435 (N_21435,N_17633,N_19282);
nand U21436 (N_21436,N_17005,N_16127);
and U21437 (N_21437,N_18996,N_18163);
xnor U21438 (N_21438,N_15890,N_16939);
or U21439 (N_21439,N_18909,N_18142);
nand U21440 (N_21440,N_15711,N_16180);
nand U21441 (N_21441,N_19791,N_16471);
or U21442 (N_21442,N_16326,N_15293);
and U21443 (N_21443,N_18887,N_17661);
or U21444 (N_21444,N_18510,N_16398);
and U21445 (N_21445,N_15493,N_18695);
nor U21446 (N_21446,N_19208,N_16790);
nor U21447 (N_21447,N_15532,N_17102);
and U21448 (N_21448,N_15808,N_15321);
xnor U21449 (N_21449,N_17393,N_18437);
xnor U21450 (N_21450,N_18916,N_19108);
or U21451 (N_21451,N_17586,N_16670);
and U21452 (N_21452,N_18986,N_15678);
nand U21453 (N_21453,N_19361,N_16705);
and U21454 (N_21454,N_17167,N_15111);
nand U21455 (N_21455,N_17737,N_15870);
xnor U21456 (N_21456,N_17268,N_16210);
or U21457 (N_21457,N_19586,N_18212);
nor U21458 (N_21458,N_18457,N_19225);
nor U21459 (N_21459,N_18506,N_19166);
or U21460 (N_21460,N_19306,N_15526);
and U21461 (N_21461,N_18511,N_17735);
nor U21462 (N_21462,N_19467,N_15982);
nor U21463 (N_21463,N_15732,N_16074);
nand U21464 (N_21464,N_15215,N_19550);
nor U21465 (N_21465,N_17696,N_18746);
xnor U21466 (N_21466,N_19381,N_18989);
xnor U21467 (N_21467,N_16563,N_15533);
nand U21468 (N_21468,N_17432,N_17490);
and U21469 (N_21469,N_17716,N_16848);
nand U21470 (N_21470,N_19470,N_16812);
and U21471 (N_21471,N_17059,N_15568);
nor U21472 (N_21472,N_18336,N_16566);
nand U21473 (N_21473,N_16634,N_19728);
or U21474 (N_21474,N_18005,N_17829);
or U21475 (N_21475,N_17935,N_19501);
nor U21476 (N_21476,N_15489,N_19526);
and U21477 (N_21477,N_19062,N_15109);
nor U21478 (N_21478,N_19934,N_15262);
nand U21479 (N_21479,N_16738,N_18767);
nor U21480 (N_21480,N_19436,N_16293);
nor U21481 (N_21481,N_15003,N_19026);
and U21482 (N_21482,N_18547,N_19689);
and U21483 (N_21483,N_19627,N_19060);
nor U21484 (N_21484,N_18478,N_19745);
or U21485 (N_21485,N_15755,N_18469);
or U21486 (N_21486,N_17147,N_16268);
nand U21487 (N_21487,N_15015,N_15241);
xnor U21488 (N_21488,N_19405,N_16077);
nor U21489 (N_21489,N_15010,N_15604);
and U21490 (N_21490,N_16557,N_19247);
and U21491 (N_21491,N_19168,N_19515);
nor U21492 (N_21492,N_15166,N_19721);
nor U21493 (N_21493,N_18041,N_15741);
nand U21494 (N_21494,N_17157,N_16574);
nand U21495 (N_21495,N_17488,N_15052);
nor U21496 (N_21496,N_19872,N_15959);
and U21497 (N_21497,N_16150,N_19033);
and U21498 (N_21498,N_18408,N_18355);
or U21499 (N_21499,N_18674,N_17556);
xor U21500 (N_21500,N_17231,N_15911);
nand U21501 (N_21501,N_18227,N_17415);
and U21502 (N_21502,N_15937,N_17204);
xor U21503 (N_21503,N_15439,N_19754);
xnor U21504 (N_21504,N_19279,N_18686);
xnor U21505 (N_21505,N_16521,N_17027);
and U21506 (N_21506,N_18373,N_19047);
nor U21507 (N_21507,N_16275,N_18102);
or U21508 (N_21508,N_18291,N_18493);
and U21509 (N_21509,N_19968,N_15263);
xor U21510 (N_21510,N_16364,N_16588);
xnor U21511 (N_21511,N_17688,N_18039);
xor U21512 (N_21512,N_17924,N_16911);
or U21513 (N_21513,N_19741,N_18162);
or U21514 (N_21514,N_19989,N_19903);
and U21515 (N_21515,N_16591,N_17306);
nand U21516 (N_21516,N_18578,N_18900);
or U21517 (N_21517,N_15666,N_15727);
nand U21518 (N_21518,N_19125,N_16422);
nor U21519 (N_21519,N_15244,N_18014);
nor U21520 (N_21520,N_19079,N_17853);
and U21521 (N_21521,N_16035,N_18206);
nand U21522 (N_21522,N_19009,N_15708);
xnor U21523 (N_21523,N_16551,N_16602);
and U21524 (N_21524,N_16713,N_16654);
nor U21525 (N_21525,N_18544,N_19190);
xnor U21526 (N_21526,N_18880,N_17440);
or U21527 (N_21527,N_19127,N_17968);
nand U21528 (N_21528,N_17326,N_15469);
nand U21529 (N_21529,N_15607,N_19625);
or U21530 (N_21530,N_19552,N_15650);
nor U21531 (N_21531,N_15523,N_15923);
or U21532 (N_21532,N_17811,N_15369);
xnor U21533 (N_21533,N_16278,N_19493);
xnor U21534 (N_21534,N_15016,N_19733);
xor U21535 (N_21535,N_17671,N_15400);
and U21536 (N_21536,N_18984,N_18522);
nor U21537 (N_21537,N_19137,N_19329);
and U21538 (N_21538,N_17920,N_17818);
or U21539 (N_21539,N_18610,N_18766);
xnor U21540 (N_21540,N_19298,N_19623);
and U21541 (N_21541,N_18772,N_17010);
and U21542 (N_21542,N_17270,N_17582);
nand U21543 (N_21543,N_17652,N_19320);
xor U21544 (N_21544,N_16244,N_15716);
nand U21545 (N_21545,N_15983,N_15611);
or U21546 (N_21546,N_17495,N_19034);
nor U21547 (N_21547,N_16507,N_18044);
nor U21548 (N_21548,N_17953,N_16239);
or U21549 (N_21549,N_19277,N_17166);
or U21550 (N_21550,N_15953,N_17374);
xor U21551 (N_21551,N_15840,N_17776);
nand U21552 (N_21552,N_19958,N_16096);
and U21553 (N_21553,N_15145,N_15751);
and U21554 (N_21554,N_16395,N_18742);
and U21555 (N_21555,N_17186,N_18152);
nand U21556 (N_21556,N_16601,N_16108);
nor U21557 (N_21557,N_15107,N_18840);
and U21558 (N_21558,N_19073,N_18160);
or U21559 (N_21559,N_17691,N_19276);
nand U21560 (N_21560,N_19415,N_15783);
or U21561 (N_21561,N_19353,N_16801);
and U21562 (N_21562,N_18167,N_17692);
xor U21563 (N_21563,N_17819,N_17603);
or U21564 (N_21564,N_16808,N_17795);
and U21565 (N_21565,N_16842,N_15419);
nor U21566 (N_21566,N_15603,N_17437);
nand U21567 (N_21567,N_16334,N_15150);
and U21568 (N_21568,N_17568,N_17919);
nor U21569 (N_21569,N_17969,N_19675);
xor U21570 (N_21570,N_15759,N_19731);
nand U21571 (N_21571,N_18517,N_15257);
nor U21572 (N_21572,N_19964,N_17512);
nand U21573 (N_21573,N_18809,N_16887);
nand U21574 (N_21574,N_17304,N_18574);
xnor U21575 (N_21575,N_15975,N_19072);
nor U21576 (N_21576,N_16302,N_18826);
nor U21577 (N_21577,N_18596,N_15483);
or U21578 (N_21578,N_15137,N_18789);
xor U21579 (N_21579,N_16132,N_15329);
nand U21580 (N_21580,N_18733,N_16661);
and U21581 (N_21581,N_15536,N_17917);
or U21582 (N_21582,N_17983,N_18138);
and U21583 (N_21583,N_16811,N_16217);
nor U21584 (N_21584,N_17471,N_15951);
xnor U21585 (N_21585,N_15294,N_18260);
nand U21586 (N_21586,N_19563,N_16024);
and U21587 (N_21587,N_18040,N_19875);
and U21588 (N_21588,N_19054,N_17774);
nand U21589 (N_21589,N_15163,N_15356);
nor U21590 (N_21590,N_17928,N_19201);
or U21591 (N_21591,N_19057,N_15944);
xnor U21592 (N_21592,N_18124,N_16604);
xnor U21593 (N_21593,N_19895,N_15502);
or U21594 (N_21594,N_17844,N_16522);
xor U21595 (N_21595,N_17115,N_18871);
and U21596 (N_21596,N_19691,N_16558);
or U21597 (N_21597,N_16381,N_15219);
nand U21598 (N_21598,N_16044,N_15134);
or U21599 (N_21599,N_18083,N_18859);
and U21600 (N_21600,N_18647,N_17008);
nand U21601 (N_21601,N_18509,N_18441);
or U21602 (N_21602,N_18279,N_19850);
xnor U21603 (N_21603,N_17612,N_18972);
xnor U21604 (N_21604,N_18150,N_19765);
xnor U21605 (N_21605,N_18448,N_17344);
and U21606 (N_21606,N_15151,N_16683);
and U21607 (N_21607,N_18110,N_17842);
nor U21608 (N_21608,N_15575,N_15472);
and U21609 (N_21609,N_16985,N_19431);
nor U21610 (N_21610,N_16815,N_19059);
nand U21611 (N_21611,N_16006,N_19896);
xnor U21612 (N_21612,N_19202,N_17300);
nor U21613 (N_21613,N_15000,N_15823);
or U21614 (N_21614,N_19114,N_19070);
and U21615 (N_21615,N_16844,N_17493);
xor U21616 (N_21616,N_19669,N_18393);
xor U21617 (N_21617,N_19946,N_15559);
and U21618 (N_21618,N_18567,N_19774);
and U21619 (N_21619,N_15835,N_18627);
and U21620 (N_21620,N_19007,N_15058);
or U21621 (N_21621,N_19424,N_19165);
nor U21622 (N_21622,N_17541,N_16651);
nand U21623 (N_21623,N_19029,N_15228);
or U21624 (N_21624,N_15541,N_19414);
and U21625 (N_21625,N_17740,N_17267);
or U21626 (N_21626,N_16069,N_16194);
and U21627 (N_21627,N_18151,N_15051);
nor U21628 (N_21628,N_15659,N_18937);
xnor U21629 (N_21629,N_17089,N_16857);
or U21630 (N_21630,N_19827,N_16082);
xor U21631 (N_21631,N_16090,N_16885);
and U21632 (N_21632,N_18047,N_19932);
or U21633 (N_21633,N_16741,N_19971);
xor U21634 (N_21634,N_17888,N_15468);
or U21635 (N_21635,N_17602,N_15626);
nor U21636 (N_21636,N_19916,N_16152);
and U21637 (N_21637,N_16120,N_18977);
and U21638 (N_21638,N_16720,N_15375);
or U21639 (N_21639,N_17709,N_15423);
xor U21640 (N_21640,N_19270,N_16870);
xnor U21641 (N_21641,N_18173,N_15737);
nand U21642 (N_21642,N_17060,N_16469);
or U21643 (N_21643,N_18740,N_18472);
nor U21644 (N_21644,N_19758,N_19440);
and U21645 (N_21645,N_19592,N_17332);
and U21646 (N_21646,N_19769,N_18687);
nand U21647 (N_21647,N_18426,N_19849);
or U21648 (N_21648,N_19772,N_18704);
or U21649 (N_21649,N_15722,N_15050);
nand U21650 (N_21650,N_16265,N_16535);
or U21651 (N_21651,N_17004,N_15670);
or U21652 (N_21652,N_16028,N_15355);
nand U21653 (N_21653,N_19013,N_17861);
or U21654 (N_21654,N_16036,N_15193);
or U21655 (N_21655,N_17670,N_15159);
and U21656 (N_21656,N_16646,N_17206);
and U21657 (N_21657,N_17768,N_18157);
and U21658 (N_21658,N_17056,N_19213);
and U21659 (N_21659,N_17042,N_15426);
xnor U21660 (N_21660,N_19680,N_17320);
or U21661 (N_21661,N_18957,N_16052);
nand U21662 (N_21662,N_17013,N_15924);
xor U21663 (N_21663,N_16161,N_16151);
nand U21664 (N_21664,N_19914,N_18808);
or U21665 (N_21665,N_19907,N_17406);
nor U21666 (N_21666,N_17305,N_15246);
nand U21667 (N_21667,N_16209,N_19113);
nand U21668 (N_21668,N_18116,N_15644);
nor U21669 (N_21669,N_16260,N_19630);
nand U21670 (N_21670,N_19991,N_18919);
nor U21671 (N_21671,N_17785,N_19116);
nand U21672 (N_21672,N_15769,N_17216);
and U21673 (N_21673,N_17256,N_17226);
nor U21674 (N_21674,N_16311,N_17570);
nand U21675 (N_21675,N_15997,N_19851);
xnor U21676 (N_21676,N_19933,N_15514);
and U21677 (N_21677,N_19602,N_15130);
nand U21678 (N_21678,N_19050,N_17192);
xnor U21679 (N_21679,N_15778,N_15954);
xor U21680 (N_21680,N_17033,N_16617);
and U21681 (N_21681,N_18771,N_18813);
xnor U21682 (N_21682,N_19037,N_18075);
nor U21683 (N_21683,N_17959,N_18632);
nor U21684 (N_21684,N_17592,N_15624);
nor U21685 (N_21685,N_17808,N_17441);
nor U21686 (N_21686,N_17190,N_19371);
or U21687 (N_21687,N_15399,N_18464);
nand U21688 (N_21688,N_18082,N_16882);
nand U21689 (N_21689,N_15971,N_19222);
nor U21690 (N_21690,N_18507,N_18187);
or U21691 (N_21691,N_16519,N_17139);
and U21692 (N_21692,N_19945,N_15415);
and U21693 (N_21693,N_18458,N_19502);
and U21694 (N_21694,N_15842,N_15710);
and U21695 (N_21695,N_15290,N_15271);
xnor U21696 (N_21696,N_15358,N_17881);
nand U21697 (N_21697,N_18497,N_17172);
nor U21698 (N_21698,N_18185,N_19067);
nor U21699 (N_21699,N_15731,N_17673);
or U21700 (N_21700,N_17431,N_19983);
and U21701 (N_21701,N_19725,N_19581);
or U21702 (N_21702,N_16513,N_19557);
xor U21703 (N_21703,N_17152,N_19028);
or U21704 (N_21704,N_18802,N_16684);
or U21705 (N_21705,N_16725,N_18581);
xnor U21706 (N_21706,N_17067,N_15458);
nor U21707 (N_21707,N_19626,N_15205);
or U21708 (N_21708,N_15135,N_17041);
nand U21709 (N_21709,N_15006,N_16621);
nor U21710 (N_21710,N_19092,N_19281);
nand U21711 (N_21711,N_15623,N_15961);
xnor U21712 (N_21712,N_17551,N_15232);
nor U21713 (N_21713,N_15413,N_16532);
nor U21714 (N_21714,N_16475,N_16622);
nand U21715 (N_21715,N_17851,N_16931);
nand U21716 (N_21716,N_16686,N_16089);
xnor U21717 (N_21717,N_18330,N_17977);
or U21718 (N_21718,N_15462,N_19777);
nand U21719 (N_21719,N_18171,N_17770);
xor U21720 (N_21720,N_15353,N_15325);
nor U21721 (N_21721,N_19251,N_16081);
or U21722 (N_21722,N_18556,N_19366);
xor U21723 (N_21723,N_18653,N_19456);
nor U21724 (N_21724,N_16100,N_17955);
or U21725 (N_21725,N_17384,N_19863);
nor U21726 (N_21726,N_18532,N_19555);
xor U21727 (N_21727,N_16517,N_17230);
nor U21728 (N_21728,N_15513,N_17874);
and U21729 (N_21729,N_18997,N_19668);
xor U21730 (N_21730,N_16500,N_17491);
nor U21731 (N_21731,N_16201,N_16474);
or U21732 (N_21732,N_15394,N_15538);
and U21733 (N_21733,N_16107,N_16462);
or U21734 (N_21734,N_17492,N_19173);
or U21735 (N_21735,N_19227,N_19697);
xnor U21736 (N_21736,N_18383,N_16252);
nand U21737 (N_21737,N_19886,N_18184);
nand U21738 (N_21738,N_16147,N_15371);
xor U21739 (N_21739,N_18685,N_15168);
xor U21740 (N_21740,N_17624,N_16285);
xnor U21741 (N_21741,N_15816,N_17369);
or U21742 (N_21742,N_16715,N_19732);
and U21743 (N_21743,N_19133,N_16682);
nand U21744 (N_21744,N_15947,N_18202);
or U21745 (N_21745,N_16025,N_18608);
and U21746 (N_21746,N_19464,N_18955);
xnor U21747 (N_21747,N_15126,N_16583);
or U21748 (N_21748,N_17940,N_17699);
nor U21749 (N_21749,N_15281,N_15481);
nand U21750 (N_21750,N_15834,N_18961);
and U21751 (N_21751,N_17734,N_16023);
nor U21752 (N_21752,N_16298,N_19399);
nor U21753 (N_21753,N_19150,N_16458);
xor U21754 (N_21754,N_15070,N_18888);
nor U21755 (N_21755,N_15165,N_15894);
nand U21756 (N_21756,N_16898,N_17562);
xor U21757 (N_21757,N_15393,N_19646);
xor U21758 (N_21758,N_16716,N_18211);
xnor U21759 (N_21759,N_17110,N_18460);
nor U21760 (N_21760,N_16520,N_16712);
xnor U21761 (N_21761,N_15018,N_18755);
xor U21762 (N_21762,N_15479,N_17676);
nor U21763 (N_21763,N_16401,N_15080);
or U21764 (N_21764,N_16099,N_17558);
xor U21765 (N_21765,N_18349,N_15139);
nand U21766 (N_21766,N_19347,N_15105);
nand U21767 (N_21767,N_19795,N_16788);
nand U21768 (N_21768,N_15424,N_15270);
nand U21769 (N_21769,N_16418,N_15750);
nand U21770 (N_21770,N_19354,N_18209);
xnor U21771 (N_21771,N_18300,N_18530);
or U21772 (N_21772,N_16926,N_18094);
nand U21773 (N_21773,N_16764,N_16378);
and U21774 (N_21774,N_15560,N_19103);
and U21775 (N_21775,N_19115,N_19969);
nand U21776 (N_21776,N_16175,N_16407);
and U21777 (N_21777,N_18980,N_18332);
or U21778 (N_21778,N_17572,N_19943);
or U21779 (N_21779,N_18568,N_15119);
nand U21780 (N_21780,N_16101,N_17064);
and U21781 (N_21781,N_15182,N_17142);
and U21782 (N_21782,N_15542,N_15747);
nand U21783 (N_21783,N_15152,N_16234);
and U21784 (N_21784,N_15081,N_18561);
and U21785 (N_21785,N_16325,N_19641);
nand U21786 (N_21786,N_18280,N_15994);
and U21787 (N_21787,N_16371,N_16950);
nand U21788 (N_21788,N_16460,N_15848);
nor U21789 (N_21789,N_17832,N_15546);
xnor U21790 (N_21790,N_18158,N_16045);
nor U21791 (N_21791,N_18287,N_19864);
nand U21792 (N_21792,N_18576,N_19041);
nor U21793 (N_21793,N_18650,N_17537);
and U21794 (N_21794,N_18357,N_19528);
xor U21795 (N_21795,N_15094,N_18814);
or U21796 (N_21796,N_19554,N_16906);
or U21797 (N_21797,N_16494,N_15252);
nor U21798 (N_21798,N_16429,N_16473);
or U21799 (N_21799,N_18688,N_16894);
or U21800 (N_21800,N_15905,N_17543);
or U21801 (N_21801,N_15099,N_19374);
nor U21802 (N_21802,N_15786,N_17580);
nor U21803 (N_21803,N_18314,N_19162);
nor U21804 (N_21804,N_19318,N_19519);
nand U21805 (N_21805,N_15958,N_17867);
nand U21806 (N_21806,N_15845,N_16966);
and U21807 (N_21807,N_16853,N_19266);
xor U21808 (N_21808,N_18273,N_19715);
xor U21809 (N_21809,N_16056,N_17298);
nand U21810 (N_21810,N_19346,N_16984);
xor U21811 (N_21811,N_15554,N_15478);
nor U21812 (N_21812,N_15467,N_19937);
nand U21813 (N_21813,N_15274,N_16273);
or U21814 (N_21814,N_16735,N_18232);
nor U21815 (N_21815,N_18175,N_16486);
or U21816 (N_21816,N_19209,N_17062);
and U21817 (N_21817,N_17931,N_15590);
xor U21818 (N_21818,N_18316,N_18800);
and U21819 (N_21819,N_17727,N_15812);
nand U21820 (N_21820,N_19486,N_16237);
or U21821 (N_21821,N_18564,N_18960);
xor U21822 (N_21822,N_19434,N_19499);
and U21823 (N_21823,N_18816,N_18963);
or U21824 (N_21824,N_15850,N_16579);
or U21825 (N_21825,N_19771,N_16595);
nor U21826 (N_21826,N_17837,N_16426);
nor U21827 (N_21827,N_19235,N_15762);
or U21828 (N_21828,N_19283,N_19084);
nand U21829 (N_21829,N_15453,N_16828);
xor U21830 (N_21830,N_16376,N_17073);
or U21831 (N_21831,N_15891,N_16823);
nor U21832 (N_21832,N_17887,N_15005);
nor U21833 (N_21833,N_15191,N_16106);
or U21834 (N_21834,N_15627,N_15941);
nor U21835 (N_21835,N_15027,N_16467);
nand U21836 (N_21836,N_17619,N_15756);
xnor U21837 (N_21837,N_17238,N_17941);
xnor U21838 (N_21838,N_18409,N_17347);
xnor U21839 (N_21839,N_19342,N_19217);
xnor U21840 (N_21840,N_19268,N_18008);
or U21841 (N_21841,N_15551,N_15520);
or U21842 (N_21842,N_17006,N_16693);
nand U21843 (N_21843,N_18600,N_17608);
nand U21844 (N_21844,N_16373,N_17594);
nor U21845 (N_21845,N_17485,N_17522);
or U21846 (N_21846,N_15864,N_18338);
nor U21847 (N_21847,N_16330,N_19242);
nor U21848 (N_21848,N_15668,N_16212);
nor U21849 (N_21849,N_19560,N_19762);
or U21850 (N_21850,N_16065,N_17476);
nor U21851 (N_21851,N_15833,N_16750);
nand U21852 (N_21852,N_19082,N_16004);
nor U21853 (N_21853,N_18288,N_16892);
or U21854 (N_21854,N_17483,N_19241);
xor U21855 (N_21855,N_19175,N_17293);
nand U21856 (N_21856,N_16657,N_17822);
xor U21857 (N_21857,N_15565,N_16833);
nand U21858 (N_21858,N_17697,N_18790);
and U21859 (N_21859,N_18714,N_17205);
and U21860 (N_21860,N_15795,N_16228);
and U21861 (N_21861,N_17665,N_15990);
nand U21862 (N_21862,N_16445,N_15883);
and U21863 (N_21863,N_18541,N_18234);
and U21864 (N_21864,N_15642,N_19740);
nand U21865 (N_21865,N_18015,N_15618);
or U21866 (N_21866,N_18760,N_15675);
xor U21867 (N_21867,N_19562,N_16736);
and U21868 (N_21868,N_18354,N_18529);
and U21869 (N_21869,N_15758,N_16995);
or U21870 (N_21870,N_16321,N_16800);
nor U21871 (N_21871,N_15047,N_15735);
or U21872 (N_21872,N_16080,N_15738);
or U21873 (N_21873,N_19687,N_19712);
xor U21874 (N_21874,N_18263,N_17002);
xor U21875 (N_21875,N_15597,N_18595);
xor U21876 (N_21876,N_18775,N_16455);
xor U21877 (N_21877,N_19422,N_19423);
nand U21878 (N_21878,N_16916,N_18197);
or U21879 (N_21879,N_15676,N_15238);
or U21880 (N_21880,N_15929,N_19761);
nor U21881 (N_21881,N_15943,N_17126);
xor U21882 (N_21882,N_18868,N_19111);
nand U21883 (N_21883,N_17096,N_18551);
xor U21884 (N_21884,N_15968,N_17003);
nor U21885 (N_21885,N_17644,N_16501);
and U21886 (N_21886,N_15378,N_17136);
xor U21887 (N_21887,N_19151,N_19376);
and U21888 (N_21888,N_18536,N_15277);
or U21889 (N_21889,N_17388,N_17678);
xnor U21890 (N_21890,N_18359,N_16104);
nand U21891 (N_21891,N_18369,N_15087);
and U21892 (N_21892,N_19334,N_18947);
and U21893 (N_21893,N_16406,N_19974);
or U21894 (N_21894,N_19044,N_16675);
or U21895 (N_21895,N_19821,N_15898);
nand U21896 (N_21896,N_17243,N_16546);
and U21897 (N_21897,N_16806,N_18365);
xor U21898 (N_21898,N_18811,N_17863);
nor U21899 (N_21899,N_18717,N_17341);
xnor U21900 (N_21900,N_16893,N_18824);
nor U21901 (N_21901,N_15189,N_19077);
xor U21902 (N_21902,N_16923,N_17574);
and U21903 (N_21903,N_17295,N_15092);
or U21904 (N_21904,N_18956,N_18592);
and U21905 (N_21905,N_15809,N_15588);
xnor U21906 (N_21906,N_19002,N_19874);
nand U21907 (N_21907,N_15973,N_18109);
nor U21908 (N_21908,N_18591,N_15057);
and U21909 (N_21909,N_18613,N_17769);
or U21910 (N_21910,N_18276,N_16611);
or U21911 (N_21911,N_16872,N_16901);
xor U21912 (N_21912,N_17717,N_18304);
nor U21913 (N_21913,N_16608,N_17860);
or U21914 (N_21914,N_15014,N_17202);
and U21915 (N_21915,N_17616,N_18801);
and U21916 (N_21916,N_19340,N_17890);
nand U21917 (N_21917,N_18549,N_16919);
and U21918 (N_21918,N_18331,N_15448);
xor U21919 (N_21919,N_19566,N_16289);
xnor U21920 (N_21920,N_18361,N_19845);
nor U21921 (N_21921,N_15685,N_18220);
and U21922 (N_21922,N_15640,N_18270);
xnor U21923 (N_21923,N_15363,N_16840);
and U21924 (N_21924,N_15687,N_18708);
and U21925 (N_21925,N_18921,N_15767);
xor U21926 (N_21926,N_16768,N_17240);
or U21927 (N_21927,N_15548,N_15116);
and U21928 (N_21928,N_18267,N_19069);
nor U21929 (N_21929,N_15585,N_16301);
nand U21930 (N_21930,N_15001,N_19205);
xor U21931 (N_21931,N_19576,N_17156);
nor U21932 (N_21932,N_17146,N_19801);
xnor U21933 (N_21933,N_18319,N_18475);
and U21934 (N_21934,N_15288,N_18720);
xor U21935 (N_21935,N_16981,N_16340);
and U21936 (N_21936,N_17187,N_18734);
nor U21937 (N_21937,N_16620,N_16009);
nand U21938 (N_21938,N_18979,N_19996);
xor U21939 (N_21939,N_17566,N_19752);
and U21940 (N_21940,N_17469,N_19393);
nor U21941 (N_21941,N_15077,N_16270);
xnor U21942 (N_21942,N_17429,N_17263);
xor U21943 (N_21943,N_16384,N_17615);
nand U21944 (N_21944,N_16478,N_16185);
xor U21945 (N_21945,N_18306,N_18643);
nor U21946 (N_21946,N_19962,N_15437);
xnor U21947 (N_21947,N_18495,N_17519);
nand U21948 (N_21948,N_17273,N_17050);
xor U21949 (N_21949,N_16701,N_19984);
nor U21950 (N_21950,N_19924,N_18896);
or U21951 (N_21951,N_15713,N_18501);
nor U21952 (N_21952,N_19027,N_15622);
xor U21953 (N_21953,N_15044,N_15949);
nand U21954 (N_21954,N_18069,N_18599);
and U21955 (N_21955,N_19427,N_16416);
xnor U21956 (N_21956,N_19365,N_16017);
nand U21957 (N_21957,N_19109,N_15837);
or U21958 (N_21958,N_19492,N_15617);
and U21959 (N_21959,N_19824,N_15269);
nand U21960 (N_21960,N_17215,N_19474);
or U21961 (N_21961,N_19210,N_18418);
nor U21962 (N_21962,N_18689,N_16173);
nand U21963 (N_21963,N_15447,N_19961);
nor U21964 (N_21964,N_15208,N_19335);
xnor U21965 (N_21965,N_15822,N_16972);
and U21966 (N_21966,N_16229,N_19500);
nand U21967 (N_21967,N_16393,N_18351);
nand U21968 (N_21968,N_16333,N_15096);
or U21969 (N_21969,N_17184,N_17444);
nor U21970 (N_21970,N_18278,N_18877);
xor U21971 (N_21971,N_17080,N_15224);
or U21972 (N_21972,N_16193,N_17460);
nand U21973 (N_21973,N_16049,N_16871);
or U21974 (N_21974,N_19458,N_17368);
or U21975 (N_21975,N_15830,N_16489);
and U21976 (N_21976,N_16909,N_19272);
nor U21977 (N_21977,N_17625,N_18998);
or U21978 (N_21978,N_16729,N_15857);
nor U21979 (N_21979,N_15996,N_15936);
nand U21980 (N_21980,N_17302,N_19587);
or U21981 (N_21981,N_16922,N_17213);
nand U21982 (N_21982,N_15073,N_19534);
xor U21983 (N_21983,N_17397,N_17079);
and U21984 (N_21984,N_18219,N_17843);
nand U21985 (N_21985,N_19841,N_16819);
nor U21986 (N_21986,N_19857,N_18432);
or U21987 (N_21987,N_18851,N_17781);
xor U21988 (N_21988,N_17112,N_17814);
or U21989 (N_21989,N_16487,N_17065);
xor U21990 (N_21990,N_19800,N_17539);
xor U21991 (N_21991,N_16064,N_15289);
or U21992 (N_21992,N_15484,N_19186);
nor U21993 (N_21993,N_19814,N_15544);
nand U21994 (N_21994,N_19957,N_16998);
or U21995 (N_21995,N_16240,N_16778);
and U21996 (N_21996,N_15435,N_17656);
or U21997 (N_21997,N_15365,N_15454);
nor U21998 (N_21998,N_17239,N_18065);
or U21999 (N_21999,N_19032,N_18709);
and U22000 (N_22000,N_16606,N_17585);
nand U22001 (N_22001,N_16638,N_19673);
nand U22002 (N_22002,N_18959,N_19785);
or U22003 (N_22003,N_18481,N_19094);
and U22004 (N_22004,N_17361,N_15600);
nor U22005 (N_22005,N_15798,N_17000);
xor U22006 (N_22006,N_17047,N_19867);
nor U22007 (N_22007,N_17514,N_17438);
xnor U22008 (N_22008,N_16580,N_19295);
or U22009 (N_22009,N_19530,N_17712);
or U22010 (N_22010,N_16184,N_17643);
and U22011 (N_22011,N_17802,N_15131);
and U22012 (N_22012,N_15564,N_17724);
and U22013 (N_22013,N_16057,N_15712);
nand U22014 (N_22014,N_18521,N_17131);
xor U22015 (N_22015,N_17623,N_18573);
xor U22016 (N_22016,N_18513,N_18147);
or U22017 (N_22017,N_19495,N_17284);
xnor U22018 (N_22018,N_16924,N_19288);
or U22019 (N_22019,N_16499,N_17812);
or U22020 (N_22020,N_16058,N_16164);
nor U22021 (N_22021,N_18554,N_15696);
and U22022 (N_22022,N_19350,N_17322);
or U22023 (N_22023,N_16162,N_15055);
or U22024 (N_22024,N_19482,N_19220);
and U22025 (N_22025,N_18078,N_18735);
nand U22026 (N_22026,N_15418,N_17605);
nand U22027 (N_22027,N_15416,N_19890);
or U22028 (N_22028,N_15645,N_16314);
and U22029 (N_22029,N_16805,N_18010);
and U22030 (N_22030,N_17098,N_15680);
and U22031 (N_22031,N_19607,N_17826);
xnor U22032 (N_22032,N_15763,N_18683);
xnor U22033 (N_22033,N_15993,N_18999);
nand U22034 (N_22034,N_15115,N_18480);
or U22035 (N_22035,N_17879,N_19182);
xnor U22036 (N_22036,N_19724,N_15351);
or U22037 (N_22037,N_15486,N_15697);
nor U22038 (N_22038,N_16977,N_15962);
xor U22039 (N_22039,N_15091,N_18550);
xnor U22040 (N_22040,N_15333,N_19927);
xor U22041 (N_22041,N_19146,N_16466);
nand U22042 (N_22042,N_18881,N_15451);
xor U22043 (N_22043,N_17453,N_19240);
and U22044 (N_22044,N_19978,N_18378);
nor U22045 (N_22045,N_16295,N_19380);
nand U22046 (N_22046,N_19061,N_16817);
or U22047 (N_22047,N_19391,N_17847);
xnor U22048 (N_22048,N_16553,N_18677);
and U22049 (N_22049,N_18248,N_19759);
xor U22050 (N_22050,N_15873,N_16881);
and U22051 (N_22051,N_18366,N_18446);
nor U22052 (N_22052,N_18502,N_19413);
and U22053 (N_22053,N_16785,N_18699);
and U22054 (N_22054,N_16112,N_19021);
xor U22055 (N_22055,N_15495,N_16446);
nor U22056 (N_22056,N_17108,N_15142);
xnor U22057 (N_22057,N_16353,N_16392);
xor U22058 (N_22058,N_18343,N_15893);
xor U22059 (N_22059,N_15701,N_19930);
xnor U22060 (N_22060,N_18983,N_17569);
or U22061 (N_22061,N_16698,N_16464);
or U22062 (N_22062,N_18857,N_19585);
nand U22063 (N_22063,N_19231,N_16413);
and U22064 (N_22064,N_17880,N_18703);
and U22065 (N_22065,N_15153,N_16506);
nand U22066 (N_22066,N_17208,N_18525);
xnor U22067 (N_22067,N_19435,N_18179);
xnor U22068 (N_22068,N_19882,N_18101);
or U22069 (N_22069,N_16839,N_17277);
nor U22070 (N_22070,N_17627,N_17362);
nor U22071 (N_22071,N_15987,N_15267);
and U22072 (N_22072,N_18286,N_19513);
nand U22073 (N_22073,N_17897,N_17864);
nand U22074 (N_22074,N_15700,N_15175);
nor U22075 (N_22075,N_15939,N_19488);
or U22076 (N_22076,N_19516,N_15578);
xnor U22077 (N_22077,N_15210,N_18307);
nand U22078 (N_22078,N_17352,N_15779);
xnor U22079 (N_22079,N_18949,N_19024);
or U22080 (N_22080,N_17961,N_15841);
nand U22081 (N_22081,N_16087,N_19450);
and U22082 (N_22082,N_16227,N_18177);
and U22083 (N_22083,N_16804,N_17385);
and U22084 (N_22084,N_17682,N_15517);
or U22085 (N_22085,N_17081,N_16452);
or U22086 (N_22086,N_19144,N_15902);
and U22087 (N_22087,N_15323,N_17560);
xnor U22088 (N_22088,N_19919,N_17317);
and U22089 (N_22089,N_15768,N_18084);
xnor U22090 (N_22090,N_18768,N_15765);
xnor U22091 (N_22091,N_17241,N_15787);
xnor U22092 (N_22092,N_18605,N_15429);
or U22093 (N_22093,N_18815,N_17451);
and U22094 (N_22094,N_18694,N_17315);
and U22095 (N_22095,N_16188,N_15406);
or U22096 (N_22096,N_16223,N_16987);
nand U22097 (N_22097,N_17513,N_19525);
nand U22098 (N_22098,N_16754,N_19967);
nor U22099 (N_22099,N_16589,N_18571);
nand U22100 (N_22100,N_18821,N_15884);
or U22101 (N_22101,N_16433,N_17076);
nor U22102 (N_22102,N_18111,N_15301);
nor U22103 (N_22103,N_15978,N_19892);
nand U22104 (N_22104,N_19736,N_15372);
and U22105 (N_22105,N_15343,N_15295);
xnor U22106 (N_22106,N_18538,N_18950);
nand U22107 (N_22107,N_18401,N_15409);
nor U22108 (N_22108,N_16825,N_19419);
nand U22109 (N_22109,N_19599,N_15392);
nor U22110 (N_22110,N_15348,N_17109);
xor U22111 (N_22111,N_18471,N_17409);
xor U22112 (N_22112,N_19102,N_18406);
or U22113 (N_22113,N_17869,N_16708);
xnor U22114 (N_22114,N_15539,N_15158);
nor U22115 (N_22115,N_17704,N_18293);
nand U22116 (N_22116,N_19837,N_18737);
nand U22117 (N_22117,N_18604,N_18033);
nand U22118 (N_22118,N_16888,N_15980);
or U22119 (N_22119,N_18494,N_17714);
nor U22120 (N_22120,N_15039,N_19030);
nor U22121 (N_22121,N_15764,N_18055);
or U22122 (N_22122,N_16598,N_18321);
and U22123 (N_22123,N_18662,N_17815);
nor U22124 (N_22124,N_19820,N_17939);
nor U22125 (N_22125,N_18987,N_16627);
or U22126 (N_22126,N_18672,N_18675);
and U22127 (N_22127,N_17708,N_17084);
xor U22128 (N_22128,N_19142,N_17400);
nor U22129 (N_22129,N_15106,N_16547);
or U22130 (N_22130,N_19558,N_15352);
or U22131 (N_22131,N_18294,N_16504);
and U22132 (N_22132,N_16691,N_18555);
nand U22133 (N_22133,N_17016,N_17214);
and U22134 (N_22134,N_17377,N_18166);
and U22135 (N_22135,N_19871,N_19737);
nor U22136 (N_22136,N_15667,N_17023);
xor U22137 (N_22137,N_15566,N_19248);
nand U22138 (N_22138,N_15896,N_16113);
nor U22139 (N_22139,N_19503,N_16747);
xnor U22140 (N_22140,N_17686,N_18045);
or U22141 (N_22141,N_15584,N_16935);
nand U22142 (N_22142,N_17324,N_16269);
xnor U22143 (N_22143,N_16706,N_19815);
xor U22144 (N_22144,N_18112,N_15177);
nor U22145 (N_22145,N_15636,N_18335);
nor U22146 (N_22146,N_17793,N_17308);
and U22147 (N_22147,N_17398,N_16752);
nand U22148 (N_22148,N_17529,N_16644);
or U22149 (N_22149,N_19481,N_17571);
nor U22150 (N_22150,N_15443,N_17542);
nor U22151 (N_22151,N_16282,N_19597);
nand U22152 (N_22152,N_15431,N_15204);
xnor U22153 (N_22153,N_19496,N_19990);
xnor U22154 (N_22154,N_19018,N_16235);
or U22155 (N_22155,N_15007,N_17998);
nor U22156 (N_22156,N_17151,N_15136);
and U22157 (N_22157,N_16356,N_19887);
nand U22158 (N_22158,N_19403,N_16917);
and U22159 (N_22159,N_15019,N_15401);
and U22160 (N_22160,N_15935,N_17746);
nand U22161 (N_22161,N_18791,N_15965);
nand U22162 (N_22162,N_15463,N_17719);
nor U22163 (N_22163,N_17163,N_19862);
nor U22164 (N_22164,N_15207,N_17701);
nand U22165 (N_22165,N_19975,N_19083);
and U22166 (N_22166,N_16710,N_17370);
nand U22167 (N_22167,N_15531,N_19016);
xnor U22168 (N_22168,N_17283,N_15247);
and U22169 (N_22169,N_17792,N_15630);
nor U22170 (N_22170,N_17461,N_19579);
or U22171 (N_22171,N_15490,N_17248);
nand U22172 (N_22172,N_16890,N_19730);
nand U22173 (N_22173,N_17651,N_19408);
and U22174 (N_22174,N_18609,N_17641);
and U22175 (N_22175,N_15069,N_15856);
or U22176 (N_22176,N_16372,N_18070);
nand U22177 (N_22177,N_15466,N_16555);
or U22178 (N_22178,N_19942,N_16518);
or U22179 (N_22179,N_15380,N_15397);
xnor U22180 (N_22180,N_15412,N_17140);
nand U22181 (N_22181,N_17193,N_18832);
nand U22182 (N_22182,N_15360,N_19931);
nand U22183 (N_22183,N_15188,N_15639);
nor U22184 (N_22184,N_18423,N_15879);
nor U22185 (N_22185,N_15141,N_19377);
xnor U22186 (N_22186,N_16186,N_19379);
nand U22187 (N_22187,N_19223,N_18362);
and U22188 (N_22188,N_19490,N_17466);
xor U22189 (N_22189,N_16346,N_18159);
nand U22190 (N_22190,N_19688,N_17340);
or U22191 (N_22191,N_18988,N_15836);
or U22192 (N_22192,N_18407,N_19267);
or U22193 (N_22193,N_18259,N_15567);
and U22194 (N_22194,N_19091,N_19569);
nor U22195 (N_22195,N_16739,N_19947);
or U22196 (N_22196,N_17288,N_15773);
nand U22197 (N_22197,N_19484,N_18951);
nor U22198 (N_22198,N_18204,N_18165);
nor U22199 (N_22199,N_19098,N_19952);
xnor U22200 (N_22200,N_19865,N_15555);
nor U22201 (N_22201,N_18784,N_16832);
nor U22202 (N_22202,N_15291,N_15197);
nand U22203 (N_22203,N_17794,N_16913);
nand U22204 (N_22204,N_17408,N_16299);
and U22205 (N_22205,N_16539,N_17805);
nor U22206 (N_22206,N_15266,N_19294);
nor U22207 (N_22207,N_17849,N_16603);
nor U22208 (N_22208,N_15948,N_19956);
xnor U22209 (N_22209,N_15123,N_15683);
nor U22210 (N_22210,N_17390,N_16928);
and U22211 (N_22211,N_15350,N_18995);
nor U22212 (N_22212,N_15282,N_19818);
and U22213 (N_22213,N_17994,N_19031);
or U22214 (N_22214,N_18242,N_17587);
and U22215 (N_22215,N_16988,N_17972);
nor U22216 (N_22216,N_16979,N_16697);
or U22217 (N_22217,N_16434,N_17713);
nor U22218 (N_22218,N_17425,N_17395);
nor U22219 (N_22219,N_19428,N_19046);
and U22220 (N_22220,N_19273,N_16060);
or U22221 (N_22221,N_15229,N_18016);
nor U22222 (N_22222,N_16889,N_16597);
xor U22223 (N_22223,N_16172,N_15602);
nand U22224 (N_22224,N_17606,N_19548);
and U22225 (N_22225,N_15916,N_15505);
nor U22226 (N_22226,N_17419,N_17858);
nand U22227 (N_22227,N_18103,N_15774);
xnor U22228 (N_22228,N_16284,N_15910);
xnor U22229 (N_22229,N_19805,N_18906);
xnor U22230 (N_22230,N_19922,N_19622);
xor U22231 (N_22231,N_17782,N_19317);
or U22232 (N_22232,N_15367,N_19610);
xor U22233 (N_22233,N_16122,N_15298);
xnor U22234 (N_22234,N_16846,N_18864);
nor U22235 (N_22235,N_16626,N_15854);
nor U22236 (N_22236,N_18323,N_19218);
or U22237 (N_22237,N_15596,N_17850);
xor U22238 (N_22238,N_16704,N_15460);
nand U22239 (N_22239,N_19727,N_16019);
nand U22240 (N_22240,N_18183,N_18451);
xnor U22241 (N_22241,N_18787,N_19375);
nor U22242 (N_22242,N_16900,N_16544);
nand U22243 (N_22243,N_19796,N_15154);
nand U22244 (N_22244,N_17410,N_18310);
nand U22245 (N_22245,N_19834,N_17896);
nand U22246 (N_22246,N_18272,N_16137);
nor U22247 (N_22247,N_16397,N_19022);
xor U22248 (N_22248,N_15881,N_15250);
or U22249 (N_22249,N_15211,N_15212);
nand U22250 (N_22250,N_19693,N_19460);
or U22251 (N_22251,N_15464,N_15691);
nor U22252 (N_22252,N_19717,N_18337);
nor U22253 (N_22253,N_15818,N_15721);
or U22254 (N_22254,N_15882,N_17165);
nor U22255 (N_22255,N_16288,N_15345);
or U22256 (N_22256,N_17196,N_18542);
xnor U22257 (N_22257,N_17613,N_16427);
nor U22258 (N_22258,N_17739,N_18180);
xnor U22259 (N_22259,N_16117,N_19853);
nor U22260 (N_22260,N_17577,N_19891);
and U22261 (N_22261,N_15059,N_19512);
nor U22262 (N_22262,N_19219,N_16607);
xnor U22263 (N_22263,N_16807,N_16176);
and U22264 (N_22264,N_19893,N_17677);
xnor U22265 (N_22265,N_17235,N_18910);
or U22266 (N_22266,N_16534,N_15698);
and U22267 (N_22267,N_19388,N_17990);
nand U22268 (N_22268,N_16276,N_15877);
nand U22269 (N_22269,N_16572,N_16905);
nand U22270 (N_22270,N_16834,N_16259);
xor U22271 (N_22271,N_17312,N_15803);
xor U22272 (N_22272,N_15853,N_18222);
or U22273 (N_22273,N_18899,N_18440);
and U22274 (N_22274,N_18474,N_16335);
xnor U22275 (N_22275,N_17936,N_19245);
nand U22276 (N_22276,N_15251,N_15201);
and U22277 (N_22277,N_19899,N_17209);
xnor U22278 (N_22278,N_17095,N_15023);
nand U22279 (N_22279,N_16274,N_16991);
nand U22280 (N_22280,N_18639,N_17711);
and U22281 (N_22281,N_18054,N_16618);
nor U22282 (N_22282,N_15040,N_16015);
nand U22283 (N_22283,N_15020,N_15897);
nand U22284 (N_22284,N_19682,N_15307);
and U22285 (N_22285,N_17609,N_16362);
or U22286 (N_22286,N_18196,N_16280);
or U22287 (N_22287,N_18468,N_15402);
nand U22288 (N_22288,N_15132,N_16592);
and U22289 (N_22289,N_19463,N_16369);
or U22290 (N_22290,N_18402,N_17910);
and U22291 (N_22291,N_19756,N_16033);
nor U22292 (N_22292,N_15880,N_17783);
xnor U22293 (N_22293,N_19019,N_16847);
or U22294 (N_22294,N_15120,N_17001);
nor U22295 (N_22295,N_19441,N_17588);
nor U22296 (N_22296,N_15515,N_17264);
nand U22297 (N_22297,N_18628,N_19107);
nand U22298 (N_22298,N_16451,N_19012);
and U22299 (N_22299,N_16524,N_15422);
nand U22300 (N_22300,N_19773,N_15312);
xor U22301 (N_22301,N_15234,N_15506);
nand U22302 (N_22302,N_16529,N_17980);
nor U22303 (N_22303,N_15799,N_17883);
or U22304 (N_22304,N_18467,N_16508);
xor U22305 (N_22305,N_17750,N_18878);
and U22306 (N_22306,N_15733,N_18853);
nor U22307 (N_22307,N_15570,N_18214);
nor U22308 (N_22308,N_19249,N_19986);
xor U22309 (N_22309,N_16167,N_19544);
or U22310 (N_22310,N_19068,N_17310);
or U22311 (N_22311,N_16952,N_19148);
xor U22312 (N_22312,N_16207,N_15875);
xor U22313 (N_22313,N_18725,N_17731);
nor U22314 (N_22314,N_16942,N_17407);
and U22315 (N_22315,N_19164,N_19232);
nor U22316 (N_22316,N_19378,N_17655);
xnor U22317 (N_22317,N_19855,N_17535);
nand U22318 (N_22318,N_16964,N_19959);
or U22319 (N_22319,N_19147,N_18136);
nand U22320 (N_22320,N_18918,N_16361);
or U22321 (N_22321,N_18873,N_17835);
nor U22322 (N_22322,N_15089,N_19629);
nor U22323 (N_22323,N_17976,N_17799);
xor U22324 (N_22324,N_18155,N_18364);
nor U22325 (N_22325,N_18602,N_19494);
xor U22326 (N_22326,N_19357,N_15440);
nor U22327 (N_22327,N_16216,N_18884);
and U22328 (N_22328,N_17100,N_16338);
and U22329 (N_22329,N_15430,N_16144);
nand U22330 (N_22330,N_16134,N_17875);
nor U22331 (N_22331,N_19261,N_18617);
xnor U22332 (N_22332,N_18453,N_19468);
and U22333 (N_22333,N_18785,N_15521);
xor U22334 (N_22334,N_18164,N_17618);
nor U22335 (N_22335,N_18447,N_18153);
and U22336 (N_22336,N_19839,N_17141);
or U22337 (N_22337,N_17358,N_17674);
or U22338 (N_22338,N_17091,N_15985);
nand U22339 (N_22339,N_19938,N_16663);
and U22340 (N_22340,N_18648,N_18841);
nor U22341 (N_22341,N_16974,N_17325);
and U22342 (N_22342,N_18011,N_19908);
or U22343 (N_22343,N_19739,N_15273);
or U22344 (N_22344,N_16051,N_15030);
nand U22345 (N_22345,N_17748,N_15977);
or U22346 (N_22346,N_19124,N_17841);
nand U22347 (N_22347,N_18057,N_15101);
nor U22348 (N_22348,N_18764,N_15272);
nor U22349 (N_22349,N_17378,N_16525);
or U22350 (N_22350,N_16600,N_18829);
xnor U22351 (N_22351,N_19793,N_19457);
or U22352 (N_22352,N_18886,N_16103);
or U22353 (N_22353,N_19269,N_16066);
xor U22354 (N_22354,N_16003,N_19260);
nor U22355 (N_22355,N_19792,N_16312);
nor U22356 (N_22356,N_17725,N_15992);
nand U22357 (N_22357,N_15445,N_16717);
nand U22358 (N_22358,N_16281,N_17124);
nand U22359 (N_22359,N_18223,N_19221);
nor U22360 (N_22360,N_17094,N_17520);
or U22361 (N_22361,N_18946,N_19389);
nand U22362 (N_22362,N_18264,N_17445);
and U22363 (N_22363,N_18724,N_18586);
or U22364 (N_22364,N_16961,N_15125);
nor U22365 (N_22365,N_19356,N_19768);
nor U22366 (N_22366,N_15715,N_16133);
or U22367 (N_22367,N_16821,N_16037);
nand U22368 (N_22368,N_19157,N_17884);
xnor U22369 (N_22369,N_15162,N_17171);
xor U22370 (N_22370,N_18611,N_19545);
or U22371 (N_22371,N_16624,N_18176);
and U22372 (N_22372,N_16029,N_17690);
and U22373 (N_22373,N_17907,N_15300);
or U22374 (N_22374,N_15231,N_15482);
or U22375 (N_22375,N_19609,N_18971);
nand U22376 (N_22376,N_16199,N_19618);
or U22377 (N_22377,N_16975,N_17501);
or U22378 (N_22378,N_17345,N_17548);
xor U22379 (N_22379,N_16357,N_15743);
nor U22380 (N_22380,N_15022,N_17054);
nor U22381 (N_22381,N_16046,N_19003);
and U22382 (N_22382,N_15995,N_17911);
nand U22383 (N_22383,N_18241,N_16561);
or U22384 (N_22384,N_16632,N_16816);
and U22385 (N_22385,N_17316,N_15963);
nand U22386 (N_22386,N_16753,N_19565);
xnor U22387 (N_22387,N_17827,N_18243);
nor U22388 (N_22388,N_18893,N_19781);
nand U22389 (N_22389,N_18892,N_19215);
and U22390 (N_22390,N_17565,N_17282);
nand U22391 (N_22391,N_15436,N_17786);
and U22392 (N_22392,N_17640,N_18425);
nor U22393 (N_22393,N_19860,N_19540);
xnor U22394 (N_22394,N_18049,N_18061);
xnor U22395 (N_22395,N_17234,N_18690);
nor U22396 (N_22396,N_17417,N_17075);
xor U22397 (N_22397,N_15303,N_15647);
nand U22398 (N_22398,N_16997,N_15067);
xnor U22399 (N_22399,N_17251,N_18367);
and U22400 (N_22400,N_17281,N_17595);
or U22401 (N_22401,N_17967,N_16542);
nor U22402 (N_22402,N_19722,N_16786);
and U22403 (N_22403,N_16231,N_16399);
and U22404 (N_22404,N_16386,N_18130);
or U22405 (N_22405,N_19880,N_16665);
or U22406 (N_22406,N_15677,N_19883);
nand U22407 (N_22407,N_18803,N_19661);
nand U22408 (N_22408,N_19395,N_16921);
or U22409 (N_22409,N_19449,N_15374);
or U22410 (N_22410,N_15867,N_19004);
and U22411 (N_22411,N_15503,N_15974);
xor U22412 (N_22412,N_19049,N_15714);
or U22413 (N_22413,N_17457,N_15461);
nor U22414 (N_22414,N_16814,N_17838);
and U22415 (N_22415,N_19751,N_16533);
or U22416 (N_22416,N_17546,N_19183);
nor U22417 (N_22417,N_19311,N_15991);
and U22418 (N_22418,N_18712,N_18257);
or U22419 (N_22419,N_18976,N_17357);
and U22420 (N_22420,N_15347,N_18528);
and U22421 (N_22421,N_19229,N_15072);
nor U22422 (N_22422,N_15433,N_17590);
and U22423 (N_22423,N_19601,N_17125);
and U22424 (N_22424,N_15587,N_19177);
xnor U22425 (N_22425,N_18944,N_16264);
xnor U22426 (N_22426,N_15217,N_18743);
nand U22427 (N_22427,N_19757,N_19410);
xnor U22428 (N_22428,N_15053,N_18931);
nor U22429 (N_22429,N_15320,N_18713);
or U22430 (N_22430,N_15133,N_15679);
xor U22431 (N_22431,N_19505,N_19658);
and U22432 (N_22432,N_16792,N_19036);
or U22433 (N_22433,N_17484,N_19369);
xor U22434 (N_22434,N_17280,N_15280);
and U22435 (N_22435,N_17086,N_15793);
nor U22436 (N_22436,N_15885,N_15744);
and U22437 (N_22437,N_19324,N_17244);
nand U22438 (N_22438,N_18630,N_17025);
and U22439 (N_22439,N_19639,N_19416);
nor U22440 (N_22440,N_16206,N_17845);
nor U22441 (N_22441,N_19979,N_16826);
nand U22442 (N_22442,N_15605,N_18119);
and U22443 (N_22443,N_19644,N_18736);
nand U22444 (N_22444,N_16156,N_19583);
or U22445 (N_22445,N_19214,N_19647);
nand U22446 (N_22446,N_19337,N_19543);
nor U22447 (N_22447,N_16032,N_17499);
nor U22448 (N_22448,N_18412,N_16160);
nor U22449 (N_22449,N_15200,N_18807);
xnor U22450 (N_22450,N_18570,N_18027);
and U22451 (N_22451,N_17946,N_17178);
xnor U22452 (N_22452,N_16310,N_19714);
and U22453 (N_22453,N_17168,N_19196);
xnor U22454 (N_22454,N_16300,N_15709);
or U22455 (N_22455,N_19382,N_15892);
nor U22456 (N_22456,N_16835,N_16795);
nand U22457 (N_22457,N_17411,N_17175);
nand U22458 (N_22458,N_19584,N_17011);
nor U22459 (N_22459,N_19185,N_15695);
nand U22460 (N_22460,N_17584,N_16242);
nand U22461 (N_22461,N_16996,N_15825);
nand U22462 (N_22462,N_16449,N_16677);
nand U22463 (N_22463,N_16594,N_15173);
nand U22464 (N_22464,N_18133,N_17975);
nor U22465 (N_22465,N_19480,N_15455);
xor U22466 (N_22466,N_17348,N_17088);
nor U22467 (N_22467,N_18194,N_15868);
nor U22468 (N_22468,N_17550,N_19066);
and U22469 (N_22469,N_17803,N_15988);
or U22470 (N_22470,N_19571,N_17232);
and U22471 (N_22471,N_15305,N_17120);
nor U22472 (N_22472,N_17343,N_18638);
and U22473 (N_22473,N_15811,N_15084);
nor U22474 (N_22474,N_15432,N_17396);
xnor U22475 (N_22475,N_16355,N_18479);
nand U22476 (N_22476,N_19696,N_17526);
nand U22477 (N_22477,N_19596,N_18850);
or U22478 (N_22478,N_16769,N_17428);
nor U22479 (N_22479,N_16177,N_16316);
nor U22480 (N_22480,N_19383,N_18656);
nor U22481 (N_22481,N_19485,N_18903);
and U22482 (N_22482,N_18968,N_19426);
and U22483 (N_22483,N_19542,N_19483);
nand U22484 (N_22484,N_16443,N_16537);
xnor U22485 (N_22485,N_16660,N_19262);
or U22486 (N_22486,N_15576,N_16438);
or U22487 (N_22487,N_19025,N_18105);
nor U22488 (N_22488,N_19056,N_18317);
xor U22489 (N_22489,N_15777,N_18372);
xnor U22490 (N_22490,N_15108,N_16169);
and U22491 (N_22491,N_16097,N_16174);
nand U22492 (N_22492,N_17426,N_17450);
nand U22493 (N_22493,N_19829,N_15861);
nor U22494 (N_22494,N_16971,N_17037);
or U22495 (N_22495,N_18519,N_19331);
or U22496 (N_22496,N_18849,N_19904);
nor U22497 (N_22497,N_15790,N_19906);
and U22498 (N_22498,N_18491,N_18874);
xnor U22499 (N_22499,N_16403,N_19786);
xor U22500 (N_22500,N_15000,N_18017);
xor U22501 (N_22501,N_17247,N_15189);
nand U22502 (N_22502,N_15739,N_17468);
xor U22503 (N_22503,N_16773,N_17548);
xor U22504 (N_22504,N_15573,N_16392);
nor U22505 (N_22505,N_17774,N_18500);
nor U22506 (N_22506,N_17075,N_18961);
or U22507 (N_22507,N_18678,N_19146);
nand U22508 (N_22508,N_17314,N_17691);
xnor U22509 (N_22509,N_18069,N_16842);
xor U22510 (N_22510,N_15639,N_19458);
xor U22511 (N_22511,N_15659,N_15450);
or U22512 (N_22512,N_15038,N_18789);
or U22513 (N_22513,N_18382,N_16243);
xnor U22514 (N_22514,N_17428,N_19275);
or U22515 (N_22515,N_19683,N_18036);
nor U22516 (N_22516,N_18899,N_18734);
nor U22517 (N_22517,N_15097,N_18310);
and U22518 (N_22518,N_15972,N_16346);
xor U22519 (N_22519,N_17270,N_19238);
and U22520 (N_22520,N_19396,N_16448);
and U22521 (N_22521,N_15890,N_15372);
xnor U22522 (N_22522,N_17214,N_16373);
nor U22523 (N_22523,N_18380,N_18261);
or U22524 (N_22524,N_17078,N_18029);
nand U22525 (N_22525,N_15655,N_18683);
nand U22526 (N_22526,N_18102,N_19120);
and U22527 (N_22527,N_17909,N_19307);
nor U22528 (N_22528,N_17669,N_18028);
nor U22529 (N_22529,N_18191,N_19876);
nor U22530 (N_22530,N_19743,N_17680);
xnor U22531 (N_22531,N_16248,N_18685);
and U22532 (N_22532,N_18832,N_18612);
or U22533 (N_22533,N_18731,N_18960);
nand U22534 (N_22534,N_18429,N_19359);
nand U22535 (N_22535,N_18435,N_15345);
nand U22536 (N_22536,N_17090,N_19822);
and U22537 (N_22537,N_16303,N_16890);
or U22538 (N_22538,N_16624,N_17792);
or U22539 (N_22539,N_17427,N_18523);
or U22540 (N_22540,N_19944,N_16726);
xor U22541 (N_22541,N_18730,N_15503);
or U22542 (N_22542,N_19472,N_16699);
xor U22543 (N_22543,N_16670,N_15007);
nand U22544 (N_22544,N_17803,N_16520);
xnor U22545 (N_22545,N_16490,N_18935);
nor U22546 (N_22546,N_18874,N_16019);
and U22547 (N_22547,N_16912,N_19084);
and U22548 (N_22548,N_17983,N_19047);
nand U22549 (N_22549,N_19193,N_17345);
xor U22550 (N_22550,N_19367,N_15397);
nor U22551 (N_22551,N_15436,N_16525);
and U22552 (N_22552,N_18441,N_19339);
nand U22553 (N_22553,N_15372,N_19908);
and U22554 (N_22554,N_17139,N_15852);
nor U22555 (N_22555,N_18894,N_15097);
nand U22556 (N_22556,N_16582,N_15135);
nand U22557 (N_22557,N_16217,N_17784);
and U22558 (N_22558,N_15515,N_17472);
or U22559 (N_22559,N_17686,N_17472);
nor U22560 (N_22560,N_15326,N_18503);
and U22561 (N_22561,N_15392,N_16978);
or U22562 (N_22562,N_16540,N_17149);
xnor U22563 (N_22563,N_19574,N_15468);
nand U22564 (N_22564,N_19041,N_18761);
and U22565 (N_22565,N_17655,N_17935);
and U22566 (N_22566,N_19012,N_18320);
nand U22567 (N_22567,N_15345,N_16008);
or U22568 (N_22568,N_16554,N_15997);
or U22569 (N_22569,N_19524,N_18538);
nand U22570 (N_22570,N_19717,N_15705);
or U22571 (N_22571,N_15103,N_15094);
nand U22572 (N_22572,N_15512,N_15712);
and U22573 (N_22573,N_15696,N_16916);
xnor U22574 (N_22574,N_18427,N_17677);
nand U22575 (N_22575,N_16929,N_16285);
nand U22576 (N_22576,N_18798,N_18057);
nand U22577 (N_22577,N_19800,N_17787);
nand U22578 (N_22578,N_17539,N_17819);
xnor U22579 (N_22579,N_15249,N_16815);
nand U22580 (N_22580,N_19696,N_17307);
or U22581 (N_22581,N_16779,N_15059);
or U22582 (N_22582,N_15382,N_17695);
xor U22583 (N_22583,N_16343,N_17973);
nand U22584 (N_22584,N_18248,N_18827);
and U22585 (N_22585,N_18288,N_15932);
nand U22586 (N_22586,N_19180,N_15863);
nor U22587 (N_22587,N_18817,N_15604);
and U22588 (N_22588,N_15505,N_15600);
xor U22589 (N_22589,N_19246,N_16939);
or U22590 (N_22590,N_15722,N_19483);
or U22591 (N_22591,N_16492,N_18786);
nand U22592 (N_22592,N_16366,N_18324);
or U22593 (N_22593,N_19441,N_18036);
or U22594 (N_22594,N_17329,N_15190);
nand U22595 (N_22595,N_16999,N_19754);
or U22596 (N_22596,N_17934,N_16329);
nand U22597 (N_22597,N_19639,N_18156);
nor U22598 (N_22598,N_15118,N_16981);
and U22599 (N_22599,N_17999,N_16406);
xor U22600 (N_22600,N_17392,N_18953);
and U22601 (N_22601,N_19461,N_16952);
xor U22602 (N_22602,N_17777,N_17211);
nor U22603 (N_22603,N_17501,N_19681);
and U22604 (N_22604,N_18904,N_17735);
nand U22605 (N_22605,N_19350,N_19416);
and U22606 (N_22606,N_19492,N_19028);
nand U22607 (N_22607,N_18563,N_15841);
xnor U22608 (N_22608,N_19355,N_16270);
xnor U22609 (N_22609,N_15630,N_17665);
nor U22610 (N_22610,N_16035,N_16123);
nor U22611 (N_22611,N_15303,N_16596);
nor U22612 (N_22612,N_18313,N_16058);
nand U22613 (N_22613,N_19255,N_16173);
and U22614 (N_22614,N_15575,N_15706);
or U22615 (N_22615,N_18050,N_15458);
or U22616 (N_22616,N_19885,N_17362);
xnor U22617 (N_22617,N_18424,N_17559);
nor U22618 (N_22618,N_17939,N_18067);
nor U22619 (N_22619,N_16646,N_16214);
nand U22620 (N_22620,N_16718,N_15958);
or U22621 (N_22621,N_17680,N_19125);
nand U22622 (N_22622,N_16216,N_15236);
or U22623 (N_22623,N_16998,N_18419);
or U22624 (N_22624,N_19316,N_17964);
xnor U22625 (N_22625,N_19528,N_15335);
nor U22626 (N_22626,N_17818,N_16830);
or U22627 (N_22627,N_18312,N_17226);
nor U22628 (N_22628,N_16189,N_18411);
or U22629 (N_22629,N_18790,N_15580);
and U22630 (N_22630,N_19669,N_19038);
and U22631 (N_22631,N_16095,N_18296);
nand U22632 (N_22632,N_17825,N_19489);
xnor U22633 (N_22633,N_17026,N_19124);
or U22634 (N_22634,N_19879,N_19976);
nand U22635 (N_22635,N_15027,N_16758);
nand U22636 (N_22636,N_18077,N_18916);
nor U22637 (N_22637,N_19140,N_19248);
xnor U22638 (N_22638,N_15296,N_19363);
nor U22639 (N_22639,N_15769,N_16966);
and U22640 (N_22640,N_17922,N_15155);
or U22641 (N_22641,N_16486,N_19864);
xor U22642 (N_22642,N_18281,N_15676);
or U22643 (N_22643,N_16904,N_19519);
or U22644 (N_22644,N_15057,N_15858);
or U22645 (N_22645,N_15285,N_17794);
nand U22646 (N_22646,N_15408,N_15875);
or U22647 (N_22647,N_18867,N_15681);
nand U22648 (N_22648,N_16772,N_16496);
and U22649 (N_22649,N_19051,N_19877);
nand U22650 (N_22650,N_16217,N_19521);
or U22651 (N_22651,N_18885,N_17625);
or U22652 (N_22652,N_15254,N_15369);
or U22653 (N_22653,N_17534,N_19020);
or U22654 (N_22654,N_15650,N_15533);
or U22655 (N_22655,N_18139,N_15363);
and U22656 (N_22656,N_17987,N_15549);
nor U22657 (N_22657,N_19374,N_18884);
nor U22658 (N_22658,N_15745,N_16696);
nand U22659 (N_22659,N_17964,N_18564);
xnor U22660 (N_22660,N_15146,N_16715);
and U22661 (N_22661,N_18545,N_15702);
and U22662 (N_22662,N_18294,N_16355);
and U22663 (N_22663,N_17831,N_19677);
and U22664 (N_22664,N_17836,N_17912);
xor U22665 (N_22665,N_17595,N_16616);
or U22666 (N_22666,N_17828,N_17933);
nand U22667 (N_22667,N_16406,N_19862);
xor U22668 (N_22668,N_17647,N_18939);
xor U22669 (N_22669,N_15356,N_19589);
nand U22670 (N_22670,N_18460,N_18372);
or U22671 (N_22671,N_17807,N_18713);
nor U22672 (N_22672,N_17668,N_19439);
nor U22673 (N_22673,N_17335,N_15680);
xor U22674 (N_22674,N_15621,N_18008);
nand U22675 (N_22675,N_15855,N_15738);
or U22676 (N_22676,N_18394,N_17964);
xnor U22677 (N_22677,N_18982,N_17382);
and U22678 (N_22678,N_15884,N_19826);
and U22679 (N_22679,N_17602,N_16787);
and U22680 (N_22680,N_19666,N_18465);
xor U22681 (N_22681,N_19018,N_17454);
xor U22682 (N_22682,N_15222,N_17603);
xor U22683 (N_22683,N_15145,N_17226);
nand U22684 (N_22684,N_19089,N_18274);
xnor U22685 (N_22685,N_16079,N_19543);
xnor U22686 (N_22686,N_17605,N_16032);
and U22687 (N_22687,N_16694,N_15387);
nor U22688 (N_22688,N_19906,N_16912);
and U22689 (N_22689,N_17415,N_19116);
and U22690 (N_22690,N_15825,N_16649);
or U22691 (N_22691,N_19584,N_17352);
nand U22692 (N_22692,N_19145,N_15156);
or U22693 (N_22693,N_18005,N_15810);
and U22694 (N_22694,N_16693,N_17470);
nor U22695 (N_22695,N_16025,N_17584);
or U22696 (N_22696,N_19293,N_16095);
nor U22697 (N_22697,N_19878,N_15535);
nor U22698 (N_22698,N_15509,N_18620);
nor U22699 (N_22699,N_18151,N_19196);
nand U22700 (N_22700,N_17286,N_18454);
or U22701 (N_22701,N_15441,N_19769);
xor U22702 (N_22702,N_15729,N_15990);
or U22703 (N_22703,N_18200,N_17569);
or U22704 (N_22704,N_19985,N_15448);
nor U22705 (N_22705,N_18633,N_19513);
xnor U22706 (N_22706,N_16217,N_15512);
or U22707 (N_22707,N_15514,N_18675);
nor U22708 (N_22708,N_16030,N_18406);
and U22709 (N_22709,N_16010,N_18918);
nand U22710 (N_22710,N_18492,N_17929);
or U22711 (N_22711,N_19887,N_15679);
or U22712 (N_22712,N_16249,N_18753);
or U22713 (N_22713,N_17371,N_18615);
and U22714 (N_22714,N_17248,N_17472);
nor U22715 (N_22715,N_15281,N_16738);
nand U22716 (N_22716,N_15858,N_17600);
nand U22717 (N_22717,N_18278,N_19303);
and U22718 (N_22718,N_17014,N_16790);
nand U22719 (N_22719,N_15890,N_19770);
nor U22720 (N_22720,N_15979,N_16442);
nor U22721 (N_22721,N_18996,N_17303);
nand U22722 (N_22722,N_16670,N_18655);
or U22723 (N_22723,N_17209,N_17094);
or U22724 (N_22724,N_16868,N_15761);
nand U22725 (N_22725,N_19755,N_16633);
nand U22726 (N_22726,N_16625,N_16673);
and U22727 (N_22727,N_17329,N_15772);
or U22728 (N_22728,N_19485,N_15122);
nand U22729 (N_22729,N_16131,N_18423);
and U22730 (N_22730,N_18493,N_17552);
xor U22731 (N_22731,N_15429,N_16170);
nor U22732 (N_22732,N_17148,N_17989);
and U22733 (N_22733,N_16538,N_18649);
or U22734 (N_22734,N_19360,N_17323);
and U22735 (N_22735,N_17325,N_15570);
xnor U22736 (N_22736,N_18040,N_17285);
or U22737 (N_22737,N_15767,N_19565);
nand U22738 (N_22738,N_15973,N_19608);
nor U22739 (N_22739,N_17515,N_17657);
nand U22740 (N_22740,N_17763,N_16874);
xnor U22741 (N_22741,N_19105,N_18909);
nor U22742 (N_22742,N_18842,N_16674);
nor U22743 (N_22743,N_17364,N_15178);
xnor U22744 (N_22744,N_17386,N_17726);
nand U22745 (N_22745,N_17446,N_15623);
nor U22746 (N_22746,N_15108,N_17179);
nand U22747 (N_22747,N_15499,N_15309);
or U22748 (N_22748,N_19960,N_15942);
nand U22749 (N_22749,N_16690,N_16753);
or U22750 (N_22750,N_15809,N_17199);
nand U22751 (N_22751,N_18859,N_18289);
nand U22752 (N_22752,N_19947,N_19394);
nand U22753 (N_22753,N_19464,N_19267);
xnor U22754 (N_22754,N_18982,N_18667);
nand U22755 (N_22755,N_18932,N_16709);
xnor U22756 (N_22756,N_18639,N_18464);
and U22757 (N_22757,N_19392,N_19333);
xor U22758 (N_22758,N_18229,N_18182);
nand U22759 (N_22759,N_17315,N_17897);
or U22760 (N_22760,N_18287,N_17417);
nor U22761 (N_22761,N_15770,N_19473);
nor U22762 (N_22762,N_19946,N_16662);
and U22763 (N_22763,N_16454,N_19484);
and U22764 (N_22764,N_15157,N_15086);
nand U22765 (N_22765,N_18983,N_16669);
nor U22766 (N_22766,N_19447,N_19285);
nand U22767 (N_22767,N_15859,N_19227);
xnor U22768 (N_22768,N_16160,N_17881);
xor U22769 (N_22769,N_15081,N_16301);
nand U22770 (N_22770,N_18979,N_17402);
nand U22771 (N_22771,N_15919,N_18728);
nand U22772 (N_22772,N_19467,N_19903);
nor U22773 (N_22773,N_18972,N_16336);
or U22774 (N_22774,N_16024,N_15944);
or U22775 (N_22775,N_18595,N_15912);
xor U22776 (N_22776,N_16826,N_17538);
and U22777 (N_22777,N_18258,N_17217);
xor U22778 (N_22778,N_16598,N_18684);
xnor U22779 (N_22779,N_15757,N_15229);
nand U22780 (N_22780,N_18954,N_19255);
nor U22781 (N_22781,N_19316,N_15868);
or U22782 (N_22782,N_18566,N_16067);
nand U22783 (N_22783,N_18131,N_16662);
nor U22784 (N_22784,N_19955,N_15958);
xnor U22785 (N_22785,N_15337,N_18627);
and U22786 (N_22786,N_15663,N_16346);
nor U22787 (N_22787,N_17511,N_17645);
nand U22788 (N_22788,N_16841,N_19279);
and U22789 (N_22789,N_15855,N_18968);
nand U22790 (N_22790,N_16986,N_16520);
and U22791 (N_22791,N_16132,N_15600);
xor U22792 (N_22792,N_17109,N_15417);
or U22793 (N_22793,N_17282,N_16996);
or U22794 (N_22794,N_17999,N_19789);
or U22795 (N_22795,N_16955,N_17928);
nor U22796 (N_22796,N_19777,N_15847);
or U22797 (N_22797,N_18570,N_18363);
xor U22798 (N_22798,N_17408,N_18546);
nand U22799 (N_22799,N_17863,N_15199);
and U22800 (N_22800,N_18418,N_18104);
xnor U22801 (N_22801,N_19700,N_16871);
nand U22802 (N_22802,N_16852,N_17427);
nor U22803 (N_22803,N_16462,N_15729);
and U22804 (N_22804,N_16009,N_15056);
xnor U22805 (N_22805,N_18169,N_16373);
xor U22806 (N_22806,N_19359,N_15603);
nand U22807 (N_22807,N_17378,N_16997);
or U22808 (N_22808,N_17826,N_19550);
nor U22809 (N_22809,N_19688,N_16197);
or U22810 (N_22810,N_17352,N_18203);
or U22811 (N_22811,N_19776,N_19344);
nor U22812 (N_22812,N_16574,N_18521);
nand U22813 (N_22813,N_19927,N_18517);
and U22814 (N_22814,N_18016,N_16453);
xor U22815 (N_22815,N_16326,N_19321);
nor U22816 (N_22816,N_19689,N_15716);
nor U22817 (N_22817,N_17332,N_17021);
nor U22818 (N_22818,N_18243,N_17053);
nor U22819 (N_22819,N_18626,N_18911);
nand U22820 (N_22820,N_15580,N_19829);
nand U22821 (N_22821,N_17214,N_16776);
xor U22822 (N_22822,N_19383,N_16861);
nand U22823 (N_22823,N_19469,N_19129);
or U22824 (N_22824,N_15299,N_17343);
and U22825 (N_22825,N_18068,N_19142);
nor U22826 (N_22826,N_19027,N_15716);
or U22827 (N_22827,N_16527,N_19652);
nor U22828 (N_22828,N_16700,N_15099);
nand U22829 (N_22829,N_15571,N_17801);
nor U22830 (N_22830,N_16956,N_15344);
and U22831 (N_22831,N_19426,N_17242);
and U22832 (N_22832,N_17992,N_15842);
or U22833 (N_22833,N_15821,N_17061);
nand U22834 (N_22834,N_19399,N_19161);
and U22835 (N_22835,N_19020,N_16865);
or U22836 (N_22836,N_18926,N_16913);
or U22837 (N_22837,N_15639,N_16521);
nor U22838 (N_22838,N_16336,N_18260);
and U22839 (N_22839,N_16360,N_17521);
nor U22840 (N_22840,N_16799,N_19041);
and U22841 (N_22841,N_16068,N_15552);
and U22842 (N_22842,N_17519,N_18687);
or U22843 (N_22843,N_15457,N_19833);
or U22844 (N_22844,N_19223,N_18617);
nand U22845 (N_22845,N_16341,N_16643);
or U22846 (N_22846,N_19886,N_18363);
nand U22847 (N_22847,N_17932,N_17981);
xor U22848 (N_22848,N_17718,N_16718);
nand U22849 (N_22849,N_15262,N_15367);
nand U22850 (N_22850,N_19848,N_17826);
nor U22851 (N_22851,N_16776,N_18299);
nand U22852 (N_22852,N_15325,N_17610);
nor U22853 (N_22853,N_17379,N_17699);
nor U22854 (N_22854,N_16587,N_19030);
xnor U22855 (N_22855,N_17363,N_19518);
xor U22856 (N_22856,N_16374,N_17265);
or U22857 (N_22857,N_16535,N_15645);
or U22858 (N_22858,N_15574,N_17024);
and U22859 (N_22859,N_19332,N_15814);
nand U22860 (N_22860,N_19739,N_17188);
nand U22861 (N_22861,N_17090,N_15170);
xor U22862 (N_22862,N_18717,N_18191);
xor U22863 (N_22863,N_16140,N_19861);
xnor U22864 (N_22864,N_17518,N_17731);
nor U22865 (N_22865,N_19089,N_17980);
xnor U22866 (N_22866,N_16714,N_17609);
nand U22867 (N_22867,N_15036,N_17967);
and U22868 (N_22868,N_15031,N_19396);
and U22869 (N_22869,N_17903,N_17004);
and U22870 (N_22870,N_17343,N_15846);
and U22871 (N_22871,N_16484,N_15561);
or U22872 (N_22872,N_19334,N_15919);
xnor U22873 (N_22873,N_16469,N_15009);
nand U22874 (N_22874,N_18526,N_19692);
or U22875 (N_22875,N_16510,N_18260);
nand U22876 (N_22876,N_15892,N_19925);
nor U22877 (N_22877,N_17541,N_18435);
or U22878 (N_22878,N_17607,N_16154);
and U22879 (N_22879,N_16623,N_18989);
and U22880 (N_22880,N_18656,N_19706);
xor U22881 (N_22881,N_18625,N_16003);
or U22882 (N_22882,N_15956,N_18019);
or U22883 (N_22883,N_17357,N_19129);
xor U22884 (N_22884,N_15011,N_19531);
or U22885 (N_22885,N_19872,N_16380);
nor U22886 (N_22886,N_18992,N_18712);
nand U22887 (N_22887,N_16941,N_16540);
and U22888 (N_22888,N_17051,N_19350);
and U22889 (N_22889,N_19315,N_16414);
nor U22890 (N_22890,N_15253,N_17419);
xnor U22891 (N_22891,N_15005,N_18562);
nand U22892 (N_22892,N_15516,N_19667);
or U22893 (N_22893,N_17031,N_15435);
nor U22894 (N_22894,N_19772,N_19285);
or U22895 (N_22895,N_17610,N_16056);
nor U22896 (N_22896,N_16573,N_15532);
nand U22897 (N_22897,N_15882,N_19676);
or U22898 (N_22898,N_16224,N_18809);
and U22899 (N_22899,N_19748,N_19081);
and U22900 (N_22900,N_17412,N_19258);
xor U22901 (N_22901,N_15866,N_19758);
or U22902 (N_22902,N_18779,N_17474);
xnor U22903 (N_22903,N_16181,N_18757);
or U22904 (N_22904,N_18583,N_18086);
nor U22905 (N_22905,N_19693,N_16737);
nor U22906 (N_22906,N_17387,N_19083);
nor U22907 (N_22907,N_15035,N_19828);
and U22908 (N_22908,N_16046,N_16095);
and U22909 (N_22909,N_19497,N_15181);
nor U22910 (N_22910,N_16618,N_19601);
nand U22911 (N_22911,N_17708,N_19795);
nand U22912 (N_22912,N_18672,N_19063);
and U22913 (N_22913,N_17776,N_15156);
or U22914 (N_22914,N_16053,N_17096);
xor U22915 (N_22915,N_16843,N_15017);
nor U22916 (N_22916,N_16927,N_18741);
nor U22917 (N_22917,N_18186,N_15525);
nand U22918 (N_22918,N_15000,N_17843);
nand U22919 (N_22919,N_16373,N_18235);
nand U22920 (N_22920,N_18996,N_17084);
nor U22921 (N_22921,N_19197,N_18055);
xor U22922 (N_22922,N_18409,N_15700);
and U22923 (N_22923,N_19358,N_15529);
nand U22924 (N_22924,N_16826,N_16503);
xor U22925 (N_22925,N_15701,N_15174);
nand U22926 (N_22926,N_15620,N_17606);
xnor U22927 (N_22927,N_18520,N_19599);
xnor U22928 (N_22928,N_18237,N_19886);
nand U22929 (N_22929,N_18389,N_18264);
nor U22930 (N_22930,N_19959,N_18859);
xor U22931 (N_22931,N_15885,N_16421);
or U22932 (N_22932,N_17907,N_15840);
and U22933 (N_22933,N_15803,N_16386);
nand U22934 (N_22934,N_18356,N_19825);
nand U22935 (N_22935,N_15168,N_17007);
nor U22936 (N_22936,N_16286,N_16554);
nand U22937 (N_22937,N_17002,N_18170);
xnor U22938 (N_22938,N_18593,N_19695);
nor U22939 (N_22939,N_17799,N_16988);
xnor U22940 (N_22940,N_19626,N_15282);
nand U22941 (N_22941,N_17980,N_16606);
nor U22942 (N_22942,N_16426,N_16194);
or U22943 (N_22943,N_18362,N_16693);
nor U22944 (N_22944,N_19326,N_19340);
nand U22945 (N_22945,N_15659,N_15906);
nand U22946 (N_22946,N_17559,N_16944);
nand U22947 (N_22947,N_19299,N_18363);
and U22948 (N_22948,N_18182,N_15376);
nand U22949 (N_22949,N_18726,N_15269);
or U22950 (N_22950,N_15595,N_15763);
and U22951 (N_22951,N_17283,N_18021);
xor U22952 (N_22952,N_16737,N_19567);
or U22953 (N_22953,N_15207,N_16601);
or U22954 (N_22954,N_19761,N_18443);
or U22955 (N_22955,N_16556,N_16117);
xnor U22956 (N_22956,N_15299,N_16675);
xor U22957 (N_22957,N_18044,N_15945);
and U22958 (N_22958,N_16388,N_15316);
nand U22959 (N_22959,N_17635,N_16334);
or U22960 (N_22960,N_19032,N_19211);
nor U22961 (N_22961,N_18582,N_19179);
xnor U22962 (N_22962,N_19185,N_16932);
nand U22963 (N_22963,N_19401,N_19136);
or U22964 (N_22964,N_19265,N_16567);
and U22965 (N_22965,N_15681,N_17749);
and U22966 (N_22966,N_19638,N_18293);
nor U22967 (N_22967,N_19392,N_19436);
xnor U22968 (N_22968,N_15318,N_15564);
nand U22969 (N_22969,N_19484,N_18126);
nand U22970 (N_22970,N_17248,N_15587);
or U22971 (N_22971,N_19561,N_18635);
nor U22972 (N_22972,N_18641,N_17220);
xor U22973 (N_22973,N_17531,N_19794);
nand U22974 (N_22974,N_15303,N_16787);
nand U22975 (N_22975,N_18438,N_18617);
nor U22976 (N_22976,N_18742,N_18676);
nand U22977 (N_22977,N_18847,N_19268);
and U22978 (N_22978,N_16377,N_19455);
nor U22979 (N_22979,N_18155,N_17086);
and U22980 (N_22980,N_18769,N_18423);
nand U22981 (N_22981,N_15553,N_19276);
or U22982 (N_22982,N_15999,N_16880);
nor U22983 (N_22983,N_18938,N_18153);
xnor U22984 (N_22984,N_15701,N_18781);
xor U22985 (N_22985,N_15625,N_17364);
and U22986 (N_22986,N_17567,N_16926);
and U22987 (N_22987,N_18320,N_18225);
or U22988 (N_22988,N_19428,N_16778);
or U22989 (N_22989,N_19259,N_18866);
xor U22990 (N_22990,N_17165,N_17462);
or U22991 (N_22991,N_17267,N_18504);
xnor U22992 (N_22992,N_15121,N_18559);
or U22993 (N_22993,N_16408,N_17320);
nand U22994 (N_22994,N_15156,N_16909);
or U22995 (N_22995,N_19213,N_16998);
and U22996 (N_22996,N_17480,N_17011);
nand U22997 (N_22997,N_19599,N_17900);
xnor U22998 (N_22998,N_15602,N_15684);
nor U22999 (N_22999,N_18327,N_18191);
nor U23000 (N_23000,N_17405,N_16448);
nand U23001 (N_23001,N_19016,N_17101);
nor U23002 (N_23002,N_16373,N_19108);
xnor U23003 (N_23003,N_18092,N_16863);
xor U23004 (N_23004,N_18890,N_16026);
or U23005 (N_23005,N_17998,N_19812);
and U23006 (N_23006,N_19767,N_15599);
nand U23007 (N_23007,N_17434,N_19774);
nand U23008 (N_23008,N_15683,N_19826);
nor U23009 (N_23009,N_15063,N_17542);
and U23010 (N_23010,N_17283,N_16271);
xnor U23011 (N_23011,N_15352,N_18431);
or U23012 (N_23012,N_15208,N_19535);
nor U23013 (N_23013,N_16203,N_15119);
and U23014 (N_23014,N_17169,N_19565);
xnor U23015 (N_23015,N_17752,N_18952);
or U23016 (N_23016,N_19851,N_17485);
nor U23017 (N_23017,N_17052,N_19382);
xnor U23018 (N_23018,N_16230,N_19847);
and U23019 (N_23019,N_15495,N_18847);
and U23020 (N_23020,N_16308,N_15418);
and U23021 (N_23021,N_19376,N_16830);
and U23022 (N_23022,N_19377,N_17904);
and U23023 (N_23023,N_18179,N_15035);
nor U23024 (N_23024,N_19168,N_18165);
or U23025 (N_23025,N_16172,N_16129);
xnor U23026 (N_23026,N_19944,N_19041);
or U23027 (N_23027,N_18647,N_16631);
nand U23028 (N_23028,N_16635,N_15168);
nor U23029 (N_23029,N_17182,N_19982);
nand U23030 (N_23030,N_16912,N_17599);
or U23031 (N_23031,N_18462,N_18650);
nand U23032 (N_23032,N_17196,N_18101);
nor U23033 (N_23033,N_15833,N_18583);
or U23034 (N_23034,N_18116,N_16613);
xor U23035 (N_23035,N_16448,N_17613);
and U23036 (N_23036,N_15983,N_18247);
nor U23037 (N_23037,N_19332,N_19882);
and U23038 (N_23038,N_16813,N_17555);
and U23039 (N_23039,N_17055,N_19291);
nor U23040 (N_23040,N_16603,N_17833);
and U23041 (N_23041,N_17765,N_18040);
and U23042 (N_23042,N_16876,N_18460);
nand U23043 (N_23043,N_19623,N_15372);
xnor U23044 (N_23044,N_17204,N_17684);
nor U23045 (N_23045,N_17946,N_19161);
nor U23046 (N_23046,N_15805,N_16861);
xnor U23047 (N_23047,N_16668,N_16813);
nor U23048 (N_23048,N_16857,N_18457);
nand U23049 (N_23049,N_18564,N_16445);
xnor U23050 (N_23050,N_17493,N_15142);
or U23051 (N_23051,N_17042,N_16229);
xnor U23052 (N_23052,N_16742,N_17548);
xor U23053 (N_23053,N_17774,N_16869);
nor U23054 (N_23054,N_16437,N_18926);
nand U23055 (N_23055,N_15947,N_16029);
or U23056 (N_23056,N_18089,N_17111);
and U23057 (N_23057,N_17280,N_18900);
nand U23058 (N_23058,N_18557,N_15798);
nand U23059 (N_23059,N_16763,N_19159);
nand U23060 (N_23060,N_17117,N_16647);
or U23061 (N_23061,N_17226,N_18575);
and U23062 (N_23062,N_15591,N_17059);
nand U23063 (N_23063,N_15725,N_16178);
xnor U23064 (N_23064,N_16857,N_15198);
nand U23065 (N_23065,N_15482,N_19951);
xnor U23066 (N_23066,N_19571,N_18122);
nor U23067 (N_23067,N_19069,N_15972);
or U23068 (N_23068,N_18728,N_19185);
nor U23069 (N_23069,N_18887,N_17112);
nor U23070 (N_23070,N_18529,N_19798);
nor U23071 (N_23071,N_15245,N_18434);
nand U23072 (N_23072,N_16973,N_17702);
and U23073 (N_23073,N_16340,N_17735);
xnor U23074 (N_23074,N_17640,N_18187);
nor U23075 (N_23075,N_18590,N_17982);
or U23076 (N_23076,N_17400,N_15429);
xnor U23077 (N_23077,N_17813,N_15870);
nor U23078 (N_23078,N_17009,N_19491);
xnor U23079 (N_23079,N_18463,N_15874);
xor U23080 (N_23080,N_15393,N_15381);
nand U23081 (N_23081,N_15790,N_16337);
or U23082 (N_23082,N_16262,N_15627);
nand U23083 (N_23083,N_16617,N_19632);
xor U23084 (N_23084,N_19757,N_17230);
xnor U23085 (N_23085,N_16052,N_16128);
or U23086 (N_23086,N_15798,N_19611);
or U23087 (N_23087,N_19994,N_18098);
nor U23088 (N_23088,N_15699,N_19088);
nand U23089 (N_23089,N_16403,N_15315);
xor U23090 (N_23090,N_16515,N_17505);
xnor U23091 (N_23091,N_17311,N_18373);
and U23092 (N_23092,N_19591,N_19149);
xnor U23093 (N_23093,N_16007,N_18910);
nor U23094 (N_23094,N_16685,N_17640);
xor U23095 (N_23095,N_18472,N_16807);
nor U23096 (N_23096,N_19868,N_16433);
or U23097 (N_23097,N_16495,N_17429);
nor U23098 (N_23098,N_17585,N_15527);
or U23099 (N_23099,N_17431,N_17490);
or U23100 (N_23100,N_16504,N_17752);
or U23101 (N_23101,N_18711,N_19774);
nor U23102 (N_23102,N_19132,N_17036);
nor U23103 (N_23103,N_16550,N_19101);
or U23104 (N_23104,N_15334,N_19948);
nand U23105 (N_23105,N_16273,N_16467);
and U23106 (N_23106,N_19742,N_17409);
and U23107 (N_23107,N_17876,N_15302);
or U23108 (N_23108,N_18658,N_16120);
xnor U23109 (N_23109,N_16675,N_16225);
nor U23110 (N_23110,N_19079,N_19482);
nand U23111 (N_23111,N_16625,N_17299);
or U23112 (N_23112,N_16842,N_18172);
nor U23113 (N_23113,N_19687,N_15162);
nor U23114 (N_23114,N_19414,N_19549);
xor U23115 (N_23115,N_18404,N_19361);
nand U23116 (N_23116,N_15798,N_18040);
xor U23117 (N_23117,N_16855,N_15806);
xor U23118 (N_23118,N_18441,N_19584);
nor U23119 (N_23119,N_17519,N_18675);
and U23120 (N_23120,N_16457,N_19071);
or U23121 (N_23121,N_16604,N_18439);
nand U23122 (N_23122,N_19864,N_17818);
nand U23123 (N_23123,N_17526,N_17922);
xor U23124 (N_23124,N_16420,N_17912);
nor U23125 (N_23125,N_18796,N_15072);
or U23126 (N_23126,N_19448,N_18429);
and U23127 (N_23127,N_19654,N_15507);
nor U23128 (N_23128,N_15347,N_18502);
and U23129 (N_23129,N_15167,N_15617);
or U23130 (N_23130,N_19773,N_16453);
or U23131 (N_23131,N_17362,N_19091);
or U23132 (N_23132,N_19515,N_15771);
or U23133 (N_23133,N_17070,N_17591);
and U23134 (N_23134,N_16696,N_15684);
xnor U23135 (N_23135,N_17122,N_19490);
or U23136 (N_23136,N_16255,N_16589);
or U23137 (N_23137,N_17881,N_18826);
xor U23138 (N_23138,N_19402,N_16814);
xor U23139 (N_23139,N_19115,N_15390);
nor U23140 (N_23140,N_15069,N_19806);
nand U23141 (N_23141,N_16213,N_17885);
nor U23142 (N_23142,N_15805,N_19433);
and U23143 (N_23143,N_18934,N_18945);
xnor U23144 (N_23144,N_17520,N_16308);
or U23145 (N_23145,N_16060,N_19884);
and U23146 (N_23146,N_15493,N_16623);
nor U23147 (N_23147,N_17301,N_16925);
or U23148 (N_23148,N_17905,N_16535);
nor U23149 (N_23149,N_18798,N_15029);
and U23150 (N_23150,N_18047,N_19243);
nor U23151 (N_23151,N_15710,N_15942);
and U23152 (N_23152,N_17754,N_17361);
nor U23153 (N_23153,N_18951,N_16086);
nand U23154 (N_23154,N_15478,N_15686);
and U23155 (N_23155,N_18683,N_16231);
or U23156 (N_23156,N_15631,N_18709);
nor U23157 (N_23157,N_17273,N_18102);
xor U23158 (N_23158,N_16536,N_18152);
or U23159 (N_23159,N_17083,N_19444);
nor U23160 (N_23160,N_18181,N_18764);
or U23161 (N_23161,N_15014,N_19602);
nor U23162 (N_23162,N_17806,N_17945);
nand U23163 (N_23163,N_18176,N_18350);
xnor U23164 (N_23164,N_19094,N_19703);
nor U23165 (N_23165,N_18519,N_15994);
nor U23166 (N_23166,N_19260,N_18623);
nand U23167 (N_23167,N_16075,N_16956);
nor U23168 (N_23168,N_18612,N_17512);
and U23169 (N_23169,N_16598,N_19440);
and U23170 (N_23170,N_17474,N_16790);
nor U23171 (N_23171,N_19679,N_19348);
or U23172 (N_23172,N_19054,N_16651);
and U23173 (N_23173,N_15579,N_19557);
xor U23174 (N_23174,N_16277,N_18110);
or U23175 (N_23175,N_19548,N_15409);
xnor U23176 (N_23176,N_16664,N_17590);
nor U23177 (N_23177,N_18523,N_16901);
or U23178 (N_23178,N_17783,N_17922);
and U23179 (N_23179,N_15380,N_19339);
and U23180 (N_23180,N_17060,N_15446);
nor U23181 (N_23181,N_19395,N_17070);
nor U23182 (N_23182,N_17588,N_19371);
or U23183 (N_23183,N_16763,N_18968);
xnor U23184 (N_23184,N_15649,N_18710);
nand U23185 (N_23185,N_16212,N_17126);
xnor U23186 (N_23186,N_17296,N_15785);
or U23187 (N_23187,N_15509,N_18916);
and U23188 (N_23188,N_18626,N_16434);
nor U23189 (N_23189,N_16765,N_15911);
nand U23190 (N_23190,N_19252,N_18058);
and U23191 (N_23191,N_15974,N_16450);
nor U23192 (N_23192,N_17940,N_18444);
nor U23193 (N_23193,N_17943,N_19618);
nor U23194 (N_23194,N_18462,N_16940);
nand U23195 (N_23195,N_18539,N_18327);
and U23196 (N_23196,N_15387,N_19155);
and U23197 (N_23197,N_17264,N_16715);
nand U23198 (N_23198,N_17779,N_18978);
xnor U23199 (N_23199,N_15161,N_16879);
and U23200 (N_23200,N_18986,N_17712);
nand U23201 (N_23201,N_16797,N_15935);
nand U23202 (N_23202,N_17196,N_16470);
nand U23203 (N_23203,N_19731,N_18858);
nor U23204 (N_23204,N_15658,N_17086);
and U23205 (N_23205,N_17625,N_15308);
or U23206 (N_23206,N_16994,N_16300);
and U23207 (N_23207,N_18150,N_16917);
or U23208 (N_23208,N_16676,N_16533);
xnor U23209 (N_23209,N_17200,N_15393);
xnor U23210 (N_23210,N_17120,N_19442);
and U23211 (N_23211,N_16249,N_19309);
nor U23212 (N_23212,N_18358,N_16478);
nand U23213 (N_23213,N_17763,N_17596);
and U23214 (N_23214,N_17751,N_15279);
nor U23215 (N_23215,N_19710,N_16150);
nand U23216 (N_23216,N_18885,N_15187);
xnor U23217 (N_23217,N_16683,N_18234);
nor U23218 (N_23218,N_17123,N_18714);
xor U23219 (N_23219,N_19241,N_17024);
nand U23220 (N_23220,N_18844,N_17010);
and U23221 (N_23221,N_17566,N_19689);
or U23222 (N_23222,N_16891,N_15495);
or U23223 (N_23223,N_16108,N_19108);
nand U23224 (N_23224,N_16317,N_19755);
and U23225 (N_23225,N_17303,N_16660);
xnor U23226 (N_23226,N_17019,N_15640);
nand U23227 (N_23227,N_18035,N_17210);
and U23228 (N_23228,N_16508,N_18334);
and U23229 (N_23229,N_16374,N_18423);
nor U23230 (N_23230,N_15971,N_18532);
or U23231 (N_23231,N_19188,N_19907);
xor U23232 (N_23232,N_19399,N_15805);
and U23233 (N_23233,N_19122,N_19608);
nor U23234 (N_23234,N_16358,N_18305);
xor U23235 (N_23235,N_16319,N_19364);
nand U23236 (N_23236,N_17315,N_16641);
and U23237 (N_23237,N_18791,N_15972);
nor U23238 (N_23238,N_17486,N_17359);
xor U23239 (N_23239,N_16026,N_17530);
nand U23240 (N_23240,N_15985,N_18416);
and U23241 (N_23241,N_15803,N_17250);
nor U23242 (N_23242,N_17988,N_16659);
xor U23243 (N_23243,N_15509,N_19920);
nand U23244 (N_23244,N_15556,N_19420);
xor U23245 (N_23245,N_15113,N_16051);
xnor U23246 (N_23246,N_18318,N_17900);
nand U23247 (N_23247,N_17701,N_16571);
nand U23248 (N_23248,N_15839,N_19583);
or U23249 (N_23249,N_17513,N_17168);
nand U23250 (N_23250,N_19573,N_18319);
xnor U23251 (N_23251,N_15411,N_15849);
xnor U23252 (N_23252,N_16736,N_18378);
nand U23253 (N_23253,N_18463,N_19605);
nor U23254 (N_23254,N_16159,N_16505);
xnor U23255 (N_23255,N_15285,N_19920);
and U23256 (N_23256,N_19292,N_17787);
nor U23257 (N_23257,N_17504,N_16592);
xnor U23258 (N_23258,N_17283,N_16769);
nand U23259 (N_23259,N_19740,N_16287);
nand U23260 (N_23260,N_15680,N_16161);
xor U23261 (N_23261,N_19132,N_17562);
xor U23262 (N_23262,N_18284,N_18663);
nand U23263 (N_23263,N_15884,N_19528);
xor U23264 (N_23264,N_19789,N_15689);
nand U23265 (N_23265,N_19537,N_15841);
and U23266 (N_23266,N_18283,N_17212);
nor U23267 (N_23267,N_15197,N_19754);
xnor U23268 (N_23268,N_18285,N_16424);
nand U23269 (N_23269,N_19146,N_16003);
nor U23270 (N_23270,N_19042,N_19421);
nor U23271 (N_23271,N_18877,N_19881);
nor U23272 (N_23272,N_18442,N_19841);
xnor U23273 (N_23273,N_19950,N_18322);
or U23274 (N_23274,N_19068,N_17201);
or U23275 (N_23275,N_18898,N_17022);
or U23276 (N_23276,N_16238,N_15861);
and U23277 (N_23277,N_19215,N_17524);
and U23278 (N_23278,N_15380,N_17796);
or U23279 (N_23279,N_18296,N_18675);
xor U23280 (N_23280,N_16674,N_15361);
nor U23281 (N_23281,N_16652,N_15281);
nand U23282 (N_23282,N_19817,N_17979);
nor U23283 (N_23283,N_19499,N_15384);
nand U23284 (N_23284,N_17258,N_17200);
nand U23285 (N_23285,N_15037,N_16868);
or U23286 (N_23286,N_18509,N_19374);
or U23287 (N_23287,N_15469,N_17168);
or U23288 (N_23288,N_18346,N_15547);
xnor U23289 (N_23289,N_16891,N_19948);
and U23290 (N_23290,N_18660,N_16248);
xor U23291 (N_23291,N_16051,N_16514);
nor U23292 (N_23292,N_19864,N_18601);
and U23293 (N_23293,N_18313,N_17505);
nor U23294 (N_23294,N_18540,N_15125);
or U23295 (N_23295,N_15370,N_19629);
nor U23296 (N_23296,N_16927,N_19952);
and U23297 (N_23297,N_15704,N_17789);
nor U23298 (N_23298,N_16376,N_19508);
xor U23299 (N_23299,N_18993,N_19271);
or U23300 (N_23300,N_19712,N_18813);
or U23301 (N_23301,N_17161,N_15464);
and U23302 (N_23302,N_17335,N_15635);
and U23303 (N_23303,N_16946,N_18600);
nand U23304 (N_23304,N_17686,N_15587);
and U23305 (N_23305,N_15754,N_18250);
and U23306 (N_23306,N_19265,N_19715);
nor U23307 (N_23307,N_18905,N_15009);
or U23308 (N_23308,N_17552,N_16559);
nor U23309 (N_23309,N_19885,N_18340);
xor U23310 (N_23310,N_19507,N_16094);
nand U23311 (N_23311,N_16857,N_15520);
xnor U23312 (N_23312,N_16331,N_15535);
or U23313 (N_23313,N_18356,N_19013);
or U23314 (N_23314,N_19721,N_17656);
nand U23315 (N_23315,N_18719,N_19234);
nand U23316 (N_23316,N_19165,N_15656);
nand U23317 (N_23317,N_19014,N_17612);
nor U23318 (N_23318,N_18557,N_15999);
nor U23319 (N_23319,N_17029,N_18023);
and U23320 (N_23320,N_15572,N_16833);
or U23321 (N_23321,N_17930,N_16847);
or U23322 (N_23322,N_19947,N_15866);
and U23323 (N_23323,N_15491,N_18293);
nand U23324 (N_23324,N_16951,N_15562);
or U23325 (N_23325,N_17547,N_15734);
xnor U23326 (N_23326,N_19454,N_19536);
nor U23327 (N_23327,N_17417,N_19130);
xor U23328 (N_23328,N_19120,N_19129);
nor U23329 (N_23329,N_16864,N_16749);
nand U23330 (N_23330,N_17739,N_19812);
nor U23331 (N_23331,N_17319,N_19364);
nand U23332 (N_23332,N_19270,N_18470);
nand U23333 (N_23333,N_15693,N_17583);
xnor U23334 (N_23334,N_19038,N_17221);
and U23335 (N_23335,N_17403,N_18410);
and U23336 (N_23336,N_18608,N_17634);
nor U23337 (N_23337,N_16777,N_15585);
and U23338 (N_23338,N_15279,N_18586);
and U23339 (N_23339,N_16836,N_16202);
and U23340 (N_23340,N_16522,N_15317);
or U23341 (N_23341,N_17554,N_16012);
xor U23342 (N_23342,N_15853,N_16971);
xnor U23343 (N_23343,N_19456,N_15912);
or U23344 (N_23344,N_18846,N_15506);
or U23345 (N_23345,N_18573,N_18529);
and U23346 (N_23346,N_19914,N_18281);
and U23347 (N_23347,N_19279,N_18754);
or U23348 (N_23348,N_19489,N_15133);
and U23349 (N_23349,N_16757,N_18954);
nor U23350 (N_23350,N_17086,N_15821);
xnor U23351 (N_23351,N_17979,N_18209);
nand U23352 (N_23352,N_17024,N_18777);
nand U23353 (N_23353,N_19597,N_17944);
or U23354 (N_23354,N_16933,N_16143);
nand U23355 (N_23355,N_17044,N_18586);
xor U23356 (N_23356,N_15569,N_17027);
or U23357 (N_23357,N_18349,N_18134);
and U23358 (N_23358,N_18575,N_19292);
or U23359 (N_23359,N_17516,N_19189);
or U23360 (N_23360,N_18595,N_19068);
nand U23361 (N_23361,N_16736,N_15530);
nand U23362 (N_23362,N_15117,N_15893);
or U23363 (N_23363,N_18326,N_18564);
nor U23364 (N_23364,N_18297,N_19258);
nor U23365 (N_23365,N_19491,N_17868);
and U23366 (N_23366,N_16596,N_17990);
nand U23367 (N_23367,N_16643,N_17844);
or U23368 (N_23368,N_16556,N_17736);
nor U23369 (N_23369,N_19397,N_18424);
nor U23370 (N_23370,N_15484,N_19523);
nor U23371 (N_23371,N_17532,N_15128);
or U23372 (N_23372,N_15270,N_19682);
xnor U23373 (N_23373,N_19503,N_16613);
nor U23374 (N_23374,N_18638,N_17244);
nor U23375 (N_23375,N_17857,N_16977);
nor U23376 (N_23376,N_19517,N_15329);
nand U23377 (N_23377,N_16348,N_19042);
nor U23378 (N_23378,N_18719,N_17939);
nand U23379 (N_23379,N_18698,N_17043);
nand U23380 (N_23380,N_18974,N_15747);
nor U23381 (N_23381,N_15839,N_18763);
or U23382 (N_23382,N_18335,N_19512);
or U23383 (N_23383,N_16041,N_18599);
nand U23384 (N_23384,N_16825,N_17182);
nor U23385 (N_23385,N_15547,N_19719);
and U23386 (N_23386,N_17109,N_19426);
xor U23387 (N_23387,N_15194,N_18177);
xnor U23388 (N_23388,N_19837,N_18505);
nand U23389 (N_23389,N_16560,N_19180);
xnor U23390 (N_23390,N_16988,N_17746);
nor U23391 (N_23391,N_18329,N_17338);
and U23392 (N_23392,N_16137,N_15427);
and U23393 (N_23393,N_19637,N_17547);
or U23394 (N_23394,N_15176,N_17427);
and U23395 (N_23395,N_17512,N_16961);
or U23396 (N_23396,N_15360,N_19553);
xnor U23397 (N_23397,N_18551,N_19509);
xnor U23398 (N_23398,N_15636,N_19713);
nand U23399 (N_23399,N_19824,N_17414);
nor U23400 (N_23400,N_19996,N_15327);
nor U23401 (N_23401,N_19669,N_18085);
nand U23402 (N_23402,N_15521,N_16074);
nand U23403 (N_23403,N_19279,N_17266);
nand U23404 (N_23404,N_19370,N_16011);
or U23405 (N_23405,N_16238,N_18256);
nor U23406 (N_23406,N_16069,N_18309);
nand U23407 (N_23407,N_18247,N_15314);
nor U23408 (N_23408,N_18516,N_19833);
and U23409 (N_23409,N_16562,N_16924);
nor U23410 (N_23410,N_15553,N_15454);
xnor U23411 (N_23411,N_17832,N_17688);
nor U23412 (N_23412,N_16896,N_19182);
xor U23413 (N_23413,N_16402,N_15177);
and U23414 (N_23414,N_19952,N_17363);
and U23415 (N_23415,N_15383,N_16026);
nand U23416 (N_23416,N_15092,N_19902);
or U23417 (N_23417,N_17920,N_17369);
nor U23418 (N_23418,N_15739,N_15890);
nor U23419 (N_23419,N_19313,N_16527);
xor U23420 (N_23420,N_18800,N_19688);
nand U23421 (N_23421,N_16946,N_17660);
xnor U23422 (N_23422,N_16017,N_15953);
xor U23423 (N_23423,N_15437,N_19572);
nor U23424 (N_23424,N_16963,N_16731);
or U23425 (N_23425,N_18514,N_15326);
nand U23426 (N_23426,N_17970,N_17417);
nand U23427 (N_23427,N_18175,N_18411);
and U23428 (N_23428,N_19666,N_17669);
nor U23429 (N_23429,N_16958,N_16758);
nor U23430 (N_23430,N_16474,N_17397);
xor U23431 (N_23431,N_17078,N_17113);
xor U23432 (N_23432,N_19937,N_17369);
and U23433 (N_23433,N_19716,N_17672);
nand U23434 (N_23434,N_16581,N_15541);
nor U23435 (N_23435,N_15536,N_18244);
and U23436 (N_23436,N_19751,N_18879);
xor U23437 (N_23437,N_18999,N_19895);
nand U23438 (N_23438,N_17568,N_15774);
xor U23439 (N_23439,N_18939,N_15323);
and U23440 (N_23440,N_18863,N_17320);
nor U23441 (N_23441,N_17020,N_15834);
xor U23442 (N_23442,N_18603,N_17581);
nor U23443 (N_23443,N_17021,N_16085);
and U23444 (N_23444,N_15414,N_16889);
or U23445 (N_23445,N_17588,N_15216);
xnor U23446 (N_23446,N_16265,N_16637);
xnor U23447 (N_23447,N_19358,N_16280);
nor U23448 (N_23448,N_16184,N_18645);
nand U23449 (N_23449,N_18071,N_18297);
and U23450 (N_23450,N_15762,N_15452);
xnor U23451 (N_23451,N_16195,N_19196);
nor U23452 (N_23452,N_17932,N_16181);
nand U23453 (N_23453,N_18732,N_18133);
or U23454 (N_23454,N_17953,N_15442);
or U23455 (N_23455,N_15335,N_15179);
nand U23456 (N_23456,N_19488,N_17691);
or U23457 (N_23457,N_17565,N_16145);
and U23458 (N_23458,N_19531,N_16875);
xnor U23459 (N_23459,N_18501,N_16722);
nor U23460 (N_23460,N_15865,N_15795);
nor U23461 (N_23461,N_16216,N_18377);
xor U23462 (N_23462,N_19047,N_17790);
or U23463 (N_23463,N_15288,N_16950);
and U23464 (N_23464,N_15462,N_15950);
nand U23465 (N_23465,N_17668,N_16885);
xor U23466 (N_23466,N_17323,N_16549);
nand U23467 (N_23467,N_19932,N_15291);
nand U23468 (N_23468,N_17192,N_18293);
nor U23469 (N_23469,N_19827,N_15567);
nor U23470 (N_23470,N_18576,N_18396);
nor U23471 (N_23471,N_17370,N_17427);
nand U23472 (N_23472,N_15976,N_16836);
and U23473 (N_23473,N_18267,N_19717);
nand U23474 (N_23474,N_15169,N_19494);
and U23475 (N_23475,N_17369,N_16855);
nand U23476 (N_23476,N_17514,N_15011);
nor U23477 (N_23477,N_16631,N_17751);
xor U23478 (N_23478,N_18183,N_18734);
nor U23479 (N_23479,N_19889,N_16410);
and U23480 (N_23480,N_15318,N_17470);
and U23481 (N_23481,N_16707,N_16518);
nor U23482 (N_23482,N_16699,N_19164);
and U23483 (N_23483,N_16449,N_15131);
or U23484 (N_23484,N_18231,N_19519);
nand U23485 (N_23485,N_19153,N_16468);
nor U23486 (N_23486,N_19289,N_18218);
xnor U23487 (N_23487,N_17434,N_19776);
and U23488 (N_23488,N_19950,N_17835);
nand U23489 (N_23489,N_16318,N_15688);
or U23490 (N_23490,N_19164,N_19725);
or U23491 (N_23491,N_15794,N_16333);
nor U23492 (N_23492,N_17111,N_15339);
xnor U23493 (N_23493,N_18973,N_19414);
nor U23494 (N_23494,N_18858,N_18974);
and U23495 (N_23495,N_15932,N_19286);
and U23496 (N_23496,N_19036,N_17130);
nor U23497 (N_23497,N_19240,N_17173);
xor U23498 (N_23498,N_17237,N_17036);
nor U23499 (N_23499,N_15009,N_15510);
or U23500 (N_23500,N_15786,N_17215);
nand U23501 (N_23501,N_16985,N_17318);
nand U23502 (N_23502,N_16868,N_15771);
nor U23503 (N_23503,N_17898,N_15337);
and U23504 (N_23504,N_18066,N_15706);
xor U23505 (N_23505,N_18980,N_17626);
xor U23506 (N_23506,N_16053,N_19563);
nand U23507 (N_23507,N_17565,N_17572);
nor U23508 (N_23508,N_17105,N_18684);
or U23509 (N_23509,N_16264,N_17555);
and U23510 (N_23510,N_19849,N_15350);
or U23511 (N_23511,N_19949,N_18566);
xnor U23512 (N_23512,N_17867,N_16675);
or U23513 (N_23513,N_19901,N_15301);
nor U23514 (N_23514,N_18795,N_19251);
or U23515 (N_23515,N_18554,N_16473);
xnor U23516 (N_23516,N_17720,N_18688);
or U23517 (N_23517,N_19006,N_15989);
and U23518 (N_23518,N_19485,N_15332);
nand U23519 (N_23519,N_16602,N_15704);
or U23520 (N_23520,N_19899,N_18810);
xor U23521 (N_23521,N_16420,N_19949);
nand U23522 (N_23522,N_18917,N_17335);
nor U23523 (N_23523,N_15056,N_19806);
nor U23524 (N_23524,N_16961,N_15915);
nand U23525 (N_23525,N_19179,N_15373);
xor U23526 (N_23526,N_18736,N_18329);
xnor U23527 (N_23527,N_16268,N_17645);
and U23528 (N_23528,N_17998,N_18133);
and U23529 (N_23529,N_19439,N_17352);
nor U23530 (N_23530,N_17180,N_18889);
and U23531 (N_23531,N_16755,N_16361);
nand U23532 (N_23532,N_19393,N_16631);
or U23533 (N_23533,N_16223,N_15160);
nor U23534 (N_23534,N_18132,N_16463);
or U23535 (N_23535,N_15334,N_19265);
nand U23536 (N_23536,N_15439,N_16087);
nand U23537 (N_23537,N_15873,N_15906);
or U23538 (N_23538,N_15071,N_16982);
nor U23539 (N_23539,N_18299,N_16190);
nand U23540 (N_23540,N_15405,N_16883);
nor U23541 (N_23541,N_16524,N_16614);
nor U23542 (N_23542,N_18366,N_15444);
xnor U23543 (N_23543,N_15085,N_18924);
or U23544 (N_23544,N_17585,N_15641);
or U23545 (N_23545,N_16130,N_18704);
nor U23546 (N_23546,N_19521,N_18023);
nand U23547 (N_23547,N_18335,N_16735);
xnor U23548 (N_23548,N_17005,N_16946);
and U23549 (N_23549,N_19070,N_19356);
nand U23550 (N_23550,N_17026,N_19613);
xnor U23551 (N_23551,N_15065,N_18876);
xor U23552 (N_23552,N_17005,N_17593);
or U23553 (N_23553,N_19428,N_19787);
and U23554 (N_23554,N_16053,N_19120);
or U23555 (N_23555,N_16581,N_15555);
nand U23556 (N_23556,N_15105,N_17359);
and U23557 (N_23557,N_16795,N_17175);
xor U23558 (N_23558,N_17103,N_18048);
or U23559 (N_23559,N_18586,N_19958);
nand U23560 (N_23560,N_16830,N_15289);
nand U23561 (N_23561,N_19918,N_16803);
or U23562 (N_23562,N_16849,N_17232);
or U23563 (N_23563,N_15082,N_19136);
and U23564 (N_23564,N_18655,N_19177);
and U23565 (N_23565,N_16086,N_19077);
nor U23566 (N_23566,N_19092,N_17172);
or U23567 (N_23567,N_16783,N_18003);
and U23568 (N_23568,N_17096,N_18936);
and U23569 (N_23569,N_15492,N_15420);
or U23570 (N_23570,N_19088,N_15184);
xnor U23571 (N_23571,N_17706,N_18295);
nor U23572 (N_23572,N_17257,N_16461);
or U23573 (N_23573,N_15089,N_19641);
xor U23574 (N_23574,N_17766,N_16444);
nor U23575 (N_23575,N_15495,N_17864);
nand U23576 (N_23576,N_18977,N_17249);
xnor U23577 (N_23577,N_17312,N_17838);
xnor U23578 (N_23578,N_19619,N_16070);
xor U23579 (N_23579,N_15758,N_15071);
nand U23580 (N_23580,N_19924,N_17333);
nand U23581 (N_23581,N_19157,N_15509);
nand U23582 (N_23582,N_18148,N_16018);
or U23583 (N_23583,N_16671,N_18282);
or U23584 (N_23584,N_17644,N_18149);
or U23585 (N_23585,N_19660,N_19771);
nor U23586 (N_23586,N_16614,N_16781);
xor U23587 (N_23587,N_18084,N_18376);
and U23588 (N_23588,N_19851,N_15513);
nor U23589 (N_23589,N_16954,N_15941);
and U23590 (N_23590,N_16773,N_17194);
xor U23591 (N_23591,N_16114,N_16735);
and U23592 (N_23592,N_18950,N_19739);
nand U23593 (N_23593,N_18923,N_17640);
nand U23594 (N_23594,N_17322,N_19052);
xor U23595 (N_23595,N_16785,N_18335);
and U23596 (N_23596,N_18432,N_15433);
nand U23597 (N_23597,N_19115,N_16117);
and U23598 (N_23598,N_18720,N_18703);
nand U23599 (N_23599,N_17806,N_18099);
or U23600 (N_23600,N_18383,N_19369);
or U23601 (N_23601,N_17980,N_16259);
and U23602 (N_23602,N_16702,N_19730);
or U23603 (N_23603,N_18742,N_15882);
nor U23604 (N_23604,N_15671,N_15641);
nor U23605 (N_23605,N_17687,N_16116);
nand U23606 (N_23606,N_19575,N_19996);
nand U23607 (N_23607,N_16817,N_17848);
nand U23608 (N_23608,N_18483,N_17389);
nand U23609 (N_23609,N_15829,N_16270);
and U23610 (N_23610,N_17513,N_16517);
xor U23611 (N_23611,N_15506,N_16289);
or U23612 (N_23612,N_18652,N_15356);
nand U23613 (N_23613,N_19705,N_17160);
nor U23614 (N_23614,N_15317,N_18025);
nand U23615 (N_23615,N_15288,N_18614);
and U23616 (N_23616,N_18545,N_17353);
nor U23617 (N_23617,N_15574,N_17793);
xnor U23618 (N_23618,N_17786,N_18558);
nand U23619 (N_23619,N_18756,N_15626);
xor U23620 (N_23620,N_15522,N_18831);
xnor U23621 (N_23621,N_17204,N_15106);
and U23622 (N_23622,N_16828,N_16797);
and U23623 (N_23623,N_15793,N_17863);
nand U23624 (N_23624,N_19904,N_16502);
nor U23625 (N_23625,N_19539,N_15578);
or U23626 (N_23626,N_17210,N_18999);
xor U23627 (N_23627,N_15451,N_19210);
or U23628 (N_23628,N_17242,N_17364);
xnor U23629 (N_23629,N_18228,N_17164);
xor U23630 (N_23630,N_17034,N_18923);
or U23631 (N_23631,N_18294,N_19909);
nand U23632 (N_23632,N_15769,N_15902);
xnor U23633 (N_23633,N_19348,N_18141);
or U23634 (N_23634,N_19594,N_17008);
or U23635 (N_23635,N_16092,N_17368);
or U23636 (N_23636,N_16581,N_19758);
nand U23637 (N_23637,N_16998,N_17954);
nor U23638 (N_23638,N_16657,N_18913);
xor U23639 (N_23639,N_16657,N_15273);
nor U23640 (N_23640,N_19175,N_19208);
nand U23641 (N_23641,N_16288,N_17102);
xor U23642 (N_23642,N_18800,N_18657);
and U23643 (N_23643,N_17133,N_18837);
nand U23644 (N_23644,N_16148,N_16859);
or U23645 (N_23645,N_19370,N_17946);
nor U23646 (N_23646,N_16332,N_17364);
nand U23647 (N_23647,N_17137,N_17187);
nor U23648 (N_23648,N_18471,N_19586);
xor U23649 (N_23649,N_18928,N_17265);
nor U23650 (N_23650,N_18671,N_17807);
or U23651 (N_23651,N_16798,N_19625);
and U23652 (N_23652,N_19205,N_19106);
nor U23653 (N_23653,N_16033,N_17223);
nand U23654 (N_23654,N_16711,N_18905);
nand U23655 (N_23655,N_15178,N_18984);
nor U23656 (N_23656,N_17016,N_17713);
and U23657 (N_23657,N_16624,N_19622);
or U23658 (N_23658,N_17552,N_15571);
xor U23659 (N_23659,N_18082,N_16446);
and U23660 (N_23660,N_18195,N_15178);
or U23661 (N_23661,N_19819,N_18800);
xnor U23662 (N_23662,N_18871,N_15856);
and U23663 (N_23663,N_16156,N_16039);
nor U23664 (N_23664,N_17215,N_17341);
or U23665 (N_23665,N_16049,N_19061);
nor U23666 (N_23666,N_17638,N_15901);
nor U23667 (N_23667,N_17122,N_19942);
nand U23668 (N_23668,N_16749,N_16209);
nor U23669 (N_23669,N_16895,N_18151);
nand U23670 (N_23670,N_17074,N_19086);
or U23671 (N_23671,N_17882,N_15138);
nor U23672 (N_23672,N_19681,N_19891);
and U23673 (N_23673,N_17346,N_15578);
or U23674 (N_23674,N_17024,N_19161);
or U23675 (N_23675,N_18832,N_16046);
nor U23676 (N_23676,N_19014,N_19681);
nand U23677 (N_23677,N_15020,N_17669);
or U23678 (N_23678,N_15928,N_15585);
and U23679 (N_23679,N_15606,N_15255);
xor U23680 (N_23680,N_17938,N_19119);
or U23681 (N_23681,N_19641,N_18683);
and U23682 (N_23682,N_19131,N_16346);
xnor U23683 (N_23683,N_15558,N_15176);
nor U23684 (N_23684,N_15778,N_18390);
nand U23685 (N_23685,N_17687,N_16055);
and U23686 (N_23686,N_18444,N_16182);
nand U23687 (N_23687,N_17141,N_19610);
or U23688 (N_23688,N_16494,N_15306);
nand U23689 (N_23689,N_16185,N_17639);
or U23690 (N_23690,N_16082,N_15181);
nor U23691 (N_23691,N_15945,N_15050);
and U23692 (N_23692,N_17789,N_19234);
and U23693 (N_23693,N_17610,N_18340);
nor U23694 (N_23694,N_15915,N_16630);
nand U23695 (N_23695,N_19147,N_18561);
and U23696 (N_23696,N_17834,N_15699);
nand U23697 (N_23697,N_17170,N_16034);
or U23698 (N_23698,N_17982,N_15887);
nor U23699 (N_23699,N_16922,N_15911);
xnor U23700 (N_23700,N_19115,N_16051);
or U23701 (N_23701,N_18098,N_17692);
nor U23702 (N_23702,N_18744,N_17896);
or U23703 (N_23703,N_16823,N_19719);
nand U23704 (N_23704,N_16414,N_17142);
and U23705 (N_23705,N_17815,N_15909);
nand U23706 (N_23706,N_19455,N_19052);
nand U23707 (N_23707,N_19438,N_15022);
or U23708 (N_23708,N_17761,N_16589);
and U23709 (N_23709,N_16965,N_18641);
or U23710 (N_23710,N_17611,N_17077);
or U23711 (N_23711,N_15251,N_19379);
and U23712 (N_23712,N_15504,N_16658);
or U23713 (N_23713,N_15518,N_18040);
or U23714 (N_23714,N_18512,N_16136);
nor U23715 (N_23715,N_18400,N_18684);
and U23716 (N_23716,N_17633,N_17026);
or U23717 (N_23717,N_19705,N_18747);
and U23718 (N_23718,N_17200,N_19514);
nor U23719 (N_23719,N_16177,N_18149);
nand U23720 (N_23720,N_15394,N_17311);
xnor U23721 (N_23721,N_16769,N_16499);
or U23722 (N_23722,N_17337,N_17410);
or U23723 (N_23723,N_19241,N_19640);
or U23724 (N_23724,N_18133,N_17211);
nand U23725 (N_23725,N_19679,N_17849);
nand U23726 (N_23726,N_16874,N_19880);
nand U23727 (N_23727,N_19336,N_15539);
and U23728 (N_23728,N_16759,N_18402);
xnor U23729 (N_23729,N_17799,N_18945);
or U23730 (N_23730,N_15731,N_15128);
xnor U23731 (N_23731,N_18814,N_18953);
or U23732 (N_23732,N_16686,N_17450);
xor U23733 (N_23733,N_16226,N_18390);
or U23734 (N_23734,N_18820,N_18622);
or U23735 (N_23735,N_17631,N_15423);
nor U23736 (N_23736,N_18037,N_16050);
or U23737 (N_23737,N_18038,N_19118);
xnor U23738 (N_23738,N_15647,N_19277);
and U23739 (N_23739,N_19405,N_17361);
or U23740 (N_23740,N_15830,N_17130);
or U23741 (N_23741,N_15222,N_18197);
and U23742 (N_23742,N_17703,N_19934);
nor U23743 (N_23743,N_18675,N_19824);
xnor U23744 (N_23744,N_17187,N_19949);
and U23745 (N_23745,N_19382,N_19826);
nand U23746 (N_23746,N_19512,N_15481);
or U23747 (N_23747,N_16435,N_17028);
xor U23748 (N_23748,N_18921,N_15784);
xnor U23749 (N_23749,N_18226,N_16351);
and U23750 (N_23750,N_16162,N_15095);
nor U23751 (N_23751,N_19423,N_16903);
nand U23752 (N_23752,N_18093,N_19681);
xor U23753 (N_23753,N_18060,N_15794);
or U23754 (N_23754,N_18886,N_16097);
xnor U23755 (N_23755,N_18431,N_16683);
and U23756 (N_23756,N_19591,N_16280);
nor U23757 (N_23757,N_15956,N_17606);
xor U23758 (N_23758,N_19731,N_18113);
nor U23759 (N_23759,N_15043,N_15703);
or U23760 (N_23760,N_18202,N_15872);
and U23761 (N_23761,N_19514,N_16689);
and U23762 (N_23762,N_19929,N_17984);
and U23763 (N_23763,N_18773,N_19052);
or U23764 (N_23764,N_16976,N_19103);
and U23765 (N_23765,N_17891,N_17873);
xor U23766 (N_23766,N_18574,N_19799);
and U23767 (N_23767,N_16831,N_19037);
or U23768 (N_23768,N_16736,N_17885);
xor U23769 (N_23769,N_17963,N_18631);
or U23770 (N_23770,N_16243,N_16591);
or U23771 (N_23771,N_16943,N_16925);
and U23772 (N_23772,N_17467,N_18528);
nor U23773 (N_23773,N_18038,N_19939);
and U23774 (N_23774,N_15924,N_18541);
xor U23775 (N_23775,N_16166,N_16957);
and U23776 (N_23776,N_19528,N_17394);
nand U23777 (N_23777,N_19057,N_16905);
xor U23778 (N_23778,N_16127,N_16345);
nand U23779 (N_23779,N_15674,N_16798);
nand U23780 (N_23780,N_19304,N_18901);
and U23781 (N_23781,N_17669,N_19789);
nor U23782 (N_23782,N_16068,N_18290);
and U23783 (N_23783,N_15439,N_15318);
nand U23784 (N_23784,N_18146,N_17075);
and U23785 (N_23785,N_19424,N_16249);
or U23786 (N_23786,N_18747,N_18691);
or U23787 (N_23787,N_17215,N_15216);
nor U23788 (N_23788,N_16024,N_19582);
nand U23789 (N_23789,N_16699,N_16917);
xor U23790 (N_23790,N_19979,N_15892);
nand U23791 (N_23791,N_15872,N_18554);
or U23792 (N_23792,N_15623,N_17406);
xor U23793 (N_23793,N_18848,N_19467);
nor U23794 (N_23794,N_16977,N_15262);
nand U23795 (N_23795,N_19239,N_16172);
or U23796 (N_23796,N_19135,N_18894);
and U23797 (N_23797,N_17424,N_19864);
nor U23798 (N_23798,N_16613,N_18441);
or U23799 (N_23799,N_17225,N_19042);
or U23800 (N_23800,N_18738,N_16218);
xor U23801 (N_23801,N_19033,N_17389);
nor U23802 (N_23802,N_19627,N_17348);
xnor U23803 (N_23803,N_18309,N_19668);
nand U23804 (N_23804,N_17388,N_19177);
or U23805 (N_23805,N_17384,N_17638);
or U23806 (N_23806,N_19627,N_16610);
xnor U23807 (N_23807,N_18805,N_15083);
nor U23808 (N_23808,N_19715,N_19694);
nand U23809 (N_23809,N_16750,N_15100);
xor U23810 (N_23810,N_18138,N_15720);
xor U23811 (N_23811,N_19848,N_17356);
or U23812 (N_23812,N_16418,N_15263);
nand U23813 (N_23813,N_19778,N_18278);
xnor U23814 (N_23814,N_17114,N_15566);
and U23815 (N_23815,N_15141,N_19240);
xnor U23816 (N_23816,N_16681,N_17751);
and U23817 (N_23817,N_19751,N_18209);
and U23818 (N_23818,N_18040,N_18277);
and U23819 (N_23819,N_17647,N_17399);
nand U23820 (N_23820,N_18974,N_17104);
or U23821 (N_23821,N_17881,N_18447);
or U23822 (N_23822,N_17411,N_17634);
or U23823 (N_23823,N_18820,N_18524);
nand U23824 (N_23824,N_17047,N_15008);
or U23825 (N_23825,N_16085,N_16015);
and U23826 (N_23826,N_17273,N_18679);
nand U23827 (N_23827,N_17954,N_16649);
nor U23828 (N_23828,N_16616,N_17573);
xor U23829 (N_23829,N_15960,N_18553);
and U23830 (N_23830,N_16521,N_15367);
nor U23831 (N_23831,N_15877,N_15058);
and U23832 (N_23832,N_18512,N_17181);
nand U23833 (N_23833,N_18341,N_15970);
and U23834 (N_23834,N_15873,N_15369);
nand U23835 (N_23835,N_17954,N_16406);
or U23836 (N_23836,N_18654,N_16846);
nand U23837 (N_23837,N_18432,N_15632);
or U23838 (N_23838,N_19170,N_15073);
or U23839 (N_23839,N_16967,N_19136);
xnor U23840 (N_23840,N_18415,N_19057);
nand U23841 (N_23841,N_19884,N_18342);
and U23842 (N_23842,N_17470,N_16249);
or U23843 (N_23843,N_17594,N_18674);
nand U23844 (N_23844,N_15188,N_19010);
or U23845 (N_23845,N_18668,N_15349);
xnor U23846 (N_23846,N_17231,N_19246);
xnor U23847 (N_23847,N_16638,N_19924);
or U23848 (N_23848,N_16884,N_16830);
or U23849 (N_23849,N_17624,N_16295);
or U23850 (N_23850,N_16414,N_18174);
or U23851 (N_23851,N_19737,N_17667);
and U23852 (N_23852,N_18956,N_17698);
and U23853 (N_23853,N_19875,N_19313);
xor U23854 (N_23854,N_19601,N_18822);
nand U23855 (N_23855,N_16679,N_16041);
or U23856 (N_23856,N_17990,N_16498);
or U23857 (N_23857,N_15734,N_16848);
nor U23858 (N_23858,N_18907,N_16807);
nor U23859 (N_23859,N_17019,N_18399);
nand U23860 (N_23860,N_19104,N_19059);
or U23861 (N_23861,N_16699,N_16517);
nand U23862 (N_23862,N_17613,N_15703);
or U23863 (N_23863,N_18810,N_17832);
or U23864 (N_23864,N_16510,N_16123);
or U23865 (N_23865,N_16363,N_16861);
or U23866 (N_23866,N_19059,N_19921);
and U23867 (N_23867,N_17645,N_18270);
or U23868 (N_23868,N_15363,N_18048);
or U23869 (N_23869,N_17224,N_19737);
and U23870 (N_23870,N_18591,N_19010);
nor U23871 (N_23871,N_19999,N_19765);
nor U23872 (N_23872,N_18115,N_16567);
and U23873 (N_23873,N_19658,N_16541);
or U23874 (N_23874,N_16234,N_19030);
nor U23875 (N_23875,N_16042,N_17867);
and U23876 (N_23876,N_17157,N_16350);
xnor U23877 (N_23877,N_17949,N_15463);
nor U23878 (N_23878,N_15285,N_16802);
or U23879 (N_23879,N_18878,N_17127);
nand U23880 (N_23880,N_18299,N_16938);
nand U23881 (N_23881,N_18624,N_18463);
and U23882 (N_23882,N_17158,N_15281);
nand U23883 (N_23883,N_19524,N_16972);
or U23884 (N_23884,N_18188,N_18483);
nor U23885 (N_23885,N_15575,N_17717);
and U23886 (N_23886,N_15618,N_16401);
or U23887 (N_23887,N_17834,N_18852);
and U23888 (N_23888,N_19048,N_18406);
and U23889 (N_23889,N_19226,N_17460);
nor U23890 (N_23890,N_16273,N_15941);
xor U23891 (N_23891,N_17063,N_18398);
or U23892 (N_23892,N_19391,N_16329);
and U23893 (N_23893,N_17093,N_17366);
xnor U23894 (N_23894,N_19661,N_15482);
nand U23895 (N_23895,N_17580,N_19929);
or U23896 (N_23896,N_19287,N_15542);
nor U23897 (N_23897,N_18885,N_18190);
nand U23898 (N_23898,N_17250,N_18200);
and U23899 (N_23899,N_18374,N_17502);
or U23900 (N_23900,N_18392,N_17953);
xor U23901 (N_23901,N_18911,N_17826);
nor U23902 (N_23902,N_17602,N_17670);
and U23903 (N_23903,N_16693,N_16085);
nor U23904 (N_23904,N_19189,N_19465);
nor U23905 (N_23905,N_15942,N_16264);
xnor U23906 (N_23906,N_15977,N_15139);
or U23907 (N_23907,N_16251,N_19581);
nor U23908 (N_23908,N_17704,N_19576);
nand U23909 (N_23909,N_19638,N_19729);
xnor U23910 (N_23910,N_16373,N_17889);
nor U23911 (N_23911,N_16719,N_17414);
nand U23912 (N_23912,N_19130,N_19976);
nor U23913 (N_23913,N_18744,N_16536);
or U23914 (N_23914,N_18952,N_15785);
or U23915 (N_23915,N_15487,N_17778);
xor U23916 (N_23916,N_17132,N_16532);
xor U23917 (N_23917,N_18336,N_16125);
xor U23918 (N_23918,N_15791,N_19485);
xnor U23919 (N_23919,N_19532,N_18849);
and U23920 (N_23920,N_17246,N_19305);
xnor U23921 (N_23921,N_16874,N_15432);
nand U23922 (N_23922,N_16098,N_16938);
and U23923 (N_23923,N_19625,N_15149);
xnor U23924 (N_23924,N_19430,N_18945);
xor U23925 (N_23925,N_16594,N_17307);
or U23926 (N_23926,N_19525,N_18196);
nor U23927 (N_23927,N_18164,N_15072);
or U23928 (N_23928,N_16363,N_16153);
and U23929 (N_23929,N_18877,N_15933);
xor U23930 (N_23930,N_16339,N_15947);
xor U23931 (N_23931,N_19381,N_15731);
and U23932 (N_23932,N_16434,N_16809);
xor U23933 (N_23933,N_18579,N_16412);
and U23934 (N_23934,N_15452,N_16039);
and U23935 (N_23935,N_15744,N_15045);
and U23936 (N_23936,N_17779,N_18721);
xor U23937 (N_23937,N_16867,N_19875);
and U23938 (N_23938,N_17271,N_16701);
or U23939 (N_23939,N_19398,N_16569);
nand U23940 (N_23940,N_17516,N_16718);
nand U23941 (N_23941,N_16336,N_18961);
nor U23942 (N_23942,N_19296,N_19937);
and U23943 (N_23943,N_16707,N_17300);
nand U23944 (N_23944,N_18237,N_19077);
xnor U23945 (N_23945,N_17753,N_16054);
and U23946 (N_23946,N_19994,N_18965);
and U23947 (N_23947,N_17453,N_15553);
or U23948 (N_23948,N_18408,N_15719);
nand U23949 (N_23949,N_15603,N_16429);
xnor U23950 (N_23950,N_17850,N_17507);
or U23951 (N_23951,N_17557,N_17606);
xnor U23952 (N_23952,N_15224,N_19377);
nand U23953 (N_23953,N_17798,N_17071);
nand U23954 (N_23954,N_17805,N_17102);
nor U23955 (N_23955,N_16928,N_15825);
nand U23956 (N_23956,N_17440,N_16988);
and U23957 (N_23957,N_17173,N_19227);
or U23958 (N_23958,N_19273,N_16793);
nand U23959 (N_23959,N_18091,N_17435);
or U23960 (N_23960,N_19387,N_17807);
nand U23961 (N_23961,N_18675,N_19674);
nor U23962 (N_23962,N_16447,N_17386);
nand U23963 (N_23963,N_19841,N_16838);
or U23964 (N_23964,N_17176,N_15220);
or U23965 (N_23965,N_17363,N_16020);
xnor U23966 (N_23966,N_15884,N_19196);
nand U23967 (N_23967,N_19827,N_19853);
and U23968 (N_23968,N_19765,N_15926);
nor U23969 (N_23969,N_16328,N_19599);
xnor U23970 (N_23970,N_17302,N_16839);
nor U23971 (N_23971,N_15043,N_19886);
xor U23972 (N_23972,N_19408,N_15448);
nand U23973 (N_23973,N_16760,N_17854);
nand U23974 (N_23974,N_18118,N_17322);
nand U23975 (N_23975,N_18830,N_19495);
or U23976 (N_23976,N_19302,N_16781);
nor U23977 (N_23977,N_19276,N_15972);
and U23978 (N_23978,N_18487,N_16650);
nand U23979 (N_23979,N_18871,N_18717);
and U23980 (N_23980,N_16965,N_17915);
xor U23981 (N_23981,N_18882,N_18663);
and U23982 (N_23982,N_15609,N_16655);
or U23983 (N_23983,N_18665,N_17306);
nand U23984 (N_23984,N_18544,N_18972);
nand U23985 (N_23985,N_16122,N_19202);
nand U23986 (N_23986,N_15147,N_19884);
xnor U23987 (N_23987,N_17077,N_18698);
and U23988 (N_23988,N_17225,N_15592);
xor U23989 (N_23989,N_17585,N_15617);
and U23990 (N_23990,N_16515,N_15871);
and U23991 (N_23991,N_15946,N_17930);
and U23992 (N_23992,N_18984,N_17677);
nand U23993 (N_23993,N_15881,N_16020);
or U23994 (N_23994,N_17616,N_15245);
and U23995 (N_23995,N_17083,N_16294);
xor U23996 (N_23996,N_17462,N_17654);
xnor U23997 (N_23997,N_17040,N_19080);
nor U23998 (N_23998,N_19247,N_17275);
xnor U23999 (N_23999,N_15690,N_18213);
and U24000 (N_24000,N_18769,N_19849);
xor U24001 (N_24001,N_16693,N_18930);
xor U24002 (N_24002,N_19593,N_18460);
or U24003 (N_24003,N_18063,N_15307);
nor U24004 (N_24004,N_19321,N_17090);
nor U24005 (N_24005,N_15750,N_16739);
nor U24006 (N_24006,N_17219,N_18293);
xnor U24007 (N_24007,N_19674,N_18512);
nor U24008 (N_24008,N_15723,N_15486);
nand U24009 (N_24009,N_19467,N_15776);
nor U24010 (N_24010,N_18348,N_18726);
nor U24011 (N_24011,N_15395,N_15867);
nand U24012 (N_24012,N_18488,N_15491);
xnor U24013 (N_24013,N_15087,N_18677);
or U24014 (N_24014,N_17078,N_19401);
or U24015 (N_24015,N_15590,N_15420);
nor U24016 (N_24016,N_16240,N_15480);
and U24017 (N_24017,N_17837,N_15505);
nor U24018 (N_24018,N_19902,N_17912);
or U24019 (N_24019,N_15175,N_16936);
or U24020 (N_24020,N_18429,N_18603);
or U24021 (N_24021,N_16568,N_18109);
and U24022 (N_24022,N_16705,N_15435);
or U24023 (N_24023,N_15389,N_19036);
nand U24024 (N_24024,N_15595,N_16502);
and U24025 (N_24025,N_15865,N_16462);
xor U24026 (N_24026,N_15779,N_18222);
and U24027 (N_24027,N_15505,N_15425);
nand U24028 (N_24028,N_15072,N_15177);
and U24029 (N_24029,N_18555,N_18687);
or U24030 (N_24030,N_15382,N_17393);
and U24031 (N_24031,N_15326,N_19411);
nor U24032 (N_24032,N_17481,N_17607);
nor U24033 (N_24033,N_16312,N_18611);
and U24034 (N_24034,N_17919,N_17065);
nand U24035 (N_24035,N_19607,N_15700);
and U24036 (N_24036,N_18101,N_19272);
nor U24037 (N_24037,N_18920,N_19241);
xor U24038 (N_24038,N_17725,N_18232);
and U24039 (N_24039,N_15575,N_19223);
nor U24040 (N_24040,N_16320,N_18657);
or U24041 (N_24041,N_16838,N_15889);
nor U24042 (N_24042,N_16321,N_17852);
or U24043 (N_24043,N_17031,N_19725);
xor U24044 (N_24044,N_19936,N_19923);
nor U24045 (N_24045,N_18085,N_15822);
nand U24046 (N_24046,N_19410,N_16351);
nor U24047 (N_24047,N_16063,N_16832);
and U24048 (N_24048,N_17030,N_19472);
nand U24049 (N_24049,N_19836,N_19659);
xnor U24050 (N_24050,N_15447,N_19084);
nand U24051 (N_24051,N_17263,N_19952);
nand U24052 (N_24052,N_16980,N_19241);
or U24053 (N_24053,N_15577,N_16184);
xor U24054 (N_24054,N_16157,N_17983);
and U24055 (N_24055,N_17042,N_19937);
nand U24056 (N_24056,N_17769,N_18112);
xnor U24057 (N_24057,N_15397,N_17143);
xor U24058 (N_24058,N_17386,N_16840);
nor U24059 (N_24059,N_16134,N_18188);
and U24060 (N_24060,N_18112,N_17529);
xor U24061 (N_24061,N_17238,N_17799);
and U24062 (N_24062,N_18195,N_16099);
or U24063 (N_24063,N_18738,N_15477);
nor U24064 (N_24064,N_17469,N_19008);
or U24065 (N_24065,N_18890,N_16826);
and U24066 (N_24066,N_17546,N_18777);
or U24067 (N_24067,N_15904,N_16791);
or U24068 (N_24068,N_18224,N_15690);
and U24069 (N_24069,N_19609,N_18996);
and U24070 (N_24070,N_16747,N_19725);
nand U24071 (N_24071,N_17107,N_19189);
nand U24072 (N_24072,N_19588,N_16279);
or U24073 (N_24073,N_19075,N_17130);
xnor U24074 (N_24074,N_16663,N_18856);
xor U24075 (N_24075,N_17667,N_16358);
nand U24076 (N_24076,N_18997,N_18709);
nor U24077 (N_24077,N_15071,N_17749);
and U24078 (N_24078,N_19241,N_17373);
or U24079 (N_24079,N_17306,N_18567);
nand U24080 (N_24080,N_15979,N_15888);
and U24081 (N_24081,N_19255,N_18388);
or U24082 (N_24082,N_19376,N_17831);
nand U24083 (N_24083,N_19974,N_15653);
nand U24084 (N_24084,N_18448,N_19579);
or U24085 (N_24085,N_15595,N_18988);
or U24086 (N_24086,N_19730,N_16378);
or U24087 (N_24087,N_15232,N_16810);
nand U24088 (N_24088,N_19995,N_18598);
and U24089 (N_24089,N_15986,N_19674);
xnor U24090 (N_24090,N_17522,N_18353);
xor U24091 (N_24091,N_16157,N_17918);
or U24092 (N_24092,N_18168,N_17155);
and U24093 (N_24093,N_19098,N_16641);
nand U24094 (N_24094,N_15647,N_16450);
nor U24095 (N_24095,N_19724,N_18981);
xor U24096 (N_24096,N_16839,N_17716);
nor U24097 (N_24097,N_17224,N_18818);
nor U24098 (N_24098,N_18334,N_17538);
xnor U24099 (N_24099,N_16833,N_18489);
nand U24100 (N_24100,N_15179,N_19609);
xor U24101 (N_24101,N_15826,N_18322);
nand U24102 (N_24102,N_18646,N_15560);
xnor U24103 (N_24103,N_18001,N_16082);
nand U24104 (N_24104,N_17621,N_17522);
nand U24105 (N_24105,N_19480,N_17866);
and U24106 (N_24106,N_18440,N_18352);
and U24107 (N_24107,N_17760,N_15405);
or U24108 (N_24108,N_19986,N_17101);
nor U24109 (N_24109,N_15593,N_19835);
nand U24110 (N_24110,N_15858,N_15361);
nand U24111 (N_24111,N_19190,N_18817);
nand U24112 (N_24112,N_15707,N_16769);
nor U24113 (N_24113,N_19916,N_16139);
nor U24114 (N_24114,N_16731,N_18540);
nand U24115 (N_24115,N_17406,N_17420);
or U24116 (N_24116,N_17284,N_15512);
nand U24117 (N_24117,N_17974,N_16257);
xor U24118 (N_24118,N_18714,N_16005);
nand U24119 (N_24119,N_17774,N_16244);
and U24120 (N_24120,N_19036,N_15158);
and U24121 (N_24121,N_19467,N_19275);
and U24122 (N_24122,N_15362,N_16709);
nor U24123 (N_24123,N_19971,N_19607);
nor U24124 (N_24124,N_19517,N_16628);
nand U24125 (N_24125,N_16085,N_15299);
and U24126 (N_24126,N_16966,N_17560);
xor U24127 (N_24127,N_16216,N_16495);
and U24128 (N_24128,N_18107,N_15302);
nor U24129 (N_24129,N_15450,N_17607);
nand U24130 (N_24130,N_15473,N_17797);
nor U24131 (N_24131,N_15094,N_15988);
and U24132 (N_24132,N_15179,N_19701);
and U24133 (N_24133,N_19616,N_19183);
and U24134 (N_24134,N_15882,N_17503);
nor U24135 (N_24135,N_18547,N_17837);
and U24136 (N_24136,N_19148,N_19872);
and U24137 (N_24137,N_16616,N_17957);
and U24138 (N_24138,N_15372,N_16193);
nand U24139 (N_24139,N_16657,N_18846);
xnor U24140 (N_24140,N_18396,N_19930);
xor U24141 (N_24141,N_17646,N_15125);
nand U24142 (N_24142,N_19433,N_15776);
nor U24143 (N_24143,N_19984,N_15047);
nand U24144 (N_24144,N_16168,N_16501);
nand U24145 (N_24145,N_16938,N_19413);
and U24146 (N_24146,N_16782,N_19781);
and U24147 (N_24147,N_16626,N_19977);
xor U24148 (N_24148,N_16701,N_18493);
nor U24149 (N_24149,N_16649,N_18991);
and U24150 (N_24150,N_18895,N_15277);
nor U24151 (N_24151,N_16673,N_17550);
or U24152 (N_24152,N_18422,N_16808);
nor U24153 (N_24153,N_16157,N_17359);
nand U24154 (N_24154,N_15184,N_16437);
or U24155 (N_24155,N_18295,N_18233);
or U24156 (N_24156,N_17719,N_18607);
nor U24157 (N_24157,N_15494,N_17447);
or U24158 (N_24158,N_15590,N_18077);
or U24159 (N_24159,N_19832,N_17659);
and U24160 (N_24160,N_19032,N_16242);
xnor U24161 (N_24161,N_17228,N_16816);
nand U24162 (N_24162,N_15713,N_15991);
nor U24163 (N_24163,N_19692,N_19787);
or U24164 (N_24164,N_17504,N_18096);
nor U24165 (N_24165,N_15219,N_19172);
nand U24166 (N_24166,N_15287,N_16156);
and U24167 (N_24167,N_15121,N_17236);
or U24168 (N_24168,N_15340,N_16235);
nand U24169 (N_24169,N_18388,N_16399);
xnor U24170 (N_24170,N_19330,N_18736);
nand U24171 (N_24171,N_15929,N_16208);
nand U24172 (N_24172,N_17699,N_16572);
nor U24173 (N_24173,N_15723,N_17355);
and U24174 (N_24174,N_19075,N_17178);
or U24175 (N_24175,N_18999,N_18531);
nor U24176 (N_24176,N_16703,N_16298);
xnor U24177 (N_24177,N_17433,N_19924);
or U24178 (N_24178,N_15547,N_18604);
xnor U24179 (N_24179,N_17571,N_17654);
and U24180 (N_24180,N_16202,N_18210);
nand U24181 (N_24181,N_17372,N_15693);
or U24182 (N_24182,N_17595,N_17983);
nand U24183 (N_24183,N_18478,N_18716);
nand U24184 (N_24184,N_19340,N_15185);
or U24185 (N_24185,N_19022,N_19117);
or U24186 (N_24186,N_17909,N_15372);
nand U24187 (N_24187,N_19677,N_16451);
xnor U24188 (N_24188,N_18825,N_16318);
or U24189 (N_24189,N_17193,N_17596);
nand U24190 (N_24190,N_16437,N_18498);
xnor U24191 (N_24191,N_15475,N_16869);
and U24192 (N_24192,N_19247,N_16202);
or U24193 (N_24193,N_18342,N_19793);
or U24194 (N_24194,N_18466,N_15170);
nor U24195 (N_24195,N_18659,N_15618);
nand U24196 (N_24196,N_16218,N_19199);
xor U24197 (N_24197,N_15864,N_19825);
or U24198 (N_24198,N_16651,N_16006);
xor U24199 (N_24199,N_18227,N_17376);
xnor U24200 (N_24200,N_19326,N_15468);
and U24201 (N_24201,N_15258,N_16345);
nor U24202 (N_24202,N_16630,N_19525);
nand U24203 (N_24203,N_18103,N_16216);
nand U24204 (N_24204,N_15603,N_18436);
or U24205 (N_24205,N_16186,N_16579);
nand U24206 (N_24206,N_16753,N_19176);
xnor U24207 (N_24207,N_17641,N_17455);
nand U24208 (N_24208,N_16247,N_17862);
and U24209 (N_24209,N_16741,N_15087);
nand U24210 (N_24210,N_19865,N_18583);
nand U24211 (N_24211,N_15031,N_15758);
or U24212 (N_24212,N_18129,N_18243);
nor U24213 (N_24213,N_15927,N_15385);
and U24214 (N_24214,N_16663,N_19205);
and U24215 (N_24215,N_16020,N_17752);
and U24216 (N_24216,N_16723,N_17736);
or U24217 (N_24217,N_16858,N_18432);
xor U24218 (N_24218,N_19377,N_18300);
nor U24219 (N_24219,N_15736,N_15181);
or U24220 (N_24220,N_15762,N_16694);
nor U24221 (N_24221,N_16223,N_17407);
nand U24222 (N_24222,N_15262,N_16490);
xor U24223 (N_24223,N_16176,N_19368);
xnor U24224 (N_24224,N_16734,N_15940);
nor U24225 (N_24225,N_18804,N_15874);
nor U24226 (N_24226,N_18597,N_18078);
nand U24227 (N_24227,N_19084,N_15696);
xnor U24228 (N_24228,N_16504,N_18955);
xor U24229 (N_24229,N_17785,N_19282);
or U24230 (N_24230,N_16220,N_16546);
or U24231 (N_24231,N_17433,N_16445);
nor U24232 (N_24232,N_15638,N_18889);
nor U24233 (N_24233,N_19881,N_18092);
or U24234 (N_24234,N_18008,N_16952);
or U24235 (N_24235,N_15985,N_16280);
or U24236 (N_24236,N_19388,N_17367);
or U24237 (N_24237,N_17529,N_15830);
nand U24238 (N_24238,N_15524,N_16116);
nor U24239 (N_24239,N_17045,N_18783);
nand U24240 (N_24240,N_17189,N_15090);
and U24241 (N_24241,N_18786,N_16493);
xor U24242 (N_24242,N_15385,N_15836);
xor U24243 (N_24243,N_18073,N_16627);
or U24244 (N_24244,N_17311,N_17756);
and U24245 (N_24245,N_17478,N_18823);
nor U24246 (N_24246,N_17894,N_16869);
or U24247 (N_24247,N_18279,N_15026);
and U24248 (N_24248,N_16207,N_16979);
and U24249 (N_24249,N_18782,N_19804);
or U24250 (N_24250,N_18870,N_17751);
and U24251 (N_24251,N_19800,N_16316);
nor U24252 (N_24252,N_15803,N_19004);
nor U24253 (N_24253,N_15816,N_18650);
or U24254 (N_24254,N_18826,N_16298);
and U24255 (N_24255,N_19538,N_17014);
or U24256 (N_24256,N_15523,N_16773);
and U24257 (N_24257,N_18036,N_16986);
xnor U24258 (N_24258,N_19455,N_15607);
nor U24259 (N_24259,N_17350,N_16834);
nor U24260 (N_24260,N_15713,N_19711);
and U24261 (N_24261,N_18639,N_16324);
nand U24262 (N_24262,N_19420,N_15382);
nand U24263 (N_24263,N_19864,N_19801);
nand U24264 (N_24264,N_19073,N_17534);
nor U24265 (N_24265,N_15826,N_18079);
xnor U24266 (N_24266,N_17846,N_19329);
nor U24267 (N_24267,N_19931,N_15535);
and U24268 (N_24268,N_17363,N_16987);
nand U24269 (N_24269,N_16516,N_19240);
nand U24270 (N_24270,N_16339,N_15218);
nand U24271 (N_24271,N_17751,N_18412);
or U24272 (N_24272,N_15472,N_17975);
or U24273 (N_24273,N_17632,N_17213);
nor U24274 (N_24274,N_17208,N_17040);
xor U24275 (N_24275,N_15074,N_18965);
nand U24276 (N_24276,N_18092,N_16748);
and U24277 (N_24277,N_19861,N_17047);
and U24278 (N_24278,N_18818,N_17833);
nand U24279 (N_24279,N_18178,N_16514);
nor U24280 (N_24280,N_19832,N_19423);
xor U24281 (N_24281,N_16195,N_17490);
nor U24282 (N_24282,N_17824,N_15174);
or U24283 (N_24283,N_16420,N_17889);
or U24284 (N_24284,N_19307,N_15703);
nor U24285 (N_24285,N_17125,N_17345);
xnor U24286 (N_24286,N_15323,N_18722);
or U24287 (N_24287,N_18055,N_17930);
nor U24288 (N_24288,N_18605,N_19237);
or U24289 (N_24289,N_16709,N_16986);
and U24290 (N_24290,N_18858,N_19411);
and U24291 (N_24291,N_15992,N_15259);
nand U24292 (N_24292,N_17596,N_19686);
xor U24293 (N_24293,N_18302,N_19940);
or U24294 (N_24294,N_15903,N_19750);
and U24295 (N_24295,N_15742,N_15789);
nor U24296 (N_24296,N_16524,N_19506);
xnor U24297 (N_24297,N_19477,N_19900);
nand U24298 (N_24298,N_16806,N_17722);
nand U24299 (N_24299,N_18097,N_19445);
and U24300 (N_24300,N_17883,N_18996);
or U24301 (N_24301,N_16860,N_15571);
or U24302 (N_24302,N_17617,N_19487);
or U24303 (N_24303,N_15869,N_17540);
or U24304 (N_24304,N_18818,N_15863);
xor U24305 (N_24305,N_17920,N_15884);
or U24306 (N_24306,N_19448,N_15040);
nor U24307 (N_24307,N_16553,N_15112);
or U24308 (N_24308,N_15522,N_15383);
xor U24309 (N_24309,N_16864,N_18337);
xor U24310 (N_24310,N_19164,N_15448);
or U24311 (N_24311,N_16619,N_19776);
xor U24312 (N_24312,N_16992,N_15937);
or U24313 (N_24313,N_15192,N_15380);
nor U24314 (N_24314,N_17875,N_18090);
nor U24315 (N_24315,N_19152,N_15026);
or U24316 (N_24316,N_16973,N_16994);
or U24317 (N_24317,N_16835,N_19042);
or U24318 (N_24318,N_17718,N_15585);
and U24319 (N_24319,N_18360,N_16641);
nor U24320 (N_24320,N_15063,N_16177);
xor U24321 (N_24321,N_19818,N_16658);
nand U24322 (N_24322,N_19029,N_17561);
xnor U24323 (N_24323,N_18961,N_19817);
nand U24324 (N_24324,N_18033,N_15693);
and U24325 (N_24325,N_15121,N_18521);
nand U24326 (N_24326,N_17452,N_18924);
nand U24327 (N_24327,N_16785,N_19365);
and U24328 (N_24328,N_17803,N_17719);
or U24329 (N_24329,N_17146,N_19757);
or U24330 (N_24330,N_17444,N_19170);
or U24331 (N_24331,N_16597,N_18455);
nor U24332 (N_24332,N_16525,N_18549);
and U24333 (N_24333,N_15411,N_15373);
xor U24334 (N_24334,N_16877,N_17770);
xnor U24335 (N_24335,N_19110,N_16932);
or U24336 (N_24336,N_19587,N_16021);
nor U24337 (N_24337,N_16456,N_15013);
nand U24338 (N_24338,N_15312,N_16883);
nand U24339 (N_24339,N_17834,N_18473);
nand U24340 (N_24340,N_16844,N_19992);
nand U24341 (N_24341,N_16371,N_19006);
nand U24342 (N_24342,N_18403,N_15314);
nand U24343 (N_24343,N_17159,N_16621);
nand U24344 (N_24344,N_18628,N_19388);
xor U24345 (N_24345,N_19019,N_19304);
nor U24346 (N_24346,N_18236,N_15813);
and U24347 (N_24347,N_17192,N_17767);
and U24348 (N_24348,N_15171,N_17880);
or U24349 (N_24349,N_18577,N_18553);
nand U24350 (N_24350,N_17558,N_18695);
and U24351 (N_24351,N_19074,N_18356);
xnor U24352 (N_24352,N_16377,N_19230);
nor U24353 (N_24353,N_19510,N_15152);
or U24354 (N_24354,N_17280,N_17892);
or U24355 (N_24355,N_18982,N_15499);
nor U24356 (N_24356,N_16134,N_16772);
nor U24357 (N_24357,N_19811,N_18707);
nand U24358 (N_24358,N_15995,N_18814);
nor U24359 (N_24359,N_18105,N_18442);
or U24360 (N_24360,N_15346,N_16401);
and U24361 (N_24361,N_19545,N_18716);
and U24362 (N_24362,N_17914,N_17493);
nand U24363 (N_24363,N_18702,N_18740);
or U24364 (N_24364,N_18770,N_18956);
nand U24365 (N_24365,N_15761,N_18197);
or U24366 (N_24366,N_18836,N_19597);
nor U24367 (N_24367,N_17898,N_15035);
nor U24368 (N_24368,N_17747,N_17436);
nand U24369 (N_24369,N_15667,N_17741);
nor U24370 (N_24370,N_16406,N_19997);
or U24371 (N_24371,N_17966,N_18007);
or U24372 (N_24372,N_19887,N_16293);
nand U24373 (N_24373,N_16705,N_18212);
or U24374 (N_24374,N_16435,N_16531);
nand U24375 (N_24375,N_19166,N_16272);
nand U24376 (N_24376,N_18951,N_16294);
nand U24377 (N_24377,N_19587,N_19920);
and U24378 (N_24378,N_19415,N_18129);
xnor U24379 (N_24379,N_17983,N_19381);
nand U24380 (N_24380,N_18190,N_19176);
xor U24381 (N_24381,N_17976,N_17401);
nor U24382 (N_24382,N_17794,N_17689);
xnor U24383 (N_24383,N_15554,N_17077);
or U24384 (N_24384,N_19213,N_19099);
and U24385 (N_24385,N_15638,N_17779);
nor U24386 (N_24386,N_18709,N_16673);
xnor U24387 (N_24387,N_16748,N_19119);
nor U24388 (N_24388,N_18103,N_17123);
nand U24389 (N_24389,N_18854,N_19340);
or U24390 (N_24390,N_18354,N_16754);
nor U24391 (N_24391,N_19708,N_19438);
or U24392 (N_24392,N_15081,N_15116);
nor U24393 (N_24393,N_15333,N_15945);
nor U24394 (N_24394,N_17480,N_16172);
and U24395 (N_24395,N_18475,N_17127);
or U24396 (N_24396,N_18138,N_19800);
nand U24397 (N_24397,N_17339,N_19909);
nor U24398 (N_24398,N_16601,N_19817);
and U24399 (N_24399,N_19192,N_16358);
xnor U24400 (N_24400,N_16339,N_19009);
nand U24401 (N_24401,N_16203,N_19475);
xnor U24402 (N_24402,N_17085,N_16414);
xor U24403 (N_24403,N_15016,N_16698);
and U24404 (N_24404,N_16864,N_18820);
nor U24405 (N_24405,N_15879,N_18653);
nor U24406 (N_24406,N_16239,N_16814);
nor U24407 (N_24407,N_15725,N_16145);
and U24408 (N_24408,N_17696,N_19973);
nor U24409 (N_24409,N_18299,N_19432);
or U24410 (N_24410,N_18027,N_17470);
xnor U24411 (N_24411,N_16215,N_17151);
or U24412 (N_24412,N_19100,N_19602);
nor U24413 (N_24413,N_15160,N_15085);
nand U24414 (N_24414,N_17317,N_16981);
nand U24415 (N_24415,N_18718,N_16793);
or U24416 (N_24416,N_19052,N_18557);
and U24417 (N_24417,N_18255,N_19997);
nor U24418 (N_24418,N_19563,N_17033);
and U24419 (N_24419,N_17921,N_17843);
nor U24420 (N_24420,N_16086,N_16495);
nor U24421 (N_24421,N_19420,N_19777);
nand U24422 (N_24422,N_17796,N_19364);
and U24423 (N_24423,N_17908,N_18225);
nand U24424 (N_24424,N_17916,N_17976);
nor U24425 (N_24425,N_19210,N_15110);
nor U24426 (N_24426,N_17250,N_19001);
nand U24427 (N_24427,N_16122,N_17128);
xor U24428 (N_24428,N_17135,N_17213);
or U24429 (N_24429,N_17470,N_19042);
nor U24430 (N_24430,N_16194,N_17672);
nand U24431 (N_24431,N_17577,N_15584);
nand U24432 (N_24432,N_16377,N_19664);
xnor U24433 (N_24433,N_19846,N_19189);
or U24434 (N_24434,N_15157,N_16454);
or U24435 (N_24435,N_19866,N_17579);
and U24436 (N_24436,N_15398,N_19325);
or U24437 (N_24437,N_16796,N_17923);
nand U24438 (N_24438,N_19259,N_16907);
nand U24439 (N_24439,N_17478,N_15006);
or U24440 (N_24440,N_19769,N_19324);
nand U24441 (N_24441,N_15853,N_16373);
and U24442 (N_24442,N_16483,N_15665);
nand U24443 (N_24443,N_15925,N_19791);
nand U24444 (N_24444,N_15545,N_17779);
or U24445 (N_24445,N_18660,N_16876);
xor U24446 (N_24446,N_18558,N_15943);
xor U24447 (N_24447,N_18632,N_16542);
or U24448 (N_24448,N_18320,N_19031);
and U24449 (N_24449,N_16812,N_15685);
and U24450 (N_24450,N_16198,N_17116);
or U24451 (N_24451,N_16518,N_16635);
nor U24452 (N_24452,N_16794,N_17810);
and U24453 (N_24453,N_19725,N_19799);
xor U24454 (N_24454,N_16921,N_17463);
nor U24455 (N_24455,N_18337,N_15486);
or U24456 (N_24456,N_19796,N_18729);
or U24457 (N_24457,N_18466,N_19140);
nor U24458 (N_24458,N_16370,N_17183);
or U24459 (N_24459,N_18217,N_15331);
nand U24460 (N_24460,N_16282,N_19259);
and U24461 (N_24461,N_15939,N_18783);
nand U24462 (N_24462,N_19055,N_17134);
xnor U24463 (N_24463,N_18188,N_18418);
and U24464 (N_24464,N_18169,N_18769);
nand U24465 (N_24465,N_18738,N_15034);
xnor U24466 (N_24466,N_19375,N_15406);
nor U24467 (N_24467,N_18732,N_15882);
nand U24468 (N_24468,N_15526,N_15933);
nor U24469 (N_24469,N_16809,N_17906);
nor U24470 (N_24470,N_18367,N_16651);
nor U24471 (N_24471,N_15878,N_17180);
and U24472 (N_24472,N_17754,N_17786);
or U24473 (N_24473,N_19916,N_15689);
or U24474 (N_24474,N_17290,N_18173);
nor U24475 (N_24475,N_16562,N_15712);
nand U24476 (N_24476,N_19171,N_16922);
nor U24477 (N_24477,N_15641,N_15566);
nand U24478 (N_24478,N_15276,N_16369);
nor U24479 (N_24479,N_15974,N_16293);
nand U24480 (N_24480,N_16622,N_15135);
nand U24481 (N_24481,N_16399,N_18834);
nand U24482 (N_24482,N_16140,N_19431);
xnor U24483 (N_24483,N_19366,N_19721);
xor U24484 (N_24484,N_15011,N_18642);
or U24485 (N_24485,N_16517,N_17841);
nand U24486 (N_24486,N_15940,N_15288);
and U24487 (N_24487,N_18171,N_17722);
or U24488 (N_24488,N_19086,N_18865);
or U24489 (N_24489,N_17798,N_18757);
nor U24490 (N_24490,N_18284,N_18033);
nand U24491 (N_24491,N_18396,N_18521);
nand U24492 (N_24492,N_15103,N_18874);
or U24493 (N_24493,N_19825,N_18353);
or U24494 (N_24494,N_15820,N_19357);
nor U24495 (N_24495,N_16241,N_19849);
or U24496 (N_24496,N_16952,N_16470);
nor U24497 (N_24497,N_18908,N_17208);
xnor U24498 (N_24498,N_16584,N_16089);
and U24499 (N_24499,N_18481,N_19977);
and U24500 (N_24500,N_18491,N_19647);
xor U24501 (N_24501,N_15403,N_15832);
xnor U24502 (N_24502,N_19273,N_15431);
xor U24503 (N_24503,N_15246,N_15153);
nand U24504 (N_24504,N_15176,N_17751);
xor U24505 (N_24505,N_16059,N_16548);
nor U24506 (N_24506,N_19334,N_18807);
nor U24507 (N_24507,N_17391,N_18096);
nand U24508 (N_24508,N_17798,N_15192);
nand U24509 (N_24509,N_19365,N_17463);
and U24510 (N_24510,N_16548,N_16029);
nand U24511 (N_24511,N_18590,N_15307);
or U24512 (N_24512,N_15955,N_15522);
nand U24513 (N_24513,N_19925,N_16920);
nor U24514 (N_24514,N_15287,N_17119);
xnor U24515 (N_24515,N_16177,N_15840);
and U24516 (N_24516,N_19574,N_18818);
xnor U24517 (N_24517,N_17783,N_15500);
or U24518 (N_24518,N_18665,N_15183);
and U24519 (N_24519,N_17002,N_18234);
or U24520 (N_24520,N_18800,N_17336);
and U24521 (N_24521,N_18069,N_16331);
or U24522 (N_24522,N_19866,N_19888);
nand U24523 (N_24523,N_17442,N_17119);
or U24524 (N_24524,N_18815,N_15741);
xor U24525 (N_24525,N_18791,N_19175);
nor U24526 (N_24526,N_16331,N_17653);
xor U24527 (N_24527,N_15120,N_18597);
xnor U24528 (N_24528,N_16979,N_16548);
or U24529 (N_24529,N_15458,N_17441);
nand U24530 (N_24530,N_18123,N_15984);
nor U24531 (N_24531,N_17948,N_15689);
nand U24532 (N_24532,N_19559,N_17982);
nand U24533 (N_24533,N_18757,N_16200);
and U24534 (N_24534,N_19095,N_17299);
and U24535 (N_24535,N_18694,N_15814);
nand U24536 (N_24536,N_15208,N_15832);
nand U24537 (N_24537,N_19915,N_15374);
or U24538 (N_24538,N_18018,N_15706);
nor U24539 (N_24539,N_16673,N_18662);
nor U24540 (N_24540,N_16688,N_19464);
nand U24541 (N_24541,N_16001,N_17585);
nor U24542 (N_24542,N_15205,N_16196);
nand U24543 (N_24543,N_19291,N_17762);
and U24544 (N_24544,N_15179,N_17534);
nand U24545 (N_24545,N_18735,N_17997);
or U24546 (N_24546,N_17625,N_17573);
and U24547 (N_24547,N_15614,N_18526);
nand U24548 (N_24548,N_19048,N_17346);
xor U24549 (N_24549,N_18906,N_18947);
nor U24550 (N_24550,N_19248,N_17388);
nand U24551 (N_24551,N_19541,N_17112);
nand U24552 (N_24552,N_19276,N_17668);
xor U24553 (N_24553,N_19801,N_17395);
nand U24554 (N_24554,N_16572,N_19264);
nand U24555 (N_24555,N_17604,N_16184);
xnor U24556 (N_24556,N_18418,N_16761);
xnor U24557 (N_24557,N_15436,N_16120);
and U24558 (N_24558,N_19661,N_16982);
xor U24559 (N_24559,N_19139,N_17148);
or U24560 (N_24560,N_16218,N_15097);
nor U24561 (N_24561,N_18475,N_19939);
nor U24562 (N_24562,N_18281,N_17715);
xor U24563 (N_24563,N_18785,N_15765);
xnor U24564 (N_24564,N_18707,N_17135);
xnor U24565 (N_24565,N_18663,N_17943);
xnor U24566 (N_24566,N_17289,N_18449);
or U24567 (N_24567,N_18691,N_16143);
or U24568 (N_24568,N_19271,N_19105);
nor U24569 (N_24569,N_18600,N_17387);
nor U24570 (N_24570,N_16308,N_19384);
nor U24571 (N_24571,N_18520,N_17416);
and U24572 (N_24572,N_16561,N_18223);
xnor U24573 (N_24573,N_16452,N_15011);
nor U24574 (N_24574,N_15395,N_17079);
or U24575 (N_24575,N_17583,N_17338);
nand U24576 (N_24576,N_18495,N_17667);
xnor U24577 (N_24577,N_19767,N_15048);
and U24578 (N_24578,N_18205,N_15299);
xnor U24579 (N_24579,N_17959,N_17747);
nand U24580 (N_24580,N_17715,N_17736);
nor U24581 (N_24581,N_15815,N_16684);
nand U24582 (N_24582,N_19484,N_15043);
or U24583 (N_24583,N_18288,N_18310);
and U24584 (N_24584,N_19124,N_16572);
nand U24585 (N_24585,N_17700,N_17960);
and U24586 (N_24586,N_15487,N_19272);
and U24587 (N_24587,N_19114,N_17566);
nand U24588 (N_24588,N_17857,N_15065);
nor U24589 (N_24589,N_19416,N_15793);
nor U24590 (N_24590,N_19609,N_15899);
xnor U24591 (N_24591,N_19090,N_15098);
or U24592 (N_24592,N_16982,N_15326);
xor U24593 (N_24593,N_15974,N_16023);
nor U24594 (N_24594,N_16671,N_16287);
nand U24595 (N_24595,N_17231,N_15215);
nor U24596 (N_24596,N_16289,N_15275);
nor U24597 (N_24597,N_19449,N_19166);
nand U24598 (N_24598,N_18157,N_15694);
and U24599 (N_24599,N_18894,N_19698);
nor U24600 (N_24600,N_17159,N_18125);
xor U24601 (N_24601,N_19058,N_17201);
nor U24602 (N_24602,N_18945,N_17484);
or U24603 (N_24603,N_15769,N_19515);
nor U24604 (N_24604,N_17492,N_16394);
xor U24605 (N_24605,N_16164,N_19527);
or U24606 (N_24606,N_17520,N_19547);
and U24607 (N_24607,N_19431,N_17641);
xnor U24608 (N_24608,N_15427,N_17150);
and U24609 (N_24609,N_17806,N_16931);
and U24610 (N_24610,N_17661,N_15447);
and U24611 (N_24611,N_18863,N_19468);
or U24612 (N_24612,N_15550,N_17711);
nor U24613 (N_24613,N_19005,N_15689);
nand U24614 (N_24614,N_19525,N_19127);
nor U24615 (N_24615,N_18938,N_15716);
nand U24616 (N_24616,N_16739,N_19581);
nand U24617 (N_24617,N_15426,N_19877);
or U24618 (N_24618,N_18247,N_17254);
and U24619 (N_24619,N_18604,N_18205);
nor U24620 (N_24620,N_19591,N_18758);
nand U24621 (N_24621,N_17755,N_18284);
or U24622 (N_24622,N_17535,N_16799);
and U24623 (N_24623,N_16358,N_15046);
and U24624 (N_24624,N_19938,N_18945);
nand U24625 (N_24625,N_17780,N_18009);
nand U24626 (N_24626,N_17699,N_16998);
and U24627 (N_24627,N_18507,N_18076);
nor U24628 (N_24628,N_16391,N_17041);
nor U24629 (N_24629,N_15886,N_17721);
and U24630 (N_24630,N_16170,N_19062);
nand U24631 (N_24631,N_17397,N_19150);
and U24632 (N_24632,N_16869,N_19035);
xnor U24633 (N_24633,N_15454,N_16678);
nor U24634 (N_24634,N_17620,N_15298);
nand U24635 (N_24635,N_18612,N_16452);
and U24636 (N_24636,N_19938,N_19206);
and U24637 (N_24637,N_16455,N_17401);
nor U24638 (N_24638,N_15013,N_19653);
or U24639 (N_24639,N_15457,N_17368);
or U24640 (N_24640,N_19910,N_19703);
xor U24641 (N_24641,N_19401,N_19326);
and U24642 (N_24642,N_18621,N_15582);
or U24643 (N_24643,N_16968,N_15751);
and U24644 (N_24644,N_15808,N_18418);
nor U24645 (N_24645,N_15934,N_15806);
xor U24646 (N_24646,N_15180,N_18058);
nand U24647 (N_24647,N_16863,N_16829);
and U24648 (N_24648,N_15876,N_18726);
nor U24649 (N_24649,N_17147,N_18754);
xnor U24650 (N_24650,N_16802,N_19694);
and U24651 (N_24651,N_15385,N_18783);
nor U24652 (N_24652,N_17467,N_19393);
or U24653 (N_24653,N_19226,N_19533);
nand U24654 (N_24654,N_18442,N_15176);
nor U24655 (N_24655,N_18999,N_18823);
nand U24656 (N_24656,N_15349,N_15151);
xor U24657 (N_24657,N_19753,N_19119);
or U24658 (N_24658,N_18522,N_17933);
and U24659 (N_24659,N_15989,N_16935);
xor U24660 (N_24660,N_18975,N_18557);
xnor U24661 (N_24661,N_19719,N_15263);
xor U24662 (N_24662,N_19357,N_17196);
nor U24663 (N_24663,N_18078,N_16071);
nor U24664 (N_24664,N_15631,N_18116);
nor U24665 (N_24665,N_15784,N_16743);
xor U24666 (N_24666,N_17751,N_16303);
nor U24667 (N_24667,N_17518,N_19341);
or U24668 (N_24668,N_15514,N_15790);
nor U24669 (N_24669,N_16864,N_18372);
nor U24670 (N_24670,N_18653,N_18861);
xor U24671 (N_24671,N_15952,N_19946);
or U24672 (N_24672,N_18479,N_15759);
and U24673 (N_24673,N_19617,N_19263);
and U24674 (N_24674,N_19382,N_19817);
and U24675 (N_24675,N_19832,N_18134);
or U24676 (N_24676,N_19117,N_15482);
nand U24677 (N_24677,N_15318,N_18228);
or U24678 (N_24678,N_18982,N_17822);
xor U24679 (N_24679,N_15023,N_19699);
nand U24680 (N_24680,N_18010,N_15524);
xnor U24681 (N_24681,N_19520,N_15042);
or U24682 (N_24682,N_17500,N_19755);
or U24683 (N_24683,N_19622,N_18511);
and U24684 (N_24684,N_16287,N_18129);
xor U24685 (N_24685,N_16674,N_18732);
nand U24686 (N_24686,N_16089,N_15433);
nand U24687 (N_24687,N_17185,N_16633);
nand U24688 (N_24688,N_15241,N_19949);
nor U24689 (N_24689,N_17730,N_18477);
nand U24690 (N_24690,N_17461,N_15104);
xor U24691 (N_24691,N_19893,N_19753);
and U24692 (N_24692,N_17310,N_15108);
and U24693 (N_24693,N_18959,N_19718);
nor U24694 (N_24694,N_15076,N_16356);
nor U24695 (N_24695,N_15629,N_16261);
nand U24696 (N_24696,N_17723,N_16692);
xnor U24697 (N_24697,N_18059,N_19367);
nand U24698 (N_24698,N_19156,N_17906);
or U24699 (N_24699,N_16929,N_15885);
nor U24700 (N_24700,N_15128,N_19078);
nor U24701 (N_24701,N_15967,N_17074);
and U24702 (N_24702,N_18226,N_15841);
or U24703 (N_24703,N_16968,N_16670);
nand U24704 (N_24704,N_15075,N_17684);
and U24705 (N_24705,N_17589,N_15321);
nor U24706 (N_24706,N_17554,N_19462);
nand U24707 (N_24707,N_16705,N_17817);
nand U24708 (N_24708,N_19215,N_18750);
and U24709 (N_24709,N_16255,N_15120);
nor U24710 (N_24710,N_18441,N_16951);
or U24711 (N_24711,N_17525,N_19726);
nand U24712 (N_24712,N_18362,N_18854);
xnor U24713 (N_24713,N_19414,N_19977);
xor U24714 (N_24714,N_19850,N_19311);
xor U24715 (N_24715,N_15102,N_19833);
or U24716 (N_24716,N_16025,N_18857);
nand U24717 (N_24717,N_18808,N_19603);
nand U24718 (N_24718,N_15947,N_16201);
nand U24719 (N_24719,N_18226,N_15092);
nand U24720 (N_24720,N_18297,N_16111);
or U24721 (N_24721,N_17260,N_17986);
xnor U24722 (N_24722,N_18037,N_18283);
xor U24723 (N_24723,N_16882,N_17432);
xor U24724 (N_24724,N_19280,N_18240);
or U24725 (N_24725,N_15738,N_15305);
or U24726 (N_24726,N_15949,N_16563);
nand U24727 (N_24727,N_19977,N_19339);
nand U24728 (N_24728,N_15059,N_18245);
nor U24729 (N_24729,N_16165,N_17829);
nand U24730 (N_24730,N_19403,N_15766);
or U24731 (N_24731,N_17083,N_18935);
or U24732 (N_24732,N_17800,N_17824);
xor U24733 (N_24733,N_16097,N_15497);
and U24734 (N_24734,N_16230,N_18353);
xor U24735 (N_24735,N_16378,N_17514);
and U24736 (N_24736,N_19430,N_18993);
nor U24737 (N_24737,N_18395,N_19186);
or U24738 (N_24738,N_19912,N_18043);
nor U24739 (N_24739,N_15951,N_16865);
nor U24740 (N_24740,N_15407,N_16592);
xnor U24741 (N_24741,N_18047,N_15116);
or U24742 (N_24742,N_19111,N_17853);
nor U24743 (N_24743,N_18976,N_19957);
nor U24744 (N_24744,N_19570,N_15920);
nor U24745 (N_24745,N_19917,N_19193);
or U24746 (N_24746,N_16576,N_15420);
nand U24747 (N_24747,N_17944,N_16495);
xnor U24748 (N_24748,N_19393,N_16520);
nand U24749 (N_24749,N_16523,N_18720);
nor U24750 (N_24750,N_15534,N_15008);
or U24751 (N_24751,N_15123,N_15507);
and U24752 (N_24752,N_16641,N_16053);
nand U24753 (N_24753,N_15158,N_18820);
nand U24754 (N_24754,N_19461,N_19884);
xnor U24755 (N_24755,N_15712,N_15971);
or U24756 (N_24756,N_16142,N_19218);
nand U24757 (N_24757,N_19979,N_19575);
nor U24758 (N_24758,N_18830,N_17267);
and U24759 (N_24759,N_16233,N_15958);
nor U24760 (N_24760,N_19173,N_19091);
nand U24761 (N_24761,N_16494,N_15304);
and U24762 (N_24762,N_18860,N_19133);
or U24763 (N_24763,N_19634,N_16346);
xnor U24764 (N_24764,N_17259,N_17467);
xnor U24765 (N_24765,N_15522,N_18846);
xor U24766 (N_24766,N_17416,N_19832);
and U24767 (N_24767,N_19594,N_15554);
or U24768 (N_24768,N_19526,N_18322);
xnor U24769 (N_24769,N_17438,N_15047);
nand U24770 (N_24770,N_15702,N_19137);
or U24771 (N_24771,N_17640,N_19917);
and U24772 (N_24772,N_18412,N_15448);
or U24773 (N_24773,N_19833,N_17344);
nor U24774 (N_24774,N_18114,N_16958);
and U24775 (N_24775,N_17952,N_17688);
nor U24776 (N_24776,N_19423,N_18925);
or U24777 (N_24777,N_18253,N_15612);
and U24778 (N_24778,N_16752,N_15395);
nand U24779 (N_24779,N_15228,N_18241);
and U24780 (N_24780,N_17994,N_16589);
or U24781 (N_24781,N_17884,N_15140);
xnor U24782 (N_24782,N_19027,N_17228);
nor U24783 (N_24783,N_18301,N_17980);
and U24784 (N_24784,N_16138,N_19956);
xnor U24785 (N_24785,N_15647,N_18050);
and U24786 (N_24786,N_15370,N_19033);
and U24787 (N_24787,N_15445,N_15237);
or U24788 (N_24788,N_17902,N_16862);
nor U24789 (N_24789,N_15988,N_18945);
xnor U24790 (N_24790,N_15381,N_16197);
and U24791 (N_24791,N_16648,N_19854);
xor U24792 (N_24792,N_16794,N_16327);
or U24793 (N_24793,N_19597,N_15030);
nor U24794 (N_24794,N_17388,N_15028);
nor U24795 (N_24795,N_16337,N_15679);
nor U24796 (N_24796,N_15782,N_16082);
xnor U24797 (N_24797,N_15263,N_19821);
nor U24798 (N_24798,N_17769,N_19889);
xnor U24799 (N_24799,N_17890,N_16577);
nor U24800 (N_24800,N_17534,N_19229);
and U24801 (N_24801,N_17760,N_16838);
nor U24802 (N_24802,N_15613,N_18261);
or U24803 (N_24803,N_18352,N_17342);
nor U24804 (N_24804,N_19548,N_15502);
nor U24805 (N_24805,N_19491,N_15618);
nand U24806 (N_24806,N_15282,N_18016);
and U24807 (N_24807,N_19779,N_17822);
and U24808 (N_24808,N_18767,N_19489);
nor U24809 (N_24809,N_18969,N_19016);
or U24810 (N_24810,N_15280,N_17069);
nor U24811 (N_24811,N_16188,N_19154);
nand U24812 (N_24812,N_19018,N_17320);
or U24813 (N_24813,N_15291,N_15552);
or U24814 (N_24814,N_17326,N_16437);
nand U24815 (N_24815,N_19736,N_16231);
nand U24816 (N_24816,N_17749,N_15224);
and U24817 (N_24817,N_16606,N_16127);
xnor U24818 (N_24818,N_16657,N_18240);
nand U24819 (N_24819,N_19496,N_15199);
xor U24820 (N_24820,N_18458,N_15694);
xor U24821 (N_24821,N_19144,N_17429);
nand U24822 (N_24822,N_18359,N_19605);
or U24823 (N_24823,N_17731,N_19135);
nand U24824 (N_24824,N_16079,N_18043);
and U24825 (N_24825,N_18668,N_16999);
nor U24826 (N_24826,N_16905,N_15699);
and U24827 (N_24827,N_17481,N_16700);
or U24828 (N_24828,N_17428,N_18267);
nand U24829 (N_24829,N_17425,N_15769);
and U24830 (N_24830,N_15539,N_18536);
or U24831 (N_24831,N_18375,N_16673);
nor U24832 (N_24832,N_17116,N_19207);
nor U24833 (N_24833,N_15336,N_19240);
nor U24834 (N_24834,N_18794,N_18305);
and U24835 (N_24835,N_15726,N_18168);
and U24836 (N_24836,N_16052,N_18498);
xor U24837 (N_24837,N_16711,N_15838);
and U24838 (N_24838,N_19492,N_15952);
or U24839 (N_24839,N_16113,N_15108);
and U24840 (N_24840,N_16676,N_19781);
xor U24841 (N_24841,N_18980,N_18491);
and U24842 (N_24842,N_17940,N_18106);
or U24843 (N_24843,N_16180,N_18117);
nand U24844 (N_24844,N_19030,N_15240);
xnor U24845 (N_24845,N_17423,N_17852);
nor U24846 (N_24846,N_17676,N_17764);
and U24847 (N_24847,N_17712,N_16530);
nor U24848 (N_24848,N_17981,N_15626);
or U24849 (N_24849,N_19326,N_17192);
nand U24850 (N_24850,N_18229,N_15079);
nor U24851 (N_24851,N_18597,N_15331);
nor U24852 (N_24852,N_19202,N_19465);
nor U24853 (N_24853,N_19779,N_17228);
nor U24854 (N_24854,N_16741,N_17701);
nand U24855 (N_24855,N_18890,N_16193);
nor U24856 (N_24856,N_17491,N_17156);
nor U24857 (N_24857,N_16601,N_18926);
nor U24858 (N_24858,N_16935,N_16782);
nor U24859 (N_24859,N_18718,N_15961);
and U24860 (N_24860,N_18788,N_18885);
or U24861 (N_24861,N_15395,N_19301);
xnor U24862 (N_24862,N_15117,N_17351);
and U24863 (N_24863,N_16669,N_17743);
xor U24864 (N_24864,N_17190,N_19563);
nor U24865 (N_24865,N_16409,N_17766);
xnor U24866 (N_24866,N_19309,N_19969);
or U24867 (N_24867,N_18656,N_19798);
or U24868 (N_24868,N_18319,N_19793);
and U24869 (N_24869,N_15526,N_18068);
xnor U24870 (N_24870,N_15208,N_18690);
nand U24871 (N_24871,N_17506,N_18601);
nor U24872 (N_24872,N_18905,N_17579);
nand U24873 (N_24873,N_17525,N_19665);
xor U24874 (N_24874,N_18183,N_15075);
or U24875 (N_24875,N_18719,N_18505);
xor U24876 (N_24876,N_15893,N_16958);
nor U24877 (N_24877,N_17163,N_17445);
nand U24878 (N_24878,N_15565,N_16676);
and U24879 (N_24879,N_16995,N_15792);
xor U24880 (N_24880,N_16832,N_19488);
nand U24881 (N_24881,N_16191,N_19897);
or U24882 (N_24882,N_18805,N_19595);
nand U24883 (N_24883,N_19531,N_17466);
or U24884 (N_24884,N_17937,N_15832);
xnor U24885 (N_24885,N_16998,N_16013);
nand U24886 (N_24886,N_16720,N_15016);
or U24887 (N_24887,N_16786,N_15296);
or U24888 (N_24888,N_18021,N_15944);
xor U24889 (N_24889,N_19404,N_16909);
or U24890 (N_24890,N_16941,N_19195);
nand U24891 (N_24891,N_18053,N_15049);
and U24892 (N_24892,N_15325,N_17558);
nor U24893 (N_24893,N_15901,N_16428);
or U24894 (N_24894,N_15275,N_19340);
and U24895 (N_24895,N_18172,N_19687);
and U24896 (N_24896,N_18840,N_15634);
nand U24897 (N_24897,N_15095,N_16391);
and U24898 (N_24898,N_17855,N_17804);
or U24899 (N_24899,N_19343,N_18611);
and U24900 (N_24900,N_15133,N_19210);
nor U24901 (N_24901,N_17672,N_18427);
nor U24902 (N_24902,N_17150,N_17830);
nor U24903 (N_24903,N_19522,N_16974);
nand U24904 (N_24904,N_16235,N_19274);
and U24905 (N_24905,N_18722,N_15832);
nor U24906 (N_24906,N_16602,N_19177);
xor U24907 (N_24907,N_19057,N_15503);
and U24908 (N_24908,N_18795,N_16789);
nand U24909 (N_24909,N_19369,N_17694);
and U24910 (N_24910,N_18011,N_16534);
nor U24911 (N_24911,N_17052,N_15962);
and U24912 (N_24912,N_16954,N_16343);
or U24913 (N_24913,N_15281,N_17284);
nor U24914 (N_24914,N_19909,N_15892);
or U24915 (N_24915,N_19628,N_18968);
and U24916 (N_24916,N_18994,N_17954);
xor U24917 (N_24917,N_16316,N_15205);
nand U24918 (N_24918,N_18265,N_15041);
and U24919 (N_24919,N_18997,N_17261);
or U24920 (N_24920,N_17611,N_15687);
nand U24921 (N_24921,N_19080,N_15472);
nand U24922 (N_24922,N_16910,N_16009);
nor U24923 (N_24923,N_19916,N_17912);
and U24924 (N_24924,N_18993,N_16990);
xor U24925 (N_24925,N_16621,N_19645);
or U24926 (N_24926,N_16750,N_17333);
nor U24927 (N_24927,N_17045,N_15751);
and U24928 (N_24928,N_19767,N_19374);
and U24929 (N_24929,N_15912,N_19790);
nand U24930 (N_24930,N_15376,N_19447);
xnor U24931 (N_24931,N_17371,N_18682);
xor U24932 (N_24932,N_15619,N_19708);
and U24933 (N_24933,N_16908,N_16961);
nand U24934 (N_24934,N_15028,N_15523);
and U24935 (N_24935,N_18255,N_16144);
xnor U24936 (N_24936,N_18451,N_15740);
or U24937 (N_24937,N_17967,N_18128);
nand U24938 (N_24938,N_19427,N_15954);
or U24939 (N_24939,N_17729,N_17967);
and U24940 (N_24940,N_18947,N_19063);
and U24941 (N_24941,N_18249,N_18428);
nor U24942 (N_24942,N_16315,N_15058);
and U24943 (N_24943,N_15731,N_15073);
and U24944 (N_24944,N_16090,N_18912);
or U24945 (N_24945,N_18840,N_18371);
nand U24946 (N_24946,N_16617,N_15866);
nand U24947 (N_24947,N_18395,N_19213);
xor U24948 (N_24948,N_18047,N_18410);
nand U24949 (N_24949,N_15793,N_18015);
nand U24950 (N_24950,N_18844,N_17688);
or U24951 (N_24951,N_16380,N_19053);
or U24952 (N_24952,N_17778,N_16819);
and U24953 (N_24953,N_15280,N_19281);
xnor U24954 (N_24954,N_18210,N_16804);
or U24955 (N_24955,N_18246,N_15466);
xor U24956 (N_24956,N_16762,N_17560);
nand U24957 (N_24957,N_17541,N_19776);
nand U24958 (N_24958,N_17325,N_19587);
xnor U24959 (N_24959,N_18107,N_17350);
and U24960 (N_24960,N_17290,N_19387);
and U24961 (N_24961,N_17225,N_17380);
or U24962 (N_24962,N_17096,N_15129);
and U24963 (N_24963,N_19735,N_17137);
and U24964 (N_24964,N_18350,N_16607);
nor U24965 (N_24965,N_19886,N_16758);
nor U24966 (N_24966,N_17199,N_16116);
xnor U24967 (N_24967,N_19236,N_15569);
and U24968 (N_24968,N_19803,N_18553);
nor U24969 (N_24969,N_19530,N_18550);
xnor U24970 (N_24970,N_17048,N_17102);
and U24971 (N_24971,N_19790,N_19570);
and U24972 (N_24972,N_15910,N_16995);
nand U24973 (N_24973,N_16684,N_19338);
nor U24974 (N_24974,N_15563,N_16074);
xnor U24975 (N_24975,N_19958,N_17907);
nand U24976 (N_24976,N_18398,N_18312);
and U24977 (N_24977,N_18378,N_15740);
or U24978 (N_24978,N_19671,N_15298);
nand U24979 (N_24979,N_15620,N_18185);
nand U24980 (N_24980,N_19295,N_18341);
and U24981 (N_24981,N_17898,N_16770);
xor U24982 (N_24982,N_16797,N_19226);
xnor U24983 (N_24983,N_18032,N_15156);
xor U24984 (N_24984,N_18868,N_15504);
and U24985 (N_24985,N_16376,N_18519);
nor U24986 (N_24986,N_19080,N_19293);
xor U24987 (N_24987,N_15945,N_15908);
xor U24988 (N_24988,N_19963,N_18820);
or U24989 (N_24989,N_18082,N_15931);
nand U24990 (N_24990,N_19869,N_19060);
or U24991 (N_24991,N_18512,N_15783);
nor U24992 (N_24992,N_19920,N_17385);
xnor U24993 (N_24993,N_17408,N_18416);
nand U24994 (N_24994,N_19296,N_16075);
and U24995 (N_24995,N_15168,N_16057);
or U24996 (N_24996,N_17403,N_19021);
and U24997 (N_24997,N_17200,N_15554);
nand U24998 (N_24998,N_17485,N_19834);
and U24999 (N_24999,N_17697,N_17918);
nand U25000 (N_25000,N_24415,N_22145);
nand U25001 (N_25001,N_23877,N_22688);
nand U25002 (N_25002,N_24474,N_24788);
xnor U25003 (N_25003,N_23338,N_22291);
or U25004 (N_25004,N_23734,N_20953);
xor U25005 (N_25005,N_21822,N_24041);
nor U25006 (N_25006,N_23359,N_21751);
nor U25007 (N_25007,N_24727,N_20160);
nand U25008 (N_25008,N_24908,N_21576);
xor U25009 (N_25009,N_24501,N_23149);
xnor U25010 (N_25010,N_21375,N_21189);
xnor U25011 (N_25011,N_24375,N_24005);
xor U25012 (N_25012,N_23876,N_23249);
and U25013 (N_25013,N_21111,N_21711);
nand U25014 (N_25014,N_21546,N_22026);
and U25015 (N_25015,N_21473,N_23054);
nand U25016 (N_25016,N_22254,N_20435);
and U25017 (N_25017,N_24113,N_21979);
xnor U25018 (N_25018,N_24530,N_23069);
xnor U25019 (N_25019,N_21208,N_20502);
or U25020 (N_25020,N_23691,N_23158);
or U25021 (N_25021,N_22125,N_22903);
nand U25022 (N_25022,N_21112,N_23469);
xor U25023 (N_25023,N_20971,N_23942);
xor U25024 (N_25024,N_23741,N_23148);
nor U25025 (N_25025,N_21191,N_20774);
nor U25026 (N_25026,N_21517,N_21521);
and U25027 (N_25027,N_23414,N_22520);
nor U25028 (N_25028,N_22282,N_20475);
nor U25029 (N_25029,N_20198,N_24196);
nor U25030 (N_25030,N_21004,N_21176);
and U25031 (N_25031,N_24019,N_22032);
or U25032 (N_25032,N_21050,N_22694);
nand U25033 (N_25033,N_20426,N_20122);
nor U25034 (N_25034,N_23535,N_21626);
and U25035 (N_25035,N_22861,N_22430);
xor U25036 (N_25036,N_20724,N_24440);
nor U25037 (N_25037,N_20617,N_23531);
xnor U25038 (N_25038,N_20811,N_21725);
nand U25039 (N_25039,N_21833,N_21364);
nand U25040 (N_25040,N_24146,N_21409);
and U25041 (N_25041,N_23366,N_21424);
nand U25042 (N_25042,N_21075,N_20392);
xnor U25043 (N_25043,N_23233,N_23996);
nor U25044 (N_25044,N_22314,N_21748);
nand U25045 (N_25045,N_23790,N_24292);
nand U25046 (N_25046,N_20308,N_23908);
and U25047 (N_25047,N_24890,N_22793);
nor U25048 (N_25048,N_22416,N_24081);
nand U25049 (N_25049,N_20894,N_23228);
nor U25050 (N_25050,N_20587,N_21228);
and U25051 (N_25051,N_24746,N_23435);
nor U25052 (N_25052,N_21824,N_21720);
nand U25053 (N_25053,N_22894,N_24793);
xor U25054 (N_25054,N_23413,N_20937);
xnor U25055 (N_25055,N_22806,N_24248);
nor U25056 (N_25056,N_20567,N_24770);
or U25057 (N_25057,N_23291,N_24157);
or U25058 (N_25058,N_24026,N_24713);
xnor U25059 (N_25059,N_20700,N_21604);
xnor U25060 (N_25060,N_23756,N_24278);
or U25061 (N_25061,N_24227,N_22042);
or U25062 (N_25062,N_21193,N_21128);
xor U25063 (N_25063,N_24955,N_21988);
xor U25064 (N_25064,N_21454,N_21172);
xor U25065 (N_25065,N_22983,N_24650);
xnor U25066 (N_25066,N_20648,N_21919);
nor U25067 (N_25067,N_20450,N_24862);
and U25068 (N_25068,N_24074,N_22098);
nor U25069 (N_25069,N_23923,N_21257);
and U25070 (N_25070,N_22030,N_21837);
and U25071 (N_25071,N_20695,N_21280);
nand U25072 (N_25072,N_20682,N_22900);
xor U25073 (N_25073,N_20792,N_22485);
and U25074 (N_25074,N_21844,N_21887);
nand U25075 (N_25075,N_22186,N_22874);
nor U25076 (N_25076,N_22528,N_22243);
and U25077 (N_25077,N_22075,N_20874);
nand U25078 (N_25078,N_20009,N_20202);
and U25079 (N_25079,N_22493,N_24023);
xnor U25080 (N_25080,N_21689,N_22086);
nor U25081 (N_25081,N_21461,N_24328);
nand U25082 (N_25082,N_20224,N_22322);
xnor U25083 (N_25083,N_21382,N_20904);
nor U25084 (N_25084,N_22035,N_21943);
nor U25085 (N_25085,N_22572,N_22500);
xnor U25086 (N_25086,N_20654,N_23855);
nor U25087 (N_25087,N_22608,N_20522);
nand U25088 (N_25088,N_21595,N_22933);
or U25089 (N_25089,N_23809,N_22206);
and U25090 (N_25090,N_23255,N_24138);
xnor U25091 (N_25091,N_23608,N_20118);
or U25092 (N_25092,N_24166,N_24472);
nor U25093 (N_25093,N_23169,N_24006);
or U25094 (N_25094,N_20425,N_21810);
xnor U25095 (N_25095,N_22686,N_23552);
xnor U25096 (N_25096,N_22061,N_24496);
or U25097 (N_25097,N_21707,N_22696);
nor U25098 (N_25098,N_23819,N_20399);
or U25099 (N_25099,N_20145,N_22454);
xor U25100 (N_25100,N_20280,N_22594);
nand U25101 (N_25101,N_21868,N_24695);
xor U25102 (N_25102,N_24542,N_23580);
or U25103 (N_25103,N_24266,N_21638);
nor U25104 (N_25104,N_20102,N_24819);
xnor U25105 (N_25105,N_21873,N_20529);
and U25106 (N_25106,N_20422,N_24447);
xnor U25107 (N_25107,N_23928,N_23579);
nand U25108 (N_25108,N_20732,N_20839);
or U25109 (N_25109,N_20570,N_24580);
nor U25110 (N_25110,N_23938,N_20593);
nor U25111 (N_25111,N_24810,N_23289);
xor U25112 (N_25112,N_24981,N_22825);
xnor U25113 (N_25113,N_21410,N_23418);
nor U25114 (N_25114,N_21324,N_21616);
nand U25115 (N_25115,N_23119,N_20469);
nand U25116 (N_25116,N_23379,N_22810);
or U25117 (N_25117,N_20061,N_23128);
xnor U25118 (N_25118,N_24611,N_20048);
xnor U25119 (N_25119,N_23680,N_20622);
or U25120 (N_25120,N_23464,N_20833);
and U25121 (N_25121,N_22490,N_20060);
or U25122 (N_25122,N_20201,N_23684);
xnor U25123 (N_25123,N_24426,N_20794);
nor U25124 (N_25124,N_23770,N_22220);
nor U25125 (N_25125,N_20349,N_24619);
xnor U25126 (N_25126,N_21483,N_23393);
nor U25127 (N_25127,N_20492,N_24025);
nand U25128 (N_25128,N_24599,N_24556);
and U25129 (N_25129,N_23997,N_21828);
nand U25130 (N_25130,N_20560,N_24978);
nor U25131 (N_25131,N_23925,N_23163);
and U25132 (N_25132,N_24697,N_21683);
and U25133 (N_25133,N_23150,N_21073);
or U25134 (N_25134,N_20454,N_22025);
nand U25135 (N_25135,N_23104,N_24263);
or U25136 (N_25136,N_22105,N_24105);
and U25137 (N_25137,N_20550,N_22928);
nor U25138 (N_25138,N_23428,N_24976);
xnor U25139 (N_25139,N_22187,N_20059);
nor U25140 (N_25140,N_23664,N_20310);
nand U25141 (N_25141,N_20443,N_20188);
and U25142 (N_25142,N_24178,N_23159);
and U25143 (N_25143,N_21853,N_20672);
xor U25144 (N_25144,N_23761,N_22228);
and U25145 (N_25145,N_23698,N_21766);
nor U25146 (N_25146,N_20505,N_21763);
xnor U25147 (N_25147,N_24336,N_24099);
nor U25148 (N_25148,N_24691,N_20026);
and U25149 (N_25149,N_22400,N_23872);
nand U25150 (N_25150,N_20736,N_24092);
and U25151 (N_25151,N_24709,N_20050);
nand U25152 (N_25152,N_22702,N_20781);
and U25153 (N_25153,N_22636,N_24271);
nand U25154 (N_25154,N_21599,N_23179);
nor U25155 (N_25155,N_20286,N_24313);
xor U25156 (N_25156,N_20271,N_22309);
or U25157 (N_25157,N_22440,N_21437);
and U25158 (N_25158,N_24663,N_21605);
or U25159 (N_25159,N_21404,N_23225);
nand U25160 (N_25160,N_20565,N_22175);
nand U25161 (N_25161,N_20254,N_21644);
or U25162 (N_25162,N_22104,N_22555);
nand U25163 (N_25163,N_20782,N_24549);
xor U25164 (N_25164,N_21515,N_20658);
nor U25165 (N_25165,N_23893,N_21484);
or U25166 (N_25166,N_22567,N_24298);
xor U25167 (N_25167,N_22837,N_20184);
or U25168 (N_25168,N_23871,N_24429);
xnor U25169 (N_25169,N_23144,N_21817);
nand U25170 (N_25170,N_24480,N_22516);
or U25171 (N_25171,N_24555,N_22634);
xnor U25172 (N_25172,N_22359,N_22022);
nand U25173 (N_25173,N_24965,N_24735);
xnor U25174 (N_25174,N_20449,N_23114);
or U25175 (N_25175,N_22496,N_21938);
nand U25176 (N_25176,N_20631,N_20734);
or U25177 (N_25177,N_23205,N_22611);
nand U25178 (N_25178,N_21504,N_24806);
nor U25179 (N_25179,N_20600,N_20663);
nand U25180 (N_25180,N_20333,N_21964);
nor U25181 (N_25181,N_21124,N_22705);
nand U25182 (N_25182,N_24596,N_24646);
nand U25183 (N_25183,N_20723,N_22949);
xnor U25184 (N_25184,N_23306,N_22934);
xnor U25185 (N_25185,N_21487,N_23007);
nor U25186 (N_25186,N_24906,N_24783);
nor U25187 (N_25187,N_24868,N_24486);
nand U25188 (N_25188,N_21586,N_22327);
xor U25189 (N_25189,N_22531,N_23536);
and U25190 (N_25190,N_22501,N_20907);
or U25191 (N_25191,N_22950,N_21282);
xnor U25192 (N_25192,N_21806,N_23351);
and U25193 (N_25193,N_20192,N_24710);
nand U25194 (N_25194,N_21167,N_21922);
and U25195 (N_25195,N_21033,N_23096);
xor U25196 (N_25196,N_22910,N_22449);
or U25197 (N_25197,N_20068,N_22722);
xor U25198 (N_25198,N_22564,N_22877);
xnor U25199 (N_25199,N_22947,N_20287);
nor U25200 (N_25200,N_23695,N_24389);
or U25201 (N_25201,N_23548,N_23426);
xor U25202 (N_25202,N_23669,N_20042);
nand U25203 (N_25203,N_21365,N_20390);
or U25204 (N_25204,N_24944,N_22732);
nor U25205 (N_25205,N_23355,N_21910);
xnor U25206 (N_25206,N_23406,N_23105);
and U25207 (N_25207,N_24667,N_24644);
and U25208 (N_25208,N_20126,N_24737);
or U25209 (N_25209,N_20519,N_22563);
or U25210 (N_25210,N_21195,N_24229);
xnor U25211 (N_25211,N_22411,N_21314);
and U25212 (N_25212,N_23701,N_22492);
or U25213 (N_25213,N_22519,N_20710);
and U25214 (N_25214,N_20470,N_20761);
nor U25215 (N_25215,N_23875,N_23717);
and U25216 (N_25216,N_24563,N_22794);
and U25217 (N_25217,N_24467,N_20832);
or U25218 (N_25218,N_24362,N_22968);
nand U25219 (N_25219,N_22617,N_20609);
nand U25220 (N_25220,N_23389,N_20787);
and U25221 (N_25221,N_21390,N_21603);
or U25222 (N_25222,N_20234,N_24546);
nor U25223 (N_25223,N_24463,N_20244);
nand U25224 (N_25224,N_23972,N_21043);
or U25225 (N_25225,N_21264,N_20455);
nand U25226 (N_25226,N_22362,N_21042);
nand U25227 (N_25227,N_20708,N_20571);
or U25228 (N_25228,N_23018,N_21578);
or U25229 (N_25229,N_24648,N_22164);
nor U25230 (N_25230,N_24679,N_24291);
nor U25231 (N_25231,N_24384,N_24121);
nor U25232 (N_25232,N_24618,N_24791);
nand U25233 (N_25233,N_22737,N_21518);
or U25234 (N_25234,N_20152,N_23222);
and U25235 (N_25235,N_24488,N_20662);
nor U25236 (N_25236,N_22868,N_21442);
and U25237 (N_25237,N_24593,N_20642);
nand U25238 (N_25238,N_23482,N_24464);
nor U25239 (N_25239,N_23374,N_23458);
nor U25240 (N_25240,N_24883,N_20999);
or U25241 (N_25241,N_20985,N_21832);
xor U25242 (N_25242,N_22799,N_20778);
xnor U25243 (N_25243,N_23141,N_21547);
nand U25244 (N_25244,N_24854,N_21165);
or U25245 (N_25245,N_21669,N_21597);
nor U25246 (N_25246,N_20934,N_24111);
or U25247 (N_25247,N_20072,N_24012);
xnor U25248 (N_25248,N_22180,N_21447);
or U25249 (N_25249,N_23600,N_21584);
and U25250 (N_25250,N_21859,N_22899);
nand U25251 (N_25251,N_21175,N_20910);
nand U25252 (N_25252,N_22885,N_23612);
nand U25253 (N_25253,N_22556,N_23733);
or U25254 (N_25254,N_21846,N_24327);
and U25255 (N_25255,N_21237,N_24176);
xnor U25256 (N_25256,N_23283,N_21946);
xnor U25257 (N_25257,N_22007,N_21631);
nor U25258 (N_25258,N_20367,N_23738);
nand U25259 (N_25259,N_22370,N_23280);
or U25260 (N_25260,N_22819,N_21592);
nand U25261 (N_25261,N_20618,N_23318);
and U25262 (N_25262,N_20339,N_22859);
nor U25263 (N_25263,N_23848,N_20191);
xor U25264 (N_25264,N_20484,N_21655);
or U25265 (N_25265,N_22984,N_22606);
nand U25266 (N_25266,N_24149,N_21642);
nand U25267 (N_25267,N_21700,N_24889);
and U25268 (N_25268,N_21322,N_22985);
nand U25269 (N_25269,N_23815,N_21607);
nor U25270 (N_25270,N_22203,N_24846);
nor U25271 (N_25271,N_22541,N_23257);
nand U25272 (N_25272,N_21855,N_21850);
nand U25273 (N_25273,N_20235,N_22585);
xor U25274 (N_25274,N_23880,N_21090);
and U25275 (N_25275,N_23879,N_20405);
nand U25276 (N_25276,N_21975,N_23336);
nand U25277 (N_25277,N_24969,N_23013);
xnor U25278 (N_25278,N_22927,N_22614);
or U25279 (N_25279,N_22765,N_21265);
and U25280 (N_25280,N_22252,N_24030);
and U25281 (N_25281,N_22162,N_24475);
or U25282 (N_25282,N_23475,N_23826);
and U25283 (N_25283,N_20967,N_21746);
nand U25284 (N_25284,N_24289,N_21106);
nand U25285 (N_25285,N_24855,N_22919);
and U25286 (N_25286,N_21849,N_24990);
nor U25287 (N_25287,N_22082,N_21469);
xor U25288 (N_25288,N_24010,N_21559);
nand U25289 (N_25289,N_23345,N_22641);
or U25290 (N_25290,N_22467,N_24346);
nand U25291 (N_25291,N_23486,N_23164);
and U25292 (N_25292,N_22160,N_21434);
xnor U25293 (N_25293,N_23040,N_24022);
nand U25294 (N_25294,N_21378,N_22721);
and U25295 (N_25295,N_24168,N_23248);
xor U25296 (N_25296,N_23705,N_21884);
and U25297 (N_25297,N_21289,N_20421);
nor U25298 (N_25298,N_23610,N_23713);
nor U25299 (N_25299,N_20942,N_24787);
xor U25300 (N_25300,N_20686,N_23524);
nor U25301 (N_25301,N_22747,N_23951);
xnor U25302 (N_25302,N_24071,N_20278);
xnor U25303 (N_25303,N_20326,N_22211);
xor U25304 (N_25304,N_20961,N_24772);
or U25305 (N_25305,N_20900,N_24562);
xnor U25306 (N_25306,N_23181,N_24274);
or U25307 (N_25307,N_21180,N_24932);
nor U25308 (N_25308,N_20429,N_22225);
nor U25309 (N_25309,N_20984,N_20580);
nor U25310 (N_25310,N_24213,N_21630);
or U25311 (N_25311,N_23990,N_23562);
and U25312 (N_25312,N_21869,N_21357);
nor U25313 (N_25313,N_24342,N_22959);
nand U25314 (N_25314,N_22194,N_21009);
xnor U25315 (N_25315,N_21952,N_22452);
nand U25316 (N_25316,N_22615,N_22196);
nor U25317 (N_25317,N_23699,N_21227);
nand U25318 (N_25318,N_21932,N_20613);
xnor U25319 (N_25319,N_21119,N_20574);
xnor U25320 (N_25320,N_20474,N_23711);
nand U25321 (N_25321,N_24171,N_22420);
and U25322 (N_25322,N_23491,N_23005);
or U25323 (N_25323,N_20065,N_24043);
or U25324 (N_25324,N_24355,N_24350);
and U25325 (N_25325,N_20211,N_21976);
and U25326 (N_25326,N_21475,N_20989);
nand U25327 (N_25327,N_20705,N_20836);
or U25328 (N_25328,N_22616,N_24454);
nor U25329 (N_25329,N_23596,N_22404);
nor U25330 (N_25330,N_23939,N_21897);
and U25331 (N_25331,N_24308,N_23934);
nor U25332 (N_25332,N_21027,N_22354);
or U25333 (N_25333,N_20243,N_24803);
xor U25334 (N_25334,N_21657,N_21980);
nor U25335 (N_25335,N_20979,N_20362);
and U25336 (N_25336,N_24239,N_20114);
and U25337 (N_25337,N_21541,N_22149);
or U25338 (N_25338,N_20269,N_20824);
nand U25339 (N_25339,N_21594,N_22808);
nor U25340 (N_25340,N_24802,N_24095);
nor U25341 (N_25341,N_24377,N_21104);
or U25342 (N_25342,N_20886,N_21813);
nor U25343 (N_25343,N_21637,N_24400);
or U25344 (N_25344,N_21336,N_24469);
nor U25345 (N_25345,N_24079,N_23341);
and U25346 (N_25346,N_21934,N_21889);
nand U25347 (N_25347,N_23403,N_20226);
xnor U25348 (N_25348,N_23811,N_23948);
xnor U25349 (N_25349,N_22391,N_21318);
nor U25350 (N_25350,N_20078,N_23259);
nor U25351 (N_25351,N_23116,N_20849);
nor U25352 (N_25352,N_23440,N_24804);
and U25353 (N_25353,N_22752,N_22860);
xnor U25354 (N_25354,N_23687,N_21574);
or U25355 (N_25355,N_24337,N_21781);
nand U25356 (N_25356,N_23207,N_23287);
xor U25357 (N_25357,N_21163,N_20557);
xnor U25358 (N_25358,N_21298,N_21005);
xor U25359 (N_25359,N_21590,N_24117);
xnor U25360 (N_25360,N_21466,N_20847);
or U25361 (N_25361,N_20891,N_23945);
and U25362 (N_25362,N_24624,N_22476);
nand U25363 (N_25363,N_24391,N_21092);
nand U25364 (N_25364,N_23613,N_20780);
nor U25365 (N_25365,N_23549,N_24869);
or U25366 (N_25366,N_24632,N_22855);
and U25367 (N_25367,N_24756,N_21639);
or U25368 (N_25368,N_24905,N_23586);
xnor U25369 (N_25369,N_21963,N_24054);
or U25370 (N_25370,N_21118,N_23523);
and U25371 (N_25371,N_22642,N_20924);
nand U25372 (N_25372,N_22648,N_23172);
nor U25373 (N_25373,N_20249,N_22344);
or U25374 (N_25374,N_22505,N_23450);
nor U25375 (N_25375,N_23268,N_24093);
nand U25376 (N_25376,N_23299,N_23512);
nor U25377 (N_25377,N_24921,N_20706);
nor U25378 (N_25378,N_20892,N_20501);
xnor U25379 (N_25379,N_22509,N_20846);
or U25380 (N_25380,N_22851,N_23437);
or U25381 (N_25381,N_21877,N_24064);
nand U25382 (N_25382,N_24161,N_20598);
and U25383 (N_25383,N_23505,N_20670);
nor U25384 (N_25384,N_23739,N_20744);
xor U25385 (N_25385,N_23391,N_24876);
and U25386 (N_25386,N_23852,N_24568);
nor U25387 (N_25387,N_20840,N_20177);
or U25388 (N_25388,N_22037,N_23653);
nand U25389 (N_25389,N_21712,N_24056);
xor U25390 (N_25390,N_20452,N_21350);
and U25391 (N_25391,N_21393,N_24148);
xor U25392 (N_25392,N_22540,N_24661);
or U25393 (N_25393,N_24107,N_22770);
xnor U25394 (N_25394,N_23585,N_20854);
xnor U25395 (N_25395,N_24143,N_20759);
nand U25396 (N_25396,N_22392,N_20796);
xnor U25397 (N_25397,N_23642,N_20375);
and U25398 (N_25398,N_22174,N_23165);
and U25399 (N_25399,N_23075,N_21485);
nor U25400 (N_25400,N_21166,N_21463);
nor U25401 (N_25401,N_22117,N_21694);
xnor U25402 (N_25402,N_24425,N_22723);
or U25403 (N_25403,N_24812,N_20116);
and U25404 (N_25404,N_20301,N_22931);
and U25405 (N_25405,N_23550,N_22464);
or U25406 (N_25406,N_20229,N_22631);
nand U25407 (N_25407,N_22446,N_24280);
or U25408 (N_25408,N_21338,N_22693);
xor U25409 (N_25409,N_23860,N_24768);
and U25410 (N_25410,N_22473,N_20966);
nand U25411 (N_25411,N_22862,N_20941);
and U25412 (N_25412,N_24457,N_23750);
and U25413 (N_25413,N_21526,N_23060);
xor U25414 (N_25414,N_24943,N_21714);
or U25415 (N_25415,N_23079,N_24027);
or U25416 (N_25416,N_20728,N_24964);
nand U25417 (N_25417,N_23762,N_24703);
or U25418 (N_25418,N_22229,N_22951);
and U25419 (N_25419,N_23218,N_23369);
nor U25420 (N_25420,N_23131,N_20380);
or U25421 (N_25421,N_22690,N_24021);
xor U25422 (N_25422,N_20094,N_20534);
nor U25423 (N_25423,N_23728,N_24655);
xor U25424 (N_25424,N_21958,N_21617);
xor U25425 (N_25425,N_24204,N_21241);
and U25426 (N_25426,N_23385,N_22457);
and U25427 (N_25427,N_20685,N_23873);
nor U25428 (N_25428,N_22118,N_24140);
or U25429 (N_25429,N_21990,N_21088);
nor U25430 (N_25430,N_23296,N_22973);
xnor U25431 (N_25431,N_21396,N_23365);
xnor U25432 (N_25432,N_23627,N_22909);
or U25433 (N_25433,N_23793,N_21293);
or U25434 (N_25434,N_23139,N_22077);
or U25435 (N_25435,N_24642,N_21986);
nand U25436 (N_25436,N_21593,N_21676);
and U25437 (N_25437,N_24075,N_22646);
xor U25438 (N_25438,N_22898,N_22155);
xor U25439 (N_25439,N_21588,N_24189);
xnor U25440 (N_25440,N_21372,N_24323);
and U25441 (N_25441,N_20751,N_20101);
xor U25442 (N_25442,N_22880,N_23102);
nand U25443 (N_25443,N_23618,N_24134);
or U25444 (N_25444,N_22198,N_22332);
or U25445 (N_25445,N_24347,N_22286);
and U25446 (N_25446,N_21544,N_23814);
nor U25447 (N_25447,N_20197,N_21621);
and U25448 (N_25448,N_23936,N_22726);
xor U25449 (N_25449,N_23161,N_22589);
xnor U25450 (N_25450,N_24476,N_22432);
nor U25451 (N_25451,N_22137,N_21784);
or U25452 (N_25452,N_20412,N_20921);
nand U25453 (N_25453,N_23722,N_22768);
nor U25454 (N_25454,N_22970,N_20493);
nor U25455 (N_25455,N_23850,N_22447);
nor U25456 (N_25456,N_20901,N_20216);
or U25457 (N_25457,N_20625,N_22188);
xor U25458 (N_25458,N_22495,N_24759);
nor U25459 (N_25459,N_22330,N_24706);
and U25460 (N_25460,N_20097,N_21558);
and U25461 (N_25461,N_23748,N_23603);
and U25462 (N_25462,N_20917,N_23078);
xnor U25463 (N_25463,N_24898,N_21087);
and U25464 (N_25464,N_20079,N_20318);
nand U25465 (N_25465,N_21506,N_23332);
xnor U25466 (N_25466,N_21779,N_22444);
xnor U25467 (N_25467,N_24369,N_21993);
or U25468 (N_25468,N_20540,N_20853);
and U25469 (N_25469,N_21039,N_23746);
nand U25470 (N_25470,N_21602,N_24966);
xor U25471 (N_25471,N_24462,N_20981);
nand U25472 (N_25472,N_21343,N_22895);
and U25473 (N_25473,N_24660,N_20543);
or U25474 (N_25474,N_20081,N_21472);
nor U25475 (N_25475,N_22121,N_21381);
xnor U25476 (N_25476,N_23375,N_21827);
and U25477 (N_25477,N_20935,N_21749);
or U25478 (N_25478,N_23087,N_20976);
xnor U25479 (N_25479,N_22337,N_21493);
nand U25480 (N_25480,N_22853,N_24009);
or U25481 (N_25481,N_23381,N_20005);
or U25482 (N_25482,N_24576,N_21913);
and U25483 (N_25483,N_21908,N_21764);
and U25484 (N_25484,N_22664,N_21918);
or U25485 (N_25485,N_22256,N_21505);
nand U25486 (N_25486,N_20204,N_23492);
and U25487 (N_25487,N_20164,N_22466);
nor U25488 (N_25488,N_24985,N_24282);
or U25489 (N_25489,N_24181,N_24318);
nor U25490 (N_25490,N_22275,N_20518);
nand U25491 (N_25491,N_23726,N_24088);
and U25492 (N_25492,N_21462,N_23224);
or U25493 (N_25493,N_20875,N_20753);
nand U25494 (N_25494,N_23666,N_22321);
xnor U25495 (N_25495,N_23769,N_24512);
or U25496 (N_25496,N_23476,N_21174);
or U25497 (N_25497,N_24749,N_21852);
and U25498 (N_25498,N_21535,N_20297);
and U25499 (N_25499,N_21534,N_24687);
and U25500 (N_25500,N_23641,N_24891);
nand U25501 (N_25501,N_21168,N_22255);
nor U25502 (N_25502,N_21701,N_20649);
and U25503 (N_25503,N_21150,N_21368);
or U25504 (N_25504,N_22475,N_21178);
nand U25505 (N_25505,N_24996,N_23663);
xor U25506 (N_25506,N_21086,N_24719);
and U25507 (N_25507,N_21640,N_24948);
nand U25508 (N_25508,N_24760,N_23584);
nand U25509 (N_25509,N_22315,N_24485);
nand U25510 (N_25510,N_24594,N_22792);
nand U25511 (N_25511,N_22913,N_24640);
or U25512 (N_25512,N_22021,N_24158);
nor U25513 (N_25513,N_23979,N_21937);
nor U25514 (N_25514,N_23964,N_21693);
nor U25515 (N_25515,N_22639,N_21614);
or U25516 (N_25516,N_20814,N_23574);
nor U25517 (N_25517,N_20456,N_22384);
and U25518 (N_25518,N_24607,N_24960);
or U25519 (N_25519,N_21263,N_24139);
and U25520 (N_25520,N_21507,N_23985);
nor U25521 (N_25521,N_21840,N_22834);
and U25522 (N_25522,N_22039,N_24110);
and U25523 (N_25523,N_21071,N_24982);
nor U25524 (N_25524,N_20641,N_24728);
nor U25525 (N_25525,N_21113,N_20135);
xor U25526 (N_25526,N_22352,N_24106);
nor U25527 (N_25527,N_22907,N_24567);
or U25528 (N_25528,N_23667,N_21863);
and U25529 (N_25529,N_23045,N_20170);
xor U25530 (N_25530,N_23329,N_20461);
or U25531 (N_25531,N_21745,N_20620);
or U25532 (N_25532,N_23753,N_21223);
nand U25533 (N_25533,N_24209,N_23787);
xnor U25534 (N_25534,N_20646,N_21194);
xnor U25535 (N_25535,N_22715,N_24917);
and U25536 (N_25536,N_24682,N_23833);
nand U25537 (N_25537,N_23136,N_21330);
or U25538 (N_25538,N_20684,N_23417);
and U25539 (N_25539,N_23842,N_22340);
or U25540 (N_25540,N_23906,N_22578);
nand U25541 (N_25541,N_24351,N_22980);
nand U25542 (N_25542,N_20496,N_23661);
nor U25543 (N_25543,N_23969,N_24717);
and U25544 (N_25544,N_20800,N_22011);
or U25545 (N_25545,N_23589,N_20596);
xnor U25546 (N_25546,N_23166,N_24344);
or U25547 (N_25547,N_23242,N_21554);
nor U25548 (N_25548,N_22748,N_23020);
nor U25549 (N_25549,N_23083,N_23773);
and U25550 (N_25550,N_21416,N_21094);
or U25551 (N_25551,N_21570,N_24073);
nor U25552 (N_25552,N_24875,N_22057);
xnor U25553 (N_25553,N_20210,N_23940);
nand U25554 (N_25554,N_22016,N_23168);
or U25555 (N_25555,N_20187,N_24299);
nor U25556 (N_25556,N_20987,N_23333);
and U25557 (N_25557,N_22991,N_24780);
nand U25558 (N_25558,N_20194,N_23189);
or U25559 (N_25559,N_24468,N_23834);
nor U25560 (N_25560,N_23958,N_21177);
nor U25561 (N_25561,N_23174,N_22633);
nand U25562 (N_25562,N_23794,N_20877);
and U25563 (N_25563,N_23595,N_22213);
nor U25564 (N_25564,N_23122,N_20623);
nor U25565 (N_25565,N_23614,N_24002);
nor U25566 (N_25566,N_20148,N_23583);
and U25567 (N_25567,N_24294,N_21083);
xor U25568 (N_25568,N_24484,N_20413);
and U25569 (N_25569,N_21994,N_24101);
and U25570 (N_25570,N_20986,N_21315);
or U25571 (N_25571,N_22356,N_22856);
nand U25572 (N_25572,N_21864,N_22857);
nor U25573 (N_25573,N_21320,N_24823);
xor U25574 (N_25574,N_20944,N_22609);
xnor U25575 (N_25575,N_24954,N_24664);
or U25576 (N_25576,N_20324,N_23448);
nor U25577 (N_25577,N_20215,N_23196);
xnor U25578 (N_25578,N_22300,N_24638);
nor U25579 (N_25579,N_21305,N_22761);
and U25580 (N_25580,N_20758,N_20312);
nand U25581 (N_25581,N_22258,N_20905);
nor U25582 (N_25582,N_20279,N_24431);
and U25583 (N_25583,N_21871,N_23547);
xor U25584 (N_25584,N_24226,N_22130);
or U25585 (N_25585,N_21432,N_24828);
or U25586 (N_25586,N_23137,N_21481);
xnor U25587 (N_25587,N_23694,N_24201);
xor U25588 (N_25588,N_24950,N_23619);
xor U25589 (N_25589,N_21252,N_23671);
nand U25590 (N_25590,N_20980,N_22650);
xnor U25591 (N_25591,N_23543,N_22489);
or U25592 (N_25592,N_21120,N_21007);
or U25593 (N_25593,N_21865,N_24242);
nand U25594 (N_25594,N_21736,N_21894);
or U25595 (N_25595,N_22524,N_23513);
xnor U25596 (N_25596,N_21609,N_22292);
or U25597 (N_25597,N_20494,N_23796);
or U25598 (N_25598,N_23922,N_20092);
xor U25599 (N_25599,N_24532,N_24290);
nor U25600 (N_25600,N_24058,N_23777);
nor U25601 (N_25601,N_20504,N_21718);
nand U25602 (N_25602,N_22944,N_23974);
nor U25603 (N_25603,N_23266,N_20487);
nor U25604 (N_25604,N_21591,N_24283);
or U25605 (N_25605,N_20605,N_20052);
nor U25606 (N_25606,N_22844,N_22525);
xor U25607 (N_25607,N_20742,N_24877);
xnor U25608 (N_25608,N_20028,N_24919);
nand U25609 (N_25609,N_23707,N_20694);
or U25610 (N_25610,N_21508,N_21903);
and U25611 (N_25611,N_20325,N_21199);
nand U25612 (N_25612,N_21201,N_21105);
or U25613 (N_25613,N_21830,N_22461);
and U25614 (N_25614,N_24609,N_23643);
nand U25615 (N_25615,N_21311,N_22724);
nand U25616 (N_25616,N_20701,N_20711);
and U25617 (N_25617,N_24137,N_23363);
and U25618 (N_25618,N_23519,N_22550);
and U25619 (N_25619,N_24152,N_21465);
and U25620 (N_25620,N_20797,N_21303);
or U25621 (N_25621,N_24370,N_20909);
nor U25622 (N_25622,N_23481,N_20992);
or U25623 (N_25623,N_23412,N_21213);
nor U25624 (N_25624,N_20586,N_20964);
nand U25625 (N_25625,N_24032,N_21956);
nor U25626 (N_25626,N_20186,N_20532);
xor U25627 (N_25627,N_22080,N_21829);
or U25628 (N_25628,N_24957,N_22334);
or U25629 (N_25629,N_20236,N_21406);
nor U25630 (N_25630,N_21209,N_22915);
or U25631 (N_25631,N_24837,N_22735);
and U25632 (N_25632,N_24312,N_21281);
and U25633 (N_25633,N_23884,N_24592);
nor U25634 (N_25634,N_20511,N_22736);
xnor U25635 (N_25635,N_20104,N_23065);
nand U25636 (N_25636,N_24881,N_24017);
xnor U25637 (N_25637,N_23094,N_24407);
nand U25638 (N_25638,N_23957,N_23763);
nand U25639 (N_25639,N_22503,N_21279);
or U25640 (N_25640,N_20423,N_20745);
nor U25641 (N_25641,N_21924,N_20093);
nor U25642 (N_25642,N_22971,N_23836);
xor U25643 (N_25643,N_22870,N_23465);
xnor U25644 (N_25644,N_24573,N_24832);
nand U25645 (N_25645,N_22866,N_22923);
and U25646 (N_25646,N_21600,N_21397);
nor U25647 (N_25647,N_23187,N_24262);
nand U25648 (N_25648,N_22534,N_22829);
nor U25649 (N_25649,N_21878,N_24544);
and U25650 (N_25650,N_24360,N_23354);
and U25651 (N_25651,N_24471,N_23021);
nor U25652 (N_25652,N_21793,N_23843);
xor U25653 (N_25653,N_24980,N_20085);
nor U25654 (N_25654,N_24688,N_24974);
nand U25655 (N_25655,N_22365,N_22543);
or U25656 (N_25656,N_24395,N_24444);
and U25657 (N_25657,N_23474,N_22733);
nor U25658 (N_25658,N_20523,N_22902);
xor U25659 (N_25659,N_23660,N_21652);
xor U25660 (N_25660,N_23560,N_23911);
or U25661 (N_25661,N_22517,N_21349);
or U25662 (N_25662,N_20653,N_21501);
and U25663 (N_25663,N_20863,N_23208);
and U25664 (N_25664,N_23135,N_22193);
and U25665 (N_25665,N_20457,N_22271);
and U25666 (N_25666,N_24845,N_23685);
or U25667 (N_25667,N_23617,N_20881);
nand U25668 (N_25668,N_20464,N_24900);
nand U25669 (N_25669,N_23988,N_20361);
xor U25670 (N_25670,N_24551,N_20741);
or U25671 (N_25671,N_20175,N_23309);
nor U25672 (N_25672,N_23752,N_24785);
nand U25673 (N_25673,N_20247,N_20870);
nor U25674 (N_25674,N_21455,N_23310);
and U25675 (N_25675,N_21186,N_23478);
xnor U25676 (N_25676,N_21002,N_20816);
and U25677 (N_25677,N_24288,N_22238);
and U25678 (N_25678,N_22839,N_21304);
and U25679 (N_25679,N_21955,N_22560);
nor U25680 (N_25680,N_22667,N_21528);
or U25681 (N_25681,N_21140,N_21037);
or U25682 (N_25682,N_24924,N_20165);
and U25683 (N_25683,N_24224,N_24211);
or U25684 (N_25684,N_24206,N_21673);
or U25685 (N_25685,N_21055,N_24702);
nand U25686 (N_25686,N_23681,N_23837);
xnor U25687 (N_25687,N_23900,N_22434);
xnor U25688 (N_25688,N_22530,N_24169);
xnor U25689 (N_25689,N_21292,N_23910);
or U25690 (N_25690,N_20430,N_24442);
xor U25691 (N_25691,N_24163,N_22008);
nor U25692 (N_25692,N_23735,N_23278);
or U25693 (N_25693,N_21783,N_21102);
xnor U25694 (N_25694,N_24507,N_23080);
or U25695 (N_25695,N_21929,N_23064);
or U25696 (N_25696,N_22443,N_20260);
nor U25697 (N_25697,N_22831,N_21068);
nor U25698 (N_25698,N_24055,N_22601);
and U25699 (N_25699,N_22879,N_21123);
or U25700 (N_25700,N_21967,N_22976);
nor U25701 (N_25701,N_24250,N_24063);
xor U25702 (N_25702,N_20389,N_24076);
and U25703 (N_25703,N_20551,N_22964);
nor U25704 (N_25704,N_23008,N_24560);
nor U25705 (N_25705,N_20926,N_24570);
nand U25706 (N_25706,N_24062,N_21951);
or U25707 (N_25707,N_23935,N_24902);
xnor U25708 (N_25708,N_22739,N_23903);
xor U25709 (N_25709,N_22990,N_20889);
and U25710 (N_25710,N_24987,N_20100);
xor U25711 (N_25711,N_23921,N_21684);
xnor U25712 (N_25712,N_23754,N_20740);
xnor U25713 (N_25713,N_23395,N_22963);
xnor U25714 (N_25714,N_23006,N_20669);
or U25715 (N_25715,N_23443,N_21022);
or U25716 (N_25716,N_20861,N_22925);
or U25717 (N_25717,N_24123,N_23275);
and U25718 (N_25718,N_23127,N_22090);
and U25719 (N_25719,N_23262,N_24977);
and U25720 (N_25720,N_21856,N_23961);
nand U25721 (N_25721,N_22158,N_23409);
xor U25722 (N_25722,N_21224,N_20556);
xor U25723 (N_25723,N_21582,N_23024);
xor U25724 (N_25724,N_20716,N_20176);
or U25725 (N_25725,N_24896,N_20403);
and U25726 (N_25726,N_21754,N_20227);
or U25727 (N_25727,N_21622,N_22408);
xnor U25728 (N_25728,N_22378,N_22048);
nor U25729 (N_25729,N_21001,N_22612);
nand U25730 (N_25730,N_21385,N_23800);
nor U25731 (N_25731,N_22395,N_23511);
and U25732 (N_25732,N_23056,N_23704);
and U25733 (N_25733,N_20664,N_20460);
nor U25734 (N_25734,N_21867,N_20002);
and U25735 (N_25735,N_23398,N_21681);
or U25736 (N_25736,N_20095,N_23343);
and U25737 (N_25737,N_24732,N_23314);
nor U25738 (N_25738,N_22795,N_23823);
xor U25739 (N_25739,N_24261,N_23975);
nor U25740 (N_25740,N_22028,N_23235);
nand U25741 (N_25741,N_24228,N_24284);
or U25742 (N_25742,N_24967,N_20897);
and U25743 (N_25743,N_24610,N_20378);
or U25744 (N_25744,N_20099,N_21841);
nor U25745 (N_25745,N_20656,N_22656);
nor U25746 (N_25746,N_23740,N_22587);
nor U25747 (N_25747,N_20441,N_23358);
nor U25748 (N_25748,N_22103,N_24829);
nand U25749 (N_25749,N_20356,N_23125);
nor U25750 (N_25750,N_24533,N_23807);
xor U25751 (N_25751,N_24654,N_22426);
and U25752 (N_25752,N_24817,N_23180);
xor U25753 (N_25753,N_20520,N_22813);
nand U25754 (N_25754,N_24458,N_24635);
and U25755 (N_25755,N_21064,N_21323);
nand U25756 (N_25756,N_24668,N_23495);
or U25757 (N_25757,N_24840,N_22997);
or U25758 (N_25758,N_20144,N_20608);
and U25759 (N_25759,N_22746,N_20765);
nor U25760 (N_25760,N_20737,N_21904);
xor U25761 (N_25761,N_24434,N_21182);
xor U25762 (N_25762,N_22649,N_24515);
and U25763 (N_25763,N_24795,N_24813);
nand U25764 (N_25764,N_20338,N_22316);
or U25765 (N_25765,N_23858,N_24716);
nor U25766 (N_25766,N_23943,N_22202);
or U25767 (N_25767,N_20386,N_21775);
nor U25768 (N_25768,N_24264,N_20083);
or U25769 (N_25769,N_20822,N_21917);
or U25770 (N_25770,N_20112,N_24649);
nand U25771 (N_25771,N_22559,N_23886);
nor U25772 (N_25772,N_23298,N_24309);
nor U25773 (N_25773,N_22730,N_22313);
and U25774 (N_25774,N_24628,N_23261);
nor U25775 (N_25775,N_23061,N_20997);
or U25776 (N_25776,N_23506,N_22975);
nand U25777 (N_25777,N_21347,N_22527);
xor U25778 (N_25778,N_20893,N_20284);
nor U25779 (N_25779,N_20433,N_22972);
nand U25780 (N_25780,N_22629,N_24322);
nor U25781 (N_25781,N_20022,N_23319);
nor U25782 (N_25782,N_22886,N_23023);
nand U25783 (N_25783,N_23422,N_24013);
xnor U25784 (N_25784,N_20762,N_23199);
and U25785 (N_25785,N_22507,N_24489);
and U25786 (N_25786,N_23588,N_24612);
or U25787 (N_25787,N_22832,N_21231);
xor U25788 (N_25788,N_20090,N_22514);
nor U25789 (N_25789,N_23847,N_22699);
or U25790 (N_25790,N_24356,N_22569);
nor U25791 (N_25791,N_23616,N_20411);
nand U25792 (N_25792,N_23865,N_24066);
or U25793 (N_25793,N_21611,N_21870);
nor U25794 (N_25794,N_22539,N_22691);
or U25795 (N_25795,N_23710,N_24675);
xnor U25796 (N_25796,N_23736,N_23404);
or U25797 (N_25797,N_20203,N_20527);
xor U25798 (N_25798,N_21732,N_23606);
or U25799 (N_25799,N_24000,N_20573);
and U25800 (N_25800,N_23567,N_20270);
xnor U25801 (N_25801,N_21259,N_21842);
xor U25802 (N_25802,N_24397,N_24569);
nand U25803 (N_25803,N_24223,N_22427);
or U25804 (N_25804,N_21251,N_21363);
nor U25805 (N_25805,N_23601,N_22018);
and U25806 (N_25806,N_23970,N_21800);
xor U25807 (N_25807,N_20259,N_24792);
or U25808 (N_25808,N_23399,N_21847);
and U25809 (N_25809,N_20678,N_20864);
nor U25810 (N_25810,N_21317,N_21705);
xor U25811 (N_25811,N_24559,N_20045);
and U25812 (N_25812,N_24338,N_23334);
or U25813 (N_25813,N_23721,N_23479);
or U25814 (N_25814,N_22766,N_22893);
nand U25815 (N_25815,N_24069,N_22123);
and U25816 (N_25816,N_24912,N_21439);
nand U25817 (N_25817,N_21826,N_23992);
nand U25818 (N_25818,N_20978,N_23253);
nor U25819 (N_25819,N_21477,N_22122);
nand U25820 (N_25820,N_22689,N_24796);
xor U25821 (N_25821,N_22491,N_22841);
and U25822 (N_25822,N_20432,N_21218);
nor U25823 (N_25823,N_20977,N_23477);
and U25824 (N_25824,N_21095,N_23411);
and U25825 (N_25825,N_20548,N_20956);
or U25826 (N_25826,N_24084,N_20472);
and U25827 (N_25827,N_22388,N_21078);
or U25828 (N_25828,N_22287,N_21057);
xor U25829 (N_25829,N_23462,N_22661);
and U25830 (N_25830,N_21511,N_23027);
xor U25831 (N_25831,N_24359,N_22679);
xnor U25832 (N_25832,N_20820,N_22264);
nand U25833 (N_25833,N_22182,N_21901);
or U25834 (N_25834,N_21351,N_22987);
xor U25835 (N_25835,N_22363,N_23630);
or U25836 (N_25836,N_22581,N_24972);
xnor U25837 (N_25837,N_21577,N_20947);
or U25838 (N_25838,N_22081,N_20858);
or U25839 (N_25839,N_21302,N_23783);
and U25840 (N_25840,N_21190,N_24482);
or U25841 (N_25841,N_22905,N_24065);
xnor U25842 (N_25842,N_21902,N_23326);
nor U25843 (N_25843,N_22072,N_20256);
and U25844 (N_25844,N_20424,N_24670);
nand U25845 (N_25845,N_22157,N_20903);
and U25846 (N_25846,N_20051,N_23252);
nor U25847 (N_25847,N_23662,N_22580);
and U25848 (N_25848,N_22423,N_21525);
or U25849 (N_25849,N_24049,N_24358);
or U25850 (N_25850,N_22040,N_22425);
nand U25851 (N_25851,N_24190,N_23272);
or U25852 (N_25852,N_22518,N_21771);
nor U25853 (N_25853,N_20306,N_23867);
xnor U25854 (N_25854,N_23026,N_22303);
or U25855 (N_25855,N_20757,N_22884);
or U25856 (N_25856,N_23388,N_23924);
nand U25857 (N_25857,N_24831,N_24658);
xor U25858 (N_25858,N_20023,N_23963);
or U25859 (N_25859,N_24236,N_24217);
xor U25860 (N_25860,N_23433,N_21386);
xor U25861 (N_25861,N_20592,N_22588);
nor U25862 (N_25862,N_22455,N_21500);
nand U25863 (N_25863,N_21370,N_24540);
xnor U25864 (N_25864,N_22470,N_21651);
or U25865 (N_25865,N_24839,N_20137);
nor U25866 (N_25866,N_22329,N_22151);
or U25867 (N_25867,N_22940,N_23816);
xor U25868 (N_25868,N_22675,N_20657);
and U25869 (N_25869,N_20232,N_21254);
and U25870 (N_25870,N_22921,N_23962);
or U25871 (N_25871,N_23434,N_22727);
or U25872 (N_25872,N_22538,N_23427);
and U25873 (N_25873,N_22557,N_24930);
xnor U25874 (N_25874,N_23604,N_22257);
and U25875 (N_25875,N_22023,N_24247);
and U25876 (N_25876,N_22219,N_23920);
and U25877 (N_25877,N_20767,N_21285);
nor U25878 (N_25878,N_22281,N_24333);
nor U25879 (N_25879,N_24122,N_23555);
nor U25880 (N_25880,N_23915,N_20289);
and U25881 (N_25881,N_21249,N_23270);
and U25882 (N_25882,N_22897,N_21453);
nand U25883 (N_25883,N_21656,N_20590);
and U25884 (N_25884,N_23778,N_23545);
and U25885 (N_25885,N_22926,N_23167);
xnor U25886 (N_25886,N_22981,N_23093);
nor U25887 (N_25887,N_24518,N_23367);
nand U25888 (N_25888,N_21861,N_21497);
nand U25889 (N_25889,N_21215,N_22221);
or U25890 (N_25890,N_20401,N_21835);
xor U25891 (N_25891,N_20809,N_22064);
nor U25892 (N_25892,N_23303,N_24305);
or U25893 (N_25893,N_22269,N_21733);
nand U25894 (N_25894,N_20000,N_23851);
or U25895 (N_25895,N_21157,N_20017);
and U25896 (N_25896,N_23101,N_24579);
xnor U25897 (N_25897,N_20969,N_21874);
nor U25898 (N_25898,N_23500,N_24873);
and U25899 (N_25899,N_21283,N_24220);
nand U25900 (N_25900,N_23780,N_21374);
and U25901 (N_25901,N_22349,N_24089);
and U25902 (N_25902,N_21698,N_20806);
and U25903 (N_25903,N_22547,N_20916);
and U25904 (N_25904,N_20117,N_20031);
or U25905 (N_25905,N_21427,N_20804);
and U25906 (N_25906,N_20830,N_21985);
or U25907 (N_25907,N_23835,N_21886);
xnor U25908 (N_25908,N_22592,N_24422);
and U25909 (N_25909,N_22346,N_21530);
nor U25910 (N_25910,N_20668,N_21125);
or U25911 (N_25911,N_22994,N_24430);
nor U25912 (N_25912,N_22240,N_23463);
xor U25913 (N_25913,N_22486,N_24773);
xor U25914 (N_25914,N_22361,N_24878);
or U25915 (N_25915,N_22708,N_24901);
nand U25916 (N_25916,N_21196,N_23644);
or U25917 (N_25917,N_22521,N_21629);
or U25918 (N_25918,N_20769,N_20420);
xnor U25919 (N_25919,N_21890,N_23686);
nor U25920 (N_25920,N_21013,N_24527);
nand U25921 (N_25921,N_23540,N_22755);
nor U25922 (N_25922,N_24899,N_22801);
or U25923 (N_25923,N_21261,N_23857);
xor U25924 (N_25924,N_20316,N_22786);
nor U25925 (N_25925,N_23845,N_23830);
nor U25926 (N_25926,N_22397,N_23471);
xor U25927 (N_25927,N_21398,N_20591);
and U25928 (N_25928,N_21325,N_22301);
or U25929 (N_25929,N_20834,N_24304);
xor U25930 (N_25930,N_22323,N_23157);
nand U25931 (N_25931,N_23264,N_23629);
and U25932 (N_25932,N_24320,N_23665);
xor U25933 (N_25933,N_23206,N_20869);
or U25934 (N_25934,N_23598,N_21032);
and U25935 (N_25935,N_21143,N_23420);
or U25936 (N_25936,N_20768,N_24473);
nor U25937 (N_25937,N_24634,N_22232);
nor U25938 (N_25938,N_23824,N_20132);
nand U25939 (N_25939,N_20179,N_20296);
or U25940 (N_25940,N_22106,N_24647);
xnor U25941 (N_25941,N_24409,N_22945);
xnor U25942 (N_25942,N_24826,N_21758);
xnor U25943 (N_25943,N_23607,N_24940);
nand U25944 (N_25944,N_22780,N_24627);
and U25945 (N_25945,N_21555,N_20127);
and U25946 (N_25946,N_21152,N_20743);
xnor U25947 (N_25947,N_22659,N_23219);
xnor U25948 (N_25948,N_22599,N_24408);
nor U25949 (N_25949,N_21423,N_21247);
xnor U25950 (N_25950,N_21192,N_22113);
xnor U25951 (N_25951,N_24897,N_21268);
and U25952 (N_25952,N_20019,N_22177);
and U25953 (N_25953,N_23891,N_24094);
xnor U25954 (N_25954,N_20612,N_22787);
and U25955 (N_25955,N_21760,N_21188);
nor U25956 (N_25956,N_20687,N_20136);
and U25957 (N_25957,N_20459,N_24371);
and U25958 (N_25958,N_22632,N_24147);
or U25959 (N_25959,N_21851,N_22584);
xor U25960 (N_25960,N_23895,N_24045);
xor U25961 (N_25961,N_21907,N_23533);
nand U25962 (N_25962,N_20581,N_24008);
or U25963 (N_25963,N_24888,N_20029);
xor U25964 (N_25964,N_20168,N_22487);
or U25965 (N_25965,N_24301,N_24565);
or U25966 (N_25966,N_21354,N_24959);
xnor U25967 (N_25967,N_24413,N_24267);
nand U25968 (N_25968,N_23197,N_24623);
xor U25969 (N_25969,N_21069,N_24525);
nand U25970 (N_25970,N_22387,N_22353);
nand U25971 (N_25971,N_21145,N_23436);
xnor U25972 (N_25972,N_20222,N_20253);
or U25973 (N_25973,N_22816,N_22955);
nor U25974 (N_25974,N_21710,N_21085);
nand U25975 (N_25975,N_23041,N_21811);
xnor U25976 (N_25976,N_23751,N_21089);
or U25977 (N_25977,N_20888,N_24029);
or U25978 (N_25978,N_24039,N_24078);
nor U25979 (N_25979,N_24956,N_22779);
and U25980 (N_25980,N_23449,N_20044);
or U25981 (N_25981,N_23798,N_20739);
xnor U25982 (N_25982,N_24450,N_22441);
or U25983 (N_25983,N_23425,N_22071);
nand U25984 (N_25984,N_22218,N_23117);
nor U25985 (N_25985,N_23507,N_22843);
xnor U25986 (N_25986,N_21327,N_22740);
nor U25987 (N_25987,N_24052,N_22262);
nand U25988 (N_25988,N_20255,N_24543);
or U25989 (N_25989,N_21753,N_23885);
nand U25990 (N_25990,N_21332,N_20512);
and U25991 (N_25991,N_23274,N_21823);
nand U25992 (N_25992,N_23263,N_21562);
nor U25993 (N_25993,N_20346,N_21983);
nand U25994 (N_25994,N_22320,N_21791);
and U25995 (N_25995,N_24844,N_20337);
xnor U25996 (N_25996,N_21158,N_20074);
and U25997 (N_25997,N_22867,N_24505);
nand U25998 (N_25998,N_22360,N_21987);
and U25999 (N_25999,N_21722,N_23091);
xnor U26000 (N_26000,N_22308,N_21450);
and U26001 (N_26001,N_21277,N_23909);
or U26002 (N_26002,N_21737,N_21419);
nor U26003 (N_26003,N_23937,N_21061);
nor U26004 (N_26004,N_20537,N_24838);
or U26005 (N_26005,N_22681,N_21821);
nand U26006 (N_26006,N_21735,N_24493);
nor U26007 (N_26007,N_20746,N_23455);
nor U26008 (N_26008,N_21564,N_20377);
nand U26009 (N_26009,N_20054,N_23123);
nor U26010 (N_26010,N_21334,N_24096);
nand U26011 (N_26011,N_20282,N_21672);
xnor U26012 (N_26012,N_23390,N_21170);
xnor U26013 (N_26013,N_23772,N_22176);
xnor U26014 (N_26014,N_20643,N_20513);
or U26015 (N_26015,N_23508,N_20212);
xor U26016 (N_26016,N_20250,N_20402);
and U26017 (N_26017,N_21624,N_20950);
and U26018 (N_26018,N_21641,N_22052);
nor U26019 (N_26019,N_23981,N_21164);
nand U26020 (N_26020,N_24199,N_20883);
or U26021 (N_26021,N_20957,N_20862);
xor U26022 (N_26022,N_23153,N_22299);
nor U26023 (N_26023,N_20344,N_21743);
or U26024 (N_26024,N_20172,N_24060);
nand U26025 (N_26025,N_24545,N_22836);
and U26026 (N_26026,N_24997,N_20055);
and U26027 (N_26027,N_21272,N_22600);
or U26028 (N_26028,N_20123,N_21703);
or U26029 (N_26029,N_21369,N_22725);
xnor U26030 (N_26030,N_20001,N_23593);
xor U26031 (N_26031,N_20973,N_20829);
or U26032 (N_26032,N_22579,N_23755);
xor U26033 (N_26033,N_21566,N_24601);
and U26034 (N_26034,N_20182,N_20726);
xnor U26035 (N_26035,N_23625,N_24872);
nor U26036 (N_26036,N_22515,N_24723);
and U26037 (N_26037,N_20647,N_23503);
or U26038 (N_26038,N_22431,N_23846);
and U26039 (N_26039,N_23805,N_22312);
nor U26040 (N_26040,N_21240,N_24598);
nor U26041 (N_26041,N_20376,N_23645);
and U26042 (N_26042,N_24858,N_23568);
xor U26043 (N_26043,N_24275,N_21809);
nor U26044 (N_26044,N_21716,N_23339);
nor U26045 (N_26045,N_23185,N_23066);
nand U26046 (N_26046,N_21912,N_20080);
or U26047 (N_26047,N_21695,N_22759);
nand U26048 (N_26048,N_21581,N_20240);
and U26049 (N_26049,N_22259,N_24566);
nand U26050 (N_26050,N_23639,N_21649);
nand U26051 (N_26051,N_22999,N_23191);
nor U26052 (N_26052,N_22497,N_20898);
nor U26053 (N_26053,N_23529,N_22067);
nand U26054 (N_26054,N_20161,N_20720);
nor U26055 (N_26055,N_24036,N_22782);
nand U26056 (N_26056,N_23615,N_20220);
nand U26057 (N_26057,N_24151,N_20801);
xnor U26058 (N_26058,N_23802,N_23251);
and U26059 (N_26059,N_24180,N_20293);
and U26060 (N_26060,N_22967,N_22288);
and U26061 (N_26061,N_21797,N_24150);
xnor U26062 (N_26062,N_23346,N_24381);
nand U26063 (N_26063,N_24003,N_23140);
xor U26064 (N_26064,N_20645,N_20707);
or U26065 (N_26065,N_23678,N_21098);
nand U26066 (N_26066,N_20041,N_24671);
nor U26067 (N_26067,N_23774,N_21928);
nor U26068 (N_26068,N_21399,N_24797);
nand U26069 (N_26069,N_24814,N_23812);
xnor U26070 (N_26070,N_21220,N_23999);
and U26071 (N_26071,N_24396,N_22418);
nor U26072 (N_26072,N_23382,N_20860);
or U26073 (N_26073,N_22545,N_22442);
xor U26074 (N_26074,N_20776,N_21435);
or U26075 (N_26075,N_24818,N_20611);
nor U26076 (N_26076,N_21717,N_21479);
or U26077 (N_26077,N_21625,N_22757);
nor U26078 (N_26078,N_24014,N_23651);
nand U26079 (N_26079,N_20855,N_23328);
nor U26080 (N_26080,N_23993,N_24988);
nand U26081 (N_26081,N_24233,N_21647);
or U26082 (N_26082,N_23350,N_21583);
nand U26083 (N_26083,N_24520,N_23043);
nor U26084 (N_26084,N_24018,N_20478);
nor U26085 (N_26085,N_24581,N_24015);
nand U26086 (N_26086,N_22677,N_20439);
xor U26087 (N_26087,N_20666,N_20221);
nor U26088 (N_26088,N_23932,N_20615);
nor U26089 (N_26089,N_24144,N_20951);
nor U26090 (N_26090,N_20134,N_22010);
nor U26091 (N_26091,N_24374,N_20007);
xor U26092 (N_26092,N_24443,N_24246);
xor U26093 (N_26093,N_24214,N_24401);
or U26094 (N_26094,N_23217,N_21557);
nor U26095 (N_26095,N_24741,N_21154);
nor U26096 (N_26096,N_23832,N_24801);
nand U26097 (N_26097,N_20610,N_21110);
or U26098 (N_26098,N_24479,N_21258);
xor U26099 (N_26099,N_22336,N_22380);
or U26100 (N_26100,N_23323,N_24277);
and U26101 (N_26101,N_21690,N_20387);
and U26102 (N_26102,N_23679,N_23534);
xnor U26103 (N_26103,N_20335,N_24822);
xnor U26104 (N_26104,N_22840,N_20882);
xor U26105 (N_26105,N_20158,N_21606);
nor U26106 (N_26106,N_23113,N_21598);
or U26107 (N_26107,N_21214,N_21008);
xnor U26108 (N_26108,N_24495,N_23890);
xor U26109 (N_26109,N_21348,N_22827);
nand U26110 (N_26110,N_23648,N_22305);
xnor U26111 (N_26111,N_22674,N_20578);
nor U26112 (N_26112,N_22460,N_22469);
and U26113 (N_26113,N_20133,N_20481);
or U26114 (N_26114,N_24763,N_24903);
and U26115 (N_26115,N_23459,N_23051);
nand U26116 (N_26116,N_21989,N_24481);
xnor U26117 (N_26117,N_22965,N_20929);
nor U26118 (N_26118,N_21838,N_23868);
nor U26119 (N_26119,N_21953,N_24852);
nand U26120 (N_26120,N_24310,N_24895);
and U26121 (N_26121,N_23480,N_23118);
nand U26122 (N_26122,N_24300,N_24128);
nand U26123 (N_26123,N_22087,N_20283);
nand U26124 (N_26124,N_22863,N_23719);
xnor U26125 (N_26125,N_21704,N_22483);
nor U26126 (N_26126,N_24884,N_24120);
nor U26127 (N_26127,N_20589,N_24109);
xnor U26128 (N_26128,N_20983,N_24816);
and U26129 (N_26129,N_21491,N_22957);
and U26130 (N_26130,N_21335,N_22946);
or U26131 (N_26131,N_23488,N_24040);
or U26132 (N_26132,N_24243,N_23986);
xnor U26133 (N_26133,N_24234,N_21056);
nand U26134 (N_26134,N_21670,N_24477);
xnor U26135 (N_26135,N_21077,N_21848);
and U26136 (N_26136,N_23840,N_24428);
nor U26137 (N_26137,N_23246,N_21346);
nor U26138 (N_26138,N_23004,N_22542);
or U26139 (N_26139,N_21235,N_22293);
or U26140 (N_26140,N_21648,N_22815);
xor U26141 (N_26141,N_23380,N_20865);
nor U26142 (N_26142,N_20398,N_24662);
nor U26143 (N_26143,N_23240,N_22821);
nor U26144 (N_26144,N_20712,N_20515);
nand U26145 (N_26145,N_21982,N_21217);
or U26146 (N_26146,N_23494,N_23984);
nor U26147 (N_26147,N_20300,N_24465);
nand U26148 (N_26148,N_24276,N_20880);
nand U26149 (N_26149,N_22662,N_23575);
or U26150 (N_26150,N_22776,N_21891);
or U26151 (N_26151,N_20932,N_23111);
nor U26152 (N_26152,N_20920,N_20162);
and U26153 (N_26153,N_24584,N_21893);
nor U26154 (N_26154,N_20294,N_24725);
nor U26155 (N_26155,N_22657,N_20735);
nor U26156 (N_26156,N_21344,N_22754);
nor U26157 (N_26157,N_24244,N_24774);
nor U26158 (N_26158,N_24414,N_23077);
nor U26159 (N_26159,N_24461,N_21151);
nand U26160 (N_26160,N_20444,N_22215);
and U26161 (N_26161,N_21198,N_21796);
and U26162 (N_26162,N_20012,N_20309);
nor U26163 (N_26163,N_24502,N_24490);
nand U26164 (N_26164,N_23841,N_22191);
or U26165 (N_26165,N_23107,N_21896);
nand U26166 (N_26166,N_20303,N_21940);
and U26167 (N_26167,N_21900,N_22417);
xor U26168 (N_26168,N_22749,N_21339);
or U26169 (N_26169,N_24240,N_20959);
or U26170 (N_26170,N_24097,N_23888);
nand U26171 (N_26171,N_24133,N_24892);
or U26172 (N_26172,N_22936,N_20167);
nand U26173 (N_26173,N_21970,N_24517);
nand U26174 (N_26174,N_23786,N_23611);
or U26175 (N_26175,N_22144,N_21709);
nand U26176 (N_26176,N_20562,N_23520);
or U26177 (N_26177,N_20209,N_21601);
xor U26178 (N_26178,N_20714,N_24436);
nand U26179 (N_26179,N_23325,N_23801);
and U26180 (N_26180,N_22802,N_20503);
nand U26181 (N_26181,N_24692,N_22437);
xnor U26182 (N_26182,N_22577,N_20715);
xnor U26183 (N_26183,N_20828,N_23048);
xor U26184 (N_26184,N_20485,N_23036);
xor U26185 (N_26185,N_22204,N_23821);
xor U26186 (N_26186,N_21452,N_20458);
xor U26187 (N_26187,N_21741,N_20818);
xor U26188 (N_26188,N_23767,N_21650);
nor U26189 (N_26189,N_22273,N_20607);
nor U26190 (N_26190,N_22482,N_23203);
and U26191 (N_26191,N_22413,N_22212);
and U26192 (N_26192,N_24448,N_20195);
and U26193 (N_26193,N_23955,N_24893);
nor U26194 (N_26194,N_21666,N_21613);
nor U26195 (N_26195,N_24789,N_23033);
and U26196 (N_26196,N_22767,N_23447);
or U26197 (N_26197,N_22707,N_23537);
and U26198 (N_26198,N_24910,N_22523);
nor U26199 (N_26199,N_21556,N_21565);
or U26200 (N_26200,N_23315,N_22386);
and U26201 (N_26201,N_22192,N_22506);
nor U26202 (N_26202,N_24553,N_22571);
and U26203 (N_26203,N_21371,N_22544);
nand U26204 (N_26204,N_24037,N_24508);
xor U26205 (N_26205,N_20857,N_23861);
and U26206 (N_26206,N_21445,N_24033);
nor U26207 (N_26207,N_21820,N_20486);
nor U26208 (N_26208,N_24790,N_23154);
xor U26209 (N_26209,N_22742,N_21959);
xor U26210 (N_26210,N_21529,N_23292);
or U26211 (N_26211,N_20644,N_24373);
nand U26212 (N_26212,N_22261,N_22568);
nor U26213 (N_26213,N_24947,N_21880);
nor U26214 (N_26214,N_24585,N_22698);
nor U26215 (N_26215,N_20341,N_24848);
nand U26216 (N_26216,N_20200,N_23609);
nand U26217 (N_26217,N_23147,N_23715);
and U26218 (N_26218,N_20363,N_21662);
xor U26219 (N_26219,N_24061,N_20674);
and U26220 (N_26220,N_20066,N_20238);
xor U26221 (N_26221,N_24863,N_22697);
nand U26222 (N_26222,N_21905,N_20273);
and U26223 (N_26223,N_21233,N_20070);
nor U26224 (N_26224,N_21776,N_20151);
and U26225 (N_26225,N_24238,N_23799);
xor U26226 (N_26226,N_21532,N_22184);
xnor U26227 (N_26227,N_23269,N_24378);
and U26228 (N_26228,N_21879,N_20106);
or U26229 (N_26229,N_20689,N_24192);
or U26230 (N_26230,N_21115,N_24742);
and U26231 (N_26231,N_21962,N_20463);
and U26232 (N_26232,N_22882,N_21014);
nand U26233 (N_26233,N_23672,N_23620);
or U26234 (N_26234,N_20482,N_22083);
xor U26235 (N_26235,N_23095,N_24938);
nand U26236 (N_26236,N_21389,N_20406);
xor U26237 (N_26237,N_24941,N_22734);
xnor U26238 (N_26238,N_23818,N_24572);
xnor U26239 (N_26239,N_20391,N_20817);
and U26240 (N_26240,N_24303,N_20844);
and U26241 (N_26241,N_23016,N_21041);
xnor U26242 (N_26242,N_22463,N_22533);
nand U26243 (N_26243,N_24156,N_21229);
and U26244 (N_26244,N_21512,N_22381);
and U26245 (N_26245,N_21345,N_20086);
or U26246 (N_26246,N_22488,N_21205);
or U26247 (N_26247,N_21030,N_20091);
nor U26248 (N_26248,N_22552,N_21183);
and U26249 (N_26249,N_20169,N_21091);
nand U26250 (N_26250,N_20572,N_21467);
nor U26251 (N_26251,N_23330,N_23190);
nand U26252 (N_26252,N_24411,N_21920);
xnor U26253 (N_26253,N_24331,N_24339);
and U26254 (N_26254,N_21036,N_22224);
xor U26255 (N_26255,N_24506,N_24126);
nor U26256 (N_26256,N_21862,N_24775);
xnor U26257 (N_26257,N_20583,N_20601);
or U26258 (N_26258,N_21052,N_23912);
nand U26259 (N_26259,N_21244,N_20876);
nor U26260 (N_26260,N_21685,N_21040);
or U26261 (N_26261,N_24343,N_22638);
xnor U26262 (N_26262,N_21927,N_23377);
xor U26263 (N_26263,N_23230,N_22135);
or U26264 (N_26264,N_22942,N_24678);
and U26265 (N_26265,N_23184,N_22001);
nor U26266 (N_26266,N_23424,N_24859);
nand U26267 (N_26267,N_21972,N_21948);
or U26268 (N_26268,N_24603,N_22554);
or U26269 (N_26269,N_24827,N_22774);
nand U26270 (N_26270,N_20624,N_24739);
nand U26271 (N_26271,N_22166,N_24574);
xnor U26272 (N_26272,N_24368,N_20089);
nand U26273 (N_26273,N_23950,N_24046);
nor U26274 (N_26274,N_20805,N_20385);
and U26275 (N_26275,N_23636,N_22666);
xor U26276 (N_26276,N_24541,N_21552);
and U26277 (N_26277,N_24885,N_21787);
and U26278 (N_26278,N_21010,N_20595);
nor U26279 (N_26279,N_20190,N_23220);
and U26280 (N_26280,N_24325,N_23882);
nand U26281 (N_26281,N_21679,N_20514);
xnor U26282 (N_26282,N_23633,N_24379);
nand U26283 (N_26283,N_20246,N_22136);
and U26284 (N_26284,N_23640,N_24453);
nor U26285 (N_26285,N_21384,N_24622);
nor U26286 (N_26286,N_22280,N_23982);
or U26287 (N_26287,N_20627,N_20171);
xnor U26288 (N_26288,N_24335,N_20659);
xor U26289 (N_26289,N_24597,N_20483);
nand U26290 (N_26290,N_20352,N_23058);
nand U26291 (N_26291,N_20887,N_20594);
nor U26292 (N_26292,N_22881,N_21136);
nand U26293 (N_26293,N_23820,N_24621);
nor U26294 (N_26294,N_20693,N_24726);
xnor U26295 (N_26295,N_23960,N_20404);
nand U26296 (N_26296,N_20103,N_22284);
and U26297 (N_26297,N_24669,N_24372);
xor U26298 (N_26298,N_20129,N_21608);
nand U26299 (N_26299,N_22325,N_20237);
or U26300 (N_26300,N_21161,N_22041);
or U26301 (N_26301,N_20524,N_22672);
and U26302 (N_26302,N_24361,N_20295);
nor U26303 (N_26303,N_22333,N_22054);
nor U26304 (N_26304,N_23522,N_24616);
or U26305 (N_26305,N_22658,N_20276);
or U26306 (N_26306,N_24600,N_21187);
or U26307 (N_26307,N_24352,N_23499);
and U26308 (N_26308,N_23581,N_24833);
nand U26309 (N_26309,N_22953,N_22383);
xnor U26310 (N_26310,N_20704,N_23682);
nor U26311 (N_26311,N_22818,N_20692);
xnor U26312 (N_26312,N_21731,N_21129);
nor U26313 (N_26313,N_21858,N_22421);
xor U26314 (N_26314,N_24953,N_24225);
nor U26315 (N_26315,N_23965,N_20105);
nor U26316 (N_26316,N_21730,N_22875);
nand U26317 (N_26317,N_20878,N_24142);
nand U26318 (N_26318,N_24207,N_22448);
nand U26319 (N_26319,N_20407,N_21333);
xnor U26320 (N_26320,N_20193,N_23994);
nor U26321 (N_26321,N_23526,N_20533);
nor U26322 (N_26322,N_23031,N_23037);
or U26323 (N_26323,N_21498,N_23360);
xnor U26324 (N_26324,N_20082,N_22849);
and U26325 (N_26325,N_22685,N_22246);
xnor U26326 (N_26326,N_23250,N_20856);
and U26327 (N_26327,N_20332,N_20939);
and U26328 (N_26328,N_21065,N_21326);
xor U26329 (N_26329,N_24968,N_24778);
xnor U26330 (N_26330,N_24665,N_21786);
nand U26331 (N_26331,N_22237,N_20825);
nand U26332 (N_26332,N_20972,N_22376);
nand U26333 (N_26333,N_24270,N_22640);
nor U26334 (N_26334,N_20360,N_22109);
nor U26335 (N_26335,N_22302,N_22100);
nor U26336 (N_26336,N_24537,N_20602);
or U26337 (N_26337,N_24676,N_21819);
and U26338 (N_26338,N_23959,N_24024);
xor U26339 (N_26339,N_22276,N_21708);
or U26340 (N_26340,N_24973,N_20314);
or U26341 (N_26341,N_21978,N_21843);
or U26342 (N_26342,N_21262,N_24127);
and U26343 (N_26343,N_23301,N_22906);
nor U26344 (N_26344,N_20374,N_21997);
nand U26345 (N_26345,N_21923,N_23416);
nor U26346 (N_26346,N_20962,N_23032);
and U26347 (N_26347,N_24925,N_22692);
nand U26348 (N_26348,N_24754,N_20541);
nand U26349 (N_26349,N_23899,N_21274);
nor U26350 (N_26350,N_21084,N_23822);
nor U26351 (N_26351,N_23284,N_20053);
and U26352 (N_26352,N_22817,N_23015);
or U26353 (N_26353,N_22036,N_22451);
nor U26354 (N_26354,N_21857,N_23788);
and U26355 (N_26355,N_20353,N_24531);
or U26356 (N_26356,N_24316,N_21906);
nor U26357 (N_26357,N_23953,N_20546);
nor U26358 (N_26358,N_21312,N_24939);
nand U26359 (N_26359,N_20251,N_22296);
and U26360 (N_26360,N_21916,N_21366);
xnor U26361 (N_26361,N_23321,N_23460);
and U26362 (N_26362,N_23729,N_24989);
nand U26363 (N_26363,N_20415,N_20489);
and U26364 (N_26364,N_23068,N_21996);
nor U26365 (N_26365,N_23288,N_21173);
and U26366 (N_26366,N_20073,N_24811);
nor U26367 (N_26367,N_22596,N_20902);
nand U26368 (N_26368,N_21286,N_23442);
or U26369 (N_26369,N_23408,N_21792);
nor U26370 (N_26370,N_22148,N_23902);
or U26371 (N_26371,N_23771,N_22179);
or U26372 (N_26372,N_22800,N_20575);
and U26373 (N_26373,N_20016,N_21360);
or U26374 (N_26374,N_24245,N_24116);
or U26375 (N_26375,N_22377,N_24051);
xnor U26376 (N_26376,N_22484,N_22095);
xor U26377 (N_26377,N_20442,N_23856);
or U26378 (N_26378,N_22084,N_22267);
nor U26379 (N_26379,N_24499,N_24221);
xor U26380 (N_26380,N_22914,N_20223);
nand U26381 (N_26381,N_21510,N_24042);
and U26382 (N_26382,N_24758,N_23072);
xor U26383 (N_26383,N_20733,N_21024);
nand U26384 (N_26384,N_21238,N_24478);
or U26385 (N_26385,N_23156,N_21373);
and U26386 (N_26386,N_23933,N_24696);
nand U26387 (N_26387,N_24886,N_22864);
or U26388 (N_26388,N_24681,N_22718);
or U26389 (N_26389,N_20731,N_20272);
nand U26390 (N_26390,N_23510,N_22935);
nand U26391 (N_26391,N_24614,N_20056);
and U26392 (N_26392,N_20499,N_22338);
or U26393 (N_26393,N_23573,N_21156);
or U26394 (N_26394,N_21739,N_23539);
or U26395 (N_26395,N_21035,N_21549);
nor U26396 (N_26396,N_21538,N_23126);
nor U26397 (N_26397,N_21169,N_22415);
xnor U26398 (N_26398,N_22347,N_22142);
nor U26399 (N_26399,N_23143,N_23423);
nor U26400 (N_26400,N_21181,N_22871);
and U26401 (N_26401,N_24626,N_23509);
nand U26402 (N_26402,N_21058,N_21977);
or U26403 (N_26403,N_24208,N_20616);
nand U26404 (N_26404,N_23869,N_23092);
and U26405 (N_26405,N_20530,N_21909);
or U26406 (N_26406,N_22070,N_23528);
nand U26407 (N_26407,N_24237,N_21471);
xnor U26408 (N_26408,N_21116,N_23657);
or U26409 (N_26409,N_22744,N_24998);
or U26410 (N_26410,N_21340,N_24159);
and U26411 (N_26411,N_20214,N_21957);
nand U26412 (N_26412,N_21403,N_22992);
or U26413 (N_26413,N_22410,N_24249);
or U26414 (N_26414,N_20952,N_23541);
nand U26415 (N_26415,N_20477,N_24643);
and U26416 (N_26416,N_24385,N_21942);
nor U26417 (N_26417,N_23124,N_23989);
nor U26418 (N_26418,N_23432,N_24509);
xnor U26419 (N_26419,N_23797,N_20497);
or U26420 (N_26420,N_23152,N_22820);
nand U26421 (N_26421,N_22593,N_20113);
nand U26422 (N_26422,N_22995,N_21245);
nor U26423 (N_26423,N_20626,N_23971);
nor U26424 (N_26424,N_20756,N_21034);
or U26425 (N_26425,N_21044,N_23216);
xnor U26426 (N_26426,N_24874,N_22883);
xnor U26427 (N_26427,N_21623,N_20130);
and U26428 (N_26428,N_22798,N_22183);
nor U26429 (N_26429,N_24865,N_20342);
xor U26430 (N_26430,N_24633,N_22924);
nand U26431 (N_26431,N_20313,N_22830);
or U26432 (N_26432,N_22889,N_23530);
xor U26433 (N_26433,N_21160,N_23542);
xnor U26434 (N_26434,N_23002,N_20006);
xnor U26435 (N_26435,N_21379,N_24269);
and U26436 (N_26436,N_20248,N_22743);
and U26437 (N_26437,N_20434,N_21619);
and U26438 (N_26438,N_22013,N_20120);
or U26439 (N_26439,N_21888,N_21802);
or U26440 (N_26440,N_21426,N_20690);
and U26441 (N_26441,N_23038,N_24637);
xor U26442 (N_26442,N_22833,N_20043);
nor U26443 (N_26443,N_23926,N_21028);
or U26444 (N_26444,N_22364,N_22068);
and U26445 (N_26445,N_20373,N_23162);
nor U26446 (N_26446,N_22168,N_24673);
or U26447 (N_26447,N_23229,N_24686);
nand U26448 (N_26448,N_22954,N_22714);
nand U26449 (N_26449,N_23592,N_20535);
nor U26450 (N_26450,N_22474,N_22771);
or U26451 (N_26451,N_20655,N_22165);
and U26452 (N_26452,N_24766,N_22458);
or U26453 (N_26453,N_24690,N_20139);
or U26454 (N_26454,N_24059,N_23907);
or U26455 (N_26455,N_22961,N_23758);
xnor U26456 (N_26456,N_23516,N_23634);
and U26457 (N_26457,N_22762,N_21772);
nor U26458 (N_26458,N_22494,N_23839);
nand U26459 (N_26459,N_22989,N_22222);
nand U26460 (N_26460,N_21243,N_22513);
nand U26461 (N_26461,N_24253,N_24183);
nand U26462 (N_26462,N_21794,N_23084);
nand U26463 (N_26463,N_21969,N_21414);
and U26464 (N_26464,N_23760,N_22939);
or U26465 (N_26465,N_20791,N_24324);
nand U26466 (N_26466,N_20835,N_21660);
xor U26467 (N_26467,N_22459,N_24993);
or U26468 (N_26468,N_22908,N_22850);
xor U26469 (N_26469,N_20827,N_21159);
or U26470 (N_26470,N_20320,N_23052);
or U26471 (N_26471,N_23949,N_20087);
or U26472 (N_26472,N_20730,N_22498);
and U26473 (N_26473,N_23376,N_20914);
or U26474 (N_26474,N_24752,N_24882);
xor U26475 (N_26475,N_21729,N_21738);
xor U26476 (N_26476,N_23775,N_20808);
nand U26477 (N_26477,N_24794,N_21633);
xnor U26478 (N_26478,N_22797,N_24319);
nor U26479 (N_26479,N_22604,N_24751);
and U26480 (N_26480,N_22153,N_22201);
or U26481 (N_26481,N_21031,N_23452);
nor U26482 (N_26482,N_22230,N_22665);
nand U26483 (N_26483,N_24659,N_23927);
and U26484 (N_26484,N_22703,N_22869);
and U26485 (N_26485,N_23044,N_23312);
and U26486 (N_26486,N_21388,N_20703);
or U26487 (N_26487,N_22996,N_22551);
xnor U26488 (N_26488,N_21103,N_21620);
nand U26489 (N_26489,N_24390,N_22335);
and U26490 (N_26490,N_23000,N_20265);
nor U26491 (N_26491,N_22602,N_21266);
or U26492 (N_26492,N_24835,N_23776);
or U26493 (N_26493,N_23602,N_24259);
xor U26494 (N_26494,N_22062,N_24441);
or U26495 (N_26495,N_24651,N_24564);
xor U26496 (N_26496,N_23759,N_21067);
and U26497 (N_26497,N_23340,N_20945);
nor U26498 (N_26498,N_21429,N_24255);
nor U26499 (N_26499,N_20763,N_22304);
xor U26500 (N_26500,N_20890,N_24781);
nor U26501 (N_26501,N_21341,N_22020);
and U26502 (N_26502,N_20010,N_21362);
nor U26503 (N_26503,N_24524,N_23009);
xor U26504 (N_26504,N_21411,N_20955);
nor U26505 (N_26505,N_21431,N_24420);
xnor U26506 (N_26506,N_22348,N_24514);
or U26507 (N_26507,N_24340,N_23394);
nand U26508 (N_26508,N_20819,N_24552);
or U26509 (N_26509,N_21933,N_23557);
nor U26510 (N_26510,N_23337,N_20879);
nor U26511 (N_26511,N_22624,N_21520);
nor U26512 (N_26512,N_22171,N_21757);
or U26513 (N_26513,N_21550,N_23466);
and U26514 (N_26514,N_20394,N_22570);
or U26515 (N_26515,N_20779,N_22429);
nand U26516 (N_26516,N_22450,N_24418);
xnor U26517 (N_26517,N_20729,N_23967);
and U26518 (N_26518,N_22409,N_23304);
nand U26519 (N_26519,N_22065,N_21359);
nand U26520 (N_26520,N_24286,N_21250);
xor U26521 (N_26521,N_23236,N_23286);
xor U26522 (N_26522,N_24779,N_21815);
nor U26523 (N_26523,N_20180,N_22339);
xnor U26524 (N_26524,N_24615,N_22159);
nor U26525 (N_26525,N_22678,N_23285);
and U26526 (N_26526,N_22673,N_21615);
or U26527 (N_26527,N_20138,N_21747);
nor U26528 (N_26528,N_21134,N_23019);
nor U26529 (N_26529,N_20131,N_21021);
xnor U26530 (N_26530,N_23901,N_21019);
nor U26531 (N_26531,N_20395,N_20196);
nand U26532 (N_26532,N_22598,N_23838);
xor U26533 (N_26533,N_22695,N_23362);
or U26534 (N_26534,N_20577,N_21456);
nor U26535 (N_26535,N_24722,N_22250);
or U26536 (N_26536,N_24575,N_20034);
or U26537 (N_26537,N_20837,N_20417);
nor U26538 (N_26538,N_24047,N_23518);
and U26539 (N_26539,N_23792,N_23456);
and U26540 (N_26540,N_21563,N_23245);
xor U26541 (N_26541,N_24295,N_24652);
nor U26542 (N_26542,N_20115,N_22783);
nand U26543 (N_26543,N_24016,N_22248);
or U26544 (N_26544,N_24701,N_23407);
nand U26545 (N_26545,N_23055,N_23808);
nand U26546 (N_26546,N_20991,N_20124);
xnor U26547 (N_26547,N_23998,N_23570);
xor U26548 (N_26548,N_24922,N_24412);
or U26549 (N_26549,N_23566,N_21495);
or U26550 (N_26550,N_22558,N_22407);
nand U26551 (N_26551,N_20257,N_22635);
nand U26552 (N_26552,N_20826,N_23387);
nor U26553 (N_26553,N_20843,N_20526);
nor U26554 (N_26554,N_20281,N_20919);
nand U26555 (N_26555,N_22788,N_23331);
or U26556 (N_26556,N_24904,N_22887);
xor U26557 (N_26557,N_24698,N_23554);
xnor U26558 (N_26558,N_21155,N_23322);
or U26559 (N_26559,N_22769,N_22078);
nand U26560 (N_26560,N_20896,N_24296);
nand U26561 (N_26561,N_21117,N_22952);
and U26562 (N_26562,N_22565,N_20841);
and U26563 (N_26563,N_20906,N_22529);
nand U26564 (N_26564,N_22310,N_22758);
and U26565 (N_26565,N_21895,N_24182);
xor U26566 (N_26566,N_21328,N_23430);
xnor U26567 (N_26567,N_21114,N_23400);
xnor U26568 (N_26568,N_21093,N_24162);
nand U26569 (N_26569,N_23743,N_21246);
xnor U26570 (N_26570,N_21076,N_22630);
nor U26571 (N_26571,N_23472,N_22912);
nand U26572 (N_26572,N_22728,N_24586);
or U26573 (N_26573,N_23001,N_21773);
nand U26574 (N_26574,N_21761,N_24521);
nor U26575 (N_26575,N_20025,N_23789);
or U26576 (N_26576,N_23273,N_20003);
nor U26577 (N_26577,N_24098,N_21674);
nand U26578 (N_26578,N_20498,N_22958);
nand U26579 (N_26579,N_22050,N_24526);
and U26580 (N_26580,N_23121,N_20476);
or U26581 (N_26581,N_23561,N_22396);
nand U26582 (N_26582,N_20384,N_23357);
nor U26583 (N_26583,N_23646,N_22141);
xor U26584 (N_26584,N_23277,N_21127);
nand U26585 (N_26585,N_21361,N_20552);
nand U26586 (N_26586,N_20400,N_20547);
or U26587 (N_26587,N_20842,N_22031);
xnor U26588 (N_26588,N_20128,N_23324);
nor U26589 (N_26589,N_21226,N_22394);
nor U26590 (N_26590,N_23133,N_22804);
and U26591 (N_26591,N_20872,N_20473);
nor U26592 (N_26592,N_23012,N_22366);
and U26593 (N_26593,N_21025,N_24118);
and U26594 (N_26594,N_22982,N_24119);
nand U26595 (N_26595,N_20263,N_21082);
nor U26596 (N_26596,N_21464,N_22845);
xor U26597 (N_26597,N_21892,N_23223);
or U26598 (N_26598,N_20638,N_23674);
nand U26599 (N_26599,N_22079,N_21207);
or U26600 (N_26600,N_24994,N_23074);
nand U26601 (N_26601,N_20885,N_24383);
nand U26602 (N_26602,N_20521,N_23706);
xnor U26603 (N_26603,N_20629,N_21029);
nand U26604 (N_26604,N_20661,N_23307);
nor U26605 (N_26605,N_20651,N_23887);
or U26606 (N_26606,N_23966,N_20096);
nand U26607 (N_26607,N_24927,N_22172);
nand U26608 (N_26608,N_21278,N_20517);
or U26609 (N_26609,N_20679,N_20264);
nand U26610 (N_26610,N_22668,N_21391);
and U26611 (N_26611,N_23676,N_24136);
and U26612 (N_26612,N_23276,N_24975);
nand U26613 (N_26613,N_23265,N_20440);
nand U26614 (N_26614,N_24091,N_24836);
nor U26615 (N_26615,N_20350,N_24729);
nor U26616 (N_26616,N_23439,N_24942);
xnor U26617 (N_26617,N_24929,N_23813);
nor U26618 (N_26618,N_21974,N_22468);
xnor U26619 (N_26619,N_20788,N_20004);
nand U26620 (N_26620,N_20327,N_21146);
nand U26621 (N_26621,N_24738,N_20848);
nor U26622 (N_26622,N_22235,N_20831);
or U26623 (N_26623,N_23757,N_24184);
nor U26624 (N_26624,N_22306,N_21812);
nor U26625 (N_26625,N_22811,N_24936);
or U26626 (N_26626,N_23003,N_22419);
xnor U26627 (N_26627,N_21543,N_21443);
xor U26628 (N_26628,N_21273,N_22197);
nor U26629 (N_26629,N_22045,N_24834);
nor U26630 (N_26630,N_23708,N_22251);
nor U26631 (N_26631,N_22626,N_23397);
or U26632 (N_26632,N_23631,N_22129);
or U26633 (N_26633,N_22398,N_23849);
or U26634 (N_26634,N_24185,N_21523);
nor U26635 (N_26635,N_23317,N_24851);
or U26636 (N_26636,N_24677,N_24191);
xnor U26637 (N_26637,N_23017,N_20738);
xor U26638 (N_26638,N_22812,N_23371);
or U26639 (N_26639,N_20652,N_22195);
or U26640 (N_26640,N_24734,N_23293);
nor U26641 (N_26641,N_22756,N_23029);
and U26642 (N_26642,N_23057,N_24348);
nor U26643 (N_26643,N_20388,N_20036);
nor U26644 (N_26644,N_23063,N_24405);
and U26645 (N_26645,N_22034,N_21805);
and U26646 (N_26646,N_21587,N_21814);
xor U26647 (N_26647,N_20328,N_20305);
or U26648 (N_26648,N_21675,N_21446);
nor U26649 (N_26649,N_20262,N_20047);
nand U26650 (N_26650,N_21692,N_22189);
or U26651 (N_26651,N_21417,N_20466);
or U26652 (N_26652,N_22785,N_24979);
nor U26653 (N_26653,N_22729,N_20181);
and U26654 (N_26654,N_22060,N_24870);
nand U26655 (N_26655,N_24935,N_23504);
and U26656 (N_26656,N_21643,N_23652);
and U26657 (N_26657,N_20576,N_22027);
or U26658 (N_26658,N_23098,N_22775);
nor U26659 (N_26659,N_22094,N_20208);
xor U26660 (N_26660,N_21062,N_23415);
xor U26661 (N_26661,N_23232,N_20049);
and U26662 (N_26662,N_20923,N_23192);
xor U26663 (N_26663,N_21448,N_21260);
nor U26664 (N_26664,N_23070,N_20785);
or U26665 (N_26665,N_23244,N_24918);
nor U26666 (N_26666,N_22373,N_22597);
and U26667 (N_26667,N_20709,N_20911);
or U26668 (N_26668,N_22789,N_22478);
or U26669 (N_26669,N_23730,N_23521);
or U26670 (N_26670,N_24086,N_23493);
and U26671 (N_26671,N_21966,N_24265);
nor U26672 (N_26672,N_24951,N_22234);
nor U26673 (N_26673,N_23115,N_20603);
nand U26674 (N_26674,N_21635,N_22424);
and U26675 (N_26675,N_24808,N_22456);
nand U26676 (N_26676,N_21799,N_20365);
nor U26677 (N_26677,N_22088,N_20821);
and U26678 (N_26678,N_24197,N_24427);
nand U26679 (N_26679,N_22878,N_22295);
or U26680 (N_26680,N_20304,N_20628);
nor U26681 (N_26681,N_20790,N_22178);
or U26682 (N_26682,N_23854,N_21677);
or U26683 (N_26683,N_24809,N_24004);
nand U26684 (N_26684,N_21230,N_21589);
nor U26685 (N_26685,N_23700,N_21818);
nor U26686 (N_26686,N_24354,N_21458);
nor U26687 (N_26687,N_23831,N_21567);
nor U26688 (N_26688,N_22096,N_21219);
xnor U26689 (N_26689,N_23129,N_22549);
nand U26690 (N_26690,N_22842,N_21596);
nand U26691 (N_26691,N_23825,N_20561);
nor U26692 (N_26692,N_20488,N_22074);
xnor U26693 (N_26693,N_22753,N_20749);
or U26694 (N_26694,N_22796,N_24693);
xor U26695 (N_26695,N_22784,N_22553);
nor U26696 (N_26696,N_24498,N_24130);
or U26697 (N_26697,N_20760,N_24205);
nor U26698 (N_26698,N_23195,N_24173);
nand U26699 (N_26699,N_21548,N_22119);
xnor U26700 (N_26700,N_22047,N_23668);
or U26701 (N_26701,N_21926,N_20544);
or U26702 (N_26702,N_22369,N_23930);
or U26703 (N_26703,N_20650,N_20032);
nand U26704 (N_26704,N_23768,N_22583);
or U26705 (N_26705,N_23438,N_20564);
and U26706 (N_26706,N_23779,N_20396);
nor U26707 (N_26707,N_23675,N_21222);
nand U26708 (N_26708,N_20938,N_23188);
or U26709 (N_26709,N_20108,N_23175);
or U26710 (N_26710,N_24230,N_21723);
nand U26711 (N_26711,N_24053,N_20218);
and U26712 (N_26712,N_22643,N_22216);
nand U26713 (N_26713,N_24577,N_23368);
nor U26714 (N_26714,N_24437,N_20364);
nand U26715 (N_26715,N_20302,N_24085);
xor U26716 (N_26716,N_21162,N_24330);
xor U26717 (N_26717,N_24393,N_21211);
nand U26718 (N_26718,N_20699,N_23898);
xor U26719 (N_26719,N_22128,N_24961);
or U26720 (N_26720,N_23703,N_23247);
nand U26721 (N_26721,N_24382,N_23461);
nand U26722 (N_26722,N_20807,N_21321);
nor U26723 (N_26723,N_24100,N_23976);
or U26724 (N_26724,N_21721,N_20343);
nand U26725 (N_26725,N_22126,N_21636);
nor U26726 (N_26726,N_24087,N_21053);
and U26727 (N_26727,N_22217,N_20467);
and U26728 (N_26728,N_20020,N_23194);
xnor U26729 (N_26729,N_23954,N_21294);
nor U26730 (N_26730,N_22242,N_21275);
and U26731 (N_26731,N_23451,N_20329);
xnor U26732 (N_26732,N_20159,N_22116);
or U26733 (N_26733,N_21394,N_20990);
xnor U26734 (N_26734,N_20154,N_22223);
or U26735 (N_26735,N_22512,N_21387);
or U26736 (N_26736,N_22546,N_24815);
nor U26737 (N_26737,N_20965,N_21045);
nor U26738 (N_26738,N_23673,N_22120);
and U26739 (N_26739,N_23670,N_22741);
nand U26740 (N_26740,N_23806,N_22719);
or U26741 (N_26741,N_20285,N_24887);
nor U26742 (N_26742,N_24699,N_23308);
or U26743 (N_26743,N_24165,N_21825);
or U26744 (N_26744,N_21480,N_22591);
nor U26745 (N_26745,N_20671,N_24195);
nor U26746 (N_26746,N_23294,N_23656);
or U26747 (N_26747,N_20414,N_23110);
xor U26748 (N_26748,N_24983,N_20146);
nand U26749 (N_26749,N_20918,N_22911);
nand U26750 (N_26750,N_22561,N_24861);
nor U26751 (N_26751,N_23177,N_24999);
nand U26752 (N_26752,N_24155,N_22389);
xnor U26753 (N_26753,N_24894,N_23913);
nor U26754 (N_26754,N_21319,N_24765);
or U26755 (N_26755,N_22414,N_23973);
nand U26756 (N_26756,N_23749,N_24251);
and U26757 (N_26757,N_20634,N_21682);
or U26758 (N_26758,N_20838,N_24394);
and U26759 (N_26759,N_20428,N_20635);
nand U26760 (N_26760,N_22073,N_23484);
xor U26761 (N_26761,N_23260,N_23731);
or U26762 (N_26762,N_20307,N_21392);
and U26763 (N_26763,N_22393,N_20884);
and U26764 (N_26764,N_20579,N_20355);
nand U26765 (N_26765,N_24068,N_23047);
or U26766 (N_26766,N_20033,N_24578);
xnor U26767 (N_26767,N_23067,N_21728);
xnor U26768 (N_26768,N_21290,N_20908);
nor U26769 (N_26769,N_22966,N_20323);
nor U26770 (N_26770,N_23344,N_22114);
nor U26771 (N_26771,N_24497,N_23559);
xor U26772 (N_26772,N_24945,N_24160);
nor U26773 (N_26773,N_21038,N_21358);
nand U26774 (N_26774,N_23571,N_20958);
xor U26775 (N_26775,N_22562,N_20088);
and U26776 (N_26776,N_22605,N_20438);
nand U26777 (N_26777,N_22405,N_20383);
or U26778 (N_26778,N_20722,N_24721);
nor U26779 (N_26779,N_20673,N_23804);
and U26780 (N_26780,N_21420,N_22085);
xor U26781 (N_26781,N_23342,N_24680);
or U26782 (N_26782,N_21915,N_23635);
nor U26783 (N_26783,N_21831,N_21492);
xor U26784 (N_26784,N_22865,N_22618);
nor U26785 (N_26785,N_23987,N_20266);
or U26786 (N_26786,N_24500,N_20311);
nand U26787 (N_26787,N_22277,N_20786);
nand U26788 (N_26788,N_24583,N_24367);
nor U26789 (N_26789,N_23947,N_21551);
nor U26790 (N_26790,N_23582,N_20974);
xnor U26791 (N_26791,N_24712,N_20528);
nor U26792 (N_26792,N_23501,N_23467);
and U26793 (N_26793,N_24620,N_23405);
nand U26794 (N_26794,N_22573,N_20538);
nor U26795 (N_26795,N_21267,N_23747);
and U26796 (N_26796,N_23527,N_21405);
or U26797 (N_26797,N_21012,N_23810);
and U26798 (N_26798,N_21097,N_20772);
nor U26799 (N_26799,N_22173,N_23313);
and U26800 (N_26800,N_20963,N_22341);
nand U26801 (N_26801,N_22846,N_21130);
nand U26802 (N_26802,N_22777,N_22943);
and U26803 (N_26803,N_20419,N_22974);
and U26804 (N_26804,N_23231,N_22056);
or U26805 (N_26805,N_20040,N_20553);
nor U26806 (N_26806,N_22379,N_20755);
nor U26807 (N_26807,N_23444,N_23108);
xor U26808 (N_26808,N_20347,N_20067);
nand U26809 (N_26809,N_24188,N_24446);
xor U26810 (N_26810,N_24433,N_22076);
or U26811 (N_26811,N_22654,N_21135);
and U26812 (N_26812,N_20770,N_20046);
nand U26813 (N_26813,N_24991,N_20871);
xnor U26814 (N_26814,N_22319,N_23421);
xnor U26815 (N_26815,N_20275,N_21137);
nor U26816 (N_26816,N_23944,N_23290);
and U26817 (N_26817,N_20525,N_21944);
nor U26818 (N_26818,N_23727,N_21284);
nand U26819 (N_26819,N_23918,N_21383);
nor U26820 (N_26820,N_21702,N_21971);
or U26821 (N_26821,N_23683,N_21376);
nor U26822 (N_26822,N_24730,N_20569);
and U26823 (N_26823,N_21680,N_23514);
or U26824 (N_26824,N_24326,N_22986);
and U26825 (N_26825,N_20783,N_23563);
nand U26826 (N_26826,N_24995,N_20676);
nor U26827 (N_26827,N_23517,N_21898);
xor U26828 (N_26828,N_22247,N_22009);
xnor U26829 (N_26829,N_20037,N_23028);
xnor U26830 (N_26830,N_21697,N_20351);
or U26831 (N_26831,N_23100,N_22436);
and U26832 (N_26832,N_24366,N_22720);
or U26833 (N_26833,N_22751,N_22112);
or U26834 (N_26834,N_21513,N_24946);
nor U26835 (N_26835,N_20142,N_23089);
or U26836 (N_26836,N_22368,N_21367);
nor U26837 (N_26837,N_21634,N_22890);
or U26838 (N_26838,N_24494,N_20868);
nor U26839 (N_26839,N_24050,N_22239);
or U26840 (N_26840,N_23828,N_21072);
or U26841 (N_26841,N_22704,N_20510);
or U26842 (N_26842,N_24849,N_22297);
nor U26843 (N_26843,N_21377,N_23030);
xor U26844 (N_26844,N_22772,N_23352);
nor U26845 (N_26845,N_20334,N_23599);
and U26846 (N_26846,N_21560,N_20252);
xor U26847 (N_26847,N_24516,N_24417);
and U26848 (N_26848,N_21451,N_21777);
nand U26849 (N_26849,N_20465,N_24398);
nor U26850 (N_26850,N_22709,N_20321);
xnor U26851 (N_26851,N_24141,N_23071);
nand U26852 (N_26852,N_21468,N_22274);
nor U26853 (N_26853,N_24219,N_23034);
nand U26854 (N_26854,N_24782,N_23383);
nor U26855 (N_26855,N_22891,N_24376);
and U26856 (N_26856,N_21236,N_24913);
xor U26857 (N_26857,N_20462,N_20793);
nand U26858 (N_26858,N_21329,N_24911);
xor U26859 (N_26859,N_21696,N_23558);
nand U26860 (N_26860,N_21719,N_23202);
and U26861 (N_26861,N_22029,N_24279);
or U26862 (N_26862,N_22566,N_21742);
nor U26863 (N_26863,N_24452,N_21780);
and U26864 (N_26864,N_22163,N_20677);
nor U26865 (N_26865,N_24048,N_22713);
nand U26866 (N_26866,N_24202,N_20949);
or U26867 (N_26867,N_20063,N_20558);
nand U26868 (N_26868,N_20336,N_21402);
nand U26869 (N_26869,N_21667,N_24132);
nand U26870 (N_26870,N_24798,N_22453);
xnor U26871 (N_26871,N_21132,N_20630);
and U26872 (N_26872,N_22089,N_22253);
or U26873 (N_26873,N_24684,N_23978);
nor U26874 (N_26874,N_22682,N_24841);
xnor U26875 (N_26875,N_21121,N_21139);
nand U26876 (N_26876,N_21699,N_24656);
and U26877 (N_26877,N_22245,N_23689);
and U26878 (N_26878,N_20867,N_23402);
nor U26879 (N_26879,N_23853,N_22063);
nor U26880 (N_26880,N_23446,N_21133);
xnor U26881 (N_26881,N_24880,N_23791);
and U26882 (N_26882,N_20748,N_24824);
nand U26883 (N_26883,N_20149,N_22241);
xor U26884 (N_26884,N_22249,N_24608);
xor U26885 (N_26885,N_21585,N_23538);
or U26886 (N_26886,N_23396,N_21999);
xnor U26887 (N_26887,N_20554,N_20147);
and U26888 (N_26888,N_24606,N_24984);
nand U26889 (N_26889,N_24860,N_24743);
xor U26890 (N_26890,N_23445,N_20718);
and U26891 (N_26891,N_23490,N_20536);
or U26892 (N_26892,N_23649,N_24821);
xnor U26893 (N_26893,N_21941,N_21352);
nand U26894 (N_26894,N_23109,N_24364);
or U26895 (N_26895,N_23384,N_21947);
nor U26896 (N_26896,N_22231,N_21949);
xnor U26897 (N_26897,N_22044,N_24630);
xnor U26898 (N_26898,N_24786,N_22358);
nor U26899 (N_26899,N_23716,N_24402);
or U26900 (N_26900,N_22433,N_22805);
or U26901 (N_26901,N_20368,N_23980);
and U26902 (N_26902,N_24866,N_24112);
or U26903 (N_26903,N_24799,N_20775);
nand U26904 (N_26904,N_23487,N_23638);
nor U26905 (N_26905,N_24321,N_20784);
xnor U26906 (N_26906,N_22053,N_23532);
and U26907 (N_26907,N_24460,N_23335);
nand U26908 (N_26908,N_20110,N_23160);
xnor U26909 (N_26909,N_20038,N_21531);
and U26910 (N_26910,N_20636,N_22960);
and U26911 (N_26911,N_23995,N_24459);
nand U26912 (N_26912,N_24492,N_21612);
and U26913 (N_26913,N_21440,N_22613);
and U26914 (N_26914,N_21845,N_22181);
nor U26915 (N_26915,N_22227,N_20166);
nand U26916 (N_26916,N_21185,N_22809);
nand U26917 (N_26917,N_22979,N_24931);
xor U26918 (N_26918,N_24554,N_23201);
nor U26919 (N_26919,N_22962,N_20940);
and U26920 (N_26920,N_21646,N_20859);
or U26921 (N_26921,N_23014,N_21066);
nor U26922 (N_26922,N_20107,N_21313);
and U26923 (N_26923,N_22773,N_20408);
xnor U26924 (N_26924,N_23941,N_20228);
xor U26925 (N_26925,N_24952,N_21171);
and U26926 (N_26926,N_20508,N_24625);
nand U26927 (N_26927,N_23688,N_24363);
xnor U26928 (N_26928,N_24179,N_20075);
or U26929 (N_26929,N_24529,N_20899);
or U26930 (N_26930,N_24103,N_20802);
xor U26931 (N_26931,N_24645,N_23243);
and U26932 (N_26932,N_21023,N_20491);
xor U26933 (N_26933,N_22683,N_22107);
nor U26934 (N_26934,N_24287,N_20777);
and U26935 (N_26935,N_20409,N_20500);
and U26936 (N_26936,N_23454,N_22244);
and U26937 (N_26937,N_24503,N_22110);
nor U26938 (N_26938,N_22445,N_22412);
xnor U26939 (N_26939,N_24683,N_22854);
nand U26940 (N_26940,N_21184,N_20506);
nand U26941 (N_26941,N_24034,N_23239);
and U26942 (N_26942,N_24174,N_22428);
or U26943 (N_26943,N_20239,N_23081);
and U26944 (N_26944,N_20011,N_23211);
nor U26945 (N_26945,N_22350,N_23862);
nor U26946 (N_26946,N_22731,N_24031);
and U26947 (N_26947,N_22403,N_21070);
and U26948 (N_26948,N_21911,N_22603);
xnor U26949 (N_26949,N_22199,N_23621);
xor U26950 (N_26950,N_23803,N_22848);
or U26951 (N_26951,N_21206,N_21486);
nand U26952 (N_26952,N_20943,N_24920);
or U26953 (N_26953,N_20928,N_23553);
xnor U26954 (N_26954,N_21921,N_23829);
nor U26955 (N_26955,N_22435,N_20606);
and U26956 (N_26956,N_22508,N_22233);
xnor U26957 (N_26957,N_20721,N_20688);
nand U26958 (N_26958,N_20946,N_20039);
nand U26959 (N_26959,N_23062,N_20098);
and U26960 (N_26960,N_20764,N_23392);
or U26961 (N_26961,N_24700,N_20233);
xnor U26962 (N_26962,N_20542,N_22977);
and U26963 (N_26963,N_23968,N_22711);
xor U26964 (N_26964,N_21645,N_21295);
and U26965 (N_26965,N_22835,N_23171);
nor U26966 (N_26966,N_21545,N_21931);
nand U26967 (N_26967,N_24547,N_24571);
nand U26968 (N_26968,N_22607,N_20789);
xor U26969 (N_26969,N_20331,N_21046);
nor U26970 (N_26970,N_22822,N_21441);
nor U26971 (N_26971,N_23238,N_20416);
nand U26972 (N_26972,N_21355,N_21316);
nor U26973 (N_26973,N_23215,N_23785);
nor U26974 (N_26974,N_23623,N_20585);
nor U26975 (N_26975,N_22628,N_21018);
and U26976 (N_26976,N_24744,N_22651);
nand U26977 (N_26977,N_23254,N_21356);
nor U26978 (N_26978,N_23564,N_20852);
xnor U26979 (N_26979,N_20207,N_24769);
and U26980 (N_26980,N_22838,N_20062);
or U26981 (N_26981,N_21216,N_24777);
and U26982 (N_26982,N_21108,N_21353);
xnor U26983 (N_26983,N_20927,N_22510);
nor U26984 (N_26984,N_20614,N_24909);
or U26985 (N_26985,N_24907,N_20480);
or U26986 (N_26986,N_23624,N_21017);
or U26987 (N_26987,N_23090,N_23654);
xor U26988 (N_26988,N_22357,N_23182);
or U26989 (N_26989,N_22208,N_23892);
xnor U26990 (N_26990,N_21618,N_21430);
and U26991 (N_26991,N_20298,N_21854);
and U26992 (N_26992,N_24590,N_24535);
xor U26993 (N_26993,N_20241,N_21740);
nor U26994 (N_26994,N_24557,N_22828);
xnor U26995 (N_26995,N_21885,N_20242);
nor U26996 (N_26996,N_22438,N_20436);
xor U26997 (N_26997,N_23302,N_24528);
or U26998 (N_26998,N_20913,N_22318);
nand U26999 (N_26999,N_20014,N_24129);
nand U27000 (N_27000,N_21664,N_22038);
xor U27001 (N_27001,N_23305,N_22205);
and U27002 (N_27002,N_20348,N_21686);
nor U27003 (N_27003,N_24928,N_23227);
xor U27004 (N_27004,N_21197,N_21654);
xnor U27005 (N_27005,N_22998,N_23889);
or U27006 (N_27006,N_20588,N_20970);
nand U27007 (N_27007,N_20637,N_22371);
xnor U27008 (N_27008,N_23874,N_22004);
nor U27009 (N_27009,N_22576,N_22169);
or U27010 (N_27010,N_21269,N_22059);
or U27011 (N_27011,N_21179,N_23311);
nand U27012 (N_27012,N_21407,N_24605);
and U27013 (N_27013,N_20077,N_20069);
nor U27014 (N_27014,N_21965,N_24080);
nand U27015 (N_27015,N_21148,N_22102);
nand U27016 (N_27016,N_22210,N_21425);
xnor U27017 (N_27017,N_23725,N_23931);
and U27018 (N_27018,N_20245,N_22043);
nand U27019 (N_27019,N_24504,N_23470);
and U27020 (N_27020,N_23353,N_20274);
nor U27021 (N_27021,N_22750,N_20982);
nand U27022 (N_27022,N_21715,N_20292);
nand U27023 (N_27023,N_20453,N_24820);
nand U27024 (N_27024,N_21628,N_21482);
nor U27025 (N_27025,N_24449,N_23745);
nand U27026 (N_27026,N_23859,N_22471);
nand U27027 (N_27027,N_23632,N_20812);
xor U27028 (N_27028,N_24254,N_21866);
and U27029 (N_27029,N_21395,N_23151);
nand U27030 (N_27030,N_24561,N_20330);
xnor U27031 (N_27031,N_20468,N_22680);
or U27032 (N_27032,N_21428,N_23173);
and U27033 (N_27033,N_23361,N_22502);
or U27034 (N_27034,N_22290,N_21212);
nand U27035 (N_27035,N_24410,N_20185);
or U27036 (N_27036,N_24550,N_22645);
xnor U27037 (N_27037,N_20968,N_21659);
xnor U27038 (N_27038,N_24131,N_20771);
nand U27039 (N_27039,N_22937,N_24971);
nor U27040 (N_27040,N_22139,N_20163);
and U27041 (N_27041,N_22622,N_21750);
or U27042 (N_27042,N_22439,N_20084);
nor U27043 (N_27043,N_23569,N_22226);
and U27044 (N_27044,N_23485,N_23897);
nor U27045 (N_27045,N_22051,N_24708);
nand U27046 (N_27046,N_20566,N_24317);
nor U27047 (N_27047,N_24926,N_24704);
and U27048 (N_27048,N_22401,N_23356);
nand U27049 (N_27049,N_22710,N_24306);
nand U27050 (N_27050,N_21769,N_24210);
and U27051 (N_27051,N_23502,N_21724);
or U27052 (N_27052,N_20795,N_22511);
xor U27053 (N_27053,N_24714,N_24125);
nand U27054 (N_27054,N_24392,N_22140);
xnor U27055 (N_27055,N_21834,N_24843);
xnor U27056 (N_27056,N_22938,N_24511);
xnor U27057 (N_27057,N_21954,N_23132);
xor U27058 (N_27058,N_21051,N_24711);
xnor U27059 (N_27059,N_24740,N_24154);
or U27060 (N_27060,N_23718,N_23498);
nand U27061 (N_27061,N_23578,N_22317);
xor U27062 (N_27062,N_21568,N_23692);
nand U27063 (N_27063,N_24421,N_24419);
and U27064 (N_27064,N_21514,N_21767);
nand U27065 (N_27065,N_20873,N_22781);
nor U27066 (N_27066,N_22803,N_21899);
nor U27067 (N_27067,N_23883,N_23146);
nand U27068 (N_27068,N_24258,N_24198);
xnor U27069 (N_27069,N_20140,N_21074);
and U27070 (N_27070,N_23349,N_21478);
or U27071 (N_27071,N_23781,N_24090);
xor U27072 (N_27072,N_21610,N_21297);
and U27073 (N_27073,N_20930,N_21380);
nor U27074 (N_27074,N_23724,N_21860);
and U27075 (N_27075,N_22687,N_21153);
xnor U27076 (N_27076,N_21200,N_23085);
and U27077 (N_27077,N_21142,N_24694);
nand U27078 (N_27078,N_20225,N_21807);
nor U27079 (N_27079,N_21081,N_21221);
and U27080 (N_27080,N_24424,N_22575);
nand U27081 (N_27081,N_21099,N_24747);
and U27082 (N_27082,N_23929,N_20379);
nor U27083 (N_27083,N_22956,N_24252);
nor U27084 (N_27084,N_23120,N_22207);
or U27085 (N_27085,N_22272,N_23693);
xor U27086 (N_27086,N_24857,N_20681);
nand U27087 (N_27087,N_23702,N_22146);
nor U27088 (N_27088,N_23419,N_22930);
or U27089 (N_27089,N_24456,N_23894);
xnor U27090 (N_27090,N_24439,N_21579);
or U27091 (N_27091,N_23723,N_21122);
xnor U27092 (N_27092,N_24423,N_20996);
xor U27093 (N_27093,N_23983,N_21519);
nor U27094 (N_27094,N_20008,N_22852);
or U27095 (N_27095,N_22526,N_21496);
nand U27096 (N_27096,N_20445,N_21875);
nor U27097 (N_27097,N_24186,N_22015);
nor U27098 (N_27098,N_23795,N_21141);
or U27099 (N_27099,N_24104,N_22858);
xor U27100 (N_27100,N_23709,N_23106);
and U27101 (N_27101,N_20369,N_21872);
and U27102 (N_27102,N_23410,N_22904);
or U27103 (N_27103,N_23576,N_21678);
nor U27104 (N_27104,N_21573,N_22652);
xnor U27105 (N_27105,N_21308,N_24268);
nand U27106 (N_27106,N_22012,N_23496);
nand U27107 (N_27107,N_21438,N_21539);
and U27108 (N_27108,N_24923,N_20933);
xor U27109 (N_27109,N_24167,N_21047);
nand U27110 (N_27110,N_23659,N_22092);
xor U27111 (N_27111,N_24657,N_21553);
nor U27112 (N_27112,N_23237,N_22896);
and U27113 (N_27113,N_20205,N_24175);
and U27114 (N_27114,N_23186,N_23035);
nand U27115 (N_27115,N_21533,N_20267);
nor U27116 (N_27116,N_21232,N_22917);
nand U27117 (N_27117,N_20975,N_20021);
nand U27118 (N_27118,N_24057,N_24761);
or U27119 (N_27119,N_24114,N_21489);
or U27120 (N_27120,N_23904,N_22826);
xnor U27121 (N_27121,N_21415,N_21998);
nand U27122 (N_27122,N_21668,N_24232);
or U27123 (N_27123,N_23556,N_24072);
or U27124 (N_27124,N_20291,N_22266);
xnor U27125 (N_27125,N_23697,N_23279);
nand U27126 (N_27126,N_21790,N_21752);
and U27127 (N_27127,N_20702,N_24639);
nand U27128 (N_27128,N_24558,N_24455);
and U27129 (N_27129,N_22091,N_20660);
nor U27130 (N_27130,N_21788,N_22066);
and U27131 (N_27131,N_22669,N_22331);
nand U27132 (N_27132,N_21476,N_21109);
xor U27133 (N_27133,N_21138,N_22147);
and U27134 (N_27134,N_22097,N_22499);
and U27135 (N_27135,N_23914,N_22760);
and U27136 (N_27136,N_22918,N_23022);
or U27137 (N_27137,N_24135,N_22143);
and U27138 (N_27138,N_23827,N_21299);
xor U27139 (N_27139,N_24582,N_24534);
or U27140 (N_27140,N_22268,N_22170);
nor U27141 (N_27141,N_21663,N_23870);
nor U27142 (N_27142,N_23178,N_21527);
nor U27143 (N_27143,N_21210,N_23587);
or U27144 (N_27144,N_23864,N_22745);
nand U27145 (N_27145,N_22289,N_20803);
nor U27146 (N_27146,N_21945,N_20866);
nor U27147 (N_27147,N_22504,N_21768);
xnor U27148 (N_27148,N_20418,N_23525);
nand U27149 (N_27149,N_24853,N_24311);
nor U27150 (N_27150,N_24591,N_21011);
or U27151 (N_27151,N_20691,N_23515);
nand U27152 (N_27152,N_24724,N_23896);
nor U27153 (N_27153,N_21935,N_20960);
nor U27154 (N_27154,N_22712,N_23226);
nor U27155 (N_27155,N_21401,N_21572);
or U27156 (N_27156,N_24145,N_21653);
nor U27157 (N_27157,N_24231,N_23010);
xnor U27158 (N_27158,N_20366,N_23212);
xnor U27159 (N_27159,N_24871,N_22093);
xnor U27160 (N_27160,N_24334,N_21580);
xnor U27161 (N_27161,N_20064,N_23817);
xnor U27162 (N_27162,N_22345,N_21060);
xor U27163 (N_27163,N_24867,N_20925);
nand U27164 (N_27164,N_22920,N_20773);
nor U27165 (N_27165,N_20559,N_22185);
nand U27166 (N_27166,N_20915,N_20667);
xor U27167 (N_27167,N_24934,N_23213);
or U27168 (N_27168,N_20447,N_24200);
or U27169 (N_27169,N_20319,N_20178);
nor U27170 (N_27170,N_24082,N_23049);
nand U27171 (N_27171,N_21079,N_21020);
nand U27172 (N_27172,N_21026,N_21882);
and U27173 (N_27173,N_22127,N_21536);
xor U27174 (N_27174,N_21726,N_24762);
or U27175 (N_27175,N_22670,N_21803);
nor U27176 (N_27176,N_22019,N_20345);
or U27177 (N_27177,N_23300,N_21144);
nand U27178 (N_27178,N_22375,N_23130);
and U27179 (N_27179,N_23905,N_23468);
or U27180 (N_27180,N_22150,N_22214);
xnor U27181 (N_27181,N_23155,N_24587);
nor U27182 (N_27182,N_23142,N_23200);
and U27183 (N_27183,N_23590,N_24028);
and U27184 (N_27184,N_22134,N_21256);
xor U27185 (N_27185,N_21961,N_21936);
and U27186 (N_27186,N_21537,N_24329);
nor U27187 (N_27187,N_20125,N_20549);
nor U27188 (N_27188,N_20936,N_23295);
nor U27189 (N_27189,N_20143,N_24513);
nor U27190 (N_27190,N_20013,N_22948);
nand U27191 (N_27191,N_24519,N_22582);
nand U27192 (N_27192,N_22190,N_20719);
xor U27193 (N_27193,N_20507,N_20639);
and U27194 (N_27194,N_24771,N_21706);
xor U27195 (N_27195,N_24755,N_23784);
nand U27196 (N_27196,N_23919,N_20799);
xnor U27197 (N_27197,N_24044,N_20071);
and U27198 (N_27198,N_23050,N_20437);
nor U27199 (N_27199,N_22406,N_21306);
or U27200 (N_27200,N_20315,N_24349);
or U27201 (N_27201,N_21126,N_23347);
nand U27202 (N_27202,N_24307,N_21239);
nand U27203 (N_27203,N_22161,N_22625);
nor U27204 (N_27204,N_22876,N_24689);
xor U27205 (N_27205,N_20479,N_23714);
xor U27206 (N_27206,N_21449,N_24842);
and U27207 (N_27207,N_24805,N_20568);
xor U27208 (N_27208,N_23497,N_23039);
xor U27209 (N_27209,N_22969,N_21502);
or U27210 (N_27210,N_22807,N_21992);
xor U27211 (N_27211,N_22017,N_24539);
xor U27212 (N_27212,N_21960,N_21310);
or U27213 (N_27213,N_23214,N_22200);
or U27214 (N_27214,N_21713,N_21300);
nor U27215 (N_27215,N_24674,N_24720);
and U27216 (N_27216,N_21688,N_20231);
or U27217 (N_27217,N_22684,N_21307);
xor U27218 (N_27218,N_24850,N_20680);
or U27219 (N_27219,N_23637,N_22590);
nand U27220 (N_27220,N_24800,N_21522);
or U27221 (N_27221,N_24212,N_24241);
nor U27222 (N_27222,N_24108,N_21801);
nand U27223 (N_27223,N_21408,N_21632);
nand U27224 (N_27224,N_21342,N_22620);
and U27225 (N_27225,N_24629,N_23076);
nor U27226 (N_27226,N_20370,N_23193);
nand U27227 (N_27227,N_24588,N_24435);
nor U27228 (N_27228,N_24536,N_21765);
or U27229 (N_27229,N_24731,N_23256);
or U27230 (N_27230,N_24705,N_22763);
and U27231 (N_27231,N_20665,N_20410);
and U27232 (N_27232,N_22014,N_20156);
or U27233 (N_27233,N_21225,N_21883);
and U27234 (N_27234,N_24380,N_21816);
nand U27235 (N_27235,N_24962,N_21490);
nor U27236 (N_27236,N_22536,N_24177);
and U27237 (N_27237,N_23977,N_24172);
nor U27238 (N_27238,N_24216,N_22647);
nor U27239 (N_27239,N_21836,N_21503);
nand U27240 (N_27240,N_22916,N_24653);
and U27241 (N_27241,N_21939,N_20173);
xor U27242 (N_27242,N_22872,N_24260);
xnor U27243 (N_27243,N_21000,N_24011);
nor U27244 (N_27244,N_23241,N_22283);
and U27245 (N_27245,N_24745,N_24613);
and U27246 (N_27246,N_23720,N_22138);
or U27247 (N_27247,N_24487,N_22351);
nand U27248 (N_27248,N_24272,N_24215);
or U27249 (N_27249,N_20427,N_23059);
nor U27250 (N_27250,N_20604,N_20993);
xor U27251 (N_27251,N_23766,N_23320);
and U27252 (N_27252,N_20121,N_20633);
or U27253 (N_27253,N_24986,N_20382);
or U27254 (N_27254,N_22132,N_20713);
xor U27255 (N_27255,N_24387,N_23956);
nand U27256 (N_27256,N_22663,N_23348);
and U27257 (N_27257,N_21149,N_20354);
nand U27258 (N_27258,N_24067,N_20024);
nor U27259 (N_27259,N_20632,N_21727);
nor U27260 (N_27260,N_24856,N_21096);
and U27261 (N_27261,N_21460,N_21288);
nand U27262 (N_27262,N_22311,N_24353);
nor U27263 (N_27263,N_23053,N_23457);
xnor U27264 (N_27264,N_23046,N_20340);
xnor U27265 (N_27265,N_23916,N_20359);
or U27266 (N_27266,N_21930,N_23267);
nor U27267 (N_27267,N_22343,N_22131);
or U27268 (N_27268,N_24470,N_20268);
xor U27269 (N_27269,N_24807,N_22402);
and U27270 (N_27270,N_23866,N_22814);
xnor U27271 (N_27271,N_24332,N_24257);
nand U27272 (N_27272,N_22382,N_22390);
nor U27273 (N_27273,N_23011,N_22717);
and U27274 (N_27274,N_24386,N_22049);
nor U27275 (N_27275,N_22101,N_22399);
and U27276 (N_27276,N_21291,N_22479);
nand U27277 (N_27277,N_20219,N_24864);
and U27278 (N_27278,N_24001,N_23626);
or U27279 (N_27279,N_20539,N_24748);
nand U27280 (N_27280,N_21658,N_22003);
and U27281 (N_27281,N_23863,N_24672);
xnor U27282 (N_27282,N_24153,N_24007);
nor U27283 (N_27283,N_22156,N_22167);
and U27284 (N_27284,N_20150,N_24164);
nor U27285 (N_27285,N_23327,N_24958);
nor U27286 (N_27286,N_21248,N_24933);
nand U27287 (N_27287,N_20058,N_21202);
nor U27288 (N_27288,N_24949,N_20157);
and U27289 (N_27289,N_22522,N_22033);
xor U27290 (N_27290,N_22929,N_22700);
nor U27291 (N_27291,N_23145,N_21063);
and U27292 (N_27292,N_24293,N_20183);
or U27293 (N_27293,N_24604,N_21734);
nor U27294 (N_27294,N_23712,N_23386);
xnor U27295 (N_27295,N_21271,N_22532);
or U27296 (N_27296,N_24733,N_24365);
xnor U27297 (N_27297,N_22537,N_24483);
nor U27298 (N_27298,N_23737,N_23086);
and U27299 (N_27299,N_23622,N_24736);
or U27300 (N_27300,N_21782,N_20922);
nor U27301 (N_27301,N_20954,N_23198);
nand U27302 (N_27302,N_20322,N_20754);
nand U27303 (N_27303,N_20727,N_22058);
or U27304 (N_27304,N_24617,N_21048);
or U27305 (N_27305,N_22901,N_20531);
or U27306 (N_27306,N_20372,N_21665);
nor U27307 (N_27307,N_23282,N_21808);
xor U27308 (N_27308,N_22324,N_20155);
nand U27309 (N_27309,N_21778,N_20174);
nand U27310 (N_27310,N_21301,N_20683);
xor U27311 (N_27311,N_24641,N_24685);
nor U27312 (N_27312,N_24510,N_20471);
xnor U27313 (N_27313,N_21054,N_20189);
xor U27314 (N_27314,N_21204,N_20823);
and U27315 (N_27315,N_22099,N_24636);
and U27316 (N_27316,N_21255,N_20381);
or U27317 (N_27317,N_23234,N_21494);
or U27318 (N_27318,N_21540,N_20584);
nand U27319 (N_27319,N_20035,N_20697);
nand U27320 (N_27320,N_24399,N_21839);
xor U27321 (N_27321,N_21444,N_23138);
and U27322 (N_27322,N_20747,N_21331);
and U27323 (N_27323,N_20213,N_20995);
nor U27324 (N_27324,N_23378,N_21981);
and U27325 (N_27325,N_24070,N_24879);
xor U27326 (N_27326,N_24538,N_22988);
xor U27327 (N_27327,N_21569,N_24077);
nand U27328 (N_27328,N_21474,N_21309);
and U27329 (N_27329,N_23546,N_21147);
and U27330 (N_27330,N_23551,N_24750);
and U27331 (N_27331,N_24297,N_21804);
and U27332 (N_27332,N_23297,N_24285);
nor U27333 (N_27333,N_21433,N_23544);
and U27334 (N_27334,N_20397,N_24707);
or U27335 (N_27335,N_22548,N_21101);
nor U27336 (N_27336,N_20015,N_24847);
and U27337 (N_27337,N_22355,N_22055);
and U27338 (N_27338,N_24281,N_20509);
xor U27339 (N_27339,N_22260,N_21413);
or U27340 (N_27340,N_23429,N_20357);
nor U27341 (N_27341,N_24235,N_20850);
and U27342 (N_27342,N_23271,N_23650);
or U27343 (N_27343,N_21571,N_20948);
xnor U27344 (N_27344,N_23097,N_24548);
xor U27345 (N_27345,N_22701,N_20206);
and U27346 (N_27346,N_22791,N_22005);
or U27347 (N_27347,N_22385,N_23473);
and U27348 (N_27348,N_20750,N_24589);
xnor U27349 (N_27349,N_20141,N_20217);
xnor U27350 (N_27350,N_24038,N_22637);
nor U27351 (N_27351,N_23209,N_21755);
xor U27352 (N_27352,N_24491,N_23572);
and U27353 (N_27353,N_20018,N_24406);
or U27354 (N_27354,N_22888,N_23742);
xor U27355 (N_27355,N_21131,N_20621);
or U27356 (N_27356,N_24035,N_24631);
xor U27357 (N_27357,N_20199,N_23453);
nor U27358 (N_27358,N_21270,N_21509);
xnor U27359 (N_27359,N_20813,N_20675);
or U27360 (N_27360,N_20988,N_23441);
nor U27361 (N_27361,N_20851,N_24937);
or U27362 (N_27362,N_20448,N_22738);
and U27363 (N_27363,N_23204,N_23025);
or U27364 (N_27364,N_20895,N_23316);
xnor U27365 (N_27365,N_23658,N_22263);
nand U27366 (N_27366,N_23878,N_20111);
nor U27367 (N_27367,N_22006,N_22847);
xor U27368 (N_27368,N_23372,N_20725);
or U27369 (N_27369,N_21691,N_21968);
nor U27370 (N_27370,N_21080,N_23210);
nand U27371 (N_27371,N_21759,N_22627);
xor U27372 (N_27372,N_24020,N_21627);
and U27373 (N_27373,N_24273,N_20030);
nand U27374 (N_27374,N_24963,N_21785);
and U27375 (N_27375,N_22465,N_22623);
nor U27376 (N_27376,N_21744,N_22133);
or U27377 (N_27377,N_21276,N_23170);
xnor U27378 (N_27378,N_22824,N_24222);
or U27379 (N_27379,N_20998,N_24757);
and U27380 (N_27380,N_20698,N_21774);
xor U27381 (N_27381,N_23690,N_20277);
nor U27382 (N_27382,N_24403,N_22790);
nor U27383 (N_27383,N_21421,N_23082);
and U27384 (N_27384,N_20931,N_21457);
or U27385 (N_27385,N_24194,N_24445);
nand U27386 (N_27386,N_22279,N_20393);
and U27387 (N_27387,N_20752,N_23099);
xor U27388 (N_27388,N_21488,N_21499);
and U27389 (N_27389,N_24776,N_22480);
nand U27390 (N_27390,N_21524,N_20563);
xor U27391 (N_27391,N_22152,N_20495);
xnor U27392 (N_27392,N_22932,N_22024);
nor U27393 (N_27393,N_22655,N_23103);
xnor U27394 (N_27394,N_21418,N_24784);
and U27395 (N_27395,N_22108,N_23134);
nand U27396 (N_27396,N_20582,N_24466);
or U27397 (N_27397,N_20597,N_21762);
or U27398 (N_27398,N_20912,N_21881);
xnor U27399 (N_27399,N_20815,N_24388);
xnor U27400 (N_27400,N_21575,N_24256);
xnor U27401 (N_27401,N_21789,N_21006);
nor U27402 (N_27402,N_21991,N_23952);
nor U27403 (N_27403,N_23881,N_24404);
xor U27404 (N_27404,N_22941,N_24970);
or U27405 (N_27405,N_23088,N_24451);
or U27406 (N_27406,N_24916,N_21203);
nor U27407 (N_27407,N_21950,N_24602);
xor U27408 (N_27408,N_23597,N_21984);
xnor U27409 (N_27409,N_22326,N_21925);
or U27410 (N_27410,N_20640,N_24764);
and U27411 (N_27411,N_24830,N_24715);
nand U27412 (N_27412,N_21876,N_20798);
and U27413 (N_27413,N_24193,N_20717);
xor U27414 (N_27414,N_21242,N_21661);
or U27415 (N_27415,N_22706,N_20076);
or U27416 (N_27416,N_22372,N_21016);
and U27417 (N_27417,N_21003,N_24438);
and U27418 (N_27418,N_22472,N_21798);
or U27419 (N_27419,N_22595,N_22574);
and U27420 (N_27420,N_21049,N_22307);
xnor U27421 (N_27421,N_21059,N_23183);
and U27422 (N_27422,N_22111,N_23677);
xnor U27423 (N_27423,N_23765,N_20027);
or U27424 (N_27424,N_22671,N_23591);
and U27425 (N_27425,N_24115,N_22209);
nand U27426 (N_27426,N_23489,N_20545);
nor U27427 (N_27427,N_21459,N_22610);
or U27428 (N_27428,N_20599,N_21516);
or U27429 (N_27429,N_24718,N_24170);
xnor U27430 (N_27430,N_22653,N_23917);
xnor U27431 (N_27431,N_20451,N_20290);
nor U27432 (N_27432,N_23483,N_22374);
or U27433 (N_27433,N_22764,N_24416);
and U27434 (N_27434,N_21436,N_20358);
xor U27435 (N_27435,N_20696,N_21015);
nand U27436 (N_27436,N_23112,N_21287);
nor U27437 (N_27437,N_20057,N_23991);
nor U27438 (N_27438,N_23577,N_23782);
xor U27439 (N_27439,N_22978,N_23042);
or U27440 (N_27440,N_22644,N_22270);
nor U27441 (N_27441,N_21687,N_22676);
xor U27442 (N_27442,N_23946,N_23258);
or U27443 (N_27443,N_24345,N_23655);
nor U27444 (N_27444,N_21795,N_21470);
nand U27445 (N_27445,N_21914,N_24767);
or U27446 (N_27446,N_20845,N_24595);
xnor U27447 (N_27447,N_23281,N_21995);
or U27448 (N_27448,N_22873,N_20446);
xnor U27449 (N_27449,N_23696,N_23605);
nor U27450 (N_27450,N_22660,N_21107);
and U27451 (N_27451,N_22422,N_24315);
nor U27452 (N_27452,N_20119,N_22124);
nand U27453 (N_27453,N_21400,N_24523);
or U27454 (N_27454,N_23647,N_22115);
nand U27455 (N_27455,N_20288,N_24083);
and U27456 (N_27456,N_24124,N_23073);
nor U27457 (N_27457,N_22298,N_24992);
or U27458 (N_27458,N_24187,N_21234);
or U27459 (N_27459,N_20258,N_20516);
nand U27460 (N_27460,N_20299,N_22621);
or U27461 (N_27461,N_21337,N_20261);
or U27462 (N_27462,N_20619,N_24357);
nand U27463 (N_27463,N_23565,N_20766);
and U27464 (N_27464,N_23594,N_23373);
or U27465 (N_27465,N_22535,N_20490);
or U27466 (N_27466,N_20317,N_23176);
or U27467 (N_27467,N_22716,N_22069);
nand U27468 (N_27468,N_22154,N_22922);
xor U27469 (N_27469,N_20109,N_24666);
xor U27470 (N_27470,N_23732,N_23401);
and U27471 (N_27471,N_21412,N_21756);
or U27472 (N_27472,N_22000,N_21561);
nand U27473 (N_27473,N_21296,N_24218);
and U27474 (N_27474,N_20810,N_22046);
nand U27475 (N_27475,N_23764,N_21973);
nor U27476 (N_27476,N_22778,N_23364);
and U27477 (N_27477,N_22586,N_24825);
and U27478 (N_27478,N_21253,N_20371);
and U27479 (N_27479,N_21422,N_22002);
and U27480 (N_27480,N_23628,N_23370);
nor U27481 (N_27481,N_24914,N_21770);
xnor U27482 (N_27482,N_24915,N_22265);
nand U27483 (N_27483,N_21671,N_22481);
nor U27484 (N_27484,N_20153,N_23744);
nor U27485 (N_27485,N_20230,N_24102);
and U27486 (N_27486,N_22462,N_22285);
and U27487 (N_27487,N_24753,N_22477);
and U27488 (N_27488,N_21542,N_22328);
nor U27489 (N_27489,N_24341,N_24314);
nand U27490 (N_27490,N_20555,N_22278);
xnor U27491 (N_27491,N_22367,N_24302);
xor U27492 (N_27492,N_21100,N_24203);
xor U27493 (N_27493,N_22342,N_20431);
nand U27494 (N_27494,N_24522,N_20994);
or U27495 (N_27495,N_23221,N_22892);
or U27496 (N_27496,N_22993,N_22294);
and U27497 (N_27497,N_22619,N_23431);
and U27498 (N_27498,N_23844,N_24432);
and U27499 (N_27499,N_22823,N_22236);
xnor U27500 (N_27500,N_22436,N_23948);
and U27501 (N_27501,N_21476,N_23726);
nor U27502 (N_27502,N_22244,N_23402);
nand U27503 (N_27503,N_23756,N_21084);
nand U27504 (N_27504,N_23392,N_22675);
xor U27505 (N_27505,N_21513,N_23764);
or U27506 (N_27506,N_22287,N_21234);
nor U27507 (N_27507,N_20169,N_23368);
or U27508 (N_27508,N_24465,N_22402);
nand U27509 (N_27509,N_24614,N_24070);
nor U27510 (N_27510,N_23881,N_23388);
xnor U27511 (N_27511,N_21596,N_23045);
or U27512 (N_27512,N_22150,N_22324);
and U27513 (N_27513,N_23903,N_23176);
and U27514 (N_27514,N_21357,N_24938);
or U27515 (N_27515,N_24841,N_22037);
xnor U27516 (N_27516,N_24816,N_21608);
nor U27517 (N_27517,N_24754,N_22822);
xnor U27518 (N_27518,N_20659,N_20929);
or U27519 (N_27519,N_21857,N_20907);
nand U27520 (N_27520,N_21238,N_21255);
nor U27521 (N_27521,N_20183,N_21243);
nor U27522 (N_27522,N_20722,N_24872);
nor U27523 (N_27523,N_21788,N_24972);
or U27524 (N_27524,N_20018,N_22741);
and U27525 (N_27525,N_21774,N_20985);
nand U27526 (N_27526,N_21630,N_23515);
nand U27527 (N_27527,N_21040,N_20349);
or U27528 (N_27528,N_20711,N_24430);
and U27529 (N_27529,N_21284,N_23999);
or U27530 (N_27530,N_23218,N_22072);
nor U27531 (N_27531,N_20902,N_22531);
nand U27532 (N_27532,N_21757,N_20191);
nor U27533 (N_27533,N_21988,N_23063);
nand U27534 (N_27534,N_23791,N_22527);
xor U27535 (N_27535,N_20964,N_24796);
xnor U27536 (N_27536,N_22293,N_20588);
nand U27537 (N_27537,N_20445,N_21623);
nor U27538 (N_27538,N_24654,N_21898);
and U27539 (N_27539,N_20767,N_21851);
nand U27540 (N_27540,N_23880,N_21148);
nor U27541 (N_27541,N_20812,N_23223);
or U27542 (N_27542,N_22102,N_23571);
or U27543 (N_27543,N_22968,N_24153);
and U27544 (N_27544,N_23213,N_22981);
and U27545 (N_27545,N_21097,N_22193);
xor U27546 (N_27546,N_24161,N_22573);
and U27547 (N_27547,N_20489,N_20741);
nor U27548 (N_27548,N_20399,N_20373);
or U27549 (N_27549,N_22988,N_24207);
xor U27550 (N_27550,N_22890,N_24711);
xor U27551 (N_27551,N_23851,N_23599);
nor U27552 (N_27552,N_23365,N_23568);
nor U27553 (N_27553,N_20036,N_20073);
or U27554 (N_27554,N_21989,N_22099);
nor U27555 (N_27555,N_22434,N_20398);
or U27556 (N_27556,N_23073,N_22849);
or U27557 (N_27557,N_20299,N_23935);
xor U27558 (N_27558,N_24456,N_21763);
and U27559 (N_27559,N_24131,N_20017);
xnor U27560 (N_27560,N_24894,N_20274);
xnor U27561 (N_27561,N_20306,N_22267);
and U27562 (N_27562,N_20316,N_20019);
nand U27563 (N_27563,N_23069,N_23601);
nor U27564 (N_27564,N_21533,N_23738);
and U27565 (N_27565,N_24829,N_20661);
nor U27566 (N_27566,N_20277,N_22409);
nor U27567 (N_27567,N_23467,N_21019);
and U27568 (N_27568,N_20552,N_22687);
xnor U27569 (N_27569,N_22493,N_20758);
nor U27570 (N_27570,N_21257,N_21493);
and U27571 (N_27571,N_23869,N_24822);
nand U27572 (N_27572,N_22862,N_21970);
xnor U27573 (N_27573,N_24050,N_23182);
nand U27574 (N_27574,N_22044,N_21897);
nand U27575 (N_27575,N_21200,N_21952);
nand U27576 (N_27576,N_21137,N_22275);
nand U27577 (N_27577,N_23660,N_21496);
nor U27578 (N_27578,N_23525,N_21402);
nor U27579 (N_27579,N_22701,N_24190);
or U27580 (N_27580,N_22141,N_24747);
and U27581 (N_27581,N_22640,N_21356);
nor U27582 (N_27582,N_20549,N_20350);
or U27583 (N_27583,N_20835,N_24454);
and U27584 (N_27584,N_22496,N_20484);
and U27585 (N_27585,N_20673,N_20244);
or U27586 (N_27586,N_20036,N_23696);
or U27587 (N_27587,N_24423,N_22322);
xnor U27588 (N_27588,N_20457,N_20648);
xnor U27589 (N_27589,N_24760,N_23169);
or U27590 (N_27590,N_20300,N_21398);
and U27591 (N_27591,N_24941,N_22586);
and U27592 (N_27592,N_20156,N_23441);
or U27593 (N_27593,N_22621,N_21429);
xor U27594 (N_27594,N_21360,N_24249);
nand U27595 (N_27595,N_24828,N_20347);
and U27596 (N_27596,N_21538,N_24034);
nand U27597 (N_27597,N_21486,N_23899);
xor U27598 (N_27598,N_21533,N_22531);
nor U27599 (N_27599,N_24691,N_20391);
or U27600 (N_27600,N_22915,N_20304);
xnor U27601 (N_27601,N_23442,N_23572);
and U27602 (N_27602,N_22026,N_22707);
xnor U27603 (N_27603,N_23472,N_21118);
nor U27604 (N_27604,N_24402,N_23576);
or U27605 (N_27605,N_21357,N_20373);
nor U27606 (N_27606,N_23272,N_23157);
xnor U27607 (N_27607,N_21927,N_22012);
nor U27608 (N_27608,N_21343,N_23448);
xor U27609 (N_27609,N_24828,N_21280);
xnor U27610 (N_27610,N_21097,N_22929);
xnor U27611 (N_27611,N_21295,N_20811);
nand U27612 (N_27612,N_23056,N_20321);
and U27613 (N_27613,N_20300,N_21390);
xor U27614 (N_27614,N_24950,N_22154);
xor U27615 (N_27615,N_20170,N_21058);
and U27616 (N_27616,N_23212,N_24960);
or U27617 (N_27617,N_21923,N_21964);
nand U27618 (N_27618,N_23499,N_22664);
nor U27619 (N_27619,N_24950,N_22614);
and U27620 (N_27620,N_20618,N_23045);
nor U27621 (N_27621,N_24777,N_20458);
xnor U27622 (N_27622,N_21614,N_22239);
or U27623 (N_27623,N_24967,N_23470);
and U27624 (N_27624,N_20433,N_24529);
xor U27625 (N_27625,N_24825,N_24349);
or U27626 (N_27626,N_23175,N_23910);
xnor U27627 (N_27627,N_22966,N_20389);
and U27628 (N_27628,N_21596,N_24812);
xnor U27629 (N_27629,N_23664,N_20419);
nor U27630 (N_27630,N_23827,N_24061);
and U27631 (N_27631,N_23606,N_24897);
xor U27632 (N_27632,N_20377,N_23332);
and U27633 (N_27633,N_23654,N_24182);
nand U27634 (N_27634,N_21032,N_20282);
or U27635 (N_27635,N_21929,N_21084);
xor U27636 (N_27636,N_24566,N_23886);
xor U27637 (N_27637,N_24713,N_23651);
and U27638 (N_27638,N_22095,N_23718);
and U27639 (N_27639,N_22513,N_21019);
and U27640 (N_27640,N_21255,N_24567);
or U27641 (N_27641,N_24964,N_21682);
xor U27642 (N_27642,N_21359,N_22294);
xnor U27643 (N_27643,N_20972,N_23154);
nand U27644 (N_27644,N_20443,N_20078);
nand U27645 (N_27645,N_20141,N_24781);
nand U27646 (N_27646,N_21116,N_21842);
nor U27647 (N_27647,N_21502,N_24339);
or U27648 (N_27648,N_21415,N_22626);
xnor U27649 (N_27649,N_24107,N_24425);
or U27650 (N_27650,N_20801,N_23064);
nor U27651 (N_27651,N_23759,N_24879);
nand U27652 (N_27652,N_24754,N_23529);
xnor U27653 (N_27653,N_21196,N_21594);
and U27654 (N_27654,N_24954,N_20110);
nor U27655 (N_27655,N_21924,N_21740);
and U27656 (N_27656,N_22488,N_22039);
xor U27657 (N_27657,N_24529,N_23810);
or U27658 (N_27658,N_23338,N_24185);
and U27659 (N_27659,N_22468,N_23271);
nor U27660 (N_27660,N_23819,N_22084);
and U27661 (N_27661,N_23284,N_23566);
nor U27662 (N_27662,N_23528,N_23950);
or U27663 (N_27663,N_24067,N_24407);
nand U27664 (N_27664,N_23024,N_23280);
nor U27665 (N_27665,N_24161,N_24268);
and U27666 (N_27666,N_20542,N_24515);
and U27667 (N_27667,N_21018,N_20776);
nand U27668 (N_27668,N_20883,N_21501);
xnor U27669 (N_27669,N_22305,N_22852);
and U27670 (N_27670,N_21555,N_23662);
nand U27671 (N_27671,N_21086,N_24990);
nor U27672 (N_27672,N_24829,N_20714);
nor U27673 (N_27673,N_23631,N_22604);
and U27674 (N_27674,N_22231,N_24587);
and U27675 (N_27675,N_20489,N_23912);
nand U27676 (N_27676,N_23852,N_21268);
or U27677 (N_27677,N_20826,N_24009);
and U27678 (N_27678,N_22654,N_24332);
and U27679 (N_27679,N_23097,N_22705);
and U27680 (N_27680,N_22353,N_24042);
nand U27681 (N_27681,N_23108,N_23654);
nor U27682 (N_27682,N_23093,N_24383);
xnor U27683 (N_27683,N_23975,N_24313);
and U27684 (N_27684,N_22044,N_20956);
and U27685 (N_27685,N_23131,N_24670);
or U27686 (N_27686,N_21764,N_24965);
nand U27687 (N_27687,N_24464,N_24205);
nor U27688 (N_27688,N_24820,N_22512);
nor U27689 (N_27689,N_24343,N_21080);
or U27690 (N_27690,N_22877,N_21206);
or U27691 (N_27691,N_21105,N_23224);
or U27692 (N_27692,N_22336,N_21216);
or U27693 (N_27693,N_24308,N_21226);
nor U27694 (N_27694,N_23545,N_21021);
xor U27695 (N_27695,N_23661,N_22546);
nand U27696 (N_27696,N_24190,N_23380);
or U27697 (N_27697,N_24120,N_23690);
or U27698 (N_27698,N_21503,N_21499);
nand U27699 (N_27699,N_24485,N_22155);
nand U27700 (N_27700,N_20055,N_24032);
nand U27701 (N_27701,N_23562,N_24208);
nor U27702 (N_27702,N_21756,N_23395);
nand U27703 (N_27703,N_24366,N_21868);
and U27704 (N_27704,N_22388,N_24515);
nand U27705 (N_27705,N_24045,N_20842);
xnor U27706 (N_27706,N_22990,N_24045);
or U27707 (N_27707,N_22163,N_24385);
and U27708 (N_27708,N_23292,N_24591);
nand U27709 (N_27709,N_21115,N_21976);
and U27710 (N_27710,N_20109,N_21880);
and U27711 (N_27711,N_23350,N_22049);
nor U27712 (N_27712,N_23774,N_20184);
and U27713 (N_27713,N_24482,N_21069);
xnor U27714 (N_27714,N_23743,N_24454);
xor U27715 (N_27715,N_21083,N_23633);
and U27716 (N_27716,N_22682,N_23525);
nand U27717 (N_27717,N_24289,N_20506);
nor U27718 (N_27718,N_24258,N_21828);
nand U27719 (N_27719,N_21804,N_24422);
nor U27720 (N_27720,N_20557,N_23071);
or U27721 (N_27721,N_22971,N_23875);
and U27722 (N_27722,N_22158,N_21937);
or U27723 (N_27723,N_20216,N_23802);
xor U27724 (N_27724,N_21403,N_21004);
xor U27725 (N_27725,N_21085,N_21966);
nand U27726 (N_27726,N_23055,N_22009);
and U27727 (N_27727,N_22349,N_22767);
nor U27728 (N_27728,N_24936,N_21583);
xor U27729 (N_27729,N_20013,N_21958);
nor U27730 (N_27730,N_24907,N_21981);
nand U27731 (N_27731,N_22221,N_24501);
and U27732 (N_27732,N_21451,N_23442);
nor U27733 (N_27733,N_22653,N_21579);
nor U27734 (N_27734,N_24236,N_22381);
nor U27735 (N_27735,N_24199,N_20879);
and U27736 (N_27736,N_21638,N_23933);
or U27737 (N_27737,N_20294,N_23488);
nand U27738 (N_27738,N_24949,N_24999);
xor U27739 (N_27739,N_20632,N_23565);
and U27740 (N_27740,N_24898,N_20584);
nand U27741 (N_27741,N_22588,N_23599);
and U27742 (N_27742,N_21710,N_22803);
and U27743 (N_27743,N_20974,N_24711);
or U27744 (N_27744,N_22117,N_21705);
and U27745 (N_27745,N_20553,N_21607);
and U27746 (N_27746,N_21069,N_24414);
and U27747 (N_27747,N_24241,N_20401);
nor U27748 (N_27748,N_24433,N_21470);
xor U27749 (N_27749,N_24375,N_22174);
nand U27750 (N_27750,N_24304,N_23750);
nand U27751 (N_27751,N_20394,N_20194);
nand U27752 (N_27752,N_23656,N_23863);
and U27753 (N_27753,N_23544,N_23742);
nor U27754 (N_27754,N_22253,N_20484);
and U27755 (N_27755,N_24153,N_20729);
nor U27756 (N_27756,N_20438,N_20147);
xor U27757 (N_27757,N_20543,N_22254);
or U27758 (N_27758,N_20793,N_24782);
and U27759 (N_27759,N_23784,N_22466);
and U27760 (N_27760,N_22281,N_21503);
xor U27761 (N_27761,N_20491,N_24899);
and U27762 (N_27762,N_22901,N_22262);
or U27763 (N_27763,N_23987,N_23214);
and U27764 (N_27764,N_21431,N_21493);
or U27765 (N_27765,N_20953,N_20793);
nand U27766 (N_27766,N_20911,N_21626);
xnor U27767 (N_27767,N_20098,N_24146);
nor U27768 (N_27768,N_21364,N_22172);
nor U27769 (N_27769,N_21462,N_23848);
xnor U27770 (N_27770,N_23581,N_22314);
nand U27771 (N_27771,N_24372,N_22282);
or U27772 (N_27772,N_22785,N_20735);
and U27773 (N_27773,N_21089,N_22289);
or U27774 (N_27774,N_22483,N_20120);
or U27775 (N_27775,N_23719,N_24905);
and U27776 (N_27776,N_24179,N_23928);
or U27777 (N_27777,N_21748,N_24451);
nand U27778 (N_27778,N_23959,N_24707);
and U27779 (N_27779,N_23952,N_24871);
nor U27780 (N_27780,N_20164,N_24894);
nand U27781 (N_27781,N_23632,N_24384);
or U27782 (N_27782,N_22142,N_24753);
nor U27783 (N_27783,N_24938,N_22446);
nor U27784 (N_27784,N_23937,N_22513);
nor U27785 (N_27785,N_23525,N_23608);
and U27786 (N_27786,N_22490,N_21512);
and U27787 (N_27787,N_23398,N_20540);
or U27788 (N_27788,N_20116,N_20589);
and U27789 (N_27789,N_23098,N_20590);
and U27790 (N_27790,N_21230,N_22056);
xor U27791 (N_27791,N_21263,N_21290);
nor U27792 (N_27792,N_22000,N_23212);
nand U27793 (N_27793,N_20714,N_24823);
nand U27794 (N_27794,N_24170,N_22628);
and U27795 (N_27795,N_23914,N_22538);
or U27796 (N_27796,N_21231,N_20912);
xor U27797 (N_27797,N_21847,N_24236);
or U27798 (N_27798,N_23538,N_22066);
and U27799 (N_27799,N_23017,N_20520);
and U27800 (N_27800,N_21836,N_21819);
and U27801 (N_27801,N_21703,N_24574);
or U27802 (N_27802,N_20607,N_23303);
or U27803 (N_27803,N_20777,N_21263);
nor U27804 (N_27804,N_23652,N_24558);
or U27805 (N_27805,N_24040,N_21868);
or U27806 (N_27806,N_24240,N_24194);
and U27807 (N_27807,N_20623,N_24663);
and U27808 (N_27808,N_24438,N_23438);
nand U27809 (N_27809,N_21312,N_20471);
xor U27810 (N_27810,N_24248,N_23274);
xor U27811 (N_27811,N_20735,N_22492);
nor U27812 (N_27812,N_20153,N_22706);
and U27813 (N_27813,N_22969,N_20294);
nor U27814 (N_27814,N_23684,N_22457);
or U27815 (N_27815,N_23662,N_22051);
nor U27816 (N_27816,N_22802,N_22135);
nand U27817 (N_27817,N_24537,N_22248);
nor U27818 (N_27818,N_21222,N_22001);
xor U27819 (N_27819,N_23778,N_20885);
nand U27820 (N_27820,N_20062,N_24705);
or U27821 (N_27821,N_22978,N_20456);
nand U27822 (N_27822,N_21846,N_24434);
nor U27823 (N_27823,N_24137,N_24926);
xnor U27824 (N_27824,N_21684,N_24336);
nand U27825 (N_27825,N_20322,N_23263);
nor U27826 (N_27826,N_22704,N_22528);
nand U27827 (N_27827,N_23296,N_22222);
or U27828 (N_27828,N_21910,N_22376);
nand U27829 (N_27829,N_23371,N_23549);
nor U27830 (N_27830,N_23523,N_20384);
or U27831 (N_27831,N_20868,N_24540);
nor U27832 (N_27832,N_21191,N_23945);
nor U27833 (N_27833,N_21490,N_22078);
nor U27834 (N_27834,N_22949,N_20222);
xnor U27835 (N_27835,N_22048,N_22056);
or U27836 (N_27836,N_23124,N_20948);
and U27837 (N_27837,N_20630,N_21544);
nor U27838 (N_27838,N_24958,N_24065);
and U27839 (N_27839,N_21446,N_24493);
and U27840 (N_27840,N_22458,N_20887);
nor U27841 (N_27841,N_21096,N_20536);
and U27842 (N_27842,N_23070,N_24594);
nor U27843 (N_27843,N_22130,N_21477);
or U27844 (N_27844,N_20141,N_21251);
and U27845 (N_27845,N_21696,N_23259);
nor U27846 (N_27846,N_20727,N_20248);
and U27847 (N_27847,N_22076,N_20632);
nor U27848 (N_27848,N_22679,N_22554);
xor U27849 (N_27849,N_23667,N_21544);
nand U27850 (N_27850,N_24360,N_21019);
or U27851 (N_27851,N_23023,N_24111);
nand U27852 (N_27852,N_22853,N_20459);
or U27853 (N_27853,N_20740,N_22574);
nor U27854 (N_27854,N_23731,N_22125);
nor U27855 (N_27855,N_22872,N_21788);
xnor U27856 (N_27856,N_22383,N_20780);
nor U27857 (N_27857,N_23855,N_23619);
xnor U27858 (N_27858,N_21022,N_23410);
xnor U27859 (N_27859,N_21644,N_22979);
nand U27860 (N_27860,N_21539,N_20148);
and U27861 (N_27861,N_20754,N_24880);
nand U27862 (N_27862,N_24335,N_24054);
and U27863 (N_27863,N_23495,N_24457);
nand U27864 (N_27864,N_22180,N_21600);
and U27865 (N_27865,N_21774,N_24341);
and U27866 (N_27866,N_22733,N_21562);
and U27867 (N_27867,N_22062,N_23071);
or U27868 (N_27868,N_21584,N_24185);
nor U27869 (N_27869,N_21600,N_24017);
or U27870 (N_27870,N_23148,N_20709);
and U27871 (N_27871,N_21854,N_22472);
xor U27872 (N_27872,N_24017,N_20076);
nand U27873 (N_27873,N_20650,N_24387);
xnor U27874 (N_27874,N_23513,N_20375);
and U27875 (N_27875,N_24265,N_20001);
nor U27876 (N_27876,N_20191,N_23799);
nand U27877 (N_27877,N_20600,N_21225);
nor U27878 (N_27878,N_22504,N_20034);
and U27879 (N_27879,N_21332,N_24498);
or U27880 (N_27880,N_24349,N_22870);
or U27881 (N_27881,N_21795,N_23081);
and U27882 (N_27882,N_22788,N_21621);
xor U27883 (N_27883,N_24998,N_21602);
xnor U27884 (N_27884,N_21471,N_21399);
and U27885 (N_27885,N_23067,N_21962);
or U27886 (N_27886,N_21073,N_20813);
nand U27887 (N_27887,N_20035,N_23282);
xor U27888 (N_27888,N_21793,N_20152);
nor U27889 (N_27889,N_21661,N_21675);
xor U27890 (N_27890,N_24863,N_21488);
nand U27891 (N_27891,N_23068,N_21736);
nor U27892 (N_27892,N_24436,N_20447);
xor U27893 (N_27893,N_22245,N_22344);
nand U27894 (N_27894,N_21291,N_23524);
xnor U27895 (N_27895,N_22126,N_21709);
or U27896 (N_27896,N_23540,N_23399);
and U27897 (N_27897,N_23181,N_20147);
nor U27898 (N_27898,N_24082,N_20994);
or U27899 (N_27899,N_20081,N_21548);
xnor U27900 (N_27900,N_21553,N_21068);
or U27901 (N_27901,N_24125,N_21666);
xnor U27902 (N_27902,N_22022,N_21920);
nand U27903 (N_27903,N_22021,N_20705);
xnor U27904 (N_27904,N_20927,N_23085);
xor U27905 (N_27905,N_22994,N_22716);
or U27906 (N_27906,N_21192,N_21958);
xor U27907 (N_27907,N_23643,N_23176);
xnor U27908 (N_27908,N_24678,N_24176);
nand U27909 (N_27909,N_22690,N_23987);
xnor U27910 (N_27910,N_21984,N_23747);
nor U27911 (N_27911,N_21366,N_21631);
or U27912 (N_27912,N_20180,N_22965);
and U27913 (N_27913,N_21667,N_23452);
or U27914 (N_27914,N_21753,N_20548);
nand U27915 (N_27915,N_21318,N_23287);
and U27916 (N_27916,N_24947,N_21710);
or U27917 (N_27917,N_20646,N_23486);
xor U27918 (N_27918,N_23521,N_20802);
and U27919 (N_27919,N_24289,N_21588);
nor U27920 (N_27920,N_20583,N_23288);
nand U27921 (N_27921,N_22973,N_20057);
xnor U27922 (N_27922,N_20285,N_24030);
nand U27923 (N_27923,N_22578,N_24915);
nor U27924 (N_27924,N_20130,N_20400);
xnor U27925 (N_27925,N_23304,N_22872);
nor U27926 (N_27926,N_24683,N_24416);
nand U27927 (N_27927,N_20627,N_23654);
or U27928 (N_27928,N_23989,N_22206);
xor U27929 (N_27929,N_21080,N_21746);
xnor U27930 (N_27930,N_20989,N_21640);
and U27931 (N_27931,N_20120,N_21757);
xor U27932 (N_27932,N_20123,N_24044);
and U27933 (N_27933,N_24665,N_21507);
nor U27934 (N_27934,N_21722,N_24353);
and U27935 (N_27935,N_24348,N_21332);
xnor U27936 (N_27936,N_22845,N_21975);
nand U27937 (N_27937,N_20553,N_22234);
or U27938 (N_27938,N_23640,N_22975);
and U27939 (N_27939,N_21322,N_24945);
or U27940 (N_27940,N_20285,N_22423);
nand U27941 (N_27941,N_20399,N_22751);
xor U27942 (N_27942,N_21867,N_22043);
nand U27943 (N_27943,N_24306,N_24412);
xor U27944 (N_27944,N_20202,N_22749);
or U27945 (N_27945,N_21749,N_23185);
or U27946 (N_27946,N_22962,N_22746);
and U27947 (N_27947,N_24833,N_22977);
xnor U27948 (N_27948,N_23520,N_21075);
or U27949 (N_27949,N_22307,N_22053);
nand U27950 (N_27950,N_22962,N_23223);
and U27951 (N_27951,N_21426,N_20724);
nand U27952 (N_27952,N_24093,N_24704);
or U27953 (N_27953,N_20896,N_22845);
nor U27954 (N_27954,N_22593,N_22130);
nor U27955 (N_27955,N_22275,N_20243);
or U27956 (N_27956,N_20408,N_24407);
and U27957 (N_27957,N_24952,N_22512);
or U27958 (N_27958,N_22663,N_21664);
and U27959 (N_27959,N_20185,N_21975);
xor U27960 (N_27960,N_22406,N_21910);
xor U27961 (N_27961,N_22344,N_20398);
nand U27962 (N_27962,N_20500,N_22346);
xnor U27963 (N_27963,N_21832,N_21238);
xor U27964 (N_27964,N_22893,N_20407);
or U27965 (N_27965,N_21536,N_21308);
and U27966 (N_27966,N_20824,N_21554);
or U27967 (N_27967,N_20040,N_21312);
xnor U27968 (N_27968,N_22085,N_24031);
xnor U27969 (N_27969,N_20667,N_23400);
nand U27970 (N_27970,N_22058,N_23662);
nor U27971 (N_27971,N_20739,N_24360);
xor U27972 (N_27972,N_24360,N_22372);
or U27973 (N_27973,N_22999,N_23703);
and U27974 (N_27974,N_22378,N_24202);
nor U27975 (N_27975,N_24802,N_20420);
or U27976 (N_27976,N_20605,N_23752);
and U27977 (N_27977,N_20499,N_21017);
or U27978 (N_27978,N_21190,N_24236);
nor U27979 (N_27979,N_23853,N_24122);
nor U27980 (N_27980,N_23605,N_24284);
and U27981 (N_27981,N_20060,N_23451);
nor U27982 (N_27982,N_21199,N_20545);
and U27983 (N_27983,N_22351,N_24512);
nand U27984 (N_27984,N_24247,N_23463);
nand U27985 (N_27985,N_23300,N_22436);
and U27986 (N_27986,N_23891,N_23934);
nor U27987 (N_27987,N_21586,N_23193);
nand U27988 (N_27988,N_24491,N_20029);
nand U27989 (N_27989,N_22216,N_23316);
and U27990 (N_27990,N_22210,N_21399);
nor U27991 (N_27991,N_21895,N_24278);
nor U27992 (N_27992,N_24516,N_23907);
and U27993 (N_27993,N_20644,N_24770);
or U27994 (N_27994,N_23093,N_22873);
xor U27995 (N_27995,N_23880,N_24564);
nand U27996 (N_27996,N_24875,N_24472);
xnor U27997 (N_27997,N_21775,N_21842);
nand U27998 (N_27998,N_22901,N_23256);
nand U27999 (N_27999,N_22979,N_22140);
and U28000 (N_28000,N_22210,N_24926);
xor U28001 (N_28001,N_23706,N_23434);
nor U28002 (N_28002,N_22475,N_23695);
nand U28003 (N_28003,N_23938,N_24691);
nor U28004 (N_28004,N_20706,N_23879);
xnor U28005 (N_28005,N_23438,N_22439);
nor U28006 (N_28006,N_22539,N_21059);
or U28007 (N_28007,N_20424,N_23152);
nor U28008 (N_28008,N_22966,N_23800);
or U28009 (N_28009,N_24339,N_23830);
xnor U28010 (N_28010,N_23148,N_23137);
nand U28011 (N_28011,N_24266,N_23925);
and U28012 (N_28012,N_23074,N_22194);
xor U28013 (N_28013,N_24231,N_22655);
or U28014 (N_28014,N_23924,N_24676);
nand U28015 (N_28015,N_20406,N_21326);
or U28016 (N_28016,N_22905,N_22733);
or U28017 (N_28017,N_23416,N_22125);
xor U28018 (N_28018,N_23166,N_24796);
xnor U28019 (N_28019,N_22117,N_22197);
and U28020 (N_28020,N_22865,N_20760);
and U28021 (N_28021,N_23311,N_22630);
nand U28022 (N_28022,N_22925,N_24604);
nand U28023 (N_28023,N_23552,N_23130);
nand U28024 (N_28024,N_23123,N_24950);
or U28025 (N_28025,N_23510,N_24796);
nand U28026 (N_28026,N_23641,N_23050);
and U28027 (N_28027,N_21952,N_24774);
or U28028 (N_28028,N_23138,N_21211);
and U28029 (N_28029,N_20404,N_23212);
nor U28030 (N_28030,N_20339,N_20825);
nand U28031 (N_28031,N_24407,N_24082);
and U28032 (N_28032,N_23658,N_24616);
nand U28033 (N_28033,N_24105,N_22723);
xnor U28034 (N_28034,N_23633,N_20264);
nor U28035 (N_28035,N_21517,N_23274);
xor U28036 (N_28036,N_21480,N_21199);
nor U28037 (N_28037,N_23489,N_23890);
or U28038 (N_28038,N_24873,N_24571);
nor U28039 (N_28039,N_23467,N_20560);
xor U28040 (N_28040,N_20155,N_20496);
xnor U28041 (N_28041,N_21111,N_24330);
nor U28042 (N_28042,N_20160,N_24622);
xor U28043 (N_28043,N_20173,N_24032);
nand U28044 (N_28044,N_24556,N_20282);
or U28045 (N_28045,N_23791,N_20382);
and U28046 (N_28046,N_23335,N_23425);
nand U28047 (N_28047,N_22660,N_23168);
or U28048 (N_28048,N_20588,N_24621);
or U28049 (N_28049,N_22513,N_24020);
or U28050 (N_28050,N_22102,N_22044);
nand U28051 (N_28051,N_22598,N_22940);
or U28052 (N_28052,N_23855,N_22390);
nand U28053 (N_28053,N_21558,N_24889);
and U28054 (N_28054,N_22745,N_23987);
nand U28055 (N_28055,N_23257,N_23387);
or U28056 (N_28056,N_20054,N_23429);
and U28057 (N_28057,N_23744,N_22424);
xnor U28058 (N_28058,N_23215,N_20604);
nor U28059 (N_28059,N_24748,N_23012);
nand U28060 (N_28060,N_23856,N_23744);
nor U28061 (N_28061,N_23927,N_23098);
nor U28062 (N_28062,N_24577,N_24906);
nand U28063 (N_28063,N_23565,N_21985);
nor U28064 (N_28064,N_21135,N_23361);
xnor U28065 (N_28065,N_22064,N_21541);
nor U28066 (N_28066,N_23059,N_22614);
and U28067 (N_28067,N_20535,N_21249);
nor U28068 (N_28068,N_23981,N_24358);
or U28069 (N_28069,N_20053,N_24542);
nand U28070 (N_28070,N_23536,N_24187);
nor U28071 (N_28071,N_23808,N_21284);
nor U28072 (N_28072,N_23573,N_24375);
xor U28073 (N_28073,N_23022,N_22607);
nor U28074 (N_28074,N_22502,N_23905);
nand U28075 (N_28075,N_20249,N_24003);
and U28076 (N_28076,N_21416,N_24726);
nand U28077 (N_28077,N_21397,N_21041);
nand U28078 (N_28078,N_23369,N_21898);
nand U28079 (N_28079,N_21290,N_24288);
nand U28080 (N_28080,N_23241,N_23792);
and U28081 (N_28081,N_20338,N_20986);
xor U28082 (N_28082,N_20492,N_21457);
or U28083 (N_28083,N_20109,N_23359);
nand U28084 (N_28084,N_22888,N_23836);
nand U28085 (N_28085,N_22593,N_21820);
nor U28086 (N_28086,N_22842,N_20856);
or U28087 (N_28087,N_22851,N_22880);
and U28088 (N_28088,N_23974,N_21845);
or U28089 (N_28089,N_21937,N_22013);
and U28090 (N_28090,N_20019,N_23503);
nor U28091 (N_28091,N_21380,N_22091);
and U28092 (N_28092,N_21282,N_23827);
and U28093 (N_28093,N_23114,N_21776);
xnor U28094 (N_28094,N_21510,N_23840);
or U28095 (N_28095,N_23440,N_21802);
or U28096 (N_28096,N_24798,N_24954);
and U28097 (N_28097,N_24061,N_20409);
xnor U28098 (N_28098,N_20822,N_24683);
nor U28099 (N_28099,N_23912,N_22385);
xnor U28100 (N_28100,N_24792,N_20670);
and U28101 (N_28101,N_20422,N_22544);
and U28102 (N_28102,N_20150,N_23188);
nor U28103 (N_28103,N_20994,N_21996);
nand U28104 (N_28104,N_22490,N_23160);
nand U28105 (N_28105,N_20286,N_23845);
and U28106 (N_28106,N_22908,N_20696);
and U28107 (N_28107,N_23070,N_21158);
and U28108 (N_28108,N_24648,N_24026);
or U28109 (N_28109,N_20684,N_23152);
and U28110 (N_28110,N_21676,N_22895);
and U28111 (N_28111,N_22837,N_24976);
and U28112 (N_28112,N_23374,N_24142);
and U28113 (N_28113,N_23720,N_22746);
and U28114 (N_28114,N_22127,N_20596);
and U28115 (N_28115,N_20555,N_20482);
nand U28116 (N_28116,N_23785,N_20935);
nor U28117 (N_28117,N_20879,N_22540);
nand U28118 (N_28118,N_22334,N_23914);
nand U28119 (N_28119,N_24921,N_24013);
xnor U28120 (N_28120,N_22655,N_21855);
nor U28121 (N_28121,N_21982,N_23533);
nand U28122 (N_28122,N_21249,N_22559);
and U28123 (N_28123,N_22851,N_20168);
and U28124 (N_28124,N_20088,N_21826);
or U28125 (N_28125,N_24138,N_20524);
and U28126 (N_28126,N_23356,N_20837);
nand U28127 (N_28127,N_24470,N_20624);
and U28128 (N_28128,N_20701,N_22966);
nor U28129 (N_28129,N_24673,N_20946);
nor U28130 (N_28130,N_24090,N_24223);
and U28131 (N_28131,N_23016,N_21892);
and U28132 (N_28132,N_21574,N_20106);
or U28133 (N_28133,N_24885,N_22668);
nor U28134 (N_28134,N_23669,N_23200);
nand U28135 (N_28135,N_23707,N_24845);
or U28136 (N_28136,N_22355,N_22348);
xnor U28137 (N_28137,N_23544,N_24910);
nand U28138 (N_28138,N_22988,N_24283);
xor U28139 (N_28139,N_22660,N_21531);
nor U28140 (N_28140,N_24838,N_20895);
nor U28141 (N_28141,N_24882,N_24017);
xnor U28142 (N_28142,N_24604,N_21306);
xnor U28143 (N_28143,N_21842,N_20831);
and U28144 (N_28144,N_24174,N_22190);
nor U28145 (N_28145,N_20515,N_24397);
nand U28146 (N_28146,N_21389,N_21781);
nand U28147 (N_28147,N_21256,N_22719);
xor U28148 (N_28148,N_20924,N_23692);
and U28149 (N_28149,N_22610,N_20303);
or U28150 (N_28150,N_20592,N_21200);
xnor U28151 (N_28151,N_22574,N_24792);
nand U28152 (N_28152,N_20564,N_20573);
and U28153 (N_28153,N_23649,N_22751);
nor U28154 (N_28154,N_20184,N_20265);
nand U28155 (N_28155,N_22174,N_20799);
nor U28156 (N_28156,N_20468,N_24493);
xor U28157 (N_28157,N_24563,N_24909);
nand U28158 (N_28158,N_22152,N_24090);
and U28159 (N_28159,N_23126,N_23369);
xor U28160 (N_28160,N_22460,N_23907);
or U28161 (N_28161,N_22685,N_20789);
xnor U28162 (N_28162,N_24746,N_23321);
or U28163 (N_28163,N_21209,N_23188);
or U28164 (N_28164,N_21164,N_24781);
and U28165 (N_28165,N_22268,N_20520);
and U28166 (N_28166,N_23802,N_21101);
nand U28167 (N_28167,N_20258,N_20422);
nand U28168 (N_28168,N_21296,N_20888);
nor U28169 (N_28169,N_24901,N_24479);
nand U28170 (N_28170,N_23158,N_22130);
or U28171 (N_28171,N_20120,N_24366);
xnor U28172 (N_28172,N_23704,N_20686);
and U28173 (N_28173,N_20314,N_20875);
and U28174 (N_28174,N_24251,N_21831);
nand U28175 (N_28175,N_21070,N_24125);
xor U28176 (N_28176,N_20512,N_20668);
or U28177 (N_28177,N_20621,N_24392);
or U28178 (N_28178,N_21166,N_22877);
nor U28179 (N_28179,N_20145,N_24607);
nand U28180 (N_28180,N_23548,N_21807);
nand U28181 (N_28181,N_23017,N_23868);
and U28182 (N_28182,N_21929,N_21293);
nor U28183 (N_28183,N_20798,N_23581);
xor U28184 (N_28184,N_21006,N_23605);
xor U28185 (N_28185,N_21736,N_22728);
and U28186 (N_28186,N_24374,N_22049);
xor U28187 (N_28187,N_24344,N_22206);
nor U28188 (N_28188,N_20089,N_21145);
or U28189 (N_28189,N_20504,N_21964);
nor U28190 (N_28190,N_22560,N_23609);
nor U28191 (N_28191,N_22247,N_22078);
nor U28192 (N_28192,N_24024,N_22985);
nand U28193 (N_28193,N_22997,N_20060);
nand U28194 (N_28194,N_21897,N_21019);
xnor U28195 (N_28195,N_23801,N_21875);
nand U28196 (N_28196,N_24146,N_21679);
and U28197 (N_28197,N_20073,N_22361);
or U28198 (N_28198,N_24607,N_21045);
nand U28199 (N_28199,N_24103,N_20137);
and U28200 (N_28200,N_24020,N_20908);
and U28201 (N_28201,N_20111,N_24139);
or U28202 (N_28202,N_23166,N_20556);
xnor U28203 (N_28203,N_24430,N_22547);
nand U28204 (N_28204,N_24523,N_22464);
nor U28205 (N_28205,N_21093,N_24810);
or U28206 (N_28206,N_22997,N_21283);
or U28207 (N_28207,N_23793,N_24528);
nand U28208 (N_28208,N_20847,N_20658);
nand U28209 (N_28209,N_21393,N_22867);
xnor U28210 (N_28210,N_21673,N_21759);
and U28211 (N_28211,N_20472,N_22980);
nor U28212 (N_28212,N_20792,N_23652);
or U28213 (N_28213,N_20152,N_21381);
nor U28214 (N_28214,N_23349,N_20557);
or U28215 (N_28215,N_22641,N_21432);
nor U28216 (N_28216,N_23350,N_23584);
nand U28217 (N_28217,N_22146,N_24611);
nand U28218 (N_28218,N_20375,N_24375);
and U28219 (N_28219,N_20968,N_20602);
or U28220 (N_28220,N_24443,N_21835);
or U28221 (N_28221,N_21816,N_24092);
nand U28222 (N_28222,N_23737,N_20524);
nand U28223 (N_28223,N_23553,N_23985);
xor U28224 (N_28224,N_24244,N_21316);
xor U28225 (N_28225,N_22915,N_21753);
nor U28226 (N_28226,N_23672,N_22259);
xnor U28227 (N_28227,N_23919,N_24194);
and U28228 (N_28228,N_21177,N_21979);
or U28229 (N_28229,N_22776,N_23455);
xor U28230 (N_28230,N_23931,N_24388);
nor U28231 (N_28231,N_23652,N_21624);
nor U28232 (N_28232,N_24949,N_24150);
nand U28233 (N_28233,N_20708,N_24969);
nand U28234 (N_28234,N_23065,N_24369);
nor U28235 (N_28235,N_22741,N_23570);
and U28236 (N_28236,N_20393,N_23474);
xor U28237 (N_28237,N_21118,N_24391);
or U28238 (N_28238,N_24136,N_21046);
or U28239 (N_28239,N_23188,N_24183);
or U28240 (N_28240,N_23326,N_21366);
nand U28241 (N_28241,N_22431,N_22504);
or U28242 (N_28242,N_24964,N_23586);
and U28243 (N_28243,N_23524,N_22517);
nand U28244 (N_28244,N_23219,N_20015);
or U28245 (N_28245,N_20172,N_20964);
or U28246 (N_28246,N_23591,N_23669);
and U28247 (N_28247,N_23118,N_21843);
nor U28248 (N_28248,N_22835,N_22406);
xor U28249 (N_28249,N_21596,N_24824);
or U28250 (N_28250,N_21842,N_20094);
or U28251 (N_28251,N_22905,N_22726);
and U28252 (N_28252,N_22025,N_24514);
nor U28253 (N_28253,N_23306,N_21107);
and U28254 (N_28254,N_24664,N_23656);
and U28255 (N_28255,N_21020,N_20471);
nor U28256 (N_28256,N_21973,N_22569);
or U28257 (N_28257,N_21075,N_24762);
xnor U28258 (N_28258,N_21444,N_22620);
xnor U28259 (N_28259,N_21910,N_24797);
nand U28260 (N_28260,N_21489,N_21252);
and U28261 (N_28261,N_21587,N_22510);
nand U28262 (N_28262,N_23426,N_20816);
or U28263 (N_28263,N_23023,N_23252);
and U28264 (N_28264,N_22676,N_22602);
and U28265 (N_28265,N_24383,N_24236);
xnor U28266 (N_28266,N_23443,N_23817);
nor U28267 (N_28267,N_21642,N_21648);
and U28268 (N_28268,N_20611,N_24174);
and U28269 (N_28269,N_20105,N_24974);
or U28270 (N_28270,N_24698,N_22468);
or U28271 (N_28271,N_21999,N_21694);
xor U28272 (N_28272,N_20992,N_22567);
nor U28273 (N_28273,N_21642,N_22883);
nor U28274 (N_28274,N_23436,N_21708);
or U28275 (N_28275,N_20625,N_23617);
nor U28276 (N_28276,N_20940,N_20192);
nor U28277 (N_28277,N_20414,N_20617);
xnor U28278 (N_28278,N_24480,N_20757);
nor U28279 (N_28279,N_21979,N_21174);
nand U28280 (N_28280,N_22976,N_20742);
nand U28281 (N_28281,N_24857,N_23992);
xor U28282 (N_28282,N_24565,N_21452);
and U28283 (N_28283,N_21657,N_24253);
and U28284 (N_28284,N_21599,N_23010);
xnor U28285 (N_28285,N_21416,N_24888);
or U28286 (N_28286,N_21723,N_21794);
nor U28287 (N_28287,N_20015,N_21682);
and U28288 (N_28288,N_22041,N_21394);
or U28289 (N_28289,N_21589,N_23577);
and U28290 (N_28290,N_20355,N_20017);
and U28291 (N_28291,N_21137,N_22653);
nand U28292 (N_28292,N_20298,N_21040);
nor U28293 (N_28293,N_21648,N_21423);
xnor U28294 (N_28294,N_20899,N_20784);
or U28295 (N_28295,N_24722,N_24770);
xor U28296 (N_28296,N_23789,N_21797);
nor U28297 (N_28297,N_23497,N_20859);
nand U28298 (N_28298,N_24519,N_20416);
xnor U28299 (N_28299,N_23268,N_24133);
or U28300 (N_28300,N_22917,N_21508);
xnor U28301 (N_28301,N_20313,N_23708);
nor U28302 (N_28302,N_22484,N_21215);
xor U28303 (N_28303,N_22769,N_22401);
and U28304 (N_28304,N_24677,N_23818);
xnor U28305 (N_28305,N_24298,N_20968);
nor U28306 (N_28306,N_20371,N_22123);
nand U28307 (N_28307,N_22413,N_20087);
xnor U28308 (N_28308,N_20934,N_20623);
xnor U28309 (N_28309,N_22237,N_21478);
xor U28310 (N_28310,N_24892,N_22203);
nand U28311 (N_28311,N_23090,N_21515);
xnor U28312 (N_28312,N_21327,N_22847);
nand U28313 (N_28313,N_23091,N_21007);
xor U28314 (N_28314,N_23638,N_20678);
and U28315 (N_28315,N_23683,N_20227);
and U28316 (N_28316,N_24995,N_20466);
or U28317 (N_28317,N_24412,N_22041);
nor U28318 (N_28318,N_21252,N_22066);
xnor U28319 (N_28319,N_22259,N_24996);
nor U28320 (N_28320,N_21003,N_22318);
xnor U28321 (N_28321,N_22318,N_23333);
nand U28322 (N_28322,N_24327,N_20210);
nor U28323 (N_28323,N_23952,N_23544);
nor U28324 (N_28324,N_20155,N_21288);
xnor U28325 (N_28325,N_23794,N_24674);
nand U28326 (N_28326,N_21197,N_20650);
xnor U28327 (N_28327,N_20616,N_24303);
nor U28328 (N_28328,N_22955,N_24082);
nor U28329 (N_28329,N_22080,N_20704);
nand U28330 (N_28330,N_21196,N_24661);
nand U28331 (N_28331,N_21068,N_21777);
nand U28332 (N_28332,N_24086,N_22075);
nand U28333 (N_28333,N_21142,N_20449);
xnor U28334 (N_28334,N_20993,N_21874);
and U28335 (N_28335,N_22144,N_24681);
nand U28336 (N_28336,N_20116,N_22895);
or U28337 (N_28337,N_23060,N_21151);
xnor U28338 (N_28338,N_21582,N_23940);
and U28339 (N_28339,N_22111,N_21508);
xnor U28340 (N_28340,N_24313,N_22057);
nor U28341 (N_28341,N_24430,N_24061);
or U28342 (N_28342,N_20545,N_23127);
and U28343 (N_28343,N_21751,N_21403);
and U28344 (N_28344,N_22664,N_21591);
nor U28345 (N_28345,N_22947,N_22874);
nand U28346 (N_28346,N_23804,N_24395);
nand U28347 (N_28347,N_24867,N_20036);
nand U28348 (N_28348,N_21789,N_24940);
nor U28349 (N_28349,N_20319,N_22077);
nand U28350 (N_28350,N_23660,N_23133);
or U28351 (N_28351,N_24590,N_24761);
nand U28352 (N_28352,N_23110,N_21239);
and U28353 (N_28353,N_24158,N_21125);
and U28354 (N_28354,N_23250,N_22355);
nor U28355 (N_28355,N_24403,N_22560);
nor U28356 (N_28356,N_24527,N_21251);
xor U28357 (N_28357,N_21711,N_20665);
xnor U28358 (N_28358,N_20007,N_20713);
nand U28359 (N_28359,N_22276,N_24231);
and U28360 (N_28360,N_24830,N_20683);
and U28361 (N_28361,N_22105,N_20555);
or U28362 (N_28362,N_21281,N_24243);
and U28363 (N_28363,N_20781,N_22859);
and U28364 (N_28364,N_23878,N_20844);
nand U28365 (N_28365,N_22082,N_21627);
xnor U28366 (N_28366,N_24458,N_21983);
and U28367 (N_28367,N_21456,N_24068);
and U28368 (N_28368,N_21996,N_23343);
nor U28369 (N_28369,N_20635,N_23862);
or U28370 (N_28370,N_21321,N_23300);
and U28371 (N_28371,N_22354,N_23496);
nand U28372 (N_28372,N_24464,N_20260);
xor U28373 (N_28373,N_24816,N_21706);
and U28374 (N_28374,N_20773,N_21903);
xor U28375 (N_28375,N_21324,N_24383);
nor U28376 (N_28376,N_20106,N_22544);
and U28377 (N_28377,N_24554,N_23020);
nand U28378 (N_28378,N_21214,N_22237);
xnor U28379 (N_28379,N_22370,N_23514);
and U28380 (N_28380,N_24355,N_24885);
or U28381 (N_28381,N_24218,N_20737);
nand U28382 (N_28382,N_22346,N_20456);
nor U28383 (N_28383,N_21652,N_23571);
nand U28384 (N_28384,N_23292,N_23315);
and U28385 (N_28385,N_24488,N_23012);
or U28386 (N_28386,N_21192,N_20121);
and U28387 (N_28387,N_23991,N_20442);
xnor U28388 (N_28388,N_24948,N_21580);
and U28389 (N_28389,N_23933,N_23708);
nor U28390 (N_28390,N_20172,N_24849);
or U28391 (N_28391,N_20730,N_22031);
or U28392 (N_28392,N_21778,N_22862);
nand U28393 (N_28393,N_22077,N_20956);
nand U28394 (N_28394,N_24408,N_21115);
nand U28395 (N_28395,N_21045,N_24840);
nor U28396 (N_28396,N_21923,N_20987);
nor U28397 (N_28397,N_24420,N_23768);
xnor U28398 (N_28398,N_22413,N_23284);
xnor U28399 (N_28399,N_20646,N_20371);
nand U28400 (N_28400,N_21042,N_23159);
nand U28401 (N_28401,N_21499,N_21982);
nand U28402 (N_28402,N_20678,N_22949);
xnor U28403 (N_28403,N_23310,N_23893);
and U28404 (N_28404,N_21723,N_21699);
or U28405 (N_28405,N_23430,N_24709);
nor U28406 (N_28406,N_22527,N_23054);
xor U28407 (N_28407,N_21135,N_20173);
or U28408 (N_28408,N_24744,N_22205);
nor U28409 (N_28409,N_21515,N_24009);
nand U28410 (N_28410,N_21650,N_21273);
nand U28411 (N_28411,N_23372,N_24386);
xnor U28412 (N_28412,N_21303,N_21975);
or U28413 (N_28413,N_23239,N_20032);
xnor U28414 (N_28414,N_22404,N_22003);
nor U28415 (N_28415,N_24961,N_23831);
or U28416 (N_28416,N_21160,N_20357);
nand U28417 (N_28417,N_21355,N_24366);
and U28418 (N_28418,N_20996,N_23661);
nor U28419 (N_28419,N_22428,N_24379);
or U28420 (N_28420,N_24532,N_20615);
nand U28421 (N_28421,N_24930,N_20354);
nor U28422 (N_28422,N_22868,N_24812);
and U28423 (N_28423,N_20214,N_21846);
xor U28424 (N_28424,N_20924,N_22604);
xor U28425 (N_28425,N_24965,N_22327);
and U28426 (N_28426,N_21069,N_24614);
nand U28427 (N_28427,N_20722,N_21465);
nand U28428 (N_28428,N_23526,N_23205);
or U28429 (N_28429,N_24295,N_20637);
and U28430 (N_28430,N_24965,N_20280);
or U28431 (N_28431,N_23776,N_23165);
xnor U28432 (N_28432,N_22531,N_24298);
nand U28433 (N_28433,N_24815,N_22162);
and U28434 (N_28434,N_22981,N_23299);
xor U28435 (N_28435,N_24332,N_22522);
xor U28436 (N_28436,N_21411,N_21264);
xnor U28437 (N_28437,N_24745,N_24810);
nor U28438 (N_28438,N_21830,N_20319);
or U28439 (N_28439,N_21776,N_22346);
nand U28440 (N_28440,N_24669,N_20892);
xnor U28441 (N_28441,N_20862,N_22931);
and U28442 (N_28442,N_20332,N_24206);
and U28443 (N_28443,N_23344,N_23558);
nor U28444 (N_28444,N_24015,N_23668);
nor U28445 (N_28445,N_22877,N_22241);
xnor U28446 (N_28446,N_23335,N_20438);
or U28447 (N_28447,N_23590,N_20704);
and U28448 (N_28448,N_21038,N_22125);
nand U28449 (N_28449,N_20130,N_23273);
xor U28450 (N_28450,N_20145,N_22315);
nor U28451 (N_28451,N_20565,N_24389);
nor U28452 (N_28452,N_24397,N_23342);
and U28453 (N_28453,N_22069,N_24752);
nand U28454 (N_28454,N_24277,N_20734);
and U28455 (N_28455,N_24750,N_22413);
xnor U28456 (N_28456,N_21083,N_20699);
nor U28457 (N_28457,N_23757,N_23538);
nor U28458 (N_28458,N_23443,N_22411);
or U28459 (N_28459,N_23874,N_23456);
xnor U28460 (N_28460,N_21945,N_20144);
and U28461 (N_28461,N_21521,N_22777);
nor U28462 (N_28462,N_23731,N_20674);
and U28463 (N_28463,N_20696,N_22686);
nand U28464 (N_28464,N_21159,N_21013);
or U28465 (N_28465,N_20447,N_23354);
xnor U28466 (N_28466,N_23843,N_21140);
or U28467 (N_28467,N_23036,N_24018);
xor U28468 (N_28468,N_22397,N_23972);
or U28469 (N_28469,N_22278,N_24083);
or U28470 (N_28470,N_23672,N_20175);
xnor U28471 (N_28471,N_21822,N_23852);
xnor U28472 (N_28472,N_22515,N_20247);
or U28473 (N_28473,N_22871,N_22304);
and U28474 (N_28474,N_23145,N_23725);
nor U28475 (N_28475,N_21958,N_23981);
nor U28476 (N_28476,N_22563,N_23779);
nand U28477 (N_28477,N_21297,N_22140);
and U28478 (N_28478,N_20045,N_23754);
nor U28479 (N_28479,N_24036,N_21134);
xnor U28480 (N_28480,N_22938,N_21880);
nor U28481 (N_28481,N_21052,N_22515);
nor U28482 (N_28482,N_21300,N_21631);
nor U28483 (N_28483,N_23275,N_23475);
and U28484 (N_28484,N_20281,N_22447);
nand U28485 (N_28485,N_21168,N_23088);
nand U28486 (N_28486,N_24062,N_23285);
and U28487 (N_28487,N_22081,N_22961);
xor U28488 (N_28488,N_20832,N_20744);
and U28489 (N_28489,N_22285,N_21382);
and U28490 (N_28490,N_23762,N_22322);
nand U28491 (N_28491,N_21912,N_20603);
xnor U28492 (N_28492,N_23991,N_23203);
xor U28493 (N_28493,N_22440,N_20059);
or U28494 (N_28494,N_21959,N_20704);
xnor U28495 (N_28495,N_21524,N_20745);
nand U28496 (N_28496,N_22988,N_20092);
and U28497 (N_28497,N_23613,N_23932);
and U28498 (N_28498,N_24454,N_21698);
nand U28499 (N_28499,N_22585,N_21429);
or U28500 (N_28500,N_22721,N_21728);
or U28501 (N_28501,N_23647,N_20728);
nor U28502 (N_28502,N_23928,N_22325);
nand U28503 (N_28503,N_23099,N_23549);
nor U28504 (N_28504,N_24472,N_22332);
xnor U28505 (N_28505,N_21170,N_20143);
or U28506 (N_28506,N_22256,N_24025);
nand U28507 (N_28507,N_20826,N_22410);
nor U28508 (N_28508,N_22377,N_23612);
nand U28509 (N_28509,N_20110,N_22987);
xnor U28510 (N_28510,N_21120,N_22124);
nor U28511 (N_28511,N_23153,N_24818);
nor U28512 (N_28512,N_20124,N_23229);
and U28513 (N_28513,N_22174,N_21564);
xnor U28514 (N_28514,N_21453,N_22896);
or U28515 (N_28515,N_22678,N_20216);
or U28516 (N_28516,N_24794,N_21051);
nor U28517 (N_28517,N_21163,N_24704);
or U28518 (N_28518,N_24196,N_24416);
nor U28519 (N_28519,N_22893,N_24483);
nand U28520 (N_28520,N_23450,N_24195);
nor U28521 (N_28521,N_23322,N_20538);
nand U28522 (N_28522,N_20403,N_24278);
nor U28523 (N_28523,N_21301,N_20305);
or U28524 (N_28524,N_21635,N_24745);
nor U28525 (N_28525,N_24531,N_22955);
and U28526 (N_28526,N_24435,N_23116);
xnor U28527 (N_28527,N_23162,N_20336);
xor U28528 (N_28528,N_20282,N_24613);
xor U28529 (N_28529,N_24553,N_24885);
and U28530 (N_28530,N_21522,N_21664);
xor U28531 (N_28531,N_23791,N_22403);
and U28532 (N_28532,N_20855,N_23653);
nand U28533 (N_28533,N_24413,N_22337);
or U28534 (N_28534,N_21208,N_21846);
or U28535 (N_28535,N_23257,N_24207);
nor U28536 (N_28536,N_22027,N_24914);
nand U28537 (N_28537,N_20483,N_20281);
nand U28538 (N_28538,N_23109,N_20788);
nand U28539 (N_28539,N_24271,N_22080);
nand U28540 (N_28540,N_21926,N_23030);
nor U28541 (N_28541,N_20802,N_22659);
xor U28542 (N_28542,N_23563,N_20880);
and U28543 (N_28543,N_21512,N_21555);
or U28544 (N_28544,N_22826,N_21955);
xor U28545 (N_28545,N_24556,N_23908);
and U28546 (N_28546,N_22557,N_20471);
or U28547 (N_28547,N_21051,N_23992);
or U28548 (N_28548,N_22807,N_22508);
nand U28549 (N_28549,N_24745,N_22206);
nor U28550 (N_28550,N_24039,N_24887);
or U28551 (N_28551,N_23068,N_20767);
and U28552 (N_28552,N_21939,N_21696);
and U28553 (N_28553,N_24458,N_22052);
and U28554 (N_28554,N_20185,N_21844);
nand U28555 (N_28555,N_22159,N_24445);
or U28556 (N_28556,N_20421,N_22783);
nor U28557 (N_28557,N_24914,N_24934);
xor U28558 (N_28558,N_20737,N_21157);
and U28559 (N_28559,N_20255,N_20935);
or U28560 (N_28560,N_24487,N_21485);
or U28561 (N_28561,N_20564,N_20813);
xor U28562 (N_28562,N_20959,N_24828);
or U28563 (N_28563,N_24011,N_21131);
or U28564 (N_28564,N_20479,N_23296);
and U28565 (N_28565,N_21829,N_24112);
and U28566 (N_28566,N_24397,N_23551);
or U28567 (N_28567,N_20473,N_21472);
or U28568 (N_28568,N_20603,N_21959);
and U28569 (N_28569,N_20882,N_21785);
or U28570 (N_28570,N_24776,N_20232);
nor U28571 (N_28571,N_20409,N_22158);
and U28572 (N_28572,N_20405,N_21904);
nor U28573 (N_28573,N_20601,N_21081);
or U28574 (N_28574,N_24612,N_23098);
nand U28575 (N_28575,N_21355,N_21189);
or U28576 (N_28576,N_24987,N_23331);
nor U28577 (N_28577,N_22568,N_21428);
or U28578 (N_28578,N_24914,N_23211);
xor U28579 (N_28579,N_20101,N_23750);
and U28580 (N_28580,N_22969,N_20686);
and U28581 (N_28581,N_24902,N_24190);
nor U28582 (N_28582,N_22904,N_20057);
xnor U28583 (N_28583,N_23378,N_22380);
nor U28584 (N_28584,N_24161,N_22921);
nand U28585 (N_28585,N_21888,N_22618);
or U28586 (N_28586,N_21721,N_24091);
and U28587 (N_28587,N_23628,N_24932);
nand U28588 (N_28588,N_22237,N_22999);
or U28589 (N_28589,N_24999,N_21278);
nand U28590 (N_28590,N_20653,N_24162);
and U28591 (N_28591,N_22105,N_22934);
or U28592 (N_28592,N_20243,N_21424);
and U28593 (N_28593,N_24170,N_22238);
and U28594 (N_28594,N_20959,N_20240);
xor U28595 (N_28595,N_21057,N_24610);
or U28596 (N_28596,N_20330,N_23905);
or U28597 (N_28597,N_21977,N_22496);
and U28598 (N_28598,N_21463,N_20190);
xor U28599 (N_28599,N_20286,N_23396);
or U28600 (N_28600,N_23501,N_22049);
and U28601 (N_28601,N_24394,N_21914);
or U28602 (N_28602,N_22240,N_24885);
or U28603 (N_28603,N_20316,N_23170);
nand U28604 (N_28604,N_24958,N_20467);
and U28605 (N_28605,N_23522,N_21573);
nand U28606 (N_28606,N_20538,N_20685);
nand U28607 (N_28607,N_22233,N_24598);
nor U28608 (N_28608,N_20531,N_23765);
nor U28609 (N_28609,N_21315,N_21161);
nand U28610 (N_28610,N_23435,N_23385);
nor U28611 (N_28611,N_20784,N_24439);
or U28612 (N_28612,N_21383,N_21049);
xnor U28613 (N_28613,N_20325,N_22335);
nor U28614 (N_28614,N_21647,N_23909);
and U28615 (N_28615,N_22419,N_24229);
and U28616 (N_28616,N_24959,N_24507);
or U28617 (N_28617,N_20849,N_20837);
nor U28618 (N_28618,N_21640,N_20187);
nor U28619 (N_28619,N_24728,N_23805);
and U28620 (N_28620,N_20767,N_21268);
xnor U28621 (N_28621,N_23034,N_20365);
and U28622 (N_28622,N_21268,N_20679);
or U28623 (N_28623,N_22605,N_24375);
nand U28624 (N_28624,N_21928,N_24755);
and U28625 (N_28625,N_21367,N_20796);
nand U28626 (N_28626,N_23432,N_23546);
or U28627 (N_28627,N_22550,N_21715);
and U28628 (N_28628,N_21127,N_21250);
nand U28629 (N_28629,N_24570,N_24396);
nor U28630 (N_28630,N_21725,N_23938);
and U28631 (N_28631,N_21688,N_22956);
nor U28632 (N_28632,N_22809,N_24823);
or U28633 (N_28633,N_24268,N_22704);
nor U28634 (N_28634,N_23492,N_24523);
and U28635 (N_28635,N_24302,N_20720);
or U28636 (N_28636,N_24340,N_22156);
xor U28637 (N_28637,N_21951,N_24734);
nor U28638 (N_28638,N_20208,N_21335);
nor U28639 (N_28639,N_20677,N_24842);
and U28640 (N_28640,N_22640,N_24258);
nor U28641 (N_28641,N_23880,N_24435);
or U28642 (N_28642,N_24658,N_20425);
nand U28643 (N_28643,N_20796,N_21985);
and U28644 (N_28644,N_21786,N_21746);
nand U28645 (N_28645,N_24642,N_23905);
and U28646 (N_28646,N_23179,N_21646);
xnor U28647 (N_28647,N_20012,N_23999);
or U28648 (N_28648,N_23965,N_20570);
and U28649 (N_28649,N_23298,N_23749);
nand U28650 (N_28650,N_22771,N_20521);
nand U28651 (N_28651,N_24665,N_23315);
and U28652 (N_28652,N_21657,N_22378);
nor U28653 (N_28653,N_24774,N_20969);
xor U28654 (N_28654,N_20248,N_21977);
nor U28655 (N_28655,N_23692,N_22421);
nand U28656 (N_28656,N_20054,N_20609);
and U28657 (N_28657,N_21787,N_20750);
and U28658 (N_28658,N_24703,N_22355);
nand U28659 (N_28659,N_22468,N_24869);
nand U28660 (N_28660,N_21459,N_23677);
and U28661 (N_28661,N_22482,N_22244);
nand U28662 (N_28662,N_24601,N_20263);
and U28663 (N_28663,N_20718,N_23328);
nor U28664 (N_28664,N_23284,N_22000);
or U28665 (N_28665,N_20047,N_21966);
nand U28666 (N_28666,N_22644,N_24278);
xor U28667 (N_28667,N_21967,N_20223);
nand U28668 (N_28668,N_20660,N_24258);
xor U28669 (N_28669,N_23031,N_21787);
xnor U28670 (N_28670,N_22733,N_20427);
and U28671 (N_28671,N_20663,N_24538);
or U28672 (N_28672,N_20024,N_20656);
and U28673 (N_28673,N_21256,N_24738);
nor U28674 (N_28674,N_22003,N_22525);
xnor U28675 (N_28675,N_20414,N_22721);
nor U28676 (N_28676,N_20582,N_22455);
or U28677 (N_28677,N_23615,N_23223);
or U28678 (N_28678,N_23665,N_22443);
and U28679 (N_28679,N_22799,N_20067);
or U28680 (N_28680,N_23322,N_20275);
xnor U28681 (N_28681,N_23613,N_20121);
and U28682 (N_28682,N_22021,N_23782);
nand U28683 (N_28683,N_20868,N_21371);
nor U28684 (N_28684,N_22616,N_22330);
or U28685 (N_28685,N_21672,N_22971);
and U28686 (N_28686,N_23442,N_20019);
or U28687 (N_28687,N_20522,N_21668);
nor U28688 (N_28688,N_21264,N_22314);
and U28689 (N_28689,N_23316,N_20659);
nor U28690 (N_28690,N_24443,N_21761);
nand U28691 (N_28691,N_23508,N_21415);
or U28692 (N_28692,N_24222,N_20239);
nor U28693 (N_28693,N_21561,N_23402);
or U28694 (N_28694,N_23540,N_23173);
nand U28695 (N_28695,N_24797,N_20610);
xor U28696 (N_28696,N_20963,N_24821);
nand U28697 (N_28697,N_22214,N_24737);
xnor U28698 (N_28698,N_23585,N_22264);
nand U28699 (N_28699,N_22095,N_21485);
nand U28700 (N_28700,N_21935,N_21458);
and U28701 (N_28701,N_22104,N_23156);
xnor U28702 (N_28702,N_24641,N_20329);
or U28703 (N_28703,N_21070,N_21699);
or U28704 (N_28704,N_22306,N_23398);
and U28705 (N_28705,N_21823,N_20546);
or U28706 (N_28706,N_20520,N_24191);
nor U28707 (N_28707,N_21153,N_20532);
and U28708 (N_28708,N_23069,N_20559);
and U28709 (N_28709,N_21672,N_21624);
nand U28710 (N_28710,N_24012,N_24946);
or U28711 (N_28711,N_21938,N_21003);
nor U28712 (N_28712,N_20619,N_22121);
or U28713 (N_28713,N_23842,N_24213);
xnor U28714 (N_28714,N_22748,N_20469);
xnor U28715 (N_28715,N_21077,N_24124);
nor U28716 (N_28716,N_23449,N_24525);
or U28717 (N_28717,N_23328,N_24954);
nand U28718 (N_28718,N_24153,N_23392);
or U28719 (N_28719,N_24823,N_21163);
xnor U28720 (N_28720,N_20410,N_22735);
and U28721 (N_28721,N_21497,N_23683);
nor U28722 (N_28722,N_24603,N_24321);
nand U28723 (N_28723,N_21448,N_20801);
xnor U28724 (N_28724,N_20678,N_24401);
xor U28725 (N_28725,N_24820,N_20592);
and U28726 (N_28726,N_23429,N_22370);
nor U28727 (N_28727,N_20521,N_22983);
nor U28728 (N_28728,N_24711,N_22218);
nor U28729 (N_28729,N_23274,N_21768);
and U28730 (N_28730,N_22609,N_22653);
and U28731 (N_28731,N_22590,N_21244);
xor U28732 (N_28732,N_20066,N_24100);
or U28733 (N_28733,N_24416,N_24719);
or U28734 (N_28734,N_23363,N_22089);
nor U28735 (N_28735,N_24431,N_22605);
xnor U28736 (N_28736,N_23765,N_24924);
and U28737 (N_28737,N_21391,N_24390);
nor U28738 (N_28738,N_22718,N_22338);
nor U28739 (N_28739,N_24363,N_22835);
or U28740 (N_28740,N_22862,N_23018);
nor U28741 (N_28741,N_23604,N_20075);
nand U28742 (N_28742,N_22078,N_24949);
nor U28743 (N_28743,N_24449,N_24676);
or U28744 (N_28744,N_22247,N_22234);
or U28745 (N_28745,N_20814,N_24410);
and U28746 (N_28746,N_22300,N_22846);
xnor U28747 (N_28747,N_20349,N_24557);
xor U28748 (N_28748,N_24559,N_21547);
xor U28749 (N_28749,N_24360,N_23676);
nand U28750 (N_28750,N_21672,N_20674);
or U28751 (N_28751,N_24351,N_20440);
xnor U28752 (N_28752,N_22867,N_23431);
nand U28753 (N_28753,N_24383,N_21838);
nand U28754 (N_28754,N_23359,N_21972);
or U28755 (N_28755,N_24412,N_23020);
or U28756 (N_28756,N_23557,N_24459);
xor U28757 (N_28757,N_23017,N_24361);
xor U28758 (N_28758,N_24581,N_22509);
and U28759 (N_28759,N_22839,N_21262);
or U28760 (N_28760,N_21248,N_20264);
nand U28761 (N_28761,N_23678,N_24682);
xnor U28762 (N_28762,N_21409,N_23396);
and U28763 (N_28763,N_21071,N_21274);
and U28764 (N_28764,N_24743,N_20797);
and U28765 (N_28765,N_20545,N_20661);
xnor U28766 (N_28766,N_23582,N_24249);
or U28767 (N_28767,N_21881,N_24381);
nor U28768 (N_28768,N_22491,N_24765);
and U28769 (N_28769,N_22344,N_20196);
xnor U28770 (N_28770,N_21148,N_22340);
and U28771 (N_28771,N_20309,N_22544);
and U28772 (N_28772,N_20698,N_22526);
xor U28773 (N_28773,N_21546,N_21583);
nor U28774 (N_28774,N_22103,N_24752);
and U28775 (N_28775,N_24462,N_20608);
or U28776 (N_28776,N_22366,N_20037);
nand U28777 (N_28777,N_23450,N_21034);
nand U28778 (N_28778,N_24895,N_21690);
or U28779 (N_28779,N_24892,N_20591);
nand U28780 (N_28780,N_23827,N_20963);
and U28781 (N_28781,N_23192,N_22220);
xor U28782 (N_28782,N_20317,N_21222);
nor U28783 (N_28783,N_22996,N_22807);
nand U28784 (N_28784,N_21056,N_24743);
and U28785 (N_28785,N_24518,N_24554);
nand U28786 (N_28786,N_24129,N_24212);
and U28787 (N_28787,N_24552,N_20604);
nor U28788 (N_28788,N_23496,N_24580);
or U28789 (N_28789,N_21952,N_24492);
or U28790 (N_28790,N_21117,N_20754);
and U28791 (N_28791,N_20545,N_23223);
nor U28792 (N_28792,N_20001,N_20000);
nand U28793 (N_28793,N_23576,N_22227);
xnor U28794 (N_28794,N_23257,N_22249);
xnor U28795 (N_28795,N_20517,N_21605);
nor U28796 (N_28796,N_20468,N_23583);
xor U28797 (N_28797,N_21452,N_21935);
and U28798 (N_28798,N_24284,N_21166);
nor U28799 (N_28799,N_24292,N_23260);
nor U28800 (N_28800,N_23421,N_21187);
nor U28801 (N_28801,N_20911,N_23512);
xnor U28802 (N_28802,N_21735,N_22874);
xor U28803 (N_28803,N_20489,N_24940);
and U28804 (N_28804,N_22597,N_23488);
nand U28805 (N_28805,N_23292,N_21292);
and U28806 (N_28806,N_20583,N_21150);
and U28807 (N_28807,N_24668,N_21407);
nand U28808 (N_28808,N_23871,N_22866);
xnor U28809 (N_28809,N_23523,N_21111);
xnor U28810 (N_28810,N_23704,N_20445);
xnor U28811 (N_28811,N_23762,N_21851);
or U28812 (N_28812,N_24525,N_24156);
nor U28813 (N_28813,N_20153,N_22631);
nand U28814 (N_28814,N_22430,N_21234);
xnor U28815 (N_28815,N_21283,N_22642);
and U28816 (N_28816,N_21784,N_22291);
xnor U28817 (N_28817,N_21061,N_23889);
nand U28818 (N_28818,N_22236,N_22776);
nand U28819 (N_28819,N_21747,N_23290);
nand U28820 (N_28820,N_24797,N_21917);
and U28821 (N_28821,N_20828,N_21033);
nand U28822 (N_28822,N_20638,N_23758);
nor U28823 (N_28823,N_20723,N_24805);
nor U28824 (N_28824,N_23302,N_20364);
nand U28825 (N_28825,N_22261,N_23178);
nand U28826 (N_28826,N_24224,N_23572);
nor U28827 (N_28827,N_22540,N_22211);
and U28828 (N_28828,N_20767,N_20121);
and U28829 (N_28829,N_23580,N_22762);
and U28830 (N_28830,N_23582,N_24115);
nor U28831 (N_28831,N_20010,N_22124);
and U28832 (N_28832,N_20967,N_20243);
xor U28833 (N_28833,N_23764,N_23210);
nand U28834 (N_28834,N_24986,N_21434);
or U28835 (N_28835,N_21501,N_21473);
and U28836 (N_28836,N_23188,N_20347);
nor U28837 (N_28837,N_24055,N_20491);
nand U28838 (N_28838,N_22904,N_20744);
nor U28839 (N_28839,N_21728,N_22406);
nand U28840 (N_28840,N_23813,N_23759);
or U28841 (N_28841,N_24527,N_24978);
xnor U28842 (N_28842,N_20370,N_21958);
and U28843 (N_28843,N_22903,N_22462);
nor U28844 (N_28844,N_20943,N_20738);
xnor U28845 (N_28845,N_24740,N_24030);
or U28846 (N_28846,N_23671,N_24564);
nand U28847 (N_28847,N_24144,N_24753);
nor U28848 (N_28848,N_23777,N_23763);
or U28849 (N_28849,N_20938,N_21476);
or U28850 (N_28850,N_21036,N_22941);
or U28851 (N_28851,N_23655,N_20030);
and U28852 (N_28852,N_21238,N_23755);
nor U28853 (N_28853,N_23253,N_23183);
xor U28854 (N_28854,N_24269,N_21629);
or U28855 (N_28855,N_22807,N_24421);
or U28856 (N_28856,N_20180,N_22851);
and U28857 (N_28857,N_22568,N_20128);
or U28858 (N_28858,N_24972,N_20276);
nand U28859 (N_28859,N_22145,N_21282);
and U28860 (N_28860,N_21461,N_20438);
or U28861 (N_28861,N_20135,N_20506);
nor U28862 (N_28862,N_24858,N_20651);
nor U28863 (N_28863,N_22275,N_20878);
nor U28864 (N_28864,N_24909,N_20135);
or U28865 (N_28865,N_24495,N_22746);
or U28866 (N_28866,N_20844,N_20294);
or U28867 (N_28867,N_20122,N_23425);
nand U28868 (N_28868,N_23035,N_20128);
and U28869 (N_28869,N_23070,N_21774);
and U28870 (N_28870,N_20745,N_20603);
and U28871 (N_28871,N_20861,N_22011);
nand U28872 (N_28872,N_21697,N_23397);
nand U28873 (N_28873,N_20819,N_20447);
and U28874 (N_28874,N_23231,N_20642);
and U28875 (N_28875,N_21377,N_22163);
nand U28876 (N_28876,N_21904,N_22724);
nand U28877 (N_28877,N_24412,N_20614);
or U28878 (N_28878,N_22077,N_22011);
or U28879 (N_28879,N_20176,N_23460);
nand U28880 (N_28880,N_20157,N_24163);
xor U28881 (N_28881,N_22695,N_22044);
xnor U28882 (N_28882,N_23265,N_23178);
and U28883 (N_28883,N_24470,N_21726);
nand U28884 (N_28884,N_21939,N_21694);
and U28885 (N_28885,N_20237,N_20276);
nor U28886 (N_28886,N_22800,N_24416);
or U28887 (N_28887,N_22005,N_23638);
or U28888 (N_28888,N_24627,N_21991);
or U28889 (N_28889,N_20566,N_21193);
xor U28890 (N_28890,N_23331,N_21742);
nand U28891 (N_28891,N_22705,N_24878);
and U28892 (N_28892,N_20906,N_21691);
and U28893 (N_28893,N_23469,N_24064);
xnor U28894 (N_28894,N_24754,N_24858);
or U28895 (N_28895,N_23068,N_21165);
or U28896 (N_28896,N_21277,N_24100);
or U28897 (N_28897,N_20657,N_21363);
and U28898 (N_28898,N_21438,N_24487);
nor U28899 (N_28899,N_22728,N_21819);
or U28900 (N_28900,N_24003,N_23384);
nand U28901 (N_28901,N_22038,N_22461);
xor U28902 (N_28902,N_22853,N_20822);
nor U28903 (N_28903,N_23600,N_24482);
or U28904 (N_28904,N_24277,N_23049);
or U28905 (N_28905,N_20655,N_21508);
or U28906 (N_28906,N_20435,N_23586);
nand U28907 (N_28907,N_24908,N_21722);
nand U28908 (N_28908,N_21963,N_20781);
nand U28909 (N_28909,N_24756,N_23120);
or U28910 (N_28910,N_20622,N_21251);
xnor U28911 (N_28911,N_22667,N_20694);
nand U28912 (N_28912,N_20358,N_23238);
or U28913 (N_28913,N_23453,N_21443);
nor U28914 (N_28914,N_20419,N_20505);
and U28915 (N_28915,N_22064,N_23062);
xnor U28916 (N_28916,N_22770,N_23395);
and U28917 (N_28917,N_20657,N_21191);
or U28918 (N_28918,N_23427,N_20159);
and U28919 (N_28919,N_24534,N_20495);
xnor U28920 (N_28920,N_23820,N_24917);
or U28921 (N_28921,N_21421,N_21589);
xor U28922 (N_28922,N_20203,N_23143);
xor U28923 (N_28923,N_20312,N_20024);
or U28924 (N_28924,N_20331,N_21205);
or U28925 (N_28925,N_22750,N_21498);
and U28926 (N_28926,N_23622,N_24604);
nand U28927 (N_28927,N_20094,N_20072);
or U28928 (N_28928,N_20343,N_20970);
nand U28929 (N_28929,N_20084,N_21944);
and U28930 (N_28930,N_21862,N_24392);
xnor U28931 (N_28931,N_21127,N_20782);
and U28932 (N_28932,N_21934,N_22010);
and U28933 (N_28933,N_23831,N_21060);
xnor U28934 (N_28934,N_23760,N_20928);
nor U28935 (N_28935,N_24546,N_24203);
and U28936 (N_28936,N_22253,N_24586);
xor U28937 (N_28937,N_22496,N_23519);
and U28938 (N_28938,N_22311,N_22307);
nor U28939 (N_28939,N_20624,N_23884);
and U28940 (N_28940,N_22113,N_21107);
nand U28941 (N_28941,N_22264,N_21747);
xnor U28942 (N_28942,N_21760,N_22728);
or U28943 (N_28943,N_20823,N_22745);
xor U28944 (N_28944,N_23465,N_24852);
nor U28945 (N_28945,N_21414,N_22919);
xnor U28946 (N_28946,N_24691,N_21420);
nand U28947 (N_28947,N_22401,N_21546);
and U28948 (N_28948,N_23576,N_20343);
nand U28949 (N_28949,N_22797,N_24382);
and U28950 (N_28950,N_21810,N_21110);
or U28951 (N_28951,N_24625,N_24066);
xor U28952 (N_28952,N_21516,N_20437);
or U28953 (N_28953,N_22361,N_22521);
nand U28954 (N_28954,N_22687,N_20165);
or U28955 (N_28955,N_21142,N_21238);
nor U28956 (N_28956,N_22472,N_24149);
or U28957 (N_28957,N_23492,N_21080);
xnor U28958 (N_28958,N_24924,N_21445);
and U28959 (N_28959,N_24605,N_24756);
and U28960 (N_28960,N_21449,N_23512);
and U28961 (N_28961,N_21790,N_22966);
and U28962 (N_28962,N_24702,N_21996);
or U28963 (N_28963,N_22260,N_24657);
nor U28964 (N_28964,N_24165,N_23597);
and U28965 (N_28965,N_24556,N_23709);
nand U28966 (N_28966,N_20446,N_22745);
or U28967 (N_28967,N_22889,N_20022);
nor U28968 (N_28968,N_22449,N_22641);
nor U28969 (N_28969,N_23013,N_20262);
nand U28970 (N_28970,N_21849,N_20796);
and U28971 (N_28971,N_22479,N_22360);
and U28972 (N_28972,N_20492,N_23583);
nand U28973 (N_28973,N_22051,N_22778);
xnor U28974 (N_28974,N_24423,N_24322);
nand U28975 (N_28975,N_23320,N_24293);
or U28976 (N_28976,N_21377,N_23825);
xnor U28977 (N_28977,N_24954,N_24603);
or U28978 (N_28978,N_23947,N_22107);
nor U28979 (N_28979,N_23427,N_23906);
and U28980 (N_28980,N_24889,N_24860);
or U28981 (N_28981,N_24289,N_20744);
nand U28982 (N_28982,N_24169,N_20107);
or U28983 (N_28983,N_22216,N_23600);
or U28984 (N_28984,N_20248,N_23577);
nor U28985 (N_28985,N_21832,N_20564);
nor U28986 (N_28986,N_23610,N_24179);
nand U28987 (N_28987,N_24997,N_21076);
and U28988 (N_28988,N_24095,N_24080);
xnor U28989 (N_28989,N_24337,N_23726);
xnor U28990 (N_28990,N_24708,N_20652);
and U28991 (N_28991,N_24387,N_22166);
xor U28992 (N_28992,N_22388,N_24023);
nand U28993 (N_28993,N_22026,N_23274);
or U28994 (N_28994,N_23317,N_23678);
xor U28995 (N_28995,N_21242,N_24682);
nand U28996 (N_28996,N_22796,N_22076);
nor U28997 (N_28997,N_24470,N_22335);
and U28998 (N_28998,N_24378,N_22871);
nor U28999 (N_28999,N_21942,N_22245);
nor U29000 (N_29000,N_21312,N_20390);
and U29001 (N_29001,N_24820,N_23101);
or U29002 (N_29002,N_23275,N_21139);
xor U29003 (N_29003,N_24364,N_21099);
xor U29004 (N_29004,N_21803,N_24677);
nand U29005 (N_29005,N_23429,N_24374);
xor U29006 (N_29006,N_22537,N_20490);
and U29007 (N_29007,N_23514,N_23559);
nand U29008 (N_29008,N_23147,N_21060);
nand U29009 (N_29009,N_20649,N_22987);
and U29010 (N_29010,N_24481,N_24551);
or U29011 (N_29011,N_20319,N_23484);
nor U29012 (N_29012,N_23434,N_23943);
and U29013 (N_29013,N_23240,N_24408);
and U29014 (N_29014,N_22011,N_23326);
nand U29015 (N_29015,N_23030,N_21951);
nor U29016 (N_29016,N_21585,N_22762);
nand U29017 (N_29017,N_21556,N_21699);
nor U29018 (N_29018,N_20065,N_23614);
nor U29019 (N_29019,N_21899,N_21949);
nor U29020 (N_29020,N_23434,N_20252);
or U29021 (N_29021,N_22499,N_24674);
or U29022 (N_29022,N_20122,N_24474);
nand U29023 (N_29023,N_23850,N_20101);
nand U29024 (N_29024,N_24623,N_22204);
nand U29025 (N_29025,N_21399,N_21048);
nand U29026 (N_29026,N_22863,N_24709);
or U29027 (N_29027,N_22986,N_22818);
and U29028 (N_29028,N_22689,N_24496);
xor U29029 (N_29029,N_22792,N_20231);
and U29030 (N_29030,N_22183,N_20677);
nor U29031 (N_29031,N_20330,N_24693);
xnor U29032 (N_29032,N_22042,N_24895);
and U29033 (N_29033,N_24145,N_21714);
and U29034 (N_29034,N_24777,N_23393);
nor U29035 (N_29035,N_21795,N_22407);
nand U29036 (N_29036,N_21314,N_24486);
xnor U29037 (N_29037,N_24971,N_23894);
or U29038 (N_29038,N_21029,N_20616);
and U29039 (N_29039,N_22024,N_22557);
or U29040 (N_29040,N_23183,N_23053);
nand U29041 (N_29041,N_23347,N_21159);
or U29042 (N_29042,N_20306,N_23878);
nand U29043 (N_29043,N_22880,N_20153);
nand U29044 (N_29044,N_24058,N_20579);
xnor U29045 (N_29045,N_24662,N_22404);
xnor U29046 (N_29046,N_20436,N_22693);
nand U29047 (N_29047,N_24910,N_23840);
or U29048 (N_29048,N_23139,N_23980);
and U29049 (N_29049,N_21089,N_24459);
nor U29050 (N_29050,N_24386,N_20180);
xnor U29051 (N_29051,N_22778,N_24023);
and U29052 (N_29052,N_21971,N_22417);
and U29053 (N_29053,N_24712,N_20228);
or U29054 (N_29054,N_20598,N_23271);
nor U29055 (N_29055,N_20675,N_21695);
or U29056 (N_29056,N_24329,N_22862);
nor U29057 (N_29057,N_21305,N_22550);
xnor U29058 (N_29058,N_24797,N_23788);
xor U29059 (N_29059,N_21616,N_21658);
and U29060 (N_29060,N_24845,N_23568);
and U29061 (N_29061,N_23469,N_24068);
nand U29062 (N_29062,N_21323,N_24171);
xnor U29063 (N_29063,N_20756,N_24090);
or U29064 (N_29064,N_22705,N_23208);
nand U29065 (N_29065,N_24931,N_24259);
or U29066 (N_29066,N_23435,N_21878);
or U29067 (N_29067,N_23765,N_24006);
nor U29068 (N_29068,N_20662,N_20902);
nand U29069 (N_29069,N_22819,N_23601);
nand U29070 (N_29070,N_20710,N_23099);
nand U29071 (N_29071,N_24428,N_20812);
xnor U29072 (N_29072,N_20382,N_20028);
and U29073 (N_29073,N_24926,N_21063);
and U29074 (N_29074,N_24003,N_20305);
nor U29075 (N_29075,N_23331,N_22881);
nand U29076 (N_29076,N_21590,N_22763);
nand U29077 (N_29077,N_24391,N_23347);
and U29078 (N_29078,N_21549,N_21118);
nand U29079 (N_29079,N_23053,N_22283);
and U29080 (N_29080,N_21302,N_21588);
nand U29081 (N_29081,N_22340,N_22443);
or U29082 (N_29082,N_24401,N_22554);
and U29083 (N_29083,N_22388,N_24862);
nor U29084 (N_29084,N_21966,N_21412);
and U29085 (N_29085,N_23560,N_20778);
nand U29086 (N_29086,N_23077,N_23392);
and U29087 (N_29087,N_20197,N_21458);
and U29088 (N_29088,N_22242,N_22003);
nand U29089 (N_29089,N_23488,N_21172);
nor U29090 (N_29090,N_22046,N_24349);
xnor U29091 (N_29091,N_22941,N_21198);
nor U29092 (N_29092,N_21229,N_22853);
xor U29093 (N_29093,N_21272,N_23511);
and U29094 (N_29094,N_20859,N_23338);
or U29095 (N_29095,N_22058,N_22987);
nand U29096 (N_29096,N_20568,N_21713);
nor U29097 (N_29097,N_20469,N_20563);
nand U29098 (N_29098,N_20059,N_20566);
and U29099 (N_29099,N_22347,N_22257);
xnor U29100 (N_29100,N_22791,N_24370);
or U29101 (N_29101,N_21756,N_22514);
xor U29102 (N_29102,N_20793,N_23182);
nand U29103 (N_29103,N_21687,N_21244);
and U29104 (N_29104,N_21774,N_24144);
nand U29105 (N_29105,N_24234,N_20309);
nor U29106 (N_29106,N_21573,N_24761);
nor U29107 (N_29107,N_23023,N_21621);
and U29108 (N_29108,N_21928,N_23574);
nor U29109 (N_29109,N_23858,N_23228);
nand U29110 (N_29110,N_23332,N_20707);
nor U29111 (N_29111,N_23261,N_22826);
nand U29112 (N_29112,N_21343,N_23267);
nand U29113 (N_29113,N_23344,N_24074);
nand U29114 (N_29114,N_20788,N_23447);
nand U29115 (N_29115,N_21699,N_23045);
xnor U29116 (N_29116,N_23057,N_23967);
nor U29117 (N_29117,N_22548,N_23179);
and U29118 (N_29118,N_22348,N_23788);
xnor U29119 (N_29119,N_22152,N_22097);
or U29120 (N_29120,N_22247,N_21124);
nand U29121 (N_29121,N_22921,N_22658);
and U29122 (N_29122,N_21514,N_20657);
or U29123 (N_29123,N_24373,N_24313);
nor U29124 (N_29124,N_23043,N_21899);
nand U29125 (N_29125,N_22496,N_22655);
and U29126 (N_29126,N_20076,N_24070);
nand U29127 (N_29127,N_22756,N_22431);
and U29128 (N_29128,N_20385,N_22445);
xnor U29129 (N_29129,N_24948,N_21662);
and U29130 (N_29130,N_23252,N_23477);
nand U29131 (N_29131,N_23318,N_24746);
nand U29132 (N_29132,N_20007,N_24846);
nor U29133 (N_29133,N_22521,N_22061);
nor U29134 (N_29134,N_20446,N_22535);
nor U29135 (N_29135,N_24155,N_20176);
nor U29136 (N_29136,N_24004,N_22447);
and U29137 (N_29137,N_24352,N_20587);
nand U29138 (N_29138,N_23823,N_21455);
xor U29139 (N_29139,N_21311,N_23161);
and U29140 (N_29140,N_22649,N_24260);
and U29141 (N_29141,N_20373,N_20356);
xor U29142 (N_29142,N_21220,N_23602);
nand U29143 (N_29143,N_23890,N_24687);
nand U29144 (N_29144,N_23258,N_23564);
and U29145 (N_29145,N_23435,N_21434);
nor U29146 (N_29146,N_22356,N_20935);
and U29147 (N_29147,N_20565,N_22618);
and U29148 (N_29148,N_24797,N_24180);
nand U29149 (N_29149,N_21692,N_24353);
nand U29150 (N_29150,N_21143,N_22624);
xor U29151 (N_29151,N_20531,N_22228);
or U29152 (N_29152,N_23235,N_21746);
nor U29153 (N_29153,N_20613,N_21162);
nor U29154 (N_29154,N_21157,N_20227);
nand U29155 (N_29155,N_21512,N_20800);
and U29156 (N_29156,N_22870,N_22880);
nor U29157 (N_29157,N_20802,N_23622);
nand U29158 (N_29158,N_21155,N_20390);
nand U29159 (N_29159,N_23650,N_22245);
xnor U29160 (N_29160,N_23419,N_20791);
or U29161 (N_29161,N_24823,N_21184);
xor U29162 (N_29162,N_22606,N_20137);
or U29163 (N_29163,N_22102,N_22886);
xor U29164 (N_29164,N_23797,N_22297);
nand U29165 (N_29165,N_22589,N_21435);
nor U29166 (N_29166,N_23353,N_21863);
nor U29167 (N_29167,N_22034,N_23948);
nand U29168 (N_29168,N_23652,N_23304);
and U29169 (N_29169,N_20052,N_21734);
xor U29170 (N_29170,N_20975,N_21842);
or U29171 (N_29171,N_22933,N_21220);
xnor U29172 (N_29172,N_24945,N_23214);
or U29173 (N_29173,N_20341,N_22597);
nor U29174 (N_29174,N_23374,N_22296);
nand U29175 (N_29175,N_20493,N_20142);
or U29176 (N_29176,N_24444,N_23670);
nor U29177 (N_29177,N_20792,N_22568);
xnor U29178 (N_29178,N_20382,N_23598);
or U29179 (N_29179,N_20777,N_23280);
or U29180 (N_29180,N_24435,N_23723);
nand U29181 (N_29181,N_22882,N_20715);
or U29182 (N_29182,N_23390,N_20721);
xor U29183 (N_29183,N_24226,N_22116);
xor U29184 (N_29184,N_20595,N_24930);
or U29185 (N_29185,N_24240,N_22201);
nand U29186 (N_29186,N_20448,N_21908);
xor U29187 (N_29187,N_20869,N_24871);
and U29188 (N_29188,N_21417,N_24853);
nor U29189 (N_29189,N_20776,N_22476);
xnor U29190 (N_29190,N_20532,N_23416);
nand U29191 (N_29191,N_22171,N_20478);
nor U29192 (N_29192,N_24970,N_20000);
xnor U29193 (N_29193,N_20507,N_23475);
xor U29194 (N_29194,N_20962,N_21017);
xor U29195 (N_29195,N_21177,N_22860);
nand U29196 (N_29196,N_24603,N_21199);
or U29197 (N_29197,N_23807,N_24403);
or U29198 (N_29198,N_20755,N_22897);
or U29199 (N_29199,N_23268,N_24058);
nor U29200 (N_29200,N_22611,N_20596);
or U29201 (N_29201,N_21305,N_20973);
xor U29202 (N_29202,N_21217,N_23300);
nor U29203 (N_29203,N_23474,N_21007);
xor U29204 (N_29204,N_21907,N_20930);
and U29205 (N_29205,N_23410,N_24850);
or U29206 (N_29206,N_22456,N_23040);
and U29207 (N_29207,N_24246,N_22238);
nand U29208 (N_29208,N_20540,N_21339);
and U29209 (N_29209,N_24149,N_23333);
and U29210 (N_29210,N_20296,N_20527);
nor U29211 (N_29211,N_22967,N_24070);
nor U29212 (N_29212,N_22903,N_22150);
and U29213 (N_29213,N_20708,N_23940);
and U29214 (N_29214,N_20702,N_20858);
and U29215 (N_29215,N_22401,N_20116);
xnor U29216 (N_29216,N_24259,N_23450);
nand U29217 (N_29217,N_22973,N_23944);
nand U29218 (N_29218,N_22098,N_20843);
and U29219 (N_29219,N_20677,N_21386);
xnor U29220 (N_29220,N_21282,N_23554);
xor U29221 (N_29221,N_23808,N_23522);
and U29222 (N_29222,N_22238,N_24444);
nand U29223 (N_29223,N_21583,N_23364);
nor U29224 (N_29224,N_21354,N_23310);
nor U29225 (N_29225,N_24591,N_20702);
and U29226 (N_29226,N_23033,N_20787);
or U29227 (N_29227,N_21831,N_22543);
xor U29228 (N_29228,N_23942,N_21542);
and U29229 (N_29229,N_23310,N_24320);
xor U29230 (N_29230,N_20880,N_20947);
xnor U29231 (N_29231,N_21158,N_21616);
and U29232 (N_29232,N_20691,N_23135);
and U29233 (N_29233,N_23864,N_22333);
xnor U29234 (N_29234,N_24034,N_23042);
and U29235 (N_29235,N_24186,N_22995);
nor U29236 (N_29236,N_24448,N_23339);
and U29237 (N_29237,N_20713,N_22730);
xnor U29238 (N_29238,N_21135,N_24259);
nor U29239 (N_29239,N_21017,N_23766);
or U29240 (N_29240,N_21335,N_22785);
nor U29241 (N_29241,N_24289,N_22862);
and U29242 (N_29242,N_22325,N_21314);
and U29243 (N_29243,N_20978,N_21879);
or U29244 (N_29244,N_24865,N_22879);
nand U29245 (N_29245,N_24625,N_22995);
or U29246 (N_29246,N_24227,N_22337);
nand U29247 (N_29247,N_23865,N_21553);
or U29248 (N_29248,N_21507,N_23206);
nand U29249 (N_29249,N_20137,N_24599);
nor U29250 (N_29250,N_24348,N_24662);
or U29251 (N_29251,N_22553,N_23970);
nand U29252 (N_29252,N_24993,N_20015);
nor U29253 (N_29253,N_23819,N_22417);
xor U29254 (N_29254,N_21421,N_20881);
xnor U29255 (N_29255,N_20644,N_22793);
and U29256 (N_29256,N_24909,N_20012);
nor U29257 (N_29257,N_22745,N_22482);
or U29258 (N_29258,N_23552,N_22153);
nor U29259 (N_29259,N_22771,N_21800);
xor U29260 (N_29260,N_22395,N_20491);
nor U29261 (N_29261,N_23218,N_21174);
xnor U29262 (N_29262,N_23228,N_22303);
and U29263 (N_29263,N_23229,N_23801);
and U29264 (N_29264,N_22243,N_20017);
xor U29265 (N_29265,N_20116,N_20633);
nor U29266 (N_29266,N_22925,N_20622);
xor U29267 (N_29267,N_21567,N_24130);
or U29268 (N_29268,N_24317,N_22205);
nand U29269 (N_29269,N_24175,N_20103);
xnor U29270 (N_29270,N_23808,N_24251);
nand U29271 (N_29271,N_22550,N_20608);
nand U29272 (N_29272,N_24976,N_21822);
nand U29273 (N_29273,N_24078,N_20222);
xor U29274 (N_29274,N_24505,N_22931);
and U29275 (N_29275,N_23172,N_21961);
or U29276 (N_29276,N_22429,N_24443);
and U29277 (N_29277,N_20644,N_20371);
nor U29278 (N_29278,N_21026,N_20187);
nor U29279 (N_29279,N_24537,N_23203);
nand U29280 (N_29280,N_23096,N_21354);
or U29281 (N_29281,N_22699,N_22746);
and U29282 (N_29282,N_22554,N_24279);
nor U29283 (N_29283,N_22767,N_24760);
nor U29284 (N_29284,N_22900,N_21527);
or U29285 (N_29285,N_24589,N_23436);
nand U29286 (N_29286,N_24442,N_22850);
xnor U29287 (N_29287,N_24033,N_23307);
nor U29288 (N_29288,N_22850,N_24266);
or U29289 (N_29289,N_24848,N_21110);
nor U29290 (N_29290,N_20514,N_22702);
nand U29291 (N_29291,N_23756,N_20634);
nor U29292 (N_29292,N_24349,N_20889);
nand U29293 (N_29293,N_24043,N_22830);
or U29294 (N_29294,N_22967,N_21539);
nand U29295 (N_29295,N_21305,N_20926);
or U29296 (N_29296,N_21405,N_20292);
and U29297 (N_29297,N_20162,N_20353);
nor U29298 (N_29298,N_21472,N_24821);
nor U29299 (N_29299,N_20695,N_20554);
nand U29300 (N_29300,N_20686,N_22197);
nand U29301 (N_29301,N_23727,N_23805);
nand U29302 (N_29302,N_20583,N_20663);
or U29303 (N_29303,N_22213,N_20462);
and U29304 (N_29304,N_21511,N_22074);
nor U29305 (N_29305,N_23808,N_23445);
and U29306 (N_29306,N_24183,N_23416);
nand U29307 (N_29307,N_21728,N_20344);
nand U29308 (N_29308,N_21867,N_22602);
nor U29309 (N_29309,N_24156,N_24974);
or U29310 (N_29310,N_24695,N_21273);
or U29311 (N_29311,N_24040,N_22324);
xnor U29312 (N_29312,N_22563,N_24185);
and U29313 (N_29313,N_20383,N_23029);
and U29314 (N_29314,N_21434,N_20368);
or U29315 (N_29315,N_21063,N_20644);
and U29316 (N_29316,N_24792,N_24222);
xnor U29317 (N_29317,N_22073,N_20913);
or U29318 (N_29318,N_21562,N_23500);
nand U29319 (N_29319,N_23015,N_22713);
nor U29320 (N_29320,N_23928,N_23422);
xor U29321 (N_29321,N_21873,N_20297);
or U29322 (N_29322,N_24655,N_22842);
nor U29323 (N_29323,N_24284,N_23086);
or U29324 (N_29324,N_24410,N_21651);
nand U29325 (N_29325,N_22855,N_20268);
xnor U29326 (N_29326,N_22662,N_22916);
or U29327 (N_29327,N_22931,N_24147);
or U29328 (N_29328,N_22352,N_22680);
nand U29329 (N_29329,N_20967,N_21959);
nand U29330 (N_29330,N_24622,N_21967);
or U29331 (N_29331,N_20762,N_24454);
or U29332 (N_29332,N_24685,N_21199);
nand U29333 (N_29333,N_23349,N_24889);
nor U29334 (N_29334,N_20527,N_21787);
and U29335 (N_29335,N_23581,N_21915);
or U29336 (N_29336,N_24084,N_21171);
nand U29337 (N_29337,N_21601,N_22856);
nand U29338 (N_29338,N_21013,N_20880);
and U29339 (N_29339,N_23242,N_23219);
nand U29340 (N_29340,N_24580,N_23637);
xnor U29341 (N_29341,N_21156,N_20787);
nor U29342 (N_29342,N_20684,N_22756);
nand U29343 (N_29343,N_22191,N_22566);
nor U29344 (N_29344,N_21605,N_21194);
nand U29345 (N_29345,N_24164,N_21294);
xor U29346 (N_29346,N_22521,N_21758);
nand U29347 (N_29347,N_23213,N_24599);
nand U29348 (N_29348,N_21243,N_22598);
nand U29349 (N_29349,N_21165,N_23309);
nand U29350 (N_29350,N_21707,N_24499);
xnor U29351 (N_29351,N_23427,N_20597);
nand U29352 (N_29352,N_22476,N_20340);
nand U29353 (N_29353,N_22917,N_20357);
nor U29354 (N_29354,N_21204,N_20348);
and U29355 (N_29355,N_24831,N_24682);
xor U29356 (N_29356,N_20482,N_20968);
nor U29357 (N_29357,N_24711,N_24035);
nor U29358 (N_29358,N_23638,N_23783);
nand U29359 (N_29359,N_24155,N_24197);
and U29360 (N_29360,N_20272,N_21560);
and U29361 (N_29361,N_22834,N_23344);
nand U29362 (N_29362,N_20289,N_23241);
nand U29363 (N_29363,N_24917,N_24450);
and U29364 (N_29364,N_20206,N_23453);
xnor U29365 (N_29365,N_20211,N_20420);
nor U29366 (N_29366,N_21457,N_24754);
xor U29367 (N_29367,N_21659,N_24612);
nand U29368 (N_29368,N_24111,N_23782);
or U29369 (N_29369,N_23811,N_21195);
or U29370 (N_29370,N_24657,N_22485);
and U29371 (N_29371,N_21325,N_23095);
nor U29372 (N_29372,N_24146,N_23158);
and U29373 (N_29373,N_23819,N_22522);
nor U29374 (N_29374,N_22916,N_20607);
xor U29375 (N_29375,N_22689,N_23005);
nand U29376 (N_29376,N_24960,N_22922);
or U29377 (N_29377,N_24324,N_21991);
or U29378 (N_29378,N_23508,N_20619);
xnor U29379 (N_29379,N_23356,N_24963);
or U29380 (N_29380,N_23583,N_23538);
xnor U29381 (N_29381,N_20186,N_21104);
nor U29382 (N_29382,N_23218,N_24700);
xor U29383 (N_29383,N_20821,N_23502);
or U29384 (N_29384,N_21782,N_21901);
and U29385 (N_29385,N_20288,N_22069);
and U29386 (N_29386,N_23775,N_23652);
xnor U29387 (N_29387,N_21785,N_21174);
xor U29388 (N_29388,N_20652,N_24382);
or U29389 (N_29389,N_23150,N_24873);
and U29390 (N_29390,N_20398,N_22065);
xor U29391 (N_29391,N_23493,N_23660);
nand U29392 (N_29392,N_23730,N_23319);
or U29393 (N_29393,N_24763,N_23840);
nand U29394 (N_29394,N_22231,N_21780);
and U29395 (N_29395,N_22969,N_24919);
xnor U29396 (N_29396,N_20272,N_23168);
nand U29397 (N_29397,N_22946,N_24970);
and U29398 (N_29398,N_22918,N_20232);
and U29399 (N_29399,N_22348,N_21611);
and U29400 (N_29400,N_20508,N_21004);
or U29401 (N_29401,N_21404,N_20819);
xnor U29402 (N_29402,N_22281,N_23508);
nor U29403 (N_29403,N_23365,N_22880);
nand U29404 (N_29404,N_22591,N_21978);
xnor U29405 (N_29405,N_22121,N_24261);
or U29406 (N_29406,N_20093,N_20758);
xor U29407 (N_29407,N_21928,N_23408);
xor U29408 (N_29408,N_24679,N_24527);
and U29409 (N_29409,N_22360,N_20056);
nand U29410 (N_29410,N_24314,N_23206);
and U29411 (N_29411,N_22688,N_21531);
nand U29412 (N_29412,N_21165,N_22549);
nor U29413 (N_29413,N_20565,N_20687);
nand U29414 (N_29414,N_21125,N_22675);
or U29415 (N_29415,N_21169,N_23584);
nand U29416 (N_29416,N_20306,N_23901);
xor U29417 (N_29417,N_22508,N_20414);
nand U29418 (N_29418,N_21294,N_23777);
xnor U29419 (N_29419,N_20884,N_23623);
nand U29420 (N_29420,N_24716,N_20920);
nor U29421 (N_29421,N_23961,N_22548);
nand U29422 (N_29422,N_24805,N_21209);
xnor U29423 (N_29423,N_20124,N_23028);
xnor U29424 (N_29424,N_24875,N_23530);
and U29425 (N_29425,N_22573,N_20321);
nand U29426 (N_29426,N_22310,N_20844);
xor U29427 (N_29427,N_22114,N_24690);
or U29428 (N_29428,N_22322,N_24501);
xor U29429 (N_29429,N_24405,N_23338);
and U29430 (N_29430,N_20198,N_23860);
nand U29431 (N_29431,N_24279,N_23932);
nor U29432 (N_29432,N_23164,N_21596);
nand U29433 (N_29433,N_21243,N_24720);
xor U29434 (N_29434,N_21973,N_20692);
or U29435 (N_29435,N_20121,N_22886);
nand U29436 (N_29436,N_21732,N_22972);
xor U29437 (N_29437,N_23299,N_24228);
nand U29438 (N_29438,N_23561,N_21526);
nor U29439 (N_29439,N_23788,N_22373);
nand U29440 (N_29440,N_23481,N_24349);
and U29441 (N_29441,N_20160,N_21209);
nand U29442 (N_29442,N_20055,N_24281);
or U29443 (N_29443,N_22368,N_22752);
nor U29444 (N_29444,N_21444,N_23567);
nand U29445 (N_29445,N_24973,N_21174);
and U29446 (N_29446,N_23726,N_21971);
xor U29447 (N_29447,N_24883,N_23294);
nand U29448 (N_29448,N_24553,N_23230);
nand U29449 (N_29449,N_22742,N_20950);
nor U29450 (N_29450,N_22373,N_23862);
and U29451 (N_29451,N_22938,N_21840);
nor U29452 (N_29452,N_23382,N_22703);
nor U29453 (N_29453,N_22954,N_24848);
or U29454 (N_29454,N_20763,N_21344);
nor U29455 (N_29455,N_21984,N_23702);
or U29456 (N_29456,N_22473,N_24529);
or U29457 (N_29457,N_24177,N_22967);
or U29458 (N_29458,N_20680,N_20926);
nand U29459 (N_29459,N_22179,N_22263);
nand U29460 (N_29460,N_22076,N_24133);
and U29461 (N_29461,N_24458,N_24586);
and U29462 (N_29462,N_22794,N_24936);
and U29463 (N_29463,N_21023,N_24009);
xor U29464 (N_29464,N_23797,N_20095);
or U29465 (N_29465,N_21861,N_22818);
nand U29466 (N_29466,N_20098,N_23012);
and U29467 (N_29467,N_21521,N_20828);
and U29468 (N_29468,N_22055,N_22389);
or U29469 (N_29469,N_24617,N_20946);
xor U29470 (N_29470,N_23197,N_24996);
nand U29471 (N_29471,N_22066,N_22685);
and U29472 (N_29472,N_24943,N_24248);
or U29473 (N_29473,N_22875,N_24609);
nand U29474 (N_29474,N_22211,N_23202);
xor U29475 (N_29475,N_21900,N_23132);
nor U29476 (N_29476,N_20877,N_20251);
xnor U29477 (N_29477,N_21671,N_21446);
nand U29478 (N_29478,N_20506,N_23674);
xnor U29479 (N_29479,N_20605,N_23800);
nor U29480 (N_29480,N_22856,N_23028);
nor U29481 (N_29481,N_20687,N_23203);
or U29482 (N_29482,N_24177,N_23131);
nor U29483 (N_29483,N_21027,N_23410);
and U29484 (N_29484,N_20716,N_23763);
or U29485 (N_29485,N_20908,N_21605);
nor U29486 (N_29486,N_22205,N_22017);
xnor U29487 (N_29487,N_21321,N_24662);
nand U29488 (N_29488,N_20847,N_23258);
or U29489 (N_29489,N_20298,N_24996);
xor U29490 (N_29490,N_24559,N_22702);
xnor U29491 (N_29491,N_24364,N_24887);
nor U29492 (N_29492,N_23608,N_20529);
nand U29493 (N_29493,N_24413,N_22033);
and U29494 (N_29494,N_21401,N_22395);
and U29495 (N_29495,N_24747,N_24119);
and U29496 (N_29496,N_20908,N_22522);
nor U29497 (N_29497,N_20032,N_21111);
nor U29498 (N_29498,N_23737,N_22338);
xnor U29499 (N_29499,N_23086,N_24921);
or U29500 (N_29500,N_22994,N_23496);
nor U29501 (N_29501,N_23399,N_23787);
or U29502 (N_29502,N_23486,N_20715);
and U29503 (N_29503,N_20843,N_24539);
nor U29504 (N_29504,N_22300,N_23918);
xor U29505 (N_29505,N_24695,N_21446);
nand U29506 (N_29506,N_23157,N_24858);
nor U29507 (N_29507,N_24594,N_24143);
xor U29508 (N_29508,N_24296,N_24108);
nor U29509 (N_29509,N_20700,N_21046);
or U29510 (N_29510,N_23614,N_21561);
or U29511 (N_29511,N_21822,N_22199);
and U29512 (N_29512,N_22552,N_24369);
xnor U29513 (N_29513,N_24556,N_23262);
nand U29514 (N_29514,N_24450,N_20773);
and U29515 (N_29515,N_24350,N_22533);
or U29516 (N_29516,N_23195,N_23931);
nand U29517 (N_29517,N_20508,N_24595);
nand U29518 (N_29518,N_21669,N_20234);
and U29519 (N_29519,N_21037,N_20786);
or U29520 (N_29520,N_21821,N_23441);
nor U29521 (N_29521,N_22293,N_24485);
nor U29522 (N_29522,N_24588,N_21272);
xnor U29523 (N_29523,N_22597,N_24373);
nand U29524 (N_29524,N_22335,N_20610);
nand U29525 (N_29525,N_24345,N_20256);
xor U29526 (N_29526,N_20712,N_24277);
nand U29527 (N_29527,N_22428,N_24576);
nor U29528 (N_29528,N_20357,N_22976);
nand U29529 (N_29529,N_23140,N_23681);
or U29530 (N_29530,N_21638,N_20365);
xnor U29531 (N_29531,N_24866,N_23850);
nor U29532 (N_29532,N_24036,N_20598);
xnor U29533 (N_29533,N_21835,N_22413);
and U29534 (N_29534,N_24202,N_24480);
and U29535 (N_29535,N_21646,N_23183);
nor U29536 (N_29536,N_22477,N_21667);
xnor U29537 (N_29537,N_20938,N_20112);
and U29538 (N_29538,N_22705,N_21326);
nor U29539 (N_29539,N_24194,N_24574);
nand U29540 (N_29540,N_20716,N_20200);
or U29541 (N_29541,N_24540,N_24750);
or U29542 (N_29542,N_20755,N_20489);
nand U29543 (N_29543,N_21610,N_20989);
nand U29544 (N_29544,N_22036,N_23959);
and U29545 (N_29545,N_22796,N_21691);
nor U29546 (N_29546,N_22909,N_24883);
xnor U29547 (N_29547,N_20023,N_21490);
nand U29548 (N_29548,N_22406,N_20664);
or U29549 (N_29549,N_23983,N_23611);
nor U29550 (N_29550,N_23517,N_24135);
xor U29551 (N_29551,N_22449,N_22414);
nor U29552 (N_29552,N_20021,N_24598);
xor U29553 (N_29553,N_23983,N_22439);
xor U29554 (N_29554,N_21796,N_22413);
or U29555 (N_29555,N_21855,N_21035);
or U29556 (N_29556,N_20710,N_20574);
nor U29557 (N_29557,N_21426,N_23962);
or U29558 (N_29558,N_23131,N_23005);
xor U29559 (N_29559,N_20564,N_24292);
or U29560 (N_29560,N_23335,N_22814);
and U29561 (N_29561,N_23099,N_20499);
xor U29562 (N_29562,N_23672,N_21708);
xor U29563 (N_29563,N_20619,N_23853);
or U29564 (N_29564,N_24119,N_22986);
xor U29565 (N_29565,N_24948,N_24601);
xor U29566 (N_29566,N_20514,N_22531);
and U29567 (N_29567,N_20043,N_21866);
and U29568 (N_29568,N_21463,N_24920);
and U29569 (N_29569,N_20709,N_21913);
xor U29570 (N_29570,N_21533,N_23754);
nor U29571 (N_29571,N_22916,N_20163);
nor U29572 (N_29572,N_24666,N_23830);
xor U29573 (N_29573,N_22269,N_22285);
nand U29574 (N_29574,N_24525,N_20185);
nand U29575 (N_29575,N_24928,N_22563);
nor U29576 (N_29576,N_21416,N_24075);
nand U29577 (N_29577,N_23823,N_20394);
nor U29578 (N_29578,N_21680,N_22498);
nand U29579 (N_29579,N_24955,N_20006);
and U29580 (N_29580,N_22704,N_22880);
or U29581 (N_29581,N_23960,N_20303);
xnor U29582 (N_29582,N_22507,N_22968);
nand U29583 (N_29583,N_24616,N_22518);
nand U29584 (N_29584,N_20854,N_24384);
nor U29585 (N_29585,N_20661,N_20477);
xor U29586 (N_29586,N_20993,N_20005);
and U29587 (N_29587,N_21569,N_21803);
nor U29588 (N_29588,N_24167,N_24709);
nand U29589 (N_29589,N_21173,N_24937);
nor U29590 (N_29590,N_20045,N_20359);
xnor U29591 (N_29591,N_22557,N_24024);
nor U29592 (N_29592,N_24292,N_23541);
xor U29593 (N_29593,N_20941,N_20557);
xnor U29594 (N_29594,N_23352,N_24692);
xor U29595 (N_29595,N_24569,N_23225);
nand U29596 (N_29596,N_21605,N_22872);
nand U29597 (N_29597,N_24157,N_22478);
or U29598 (N_29598,N_22223,N_21403);
nor U29599 (N_29599,N_20275,N_22534);
or U29600 (N_29600,N_23467,N_20508);
nand U29601 (N_29601,N_21745,N_20164);
xor U29602 (N_29602,N_23538,N_22297);
and U29603 (N_29603,N_20257,N_20566);
xor U29604 (N_29604,N_22196,N_23806);
and U29605 (N_29605,N_21054,N_22708);
and U29606 (N_29606,N_24705,N_24198);
nor U29607 (N_29607,N_22921,N_24532);
xor U29608 (N_29608,N_23388,N_24158);
and U29609 (N_29609,N_23929,N_22720);
nor U29610 (N_29610,N_22928,N_22795);
nand U29611 (N_29611,N_24007,N_21930);
xor U29612 (N_29612,N_20780,N_23431);
xor U29613 (N_29613,N_20505,N_24881);
xor U29614 (N_29614,N_24472,N_23503);
nor U29615 (N_29615,N_21949,N_22185);
nand U29616 (N_29616,N_23630,N_23741);
nor U29617 (N_29617,N_24862,N_20184);
nand U29618 (N_29618,N_20700,N_23988);
or U29619 (N_29619,N_23875,N_20344);
xnor U29620 (N_29620,N_23885,N_22479);
nor U29621 (N_29621,N_22179,N_23975);
or U29622 (N_29622,N_24048,N_22909);
and U29623 (N_29623,N_22026,N_23284);
or U29624 (N_29624,N_20809,N_21091);
xnor U29625 (N_29625,N_24094,N_20626);
nor U29626 (N_29626,N_23541,N_24249);
or U29627 (N_29627,N_21395,N_24712);
and U29628 (N_29628,N_21922,N_21545);
and U29629 (N_29629,N_22792,N_21969);
nand U29630 (N_29630,N_20308,N_21469);
or U29631 (N_29631,N_22107,N_22599);
nand U29632 (N_29632,N_20583,N_24216);
nand U29633 (N_29633,N_21946,N_20366);
nand U29634 (N_29634,N_20600,N_20470);
and U29635 (N_29635,N_23413,N_20989);
xor U29636 (N_29636,N_21132,N_23607);
and U29637 (N_29637,N_21359,N_20372);
and U29638 (N_29638,N_23080,N_21657);
and U29639 (N_29639,N_21205,N_24771);
and U29640 (N_29640,N_21574,N_24848);
nand U29641 (N_29641,N_20686,N_22332);
or U29642 (N_29642,N_20376,N_20651);
or U29643 (N_29643,N_22828,N_20009);
xor U29644 (N_29644,N_22324,N_24724);
nand U29645 (N_29645,N_24012,N_24324);
or U29646 (N_29646,N_20745,N_23045);
nor U29647 (N_29647,N_20782,N_20101);
nand U29648 (N_29648,N_23281,N_20241);
xor U29649 (N_29649,N_21669,N_20724);
xor U29650 (N_29650,N_20903,N_22993);
xnor U29651 (N_29651,N_21834,N_20300);
xnor U29652 (N_29652,N_22255,N_24362);
and U29653 (N_29653,N_21558,N_23446);
or U29654 (N_29654,N_21166,N_20742);
or U29655 (N_29655,N_23602,N_22762);
nor U29656 (N_29656,N_21983,N_22028);
xnor U29657 (N_29657,N_21449,N_20906);
xor U29658 (N_29658,N_24318,N_24202);
xnor U29659 (N_29659,N_21384,N_24364);
and U29660 (N_29660,N_24737,N_20249);
and U29661 (N_29661,N_21420,N_24150);
and U29662 (N_29662,N_21380,N_21061);
xor U29663 (N_29663,N_24789,N_20025);
xor U29664 (N_29664,N_20398,N_20547);
and U29665 (N_29665,N_23844,N_24443);
nand U29666 (N_29666,N_21069,N_20715);
or U29667 (N_29667,N_21842,N_23305);
xnor U29668 (N_29668,N_21914,N_21954);
or U29669 (N_29669,N_23661,N_24716);
or U29670 (N_29670,N_23108,N_22604);
nand U29671 (N_29671,N_23565,N_21633);
nor U29672 (N_29672,N_21403,N_20239);
nor U29673 (N_29673,N_22690,N_20544);
and U29674 (N_29674,N_20864,N_20596);
or U29675 (N_29675,N_20202,N_21138);
nor U29676 (N_29676,N_21326,N_21347);
and U29677 (N_29677,N_20367,N_24321);
xnor U29678 (N_29678,N_23703,N_24162);
nand U29679 (N_29679,N_20148,N_24170);
nor U29680 (N_29680,N_20832,N_23120);
nand U29681 (N_29681,N_24140,N_20654);
xnor U29682 (N_29682,N_24848,N_21984);
nor U29683 (N_29683,N_22810,N_21080);
nor U29684 (N_29684,N_24855,N_21406);
xnor U29685 (N_29685,N_23012,N_21363);
nor U29686 (N_29686,N_24125,N_23271);
xnor U29687 (N_29687,N_21085,N_24615);
xnor U29688 (N_29688,N_23069,N_21842);
nor U29689 (N_29689,N_20800,N_22273);
nand U29690 (N_29690,N_22966,N_23827);
xnor U29691 (N_29691,N_23424,N_23864);
xnor U29692 (N_29692,N_20327,N_21739);
or U29693 (N_29693,N_22515,N_21405);
nand U29694 (N_29694,N_20943,N_23572);
nand U29695 (N_29695,N_23857,N_24131);
or U29696 (N_29696,N_21213,N_23599);
or U29697 (N_29697,N_24053,N_24550);
xor U29698 (N_29698,N_23678,N_23545);
nand U29699 (N_29699,N_23654,N_21646);
or U29700 (N_29700,N_20133,N_24528);
nand U29701 (N_29701,N_20855,N_22731);
nor U29702 (N_29702,N_20267,N_20378);
and U29703 (N_29703,N_22181,N_20258);
xor U29704 (N_29704,N_23546,N_24714);
nand U29705 (N_29705,N_22240,N_21441);
nor U29706 (N_29706,N_23666,N_23159);
nor U29707 (N_29707,N_23895,N_23466);
and U29708 (N_29708,N_21441,N_23018);
nand U29709 (N_29709,N_23541,N_20680);
xnor U29710 (N_29710,N_24455,N_23126);
xnor U29711 (N_29711,N_24433,N_21034);
or U29712 (N_29712,N_21847,N_24437);
and U29713 (N_29713,N_24701,N_23978);
nor U29714 (N_29714,N_22409,N_24800);
nor U29715 (N_29715,N_21138,N_23921);
or U29716 (N_29716,N_20792,N_20674);
nor U29717 (N_29717,N_21489,N_24464);
and U29718 (N_29718,N_21475,N_22212);
nand U29719 (N_29719,N_21115,N_23278);
or U29720 (N_29720,N_24114,N_23077);
nand U29721 (N_29721,N_24897,N_24600);
and U29722 (N_29722,N_21387,N_21364);
or U29723 (N_29723,N_23680,N_21277);
or U29724 (N_29724,N_20456,N_22318);
xnor U29725 (N_29725,N_21872,N_24500);
nor U29726 (N_29726,N_20910,N_24106);
and U29727 (N_29727,N_24320,N_21550);
or U29728 (N_29728,N_22414,N_23179);
nand U29729 (N_29729,N_22434,N_21027);
nand U29730 (N_29730,N_20658,N_23275);
nand U29731 (N_29731,N_22067,N_22840);
nor U29732 (N_29732,N_22779,N_23591);
nor U29733 (N_29733,N_23690,N_20720);
nor U29734 (N_29734,N_23776,N_21912);
xnor U29735 (N_29735,N_24057,N_20522);
nand U29736 (N_29736,N_23881,N_23084);
nand U29737 (N_29737,N_21821,N_20488);
or U29738 (N_29738,N_21649,N_20384);
and U29739 (N_29739,N_23427,N_22085);
nand U29740 (N_29740,N_20658,N_24910);
or U29741 (N_29741,N_22223,N_21581);
nor U29742 (N_29742,N_21670,N_20887);
or U29743 (N_29743,N_22298,N_23852);
nand U29744 (N_29744,N_21666,N_21070);
xor U29745 (N_29745,N_20461,N_22508);
xor U29746 (N_29746,N_20348,N_24054);
or U29747 (N_29747,N_24131,N_20403);
nor U29748 (N_29748,N_23862,N_24971);
or U29749 (N_29749,N_23877,N_21411);
or U29750 (N_29750,N_20904,N_20311);
nand U29751 (N_29751,N_21513,N_20588);
xor U29752 (N_29752,N_24708,N_20521);
xor U29753 (N_29753,N_23633,N_24866);
or U29754 (N_29754,N_23785,N_21435);
nor U29755 (N_29755,N_24902,N_22366);
nor U29756 (N_29756,N_21070,N_24787);
xor U29757 (N_29757,N_23577,N_23812);
nor U29758 (N_29758,N_20372,N_24388);
xnor U29759 (N_29759,N_20411,N_24623);
nor U29760 (N_29760,N_24054,N_24297);
nor U29761 (N_29761,N_23743,N_24067);
and U29762 (N_29762,N_23620,N_24977);
or U29763 (N_29763,N_20759,N_20546);
nor U29764 (N_29764,N_21354,N_24606);
xor U29765 (N_29765,N_22599,N_23319);
nand U29766 (N_29766,N_21215,N_24799);
xnor U29767 (N_29767,N_23715,N_20096);
or U29768 (N_29768,N_23937,N_24658);
nand U29769 (N_29769,N_22540,N_23085);
and U29770 (N_29770,N_23245,N_22178);
xor U29771 (N_29771,N_23520,N_21005);
nor U29772 (N_29772,N_23600,N_21243);
nand U29773 (N_29773,N_21856,N_21081);
xnor U29774 (N_29774,N_20596,N_23251);
xnor U29775 (N_29775,N_20032,N_21467);
xnor U29776 (N_29776,N_24093,N_21654);
and U29777 (N_29777,N_22191,N_23290);
nor U29778 (N_29778,N_21839,N_22156);
or U29779 (N_29779,N_22666,N_24886);
and U29780 (N_29780,N_24333,N_20702);
or U29781 (N_29781,N_21081,N_24488);
and U29782 (N_29782,N_23043,N_22676);
or U29783 (N_29783,N_21662,N_20354);
nand U29784 (N_29784,N_20584,N_22113);
nor U29785 (N_29785,N_24121,N_24463);
nand U29786 (N_29786,N_21047,N_23430);
and U29787 (N_29787,N_22176,N_21332);
nor U29788 (N_29788,N_20390,N_23752);
nor U29789 (N_29789,N_20159,N_23811);
or U29790 (N_29790,N_24060,N_21235);
nor U29791 (N_29791,N_24850,N_21463);
nor U29792 (N_29792,N_20280,N_24714);
and U29793 (N_29793,N_20028,N_21837);
or U29794 (N_29794,N_21507,N_21222);
xnor U29795 (N_29795,N_20040,N_22204);
and U29796 (N_29796,N_23943,N_23877);
nor U29797 (N_29797,N_20427,N_20925);
and U29798 (N_29798,N_21662,N_20297);
or U29799 (N_29799,N_23095,N_24053);
nand U29800 (N_29800,N_22685,N_21742);
nor U29801 (N_29801,N_20456,N_23044);
or U29802 (N_29802,N_24020,N_24690);
nor U29803 (N_29803,N_23955,N_22340);
nand U29804 (N_29804,N_24578,N_23773);
or U29805 (N_29805,N_24686,N_21781);
or U29806 (N_29806,N_21164,N_20849);
nand U29807 (N_29807,N_24435,N_20121);
and U29808 (N_29808,N_21257,N_20352);
nand U29809 (N_29809,N_22884,N_24071);
nand U29810 (N_29810,N_20878,N_21964);
xnor U29811 (N_29811,N_20704,N_20248);
or U29812 (N_29812,N_20993,N_23168);
xor U29813 (N_29813,N_24377,N_24470);
nor U29814 (N_29814,N_20361,N_22906);
or U29815 (N_29815,N_24107,N_22618);
xor U29816 (N_29816,N_23478,N_22407);
nand U29817 (N_29817,N_22145,N_20558);
or U29818 (N_29818,N_23386,N_24970);
or U29819 (N_29819,N_21337,N_20524);
nand U29820 (N_29820,N_23907,N_20636);
xnor U29821 (N_29821,N_23271,N_21231);
nor U29822 (N_29822,N_22802,N_20978);
nor U29823 (N_29823,N_22945,N_23339);
nand U29824 (N_29824,N_20380,N_23892);
and U29825 (N_29825,N_20940,N_23933);
xnor U29826 (N_29826,N_22644,N_23207);
and U29827 (N_29827,N_23868,N_24335);
nor U29828 (N_29828,N_21059,N_22221);
and U29829 (N_29829,N_23564,N_21817);
nor U29830 (N_29830,N_22376,N_24192);
nand U29831 (N_29831,N_22050,N_21353);
xnor U29832 (N_29832,N_22916,N_22535);
or U29833 (N_29833,N_24832,N_20180);
and U29834 (N_29834,N_23012,N_22211);
and U29835 (N_29835,N_20390,N_23135);
xnor U29836 (N_29836,N_20898,N_24224);
xor U29837 (N_29837,N_21136,N_21107);
xnor U29838 (N_29838,N_23847,N_22110);
xor U29839 (N_29839,N_21976,N_22259);
or U29840 (N_29840,N_22791,N_21841);
and U29841 (N_29841,N_24669,N_21256);
nand U29842 (N_29842,N_21432,N_24274);
nand U29843 (N_29843,N_20109,N_22839);
nor U29844 (N_29844,N_24282,N_23438);
or U29845 (N_29845,N_21753,N_24621);
or U29846 (N_29846,N_23542,N_22314);
and U29847 (N_29847,N_21763,N_22076);
or U29848 (N_29848,N_20876,N_20480);
nor U29849 (N_29849,N_22040,N_22818);
or U29850 (N_29850,N_23536,N_21411);
nor U29851 (N_29851,N_21144,N_23991);
or U29852 (N_29852,N_22562,N_20685);
nand U29853 (N_29853,N_21626,N_23436);
and U29854 (N_29854,N_24012,N_20181);
or U29855 (N_29855,N_24669,N_22821);
xnor U29856 (N_29856,N_20177,N_24180);
xnor U29857 (N_29857,N_23429,N_22551);
nor U29858 (N_29858,N_22098,N_23912);
nor U29859 (N_29859,N_22057,N_20311);
nand U29860 (N_29860,N_22628,N_21634);
nor U29861 (N_29861,N_22810,N_24346);
nor U29862 (N_29862,N_22316,N_24418);
nor U29863 (N_29863,N_20577,N_20993);
nand U29864 (N_29864,N_24557,N_21604);
xnor U29865 (N_29865,N_23840,N_23310);
or U29866 (N_29866,N_22838,N_24036);
xor U29867 (N_29867,N_22137,N_21931);
nor U29868 (N_29868,N_22378,N_22229);
or U29869 (N_29869,N_24837,N_21162);
or U29870 (N_29870,N_22600,N_22627);
nor U29871 (N_29871,N_22388,N_22544);
nand U29872 (N_29872,N_21738,N_23605);
or U29873 (N_29873,N_22150,N_21147);
or U29874 (N_29874,N_21893,N_20811);
or U29875 (N_29875,N_21469,N_24884);
and U29876 (N_29876,N_20483,N_21929);
nand U29877 (N_29877,N_23653,N_20232);
or U29878 (N_29878,N_21282,N_22148);
xnor U29879 (N_29879,N_24163,N_20703);
nor U29880 (N_29880,N_20830,N_20761);
nand U29881 (N_29881,N_22586,N_20095);
and U29882 (N_29882,N_20228,N_20270);
xor U29883 (N_29883,N_24987,N_22631);
nand U29884 (N_29884,N_21751,N_21293);
or U29885 (N_29885,N_20601,N_22681);
or U29886 (N_29886,N_21335,N_22207);
or U29887 (N_29887,N_22585,N_23296);
nor U29888 (N_29888,N_23241,N_24288);
xnor U29889 (N_29889,N_20375,N_24885);
xnor U29890 (N_29890,N_20728,N_24730);
nand U29891 (N_29891,N_24190,N_24132);
xnor U29892 (N_29892,N_23482,N_21133);
nor U29893 (N_29893,N_21160,N_22328);
xor U29894 (N_29894,N_22562,N_20834);
or U29895 (N_29895,N_21837,N_21979);
nor U29896 (N_29896,N_23285,N_21148);
nand U29897 (N_29897,N_21505,N_23360);
xnor U29898 (N_29898,N_23056,N_22179);
xnor U29899 (N_29899,N_22123,N_20430);
nor U29900 (N_29900,N_21629,N_22781);
nor U29901 (N_29901,N_23055,N_20036);
nor U29902 (N_29902,N_21239,N_24546);
xnor U29903 (N_29903,N_21370,N_22611);
and U29904 (N_29904,N_22569,N_23938);
or U29905 (N_29905,N_20130,N_22372);
nand U29906 (N_29906,N_22262,N_21309);
xnor U29907 (N_29907,N_24122,N_20379);
or U29908 (N_29908,N_20851,N_23478);
xnor U29909 (N_29909,N_20067,N_24620);
nand U29910 (N_29910,N_23321,N_24188);
xor U29911 (N_29911,N_21371,N_23529);
nand U29912 (N_29912,N_21363,N_24884);
xnor U29913 (N_29913,N_21653,N_21179);
nor U29914 (N_29914,N_22579,N_21215);
nor U29915 (N_29915,N_22293,N_21726);
nand U29916 (N_29916,N_24136,N_23421);
or U29917 (N_29917,N_23660,N_21373);
and U29918 (N_29918,N_22735,N_23646);
nor U29919 (N_29919,N_23711,N_23277);
and U29920 (N_29920,N_22318,N_20813);
nand U29921 (N_29921,N_22979,N_21042);
and U29922 (N_29922,N_24869,N_23878);
or U29923 (N_29923,N_23292,N_20697);
xnor U29924 (N_29924,N_23393,N_22706);
nor U29925 (N_29925,N_24772,N_22357);
or U29926 (N_29926,N_21043,N_20126);
or U29927 (N_29927,N_23059,N_23116);
and U29928 (N_29928,N_21558,N_23501);
nor U29929 (N_29929,N_20944,N_24014);
or U29930 (N_29930,N_21194,N_20091);
nand U29931 (N_29931,N_22197,N_23725);
nand U29932 (N_29932,N_20862,N_20540);
and U29933 (N_29933,N_23566,N_23629);
nor U29934 (N_29934,N_22483,N_21475);
xor U29935 (N_29935,N_24165,N_22698);
or U29936 (N_29936,N_23885,N_21444);
nand U29937 (N_29937,N_20111,N_21697);
and U29938 (N_29938,N_20170,N_23002);
nand U29939 (N_29939,N_22927,N_23920);
nand U29940 (N_29940,N_21514,N_24678);
or U29941 (N_29941,N_20337,N_24968);
nor U29942 (N_29942,N_22781,N_22786);
and U29943 (N_29943,N_22541,N_21191);
or U29944 (N_29944,N_20456,N_20124);
or U29945 (N_29945,N_24333,N_20556);
and U29946 (N_29946,N_23003,N_20550);
or U29947 (N_29947,N_24330,N_24345);
or U29948 (N_29948,N_20239,N_23325);
or U29949 (N_29949,N_20374,N_24242);
and U29950 (N_29950,N_22766,N_24440);
nor U29951 (N_29951,N_24991,N_20200);
xnor U29952 (N_29952,N_21252,N_21260);
and U29953 (N_29953,N_21996,N_24501);
xnor U29954 (N_29954,N_21667,N_21622);
nand U29955 (N_29955,N_20733,N_21191);
nor U29956 (N_29956,N_23919,N_20099);
nand U29957 (N_29957,N_21548,N_23678);
nand U29958 (N_29958,N_24523,N_20044);
nor U29959 (N_29959,N_23558,N_21086);
xor U29960 (N_29960,N_22508,N_23465);
xor U29961 (N_29961,N_21465,N_21073);
nor U29962 (N_29962,N_24891,N_23460);
nor U29963 (N_29963,N_23262,N_20720);
xnor U29964 (N_29964,N_23598,N_20139);
nand U29965 (N_29965,N_22323,N_23681);
nor U29966 (N_29966,N_22273,N_20844);
or U29967 (N_29967,N_21006,N_24280);
nand U29968 (N_29968,N_23924,N_24548);
or U29969 (N_29969,N_23203,N_20449);
xnor U29970 (N_29970,N_20613,N_24177);
xnor U29971 (N_29971,N_22932,N_22510);
nand U29972 (N_29972,N_20799,N_24119);
xor U29973 (N_29973,N_21958,N_21770);
and U29974 (N_29974,N_22826,N_23884);
xnor U29975 (N_29975,N_22233,N_20353);
or U29976 (N_29976,N_22781,N_20887);
xnor U29977 (N_29977,N_21905,N_23296);
and U29978 (N_29978,N_23043,N_24005);
nor U29979 (N_29979,N_24519,N_22935);
nor U29980 (N_29980,N_24345,N_23399);
xor U29981 (N_29981,N_21662,N_22982);
nor U29982 (N_29982,N_23133,N_20980);
and U29983 (N_29983,N_21005,N_22232);
nor U29984 (N_29984,N_24204,N_20744);
and U29985 (N_29985,N_22389,N_21344);
and U29986 (N_29986,N_22879,N_22615);
or U29987 (N_29987,N_20252,N_22948);
nand U29988 (N_29988,N_24961,N_22335);
and U29989 (N_29989,N_22598,N_24541);
and U29990 (N_29990,N_21990,N_24488);
nor U29991 (N_29991,N_20654,N_21206);
xor U29992 (N_29992,N_21398,N_21737);
or U29993 (N_29993,N_23696,N_20812);
and U29994 (N_29994,N_21067,N_20630);
or U29995 (N_29995,N_23921,N_23971);
or U29996 (N_29996,N_24544,N_23075);
or U29997 (N_29997,N_20836,N_20801);
or U29998 (N_29998,N_23302,N_24861);
or U29999 (N_29999,N_22462,N_20709);
xnor U30000 (N_30000,N_25777,N_28661);
or U30001 (N_30001,N_29462,N_29327);
xnor U30002 (N_30002,N_25700,N_27095);
xor U30003 (N_30003,N_29384,N_29207);
and U30004 (N_30004,N_25229,N_27894);
nor U30005 (N_30005,N_27043,N_28724);
nor U30006 (N_30006,N_27534,N_26388);
and U30007 (N_30007,N_25952,N_28726);
and U30008 (N_30008,N_29668,N_25606);
nor U30009 (N_30009,N_25261,N_27411);
and U30010 (N_30010,N_29536,N_29979);
xor U30011 (N_30011,N_25825,N_29538);
nor U30012 (N_30012,N_25356,N_28597);
nand U30013 (N_30013,N_29801,N_28966);
or U30014 (N_30014,N_27319,N_29274);
and U30015 (N_30015,N_28808,N_27333);
or U30016 (N_30016,N_29928,N_26837);
nor U30017 (N_30017,N_29755,N_26827);
nand U30018 (N_30018,N_28954,N_29263);
xnor U30019 (N_30019,N_29751,N_26328);
or U30020 (N_30020,N_26230,N_27617);
xnor U30021 (N_30021,N_29276,N_25631);
nand U30022 (N_30022,N_27941,N_26899);
nand U30023 (N_30023,N_29165,N_29865);
and U30024 (N_30024,N_29839,N_26864);
or U30025 (N_30025,N_27010,N_29267);
or U30026 (N_30026,N_28865,N_25774);
xor U30027 (N_30027,N_28589,N_28314);
nand U30028 (N_30028,N_29265,N_27834);
nand U30029 (N_30029,N_25466,N_29308);
xnor U30030 (N_30030,N_26287,N_25561);
or U30031 (N_30031,N_27357,N_28605);
xor U30032 (N_30032,N_27205,N_25255);
nor U30033 (N_30033,N_25844,N_28557);
and U30034 (N_30034,N_26194,N_27315);
nand U30035 (N_30035,N_27803,N_29737);
or U30036 (N_30036,N_29437,N_28941);
and U30037 (N_30037,N_27076,N_25820);
and U30038 (N_30038,N_28623,N_26763);
or U30039 (N_30039,N_27830,N_26876);
and U30040 (N_30040,N_25563,N_27732);
nor U30041 (N_30041,N_27512,N_29799);
or U30042 (N_30042,N_27546,N_25724);
nor U30043 (N_30043,N_28218,N_27037);
or U30044 (N_30044,N_26882,N_27194);
xor U30045 (N_30045,N_25522,N_25436);
nor U30046 (N_30046,N_25891,N_25908);
nor U30047 (N_30047,N_29466,N_25664);
and U30048 (N_30048,N_26771,N_29117);
xor U30049 (N_30049,N_27906,N_26814);
nor U30050 (N_30050,N_25934,N_29168);
and U30051 (N_30051,N_27405,N_28626);
and U30052 (N_30052,N_28430,N_25000);
nor U30053 (N_30053,N_29102,N_25787);
xor U30054 (N_30054,N_29515,N_26874);
or U30055 (N_30055,N_29337,N_26207);
xnor U30056 (N_30056,N_26891,N_26791);
nor U30057 (N_30057,N_29509,N_27460);
xnor U30058 (N_30058,N_29348,N_28097);
or U30059 (N_30059,N_28518,N_27925);
and U30060 (N_30060,N_28801,N_25176);
and U30061 (N_30061,N_29615,N_29461);
nand U30062 (N_30062,N_26485,N_27932);
nand U30063 (N_30063,N_29224,N_29100);
nor U30064 (N_30064,N_28025,N_25720);
nor U30065 (N_30065,N_28447,N_27792);
or U30066 (N_30066,N_28418,N_27376);
nand U30067 (N_30067,N_28442,N_26175);
xor U30068 (N_30068,N_25275,N_25299);
and U30069 (N_30069,N_28168,N_27623);
xnor U30070 (N_30070,N_26359,N_29763);
nor U30071 (N_30071,N_29077,N_25168);
nand U30072 (N_30072,N_25317,N_29858);
nand U30073 (N_30073,N_29873,N_27047);
xor U30074 (N_30074,N_29387,N_25003);
and U30075 (N_30075,N_28863,N_26753);
nor U30076 (N_30076,N_28743,N_26502);
or U30077 (N_30077,N_27438,N_27624);
nor U30078 (N_30078,N_26866,N_26020);
and U30079 (N_30079,N_29402,N_27400);
and U30080 (N_30080,N_26664,N_28227);
and U30081 (N_30081,N_27498,N_29085);
or U30082 (N_30082,N_28343,N_28551);
nand U30083 (N_30083,N_28593,N_28830);
or U30084 (N_30084,N_27513,N_26167);
and U30085 (N_30085,N_26636,N_27694);
nor U30086 (N_30086,N_26657,N_25671);
and U30087 (N_30087,N_29345,N_25349);
xor U30088 (N_30088,N_25185,N_29604);
nor U30089 (N_30089,N_28038,N_27998);
nor U30090 (N_30090,N_26021,N_26695);
or U30091 (N_30091,N_28531,N_27589);
xnor U30092 (N_30092,N_29579,N_28262);
or U30093 (N_30093,N_27819,N_28364);
xnor U30094 (N_30094,N_27297,N_27298);
or U30095 (N_30095,N_27256,N_28750);
nand U30096 (N_30096,N_28883,N_27207);
nand U30097 (N_30097,N_25867,N_28799);
and U30098 (N_30098,N_25402,N_25604);
xnor U30099 (N_30099,N_28056,N_26419);
or U30100 (N_30100,N_27280,N_29380);
and U30101 (N_30101,N_29527,N_29614);
nor U30102 (N_30102,N_27358,N_25854);
or U30103 (N_30103,N_25348,N_29496);
nor U30104 (N_30104,N_28765,N_27288);
nor U30105 (N_30105,N_29225,N_29699);
xor U30106 (N_30106,N_28760,N_28127);
nand U30107 (N_30107,N_29857,N_25379);
or U30108 (N_30108,N_28712,N_25374);
nand U30109 (N_30109,N_27885,N_26652);
xnor U30110 (N_30110,N_26555,N_26023);
xnor U30111 (N_30111,N_26311,N_27011);
nor U30112 (N_30112,N_25068,N_28681);
nand U30113 (N_30113,N_26660,N_26093);
or U30114 (N_30114,N_28394,N_25605);
xor U30115 (N_30115,N_25884,N_29130);
nand U30116 (N_30116,N_29004,N_28942);
nor U30117 (N_30117,N_26169,N_28274);
or U30118 (N_30118,N_28031,N_25096);
and U30119 (N_30119,N_29269,N_27106);
xnor U30120 (N_30120,N_26514,N_25449);
nand U30121 (N_30121,N_26275,N_27214);
nor U30122 (N_30122,N_27223,N_28142);
nand U30123 (N_30123,N_27957,N_28854);
nor U30124 (N_30124,N_27414,N_25084);
or U30125 (N_30125,N_28202,N_26966);
nor U30126 (N_30126,N_28848,N_26599);
nor U30127 (N_30127,N_26844,N_25417);
and U30128 (N_30128,N_27377,N_28028);
nand U30129 (N_30129,N_26812,N_26310);
nand U30130 (N_30130,N_27407,N_25395);
or U30131 (N_30131,N_27350,N_29984);
xnor U30132 (N_30132,N_27691,N_27616);
nand U30133 (N_30133,N_29322,N_25221);
or U30134 (N_30134,N_29576,N_26174);
or U30135 (N_30135,N_28466,N_27329);
nand U30136 (N_30136,N_25918,N_26649);
nand U30137 (N_30137,N_27393,N_28565);
nand U30138 (N_30138,N_27439,N_28018);
and U30139 (N_30139,N_28894,N_26718);
and U30140 (N_30140,N_26561,N_26339);
or U30141 (N_30141,N_26639,N_29342);
and U30142 (N_30142,N_29143,N_27591);
or U30143 (N_30143,N_28363,N_27521);
and U30144 (N_30144,N_29864,N_26429);
nand U30145 (N_30145,N_29415,N_25656);
nor U30146 (N_30146,N_26984,N_27192);
nand U30147 (N_30147,N_27781,N_28051);
nand U30148 (N_30148,N_25063,N_25476);
nand U30149 (N_30149,N_27917,N_26115);
nand U30150 (N_30150,N_28833,N_28767);
and U30151 (N_30151,N_29052,N_25640);
xnor U30152 (N_30152,N_28437,N_27689);
nand U30153 (N_30153,N_26210,N_27481);
or U30154 (N_30154,N_29053,N_27212);
and U30155 (N_30155,N_26790,N_25070);
xnor U30156 (N_30156,N_28775,N_28369);
nor U30157 (N_30157,N_27286,N_29486);
and U30158 (N_30158,N_27155,N_25312);
nand U30159 (N_30159,N_28293,N_26831);
or U30160 (N_30160,N_29757,N_27867);
nor U30161 (N_30161,N_26407,N_29567);
or U30162 (N_30162,N_25965,N_29043);
or U30163 (N_30163,N_27502,N_27126);
and U30164 (N_30164,N_25623,N_29317);
and U30165 (N_30165,N_28719,N_28371);
xor U30166 (N_30166,N_26982,N_28278);
nor U30167 (N_30167,N_27361,N_27662);
and U30168 (N_30168,N_28332,N_27324);
nor U30169 (N_30169,N_29859,N_29927);
nor U30170 (N_30170,N_28123,N_28326);
nand U30171 (N_30171,N_27704,N_28609);
and U30172 (N_30172,N_28501,N_25574);
or U30173 (N_30173,N_27908,N_25400);
nor U30174 (N_30174,N_26289,N_26838);
or U30175 (N_30175,N_27699,N_26641);
nor U30176 (N_30176,N_25532,N_27461);
nor U30177 (N_30177,N_29047,N_28581);
nor U30178 (N_30178,N_26687,N_26968);
or U30179 (N_30179,N_28819,N_25986);
xor U30180 (N_30180,N_25154,N_26246);
xnor U30181 (N_30181,N_27038,N_28722);
xor U30182 (N_30182,N_27654,N_27339);
nor U30183 (N_30183,N_27936,N_29103);
or U30184 (N_30184,N_28720,N_29075);
nor U30185 (N_30185,N_29718,N_26049);
nand U30186 (N_30186,N_25558,N_25830);
and U30187 (N_30187,N_25383,N_29151);
and U30188 (N_30188,N_26694,N_25872);
and U30189 (N_30189,N_28292,N_29273);
xnor U30190 (N_30190,N_29526,N_27462);
xnor U30191 (N_30191,N_29012,N_28596);
nand U30192 (N_30192,N_27167,N_27557);
and U30193 (N_30193,N_26726,N_25603);
nand U30194 (N_30194,N_28105,N_25839);
nand U30195 (N_30195,N_29157,N_26281);
or U30196 (N_30196,N_28417,N_25242);
nand U30197 (N_30197,N_27531,N_28246);
or U30198 (N_30198,N_28185,N_29350);
nand U30199 (N_30199,N_25899,N_25688);
and U30200 (N_30200,N_26821,N_28617);
nand U30201 (N_30201,N_26819,N_29636);
nand U30202 (N_30202,N_25060,N_26676);
nand U30203 (N_30203,N_29943,N_28256);
and U30204 (N_30204,N_28691,N_27943);
nor U30205 (N_30205,N_25314,N_25005);
nor U30206 (N_30206,N_26393,N_26160);
xnor U30207 (N_30207,N_27385,N_27950);
and U30208 (N_30208,N_29769,N_26408);
and U30209 (N_30209,N_25306,N_28996);
nor U30210 (N_30210,N_28555,N_26569);
and U30211 (N_30211,N_27570,N_26648);
and U30212 (N_30212,N_26209,N_29236);
nor U30213 (N_30213,N_28662,N_25661);
nand U30214 (N_30214,N_26723,N_25578);
nor U30215 (N_30215,N_27174,N_28040);
or U30216 (N_30216,N_28283,N_28853);
nand U30217 (N_30217,N_27595,N_25159);
nand U30218 (N_30218,N_26574,N_26430);
nand U30219 (N_30219,N_28825,N_28120);
nand U30220 (N_30220,N_25035,N_27535);
xor U30221 (N_30221,N_27145,N_29732);
nand U30222 (N_30222,N_26884,N_28070);
nor U30223 (N_30223,N_28360,N_28911);
xnor U30224 (N_30224,N_29639,N_29583);
nand U30225 (N_30225,N_29982,N_29907);
nor U30226 (N_30226,N_25812,N_26645);
or U30227 (N_30227,N_25619,N_27356);
xor U30228 (N_30228,N_26559,N_26143);
and U30229 (N_30229,N_27431,N_27912);
or U30230 (N_30230,N_26607,N_25556);
xnor U30231 (N_30231,N_26205,N_29280);
xnor U30232 (N_30232,N_26562,N_28382);
or U30233 (N_30233,N_25654,N_25498);
nor U30234 (N_30234,N_28378,N_26098);
or U30235 (N_30235,N_26251,N_28194);
and U30236 (N_30236,N_26589,N_27486);
or U30237 (N_30237,N_29998,N_28812);
or U30238 (N_30238,N_28098,N_28864);
and U30239 (N_30239,N_26202,N_29860);
and U30240 (N_30240,N_27711,N_25523);
and U30241 (N_30241,N_28672,N_25978);
xnor U30242 (N_30242,N_26683,N_25113);
nor U30243 (N_30243,N_26877,N_29039);
and U30244 (N_30244,N_29054,N_27232);
nor U30245 (N_30245,N_26147,N_29533);
xnor U30246 (N_30246,N_27060,N_27386);
and U30247 (N_30247,N_27284,N_29563);
nor U30248 (N_30248,N_29909,N_26266);
nor U30249 (N_30249,N_29803,N_29925);
xor U30250 (N_30250,N_28043,N_25819);
nor U30251 (N_30251,N_27861,N_28297);
and U30252 (N_30252,N_28113,N_28682);
or U30253 (N_30253,N_26799,N_28352);
or U30254 (N_30254,N_25336,N_29204);
xnor U30255 (N_30255,N_27408,N_25906);
nand U30256 (N_30256,N_29477,N_25411);
nor U30257 (N_30257,N_29036,N_27544);
nand U30258 (N_30258,N_26856,N_27345);
nand U30259 (N_30259,N_26456,N_26498);
xnor U30260 (N_30260,N_26451,N_26854);
or U30261 (N_30261,N_29712,N_26253);
or U30262 (N_30262,N_25738,N_25576);
nor U30263 (N_30263,N_27472,N_28699);
xnor U30264 (N_30264,N_26119,N_28636);
and U30265 (N_30265,N_29875,N_26046);
nor U30266 (N_30266,N_29593,N_27003);
xor U30267 (N_30267,N_25297,N_25415);
xnor U30268 (N_30268,N_26390,N_28665);
or U30269 (N_30269,N_27142,N_29890);
nor U30270 (N_30270,N_25352,N_26371);
xor U30271 (N_30271,N_25325,N_27923);
and U30272 (N_30272,N_28348,N_27731);
nand U30273 (N_30273,N_25740,N_26022);
or U30274 (N_30274,N_27419,N_29459);
and U30275 (N_30275,N_25589,N_26826);
or U30276 (N_30276,N_27208,N_25055);
or U30277 (N_30277,N_25265,N_25303);
xnor U30278 (N_30278,N_27237,N_26432);
and U30279 (N_30279,N_28616,N_27716);
xor U30280 (N_30280,N_28413,N_27177);
xor U30281 (N_30281,N_29768,N_26547);
or U30282 (N_30282,N_25246,N_28530);
nor U30283 (N_30283,N_27636,N_29715);
nor U30284 (N_30284,N_26212,N_27020);
and U30285 (N_30285,N_27480,N_28446);
xor U30286 (N_30286,N_26280,N_26531);
and U30287 (N_30287,N_25646,N_29561);
and U30288 (N_30288,N_29885,N_27353);
or U30289 (N_30289,N_28091,N_27737);
nand U30290 (N_30290,N_27575,N_28696);
nor U30291 (N_30291,N_26025,N_28154);
nand U30292 (N_30292,N_28885,N_26192);
and U30293 (N_30293,N_29167,N_29005);
or U30294 (N_30294,N_26383,N_26374);
nand U30295 (N_30295,N_28429,N_27606);
or U30296 (N_30296,N_25503,N_25858);
nor U30297 (N_30297,N_29884,N_27703);
or U30298 (N_30298,N_27226,N_26697);
or U30299 (N_30299,N_26992,N_27228);
xor U30300 (N_30300,N_28462,N_25600);
xor U30301 (N_30301,N_26235,N_25860);
nor U30302 (N_30302,N_28167,N_27227);
nand U30303 (N_30303,N_29163,N_28376);
and U30304 (N_30304,N_26001,N_27225);
or U30305 (N_30305,N_25416,N_25681);
xnor U30306 (N_30306,N_27701,N_26708);
nand U30307 (N_30307,N_29525,N_27783);
and U30308 (N_30308,N_25694,N_26646);
xor U30309 (N_30309,N_27437,N_26448);
nor U30310 (N_30310,N_25726,N_29050);
and U30311 (N_30311,N_27734,N_29571);
nand U30312 (N_30312,N_29772,N_26788);
and U30313 (N_30313,N_27264,N_26983);
nor U30314 (N_30314,N_29430,N_28008);
xnor U30315 (N_30315,N_27963,N_29046);
nor U30316 (N_30316,N_28667,N_28611);
or U30317 (N_30317,N_27257,N_29625);
nor U30318 (N_30318,N_25827,N_25288);
nor U30319 (N_30319,N_27631,N_25123);
nor U30320 (N_30320,N_29694,N_26947);
nor U30321 (N_30321,N_27960,N_27346);
and U30322 (N_30322,N_27000,N_25732);
nand U30323 (N_30323,N_25041,N_27379);
xnor U30324 (N_30324,N_29640,N_27667);
xnor U30325 (N_30325,N_27176,N_29521);
xnor U30326 (N_30326,N_25541,N_28859);
and U30327 (N_30327,N_29988,N_28355);
xor U30328 (N_30328,N_28508,N_27554);
xor U30329 (N_30329,N_27794,N_25450);
or U30330 (N_30330,N_28958,N_28540);
and U30331 (N_30331,N_29110,N_27231);
nor U30332 (N_30332,N_25057,N_27844);
and U30333 (N_30333,N_25873,N_28721);
xor U30334 (N_30334,N_27373,N_28546);
nand U30335 (N_30335,N_28368,N_28450);
or U30336 (N_30336,N_29662,N_25492);
xnor U30337 (N_30337,N_28434,N_27072);
and U30338 (N_30338,N_25911,N_26523);
nor U30339 (N_30339,N_26358,N_29968);
and U30340 (N_30340,N_25943,N_25817);
and U30341 (N_30341,N_25283,N_27249);
nor U30342 (N_30342,N_27161,N_28261);
nand U30343 (N_30343,N_25923,N_25272);
nand U30344 (N_30344,N_26997,N_29920);
nand U30345 (N_30345,N_26367,N_29433);
or U30346 (N_30346,N_27166,N_28713);
or U30347 (N_30347,N_28505,N_27395);
and U30348 (N_30348,N_27607,N_29516);
nor U30349 (N_30349,N_28993,N_25514);
nor U30350 (N_30350,N_29002,N_25669);
and U30351 (N_30351,N_29467,N_25230);
xnor U30352 (N_30352,N_28024,N_27447);
nor U30353 (N_30353,N_25678,N_27533);
xor U30354 (N_30354,N_26481,N_29631);
nor U30355 (N_30355,N_28562,N_26948);
nor U30356 (N_30356,N_27100,N_25611);
or U30357 (N_30357,N_29827,N_27418);
and U30358 (N_30358,N_29861,N_27215);
xor U30359 (N_30359,N_29196,N_26590);
and U30360 (N_30360,N_25804,N_25422);
xor U30361 (N_30361,N_25329,N_25781);
nand U30362 (N_30362,N_28519,N_26270);
or U30363 (N_30363,N_29818,N_27242);
nor U30364 (N_30364,N_26693,N_25194);
xor U30365 (N_30365,N_27629,N_27222);
or U30366 (N_30366,N_25008,N_26824);
or U30367 (N_30367,N_25107,N_29155);
or U30368 (N_30368,N_29959,N_28301);
or U30369 (N_30369,N_25291,N_29293);
and U30370 (N_30370,N_28693,N_26297);
xor U30371 (N_30371,N_29644,N_29019);
and U30372 (N_30372,N_29185,N_25213);
xor U30373 (N_30373,N_29418,N_28882);
or U30374 (N_30374,N_29993,N_25225);
or U30375 (N_30375,N_27069,N_28473);
xor U30376 (N_30376,N_25909,N_29739);
and U30377 (N_30377,N_28082,N_26184);
or U30378 (N_30378,N_28305,N_28836);
nor U30379 (N_30379,N_29822,N_26406);
nand U30380 (N_30380,N_29068,N_28298);
nand U30381 (N_30381,N_27736,N_25292);
nor U30382 (N_30382,N_25608,N_26786);
xnor U30383 (N_30383,N_27334,N_26794);
nor U30384 (N_30384,N_28844,N_26351);
nand U30385 (N_30385,N_27907,N_28736);
xnor U30386 (N_30386,N_29596,N_28211);
xnor U30387 (N_30387,N_25174,N_27262);
and U30388 (N_30388,N_28248,N_26105);
and U30389 (N_30389,N_28487,N_26191);
xor U30390 (N_30390,N_25684,N_26684);
and U30391 (N_30391,N_28026,N_25384);
nand U30392 (N_30392,N_28016,N_26166);
or U30393 (N_30393,N_28648,N_28401);
xor U30394 (N_30394,N_29227,N_25783);
nand U30395 (N_30395,N_27578,N_25001);
and U30396 (N_30396,N_28822,N_27050);
xor U30397 (N_30397,N_27919,N_25805);
and U30398 (N_30398,N_27160,N_28642);
xor U30399 (N_30399,N_29323,N_26520);
xnor U30400 (N_30400,N_25036,N_29949);
xor U30401 (N_30401,N_28992,N_25548);
nor U30402 (N_30402,N_26142,N_25266);
or U30403 (N_30403,N_29378,N_26721);
nor U30404 (N_30404,N_27748,N_29200);
xnor U30405 (N_30405,N_29534,N_28938);
xnor U30406 (N_30406,N_25431,N_25565);
xor U30407 (N_30407,N_28550,N_25011);
and U30408 (N_30408,N_25407,N_27260);
xor U30409 (N_30409,N_25616,N_28689);
or U30410 (N_30410,N_25637,N_26681);
nand U30411 (N_30411,N_28214,N_27233);
xnor U30412 (N_30412,N_26491,N_29926);
nand U30413 (N_30413,N_27383,N_26748);
nor U30414 (N_30414,N_27469,N_25069);
or U30415 (N_30415,N_28432,N_26344);
or U30416 (N_30416,N_26817,N_28441);
and U30417 (N_30417,N_25543,N_25151);
xor U30418 (N_30418,N_25226,N_29695);
xor U30419 (N_30419,N_28579,N_29406);
or U30420 (N_30420,N_29125,N_29748);
or U30421 (N_30421,N_25105,N_26350);
or U30422 (N_30422,N_26099,N_29658);
nor U30423 (N_30423,N_26172,N_27702);
nand U30424 (N_30424,N_25403,N_28110);
nor U30425 (N_30425,N_27574,N_26686);
nand U30426 (N_30426,N_27832,N_28884);
xnor U30427 (N_30427,N_26039,N_27848);
and U30428 (N_30428,N_26910,N_25094);
nand U30429 (N_30429,N_27496,N_27332);
nand U30430 (N_30430,N_25304,N_25855);
or U30431 (N_30431,N_29082,N_28732);
xnor U30432 (N_30432,N_27505,N_25301);
or U30433 (N_30433,N_25128,N_27620);
or U30434 (N_30434,N_25878,N_28621);
or U30435 (N_30435,N_27434,N_29417);
nand U30436 (N_30436,N_28321,N_28128);
and U30437 (N_30437,N_27688,N_26965);
xnor U30438 (N_30438,N_25289,N_26907);
nand U30439 (N_30439,N_25461,N_27077);
xnor U30440 (N_30440,N_29436,N_25191);
nand U30441 (N_30441,N_25975,N_25966);
or U30442 (N_30442,N_29425,N_28937);
nand U30443 (N_30443,N_28236,N_26033);
nand U30444 (N_30444,N_29111,N_29630);
xnor U30445 (N_30445,N_29066,N_26576);
nor U30446 (N_30446,N_27934,N_28520);
xnor U30447 (N_30447,N_29038,N_25212);
xnor U30448 (N_30448,N_27780,N_29577);
nor U30449 (N_30449,N_26106,N_25347);
and U30450 (N_30450,N_29735,N_27797);
xor U30451 (N_30451,N_26624,N_25928);
or U30452 (N_30452,N_29215,N_29281);
nor U30453 (N_30453,N_27149,N_25220);
nand U30454 (N_30454,N_25357,N_25840);
and U30455 (N_30455,N_27399,N_28212);
nor U30456 (N_30456,N_28300,N_29776);
nand U30457 (N_30457,N_28643,N_28482);
and U30458 (N_30458,N_26847,N_29234);
nor U30459 (N_30459,N_28828,N_29217);
and U30460 (N_30460,N_25367,N_28917);
or U30461 (N_30461,N_26034,N_26593);
or U30462 (N_30462,N_29830,N_25927);
xor U30463 (N_30463,N_29744,N_28498);
nand U30464 (N_30464,N_28975,N_25744);
and U30465 (N_30465,N_26307,N_26525);
or U30466 (N_30466,N_26571,N_26752);
xnor U30467 (N_30467,N_28356,N_28152);
or U30468 (N_30468,N_28535,N_28905);
or U30469 (N_30469,N_29128,N_25948);
or U30470 (N_30470,N_28181,N_29341);
nor U30471 (N_30471,N_26606,N_28471);
nor U30472 (N_30472,N_27436,N_25657);
xor U30473 (N_30473,N_27403,N_28655);
nand U30474 (N_30474,N_25922,N_28273);
xor U30475 (N_30475,N_29693,N_25210);
and U30476 (N_30476,N_29874,N_27443);
and U30477 (N_30477,N_27313,N_26321);
xor U30478 (N_30478,N_25027,N_26878);
xnor U30479 (N_30479,N_25064,N_25012);
xnor U30480 (N_30480,N_27898,N_28916);
and U30481 (N_30481,N_26846,N_25144);
and U30482 (N_30482,N_29656,N_27985);
and U30483 (N_30483,N_27955,N_25883);
or U30484 (N_30484,N_29432,N_29866);
nand U30485 (N_30485,N_25760,N_26988);
nor U30486 (N_30486,N_29092,N_29134);
xor U30487 (N_30487,N_26170,N_26696);
nor U30488 (N_30488,N_25689,N_26830);
nand U30489 (N_30489,N_26078,N_26613);
xnor U30490 (N_30490,N_26735,N_26053);
and U30491 (N_30491,N_28964,N_25542);
nor U30492 (N_30492,N_25389,N_28687);
xnor U30493 (N_30493,N_27980,N_26626);
or U30494 (N_30494,N_26024,N_29319);
nand U30495 (N_30495,N_25248,N_27644);
nor U30496 (N_30496,N_28092,N_29249);
xnor U30497 (N_30497,N_28945,N_29315);
nand U30498 (N_30498,N_25832,N_27918);
nor U30499 (N_30499,N_25765,N_29981);
nand U30500 (N_30500,N_27922,N_26101);
nor U30501 (N_30501,N_27349,N_28328);
nand U30502 (N_30502,N_29014,N_28561);
or U30503 (N_30503,N_25963,N_25940);
and U30504 (N_30504,N_25345,N_28683);
xor U30505 (N_30505,N_28872,N_25121);
nor U30506 (N_30506,N_27576,N_29410);
and U30507 (N_30507,N_26811,N_29401);
and U30508 (N_30508,N_27369,N_27793);
xnor U30509 (N_30509,N_27893,N_25753);
xor U30510 (N_30510,N_26783,N_29191);
or U30511 (N_30511,N_26442,N_25701);
and U30512 (N_30512,N_25773,N_28838);
xor U30513 (N_30513,N_27862,N_26500);
or U30514 (N_30514,N_27787,N_25486);
xnor U30515 (N_30515,N_29541,N_29964);
or U30516 (N_30516,N_27785,N_28050);
or U30517 (N_30517,N_26237,N_25711);
and U30518 (N_30518,N_29934,N_25766);
and U30519 (N_30519,N_28839,N_26833);
nand U30520 (N_30520,N_27240,N_26415);
xor U30521 (N_30521,N_27596,N_29148);
and U30522 (N_30522,N_27401,N_27739);
nor U30523 (N_30523,N_27657,N_25447);
and U30524 (N_30524,N_27398,N_28503);
or U30525 (N_30525,N_25098,N_27099);
nor U30526 (N_30526,N_28490,N_29646);
xnor U30527 (N_30527,N_25153,N_29069);
or U30528 (N_30528,N_27992,N_27068);
nor U30529 (N_30529,N_29336,N_29194);
and U30530 (N_30530,N_28398,N_29228);
nor U30531 (N_30531,N_29040,N_28096);
nand U30532 (N_30532,N_27761,N_25481);
or U30533 (N_30533,N_25278,N_26206);
or U30534 (N_30534,N_28592,N_29363);
nor U30535 (N_30535,N_26879,N_26976);
xor U30536 (N_30536,N_27150,N_29216);
nand U30537 (N_30537,N_29553,N_29011);
xor U30538 (N_30538,N_28048,N_28318);
and U30539 (N_30539,N_25066,N_27969);
nand U30540 (N_30540,N_28061,N_25862);
and U30541 (N_30541,N_26480,N_27900);
and U30542 (N_30542,N_25841,N_27827);
nand U30543 (N_30543,N_29507,N_25023);
or U30544 (N_30544,N_27782,N_26197);
or U30545 (N_30545,N_26127,N_25933);
xor U30546 (N_30546,N_29923,N_27952);
or U30547 (N_30547,N_25205,N_26369);
or U30548 (N_30548,N_27859,N_28419);
xnor U30549 (N_30549,N_25628,N_27359);
nand U30550 (N_30550,N_25980,N_29219);
and U30551 (N_30551,N_27805,N_27064);
nor U30552 (N_30552,N_26551,N_26869);
and U30553 (N_30553,N_27216,N_27118);
nor U30554 (N_30554,N_25998,N_26014);
xnor U30555 (N_30555,N_25218,N_27742);
and U30556 (N_30556,N_28586,N_27630);
nor U30557 (N_30557,N_25155,N_28762);
or U30558 (N_30558,N_26154,N_27234);
xor U30559 (N_30559,N_27668,N_26587);
and U30560 (N_30560,N_29550,N_29392);
xnor U30561 (N_30561,N_29605,N_27509);
xor U30562 (N_30562,N_25393,N_28752);
xnor U30563 (N_30563,N_26010,N_27170);
nand U30564 (N_30564,N_29876,N_29848);
xnor U30565 (N_30565,N_28336,N_27279);
and U30566 (N_30566,N_26440,N_26689);
xor U30567 (N_30567,N_29223,N_25667);
xnor U30568 (N_30568,N_25881,N_25800);
or U30569 (N_30569,N_28232,N_29369);
nand U30570 (N_30570,N_29377,N_28416);
nor U30571 (N_30571,N_28093,N_26019);
nor U30572 (N_30572,N_29733,N_27507);
xor U30573 (N_30573,N_28306,N_28630);
xnor U30574 (N_30574,N_28426,N_26777);
nor U30575 (N_30575,N_25511,N_28303);
nand U30576 (N_30576,N_28133,N_29547);
nor U30577 (N_30577,N_27080,N_26719);
nor U30578 (N_30578,N_26454,N_27802);
xnor U30579 (N_30579,N_28650,N_28361);
xnor U30580 (N_30580,N_29501,N_25690);
nor U30581 (N_30581,N_29118,N_27101);
or U30582 (N_30582,N_25953,N_25950);
nand U30583 (N_30583,N_25512,N_26277);
or U30584 (N_30584,N_26215,N_27001);
nand U30585 (N_30585,N_27660,N_29844);
and U30586 (N_30586,N_26772,N_25067);
nand U30587 (N_30587,N_29049,N_28488);
nand U30588 (N_30588,N_29511,N_25544);
nand U30589 (N_30589,N_28308,N_26465);
and U30590 (N_30590,N_29373,N_27600);
nor U30591 (N_30591,N_28787,N_26190);
xor U30592 (N_30592,N_29891,N_26221);
xnor U30593 (N_30593,N_29655,N_27023);
nand U30594 (N_30594,N_29442,N_25540);
xnor U30595 (N_30595,N_27890,N_25741);
nor U30596 (N_30596,N_25441,N_27762);
and U30597 (N_30597,N_28150,N_28747);
nand U30598 (N_30598,N_26490,N_28270);
nor U30599 (N_30599,N_26509,N_27613);
nor U30600 (N_30600,N_29967,N_27028);
and U30601 (N_30601,N_28922,N_27019);
nand U30602 (N_30602,N_25095,N_26203);
nor U30603 (N_30603,N_26806,N_28965);
xor U30604 (N_30604,N_28845,N_29688);
nor U30605 (N_30605,N_28913,N_26135);
xor U30606 (N_30606,N_28465,N_26659);
xor U30607 (N_30607,N_29379,N_29612);
or U30608 (N_30608,N_26943,N_25318);
or U30609 (N_30609,N_27290,N_25531);
nor U30610 (N_30610,N_29492,N_25530);
xor U30611 (N_30611,N_28404,N_25088);
or U30612 (N_30612,N_26519,N_26921);
xor U30613 (N_30613,N_25136,N_28569);
nor U30614 (N_30614,N_26469,N_28532);
nand U30615 (N_30615,N_25320,N_28006);
and U30616 (N_30616,N_27677,N_25560);
and U30617 (N_30617,N_26424,N_25264);
xor U30618 (N_30618,N_26730,N_26710);
xor U30619 (N_30619,N_28639,N_25851);
nand U30620 (N_30620,N_29295,N_28659);
xor U30621 (N_30621,N_26436,N_26400);
or U30622 (N_30622,N_26052,N_25274);
or U30623 (N_30623,N_25902,N_28989);
nor U30624 (N_30624,N_29602,N_25127);
nand U30625 (N_30625,N_26535,N_29621);
nand U30626 (N_30626,N_26558,N_28111);
xor U30627 (N_30627,N_27706,N_29514);
nor U30628 (N_30628,N_26435,N_29824);
and U30629 (N_30629,N_25047,N_29540);
nor U30630 (N_30630,N_25117,N_25146);
nand U30631 (N_30631,N_29086,N_26144);
and U30632 (N_30632,N_29242,N_26756);
or U30633 (N_30633,N_28027,N_27241);
or U30634 (N_30634,N_25979,N_29241);
xor U30635 (N_30635,N_29420,N_25162);
nor U30636 (N_30636,N_26912,N_29791);
nor U30637 (N_30637,N_27348,N_29843);
nand U30638 (N_30638,N_26336,N_29641);
and U30639 (N_30639,N_29285,N_27347);
xnor U30640 (N_30640,N_27396,N_26217);
and U30641 (N_30641,N_26953,N_27566);
xnor U30642 (N_30642,N_27966,N_27806);
or U30643 (N_30643,N_26896,N_29186);
nand U30644 (N_30644,N_29141,N_26873);
xor U30645 (N_30645,N_27627,N_26259);
nand U30646 (N_30646,N_27012,N_25959);
or U30647 (N_30647,N_27244,N_29798);
xor U30648 (N_30648,N_26460,N_28940);
or U30649 (N_30649,N_29268,N_26441);
xor U30650 (N_30650,N_27756,N_28694);
nor U30651 (N_30651,N_25237,N_29962);
and U30652 (N_30652,N_25536,N_27989);
or U30653 (N_30653,N_27454,N_29838);
or U30654 (N_30654,N_27081,N_28521);
xor U30655 (N_30655,N_27961,N_25324);
xnor U30656 (N_30656,N_26495,N_27308);
or U30657 (N_30657,N_25187,N_28702);
xnor U30658 (N_30658,N_28357,N_25771);
nor U30659 (N_30659,N_27094,N_29508);
xnor U30660 (N_30660,N_25494,N_27871);
and U30661 (N_30661,N_28225,N_26453);
nor U30662 (N_30662,N_27499,N_26118);
and U30663 (N_30663,N_27759,N_27267);
nor U30664 (N_30664,N_27845,N_25179);
and U30665 (N_30665,N_25717,N_26774);
nor U30666 (N_30666,N_26985,N_28013);
nor U30667 (N_30667,N_26361,N_26619);
xnor U30668 (N_30668,N_28329,N_26533);
nand U30669 (N_30669,N_25445,N_25696);
nand U30670 (N_30670,N_28991,N_26632);
or U30671 (N_30671,N_26055,N_25951);
nand U30672 (N_30672,N_28784,N_28235);
nand U30673 (N_30673,N_27270,N_25794);
nand U30674 (N_30674,N_27131,N_26009);
nand U30675 (N_30675,N_28081,N_26095);
xor U30676 (N_30676,N_26653,N_29291);
nand U30677 (N_30677,N_28806,N_26541);
and U30678 (N_30678,N_27311,N_26724);
xor U30679 (N_30679,N_29747,N_28962);
and U30680 (N_30680,N_29917,N_26546);
nand U30681 (N_30681,N_29581,N_28594);
nand U30682 (N_30682,N_27274,N_28493);
and U30683 (N_30683,N_27673,N_26995);
nor U30684 (N_30684,N_29316,N_25426);
nand U30685 (N_30685,N_28563,N_27110);
nor U30686 (N_30686,N_27927,N_25968);
nor U30687 (N_30687,N_27448,N_27183);
and U30688 (N_30688,N_28779,N_25864);
and U30689 (N_30689,N_25809,N_26075);
xor U30690 (N_30690,N_25874,N_25789);
nand U30691 (N_30691,N_28095,N_28956);
or U30692 (N_30692,N_29403,N_26868);
or U30693 (N_30693,N_27740,N_25723);
xor U30694 (N_30694,N_26527,N_27171);
or U30695 (N_30695,N_28162,N_25799);
nor U30696 (N_30696,N_28652,N_28021);
nand U30697 (N_30697,N_25421,N_28327);
and U30698 (N_30698,N_27258,N_28705);
xnor U30699 (N_30699,N_27213,N_28279);
nand U30700 (N_30700,N_26577,N_25037);
xor U30701 (N_30701,N_27994,N_29956);
nor U30702 (N_30702,N_28849,N_25206);
xnor U30703 (N_30703,N_27303,N_27129);
and U30704 (N_30704,N_28406,N_25170);
xor U30705 (N_30705,N_25224,N_27580);
and U30706 (N_30706,N_29600,N_28601);
nand U30707 (N_30707,N_25676,N_26886);
nand U30708 (N_30708,N_28015,N_29840);
nor U30709 (N_30709,N_26544,N_25734);
and U30710 (N_30710,N_28804,N_28727);
nor U30711 (N_30711,N_28289,N_29407);
nor U30712 (N_30712,N_27836,N_28220);
and U30713 (N_30713,N_26940,N_26300);
or U30714 (N_30714,N_28982,N_25612);
and U30715 (N_30715,N_26355,N_26410);
or U30716 (N_30716,N_26278,N_28287);
or U30717 (N_30717,N_27191,N_26820);
or U30718 (N_30718,N_29455,N_27665);
and U30719 (N_30719,N_29318,N_25983);
and U30720 (N_30720,N_27248,N_28831);
xor U30721 (N_30721,N_27920,N_25655);
xnor U30722 (N_30722,N_29609,N_29334);
xnor U30723 (N_30723,N_29590,N_25956);
nor U30724 (N_30724,N_28019,N_26510);
xor U30725 (N_30725,N_28219,N_25381);
xor U30726 (N_30726,N_28866,N_25903);
or U30727 (N_30727,N_26360,N_27482);
or U30728 (N_30728,N_26567,N_29260);
and U30729 (N_30729,N_25216,N_26475);
or U30730 (N_30730,N_26642,N_26479);
nor U30731 (N_30731,N_28411,N_29564);
or U30732 (N_30732,N_26853,N_29788);
nor U30733 (N_30733,N_25173,N_26027);
nand U30734 (N_30734,N_25824,N_25368);
and U30735 (N_30735,N_27265,N_29676);
xor U30736 (N_30736,N_27869,N_25111);
and U30737 (N_30737,N_28384,N_25643);
nor U30738 (N_30738,N_29505,N_28921);
nor U30739 (N_30739,N_27330,N_27820);
nor U30740 (N_30740,N_26303,N_28739);
nand U30741 (N_30741,N_25699,N_25529);
or U30742 (N_30742,N_27465,N_29124);
xor U30743 (N_30743,N_26030,N_26885);
and U30744 (N_30744,N_27928,N_28475);
nor U30745 (N_30745,N_25905,N_29032);
nor U30746 (N_30746,N_26492,N_28939);
nor U30747 (N_30747,N_26265,N_26929);
and U30748 (N_30748,N_25026,N_29331);
xor U30749 (N_30749,N_26620,N_28645);
nand U30750 (N_30750,N_25437,N_26496);
nor U30751 (N_30751,N_27083,N_26581);
nand U30752 (N_30752,N_29065,N_29601);
nand U30753 (N_30753,N_27005,N_27945);
nor U30754 (N_30754,N_26640,N_25158);
and U30755 (N_30755,N_25808,N_26580);
and U30756 (N_30756,N_27058,N_28479);
nor U30757 (N_30757,N_25505,N_25907);
xnor U30758 (N_30758,N_29473,N_25836);
xor U30759 (N_30759,N_26871,N_28409);
nor U30760 (N_30760,N_29504,N_27973);
or U30761 (N_30761,N_27491,N_28102);
nand U30762 (N_30762,N_29673,N_26897);
or U30763 (N_30763,N_25702,N_29376);
nor U30764 (N_30764,N_27091,N_25363);
or U30765 (N_30765,N_25784,N_29449);
nor U30766 (N_30766,N_28778,N_25490);
and U30767 (N_30767,N_29500,N_29548);
or U30768 (N_30768,N_29696,N_27750);
or U30769 (N_30769,N_27172,N_27370);
nor U30770 (N_30770,N_26566,N_28793);
or U30771 (N_30771,N_25468,N_25112);
and U30772 (N_30772,N_26919,N_26296);
xor U30773 (N_30773,N_27420,N_25757);
xor U30774 (N_30774,N_27501,N_26993);
and U30775 (N_30775,N_25024,N_27429);
and U30776 (N_30776,N_29391,N_29288);
or U30777 (N_30777,N_25252,N_28548);
and U30778 (N_30778,N_28144,N_29664);
nor U30779 (N_30779,N_26036,N_26159);
xor U30780 (N_30780,N_28502,N_29717);
and U30781 (N_30781,N_27133,N_27831);
xor U30782 (N_30782,N_28695,N_29247);
xnor U30783 (N_30783,N_25735,N_25647);
or U30784 (N_30784,N_26722,N_29329);
xor U30785 (N_30785,N_27634,N_28156);
nand U30786 (N_30786,N_27938,N_28231);
or U30787 (N_30787,N_26970,N_28052);
and U30788 (N_30788,N_28089,N_26179);
nor U30789 (N_30789,N_29719,N_26754);
nand U30790 (N_30790,N_25479,N_25607);
and U30791 (N_30791,N_29015,N_25249);
nand U30792 (N_30792,N_27884,N_28099);
and U30793 (N_30793,N_29726,N_26883);
nand U30794 (N_30794,N_28977,N_26630);
nand U30795 (N_30795,N_28800,N_26603);
nor U30796 (N_30796,N_28788,N_28783);
or U30797 (N_30797,N_26742,N_26860);
xor U30798 (N_30798,N_26346,N_26563);
and U30799 (N_30799,N_28041,N_27354);
and U30800 (N_30800,N_26540,N_27433);
nand U30801 (N_30801,N_25016,N_28670);
xnor U30802 (N_30802,N_26954,N_28299);
nand U30803 (N_30803,N_28193,N_28742);
nand U30804 (N_30804,N_25473,N_26612);
or U30805 (N_30805,N_26422,N_28047);
or U30806 (N_30806,N_25502,N_25835);
nor U30807 (N_30807,N_27573,N_25126);
nand U30808 (N_30808,N_27522,N_27982);
nand U30809 (N_30809,N_29184,N_27758);
nor U30810 (N_30810,N_28458,N_28770);
and U30811 (N_30811,N_27154,N_25893);
and U30812 (N_30812,N_27467,N_25828);
and U30813 (N_30813,N_25811,N_26338);
and U30814 (N_30814,N_26365,N_29259);
or U30815 (N_30815,N_25424,N_26072);
and U30816 (N_30816,N_25193,N_26056);
nand U30817 (N_30817,N_29007,N_26155);
xnor U30818 (N_30818,N_25458,N_29290);
xor U30819 (N_30819,N_28957,N_28108);
nor U30820 (N_30820,N_27775,N_28595);
and U30821 (N_30821,N_29978,N_28242);
nor U30822 (N_30822,N_27881,N_27340);
xor U30823 (N_30823,N_27579,N_26074);
xor U30824 (N_30824,N_26727,N_25926);
and U30825 (N_30825,N_27784,N_29812);
xor U30826 (N_30826,N_29368,N_28635);
or U30827 (N_30827,N_25195,N_27903);
nand U30828 (N_30828,N_26585,N_26635);
nand U30829 (N_30829,N_29470,N_26048);
and U30830 (N_30830,N_26082,N_26704);
nor U30831 (N_30831,N_25597,N_25613);
and U30832 (N_30832,N_26617,N_26168);
xor U30833 (N_30833,N_28846,N_29427);
nor U30834 (N_30834,N_28049,N_26627);
nor U30835 (N_30835,N_25843,N_28673);
nor U30836 (N_30836,N_25446,N_28582);
xnor U30837 (N_30837,N_27435,N_25108);
xnor U30838 (N_30838,N_26731,N_26378);
xor U30839 (N_30839,N_26079,N_25223);
nand U30840 (N_30840,N_29723,N_26776);
or U30841 (N_30841,N_28180,N_28817);
nand U30842 (N_30842,N_29503,N_26548);
and U30843 (N_30843,N_25250,N_26482);
or U30844 (N_30844,N_25845,N_26322);
or U30845 (N_30845,N_25156,N_29879);
or U30846 (N_30846,N_26792,N_28340);
nor U30847 (N_30847,N_28723,N_29448);
nand U30848 (N_30848,N_26946,N_25409);
or U30849 (N_30849,N_26294,N_29067);
xnor U30850 (N_30850,N_26250,N_28310);
xnor U30851 (N_30851,N_27818,N_27678);
nor U30852 (N_30852,N_28809,N_27997);
nand U30853 (N_30853,N_26937,N_29287);
nand U30854 (N_30854,N_29560,N_25148);
or U30855 (N_30855,N_26396,N_27057);
and U30856 (N_30856,N_28930,N_27104);
xor U30857 (N_30857,N_29144,N_27141);
xnor U30858 (N_30858,N_29811,N_28137);
and U30859 (N_30859,N_27585,N_27053);
nor U30860 (N_30860,N_25742,N_26218);
nand U30861 (N_30861,N_25295,N_29344);
and U30862 (N_30862,N_29476,N_25222);
nand U30863 (N_30863,N_27128,N_26644);
or U30864 (N_30864,N_25868,N_29233);
nand U30865 (N_30865,N_25271,N_29782);
nand U30866 (N_30866,N_26634,N_25059);
or U30867 (N_30867,N_25413,N_29953);
nor U30868 (N_30868,N_25638,N_28706);
xnor U30869 (N_30869,N_26904,N_26605);
nand U30870 (N_30870,N_27200,N_26598);
or U30871 (N_30871,N_29780,N_27463);
and U30872 (N_30872,N_28174,N_26291);
nand U30873 (N_30873,N_29936,N_25438);
nor U30874 (N_30874,N_28347,N_26651);
xnor U30875 (N_30875,N_29304,N_27102);
nor U30876 (N_30876,N_25570,N_27542);
nor U30877 (N_30877,N_27708,N_28583);
and U30878 (N_30878,N_28164,N_25995);
nor U30879 (N_30879,N_27725,N_28679);
xnor U30880 (N_30880,N_26909,N_27275);
or U30881 (N_30881,N_27009,N_27471);
and U30882 (N_30882,N_29980,N_27415);
nand U30883 (N_30883,N_29555,N_26770);
nand U30884 (N_30884,N_25103,N_29899);
nand U30885 (N_30885,N_28820,N_28309);
nand U30886 (N_30886,N_29372,N_28187);
and U30887 (N_30887,N_26505,N_29272);
or U30888 (N_30888,N_27459,N_27475);
and U30889 (N_30889,N_28072,N_29740);
or U30890 (N_30890,N_25610,N_26462);
xor U30891 (N_30891,N_29554,N_28171);
nor U30892 (N_30892,N_29974,N_25535);
nand U30893 (N_30893,N_27307,N_26187);
nand U30894 (N_30894,N_25731,N_27538);
xor U30895 (N_30895,N_25244,N_29721);
nor U30896 (N_30896,N_28143,N_28827);
nor U30897 (N_30897,N_28543,N_29238);
nand U30898 (N_30898,N_26658,N_25102);
xor U30899 (N_30899,N_25182,N_29299);
nand U30900 (N_30900,N_25931,N_25030);
nor U30901 (N_30901,N_29828,N_25457);
xor U30902 (N_30902,N_25474,N_29048);
nor U30903 (N_30903,N_27440,N_26341);
xnor U30904 (N_30904,N_25586,N_27828);
or U30905 (N_30905,N_27514,N_29298);
or U30906 (N_30906,N_28692,N_27096);
or U30907 (N_30907,N_26051,N_25880);
nor U30908 (N_30908,N_25533,N_25510);
or U30909 (N_30909,N_28063,N_28275);
xnor U30910 (N_30910,N_27045,N_25165);
nor U30911 (N_30911,N_28438,N_25263);
xnor U30912 (N_30912,N_28088,N_28059);
nand U30913 (N_30913,N_27220,N_25480);
nand U30914 (N_30914,N_25686,N_29123);
and U30915 (N_30915,N_29808,N_28728);
nor U30916 (N_30916,N_28400,N_27626);
nor U30917 (N_30917,N_29922,N_27829);
nor U30918 (N_30918,N_29453,N_25624);
nor U30919 (N_30919,N_28842,N_25062);
xor U30920 (N_30920,N_28810,N_26611);
or U30921 (N_30921,N_28077,N_26974);
or U30922 (N_30922,N_25672,N_26140);
or U30923 (N_30923,N_25375,N_27962);
nor U30924 (N_30924,N_28553,N_27795);
and U30925 (N_30925,N_28380,N_25635);
nor U30926 (N_30926,N_27428,N_29126);
nor U30927 (N_30927,N_26399,N_27197);
nor U30928 (N_30928,N_25775,N_27305);
or U30929 (N_30929,N_29971,N_29837);
nand U30930 (N_30930,N_28177,N_25360);
or U30931 (N_30931,N_28222,N_26240);
and U30932 (N_30932,N_28870,N_25214);
or U30933 (N_30933,N_27203,N_27892);
nand U30934 (N_30934,N_26739,N_25621);
or U30935 (N_30935,N_29754,N_27592);
and U30936 (N_30936,N_27967,N_29306);
or U30937 (N_30937,N_25477,N_28680);
nand U30938 (N_30938,N_27520,N_25564);
and U30939 (N_30939,N_29365,N_29301);
xor U30940 (N_30940,N_25592,N_26582);
nand U30941 (N_30941,N_28036,N_26625);
nor U30942 (N_30942,N_28947,N_26000);
or U30943 (N_30943,N_26493,N_25659);
and U30944 (N_30944,N_26950,N_27087);
nand U30945 (N_30945,N_26330,N_29332);
xnor U30946 (N_30946,N_29686,N_26041);
xor U30947 (N_30947,N_26256,N_25882);
nor U30948 (N_30948,N_25235,N_25184);
xnor U30949 (N_30949,N_26655,N_26832);
nand U30950 (N_30950,N_29140,N_27230);
and U30951 (N_30951,N_27033,N_29565);
and U30952 (N_30952,N_29078,N_27352);
or U30953 (N_30953,N_28534,N_27873);
or U30954 (N_30954,N_26201,N_27976);
nor U30955 (N_30955,N_28851,N_28600);
nand U30956 (N_30956,N_29589,N_26743);
nor U30957 (N_30957,N_29497,N_26138);
or U30958 (N_30958,N_25818,N_28560);
nand U30959 (N_30959,N_27584,N_27766);
nor U30960 (N_30960,N_26768,N_27235);
nand U30961 (N_30961,N_27916,N_27061);
or U30962 (N_30962,N_26452,N_25044);
xnor U30963 (N_30963,N_28381,N_28265);
xnor U30964 (N_30964,N_26043,N_28112);
or U30965 (N_30965,N_27406,N_27067);
nor U30966 (N_30966,N_29820,N_25630);
and U30967 (N_30967,N_28179,N_25752);
or U30968 (N_30968,N_25721,N_28374);
or U30969 (N_30969,N_29346,N_25942);
nand U30970 (N_30970,N_28731,N_29628);
or U30971 (N_30971,N_29409,N_27625);
or U30972 (N_30972,N_29480,N_26916);
nand U30973 (N_30973,N_28688,N_29164);
nand U30974 (N_30974,N_28463,N_27004);
xor U30975 (N_30975,N_25110,N_25945);
xor U30976 (N_30976,N_25465,N_25253);
or U30977 (N_30977,N_26744,N_26959);
xnor U30978 (N_30978,N_27199,N_28062);
nand U30979 (N_30979,N_25894,N_27760);
or U30980 (N_30980,N_28383,N_29831);
xnor U30981 (N_30981,N_28022,N_27054);
and U30982 (N_30982,N_27964,N_29495);
nor U30983 (N_30983,N_26766,N_25896);
xor U30984 (N_30984,N_28107,N_28345);
and U30985 (N_30985,N_29154,N_27317);
nand U30986 (N_30986,N_27423,N_26914);
or U30987 (N_30987,N_29355,N_29398);
nor U30988 (N_30988,N_28280,N_29098);
or U30989 (N_30989,N_27540,N_26243);
nand U30990 (N_30990,N_28632,N_26690);
nor U30991 (N_30991,N_28886,N_27944);
xor U30992 (N_30992,N_25310,N_27939);
xnor U30993 (N_30993,N_29996,N_29674);
nand U30994 (N_30994,N_26120,N_29314);
xor U30995 (N_30995,N_26643,N_29706);
nand U30996 (N_30996,N_29404,N_25602);
or U30997 (N_30997,N_26471,N_28933);
nor U30998 (N_30998,N_25786,N_25581);
xnor U30999 (N_30999,N_29472,N_29063);
nand U31000 (N_31000,N_26803,N_27870);
xnor U31001 (N_31001,N_27325,N_26859);
and U31002 (N_31002,N_29991,N_25190);
xor U31003 (N_31003,N_26065,N_26797);
xor U31004 (N_31004,N_27763,N_25256);
xnor U31005 (N_31005,N_26332,N_29770);
xor U31006 (N_31006,N_25890,N_26038);
nor U31007 (N_31007,N_29311,N_25961);
or U31008 (N_31008,N_25691,N_28898);
or U31009 (N_31009,N_28379,N_26848);
nand U31010 (N_31010,N_29097,N_28573);
xnor U31011 (N_31011,N_28829,N_27728);
nand U31012 (N_31012,N_28155,N_29326);
nand U31013 (N_31013,N_29562,N_25580);
or U31014 (N_31014,N_25487,N_26999);
nand U31015 (N_31015,N_26331,N_28341);
xor U31016 (N_31016,N_26740,N_28131);
nor U31017 (N_31017,N_26892,N_25321);
and U31018 (N_31018,N_28461,N_25313);
nor U31019 (N_31019,N_25938,N_27105);
nand U31020 (N_31020,N_26474,N_27476);
or U31021 (N_31021,N_25692,N_26260);
or U31022 (N_31022,N_27524,N_28772);
and U31023 (N_31023,N_26439,N_29354);
nor U31024 (N_31024,N_28334,N_27747);
xor U31025 (N_31025,N_28850,N_26779);
xnor U31026 (N_31026,N_29595,N_27107);
xnor U31027 (N_31027,N_26008,N_29896);
nor U31028 (N_31028,N_25464,N_28203);
and U31029 (N_31029,N_26327,N_26418);
nor U31030 (N_31030,N_25196,N_26762);
or U31031 (N_31031,N_26670,N_25639);
xnor U31032 (N_31032,N_26996,N_29009);
xnor U31033 (N_31033,N_25814,N_27745);
xnor U31034 (N_31034,N_27458,N_29389);
and U31035 (N_31035,N_28578,N_27421);
xor U31036 (N_31036,N_27337,N_29159);
nand U31037 (N_31037,N_27674,N_26952);
nor U31038 (N_31038,N_27690,N_28119);
and U31039 (N_31039,N_26729,N_28480);
nor U31040 (N_31040,N_26401,N_26862);
and U31041 (N_31041,N_29208,N_26836);
xor U31042 (N_31042,N_25262,N_28069);
nor U31043 (N_31043,N_28678,N_27547);
xor U31044 (N_31044,N_25315,N_29910);
nand U31045 (N_31045,N_27622,N_27209);
nand U31046 (N_31046,N_29919,N_26828);
and U31047 (N_31047,N_25364,N_29659);
xor U31048 (N_31048,N_26282,N_26185);
xnor U31049 (N_31049,N_28768,N_26979);
xnor U31050 (N_31050,N_27891,N_25472);
or U31051 (N_31051,N_26596,N_28763);
and U31052 (N_31052,N_27034,N_29594);
nor U31053 (N_31053,N_25708,N_26945);
nor U31054 (N_31054,N_27709,N_29027);
xnor U31055 (N_31055,N_29447,N_27236);
xor U31056 (N_31056,N_28130,N_25134);
or U31057 (N_31057,N_26662,N_29761);
and U31058 (N_31058,N_28140,N_29440);
and U31059 (N_31059,N_25408,N_27651);
and U31060 (N_31060,N_27754,N_28733);
xor U31061 (N_31061,N_29214,N_26650);
nor U31062 (N_31062,N_28436,N_26007);
or U31063 (N_31063,N_29778,N_29226);
nand U31064 (N_31064,N_25598,N_25201);
nor U31065 (N_31065,N_27363,N_28606);
nor U31066 (N_31066,N_29270,N_28741);
nor U31067 (N_31067,N_26706,N_29887);
nor U31068 (N_31068,N_29904,N_27125);
xnor U31069 (N_31069,N_27664,N_29142);
xnor U31070 (N_31070,N_25484,N_29648);
and U31071 (N_31071,N_28668,N_27073);
nand U31072 (N_31072,N_29588,N_26591);
xnor U31073 (N_31073,N_28651,N_26445);
xor U31074 (N_31074,N_26707,N_28572);
nand U31075 (N_31075,N_25791,N_26583);
or U31076 (N_31076,N_28567,N_26780);
or U31077 (N_31077,N_29256,N_28802);
nand U31078 (N_31078,N_26503,N_27864);
or U31079 (N_31079,N_26113,N_27051);
nor U31080 (N_31080,N_25429,N_29173);
or U31081 (N_31081,N_29423,N_29371);
and U31082 (N_31082,N_25954,N_29364);
nor U31083 (N_31083,N_28312,N_26526);
or U31084 (N_31084,N_27282,N_25152);
nand U31085 (N_31085,N_28147,N_25585);
nand U31086 (N_31086,N_29677,N_29016);
nand U31087 (N_31087,N_29846,N_28618);
or U31088 (N_31088,N_27374,N_25302);
or U31089 (N_31089,N_26081,N_29683);
and U31090 (N_31090,N_28823,N_25719);
or U31091 (N_31091,N_27854,N_26254);
or U31092 (N_31092,N_26323,N_26518);
nor U31093 (N_31093,N_28241,N_29411);
or U31094 (N_31094,N_27389,N_25929);
xor U31095 (N_31095,N_28570,N_29248);
nor U31096 (N_31096,N_26455,N_25167);
nand U31097 (N_31097,N_25913,N_27556);
xor U31098 (N_31098,N_27888,N_25455);
nand U31099 (N_31099,N_29506,N_28330);
or U31100 (N_31100,N_26425,N_26903);
xor U31101 (N_31101,N_25770,N_27291);
nor U31102 (N_31102,N_27561,N_28367);
nand U31103 (N_31103,N_27713,N_26486);
nor U31104 (N_31104,N_29975,N_29924);
xor U31105 (N_31105,N_29892,N_26345);
or U31106 (N_31106,N_25652,N_25022);
nand U31107 (N_31107,N_28615,N_26781);
or U31108 (N_31108,N_26416,N_27323);
or U31109 (N_31109,N_27510,N_25559);
nor U31110 (N_31110,N_28657,N_27560);
nor U31111 (N_31111,N_25594,N_28178);
xnor U31112 (N_31112,N_26720,N_28604);
nand U31113 (N_31113,N_26196,N_27608);
xnor U31114 (N_31114,N_27588,N_26320);
nand U31115 (N_31115,N_27412,N_27134);
xor U31116 (N_31116,N_28323,N_28453);
xor U31117 (N_31117,N_27124,N_29531);
or U31118 (N_31118,N_25236,N_25626);
or U31119 (N_31119,N_28338,N_29045);
nand U31120 (N_31120,N_25404,N_25054);
xor U31121 (N_31121,N_29324,N_26538);
or U31122 (N_31122,N_27839,N_25790);
nor U31123 (N_31123,N_28753,N_27484);
and U31124 (N_31124,N_29499,N_28319);
xor U31125 (N_31125,N_25425,N_26377);
and U31126 (N_31126,N_29574,N_27995);
nor U31127 (N_31127,N_28697,N_27897);
xor U31128 (N_31128,N_29537,N_26040);
and U31129 (N_31129,N_26459,N_29932);
and U31130 (N_31130,N_25653,N_27814);
or U31131 (N_31131,N_28874,N_28469);
and U31132 (N_31132,N_27365,N_26162);
and U31133 (N_31133,N_25780,N_27084);
nand U31134 (N_31134,N_25519,N_28909);
nor U31135 (N_31135,N_27259,N_25716);
xor U31136 (N_31136,N_26588,N_28641);
nor U31137 (N_31137,N_27856,N_25175);
and U31138 (N_31138,N_26464,N_28781);
nor U31139 (N_31139,N_26035,N_28510);
nor U31140 (N_31140,N_26674,N_27085);
or U31141 (N_31141,N_26088,N_27874);
nor U31142 (N_31142,N_25161,N_26409);
nor U31143 (N_31143,N_29889,N_27285);
nor U31144 (N_31144,N_28259,N_28067);
nand U31145 (N_31145,N_28912,N_26782);
or U31146 (N_31146,N_29897,N_26841);
or U31147 (N_31147,N_27889,N_28448);
nand U31148 (N_31148,N_25471,N_29396);
xnor U31149 (N_31149,N_29653,N_28010);
nor U31150 (N_31150,N_27113,N_25515);
or U31151 (N_31151,N_29257,N_29468);
nand U31152 (N_31152,N_28464,N_27092);
nor U31153 (N_31153,N_28444,N_25469);
nor U31154 (N_31154,N_26325,N_29813);
nor U31155 (N_31155,N_27074,N_28423);
nor U31156 (N_31156,N_29895,N_26809);
and U31157 (N_31157,N_26405,N_28483);
and U31158 (N_31158,N_26421,N_29160);
or U31159 (N_31159,N_27152,N_26506);
xnor U31160 (N_31160,N_29965,N_28191);
xor U31161 (N_31161,N_27202,N_29137);
nand U31162 (N_31162,N_27371,N_25736);
nand U31163 (N_31163,N_25955,N_28408);
nand U31164 (N_31164,N_28315,N_25577);
nand U31165 (N_31165,N_26443,N_28002);
xnor U31166 (N_31166,N_27647,N_28666);
nor U31167 (N_31167,N_29905,N_25557);
nand U31168 (N_31168,N_26366,N_28685);
xnor U31169 (N_31169,N_27880,N_25058);
nor U31170 (N_31170,N_26225,N_29552);
nand U31171 (N_31171,N_25865,N_25033);
xor U31172 (N_31172,N_26709,N_28422);
nor U31173 (N_31173,N_25129,N_25693);
and U31174 (N_31174,N_28281,N_27602);
nor U31175 (N_31175,N_27697,N_29303);
xor U31176 (N_31176,N_29773,N_28805);
or U31177 (N_31177,N_25705,N_28985);
xor U31178 (N_31178,N_28590,N_29382);
nor U31179 (N_31179,N_25837,N_27404);
or U31180 (N_31180,N_25018,N_29787);
xnor U31181 (N_31181,N_27650,N_26063);
or U31182 (N_31182,N_29367,N_26005);
nor U31183 (N_31183,N_28587,N_27661);
and U31184 (N_31184,N_26688,N_29881);
nor U31185 (N_31185,N_27799,N_26543);
and U31186 (N_31186,N_29794,N_26601);
and U31187 (N_31187,N_26573,N_25863);
and U31188 (N_31188,N_27841,N_26761);
or U31189 (N_31189,N_26552,N_26397);
nor U31190 (N_31190,N_25072,N_29175);
or U31191 (N_31191,N_25755,N_29243);
nand U31192 (N_31192,N_26091,N_25972);
xnor U31193 (N_31193,N_26204,N_25782);
nor U31194 (N_31194,N_27971,N_26949);
xor U31195 (N_31195,N_26211,N_27417);
and U31196 (N_31196,N_25135,N_28230);
xnor U31197 (N_31197,N_28513,N_27993);
nor U31198 (N_31198,N_25475,N_27649);
nor U31199 (N_31199,N_27327,N_25396);
nand U31200 (N_31200,N_28971,N_25268);
xnor U31201 (N_31201,N_29158,N_28337);
or U31202 (N_31202,N_26928,N_25660);
xor U31203 (N_31203,N_27245,N_28146);
and U31204 (N_31204,N_29578,N_25797);
nor U31205 (N_31205,N_25427,N_27899);
or U31206 (N_31206,N_29878,N_28871);
xnor U31207 (N_31207,N_25969,N_25015);
nor U31208 (N_31208,N_26737,N_28826);
nand U31209 (N_31209,N_29183,N_28714);
or U31210 (N_31210,N_29633,N_29635);
xnor U31211 (N_31211,N_27002,N_25698);
and U31212 (N_31212,N_29660,N_26006);
nand U31213 (N_31213,N_29058,N_29457);
xnor U31214 (N_31214,N_25171,N_29781);
xor U31215 (N_31215,N_27445,N_25233);
xor U31216 (N_31216,N_28190,N_29692);
xor U31217 (N_31217,N_29741,N_25104);
nor U31218 (N_31218,N_28157,N_28545);
nand U31219 (N_31219,N_27648,N_27362);
and U31220 (N_31220,N_28079,N_25002);
and U31221 (N_31221,N_27027,N_25807);
and U31222 (N_31222,N_26522,N_26677);
nor U31223 (N_31223,N_27493,N_28145);
xnor U31224 (N_31224,N_26592,N_28704);
nor U31225 (N_31225,N_27676,N_25241);
or U31226 (N_31226,N_27119,N_25142);
or U31227 (N_31227,N_29206,N_26245);
nor U31228 (N_31228,N_25936,N_27523);
and U31229 (N_31229,N_26990,N_25888);
xnor U31230 (N_31230,N_29093,N_29703);
and U31231 (N_31231,N_28151,N_29643);
or U31232 (N_31232,N_29474,N_27487);
xnor U31233 (N_31233,N_27195,N_27605);
nand U31234 (N_31234,N_27295,N_28004);
xnor U31235 (N_31235,N_26661,N_27914);
and U31236 (N_31236,N_27375,N_25981);
or U31237 (N_31237,N_29869,N_26629);
xor U31238 (N_31238,N_29062,N_26801);
and U31239 (N_31239,N_25009,N_25590);
nor U31240 (N_31240,N_28929,N_26851);
nor U31241 (N_31241,N_26044,N_27679);
and U31242 (N_31242,N_25177,N_25354);
xnor U31243 (N_31243,N_26329,N_25378);
or U31244 (N_31244,N_28612,N_26898);
nor U31245 (N_31245,N_29758,N_29056);
nor U31246 (N_31246,N_28986,N_28134);
xnor U31247 (N_31247,N_28001,N_27466);
or U31248 (N_31248,N_26354,N_26608);
nor U31249 (N_31249,N_27729,N_29343);
nand U31250 (N_31250,N_25046,N_26609);
or U31251 (N_31251,N_27065,N_28169);
xnor U31252 (N_31252,N_26565,N_29800);
xnor U31253 (N_31253,N_25526,N_28984);
and U31254 (N_31254,N_27804,N_28263);
xnor U31255 (N_31255,N_28868,N_28124);
nand U31256 (N_31256,N_29297,N_26501);
nor U31257 (N_31257,N_25538,N_25087);
and U31258 (N_31258,N_25572,N_27185);
nand U31259 (N_31259,N_26537,N_25076);
and U31260 (N_31260,N_28362,N_25361);
xor U31261 (N_31261,N_29931,N_27895);
nor U31262 (N_31262,N_28771,N_27581);
nand U31263 (N_31263,N_26103,N_25587);
nor U31264 (N_31264,N_25259,N_27049);
xnor U31265 (N_31265,N_29246,N_28407);
or U31266 (N_31266,N_28746,N_27730);
nand U31267 (N_31267,N_29825,N_26177);
nor U31268 (N_31268,N_28791,N_29546);
or U31269 (N_31269,N_27764,N_25029);
or U31270 (N_31270,N_27564,N_26261);
or U31271 (N_31271,N_28533,N_25043);
nor U31272 (N_31272,N_27527,N_27822);
nand U31273 (N_31273,N_26967,N_28294);
nor U31274 (N_31274,N_26342,N_27807);
xor U31275 (N_31275,N_26286,N_26935);
nor U31276 (N_31276,N_28428,N_29983);
nor U31277 (N_31277,N_27872,N_28640);
xor U31278 (N_31278,N_29627,N_28983);
or U31279 (N_31279,N_28751,N_29484);
nand U31280 (N_31280,N_28559,N_29107);
xor U31281 (N_31281,N_29351,N_28512);
nor U31282 (N_31282,N_29736,N_28007);
nand U31283 (N_31283,N_29720,N_26272);
nand U31284 (N_31284,N_28935,N_25432);
or U31285 (N_31285,N_27810,N_25762);
xor U31286 (N_31286,N_25886,N_27905);
and U31287 (N_31287,N_26813,N_27470);
nor U31288 (N_31288,N_27153,N_27446);
xor U31289 (N_31289,N_26668,N_28847);
xnor U31290 (N_31290,N_29592,N_28237);
and U31291 (N_31291,N_29172,N_28229);
nand U31292 (N_31292,N_27425,N_28201);
xnor U31293 (N_31293,N_25524,N_28268);
nand U31294 (N_31294,N_27456,N_28186);
nor U31295 (N_31295,N_26061,N_29000);
nor U31296 (N_31296,N_26512,N_27598);
and U31297 (N_31297,N_25967,N_27979);
nor U31298 (N_31298,N_26545,N_29104);
nor U31299 (N_31299,N_29826,N_28250);
and U31300 (N_31300,N_29240,N_28086);
xor U31301 (N_31301,N_28240,N_26241);
nor U31302 (N_31302,N_29842,N_28257);
xnor U31303 (N_31303,N_27042,N_29153);
xor U31304 (N_31304,N_26816,N_25420);
xnor U31305 (N_31305,N_29114,N_28891);
nor U31306 (N_31306,N_25970,N_27680);
nand U31307 (N_31307,N_25848,N_27879);
or U31308 (N_31308,N_27714,N_25323);
or U31309 (N_31309,N_27017,N_27715);
or U31310 (N_31310,N_29666,N_25192);
or U31311 (N_31311,N_29388,N_25568);
nand U31312 (N_31312,N_26539,N_27489);
and U31313 (N_31313,N_29832,N_28311);
nand U31314 (N_31314,N_26663,N_29478);
and U31315 (N_31315,N_29746,N_28494);
xnor U31316 (N_31316,N_28698,N_28878);
or U31317 (N_31317,N_29454,N_25999);
or U31318 (N_31318,N_27066,N_29335);
and U31319 (N_31319,N_26236,N_25651);
xor U31320 (N_31320,N_27515,N_29112);
nor U31321 (N_31321,N_26404,N_29413);
or U31322 (N_31322,N_29663,N_28990);
nor U31323 (N_31323,N_25743,N_28170);
nor U31324 (N_31324,N_25525,N_28676);
nand U31325 (N_31325,N_27335,N_27815);
nand U31326 (N_31326,N_26107,N_26458);
and U31327 (N_31327,N_25796,N_28832);
and U31328 (N_31328,N_26513,N_27384);
and U31329 (N_31329,N_28999,N_25562);
and U31330 (N_31330,N_25166,N_29383);
or U31331 (N_31331,N_26417,N_27911);
xor U31332 (N_31332,N_28125,N_29076);
or U31333 (N_31333,N_26131,N_28210);
xor U31334 (N_31334,N_25582,N_27517);
and U31335 (N_31335,N_26226,N_25877);
xnor U31336 (N_31336,N_28285,N_29912);
nand U31337 (N_31337,N_27204,N_26302);
nor U31338 (N_31338,N_25745,N_27474);
nor U31339 (N_31339,N_26438,N_25362);
nor U31340 (N_31340,N_27143,N_25555);
and U31341 (N_31341,N_28073,N_25143);
or U31342 (N_31342,N_27953,N_25772);
nor U31343 (N_31343,N_26672,N_25829);
xor U31344 (N_31344,N_25552,N_27368);
nor U31345 (N_31345,N_27464,N_25200);
nand U31346 (N_31346,N_25683,N_25372);
nor U31347 (N_31347,N_27062,N_28183);
nor U31348 (N_31348,N_26472,N_27302);
nand U31349 (N_31349,N_28711,N_25990);
nand U31350 (N_31350,N_25718,N_25386);
or U31351 (N_31351,N_26247,N_27850);
nand U31352 (N_31352,N_25537,N_28258);
nand U31353 (N_31353,N_28078,N_29935);
nand U31354 (N_31354,N_29017,N_26675);
nor U31355 (N_31355,N_25826,N_28224);
and U31356 (N_31356,N_27180,N_28058);
or U31357 (N_31357,N_27970,N_27041);
or U31358 (N_31358,N_29894,N_26121);
and U31359 (N_31359,N_25124,N_29914);
or U31360 (N_31360,N_28858,N_25418);
or U31361 (N_31361,N_25392,N_27786);
xnor U31362 (N_31362,N_26887,N_28208);
nand U31363 (N_31363,N_26228,N_25039);
nand U31364 (N_31364,N_29880,N_25085);
nand U31365 (N_31365,N_25769,N_25056);
or U31366 (N_31366,N_29584,N_26370);
nand U31367 (N_31367,N_28625,N_29940);
or U31368 (N_31368,N_26530,N_25286);
or U31369 (N_31369,N_29994,N_25670);
or U31370 (N_31370,N_28796,N_28934);
nor U31371 (N_31371,N_29558,N_27219);
nor U31372 (N_31372,N_28737,N_28182);
nand U31373 (N_31373,N_27272,N_25334);
nor U31374 (N_31374,N_25351,N_27618);
or U31375 (N_31375,N_27318,N_28575);
and U31376 (N_31376,N_28794,N_26747);
or U31377 (N_31377,N_26773,N_29471);
or U31378 (N_31378,N_25125,N_29031);
xor U31379 (N_31379,N_27770,N_29400);
or U31380 (N_31380,N_27611,N_29642);
and U31381 (N_31381,N_26264,N_29566);
nand U31382 (N_31382,N_29862,N_26917);
or U31383 (N_31383,N_26279,N_27877);
nand U31384 (N_31384,N_26732,N_28198);
nand U31385 (N_31385,N_28571,N_28166);
and U31386 (N_31386,N_25921,N_27211);
nand U31387 (N_31387,N_27569,N_25342);
nand U31388 (N_31388,N_26875,N_26554);
xnor U31389 (N_31389,N_26987,N_27007);
xor U31390 (N_31390,N_27981,N_28757);
xnor U31391 (N_31391,N_27320,N_27593);
or U31392 (N_31392,N_28492,N_27140);
nand U31393 (N_31393,N_27883,N_29760);
xnor U31394 (N_31394,N_28129,N_28629);
nor U31395 (N_31395,N_25697,N_25750);
and U31396 (N_31396,N_27422,N_26938);
nor U31397 (N_31397,N_29913,N_28638);
nand U31398 (N_31398,N_27477,N_28296);
nand U31399 (N_31399,N_26389,N_29523);
and U31400 (N_31400,N_28907,N_29610);
xor U31401 (N_31401,N_26248,N_28995);
nor U31402 (N_31402,N_27268,N_27336);
or U31403 (N_31403,N_27882,N_29255);
or U31404 (N_31404,N_26701,N_28774);
nand U31405 (N_31405,N_28903,N_26288);
or U31406 (N_31406,N_29201,N_25050);
nor U31407 (N_31407,N_28149,N_26757);
and U31408 (N_31408,N_26363,N_27768);
or U31409 (N_31409,N_28710,N_25579);
xnor U31410 (N_31410,N_29366,N_25641);
and U31411 (N_31411,N_28881,N_25712);
nand U31412 (N_31412,N_28782,N_28320);
xor U31413 (N_31413,N_28389,N_28317);
xnor U31414 (N_31414,N_28960,N_25971);
nand U31415 (N_31415,N_28176,N_28923);
nand U31416 (N_31416,N_28054,N_28979);
xnor U31417 (N_31417,N_28083,N_25958);
nor U31418 (N_31418,N_26669,N_26750);
xor U31419 (N_31419,N_28467,N_26066);
and U31420 (N_31420,N_28387,N_26905);
nand U31421 (N_31421,N_28908,N_26060);
nor U31422 (N_31422,N_27186,N_25287);
xnor U31423 (N_31423,N_27959,N_25759);
or U31424 (N_31424,N_26913,N_26306);
nor U31425 (N_31425,N_25366,N_26373);
or U31426 (N_31426,N_29237,N_27833);
nor U31427 (N_31427,N_26457,N_29580);
nand U31428 (N_31428,N_28000,N_29749);
xnor U31429 (N_31429,N_28576,N_28653);
xor U31430 (N_31430,N_27550,N_26412);
or U31431 (N_31431,N_27933,N_27253);
and U31432 (N_31432,N_28998,N_25198);
and U31433 (N_31433,N_26507,N_26895);
nand U31434 (N_31434,N_25709,N_26477);
and U31435 (N_31435,N_27868,N_25982);
nor U31436 (N_31436,N_28902,N_26751);
nor U31437 (N_31437,N_28322,N_28988);
and U31438 (N_31438,N_25666,N_29279);
nand U31439 (N_31439,N_28776,N_29709);
and U31440 (N_31440,N_29485,N_26586);
nand U31441 (N_31441,N_28267,N_27193);
or U31442 (N_31442,N_27548,N_28880);
and U31443 (N_31443,N_27221,N_26977);
nor U31444 (N_31444,N_26104,N_27306);
xor U31445 (N_31445,N_27341,N_25910);
xor U31446 (N_31446,N_28060,N_29937);
nand U31447 (N_31447,N_27139,N_26340);
and U31448 (N_31448,N_26293,N_25685);
and U31449 (N_31449,N_28353,N_28122);
xnor U31450 (N_31450,N_28053,N_28046);
nor U31451 (N_31451,N_29853,N_26805);
nor U31452 (N_31452,N_27316,N_28011);
nor U31453 (N_31453,N_27996,N_28718);
or U31454 (N_31454,N_29033,N_25282);
and U31455 (N_31455,N_26638,N_29094);
and U31456 (N_31456,N_25973,N_29356);
nand U31457 (N_31457,N_25020,N_25131);
nand U31458 (N_31458,N_25116,N_27597);
xor U31459 (N_31459,N_27842,N_28910);
or U31460 (N_31460,N_25778,N_29559);
nor U31461 (N_31461,N_29836,N_29037);
nor U31462 (N_31462,N_26129,N_25815);
nor U31463 (N_31463,N_27669,N_29933);
and U31464 (N_31464,N_29863,N_28759);
nor U31465 (N_31465,N_29210,N_25793);
nor U31466 (N_31466,N_26139,N_29519);
nand U31467 (N_31467,N_29328,N_29867);
xnor U31468 (N_31468,N_29482,N_25673);
xor U31469 (N_31469,N_29823,N_27366);
or U31470 (N_31470,N_27198,N_28204);
nor U31471 (N_31471,N_25042,N_27777);
and U31472 (N_31472,N_25846,N_27251);
and U31473 (N_31473,N_27382,N_28816);
and U31474 (N_31474,N_27503,N_25707);
nor U31475 (N_31475,N_26165,N_29586);
or U31476 (N_31476,N_29888,N_29171);
nor U31477 (N_31477,N_26560,N_26309);
or U31478 (N_31478,N_26395,N_27991);
nand U31479 (N_31479,N_28818,N_25915);
nand U31480 (N_31480,N_26499,N_28254);
nor U31481 (N_31481,N_28217,N_26845);
or U31482 (N_31482,N_26800,N_25322);
nand U31483 (N_31483,N_27312,N_26164);
and U31484 (N_31484,N_28584,N_29339);
xnor U31485 (N_31485,N_27416,N_26931);
and U31486 (N_31486,N_28901,N_25038);
and U31487 (N_31487,N_28264,N_27518);
and U31488 (N_31488,N_28372,N_25875);
and U31489 (N_31489,N_27852,N_29312);
xor U31490 (N_31490,N_28439,N_26137);
nor U31491 (N_31491,N_28932,N_29218);
or U31492 (N_31492,N_26784,N_26758);
and U31493 (N_31493,N_28754,N_26379);
and U31494 (N_31494,N_26467,N_29966);
or U31495 (N_31495,N_25962,N_28388);
and U31496 (N_31496,N_25369,N_26962);
and U31497 (N_31497,N_29177,N_28860);
nor U31498 (N_31498,N_27876,N_26449);
or U31499 (N_31499,N_27032,N_29245);
xnor U31500 (N_31500,N_27273,N_27838);
or U31501 (N_31501,N_27849,N_25813);
or U31502 (N_31502,N_27788,N_27108);
nor U31503 (N_31503,N_29030,N_28764);
and U31504 (N_31504,N_28552,N_27586);
nor U31505 (N_31505,N_25013,N_25339);
xnor U31506 (N_31506,N_29520,N_27769);
xor U31507 (N_31507,N_29570,N_26557);
or U31508 (N_31508,N_28821,N_27165);
nand U31509 (N_31509,N_29809,N_27587);
or U31510 (N_31510,N_26427,N_25442);
or U31511 (N_31511,N_26317,N_27255);
or U31512 (N_31512,N_29156,N_27565);
xnor U31513 (N_31513,N_27314,N_29399);
nand U31514 (N_31514,N_27722,N_27956);
nor U31515 (N_31515,N_26028,N_26413);
nand U31516 (N_31516,N_25985,N_29597);
nor U31517 (N_31517,N_29152,N_25164);
nor U31518 (N_31518,N_29765,N_26252);
or U31519 (N_31519,N_29807,N_28331);
or U31520 (N_31520,N_27865,N_29946);
or U31521 (N_31521,N_26528,N_25061);
and U31522 (N_31522,N_26110,N_29023);
and U31523 (N_31523,N_27800,N_27397);
or U31524 (N_31524,N_29972,N_25527);
nor U31525 (N_31525,N_27583,N_25715);
nand U31526 (N_31526,N_26711,N_25370);
or U31527 (N_31527,N_25935,N_29071);
or U31528 (N_31528,N_25528,N_28489);
xnor U31529 (N_31529,N_29057,N_28020);
nand U31530 (N_31530,N_25343,N_26234);
nor U31531 (N_31531,N_26692,N_29976);
and U31532 (N_31532,N_26924,N_27666);
xor U31533 (N_31533,N_25704,N_29079);
nor U31534 (N_31534,N_29557,N_26717);
nor U31535 (N_31535,N_26274,N_25028);
xnor U31536 (N_31536,N_29902,N_27450);
nand U31537 (N_31537,N_25337,N_28158);
xnor U31538 (N_31538,N_29133,N_29008);
nor U31539 (N_31539,N_25300,N_28950);
and U31540 (N_31540,N_25648,N_27942);
or U31541 (N_31541,N_26628,N_27525);
or U31542 (N_31542,N_29624,N_29690);
and U31543 (N_31543,N_26152,N_27082);
and U31544 (N_31544,N_28136,N_29815);
xor U31545 (N_31545,N_29632,N_27289);
xnor U31546 (N_31546,N_25534,N_26151);
nor U31547 (N_31547,N_28333,N_28528);
xor U31548 (N_31548,N_26188,N_29444);
nand U31549 (N_31549,N_28856,N_26840);
nor U31550 (N_31550,N_28153,N_27132);
xnor U31551 (N_31551,N_26521,N_28121);
and U31552 (N_31552,N_26123,N_28249);
nand U31553 (N_31553,N_29512,N_25169);
nor U31554 (N_31554,N_25232,N_27075);
nand U31555 (N_31555,N_25833,N_28064);
xor U31556 (N_31556,N_28269,N_26111);
nor U31557 (N_31557,N_26680,N_25077);
nor U31558 (N_31558,N_26163,N_27452);
and U31559 (N_31559,N_27351,N_29145);
xnor U31560 (N_31560,N_25779,N_28522);
nand U31561 (N_31561,N_28375,N_29714);
xnor U31562 (N_31562,N_29810,N_29091);
and U31563 (N_31563,N_28349,N_26112);
or U31564 (N_31564,N_25141,N_25376);
or U31565 (N_31565,N_29657,N_27146);
nor U31566 (N_31566,N_26062,N_28547);
nand U31567 (N_31567,N_27287,N_29992);
xnor U31568 (N_31568,N_26787,N_26268);
nor U31569 (N_31569,N_28598,N_26802);
xor U31570 (N_31570,N_29235,N_29405);
nand U31571 (N_31571,N_27949,N_28066);
nor U31572 (N_31572,N_28973,N_29752);
and U31573 (N_31573,N_27276,N_29790);
or U31574 (N_31574,N_29250,N_27855);
nor U31575 (N_31575,N_29199,N_27342);
nand U31576 (N_31576,N_27801,N_26532);
or U31577 (N_31577,N_25988,N_29568);
or U31578 (N_31578,N_25353,N_27112);
and U31579 (N_31579,N_29915,N_28313);
or U31580 (N_31580,N_29685,N_26829);
xnor U31581 (N_31581,N_25976,N_27696);
nor U31582 (N_31582,N_25816,N_25919);
and U31583 (N_31583,N_28949,N_25591);
and U31584 (N_31584,N_28619,N_25021);
nor U31585 (N_31585,N_26242,N_26597);
xor U31586 (N_31586,N_28039,N_26195);
or U31587 (N_31587,N_29003,N_29493);
nand U31588 (N_31588,N_27719,N_29020);
and U31589 (N_31589,N_26269,N_27442);
nor U31590 (N_31590,N_28260,N_29494);
nor U31591 (N_31591,N_26273,N_28786);
nand U31592 (N_31592,N_29929,N_26908);
and U31593 (N_31593,N_28717,N_27494);
xor U31594 (N_31594,N_28243,N_26463);
xor U31595 (N_31595,N_26357,N_26673);
xor U31596 (N_31596,N_25912,N_25341);
nor U31597 (N_31597,N_29487,N_29289);
or U31598 (N_31598,N_29729,N_25199);
nor U31599 (N_31599,N_27741,N_26381);
and U31600 (N_31600,N_29340,N_29623);
xnor U31601 (N_31601,N_26852,N_28165);
xor U31602 (N_31602,N_26124,N_28622);
nand U31603 (N_31603,N_27182,N_29491);
and U31604 (N_31604,N_26715,N_25964);
nor U31605 (N_31605,N_26789,N_25879);
and U31606 (N_31606,N_25326,N_25456);
or U31607 (N_31607,N_29489,N_27500);
xor U31608 (N_31608,N_29182,N_28393);
nor U31609 (N_31609,N_29543,N_28896);
and U31610 (N_31610,N_27999,N_27014);
nor U31611 (N_31611,N_28738,N_25900);
and U31612 (N_31612,N_26392,N_29282);
nand U31613 (N_31613,N_27006,N_25231);
nand U31614 (N_31614,N_28316,N_29129);
nand U31615 (N_31615,N_26450,N_29231);
nand U31616 (N_31616,N_28342,N_25823);
nand U31617 (N_31617,N_26096,N_27026);
and U31618 (N_31618,N_27488,N_28003);
or U31619 (N_31619,N_26403,N_28994);
and U31620 (N_31620,N_26623,N_28789);
or U31621 (N_31621,N_27840,N_26594);
or U31622 (N_31622,N_26461,N_25189);
or U31623 (N_31623,N_26153,N_27115);
and U31624 (N_31624,N_29517,N_25500);
nor U31625 (N_31625,N_25649,N_25051);
and U31626 (N_31626,N_26900,N_26515);
nor U31627 (N_31627,N_28455,N_27380);
or U31628 (N_31628,N_26016,N_27886);
xor U31629 (N_31629,N_25546,N_27718);
or U31630 (N_31630,N_27497,N_29181);
xnor U31631 (N_31631,N_27224,N_29275);
nor U31632 (N_31632,N_27958,N_25462);
and U31633 (N_31633,N_26276,N_27455);
nand U31634 (N_31634,N_28377,N_29161);
nor U31635 (N_31635,N_26728,N_29698);
and U31636 (N_31636,N_29645,N_27926);
xnor U31637 (N_31637,N_28115,N_26089);
nor U31638 (N_31638,N_26504,N_25053);
nand U31639 (N_31639,N_27394,N_25419);
nor U31640 (N_31640,N_26880,N_25412);
xor U31641 (N_31641,N_27039,N_28660);
nor U31642 (N_31642,N_28748,N_26290);
xnor U31643 (N_31643,N_29678,N_25090);
nor U31644 (N_31644,N_28523,N_26618);
nand U31645 (N_31645,N_25071,N_28199);
nand U31646 (N_31646,N_27453,N_28766);
and U31647 (N_31647,N_28675,N_25122);
or U31648 (N_31648,N_27614,N_27444);
nand U31649 (N_31649,N_28431,N_25650);
nand U31650 (N_31650,N_28690,N_27937);
nand U31651 (N_31651,N_27424,N_25281);
or U31652 (N_31652,N_28207,N_26208);
nor U31653 (N_31653,N_28118,N_26769);
nand U31654 (N_31654,N_25276,N_28044);
nor U31655 (N_31655,N_26867,N_29347);
nand U31656 (N_31656,N_28223,N_27093);
and U31657 (N_31657,N_28931,N_27378);
nor U31658 (N_31658,N_25025,N_29767);
or U31659 (N_31659,N_27055,N_27117);
nand U31660 (N_31660,N_27774,N_25703);
nor U31661 (N_31661,N_25350,N_29434);
xor U31662 (N_31662,N_25247,N_25380);
nor U31663 (N_31663,N_27642,N_29034);
nand U31664 (N_31664,N_25311,N_26158);
nor U31665 (N_31665,N_29669,N_25083);
nor U31666 (N_31666,N_27809,N_26850);
nand U31667 (N_31667,N_26930,N_29728);
nand U31668 (N_31668,N_28566,N_29021);
nor U31669 (N_31669,N_29307,N_28033);
or U31670 (N_31670,N_27735,N_25305);
nand U31671 (N_31671,N_27252,N_25207);
nor U31672 (N_31672,N_27853,N_28644);
or U31673 (N_31673,N_25573,N_26476);
nor U31674 (N_31674,N_26971,N_25785);
and U31675 (N_31675,N_26951,N_27029);
nand U31676 (N_31676,N_29209,N_27344);
xnor U31677 (N_31677,N_28302,N_25273);
or U31678 (N_31678,N_25277,N_25398);
xor U31679 (N_31679,N_29358,N_25725);
nor U31680 (N_31680,N_26633,N_27929);
xor U31681 (N_31681,N_27812,N_26292);
xor U31682 (N_31682,N_25857,N_29044);
and U31683 (N_31683,N_26604,N_28674);
or U31684 (N_31684,N_25401,N_29169);
nand U31685 (N_31685,N_27603,N_25662);
nor U31686 (N_31686,N_26487,N_29131);
nor U31687 (N_31687,N_26257,N_29271);
nor U31688 (N_31688,N_29704,N_26570);
nand U31689 (N_31689,N_26233,N_25806);
nor U31690 (N_31690,N_29121,N_27875);
xnor U31691 (N_31691,N_29132,N_25145);
or U31692 (N_31692,N_27409,N_26263);
nor U31693 (N_31693,N_26283,N_27909);
xnor U31694 (N_31694,N_25296,N_26219);
nand U31695 (N_31695,N_27338,N_27088);
or U31696 (N_31696,N_25089,N_25885);
or U31697 (N_31697,N_29119,N_29783);
or U31698 (N_31698,N_27162,N_25414);
and U31699 (N_31699,N_26176,N_29724);
or U31700 (N_31700,N_27441,N_29221);
or U31701 (N_31701,N_29775,N_27473);
nor U31702 (N_31702,N_28959,N_29120);
xnor U31703 (N_31703,N_26316,N_29986);
and U31704 (N_31704,N_27974,N_29766);
nor U31705 (N_31705,N_29852,N_29080);
nand U31706 (N_31706,N_29938,N_29193);
or U31707 (N_31707,N_25506,N_29359);
nand U31708 (N_31708,N_26579,N_28608);
or U31709 (N_31709,N_27824,N_26553);
nor U31710 (N_31710,N_28972,N_26130);
or U31711 (N_31711,N_28065,N_29178);
and U31712 (N_31712,N_29113,N_26431);
or U31713 (N_31713,N_29944,N_29999);
and U31714 (N_31714,N_29665,N_25228);
xnor U31715 (N_31715,N_25202,N_26870);
and U31716 (N_31716,N_29261,N_29961);
or U31717 (N_31717,N_29725,N_29490);
or U31718 (N_31718,N_25509,N_28391);
nand U31719 (N_31719,N_27048,N_27577);
nor U31720 (N_31720,N_25989,N_27121);
xnor U31721 (N_31721,N_25549,N_27601);
nor U31722 (N_31722,N_26765,N_28032);
nor U31723 (N_31723,N_25293,N_29941);
xnor U31724 (N_31724,N_25270,N_27727);
xnor U31725 (N_31725,N_25290,N_25082);
nor U31726 (N_31726,N_26086,N_27046);
or U31727 (N_31727,N_27749,N_29950);
nor U31728 (N_31728,N_28899,N_26934);
and U31729 (N_31729,N_25539,N_27296);
nand U31730 (N_31730,N_28160,N_25748);
nand U31731 (N_31731,N_26865,N_26037);
and U31732 (N_31732,N_29283,N_25991);
nand U31733 (N_31733,N_27151,N_27559);
xor U31734 (N_31734,N_28189,N_25101);
nand U31735 (N_31735,N_29960,N_28946);
or U31736 (N_31736,N_25801,N_28515);
or U31737 (N_31737,N_25617,N_28104);
xnor U31738 (N_31738,N_25215,N_27590);
xor U31739 (N_31739,N_25520,N_27672);
nand U31740 (N_31740,N_26810,N_27430);
or U31741 (N_31741,N_26918,N_25406);
and U31742 (N_31742,N_29463,N_28076);
xnor U31743 (N_31743,N_25687,N_25285);
xnor U31744 (N_31744,N_29591,N_27846);
and U31745 (N_31745,N_29814,N_27391);
nor U31746 (N_31746,N_29313,N_28628);
nor U31747 (N_31747,N_25620,N_27277);
xor U31748 (N_31748,N_29955,N_27771);
nor U31749 (N_31749,N_28875,N_25080);
and U31750 (N_31750,N_27519,N_26568);
nand U31751 (N_31751,N_28889,N_27238);
and U31752 (N_31752,N_29018,N_27188);
or U31753 (N_31753,N_27168,N_28631);
nor U31754 (N_31754,N_29786,N_29441);
and U31755 (N_31755,N_25677,N_26031);
or U31756 (N_31756,N_25451,N_29995);
nand U31757 (N_31757,N_25208,N_27247);
or U31758 (N_31758,N_25217,N_28148);
xnor U31759 (N_31759,N_27721,N_27410);
nand U31760 (N_31760,N_25925,N_27816);
or U31761 (N_31761,N_28424,N_27779);
and U31762 (N_31762,N_28468,N_28634);
xor U31763 (N_31763,N_26807,N_26076);
and U31764 (N_31764,N_27685,N_25439);
xor U31765 (N_31765,N_29109,N_28139);
nor U31766 (N_31766,N_29222,N_26071);
and U31767 (N_31767,N_25663,N_29572);
xor U31768 (N_31768,N_26180,N_27825);
xnor U31769 (N_31769,N_26808,N_25470);
and U31770 (N_31770,N_27568,N_27516);
xor U31771 (N_31771,N_26070,N_28504);
and U31772 (N_31772,N_25203,N_28841);
nand U31773 (N_31773,N_28637,N_27071);
or U31774 (N_31774,N_27656,N_27835);
nand U31775 (N_31775,N_29393,N_26578);
nor U31776 (N_31776,N_25551,N_28295);
and U31777 (N_31777,N_27301,N_29845);
nand U31778 (N_31778,N_28344,N_25034);
nor U31779 (N_31779,N_27863,N_29906);
or U31780 (N_31780,N_28708,N_26084);
xnor U31781 (N_31781,N_28366,N_26610);
or U31782 (N_31782,N_27184,N_28633);
and U31783 (N_31783,N_27983,N_29390);
xnor U31784 (N_31784,N_28290,N_27271);
nand U31785 (N_31785,N_29294,N_28080);
or U31786 (N_31786,N_26738,N_25385);
and U31787 (N_31787,N_27682,N_26384);
nand U31788 (N_31788,N_27432,N_28460);
xnor U31789 (N_31789,N_25130,N_28564);
nand U31790 (N_31790,N_26326,N_29738);
or U31791 (N_31791,N_29083,N_26963);
xor U31792 (N_31792,N_25234,N_29599);
nor U31793 (N_31793,N_29443,N_25460);
nand U31794 (N_31794,N_29090,N_25183);
and U31795 (N_31795,N_29877,N_28184);
xnor U31796 (N_31796,N_28663,N_26825);
nand U31797 (N_31797,N_29286,N_29292);
nand U31798 (N_31798,N_26497,N_25997);
nor U31799 (N_31799,N_25625,N_26364);
nand U31800 (N_31800,N_26216,N_26725);
or U31801 (N_31801,N_29211,N_26231);
nand U31802 (N_31802,N_27013,N_25932);
nor U31803 (N_31803,N_26298,N_28470);
xor U31804 (N_31804,N_28173,N_29060);
nand U31805 (N_31805,N_28114,N_28658);
nor U31806 (N_31806,N_26125,N_29870);
xnor U31807 (N_31807,N_25346,N_27157);
or U31808 (N_31808,N_26224,N_27206);
xnor U31809 (N_31809,N_25810,N_28410);
nand U31810 (N_31810,N_29073,N_25359);
xnor U31811 (N_31811,N_27707,N_29481);
nand U31812 (N_31812,N_25838,N_28541);
and U31813 (N_31813,N_27808,N_29305);
and U31814 (N_31814,N_26003,N_26549);
nand U31815 (N_31815,N_29716,N_28924);
nand U31816 (N_31816,N_25987,N_28397);
or U31817 (N_31817,N_28094,N_29375);
and U31818 (N_31818,N_29397,N_25916);
or U31819 (N_31819,N_26334,N_28815);
or U31820 (N_31820,N_25355,N_26759);
xor U31821 (N_31821,N_28197,N_28756);
xnor U31822 (N_31822,N_26132,N_29127);
nor U31823 (N_31823,N_29213,N_27687);
or U31824 (N_31824,N_28969,N_25045);
or U31825 (N_31825,N_29829,N_26083);
and U31826 (N_31826,N_25901,N_26647);
xor U31827 (N_31827,N_28814,N_25485);
and U31828 (N_31828,N_28325,N_27698);
nand U31829 (N_31829,N_28350,N_29138);
nand U31830 (N_31830,N_27924,N_27021);
xor U31831 (N_31831,N_28887,N_25714);
or U31832 (N_31832,N_28873,N_29081);
nor U31833 (N_31833,N_25550,N_26193);
nor U31834 (N_31834,N_27495,N_29850);
xnor U31835 (N_31835,N_26362,N_27902);
nor U31836 (N_31836,N_28536,N_26712);
xor U31837 (N_31837,N_26353,N_28023);
nor U31838 (N_31838,N_29868,N_26108);
or U31839 (N_31839,N_25452,N_28599);
nor U31840 (N_31840,N_25491,N_29582);
nand U31841 (N_31841,N_25004,N_27309);
and U31842 (N_31842,N_29446,N_29149);
or U31843 (N_31843,N_26375,N_28163);
or U31844 (N_31844,N_28684,N_29851);
and U31845 (N_31845,N_26045,N_26667);
nor U31846 (N_31846,N_28085,N_29408);
or U31847 (N_31847,N_27189,N_25513);
or U31848 (N_31848,N_26173,N_27390);
nand U31849 (N_31849,N_26517,N_28485);
xor U31850 (N_31850,N_27700,N_26026);
nor U31851 (N_31851,N_28215,N_25109);
xor U31852 (N_31852,N_26387,N_28524);
or U31853 (N_31853,N_27663,N_25870);
or U31854 (N_31854,N_29438,N_29713);
nand U31855 (N_31855,N_28919,N_28558);
nor U31856 (N_31856,N_28769,N_28890);
or U31857 (N_31857,N_28610,N_26391);
xnor U31858 (N_31858,N_25279,N_26222);
nor U31859 (N_31859,N_27951,N_25239);
nor U31860 (N_31860,N_28252,N_28943);
nand U31861 (N_31861,N_27599,N_29948);
nor U31862 (N_31862,N_27449,N_28944);
nor U31863 (N_31863,N_25091,N_29192);
nor U31864 (N_31864,N_25892,N_26349);
and U31865 (N_31865,N_26600,N_29804);
xnor U31866 (N_31866,N_28987,N_29819);
xnor U31867 (N_31867,N_27402,N_28451);
or U31868 (N_31868,N_26815,N_29254);
or U31869 (N_31869,N_26004,N_28686);
xor U31870 (N_31870,N_29872,N_29672);
and U31871 (N_31871,N_26200,N_25949);
or U31872 (N_31872,N_28725,N_25074);
and U31873 (N_31873,N_26262,N_27641);
nor U31874 (N_31874,N_28588,N_29320);
and U31875 (N_31875,N_28734,N_29701);
nand U31876 (N_31876,N_28664,N_29743);
and U31877 (N_31877,N_27878,N_25682);
or U31878 (N_31878,N_27778,N_27935);
or U31879 (N_31879,N_29381,N_25904);
or U31880 (N_31880,N_28824,N_26255);
and U31881 (N_31881,N_28852,N_28897);
and U31882 (N_31882,N_27582,N_26117);
or U31883 (N_31883,N_29146,N_25856);
nand U31884 (N_31884,N_28669,N_27229);
or U31885 (N_31885,N_28014,N_25754);
or U31886 (N_31886,N_29883,N_25079);
and U31887 (N_31887,N_27790,N_28195);
and U31888 (N_31888,N_29882,N_29174);
nand U31889 (N_31889,N_29973,N_29416);
and U31890 (N_31890,N_25204,N_27035);
xor U31891 (N_31891,N_27930,N_25645);
xor U31892 (N_31892,N_29529,N_26411);
xnor U31893 (N_31893,N_29607,N_27018);
and U31894 (N_31894,N_26699,N_29707);
xor U31895 (N_31895,N_25294,N_26189);
and U31896 (N_31896,N_25992,N_29189);
xnor U31897 (N_31897,N_28797,N_28161);
nor U31898 (N_31898,N_27541,N_27090);
xor U31899 (N_31899,N_28862,N_27866);
and U31900 (N_31900,N_26529,N_26760);
xor U31901 (N_31901,N_29357,N_26823);
nor U31902 (N_31902,N_26483,N_28087);
nand U31903 (N_31903,N_29708,N_27070);
or U31904 (N_31904,N_25567,N_25508);
or U31905 (N_31905,N_25803,N_29136);
nand U31906 (N_31906,N_29963,N_27549);
and U31907 (N_31907,N_28339,N_28284);
nor U31908 (N_31908,N_26849,N_25802);
nor U31909 (N_31909,N_29637,N_29042);
nand U31910 (N_31910,N_25410,N_28716);
nand U31911 (N_31911,N_26861,N_29530);
xnor U31912 (N_31912,N_29195,N_27511);
nor U31913 (N_31913,N_28445,N_28071);
and U31914 (N_31914,N_26839,N_28980);
or U31915 (N_31915,N_29997,N_26047);
nor U31916 (N_31916,N_25211,N_25944);
xor U31917 (N_31917,N_29689,N_26679);
and U31918 (N_31918,N_26926,N_25280);
or U31919 (N_31919,N_25298,N_29051);
nor U31920 (N_31920,N_27683,N_29792);
xor U31921 (N_31921,N_28974,N_26402);
nor U31922 (N_31922,N_26920,N_27652);
and U31923 (N_31923,N_26394,N_28835);
nand U31924 (N_31924,N_29731,N_27163);
and U31925 (N_31925,N_28477,N_28920);
xor U31926 (N_31926,N_26433,N_25309);
nand U31927 (N_31927,N_27328,N_25434);
or U31928 (N_31928,N_25219,N_28244);
or U31929 (N_31929,N_28277,N_27201);
nand U31930 (N_31930,N_26032,N_26182);
xor U31931 (N_31931,N_28811,N_28100);
and U31932 (N_31932,N_25729,N_26223);
xnor U31933 (N_31933,N_28967,N_28654);
nand U31934 (N_31934,N_29841,N_28412);
or U31935 (N_31935,N_27633,N_25260);
xor U31936 (N_31936,N_29026,N_28549);
nand U31937 (N_31937,N_27621,N_26186);
nor U31938 (N_31938,N_26778,N_26893);
xor U31939 (N_31939,N_27612,N_27563);
nand U31940 (N_31940,N_29198,N_28068);
and U31941 (N_31941,N_29456,N_29722);
xnor U31942 (N_31942,N_29649,N_27543);
nand U31943 (N_31943,N_28405,N_27553);
xnor U31944 (N_31944,N_25097,N_25767);
nor U31945 (N_31945,N_25849,N_25554);
and U31946 (N_31946,N_26426,N_26090);
or U31947 (N_31947,N_29796,N_29353);
nand U31948 (N_31948,N_29277,N_29886);
nand U31949 (N_31949,N_25644,N_26352);
and U31950 (N_31950,N_27860,N_28893);
and U31951 (N_31951,N_27910,N_26902);
xor U31952 (N_31952,N_29064,N_28012);
nor U31953 (N_31953,N_28035,N_25737);
nor U31954 (N_31954,N_29802,N_29617);
xor U31955 (N_31955,N_29176,N_28351);
xor U31956 (N_31956,N_27024,N_25499);
or U31957 (N_31957,N_26380,N_28647);
nand U31958 (N_31958,N_27040,N_27483);
xnor U31959 (N_31959,N_25727,N_28795);
nor U31960 (N_31960,N_28542,N_26958);
or U31961 (N_31961,N_28785,N_29460);
or U31962 (N_31962,N_27144,N_26183);
nor U31963 (N_31963,N_27127,N_29424);
nand U31964 (N_31964,N_25842,N_29603);
xnor U31965 (N_31965,N_27147,N_25941);
and U31966 (N_31966,N_27008,N_25618);
and U31967 (N_31967,N_26631,N_28529);
or U31968 (N_31968,N_28497,N_25642);
or U31969 (N_31969,N_26368,N_28773);
nor U31970 (N_31970,N_26858,N_25947);
or U31971 (N_31971,N_28291,N_27364);
xnor U31972 (N_31972,N_29893,N_29680);
or U31973 (N_31973,N_28526,N_29220);
nand U31974 (N_31974,N_25706,N_25138);
xnor U31975 (N_31975,N_27638,N_29498);
xnor U31976 (N_31976,N_28701,N_29251);
xor U31977 (N_31977,N_26656,N_25172);
xor U31978 (N_31978,N_25679,N_25433);
nand U31979 (N_31979,N_29742,N_25889);
xnor U31980 (N_31980,N_26888,N_28029);
or U31981 (N_31981,N_27492,N_28228);
xor U31982 (N_31982,N_29620,N_28055);
or U31983 (N_31983,N_28514,N_27130);
or U31984 (N_31984,N_25914,N_26915);
nand U31985 (N_31985,N_28286,N_29302);
nand U31986 (N_31986,N_29452,N_29569);
and U31987 (N_31987,N_28454,N_27717);
xnor U31988 (N_31988,N_27098,N_29330);
xnor U31989 (N_31989,N_25627,N_26516);
nor U31990 (N_31990,N_29374,N_26017);
and U31991 (N_31991,N_25850,N_25751);
and U31992 (N_31992,N_29756,N_27755);
xor U31993 (N_31993,N_26942,N_27789);
and U31994 (N_31994,N_29061,N_26700);
nand U31995 (N_31995,N_26080,N_29179);
nand U31996 (N_31996,N_25344,N_28373);
nor U31997 (N_31997,N_28484,N_29667);
or U31998 (N_31998,N_26213,N_26925);
nor U31999 (N_31999,N_27692,N_26069);
xnor U32000 (N_32000,N_28568,N_27643);
xor U32001 (N_32001,N_27798,N_25188);
nand U32002 (N_32002,N_29166,N_27705);
nor U32003 (N_32003,N_29687,N_28516);
xnor U32004 (N_32004,N_25898,N_26064);
or U32005 (N_32005,N_29264,N_29338);
nor U32006 (N_32006,N_28981,N_27947);
and U32007 (N_32007,N_25377,N_27640);
nor U32008 (N_32008,N_26414,N_27173);
xor U32009 (N_32009,N_29325,N_26746);
or U32010 (N_32010,N_28602,N_26312);
xor U32011 (N_32011,N_29816,N_26171);
nand U32012 (N_32012,N_25599,N_27427);
or U32013 (N_32013,N_27693,N_26536);
xor U32014 (N_32014,N_29539,N_27331);
or U32015 (N_32015,N_28396,N_26227);
nor U32016 (N_32016,N_28042,N_29429);
nand U32017 (N_32017,N_26136,N_29197);
xnor U32018 (N_32018,N_26295,N_25133);
or U32019 (N_32019,N_27837,N_29419);
xnor U32020 (N_32020,N_29284,N_26745);
xnor U32021 (N_32021,N_28556,N_29575);
xnor U32022 (N_32022,N_26956,N_29170);
nand U32023 (N_32023,N_25960,N_29750);
nor U32024 (N_32024,N_26067,N_27097);
nor U32025 (N_32025,N_25517,N_29556);
or U32026 (N_32026,N_29116,N_27532);
xor U32027 (N_32027,N_29395,N_25636);
nand U32028 (N_32028,N_29622,N_28506);
and U32029 (N_32029,N_25115,N_25993);
xnor U32030 (N_32030,N_28976,N_27031);
nand U32031 (N_32031,N_28324,N_26249);
or U32032 (N_32032,N_28613,N_25593);
nor U32033 (N_32033,N_25489,N_27940);
and U32034 (N_32034,N_26484,N_27079);
nor U32035 (N_32035,N_29278,N_28402);
nand U32036 (N_32036,N_28433,N_25984);
or U32037 (N_32037,N_25713,N_25675);
nor U32038 (N_32038,N_26975,N_29855);
xor U32039 (N_32039,N_26654,N_27078);
nand U32040 (N_32040,N_26542,N_29095);
nor U32041 (N_32041,N_28892,N_29439);
nor U32042 (N_32042,N_29431,N_28936);
xor U32043 (N_32043,N_26986,N_29262);
nand U32044 (N_32044,N_28703,N_26097);
xor U32045 (N_32045,N_28057,N_25453);
and U32046 (N_32046,N_28481,N_27594);
xnor U32047 (N_32047,N_25405,N_28857);
or U32048 (N_32048,N_28491,N_26013);
and U32049 (N_32049,N_28103,N_28354);
xnor U32050 (N_32050,N_28715,N_29618);
or U32051 (N_32051,N_27738,N_28926);
or U32052 (N_32052,N_27217,N_28175);
or U32053 (N_32053,N_27609,N_26989);
xnor U32054 (N_32054,N_26068,N_25521);
nor U32055 (N_32055,N_27646,N_26534);
xor U32056 (N_32056,N_26109,N_28745);
and U32057 (N_32057,N_27254,N_27796);
nor U32058 (N_32058,N_29524,N_26665);
nor U32059 (N_32059,N_28255,N_26050);
nand U32060 (N_32060,N_25930,N_29252);
or U32061 (N_32061,N_26703,N_27567);
xor U32062 (N_32062,N_25795,N_26564);
nor U32063 (N_32063,N_25957,N_28132);
and U32064 (N_32064,N_28399,N_26614);
and U32065 (N_32065,N_29697,N_29806);
xnor U32066 (N_32066,N_26478,N_29918);
nor U32067 (N_32067,N_26550,N_27485);
nand U32068 (N_32068,N_25258,N_29730);
nor U32069 (N_32069,N_25032,N_27552);
nand U32070 (N_32070,N_29135,N_29386);
and U32071 (N_32071,N_26145,N_26922);
or U32072 (N_32072,N_28927,N_25571);
nor U32073 (N_32073,N_28253,N_27632);
xor U32074 (N_32074,N_29522,N_25920);
and U32075 (N_32075,N_28304,N_29762);
or U32076 (N_32076,N_26671,N_27658);
or U32077 (N_32077,N_27536,N_26957);
or U32078 (N_32078,N_29651,N_26299);
or U32079 (N_32079,N_28554,N_28527);
or U32080 (N_32080,N_29671,N_28017);
and U32081 (N_32081,N_29421,N_27823);
or U32082 (N_32082,N_25040,N_28537);
and U32083 (N_32083,N_25463,N_29795);
nand U32084 (N_32084,N_26637,N_26939);
or U32085 (N_32085,N_28251,N_26148);
nand U32086 (N_32086,N_25099,N_29370);
and U32087 (N_32087,N_27530,N_28459);
and U32088 (N_32088,N_28074,N_26100);
xnor U32089 (N_32089,N_29445,N_28138);
or U32090 (N_32090,N_28627,N_27723);
and U32091 (N_32091,N_28968,N_27813);
and U32092 (N_32092,N_25149,N_29606);
nand U32093 (N_32093,N_28370,N_25584);
or U32094 (N_32094,N_29010,N_26621);
and U32095 (N_32095,N_27056,N_29650);
xor U32096 (N_32096,N_27671,N_26305);
nand U32097 (N_32097,N_25730,N_25448);
nor U32098 (N_32098,N_29212,N_28614);
and U32099 (N_32099,N_26198,N_28452);
nor U32100 (N_32100,N_28288,N_28798);
xnor U32101 (N_32101,N_26936,N_26980);
xor U32102 (N_32102,N_28869,N_28803);
nor U32103 (N_32103,N_27904,N_27968);
nor U32104 (N_32104,N_26178,N_28443);
nand U32105 (N_32105,N_25977,N_25776);
and U32106 (N_32106,N_28997,N_25834);
and U32107 (N_32107,N_27896,N_28511);
xnor U32108 (N_32108,N_26736,N_27508);
and U32109 (N_32109,N_26572,N_29634);
xor U32110 (N_32110,N_25495,N_29072);
or U32111 (N_32111,N_26927,N_28414);
or U32112 (N_32112,N_25075,N_28109);
nand U32113 (N_32113,N_27190,N_27479);
and U32114 (N_32114,N_29022,N_26157);
and U32115 (N_32115,N_26842,N_25866);
nand U32116 (N_32116,N_26337,N_27686);
xor U32117 (N_32117,N_29784,N_29764);
or U32118 (N_32118,N_28276,N_27158);
nand U32119 (N_32119,N_27388,N_29847);
nor U32120 (N_32120,N_26682,N_27468);
nand U32121 (N_32121,N_29957,N_27639);
or U32122 (N_32122,N_29990,N_28172);
nand U32123 (N_32123,N_28607,N_29549);
nand U32124 (N_32124,N_26058,N_29518);
nand U32125 (N_32125,N_29682,N_27278);
or U32126 (N_32126,N_25394,N_29916);
and U32127 (N_32127,N_25017,N_25331);
or U32128 (N_32128,N_27114,N_25746);
nor U32129 (N_32129,N_26444,N_28425);
or U32130 (N_32130,N_28963,N_29785);
or U32131 (N_32131,N_27931,N_29789);
and U32132 (N_32132,N_28266,N_28574);
or U32133 (N_32133,N_27392,N_29309);
xor U32134 (N_32134,N_27413,N_25939);
or U32135 (N_32135,N_27281,N_25504);
xnor U32136 (N_32136,N_28671,N_26698);
and U32137 (N_32137,N_26181,N_29911);
nand U32138 (N_32138,N_28509,N_27551);
xor U32139 (N_32139,N_28478,N_27710);
xor U32140 (N_32140,N_28090,N_28792);
or U32141 (N_32141,N_29479,N_28188);
and U32142 (N_32142,N_27901,N_29901);
and U32143 (N_32143,N_29528,N_26301);
xor U32144 (N_32144,N_28392,N_27293);
nor U32145 (N_32145,N_28925,N_28620);
xor U32146 (N_32146,N_27218,N_27367);
xor U32147 (N_32147,N_27726,N_28834);
nand U32148 (N_32148,N_27655,N_26872);
nor U32149 (N_32149,N_27355,N_27321);
nand U32150 (N_32150,N_29705,N_25010);
or U32151 (N_32151,N_28777,N_29239);
xnor U32152 (N_32152,N_28272,N_26785);
nand U32153 (N_32153,N_29619,N_25887);
nand U32154 (N_32154,N_27545,N_29661);
nand U32155 (N_32155,N_27326,N_29013);
or U32156 (N_32156,N_26981,N_28282);
xor U32157 (N_32157,N_25209,N_28421);
xnor U32158 (N_32158,N_29266,N_28045);
xnor U32159 (N_32159,N_27857,N_25994);
and U32160 (N_32160,N_28034,N_26798);
or U32161 (N_32161,N_27776,N_26998);
or U32162 (N_32162,N_28740,N_29469);
xor U32163 (N_32163,N_27921,N_25792);
nand U32164 (N_32164,N_26267,N_26126);
nor U32165 (N_32165,N_29422,N_29903);
and U32166 (N_32166,N_25444,N_28359);
nand U32167 (N_32167,N_26356,N_28200);
nand U32168 (N_32168,N_27159,N_29059);
xor U32169 (N_32169,N_26214,N_25428);
or U32170 (N_32170,N_28239,N_29451);
nand U32171 (N_32171,N_27122,N_26057);
nand U32172 (N_32172,N_25140,N_26285);
nor U32173 (N_32173,N_29771,N_25391);
xor U32174 (N_32174,N_27681,N_28603);
or U32175 (N_32175,N_27604,N_29115);
and U32176 (N_32176,N_25622,N_26835);
and U32177 (N_32177,N_26232,N_26894);
nand U32178 (N_32178,N_28440,N_28271);
xnor U32179 (N_32179,N_25728,N_26488);
xor U32180 (N_32180,N_26042,N_26156);
or U32181 (N_32181,N_26775,N_28135);
and U32182 (N_32182,N_26678,N_26087);
nand U32183 (N_32183,N_29362,N_25847);
or U32184 (N_32184,N_29544,N_29188);
nor U32185 (N_32185,N_28591,N_27457);
or U32186 (N_32186,N_29921,N_25049);
and U32187 (N_32187,N_26972,N_25269);
nand U32188 (N_32188,N_25633,N_29942);
nand U32189 (N_32189,N_29977,N_26382);
nor U32190 (N_32190,N_26941,N_25996);
nand U32191 (N_32191,N_26018,N_26713);
and U32192 (N_32192,N_29310,N_26749);
xor U32193 (N_32193,N_26146,N_26556);
and U32194 (N_32194,N_25254,N_26244);
nand U32195 (N_32195,N_26313,N_26843);
or U32196 (N_32196,N_28755,N_28030);
nor U32197 (N_32197,N_25227,N_29777);
or U32198 (N_32198,N_27526,N_25575);
nand U32199 (N_32199,N_29587,N_28358);
and U32200 (N_32200,N_26239,N_26973);
nor U32201 (N_32201,N_28749,N_25423);
nor U32202 (N_32202,N_28544,N_29626);
nand U32203 (N_32203,N_28915,N_29654);
xor U32204 (N_32204,N_26398,N_25430);
nor U32205 (N_32205,N_26855,N_26468);
and U32206 (N_32206,N_27156,N_25086);
nand U32207 (N_32207,N_29545,N_29187);
and U32208 (N_32208,N_27712,N_25358);
xor U32209 (N_32209,N_28861,N_29360);
or U32210 (N_32210,N_25632,N_28009);
nand U32211 (N_32211,N_27103,N_26122);
nand U32212 (N_32212,N_29232,N_26804);
and U32213 (N_32213,N_29253,N_26333);
and U32214 (N_32214,N_25859,N_25764);
nor U32215 (N_32215,N_26960,N_26602);
xnor U32216 (N_32216,N_25665,N_25798);
and U32217 (N_32217,N_26734,N_27504);
xor U32218 (N_32218,N_25831,N_26012);
and U32219 (N_32219,N_26447,N_26094);
and U32220 (N_32220,N_25566,N_29745);
nand U32221 (N_32221,N_29616,N_29710);
xor U32222 (N_32222,N_28900,N_25382);
xor U32223 (N_32223,N_25516,N_27684);
and U32224 (N_32224,N_25861,N_27653);
and U32225 (N_32225,N_29088,N_26134);
nand U32226 (N_32226,N_25137,N_26324);
xnor U32227 (N_32227,N_27744,N_28496);
or U32228 (N_32228,N_27978,N_27558);
xor U32229 (N_32229,N_25518,N_27022);
or U32230 (N_32230,N_27175,N_25974);
nor U32231 (N_32231,N_26890,N_29969);
or U32232 (N_32232,N_26116,N_28914);
and U32233 (N_32233,N_29333,N_29150);
nand U32234 (N_32234,N_27821,N_27016);
xnor U32235 (N_32235,N_27791,N_25251);
nor U32236 (N_32236,N_25493,N_26622);
xnor U32237 (N_32237,N_28855,N_27753);
xnor U32238 (N_32238,N_25073,N_27555);
xnor U32239 (N_32239,N_26705,N_25335);
nand U32240 (N_32240,N_26470,N_25388);
or U32241 (N_32241,N_25163,N_27148);
or U32242 (N_32242,N_25869,N_25588);
or U32243 (N_32243,N_29945,N_27695);
nand U32244 (N_32244,N_28116,N_25147);
nor U32245 (N_32245,N_28474,N_26141);
nand U32246 (N_32246,N_26714,N_28877);
nor U32247 (N_32247,N_27851,N_29006);
and U32248 (N_32248,N_29638,N_28580);
nor U32249 (N_32249,N_29985,N_25614);
nand U32250 (N_32250,N_29230,N_26258);
or U32251 (N_32251,N_25852,N_29585);
xor U32252 (N_32252,N_26964,N_28476);
xor U32253 (N_32253,N_27743,N_28952);
or U32254 (N_32254,N_27239,N_25695);
xnor U32255 (N_32255,N_29352,N_26220);
and U32256 (N_32256,N_28837,N_28472);
or U32257 (N_32257,N_27135,N_29542);
nor U32258 (N_32258,N_27120,N_29930);
nor U32259 (N_32259,N_28539,N_28970);
or U32260 (N_32260,N_28390,N_29833);
and U32261 (N_32261,N_26901,N_26615);
and U32262 (N_32262,N_27972,N_27086);
and U32263 (N_32263,N_28955,N_29753);
nand U32264 (N_32264,N_25501,N_26911);
xor U32265 (N_32265,N_27724,N_27767);
nor U32266 (N_32266,N_28807,N_28206);
nand U32267 (N_32267,N_28449,N_25763);
xor U32268 (N_32268,N_26466,N_29608);
xnor U32269 (N_32269,N_29951,N_26102);
xor U32270 (N_32270,N_27757,N_28196);
nand U32271 (N_32271,N_27773,N_28735);
xor U32272 (N_32272,N_29849,N_25333);
nand U32273 (N_32273,N_29035,N_27322);
and U32274 (N_32274,N_27196,N_25601);
nand U32275 (N_32275,N_27817,N_29162);
xnor U32276 (N_32276,N_28209,N_25373);
or U32277 (N_32277,N_27116,N_26906);
nor U32278 (N_32278,N_27187,N_26319);
and U32279 (N_32279,N_25454,N_27136);
or U32280 (N_32280,N_26238,N_26015);
nand U32281 (N_32281,N_25758,N_27109);
nor U32282 (N_32282,N_29598,N_28101);
nand U32283 (N_32283,N_29001,N_25853);
nand U32284 (N_32284,N_27946,N_29805);
xor U32285 (N_32285,N_25876,N_25100);
nand U32286 (N_32286,N_27610,N_27360);
xor U32287 (N_32287,N_25553,N_28335);
xor U32288 (N_32288,N_29513,N_29139);
and U32289 (N_32289,N_25710,N_25397);
and U32290 (N_32290,N_27243,N_29029);
xnor U32291 (N_32291,N_28346,N_27387);
xnor U32292 (N_32292,N_29702,N_27137);
xnor U32293 (N_32293,N_25308,N_25390);
and U32294 (N_32294,N_27490,N_29229);
xnor U32295 (N_32295,N_28876,N_25749);
nor U32296 (N_32296,N_26494,N_29414);
or U32297 (N_32297,N_29573,N_28538);
or U32298 (N_32298,N_26575,N_27169);
nor U32299 (N_32299,N_26991,N_29711);
nor U32300 (N_32300,N_29611,N_29025);
nor U32301 (N_32301,N_26114,N_29055);
or U32302 (N_32302,N_28895,N_25078);
nor U32303 (N_32303,N_28084,N_29774);
or U32304 (N_32304,N_25871,N_29106);
and U32305 (N_32305,N_26314,N_27478);
xor U32306 (N_32306,N_26767,N_27990);
or U32307 (N_32307,N_27847,N_29024);
nand U32308 (N_32308,N_27250,N_28117);
and U32309 (N_32309,N_25330,N_27562);
or U32310 (N_32310,N_25019,N_29970);
nand U32311 (N_32311,N_29793,N_29349);
xor U32312 (N_32312,N_26420,N_25483);
nand U32313 (N_32313,N_28709,N_25399);
nor U32314 (N_32314,N_26161,N_27178);
nand U32315 (N_32315,N_29647,N_29084);
xor U32316 (N_32316,N_29779,N_25114);
and U32317 (N_32317,N_28624,N_27670);
or U32318 (N_32318,N_25387,N_27372);
nor U32319 (N_32319,N_29028,N_25583);
and U32320 (N_32320,N_28677,N_25307);
or U32321 (N_32321,N_26054,N_27977);
xnor U32322 (N_32322,N_25768,N_26969);
xnor U32323 (N_32323,N_25569,N_29258);
nor U32324 (N_32324,N_25186,N_25316);
xnor U32325 (N_32325,N_28507,N_25467);
xor U32326 (N_32326,N_28585,N_29535);
nor U32327 (N_32327,N_27811,N_29074);
and U32328 (N_32328,N_29105,N_27089);
xnor U32329 (N_32329,N_26793,N_25340);
nand U32330 (N_32330,N_29691,N_25048);
or U32331 (N_32331,N_25595,N_26372);
xnor U32332 (N_32332,N_29684,N_29908);
and U32333 (N_32333,N_28486,N_25031);
and U32334 (N_32334,N_28780,N_29385);
or U32335 (N_32335,N_25435,N_25014);
or U32336 (N_32336,N_25674,N_25733);
xnor U32337 (N_32337,N_25257,N_26446);
xnor U32338 (N_32338,N_28126,N_29101);
nor U32339 (N_32339,N_27299,N_29190);
or U32340 (N_32340,N_27179,N_28385);
nand U32341 (N_32341,N_26428,N_25507);
xor U32342 (N_32342,N_27528,N_25092);
xnor U32343 (N_32343,N_25081,N_25609);
and U32344 (N_32344,N_29435,N_26437);
xnor U32345 (N_32345,N_29952,N_27720);
and U32346 (N_32346,N_27619,N_29428);
or U32347 (N_32347,N_26149,N_28247);
nand U32348 (N_32348,N_28978,N_25267);
xnor U32349 (N_32349,N_29483,N_27426);
and U32350 (N_32350,N_26923,N_28867);
xnor U32351 (N_32351,N_26822,N_29821);
nand U32352 (N_32352,N_25788,N_28234);
and U32353 (N_32353,N_26073,N_26002);
xor U32354 (N_32354,N_26315,N_29675);
nor U32355 (N_32355,N_28005,N_28245);
nor U32356 (N_32356,N_26932,N_26889);
nand U32357 (N_32357,N_27138,N_26376);
nand U32358 (N_32358,N_29089,N_28646);
nor U32359 (N_32359,N_29450,N_27637);
nand U32360 (N_32360,N_28159,N_27954);
nand U32361 (N_32361,N_28075,N_25328);
nand U32362 (N_32362,N_25284,N_28037);
nor U32363 (N_32363,N_25371,N_29108);
xor U32364 (N_32364,N_26933,N_25197);
nand U32365 (N_32365,N_27246,N_26508);
nand U32366 (N_32366,N_27181,N_28106);
xor U32367 (N_32367,N_25093,N_25150);
and U32368 (N_32368,N_27261,N_29989);
nand U32369 (N_32369,N_26834,N_27210);
nor U32370 (N_32370,N_25327,N_29296);
and U32371 (N_32371,N_26133,N_28928);
nand U32372 (N_32372,N_26994,N_25668);
or U32373 (N_32373,N_25119,N_29652);
and U32374 (N_32374,N_28141,N_29465);
or U32375 (N_32375,N_29670,N_27987);
xor U32376 (N_32376,N_27948,N_25924);
and U32377 (N_32377,N_27675,N_29475);
or U32378 (N_32378,N_29898,N_25181);
or U32379 (N_32379,N_27294,N_25440);
xor U32380 (N_32380,N_29096,N_29679);
nand U32381 (N_32381,N_29488,N_28457);
xor U32382 (N_32382,N_25917,N_26795);
nand U32383 (N_32383,N_25658,N_26716);
nor U32384 (N_32384,N_29900,N_28395);
nand U32385 (N_32385,N_27915,N_28904);
or U32386 (N_32386,N_27858,N_27746);
xor U32387 (N_32387,N_25739,N_28761);
or U32388 (N_32388,N_28758,N_27537);
xor U32389 (N_32389,N_27263,N_27015);
and U32390 (N_32390,N_25634,N_27733);
nor U32391 (N_32391,N_29700,N_27913);
or U32392 (N_32392,N_28495,N_29734);
nor U32393 (N_32393,N_28525,N_28888);
nand U32394 (N_32394,N_28649,N_29987);
and U32395 (N_32395,N_26347,N_25545);
xnor U32396 (N_32396,N_25761,N_26473);
and U32397 (N_32397,N_27506,N_26978);
and U32398 (N_32398,N_25722,N_25547);
or U32399 (N_32399,N_29321,N_26796);
and U32400 (N_32400,N_25629,N_25897);
nor U32401 (N_32401,N_28951,N_29205);
nor U32402 (N_32402,N_26489,N_27123);
xnor U32403 (N_32403,N_25496,N_28365);
or U32404 (N_32404,N_25478,N_26511);
or U32405 (N_32405,N_25497,N_27645);
and U32406 (N_32406,N_26955,N_29300);
xor U32407 (N_32407,N_27292,N_29087);
xor U32408 (N_32408,N_29835,N_26423);
and U32409 (N_32409,N_29147,N_26029);
nor U32410 (N_32410,N_27635,N_29834);
xnor U32411 (N_32411,N_28700,N_26818);
nor U32412 (N_32412,N_29871,N_26304);
or U32413 (N_32413,N_29797,N_27269);
nor U32414 (N_32414,N_25332,N_25821);
and U32415 (N_32415,N_29727,N_27572);
xnor U32416 (N_32416,N_25443,N_27539);
or U32417 (N_32417,N_28813,N_26944);
and U32418 (N_32418,N_28435,N_29122);
nand U32419 (N_32419,N_29510,N_29532);
nand U32420 (N_32420,N_25240,N_27986);
nand U32421 (N_32421,N_27988,N_25596);
xnor U32422 (N_32422,N_25007,N_29464);
nor U32423 (N_32423,N_29244,N_27063);
nor U32424 (N_32424,N_26764,N_27752);
and U32425 (N_32425,N_26741,N_29629);
nor U32426 (N_32426,N_28500,N_25006);
nor U32427 (N_32427,N_28906,N_28953);
or U32428 (N_32428,N_26691,N_28879);
nand U32429 (N_32429,N_29180,N_28918);
nand U32430 (N_32430,N_29856,N_26616);
and U32431 (N_32431,N_29426,N_27451);
and U32432 (N_32432,N_25180,N_26386);
xnor U32433 (N_32433,N_26335,N_26733);
and U32434 (N_32434,N_25937,N_27965);
and U32435 (N_32435,N_25245,N_27164);
nand U32436 (N_32436,N_29681,N_28233);
xnor U32437 (N_32437,N_27887,N_27030);
nand U32438 (N_32438,N_28961,N_25319);
nand U32439 (N_32439,N_27283,N_29099);
nor U32440 (N_32440,N_28307,N_29502);
nor U32441 (N_32441,N_28192,N_25756);
xor U32442 (N_32442,N_26524,N_25118);
nand U32443 (N_32443,N_27843,N_29613);
and U32444 (N_32444,N_27628,N_25065);
xnor U32445 (N_32445,N_25365,N_26348);
or U32446 (N_32446,N_29394,N_25822);
and U32447 (N_32447,N_27659,N_28427);
and U32448 (N_32448,N_28386,N_26284);
nand U32449 (N_32449,N_25132,N_25680);
nor U32450 (N_32450,N_27984,N_27059);
nand U32451 (N_32451,N_25139,N_28205);
and U32452 (N_32452,N_27381,N_27052);
nand U32453 (N_32453,N_26271,N_28577);
nand U32454 (N_32454,N_28790,N_27111);
nor U32455 (N_32455,N_29070,N_29958);
and U32456 (N_32456,N_26666,N_26011);
xnor U32457 (N_32457,N_29954,N_29947);
or U32458 (N_32458,N_29939,N_26229);
xor U32459 (N_32459,N_26961,N_27826);
nor U32460 (N_32460,N_27300,N_26755);
or U32461 (N_32461,N_28744,N_29361);
and U32462 (N_32462,N_28456,N_26685);
nand U32463 (N_32463,N_28403,N_25238);
nor U32464 (N_32464,N_28420,N_26385);
and U32465 (N_32465,N_27975,N_28730);
xnor U32466 (N_32466,N_27765,N_29202);
xnor U32467 (N_32467,N_26595,N_29759);
nor U32468 (N_32468,N_29817,N_28221);
and U32469 (N_32469,N_25106,N_27044);
and U32470 (N_32470,N_25488,N_26199);
xnor U32471 (N_32471,N_25052,N_25747);
nand U32472 (N_32472,N_29412,N_27343);
or U32473 (N_32473,N_27751,N_28415);
nand U32474 (N_32474,N_27529,N_27310);
and U32475 (N_32475,N_27615,N_25615);
and U32476 (N_32476,N_26702,N_25946);
and U32477 (N_32477,N_27304,N_25178);
nand U32478 (N_32478,N_28499,N_27036);
xor U32479 (N_32479,N_26150,N_28226);
xor U32480 (N_32480,N_26059,N_28216);
xor U32481 (N_32481,N_26128,N_25243);
or U32482 (N_32482,N_27772,N_26077);
nor U32483 (N_32483,N_27025,N_29203);
nor U32484 (N_32484,N_28840,N_29458);
or U32485 (N_32485,N_26881,N_26584);
xnor U32486 (N_32486,N_26308,N_25160);
and U32487 (N_32487,N_29854,N_26863);
and U32488 (N_32488,N_28238,N_28707);
and U32489 (N_32489,N_25120,N_26085);
xor U32490 (N_32490,N_28213,N_26318);
xnor U32491 (N_32491,N_25895,N_29551);
or U32492 (N_32492,N_28656,N_28517);
and U32493 (N_32493,N_25459,N_26857);
nand U32494 (N_32494,N_25157,N_28948);
xnor U32495 (N_32495,N_25482,N_26434);
nor U32496 (N_32496,N_26092,N_28843);
xnor U32497 (N_32497,N_29041,N_26343);
nand U32498 (N_32498,N_27266,N_28729);
xnor U32499 (N_32499,N_25338,N_27571);
nand U32500 (N_32500,N_29344,N_29737);
or U32501 (N_32501,N_25356,N_25913);
nand U32502 (N_32502,N_29259,N_29670);
nand U32503 (N_32503,N_28984,N_26918);
and U32504 (N_32504,N_26177,N_27159);
nor U32505 (N_32505,N_26471,N_27656);
nand U32506 (N_32506,N_25650,N_25198);
xnor U32507 (N_32507,N_26525,N_28488);
nand U32508 (N_32508,N_25411,N_27619);
nor U32509 (N_32509,N_29232,N_28993);
nand U32510 (N_32510,N_25654,N_27332);
nor U32511 (N_32511,N_25633,N_26370);
and U32512 (N_32512,N_28748,N_29001);
or U32513 (N_32513,N_26887,N_25348);
or U32514 (N_32514,N_28823,N_28465);
and U32515 (N_32515,N_29873,N_26245);
and U32516 (N_32516,N_25814,N_29882);
nor U32517 (N_32517,N_27609,N_26588);
or U32518 (N_32518,N_25097,N_29047);
or U32519 (N_32519,N_28933,N_26175);
nor U32520 (N_32520,N_28111,N_28128);
xnor U32521 (N_32521,N_27309,N_26793);
and U32522 (N_32522,N_25112,N_29792);
nor U32523 (N_32523,N_29199,N_25873);
nand U32524 (N_32524,N_26925,N_28450);
and U32525 (N_32525,N_27810,N_28517);
or U32526 (N_32526,N_25425,N_27296);
and U32527 (N_32527,N_26516,N_25546);
or U32528 (N_32528,N_28567,N_29497);
nand U32529 (N_32529,N_29877,N_25386);
or U32530 (N_32530,N_29897,N_27636);
and U32531 (N_32531,N_28117,N_26892);
xnor U32532 (N_32532,N_29386,N_29743);
or U32533 (N_32533,N_27462,N_27214);
nand U32534 (N_32534,N_29169,N_29065);
nand U32535 (N_32535,N_29611,N_28216);
xor U32536 (N_32536,N_28829,N_27114);
nand U32537 (N_32537,N_27319,N_27882);
nor U32538 (N_32538,N_29206,N_29909);
and U32539 (N_32539,N_27465,N_28195);
nand U32540 (N_32540,N_26696,N_27448);
nand U32541 (N_32541,N_26150,N_25686);
nand U32542 (N_32542,N_26628,N_26525);
or U32543 (N_32543,N_26689,N_28900);
nand U32544 (N_32544,N_29110,N_26029);
or U32545 (N_32545,N_25084,N_28984);
nand U32546 (N_32546,N_28986,N_26473);
nor U32547 (N_32547,N_28978,N_27317);
or U32548 (N_32548,N_27613,N_27954);
and U32549 (N_32549,N_26143,N_29830);
or U32550 (N_32550,N_25531,N_25187);
xor U32551 (N_32551,N_27613,N_28561);
xor U32552 (N_32552,N_29600,N_27756);
nor U32553 (N_32553,N_28897,N_28775);
nand U32554 (N_32554,N_29118,N_27299);
xnor U32555 (N_32555,N_27142,N_29461);
and U32556 (N_32556,N_25943,N_26618);
nor U32557 (N_32557,N_28261,N_27528);
nor U32558 (N_32558,N_25293,N_25278);
or U32559 (N_32559,N_29851,N_25753);
and U32560 (N_32560,N_29163,N_27934);
and U32561 (N_32561,N_25299,N_29301);
nor U32562 (N_32562,N_29514,N_29342);
nand U32563 (N_32563,N_26397,N_25812);
nor U32564 (N_32564,N_28249,N_27956);
nor U32565 (N_32565,N_28145,N_27429);
xor U32566 (N_32566,N_25189,N_25644);
and U32567 (N_32567,N_28756,N_27457);
and U32568 (N_32568,N_27752,N_28986);
or U32569 (N_32569,N_26272,N_29776);
or U32570 (N_32570,N_26213,N_29418);
and U32571 (N_32571,N_25867,N_26172);
nand U32572 (N_32572,N_28082,N_26062);
nor U32573 (N_32573,N_25708,N_25915);
and U32574 (N_32574,N_26587,N_26766);
xnor U32575 (N_32575,N_29806,N_26355);
nand U32576 (N_32576,N_29033,N_29114);
xnor U32577 (N_32577,N_28589,N_28237);
nor U32578 (N_32578,N_25948,N_29435);
xnor U32579 (N_32579,N_28696,N_28153);
and U32580 (N_32580,N_29617,N_26863);
nand U32581 (N_32581,N_28097,N_29480);
xor U32582 (N_32582,N_26716,N_25097);
or U32583 (N_32583,N_27365,N_25431);
and U32584 (N_32584,N_26213,N_27210);
xnor U32585 (N_32585,N_26140,N_28615);
and U32586 (N_32586,N_29875,N_26727);
nor U32587 (N_32587,N_29041,N_25215);
nor U32588 (N_32588,N_29334,N_27517);
nand U32589 (N_32589,N_26610,N_28829);
nand U32590 (N_32590,N_26477,N_28468);
nor U32591 (N_32591,N_26222,N_29849);
nand U32592 (N_32592,N_28930,N_26730);
nand U32593 (N_32593,N_27237,N_29968);
and U32594 (N_32594,N_26729,N_29262);
nand U32595 (N_32595,N_26912,N_29279);
and U32596 (N_32596,N_28523,N_27338);
and U32597 (N_32597,N_27094,N_27660);
or U32598 (N_32598,N_26714,N_29237);
or U32599 (N_32599,N_28392,N_29822);
nand U32600 (N_32600,N_25375,N_25004);
nor U32601 (N_32601,N_26716,N_29033);
nand U32602 (N_32602,N_28197,N_28155);
xnor U32603 (N_32603,N_27899,N_25896);
or U32604 (N_32604,N_29218,N_29038);
xnor U32605 (N_32605,N_28814,N_29630);
or U32606 (N_32606,N_27072,N_28643);
and U32607 (N_32607,N_25496,N_27379);
or U32608 (N_32608,N_25470,N_27453);
nand U32609 (N_32609,N_29565,N_29744);
nor U32610 (N_32610,N_27980,N_29718);
xnor U32611 (N_32611,N_26181,N_28917);
nand U32612 (N_32612,N_26688,N_25743);
or U32613 (N_32613,N_29681,N_25665);
or U32614 (N_32614,N_28803,N_29406);
or U32615 (N_32615,N_26311,N_28000);
or U32616 (N_32616,N_27276,N_27148);
xnor U32617 (N_32617,N_27407,N_27899);
nand U32618 (N_32618,N_28798,N_27340);
and U32619 (N_32619,N_25213,N_28637);
nor U32620 (N_32620,N_26130,N_25098);
nand U32621 (N_32621,N_26358,N_26916);
and U32622 (N_32622,N_28541,N_28106);
and U32623 (N_32623,N_29339,N_29103);
nor U32624 (N_32624,N_26588,N_26156);
and U32625 (N_32625,N_26991,N_28876);
and U32626 (N_32626,N_29590,N_27887);
and U32627 (N_32627,N_26326,N_25466);
and U32628 (N_32628,N_26639,N_29055);
nor U32629 (N_32629,N_29205,N_26474);
and U32630 (N_32630,N_26617,N_26642);
nand U32631 (N_32631,N_27662,N_27219);
nor U32632 (N_32632,N_25070,N_27570);
nand U32633 (N_32633,N_28767,N_25923);
nand U32634 (N_32634,N_27432,N_29040);
xor U32635 (N_32635,N_25980,N_26945);
and U32636 (N_32636,N_28946,N_28997);
or U32637 (N_32637,N_27369,N_29470);
and U32638 (N_32638,N_27715,N_28099);
or U32639 (N_32639,N_25038,N_26236);
xor U32640 (N_32640,N_27297,N_25399);
nor U32641 (N_32641,N_29424,N_25087);
nand U32642 (N_32642,N_27501,N_26952);
and U32643 (N_32643,N_27708,N_26277);
nand U32644 (N_32644,N_26080,N_28544);
and U32645 (N_32645,N_25335,N_25052);
nor U32646 (N_32646,N_29645,N_29397);
and U32647 (N_32647,N_26419,N_27840);
nor U32648 (N_32648,N_29768,N_25457);
or U32649 (N_32649,N_29362,N_27501);
xnor U32650 (N_32650,N_27721,N_27141);
or U32651 (N_32651,N_27851,N_28648);
nand U32652 (N_32652,N_26458,N_27695);
nand U32653 (N_32653,N_27008,N_29692);
xnor U32654 (N_32654,N_29133,N_28998);
or U32655 (N_32655,N_25531,N_29687);
nor U32656 (N_32656,N_26424,N_27833);
nor U32657 (N_32657,N_27216,N_25994);
or U32658 (N_32658,N_26967,N_28413);
xnor U32659 (N_32659,N_25115,N_26190);
and U32660 (N_32660,N_26038,N_27957);
and U32661 (N_32661,N_27387,N_29785);
nand U32662 (N_32662,N_29756,N_27780);
nor U32663 (N_32663,N_25996,N_27694);
xnor U32664 (N_32664,N_26982,N_29748);
xnor U32665 (N_32665,N_27264,N_27454);
and U32666 (N_32666,N_29641,N_28847);
nand U32667 (N_32667,N_27696,N_26073);
or U32668 (N_32668,N_27180,N_25596);
and U32669 (N_32669,N_29569,N_28500);
nor U32670 (N_32670,N_29963,N_28236);
nor U32671 (N_32671,N_29731,N_25513);
nand U32672 (N_32672,N_29061,N_25100);
xor U32673 (N_32673,N_29340,N_25628);
nand U32674 (N_32674,N_28115,N_26528);
xnor U32675 (N_32675,N_29082,N_27013);
nor U32676 (N_32676,N_29846,N_26897);
xnor U32677 (N_32677,N_27001,N_29069);
nand U32678 (N_32678,N_25074,N_29169);
or U32679 (N_32679,N_27158,N_27316);
nand U32680 (N_32680,N_26736,N_28424);
or U32681 (N_32681,N_28767,N_29601);
and U32682 (N_32682,N_26977,N_28025);
xor U32683 (N_32683,N_27674,N_29564);
or U32684 (N_32684,N_26534,N_29322);
nor U32685 (N_32685,N_28639,N_29684);
xnor U32686 (N_32686,N_28426,N_27747);
and U32687 (N_32687,N_29713,N_26849);
and U32688 (N_32688,N_26458,N_26001);
nor U32689 (N_32689,N_27727,N_29560);
or U32690 (N_32690,N_27261,N_29854);
nor U32691 (N_32691,N_25035,N_25365);
or U32692 (N_32692,N_25529,N_26727);
xnor U32693 (N_32693,N_26110,N_28525);
and U32694 (N_32694,N_25735,N_25589);
xnor U32695 (N_32695,N_26525,N_26855);
and U32696 (N_32696,N_26866,N_27252);
xnor U32697 (N_32697,N_25315,N_28029);
and U32698 (N_32698,N_29604,N_27041);
nand U32699 (N_32699,N_28832,N_26994);
or U32700 (N_32700,N_26996,N_25210);
and U32701 (N_32701,N_28804,N_28792);
nor U32702 (N_32702,N_29018,N_29706);
nand U32703 (N_32703,N_26731,N_27148);
or U32704 (N_32704,N_28742,N_25836);
or U32705 (N_32705,N_26009,N_29934);
nand U32706 (N_32706,N_29312,N_25765);
xor U32707 (N_32707,N_28065,N_29512);
xor U32708 (N_32708,N_26661,N_29755);
nor U32709 (N_32709,N_25659,N_27217);
or U32710 (N_32710,N_25664,N_28736);
and U32711 (N_32711,N_27264,N_26827);
xor U32712 (N_32712,N_25391,N_25371);
and U32713 (N_32713,N_29508,N_28777);
nor U32714 (N_32714,N_28182,N_28581);
and U32715 (N_32715,N_25547,N_26080);
and U32716 (N_32716,N_25195,N_25972);
nor U32717 (N_32717,N_29503,N_27950);
xnor U32718 (N_32718,N_29342,N_28658);
and U32719 (N_32719,N_25484,N_28206);
or U32720 (N_32720,N_27172,N_27838);
xor U32721 (N_32721,N_29031,N_29090);
nor U32722 (N_32722,N_28068,N_29358);
or U32723 (N_32723,N_28154,N_29808);
nor U32724 (N_32724,N_26036,N_25389);
nor U32725 (N_32725,N_28864,N_28998);
nand U32726 (N_32726,N_29662,N_27132);
and U32727 (N_32727,N_28533,N_27186);
or U32728 (N_32728,N_26498,N_29636);
or U32729 (N_32729,N_27067,N_25797);
and U32730 (N_32730,N_28193,N_27855);
nand U32731 (N_32731,N_28323,N_25172);
and U32732 (N_32732,N_29954,N_27860);
and U32733 (N_32733,N_28064,N_29013);
xor U32734 (N_32734,N_25894,N_28610);
nor U32735 (N_32735,N_27547,N_27103);
or U32736 (N_32736,N_26079,N_25106);
or U32737 (N_32737,N_26033,N_26817);
nand U32738 (N_32738,N_26651,N_28017);
or U32739 (N_32739,N_27724,N_26844);
and U32740 (N_32740,N_27967,N_28385);
nor U32741 (N_32741,N_27877,N_26249);
nor U32742 (N_32742,N_25255,N_27960);
nor U32743 (N_32743,N_27963,N_29493);
nand U32744 (N_32744,N_25132,N_25732);
nor U32745 (N_32745,N_28842,N_27802);
nand U32746 (N_32746,N_27043,N_25797);
nand U32747 (N_32747,N_28115,N_27634);
xor U32748 (N_32748,N_27263,N_27276);
or U32749 (N_32749,N_26184,N_28240);
xor U32750 (N_32750,N_27036,N_25603);
nor U32751 (N_32751,N_28845,N_26916);
nor U32752 (N_32752,N_25827,N_28179);
xor U32753 (N_32753,N_26669,N_29486);
nor U32754 (N_32754,N_25357,N_27019);
nor U32755 (N_32755,N_26957,N_26684);
nor U32756 (N_32756,N_29308,N_27326);
nand U32757 (N_32757,N_28595,N_26878);
or U32758 (N_32758,N_27534,N_27055);
or U32759 (N_32759,N_29508,N_27941);
or U32760 (N_32760,N_26959,N_28026);
or U32761 (N_32761,N_28106,N_27726);
nand U32762 (N_32762,N_27904,N_27675);
nor U32763 (N_32763,N_26177,N_27317);
xor U32764 (N_32764,N_27381,N_29655);
and U32765 (N_32765,N_29448,N_27559);
nand U32766 (N_32766,N_29258,N_25133);
xnor U32767 (N_32767,N_29103,N_29815);
nand U32768 (N_32768,N_28671,N_29086);
and U32769 (N_32769,N_26567,N_28988);
or U32770 (N_32770,N_28784,N_28175);
nor U32771 (N_32771,N_29466,N_27465);
xnor U32772 (N_32772,N_25102,N_27043);
nor U32773 (N_32773,N_28751,N_29263);
nand U32774 (N_32774,N_28800,N_28476);
xor U32775 (N_32775,N_29878,N_28548);
and U32776 (N_32776,N_26367,N_27648);
and U32777 (N_32777,N_26806,N_26488);
xnor U32778 (N_32778,N_27171,N_25931);
nand U32779 (N_32779,N_29956,N_27608);
and U32780 (N_32780,N_25827,N_26433);
or U32781 (N_32781,N_27221,N_29988);
and U32782 (N_32782,N_28104,N_25077);
or U32783 (N_32783,N_28470,N_28453);
nor U32784 (N_32784,N_29053,N_29475);
and U32785 (N_32785,N_28128,N_27930);
nand U32786 (N_32786,N_29067,N_28248);
nand U32787 (N_32787,N_29606,N_25717);
and U32788 (N_32788,N_27938,N_29710);
or U32789 (N_32789,N_26121,N_27068);
xor U32790 (N_32790,N_25143,N_29014);
xor U32791 (N_32791,N_29845,N_28016);
xnor U32792 (N_32792,N_28321,N_29892);
nand U32793 (N_32793,N_29182,N_29964);
nor U32794 (N_32794,N_26020,N_25842);
xnor U32795 (N_32795,N_26542,N_26148);
nand U32796 (N_32796,N_26737,N_27294);
xnor U32797 (N_32797,N_28318,N_29535);
or U32798 (N_32798,N_28971,N_28547);
and U32799 (N_32799,N_27033,N_25734);
or U32800 (N_32800,N_27304,N_28141);
or U32801 (N_32801,N_29024,N_27253);
xnor U32802 (N_32802,N_25792,N_29981);
and U32803 (N_32803,N_25367,N_28851);
and U32804 (N_32804,N_26350,N_28426);
and U32805 (N_32805,N_26685,N_29100);
nand U32806 (N_32806,N_29999,N_29049);
nand U32807 (N_32807,N_26104,N_25054);
or U32808 (N_32808,N_28899,N_28448);
and U32809 (N_32809,N_26602,N_29206);
or U32810 (N_32810,N_29086,N_28905);
nand U32811 (N_32811,N_26298,N_26407);
nand U32812 (N_32812,N_29220,N_25523);
nand U32813 (N_32813,N_25264,N_25185);
nor U32814 (N_32814,N_27199,N_27579);
xor U32815 (N_32815,N_28033,N_28813);
xor U32816 (N_32816,N_25664,N_29249);
nor U32817 (N_32817,N_26431,N_25448);
nand U32818 (N_32818,N_28920,N_25002);
or U32819 (N_32819,N_29859,N_26024);
or U32820 (N_32820,N_27927,N_29593);
nand U32821 (N_32821,N_28813,N_25664);
nand U32822 (N_32822,N_29516,N_25269);
nand U32823 (N_32823,N_29824,N_29168);
xnor U32824 (N_32824,N_29265,N_27476);
nand U32825 (N_32825,N_27348,N_28898);
nand U32826 (N_32826,N_26674,N_26931);
and U32827 (N_32827,N_26686,N_26774);
or U32828 (N_32828,N_28832,N_25606);
nand U32829 (N_32829,N_27638,N_26053);
and U32830 (N_32830,N_26549,N_26650);
xor U32831 (N_32831,N_25258,N_25737);
and U32832 (N_32832,N_27049,N_29590);
xnor U32833 (N_32833,N_25167,N_29269);
nand U32834 (N_32834,N_27265,N_28864);
xor U32835 (N_32835,N_29311,N_26546);
nand U32836 (N_32836,N_28070,N_29339);
nand U32837 (N_32837,N_25619,N_27422);
nand U32838 (N_32838,N_27952,N_29326);
xnor U32839 (N_32839,N_29266,N_27528);
or U32840 (N_32840,N_25962,N_29876);
and U32841 (N_32841,N_26801,N_27730);
or U32842 (N_32842,N_28342,N_26985);
or U32843 (N_32843,N_26014,N_27776);
or U32844 (N_32844,N_27947,N_29970);
nand U32845 (N_32845,N_26563,N_25243);
or U32846 (N_32846,N_27117,N_26485);
or U32847 (N_32847,N_26957,N_27443);
nor U32848 (N_32848,N_27260,N_26547);
xnor U32849 (N_32849,N_28816,N_25878);
nor U32850 (N_32850,N_26085,N_27749);
xor U32851 (N_32851,N_29485,N_25494);
and U32852 (N_32852,N_26319,N_25828);
nand U32853 (N_32853,N_27139,N_29995);
nor U32854 (N_32854,N_28385,N_25341);
xor U32855 (N_32855,N_25422,N_26970);
nor U32856 (N_32856,N_29249,N_26511);
or U32857 (N_32857,N_25185,N_25337);
xor U32858 (N_32858,N_26319,N_27587);
and U32859 (N_32859,N_27872,N_29098);
xnor U32860 (N_32860,N_25809,N_29963);
or U32861 (N_32861,N_28810,N_29480);
xor U32862 (N_32862,N_27825,N_27916);
xor U32863 (N_32863,N_26923,N_26604);
or U32864 (N_32864,N_25801,N_26193);
or U32865 (N_32865,N_28848,N_26251);
nor U32866 (N_32866,N_25521,N_27113);
nor U32867 (N_32867,N_25376,N_29457);
or U32868 (N_32868,N_25785,N_26866);
and U32869 (N_32869,N_26489,N_29023);
and U32870 (N_32870,N_29558,N_25306);
and U32871 (N_32871,N_27386,N_26568);
nand U32872 (N_32872,N_25583,N_29289);
xor U32873 (N_32873,N_28775,N_28137);
and U32874 (N_32874,N_28915,N_29705);
nand U32875 (N_32875,N_29130,N_28176);
nand U32876 (N_32876,N_28967,N_26072);
xnor U32877 (N_32877,N_27373,N_28265);
and U32878 (N_32878,N_29352,N_27293);
nand U32879 (N_32879,N_27154,N_29992);
and U32880 (N_32880,N_29641,N_25828);
or U32881 (N_32881,N_27588,N_29993);
nor U32882 (N_32882,N_27930,N_26867);
xnor U32883 (N_32883,N_28856,N_27421);
nand U32884 (N_32884,N_28459,N_29634);
xnor U32885 (N_32885,N_29116,N_26412);
and U32886 (N_32886,N_25077,N_28784);
nand U32887 (N_32887,N_27813,N_25291);
or U32888 (N_32888,N_26298,N_27390);
nor U32889 (N_32889,N_26426,N_25714);
and U32890 (N_32890,N_27736,N_27956);
or U32891 (N_32891,N_25651,N_25500);
nor U32892 (N_32892,N_26308,N_27904);
or U32893 (N_32893,N_29809,N_29530);
nand U32894 (N_32894,N_29895,N_29059);
or U32895 (N_32895,N_25801,N_25969);
or U32896 (N_32896,N_25945,N_27103);
xor U32897 (N_32897,N_28559,N_29552);
or U32898 (N_32898,N_25378,N_25874);
and U32899 (N_32899,N_26486,N_29822);
nand U32900 (N_32900,N_28136,N_27687);
xor U32901 (N_32901,N_26076,N_27924);
or U32902 (N_32902,N_29435,N_26488);
and U32903 (N_32903,N_27627,N_25564);
or U32904 (N_32904,N_25736,N_26889);
nand U32905 (N_32905,N_26423,N_29308);
nand U32906 (N_32906,N_28897,N_29179);
or U32907 (N_32907,N_25908,N_29345);
nor U32908 (N_32908,N_26207,N_26901);
nor U32909 (N_32909,N_28059,N_27354);
and U32910 (N_32910,N_27681,N_29933);
and U32911 (N_32911,N_27150,N_27792);
nor U32912 (N_32912,N_26242,N_29665);
xnor U32913 (N_32913,N_28386,N_29580);
nor U32914 (N_32914,N_29244,N_25995);
nand U32915 (N_32915,N_29843,N_28889);
nand U32916 (N_32916,N_27901,N_27094);
or U32917 (N_32917,N_25354,N_26073);
and U32918 (N_32918,N_27140,N_26399);
nand U32919 (N_32919,N_25627,N_25162);
nand U32920 (N_32920,N_26911,N_28393);
or U32921 (N_32921,N_25012,N_27745);
or U32922 (N_32922,N_27637,N_25055);
xor U32923 (N_32923,N_27886,N_26210);
and U32924 (N_32924,N_28584,N_28888);
xnor U32925 (N_32925,N_25664,N_28341);
nor U32926 (N_32926,N_27649,N_27410);
or U32927 (N_32927,N_26213,N_25977);
nor U32928 (N_32928,N_25857,N_29446);
or U32929 (N_32929,N_26565,N_25265);
and U32930 (N_32930,N_29780,N_27008);
nand U32931 (N_32931,N_25039,N_26490);
or U32932 (N_32932,N_25841,N_26103);
xor U32933 (N_32933,N_27430,N_25623);
xor U32934 (N_32934,N_26828,N_25080);
nor U32935 (N_32935,N_28925,N_28884);
and U32936 (N_32936,N_26946,N_28788);
nand U32937 (N_32937,N_25655,N_29471);
xnor U32938 (N_32938,N_27309,N_28242);
nor U32939 (N_32939,N_26123,N_27338);
nand U32940 (N_32940,N_28111,N_26841);
xor U32941 (N_32941,N_27711,N_29917);
nor U32942 (N_32942,N_26502,N_27873);
or U32943 (N_32943,N_27057,N_25623);
nor U32944 (N_32944,N_29254,N_29150);
nand U32945 (N_32945,N_29523,N_27848);
xor U32946 (N_32946,N_25995,N_29074);
and U32947 (N_32947,N_28832,N_28678);
or U32948 (N_32948,N_26070,N_25221);
nand U32949 (N_32949,N_29460,N_27036);
and U32950 (N_32950,N_27209,N_29758);
and U32951 (N_32951,N_25219,N_25244);
xor U32952 (N_32952,N_29750,N_26644);
and U32953 (N_32953,N_25169,N_25154);
nand U32954 (N_32954,N_25010,N_26665);
and U32955 (N_32955,N_26448,N_27021);
xor U32956 (N_32956,N_25387,N_26659);
and U32957 (N_32957,N_27764,N_27263);
or U32958 (N_32958,N_27090,N_25725);
or U32959 (N_32959,N_26367,N_29628);
and U32960 (N_32960,N_27287,N_27352);
xnor U32961 (N_32961,N_25142,N_28895);
and U32962 (N_32962,N_27302,N_26120);
xor U32963 (N_32963,N_29334,N_28251);
or U32964 (N_32964,N_29655,N_27789);
and U32965 (N_32965,N_25813,N_29636);
xnor U32966 (N_32966,N_26406,N_28483);
xor U32967 (N_32967,N_28265,N_25836);
or U32968 (N_32968,N_29782,N_29491);
and U32969 (N_32969,N_28999,N_25128);
and U32970 (N_32970,N_29731,N_29510);
or U32971 (N_32971,N_26325,N_25214);
or U32972 (N_32972,N_25001,N_25245);
nand U32973 (N_32973,N_27249,N_26644);
xor U32974 (N_32974,N_27312,N_26234);
xnor U32975 (N_32975,N_29375,N_28229);
and U32976 (N_32976,N_28464,N_29263);
and U32977 (N_32977,N_25705,N_28968);
xor U32978 (N_32978,N_25322,N_25571);
or U32979 (N_32979,N_28346,N_28141);
nor U32980 (N_32980,N_25102,N_29590);
and U32981 (N_32981,N_26822,N_25714);
and U32982 (N_32982,N_25653,N_25922);
or U32983 (N_32983,N_28579,N_29505);
and U32984 (N_32984,N_26991,N_29860);
nor U32985 (N_32985,N_27741,N_27499);
or U32986 (N_32986,N_29900,N_28268);
xor U32987 (N_32987,N_25857,N_28209);
nand U32988 (N_32988,N_28668,N_29859);
xor U32989 (N_32989,N_29153,N_27107);
and U32990 (N_32990,N_29086,N_25432);
xnor U32991 (N_32991,N_27142,N_28629);
nor U32992 (N_32992,N_28051,N_25946);
or U32993 (N_32993,N_25817,N_28823);
or U32994 (N_32994,N_26657,N_26382);
nand U32995 (N_32995,N_29077,N_25203);
or U32996 (N_32996,N_29080,N_28940);
nor U32997 (N_32997,N_25656,N_25557);
and U32998 (N_32998,N_29152,N_28985);
and U32999 (N_32999,N_29891,N_27395);
and U33000 (N_33000,N_27582,N_26179);
nand U33001 (N_33001,N_29715,N_26037);
nand U33002 (N_33002,N_27839,N_28117);
or U33003 (N_33003,N_28438,N_27322);
and U33004 (N_33004,N_26066,N_29549);
nor U33005 (N_33005,N_29524,N_27708);
nand U33006 (N_33006,N_26534,N_25884);
or U33007 (N_33007,N_26431,N_26768);
nor U33008 (N_33008,N_26143,N_28738);
nand U33009 (N_33009,N_28246,N_25457);
nor U33010 (N_33010,N_26348,N_26689);
nand U33011 (N_33011,N_27655,N_28042);
and U33012 (N_33012,N_25941,N_27375);
and U33013 (N_33013,N_29950,N_26882);
nand U33014 (N_33014,N_28864,N_27361);
or U33015 (N_33015,N_25667,N_26076);
or U33016 (N_33016,N_29585,N_27178);
nand U33017 (N_33017,N_25730,N_25453);
xnor U33018 (N_33018,N_25278,N_28264);
or U33019 (N_33019,N_27076,N_29650);
nand U33020 (N_33020,N_27452,N_28836);
and U33021 (N_33021,N_29232,N_26723);
nand U33022 (N_33022,N_25463,N_26493);
nor U33023 (N_33023,N_29093,N_28268);
or U33024 (N_33024,N_28147,N_28061);
xnor U33025 (N_33025,N_27172,N_25401);
xor U33026 (N_33026,N_29908,N_26374);
nor U33027 (N_33027,N_27484,N_27322);
or U33028 (N_33028,N_26035,N_28252);
xnor U33029 (N_33029,N_28661,N_27970);
nor U33030 (N_33030,N_28897,N_25903);
and U33031 (N_33031,N_27581,N_29828);
nor U33032 (N_33032,N_25127,N_29104);
nor U33033 (N_33033,N_29122,N_27570);
nand U33034 (N_33034,N_28215,N_28948);
nor U33035 (N_33035,N_26308,N_29266);
nand U33036 (N_33036,N_29115,N_28279);
or U33037 (N_33037,N_29080,N_26775);
nor U33038 (N_33038,N_28752,N_27303);
and U33039 (N_33039,N_25321,N_29969);
nand U33040 (N_33040,N_27789,N_26570);
nand U33041 (N_33041,N_26612,N_25941);
or U33042 (N_33042,N_29715,N_28439);
or U33043 (N_33043,N_28674,N_25794);
and U33044 (N_33044,N_28698,N_26577);
or U33045 (N_33045,N_27582,N_28381);
and U33046 (N_33046,N_27265,N_26065);
or U33047 (N_33047,N_27574,N_27258);
nor U33048 (N_33048,N_25720,N_27845);
or U33049 (N_33049,N_28341,N_28154);
nand U33050 (N_33050,N_26044,N_26814);
nor U33051 (N_33051,N_28029,N_28470);
or U33052 (N_33052,N_28059,N_29978);
and U33053 (N_33053,N_26929,N_29935);
nand U33054 (N_33054,N_27343,N_26675);
nand U33055 (N_33055,N_29340,N_28543);
or U33056 (N_33056,N_29938,N_28065);
or U33057 (N_33057,N_26828,N_28642);
nor U33058 (N_33058,N_25387,N_28857);
and U33059 (N_33059,N_29176,N_27180);
nand U33060 (N_33060,N_27474,N_29322);
and U33061 (N_33061,N_25436,N_27002);
xnor U33062 (N_33062,N_26146,N_26447);
nand U33063 (N_33063,N_28485,N_26987);
or U33064 (N_33064,N_29764,N_28419);
nor U33065 (N_33065,N_25528,N_27516);
and U33066 (N_33066,N_28554,N_25647);
or U33067 (N_33067,N_29699,N_25910);
or U33068 (N_33068,N_25786,N_26163);
nand U33069 (N_33069,N_26220,N_25099);
nor U33070 (N_33070,N_27578,N_26358);
or U33071 (N_33071,N_28866,N_29001);
nand U33072 (N_33072,N_27237,N_28843);
and U33073 (N_33073,N_25575,N_28138);
or U33074 (N_33074,N_29336,N_27790);
nand U33075 (N_33075,N_29938,N_28255);
or U33076 (N_33076,N_29771,N_29206);
nor U33077 (N_33077,N_25756,N_28464);
nor U33078 (N_33078,N_28359,N_27626);
or U33079 (N_33079,N_27339,N_28864);
xnor U33080 (N_33080,N_25528,N_28014);
and U33081 (N_33081,N_27418,N_28842);
nor U33082 (N_33082,N_25570,N_28235);
xnor U33083 (N_33083,N_27942,N_29926);
nor U33084 (N_33084,N_26553,N_25031);
nor U33085 (N_33085,N_26222,N_29556);
nor U33086 (N_33086,N_26186,N_29553);
and U33087 (N_33087,N_28851,N_26471);
nand U33088 (N_33088,N_28274,N_27465);
and U33089 (N_33089,N_28906,N_28771);
xnor U33090 (N_33090,N_28497,N_28462);
xnor U33091 (N_33091,N_29097,N_29554);
nand U33092 (N_33092,N_27559,N_28631);
and U33093 (N_33093,N_28157,N_27505);
xor U33094 (N_33094,N_25633,N_28258);
or U33095 (N_33095,N_29962,N_29532);
nand U33096 (N_33096,N_27252,N_27938);
nor U33097 (N_33097,N_26019,N_28010);
xnor U33098 (N_33098,N_27674,N_29955);
nor U33099 (N_33099,N_28810,N_27735);
or U33100 (N_33100,N_25865,N_25802);
nor U33101 (N_33101,N_28295,N_29585);
or U33102 (N_33102,N_27396,N_26216);
nand U33103 (N_33103,N_25134,N_29295);
xor U33104 (N_33104,N_25999,N_29588);
or U33105 (N_33105,N_27216,N_26239);
nand U33106 (N_33106,N_26488,N_28698);
xor U33107 (N_33107,N_25445,N_28091);
and U33108 (N_33108,N_26066,N_25493);
nand U33109 (N_33109,N_26443,N_28067);
and U33110 (N_33110,N_26349,N_28351);
xnor U33111 (N_33111,N_28673,N_28112);
nor U33112 (N_33112,N_29150,N_28705);
and U33113 (N_33113,N_27394,N_26766);
nand U33114 (N_33114,N_28521,N_26171);
xor U33115 (N_33115,N_27974,N_25239);
nand U33116 (N_33116,N_25157,N_28270);
and U33117 (N_33117,N_27054,N_29704);
nor U33118 (N_33118,N_29712,N_25501);
nand U33119 (N_33119,N_28410,N_25973);
nor U33120 (N_33120,N_27149,N_25663);
nor U33121 (N_33121,N_28054,N_25290);
nand U33122 (N_33122,N_29064,N_29609);
nand U33123 (N_33123,N_27066,N_25836);
nor U33124 (N_33124,N_28124,N_25353);
or U33125 (N_33125,N_25047,N_25958);
or U33126 (N_33126,N_29633,N_27123);
nand U33127 (N_33127,N_27725,N_26462);
and U33128 (N_33128,N_29149,N_25241);
and U33129 (N_33129,N_27394,N_26910);
nand U33130 (N_33130,N_28185,N_26002);
and U33131 (N_33131,N_25129,N_25427);
or U33132 (N_33132,N_26867,N_26216);
nand U33133 (N_33133,N_25613,N_25026);
or U33134 (N_33134,N_27494,N_26581);
xnor U33135 (N_33135,N_29868,N_26540);
nor U33136 (N_33136,N_25201,N_25113);
nor U33137 (N_33137,N_28238,N_26203);
or U33138 (N_33138,N_29219,N_28474);
nand U33139 (N_33139,N_27206,N_27626);
xnor U33140 (N_33140,N_26934,N_28768);
xnor U33141 (N_33141,N_26790,N_26384);
nor U33142 (N_33142,N_26668,N_25645);
xor U33143 (N_33143,N_28379,N_26943);
xnor U33144 (N_33144,N_28667,N_26941);
nor U33145 (N_33145,N_26726,N_28199);
nor U33146 (N_33146,N_26222,N_28765);
or U33147 (N_33147,N_27216,N_25221);
xor U33148 (N_33148,N_25765,N_25111);
and U33149 (N_33149,N_28634,N_29513);
or U33150 (N_33150,N_28731,N_29969);
or U33151 (N_33151,N_28212,N_27436);
and U33152 (N_33152,N_26279,N_26870);
nand U33153 (N_33153,N_26082,N_26312);
or U33154 (N_33154,N_29399,N_29152);
xor U33155 (N_33155,N_25843,N_27310);
nand U33156 (N_33156,N_27729,N_28149);
nor U33157 (N_33157,N_25377,N_27494);
or U33158 (N_33158,N_28436,N_28431);
or U33159 (N_33159,N_26789,N_29575);
nand U33160 (N_33160,N_25846,N_29850);
and U33161 (N_33161,N_26135,N_26947);
nor U33162 (N_33162,N_25112,N_25178);
or U33163 (N_33163,N_28102,N_25101);
xnor U33164 (N_33164,N_29889,N_29361);
nor U33165 (N_33165,N_25890,N_25228);
nor U33166 (N_33166,N_25138,N_29862);
nor U33167 (N_33167,N_26125,N_27308);
or U33168 (N_33168,N_25790,N_29945);
and U33169 (N_33169,N_29481,N_27694);
and U33170 (N_33170,N_25607,N_27886);
and U33171 (N_33171,N_28779,N_26074);
and U33172 (N_33172,N_26609,N_26539);
xor U33173 (N_33173,N_27890,N_26377);
xor U33174 (N_33174,N_27600,N_26582);
or U33175 (N_33175,N_25052,N_26337);
nor U33176 (N_33176,N_26809,N_27678);
xnor U33177 (N_33177,N_29864,N_25053);
nor U33178 (N_33178,N_28273,N_26217);
nor U33179 (N_33179,N_25881,N_27965);
xnor U33180 (N_33180,N_28562,N_26663);
and U33181 (N_33181,N_26220,N_28095);
or U33182 (N_33182,N_25278,N_28257);
and U33183 (N_33183,N_29942,N_29462);
or U33184 (N_33184,N_28252,N_26388);
and U33185 (N_33185,N_27417,N_29710);
nor U33186 (N_33186,N_26153,N_27447);
or U33187 (N_33187,N_29487,N_26979);
nand U33188 (N_33188,N_26314,N_25559);
xor U33189 (N_33189,N_29694,N_25806);
nand U33190 (N_33190,N_25665,N_29686);
or U33191 (N_33191,N_28923,N_26762);
and U33192 (N_33192,N_29748,N_26702);
nor U33193 (N_33193,N_28106,N_29664);
or U33194 (N_33194,N_28722,N_25779);
and U33195 (N_33195,N_26559,N_25870);
and U33196 (N_33196,N_25156,N_25447);
and U33197 (N_33197,N_26709,N_28800);
nor U33198 (N_33198,N_28115,N_29460);
or U33199 (N_33199,N_27156,N_27128);
and U33200 (N_33200,N_26722,N_29736);
and U33201 (N_33201,N_29572,N_27460);
or U33202 (N_33202,N_26840,N_27871);
nor U33203 (N_33203,N_25174,N_28819);
nor U33204 (N_33204,N_27901,N_26087);
or U33205 (N_33205,N_25657,N_25557);
and U33206 (N_33206,N_27493,N_26826);
xnor U33207 (N_33207,N_27225,N_27307);
xnor U33208 (N_33208,N_25912,N_28568);
nor U33209 (N_33209,N_26786,N_28704);
and U33210 (N_33210,N_26628,N_25510);
nor U33211 (N_33211,N_29214,N_27968);
and U33212 (N_33212,N_28636,N_29770);
nand U33213 (N_33213,N_29459,N_28941);
or U33214 (N_33214,N_28410,N_27276);
xnor U33215 (N_33215,N_27030,N_29890);
nand U33216 (N_33216,N_26274,N_27275);
or U33217 (N_33217,N_28308,N_25465);
or U33218 (N_33218,N_27352,N_25480);
nor U33219 (N_33219,N_25137,N_26979);
nor U33220 (N_33220,N_28999,N_25794);
and U33221 (N_33221,N_26147,N_29088);
or U33222 (N_33222,N_28164,N_27927);
nand U33223 (N_33223,N_27671,N_26537);
nor U33224 (N_33224,N_28975,N_28139);
nor U33225 (N_33225,N_29851,N_26657);
and U33226 (N_33226,N_25593,N_29548);
nor U33227 (N_33227,N_26549,N_26985);
xnor U33228 (N_33228,N_29406,N_28539);
nand U33229 (N_33229,N_29752,N_27497);
nor U33230 (N_33230,N_28291,N_27650);
xor U33231 (N_33231,N_26668,N_25697);
or U33232 (N_33232,N_27239,N_25441);
nor U33233 (N_33233,N_28064,N_26900);
nor U33234 (N_33234,N_27218,N_25293);
nand U33235 (N_33235,N_26490,N_28002);
and U33236 (N_33236,N_28258,N_29291);
or U33237 (N_33237,N_27483,N_26729);
or U33238 (N_33238,N_25069,N_29274);
xnor U33239 (N_33239,N_29031,N_25060);
nor U33240 (N_33240,N_25734,N_25545);
xor U33241 (N_33241,N_27106,N_26515);
and U33242 (N_33242,N_26788,N_29354);
or U33243 (N_33243,N_27545,N_28707);
xor U33244 (N_33244,N_27150,N_26344);
nor U33245 (N_33245,N_28945,N_27464);
or U33246 (N_33246,N_26019,N_27323);
or U33247 (N_33247,N_25855,N_29678);
xnor U33248 (N_33248,N_26189,N_26230);
and U33249 (N_33249,N_25702,N_26769);
xor U33250 (N_33250,N_28844,N_28954);
nor U33251 (N_33251,N_26054,N_25232);
and U33252 (N_33252,N_27876,N_28030);
and U33253 (N_33253,N_27445,N_28579);
or U33254 (N_33254,N_25988,N_26951);
nand U33255 (N_33255,N_29965,N_27360);
and U33256 (N_33256,N_29863,N_25723);
nor U33257 (N_33257,N_26555,N_25199);
xor U33258 (N_33258,N_29233,N_28321);
and U33259 (N_33259,N_27559,N_29782);
nor U33260 (N_33260,N_26638,N_27190);
nand U33261 (N_33261,N_26298,N_29320);
and U33262 (N_33262,N_29692,N_28574);
and U33263 (N_33263,N_29253,N_28405);
xnor U33264 (N_33264,N_26500,N_26387);
nand U33265 (N_33265,N_27270,N_29136);
or U33266 (N_33266,N_28001,N_29094);
nor U33267 (N_33267,N_28436,N_27432);
nor U33268 (N_33268,N_26683,N_27784);
nand U33269 (N_33269,N_29361,N_25655);
nand U33270 (N_33270,N_27274,N_25976);
nor U33271 (N_33271,N_25373,N_27778);
nand U33272 (N_33272,N_27899,N_29790);
nor U33273 (N_33273,N_26481,N_26118);
xor U33274 (N_33274,N_27196,N_29419);
and U33275 (N_33275,N_25713,N_26299);
and U33276 (N_33276,N_26718,N_27685);
or U33277 (N_33277,N_26946,N_27895);
or U33278 (N_33278,N_27209,N_28640);
nor U33279 (N_33279,N_28597,N_26975);
nand U33280 (N_33280,N_26625,N_27451);
or U33281 (N_33281,N_25836,N_26853);
nand U33282 (N_33282,N_29410,N_28000);
nor U33283 (N_33283,N_25762,N_26593);
nand U33284 (N_33284,N_27625,N_29316);
nor U33285 (N_33285,N_29335,N_25438);
nor U33286 (N_33286,N_27944,N_26982);
and U33287 (N_33287,N_25520,N_26177);
nand U33288 (N_33288,N_28300,N_25748);
and U33289 (N_33289,N_29974,N_29041);
nor U33290 (N_33290,N_25816,N_25896);
nor U33291 (N_33291,N_25349,N_27968);
xnor U33292 (N_33292,N_25690,N_28298);
and U33293 (N_33293,N_29204,N_25439);
xnor U33294 (N_33294,N_26945,N_25006);
xnor U33295 (N_33295,N_29523,N_26528);
nand U33296 (N_33296,N_25476,N_29843);
xor U33297 (N_33297,N_26266,N_29492);
nor U33298 (N_33298,N_26109,N_26419);
nand U33299 (N_33299,N_26849,N_29820);
nand U33300 (N_33300,N_29086,N_26812);
and U33301 (N_33301,N_26643,N_27261);
xor U33302 (N_33302,N_25610,N_25950);
nand U33303 (N_33303,N_28765,N_29176);
or U33304 (N_33304,N_27981,N_28886);
xnor U33305 (N_33305,N_25295,N_29222);
or U33306 (N_33306,N_25258,N_27400);
nor U33307 (N_33307,N_28461,N_27050);
and U33308 (N_33308,N_28547,N_29864);
nor U33309 (N_33309,N_29219,N_25542);
nand U33310 (N_33310,N_27646,N_28561);
nor U33311 (N_33311,N_28880,N_25322);
nor U33312 (N_33312,N_27114,N_29680);
nand U33313 (N_33313,N_26458,N_28350);
nor U33314 (N_33314,N_28846,N_26672);
or U33315 (N_33315,N_28965,N_27383);
nor U33316 (N_33316,N_25897,N_29209);
xor U33317 (N_33317,N_29755,N_29552);
nand U33318 (N_33318,N_28954,N_26505);
nand U33319 (N_33319,N_27570,N_26242);
xor U33320 (N_33320,N_27825,N_27711);
or U33321 (N_33321,N_25158,N_29896);
nand U33322 (N_33322,N_25205,N_29104);
nand U33323 (N_33323,N_29983,N_25755);
or U33324 (N_33324,N_29371,N_27666);
or U33325 (N_33325,N_28422,N_29887);
nand U33326 (N_33326,N_28657,N_26165);
nor U33327 (N_33327,N_28367,N_26949);
nor U33328 (N_33328,N_28333,N_25410);
nand U33329 (N_33329,N_25628,N_27438);
or U33330 (N_33330,N_27360,N_25122);
and U33331 (N_33331,N_26047,N_28396);
xor U33332 (N_33332,N_26735,N_27367);
and U33333 (N_33333,N_25742,N_26477);
and U33334 (N_33334,N_28898,N_25437);
and U33335 (N_33335,N_27399,N_29106);
xor U33336 (N_33336,N_28695,N_27682);
or U33337 (N_33337,N_27145,N_28467);
and U33338 (N_33338,N_27243,N_25397);
and U33339 (N_33339,N_26339,N_29635);
nor U33340 (N_33340,N_27775,N_25217);
nand U33341 (N_33341,N_29586,N_27841);
and U33342 (N_33342,N_25408,N_26372);
and U33343 (N_33343,N_26222,N_25881);
and U33344 (N_33344,N_29501,N_29212);
nor U33345 (N_33345,N_25749,N_27270);
and U33346 (N_33346,N_26491,N_26243);
nor U33347 (N_33347,N_26437,N_28687);
nand U33348 (N_33348,N_25711,N_27475);
and U33349 (N_33349,N_27091,N_26701);
and U33350 (N_33350,N_26044,N_28259);
and U33351 (N_33351,N_25411,N_29018);
and U33352 (N_33352,N_25386,N_26042);
xnor U33353 (N_33353,N_26147,N_28562);
nor U33354 (N_33354,N_27123,N_26989);
nand U33355 (N_33355,N_28303,N_28228);
xor U33356 (N_33356,N_28038,N_26206);
and U33357 (N_33357,N_28365,N_25871);
nand U33358 (N_33358,N_28568,N_25647);
nand U33359 (N_33359,N_25699,N_26973);
xor U33360 (N_33360,N_25665,N_29205);
and U33361 (N_33361,N_25495,N_27593);
and U33362 (N_33362,N_28452,N_29243);
and U33363 (N_33363,N_28401,N_28021);
or U33364 (N_33364,N_27616,N_27234);
or U33365 (N_33365,N_26524,N_27493);
and U33366 (N_33366,N_29479,N_26973);
nand U33367 (N_33367,N_27515,N_29368);
xor U33368 (N_33368,N_26255,N_28222);
or U33369 (N_33369,N_25129,N_28319);
nand U33370 (N_33370,N_29862,N_29486);
nand U33371 (N_33371,N_26772,N_27430);
nand U33372 (N_33372,N_29527,N_28862);
xor U33373 (N_33373,N_25696,N_26782);
nor U33374 (N_33374,N_27304,N_29054);
xor U33375 (N_33375,N_28689,N_27783);
or U33376 (N_33376,N_29691,N_27341);
nand U33377 (N_33377,N_29577,N_29432);
or U33378 (N_33378,N_29293,N_27990);
nand U33379 (N_33379,N_27882,N_27087);
xor U33380 (N_33380,N_25896,N_28713);
nor U33381 (N_33381,N_25702,N_28594);
or U33382 (N_33382,N_25320,N_28091);
and U33383 (N_33383,N_27324,N_25809);
nand U33384 (N_33384,N_28854,N_28669);
nand U33385 (N_33385,N_26532,N_29406);
and U33386 (N_33386,N_29613,N_28957);
xor U33387 (N_33387,N_27482,N_26995);
nor U33388 (N_33388,N_26850,N_27718);
or U33389 (N_33389,N_28023,N_25393);
nand U33390 (N_33390,N_28738,N_25754);
or U33391 (N_33391,N_28684,N_25635);
xnor U33392 (N_33392,N_29757,N_26951);
or U33393 (N_33393,N_25587,N_26317);
nand U33394 (N_33394,N_26614,N_28098);
nor U33395 (N_33395,N_29051,N_27230);
or U33396 (N_33396,N_29309,N_29005);
and U33397 (N_33397,N_27191,N_27182);
nor U33398 (N_33398,N_28171,N_25546);
nand U33399 (N_33399,N_25894,N_26315);
xor U33400 (N_33400,N_25363,N_25013);
xor U33401 (N_33401,N_27794,N_25603);
or U33402 (N_33402,N_25792,N_28327);
and U33403 (N_33403,N_28969,N_26895);
or U33404 (N_33404,N_26447,N_26591);
xor U33405 (N_33405,N_28284,N_28657);
xnor U33406 (N_33406,N_26974,N_29391);
nor U33407 (N_33407,N_27658,N_27304);
or U33408 (N_33408,N_28139,N_26498);
or U33409 (N_33409,N_28829,N_26426);
xnor U33410 (N_33410,N_28019,N_28301);
nor U33411 (N_33411,N_26368,N_28113);
nor U33412 (N_33412,N_25760,N_26997);
nand U33413 (N_33413,N_29213,N_27921);
nand U33414 (N_33414,N_25295,N_29893);
xnor U33415 (N_33415,N_25837,N_28496);
nand U33416 (N_33416,N_28514,N_26235);
nor U33417 (N_33417,N_26415,N_29983);
xor U33418 (N_33418,N_28166,N_26014);
or U33419 (N_33419,N_25501,N_26708);
xnor U33420 (N_33420,N_26785,N_28764);
xor U33421 (N_33421,N_28014,N_26592);
and U33422 (N_33422,N_29025,N_26488);
nand U33423 (N_33423,N_29602,N_25146);
xnor U33424 (N_33424,N_28164,N_29944);
or U33425 (N_33425,N_28926,N_26385);
and U33426 (N_33426,N_28091,N_25572);
or U33427 (N_33427,N_28266,N_29216);
and U33428 (N_33428,N_29588,N_26008);
or U33429 (N_33429,N_26054,N_26791);
xnor U33430 (N_33430,N_26985,N_25732);
and U33431 (N_33431,N_27347,N_27606);
nand U33432 (N_33432,N_27543,N_27077);
nand U33433 (N_33433,N_29955,N_28602);
nor U33434 (N_33434,N_28982,N_29590);
nand U33435 (N_33435,N_26376,N_28956);
xor U33436 (N_33436,N_26357,N_27614);
nor U33437 (N_33437,N_27563,N_27296);
and U33438 (N_33438,N_28634,N_29114);
and U33439 (N_33439,N_26018,N_27889);
and U33440 (N_33440,N_25214,N_26976);
nor U33441 (N_33441,N_28769,N_26088);
or U33442 (N_33442,N_29305,N_25485);
xor U33443 (N_33443,N_25102,N_25098);
nand U33444 (N_33444,N_28687,N_25228);
and U33445 (N_33445,N_25251,N_25685);
and U33446 (N_33446,N_28927,N_27878);
and U33447 (N_33447,N_26556,N_29041);
and U33448 (N_33448,N_25280,N_26101);
or U33449 (N_33449,N_25989,N_25626);
xor U33450 (N_33450,N_25761,N_28957);
and U33451 (N_33451,N_26023,N_26360);
nor U33452 (N_33452,N_27310,N_25887);
and U33453 (N_33453,N_28958,N_28693);
or U33454 (N_33454,N_27874,N_26499);
or U33455 (N_33455,N_26607,N_27587);
xnor U33456 (N_33456,N_25621,N_25959);
xor U33457 (N_33457,N_26373,N_26568);
and U33458 (N_33458,N_25661,N_25369);
nor U33459 (N_33459,N_26339,N_27658);
nand U33460 (N_33460,N_28878,N_29154);
xnor U33461 (N_33461,N_28559,N_25510);
nor U33462 (N_33462,N_28926,N_28655);
and U33463 (N_33463,N_26871,N_26932);
or U33464 (N_33464,N_29208,N_26208);
nor U33465 (N_33465,N_25824,N_26088);
and U33466 (N_33466,N_28606,N_27284);
nand U33467 (N_33467,N_29021,N_27743);
xor U33468 (N_33468,N_29977,N_28883);
nand U33469 (N_33469,N_27705,N_26097);
xor U33470 (N_33470,N_26678,N_29510);
nand U33471 (N_33471,N_28164,N_25224);
nor U33472 (N_33472,N_25518,N_25765);
and U33473 (N_33473,N_26312,N_27092);
nand U33474 (N_33474,N_25632,N_28509);
nand U33475 (N_33475,N_28486,N_27006);
nand U33476 (N_33476,N_26801,N_26427);
or U33477 (N_33477,N_28110,N_27909);
and U33478 (N_33478,N_27117,N_28386);
nor U33479 (N_33479,N_25381,N_27559);
xor U33480 (N_33480,N_25111,N_25377);
xor U33481 (N_33481,N_27338,N_28560);
and U33482 (N_33482,N_29889,N_26935);
or U33483 (N_33483,N_28168,N_28150);
nand U33484 (N_33484,N_29207,N_26637);
or U33485 (N_33485,N_28716,N_25687);
xnor U33486 (N_33486,N_25337,N_25027);
nor U33487 (N_33487,N_28741,N_26091);
nor U33488 (N_33488,N_25728,N_27186);
xnor U33489 (N_33489,N_27853,N_26320);
nand U33490 (N_33490,N_27679,N_28184);
and U33491 (N_33491,N_25702,N_27137);
and U33492 (N_33492,N_25894,N_27767);
or U33493 (N_33493,N_29232,N_28864);
nor U33494 (N_33494,N_28901,N_27508);
nor U33495 (N_33495,N_27221,N_25631);
nand U33496 (N_33496,N_26194,N_25344);
xnor U33497 (N_33497,N_29863,N_25497);
xor U33498 (N_33498,N_27646,N_28578);
nor U33499 (N_33499,N_25981,N_25178);
xor U33500 (N_33500,N_29723,N_29898);
or U33501 (N_33501,N_26694,N_26923);
and U33502 (N_33502,N_29223,N_28098);
and U33503 (N_33503,N_29288,N_27135);
nand U33504 (N_33504,N_26059,N_28811);
nand U33505 (N_33505,N_28106,N_29926);
xnor U33506 (N_33506,N_28667,N_27598);
nand U33507 (N_33507,N_29810,N_29141);
nand U33508 (N_33508,N_29208,N_27365);
nor U33509 (N_33509,N_25780,N_29078);
xnor U33510 (N_33510,N_27167,N_26707);
and U33511 (N_33511,N_25334,N_28472);
nor U33512 (N_33512,N_29840,N_25487);
xor U33513 (N_33513,N_29056,N_27550);
nand U33514 (N_33514,N_28197,N_29558);
nor U33515 (N_33515,N_28498,N_28701);
or U33516 (N_33516,N_26503,N_29978);
or U33517 (N_33517,N_28209,N_25732);
nor U33518 (N_33518,N_28960,N_27575);
nand U33519 (N_33519,N_29315,N_27615);
or U33520 (N_33520,N_25954,N_28477);
or U33521 (N_33521,N_28478,N_27098);
nor U33522 (N_33522,N_25996,N_27252);
and U33523 (N_33523,N_27973,N_28131);
nand U33524 (N_33524,N_28087,N_29519);
and U33525 (N_33525,N_26911,N_27302);
nor U33526 (N_33526,N_29001,N_25141);
nor U33527 (N_33527,N_27793,N_25948);
nor U33528 (N_33528,N_29634,N_25477);
and U33529 (N_33529,N_29532,N_29975);
and U33530 (N_33530,N_29280,N_28159);
and U33531 (N_33531,N_28713,N_26953);
nand U33532 (N_33532,N_29201,N_28994);
nand U33533 (N_33533,N_28625,N_29793);
and U33534 (N_33534,N_28977,N_29242);
and U33535 (N_33535,N_29165,N_25785);
nor U33536 (N_33536,N_28721,N_29524);
xnor U33537 (N_33537,N_29237,N_26190);
xor U33538 (N_33538,N_26568,N_25941);
or U33539 (N_33539,N_25806,N_29686);
and U33540 (N_33540,N_29106,N_28284);
nor U33541 (N_33541,N_27739,N_27308);
or U33542 (N_33542,N_28661,N_29140);
and U33543 (N_33543,N_25252,N_28498);
nand U33544 (N_33544,N_26070,N_29791);
nor U33545 (N_33545,N_26796,N_25504);
and U33546 (N_33546,N_27663,N_29852);
nor U33547 (N_33547,N_25626,N_25051);
nand U33548 (N_33548,N_26078,N_25303);
xnor U33549 (N_33549,N_29917,N_28757);
nor U33550 (N_33550,N_29469,N_27854);
nor U33551 (N_33551,N_27838,N_28337);
xnor U33552 (N_33552,N_28537,N_29565);
nor U33553 (N_33553,N_27747,N_25986);
xor U33554 (N_33554,N_28884,N_26488);
xor U33555 (N_33555,N_28558,N_25083);
nor U33556 (N_33556,N_25234,N_27469);
nand U33557 (N_33557,N_29976,N_27679);
nor U33558 (N_33558,N_29066,N_25549);
xnor U33559 (N_33559,N_28063,N_29895);
xnor U33560 (N_33560,N_29368,N_25291);
or U33561 (N_33561,N_26099,N_27908);
and U33562 (N_33562,N_29356,N_29081);
nor U33563 (N_33563,N_25100,N_25753);
or U33564 (N_33564,N_29307,N_25114);
nor U33565 (N_33565,N_29830,N_26891);
nand U33566 (N_33566,N_26377,N_29600);
nor U33567 (N_33567,N_27863,N_25695);
or U33568 (N_33568,N_25931,N_26779);
or U33569 (N_33569,N_28553,N_29857);
or U33570 (N_33570,N_25560,N_28161);
nand U33571 (N_33571,N_28694,N_29610);
or U33572 (N_33572,N_28585,N_26528);
xnor U33573 (N_33573,N_27758,N_28850);
nor U33574 (N_33574,N_29786,N_26382);
or U33575 (N_33575,N_25698,N_29727);
xor U33576 (N_33576,N_25525,N_28930);
and U33577 (N_33577,N_26241,N_28970);
nand U33578 (N_33578,N_25856,N_26831);
nor U33579 (N_33579,N_28019,N_29520);
xnor U33580 (N_33580,N_26344,N_25099);
or U33581 (N_33581,N_29499,N_25644);
nand U33582 (N_33582,N_25538,N_27664);
or U33583 (N_33583,N_25733,N_27687);
and U33584 (N_33584,N_26788,N_26043);
nand U33585 (N_33585,N_29249,N_28632);
nand U33586 (N_33586,N_29557,N_27012);
xor U33587 (N_33587,N_25894,N_29288);
xor U33588 (N_33588,N_29738,N_28433);
nand U33589 (N_33589,N_29261,N_26878);
nand U33590 (N_33590,N_26029,N_26812);
or U33591 (N_33591,N_28383,N_26923);
xnor U33592 (N_33592,N_27048,N_28842);
and U33593 (N_33593,N_27411,N_28799);
and U33594 (N_33594,N_27550,N_28784);
nor U33595 (N_33595,N_27820,N_26867);
xor U33596 (N_33596,N_29611,N_25092);
nand U33597 (N_33597,N_28883,N_26876);
and U33598 (N_33598,N_26690,N_26453);
nor U33599 (N_33599,N_27036,N_29501);
nand U33600 (N_33600,N_28743,N_28054);
xnor U33601 (N_33601,N_26201,N_28423);
nor U33602 (N_33602,N_29023,N_27453);
nand U33603 (N_33603,N_29515,N_27161);
or U33604 (N_33604,N_28512,N_27664);
and U33605 (N_33605,N_29516,N_29546);
xor U33606 (N_33606,N_25007,N_25171);
or U33607 (N_33607,N_25707,N_29172);
nor U33608 (N_33608,N_27524,N_27458);
nand U33609 (N_33609,N_29870,N_29106);
and U33610 (N_33610,N_29446,N_28978);
xor U33611 (N_33611,N_25011,N_25624);
nand U33612 (N_33612,N_25414,N_27452);
or U33613 (N_33613,N_26628,N_27139);
xor U33614 (N_33614,N_27355,N_28873);
xnor U33615 (N_33615,N_28202,N_29402);
nor U33616 (N_33616,N_28914,N_28208);
nor U33617 (N_33617,N_27495,N_27883);
nor U33618 (N_33618,N_28824,N_26149);
nor U33619 (N_33619,N_27302,N_26483);
and U33620 (N_33620,N_27754,N_27661);
and U33621 (N_33621,N_25160,N_28291);
nand U33622 (N_33622,N_25721,N_29358);
and U33623 (N_33623,N_29393,N_27587);
or U33624 (N_33624,N_26563,N_27634);
nor U33625 (N_33625,N_27943,N_27825);
or U33626 (N_33626,N_29149,N_25691);
nor U33627 (N_33627,N_28245,N_26933);
or U33628 (N_33628,N_27924,N_29682);
and U33629 (N_33629,N_28069,N_29151);
nand U33630 (N_33630,N_25467,N_27633);
nor U33631 (N_33631,N_25490,N_25414);
nand U33632 (N_33632,N_26047,N_28903);
xor U33633 (N_33633,N_29776,N_27940);
or U33634 (N_33634,N_25231,N_29411);
nand U33635 (N_33635,N_28230,N_25774);
xor U33636 (N_33636,N_26719,N_25329);
xnor U33637 (N_33637,N_26279,N_29462);
and U33638 (N_33638,N_27897,N_28828);
xor U33639 (N_33639,N_29835,N_27721);
nand U33640 (N_33640,N_29202,N_28550);
nand U33641 (N_33641,N_29506,N_26192);
xor U33642 (N_33642,N_26012,N_27415);
and U33643 (N_33643,N_29534,N_28325);
or U33644 (N_33644,N_27872,N_29556);
and U33645 (N_33645,N_25037,N_29597);
nand U33646 (N_33646,N_28072,N_27152);
xor U33647 (N_33647,N_27384,N_25462);
xnor U33648 (N_33648,N_25317,N_25557);
nor U33649 (N_33649,N_29985,N_29908);
and U33650 (N_33650,N_29216,N_26140);
xor U33651 (N_33651,N_26933,N_26716);
nand U33652 (N_33652,N_26438,N_26379);
nand U33653 (N_33653,N_28302,N_28661);
or U33654 (N_33654,N_29594,N_28518);
or U33655 (N_33655,N_26063,N_29418);
nand U33656 (N_33656,N_29410,N_26817);
and U33657 (N_33657,N_29487,N_29775);
xnor U33658 (N_33658,N_27652,N_25252);
or U33659 (N_33659,N_28187,N_27760);
nor U33660 (N_33660,N_29164,N_28756);
and U33661 (N_33661,N_28681,N_28845);
and U33662 (N_33662,N_27005,N_26398);
xor U33663 (N_33663,N_26003,N_27309);
xor U33664 (N_33664,N_29025,N_28693);
nand U33665 (N_33665,N_27639,N_28783);
xor U33666 (N_33666,N_26570,N_29342);
nor U33667 (N_33667,N_27203,N_29784);
nand U33668 (N_33668,N_27361,N_26849);
nor U33669 (N_33669,N_25338,N_27179);
nor U33670 (N_33670,N_27491,N_27952);
nand U33671 (N_33671,N_25833,N_25922);
nor U33672 (N_33672,N_27518,N_25307);
or U33673 (N_33673,N_25428,N_25455);
nor U33674 (N_33674,N_26011,N_29365);
or U33675 (N_33675,N_28700,N_28874);
and U33676 (N_33676,N_28986,N_29521);
xor U33677 (N_33677,N_26462,N_26779);
nor U33678 (N_33678,N_28285,N_28931);
nand U33679 (N_33679,N_25818,N_27952);
nand U33680 (N_33680,N_25934,N_29013);
xor U33681 (N_33681,N_26326,N_27604);
or U33682 (N_33682,N_27139,N_25181);
and U33683 (N_33683,N_29957,N_27873);
xnor U33684 (N_33684,N_25715,N_28282);
xor U33685 (N_33685,N_28927,N_28349);
xor U33686 (N_33686,N_28482,N_28311);
xnor U33687 (N_33687,N_25785,N_28025);
nand U33688 (N_33688,N_28306,N_28549);
and U33689 (N_33689,N_25410,N_28315);
nand U33690 (N_33690,N_26647,N_27201);
nand U33691 (N_33691,N_28993,N_27063);
nor U33692 (N_33692,N_26760,N_26386);
or U33693 (N_33693,N_26345,N_29530);
or U33694 (N_33694,N_25438,N_27980);
and U33695 (N_33695,N_26236,N_29361);
and U33696 (N_33696,N_28890,N_26790);
or U33697 (N_33697,N_29331,N_29930);
nand U33698 (N_33698,N_25352,N_26978);
or U33699 (N_33699,N_25869,N_29991);
nor U33700 (N_33700,N_25589,N_29801);
xor U33701 (N_33701,N_26557,N_25134);
nand U33702 (N_33702,N_28658,N_27047);
nor U33703 (N_33703,N_26918,N_28548);
xnor U33704 (N_33704,N_28556,N_25919);
and U33705 (N_33705,N_29701,N_27424);
and U33706 (N_33706,N_27274,N_28750);
nand U33707 (N_33707,N_27671,N_27995);
nand U33708 (N_33708,N_27657,N_25710);
nor U33709 (N_33709,N_27391,N_27434);
or U33710 (N_33710,N_28042,N_26054);
nand U33711 (N_33711,N_27943,N_26899);
nand U33712 (N_33712,N_25126,N_28334);
nand U33713 (N_33713,N_25876,N_27291);
xnor U33714 (N_33714,N_26421,N_28475);
and U33715 (N_33715,N_27081,N_27490);
and U33716 (N_33716,N_26025,N_29416);
nor U33717 (N_33717,N_25012,N_28410);
nor U33718 (N_33718,N_28636,N_27818);
nor U33719 (N_33719,N_27207,N_25375);
xor U33720 (N_33720,N_26103,N_28665);
nand U33721 (N_33721,N_29524,N_28372);
and U33722 (N_33722,N_28146,N_26401);
and U33723 (N_33723,N_29659,N_25134);
xnor U33724 (N_33724,N_28112,N_27862);
or U33725 (N_33725,N_27140,N_27488);
or U33726 (N_33726,N_28446,N_25728);
nor U33727 (N_33727,N_25435,N_27075);
or U33728 (N_33728,N_29323,N_29611);
and U33729 (N_33729,N_28810,N_26801);
or U33730 (N_33730,N_29210,N_28752);
xor U33731 (N_33731,N_28183,N_27655);
or U33732 (N_33732,N_28245,N_27335);
and U33733 (N_33733,N_26501,N_26312);
nor U33734 (N_33734,N_26335,N_26371);
and U33735 (N_33735,N_28883,N_25036);
xor U33736 (N_33736,N_26912,N_25111);
or U33737 (N_33737,N_27979,N_28997);
nor U33738 (N_33738,N_28294,N_28859);
xnor U33739 (N_33739,N_28709,N_29861);
and U33740 (N_33740,N_25879,N_25770);
nor U33741 (N_33741,N_26461,N_26542);
or U33742 (N_33742,N_25544,N_27315);
or U33743 (N_33743,N_27980,N_26889);
or U33744 (N_33744,N_26614,N_27440);
and U33745 (N_33745,N_25812,N_27725);
nor U33746 (N_33746,N_26237,N_27296);
nand U33747 (N_33747,N_26149,N_28243);
nor U33748 (N_33748,N_26289,N_29791);
nand U33749 (N_33749,N_26638,N_25929);
xor U33750 (N_33750,N_29867,N_26426);
nor U33751 (N_33751,N_27373,N_25451);
nor U33752 (N_33752,N_26998,N_29728);
or U33753 (N_33753,N_27531,N_26109);
xnor U33754 (N_33754,N_29584,N_28636);
xnor U33755 (N_33755,N_28424,N_27823);
nand U33756 (N_33756,N_29735,N_28015);
and U33757 (N_33757,N_25228,N_27374);
xnor U33758 (N_33758,N_29144,N_28179);
and U33759 (N_33759,N_29370,N_29120);
and U33760 (N_33760,N_25392,N_27545);
xnor U33761 (N_33761,N_28640,N_25251);
and U33762 (N_33762,N_28451,N_29835);
xor U33763 (N_33763,N_26624,N_25124);
or U33764 (N_33764,N_27994,N_27502);
and U33765 (N_33765,N_29401,N_28127);
nand U33766 (N_33766,N_25312,N_29586);
nor U33767 (N_33767,N_25802,N_28490);
nand U33768 (N_33768,N_29078,N_28089);
xnor U33769 (N_33769,N_28342,N_29811);
xnor U33770 (N_33770,N_26345,N_29204);
or U33771 (N_33771,N_26541,N_25273);
xor U33772 (N_33772,N_25841,N_28920);
and U33773 (N_33773,N_27753,N_28148);
or U33774 (N_33774,N_26849,N_27182);
xnor U33775 (N_33775,N_28552,N_27895);
and U33776 (N_33776,N_25708,N_29207);
and U33777 (N_33777,N_25332,N_26815);
nor U33778 (N_33778,N_29696,N_26045);
and U33779 (N_33779,N_28166,N_28018);
xnor U33780 (N_33780,N_28029,N_29983);
and U33781 (N_33781,N_27567,N_27009);
and U33782 (N_33782,N_28657,N_26771);
nor U33783 (N_33783,N_28068,N_28015);
nor U33784 (N_33784,N_28903,N_28028);
and U33785 (N_33785,N_25101,N_29840);
nand U33786 (N_33786,N_28588,N_25919);
or U33787 (N_33787,N_28426,N_29485);
and U33788 (N_33788,N_26668,N_25795);
and U33789 (N_33789,N_25478,N_29907);
nand U33790 (N_33790,N_26945,N_29394);
nor U33791 (N_33791,N_26301,N_27879);
or U33792 (N_33792,N_26911,N_25543);
and U33793 (N_33793,N_25877,N_26140);
nand U33794 (N_33794,N_28674,N_27590);
and U33795 (N_33795,N_29916,N_28730);
nor U33796 (N_33796,N_29653,N_27379);
nand U33797 (N_33797,N_29551,N_26897);
and U33798 (N_33798,N_27518,N_26126);
xor U33799 (N_33799,N_28061,N_27957);
nand U33800 (N_33800,N_25511,N_27125);
or U33801 (N_33801,N_26470,N_26969);
and U33802 (N_33802,N_25732,N_28360);
nor U33803 (N_33803,N_28213,N_28205);
nor U33804 (N_33804,N_26169,N_28915);
or U33805 (N_33805,N_27031,N_29596);
nand U33806 (N_33806,N_26679,N_25438);
or U33807 (N_33807,N_29662,N_27066);
and U33808 (N_33808,N_25955,N_26857);
nand U33809 (N_33809,N_25565,N_26869);
and U33810 (N_33810,N_28368,N_26867);
and U33811 (N_33811,N_27759,N_25884);
nand U33812 (N_33812,N_25630,N_26911);
nand U33813 (N_33813,N_29727,N_28939);
or U33814 (N_33814,N_29378,N_29749);
xnor U33815 (N_33815,N_27505,N_25471);
or U33816 (N_33816,N_27598,N_28709);
xor U33817 (N_33817,N_26792,N_27711);
and U33818 (N_33818,N_25577,N_29870);
xnor U33819 (N_33819,N_25524,N_25801);
and U33820 (N_33820,N_29248,N_26907);
nor U33821 (N_33821,N_25776,N_26315);
nor U33822 (N_33822,N_29592,N_25089);
and U33823 (N_33823,N_29691,N_29684);
nor U33824 (N_33824,N_26514,N_25035);
and U33825 (N_33825,N_28189,N_27035);
or U33826 (N_33826,N_29272,N_25108);
or U33827 (N_33827,N_26438,N_27127);
or U33828 (N_33828,N_28258,N_29401);
nand U33829 (N_33829,N_27372,N_26954);
nor U33830 (N_33830,N_29708,N_28437);
nand U33831 (N_33831,N_27474,N_28701);
xnor U33832 (N_33832,N_28712,N_29658);
nor U33833 (N_33833,N_29429,N_25492);
xnor U33834 (N_33834,N_25411,N_25607);
and U33835 (N_33835,N_29776,N_29585);
xnor U33836 (N_33836,N_26666,N_26615);
and U33837 (N_33837,N_29775,N_27128);
nand U33838 (N_33838,N_25488,N_26894);
xnor U33839 (N_33839,N_26025,N_28189);
or U33840 (N_33840,N_28477,N_26314);
nor U33841 (N_33841,N_28971,N_26774);
or U33842 (N_33842,N_28012,N_28617);
and U33843 (N_33843,N_28549,N_25513);
xor U33844 (N_33844,N_27115,N_26141);
nor U33845 (N_33845,N_28053,N_27875);
and U33846 (N_33846,N_26818,N_25637);
and U33847 (N_33847,N_27101,N_27245);
and U33848 (N_33848,N_27857,N_29838);
and U33849 (N_33849,N_25786,N_27682);
or U33850 (N_33850,N_29962,N_28235);
nand U33851 (N_33851,N_26508,N_25273);
nand U33852 (N_33852,N_28005,N_27181);
nor U33853 (N_33853,N_25207,N_29859);
nor U33854 (N_33854,N_27901,N_28184);
nand U33855 (N_33855,N_25189,N_25635);
or U33856 (N_33856,N_27853,N_29925);
xnor U33857 (N_33857,N_26395,N_26490);
or U33858 (N_33858,N_27465,N_26560);
and U33859 (N_33859,N_26985,N_29474);
or U33860 (N_33860,N_26103,N_25251);
xnor U33861 (N_33861,N_29791,N_25166);
or U33862 (N_33862,N_26047,N_25227);
and U33863 (N_33863,N_28420,N_27333);
nor U33864 (N_33864,N_29451,N_28481);
and U33865 (N_33865,N_26889,N_29310);
xnor U33866 (N_33866,N_28234,N_27015);
and U33867 (N_33867,N_26869,N_29633);
xor U33868 (N_33868,N_27667,N_27227);
nor U33869 (N_33869,N_27610,N_28379);
nand U33870 (N_33870,N_26290,N_26933);
or U33871 (N_33871,N_25994,N_25651);
and U33872 (N_33872,N_26149,N_28902);
or U33873 (N_33873,N_25877,N_25744);
nor U33874 (N_33874,N_27277,N_27684);
nand U33875 (N_33875,N_25221,N_27643);
xnor U33876 (N_33876,N_28572,N_26208);
and U33877 (N_33877,N_29201,N_26010);
nand U33878 (N_33878,N_27179,N_29587);
or U33879 (N_33879,N_25582,N_29006);
or U33880 (N_33880,N_25805,N_25539);
nand U33881 (N_33881,N_29837,N_26349);
or U33882 (N_33882,N_25154,N_27365);
nor U33883 (N_33883,N_29790,N_29068);
nand U33884 (N_33884,N_28575,N_28536);
or U33885 (N_33885,N_29871,N_28435);
xor U33886 (N_33886,N_25562,N_25901);
xnor U33887 (N_33887,N_25115,N_26602);
nor U33888 (N_33888,N_29471,N_25842);
xnor U33889 (N_33889,N_28766,N_27432);
nor U33890 (N_33890,N_25845,N_28187);
nand U33891 (N_33891,N_27739,N_29074);
and U33892 (N_33892,N_27118,N_28412);
nor U33893 (N_33893,N_29909,N_27276);
xnor U33894 (N_33894,N_29501,N_27449);
xnor U33895 (N_33895,N_26273,N_25450);
and U33896 (N_33896,N_25516,N_29569);
nand U33897 (N_33897,N_26963,N_25976);
xnor U33898 (N_33898,N_29901,N_28166);
nor U33899 (N_33899,N_27110,N_28419);
nor U33900 (N_33900,N_27122,N_27958);
or U33901 (N_33901,N_26581,N_28692);
and U33902 (N_33902,N_25732,N_28577);
xor U33903 (N_33903,N_29782,N_28015);
or U33904 (N_33904,N_28415,N_25748);
and U33905 (N_33905,N_29373,N_27504);
and U33906 (N_33906,N_27755,N_27531);
nor U33907 (N_33907,N_27149,N_25103);
and U33908 (N_33908,N_27044,N_28400);
xnor U33909 (N_33909,N_25282,N_25166);
nand U33910 (N_33910,N_28016,N_25461);
nand U33911 (N_33911,N_27311,N_28873);
or U33912 (N_33912,N_29376,N_26937);
nor U33913 (N_33913,N_25594,N_25132);
or U33914 (N_33914,N_29243,N_29305);
xnor U33915 (N_33915,N_26815,N_27538);
or U33916 (N_33916,N_25591,N_26920);
and U33917 (N_33917,N_29951,N_29988);
nand U33918 (N_33918,N_27977,N_27869);
and U33919 (N_33919,N_25340,N_29644);
nand U33920 (N_33920,N_26779,N_27863);
or U33921 (N_33921,N_28852,N_25781);
nor U33922 (N_33922,N_28118,N_27886);
xnor U33923 (N_33923,N_28282,N_29793);
or U33924 (N_33924,N_29904,N_27486);
and U33925 (N_33925,N_28908,N_29413);
and U33926 (N_33926,N_26558,N_29495);
and U33927 (N_33927,N_29178,N_29258);
nand U33928 (N_33928,N_28963,N_26177);
nand U33929 (N_33929,N_25416,N_26720);
nor U33930 (N_33930,N_29197,N_28152);
nor U33931 (N_33931,N_29511,N_25449);
nand U33932 (N_33932,N_26977,N_29574);
nor U33933 (N_33933,N_25563,N_26187);
xor U33934 (N_33934,N_28327,N_26663);
nor U33935 (N_33935,N_29368,N_27798);
nor U33936 (N_33936,N_28521,N_29614);
xor U33937 (N_33937,N_27569,N_25256);
and U33938 (N_33938,N_28545,N_26760);
nor U33939 (N_33939,N_29777,N_25689);
and U33940 (N_33940,N_29539,N_27325);
and U33941 (N_33941,N_26812,N_27540);
xnor U33942 (N_33942,N_28728,N_29675);
nand U33943 (N_33943,N_26611,N_29610);
xnor U33944 (N_33944,N_26692,N_29886);
or U33945 (N_33945,N_25714,N_26992);
and U33946 (N_33946,N_28521,N_28623);
xnor U33947 (N_33947,N_28113,N_26660);
or U33948 (N_33948,N_26014,N_25639);
nor U33949 (N_33949,N_29598,N_25476);
xor U33950 (N_33950,N_26785,N_28925);
and U33951 (N_33951,N_26518,N_27011);
nand U33952 (N_33952,N_28256,N_26645);
nor U33953 (N_33953,N_26523,N_25500);
nor U33954 (N_33954,N_27324,N_25636);
or U33955 (N_33955,N_27611,N_28447);
or U33956 (N_33956,N_25163,N_26492);
and U33957 (N_33957,N_25800,N_29507);
or U33958 (N_33958,N_29066,N_26590);
and U33959 (N_33959,N_29918,N_27826);
nand U33960 (N_33960,N_29242,N_26797);
and U33961 (N_33961,N_28848,N_29082);
xor U33962 (N_33962,N_26434,N_28569);
nor U33963 (N_33963,N_25497,N_27662);
and U33964 (N_33964,N_29875,N_26204);
nor U33965 (N_33965,N_28977,N_25565);
and U33966 (N_33966,N_29547,N_29162);
or U33967 (N_33967,N_28059,N_25054);
or U33968 (N_33968,N_28868,N_25705);
or U33969 (N_33969,N_28862,N_26578);
and U33970 (N_33970,N_26016,N_28058);
or U33971 (N_33971,N_29785,N_25590);
and U33972 (N_33972,N_29561,N_26932);
xor U33973 (N_33973,N_25406,N_28076);
xnor U33974 (N_33974,N_25099,N_25274);
or U33975 (N_33975,N_26026,N_27586);
nand U33976 (N_33976,N_25548,N_26703);
xor U33977 (N_33977,N_27586,N_25037);
nor U33978 (N_33978,N_26655,N_28111);
and U33979 (N_33979,N_26249,N_25039);
xor U33980 (N_33980,N_26569,N_28452);
nor U33981 (N_33981,N_28885,N_26717);
or U33982 (N_33982,N_27075,N_25673);
and U33983 (N_33983,N_26779,N_29799);
xnor U33984 (N_33984,N_25347,N_28576);
xor U33985 (N_33985,N_26876,N_28970);
and U33986 (N_33986,N_28112,N_28865);
or U33987 (N_33987,N_27747,N_28544);
and U33988 (N_33988,N_28014,N_29752);
and U33989 (N_33989,N_29677,N_25564);
and U33990 (N_33990,N_27346,N_26635);
nor U33991 (N_33991,N_29200,N_28691);
xor U33992 (N_33992,N_27213,N_26747);
or U33993 (N_33993,N_29432,N_25237);
nor U33994 (N_33994,N_25326,N_29147);
xor U33995 (N_33995,N_29011,N_27533);
nor U33996 (N_33996,N_28846,N_26702);
nand U33997 (N_33997,N_29984,N_26884);
or U33998 (N_33998,N_29689,N_29494);
xor U33999 (N_33999,N_29770,N_27415);
xor U34000 (N_34000,N_26373,N_28105);
and U34001 (N_34001,N_29306,N_26953);
or U34002 (N_34002,N_27136,N_25729);
and U34003 (N_34003,N_26159,N_28728);
nor U34004 (N_34004,N_27462,N_27567);
nand U34005 (N_34005,N_25430,N_26250);
and U34006 (N_34006,N_28274,N_29508);
and U34007 (N_34007,N_25127,N_25906);
xor U34008 (N_34008,N_29835,N_29769);
nand U34009 (N_34009,N_27496,N_29784);
xor U34010 (N_34010,N_28335,N_29711);
xnor U34011 (N_34011,N_29757,N_29265);
nand U34012 (N_34012,N_28901,N_28470);
or U34013 (N_34013,N_25895,N_25797);
and U34014 (N_34014,N_28951,N_29402);
nor U34015 (N_34015,N_27440,N_26761);
nor U34016 (N_34016,N_25094,N_26590);
xnor U34017 (N_34017,N_29476,N_25660);
and U34018 (N_34018,N_28359,N_28673);
or U34019 (N_34019,N_28339,N_26265);
and U34020 (N_34020,N_26314,N_29041);
nand U34021 (N_34021,N_28254,N_25070);
xor U34022 (N_34022,N_26274,N_27416);
and U34023 (N_34023,N_26554,N_27838);
nand U34024 (N_34024,N_25930,N_28737);
nand U34025 (N_34025,N_28480,N_28333);
nand U34026 (N_34026,N_29147,N_26537);
or U34027 (N_34027,N_26157,N_27802);
xnor U34028 (N_34028,N_26521,N_28880);
or U34029 (N_34029,N_26636,N_28535);
nand U34030 (N_34030,N_25284,N_28904);
xnor U34031 (N_34031,N_25915,N_27168);
xnor U34032 (N_34032,N_28977,N_25717);
or U34033 (N_34033,N_26705,N_25419);
nor U34034 (N_34034,N_27953,N_26810);
and U34035 (N_34035,N_27168,N_28554);
xnor U34036 (N_34036,N_28307,N_29962);
and U34037 (N_34037,N_29864,N_28860);
and U34038 (N_34038,N_25528,N_28892);
or U34039 (N_34039,N_29468,N_26235);
or U34040 (N_34040,N_25011,N_25645);
or U34041 (N_34041,N_26558,N_26678);
nor U34042 (N_34042,N_28893,N_28298);
xor U34043 (N_34043,N_25914,N_27606);
nor U34044 (N_34044,N_29223,N_25917);
and U34045 (N_34045,N_25066,N_29178);
or U34046 (N_34046,N_28244,N_25136);
xor U34047 (N_34047,N_29928,N_27279);
xor U34048 (N_34048,N_27748,N_25419);
nor U34049 (N_34049,N_27703,N_28311);
xor U34050 (N_34050,N_29066,N_25462);
and U34051 (N_34051,N_27147,N_28435);
nand U34052 (N_34052,N_26011,N_27664);
nor U34053 (N_34053,N_26528,N_29565);
nor U34054 (N_34054,N_25204,N_27991);
xor U34055 (N_34055,N_25284,N_27761);
or U34056 (N_34056,N_28143,N_28993);
and U34057 (N_34057,N_27342,N_25761);
xor U34058 (N_34058,N_26837,N_27518);
and U34059 (N_34059,N_29675,N_28600);
or U34060 (N_34060,N_27138,N_29665);
nand U34061 (N_34061,N_28618,N_25560);
xnor U34062 (N_34062,N_29327,N_27705);
or U34063 (N_34063,N_27310,N_28538);
nand U34064 (N_34064,N_27935,N_29490);
or U34065 (N_34065,N_28368,N_27510);
xnor U34066 (N_34066,N_28661,N_27984);
and U34067 (N_34067,N_28082,N_29576);
nor U34068 (N_34068,N_27316,N_27206);
and U34069 (N_34069,N_26797,N_25857);
or U34070 (N_34070,N_27644,N_25002);
or U34071 (N_34071,N_27527,N_27719);
or U34072 (N_34072,N_27163,N_28214);
and U34073 (N_34073,N_27966,N_29516);
or U34074 (N_34074,N_27811,N_26737);
and U34075 (N_34075,N_25795,N_27330);
nor U34076 (N_34076,N_28863,N_28788);
nand U34077 (N_34077,N_29779,N_29770);
and U34078 (N_34078,N_26214,N_29771);
nor U34079 (N_34079,N_29520,N_25214);
nor U34080 (N_34080,N_26285,N_27583);
xnor U34081 (N_34081,N_25932,N_26351);
nor U34082 (N_34082,N_29165,N_29408);
xnor U34083 (N_34083,N_26322,N_29366);
or U34084 (N_34084,N_25383,N_27457);
xor U34085 (N_34085,N_27274,N_28165);
and U34086 (N_34086,N_25024,N_28479);
nand U34087 (N_34087,N_27935,N_26712);
nor U34088 (N_34088,N_27550,N_26493);
nor U34089 (N_34089,N_26444,N_28844);
and U34090 (N_34090,N_26318,N_25959);
nor U34091 (N_34091,N_25226,N_29166);
xor U34092 (N_34092,N_27313,N_27670);
or U34093 (N_34093,N_25588,N_28874);
nor U34094 (N_34094,N_26856,N_25151);
or U34095 (N_34095,N_25365,N_25658);
nor U34096 (N_34096,N_28001,N_29933);
or U34097 (N_34097,N_27835,N_27063);
or U34098 (N_34098,N_25724,N_26003);
or U34099 (N_34099,N_29233,N_26989);
nand U34100 (N_34100,N_28074,N_28241);
or U34101 (N_34101,N_29968,N_27301);
nand U34102 (N_34102,N_27880,N_29370);
or U34103 (N_34103,N_25884,N_29150);
nand U34104 (N_34104,N_25488,N_26970);
nor U34105 (N_34105,N_26727,N_26582);
and U34106 (N_34106,N_25728,N_29591);
nor U34107 (N_34107,N_26514,N_29862);
xor U34108 (N_34108,N_27413,N_25420);
nor U34109 (N_34109,N_26326,N_29034);
or U34110 (N_34110,N_29452,N_26712);
or U34111 (N_34111,N_25941,N_25496);
and U34112 (N_34112,N_28183,N_28900);
or U34113 (N_34113,N_26929,N_25050);
and U34114 (N_34114,N_29198,N_28191);
and U34115 (N_34115,N_25507,N_27169);
nand U34116 (N_34116,N_29619,N_26836);
nand U34117 (N_34117,N_28022,N_28095);
nor U34118 (N_34118,N_28049,N_27695);
and U34119 (N_34119,N_26659,N_26048);
and U34120 (N_34120,N_26548,N_28553);
xnor U34121 (N_34121,N_29331,N_29380);
and U34122 (N_34122,N_27272,N_25723);
nor U34123 (N_34123,N_27721,N_29712);
nand U34124 (N_34124,N_28856,N_29613);
nor U34125 (N_34125,N_27529,N_26038);
and U34126 (N_34126,N_27369,N_26185);
or U34127 (N_34127,N_28904,N_28966);
xor U34128 (N_34128,N_26414,N_27949);
or U34129 (N_34129,N_26196,N_27759);
nand U34130 (N_34130,N_25383,N_26625);
or U34131 (N_34131,N_27718,N_25411);
nor U34132 (N_34132,N_28278,N_28579);
xnor U34133 (N_34133,N_26498,N_25786);
or U34134 (N_34134,N_25122,N_27533);
or U34135 (N_34135,N_26752,N_25047);
or U34136 (N_34136,N_25883,N_26531);
nand U34137 (N_34137,N_27559,N_25328);
nand U34138 (N_34138,N_26246,N_25647);
nor U34139 (N_34139,N_28632,N_25940);
nor U34140 (N_34140,N_27521,N_28429);
or U34141 (N_34141,N_25400,N_26749);
xnor U34142 (N_34142,N_25203,N_29016);
and U34143 (N_34143,N_25016,N_26774);
and U34144 (N_34144,N_25116,N_26621);
and U34145 (N_34145,N_28466,N_25491);
and U34146 (N_34146,N_27793,N_26439);
and U34147 (N_34147,N_25626,N_28076);
nor U34148 (N_34148,N_29753,N_28615);
nor U34149 (N_34149,N_25327,N_27019);
nand U34150 (N_34150,N_29376,N_25320);
or U34151 (N_34151,N_29066,N_28069);
or U34152 (N_34152,N_29616,N_28947);
nand U34153 (N_34153,N_27449,N_27461);
xnor U34154 (N_34154,N_25903,N_27052);
xor U34155 (N_34155,N_28999,N_29994);
nor U34156 (N_34156,N_29110,N_27576);
xnor U34157 (N_34157,N_28377,N_26799);
nand U34158 (N_34158,N_27459,N_25198);
and U34159 (N_34159,N_28660,N_25863);
nor U34160 (N_34160,N_29008,N_26860);
nor U34161 (N_34161,N_28637,N_26681);
and U34162 (N_34162,N_26113,N_26238);
xnor U34163 (N_34163,N_29325,N_27083);
nand U34164 (N_34164,N_27342,N_29221);
xor U34165 (N_34165,N_25146,N_26217);
nand U34166 (N_34166,N_25575,N_27833);
or U34167 (N_34167,N_26602,N_28779);
nand U34168 (N_34168,N_28899,N_25854);
nor U34169 (N_34169,N_26998,N_27614);
nor U34170 (N_34170,N_27181,N_28192);
nand U34171 (N_34171,N_29131,N_26702);
or U34172 (N_34172,N_28864,N_27591);
xnor U34173 (N_34173,N_26483,N_27572);
nand U34174 (N_34174,N_26472,N_27733);
xor U34175 (N_34175,N_28068,N_25433);
nor U34176 (N_34176,N_25049,N_29969);
nand U34177 (N_34177,N_26241,N_27032);
nand U34178 (N_34178,N_25951,N_27637);
or U34179 (N_34179,N_28183,N_27641);
nand U34180 (N_34180,N_29963,N_26241);
xnor U34181 (N_34181,N_29562,N_25109);
nor U34182 (N_34182,N_27111,N_29061);
or U34183 (N_34183,N_27736,N_28189);
nor U34184 (N_34184,N_26186,N_26300);
nand U34185 (N_34185,N_25568,N_29443);
nand U34186 (N_34186,N_26603,N_25584);
or U34187 (N_34187,N_25990,N_29287);
and U34188 (N_34188,N_28020,N_25669);
xnor U34189 (N_34189,N_26805,N_26088);
nand U34190 (N_34190,N_29315,N_25594);
xor U34191 (N_34191,N_26394,N_27221);
and U34192 (N_34192,N_26847,N_25632);
and U34193 (N_34193,N_27549,N_26993);
or U34194 (N_34194,N_26666,N_29444);
nand U34195 (N_34195,N_28002,N_27833);
xor U34196 (N_34196,N_25797,N_28639);
nor U34197 (N_34197,N_25203,N_26699);
nand U34198 (N_34198,N_26851,N_25636);
nor U34199 (N_34199,N_26315,N_25610);
nand U34200 (N_34200,N_26174,N_25272);
or U34201 (N_34201,N_25845,N_25822);
or U34202 (N_34202,N_26406,N_26464);
xnor U34203 (N_34203,N_29520,N_27958);
xnor U34204 (N_34204,N_26111,N_25675);
nor U34205 (N_34205,N_28458,N_27998);
and U34206 (N_34206,N_28469,N_27225);
and U34207 (N_34207,N_27361,N_28048);
and U34208 (N_34208,N_28620,N_29512);
and U34209 (N_34209,N_29018,N_28557);
nor U34210 (N_34210,N_25276,N_28379);
nand U34211 (N_34211,N_26897,N_27893);
or U34212 (N_34212,N_29636,N_26924);
and U34213 (N_34213,N_25881,N_28840);
xor U34214 (N_34214,N_26134,N_26981);
and U34215 (N_34215,N_26499,N_29068);
or U34216 (N_34216,N_26038,N_27944);
xor U34217 (N_34217,N_28937,N_26661);
nor U34218 (N_34218,N_29126,N_26586);
xnor U34219 (N_34219,N_28365,N_29976);
and U34220 (N_34220,N_28376,N_25342);
and U34221 (N_34221,N_29051,N_26859);
nor U34222 (N_34222,N_28666,N_26810);
xor U34223 (N_34223,N_28734,N_26392);
nor U34224 (N_34224,N_28094,N_26389);
nor U34225 (N_34225,N_28163,N_25760);
nand U34226 (N_34226,N_27666,N_29632);
nor U34227 (N_34227,N_27560,N_26031);
nor U34228 (N_34228,N_29696,N_27937);
or U34229 (N_34229,N_29212,N_26216);
or U34230 (N_34230,N_28854,N_25952);
and U34231 (N_34231,N_27633,N_28495);
and U34232 (N_34232,N_26533,N_27819);
nand U34233 (N_34233,N_29279,N_29609);
nor U34234 (N_34234,N_29639,N_26390);
and U34235 (N_34235,N_25058,N_28450);
nand U34236 (N_34236,N_29791,N_29184);
nor U34237 (N_34237,N_28721,N_28447);
or U34238 (N_34238,N_28086,N_26885);
xor U34239 (N_34239,N_29049,N_25457);
nand U34240 (N_34240,N_26972,N_28310);
xor U34241 (N_34241,N_29744,N_27196);
nor U34242 (N_34242,N_25222,N_27985);
nor U34243 (N_34243,N_26176,N_29004);
or U34244 (N_34244,N_29042,N_25135);
nor U34245 (N_34245,N_28360,N_26621);
nand U34246 (N_34246,N_26601,N_26110);
xnor U34247 (N_34247,N_29398,N_27646);
xor U34248 (N_34248,N_27490,N_27487);
or U34249 (N_34249,N_25368,N_25561);
nor U34250 (N_34250,N_27039,N_25983);
and U34251 (N_34251,N_25664,N_26804);
nand U34252 (N_34252,N_27509,N_26931);
nor U34253 (N_34253,N_25524,N_25313);
and U34254 (N_34254,N_27330,N_27038);
nor U34255 (N_34255,N_27747,N_28861);
xor U34256 (N_34256,N_28452,N_26547);
and U34257 (N_34257,N_25985,N_26072);
nor U34258 (N_34258,N_25326,N_29023);
and U34259 (N_34259,N_29701,N_26018);
or U34260 (N_34260,N_27111,N_29946);
and U34261 (N_34261,N_29629,N_28020);
nor U34262 (N_34262,N_28317,N_27357);
or U34263 (N_34263,N_29816,N_25484);
nor U34264 (N_34264,N_29657,N_26034);
nand U34265 (N_34265,N_26199,N_28177);
nand U34266 (N_34266,N_29231,N_27349);
or U34267 (N_34267,N_28794,N_25015);
nand U34268 (N_34268,N_27387,N_25745);
nand U34269 (N_34269,N_27397,N_26705);
or U34270 (N_34270,N_26900,N_25730);
xnor U34271 (N_34271,N_28921,N_28918);
and U34272 (N_34272,N_29886,N_25884);
or U34273 (N_34273,N_28031,N_29406);
nand U34274 (N_34274,N_28385,N_27623);
nor U34275 (N_34275,N_25623,N_26765);
xor U34276 (N_34276,N_29416,N_26040);
or U34277 (N_34277,N_27468,N_26741);
nor U34278 (N_34278,N_25617,N_29381);
xnor U34279 (N_34279,N_28585,N_28159);
xnor U34280 (N_34280,N_28233,N_25236);
xor U34281 (N_34281,N_28326,N_29636);
and U34282 (N_34282,N_25650,N_26442);
xor U34283 (N_34283,N_28732,N_25377);
nand U34284 (N_34284,N_26475,N_25273);
nand U34285 (N_34285,N_26525,N_29984);
xnor U34286 (N_34286,N_25989,N_26263);
xor U34287 (N_34287,N_25598,N_26925);
or U34288 (N_34288,N_29682,N_27299);
or U34289 (N_34289,N_29559,N_29417);
xor U34290 (N_34290,N_27222,N_27705);
nor U34291 (N_34291,N_29255,N_29191);
or U34292 (N_34292,N_27070,N_25443);
nand U34293 (N_34293,N_29824,N_25208);
or U34294 (N_34294,N_26515,N_26330);
nand U34295 (N_34295,N_27699,N_25599);
nor U34296 (N_34296,N_25892,N_26741);
or U34297 (N_34297,N_29260,N_25322);
nand U34298 (N_34298,N_26883,N_25752);
xor U34299 (N_34299,N_29740,N_29250);
or U34300 (N_34300,N_29458,N_25960);
and U34301 (N_34301,N_25446,N_27799);
nor U34302 (N_34302,N_29863,N_26756);
xnor U34303 (N_34303,N_26619,N_28539);
nand U34304 (N_34304,N_29876,N_29272);
or U34305 (N_34305,N_29072,N_25762);
xnor U34306 (N_34306,N_25406,N_25019);
nor U34307 (N_34307,N_29452,N_27110);
xor U34308 (N_34308,N_27385,N_25550);
xnor U34309 (N_34309,N_25524,N_25375);
nand U34310 (N_34310,N_26711,N_26320);
and U34311 (N_34311,N_25760,N_25714);
nand U34312 (N_34312,N_27613,N_25322);
nor U34313 (N_34313,N_26122,N_27557);
xnor U34314 (N_34314,N_29975,N_29613);
nand U34315 (N_34315,N_27712,N_25027);
and U34316 (N_34316,N_27401,N_26073);
nand U34317 (N_34317,N_28158,N_29175);
and U34318 (N_34318,N_26481,N_26220);
or U34319 (N_34319,N_29131,N_26606);
or U34320 (N_34320,N_29207,N_28071);
xor U34321 (N_34321,N_29864,N_28909);
or U34322 (N_34322,N_27858,N_27793);
nand U34323 (N_34323,N_25745,N_28874);
nand U34324 (N_34324,N_28004,N_28512);
or U34325 (N_34325,N_25212,N_28186);
xnor U34326 (N_34326,N_27044,N_29829);
nor U34327 (N_34327,N_29507,N_27416);
nor U34328 (N_34328,N_27946,N_28436);
or U34329 (N_34329,N_26056,N_27723);
nor U34330 (N_34330,N_25516,N_25303);
xnor U34331 (N_34331,N_28739,N_29039);
or U34332 (N_34332,N_29548,N_26703);
nand U34333 (N_34333,N_26918,N_25586);
nand U34334 (N_34334,N_27981,N_27416);
and U34335 (N_34335,N_26854,N_28183);
nand U34336 (N_34336,N_28819,N_29262);
nor U34337 (N_34337,N_26681,N_29415);
and U34338 (N_34338,N_26863,N_27316);
nand U34339 (N_34339,N_26200,N_25099);
and U34340 (N_34340,N_29194,N_28684);
xnor U34341 (N_34341,N_29476,N_28770);
nor U34342 (N_34342,N_29400,N_26379);
nor U34343 (N_34343,N_29138,N_26606);
or U34344 (N_34344,N_28975,N_26766);
xnor U34345 (N_34345,N_28318,N_26972);
or U34346 (N_34346,N_29668,N_27102);
nand U34347 (N_34347,N_26183,N_28438);
nor U34348 (N_34348,N_29544,N_27122);
xnor U34349 (N_34349,N_25139,N_27044);
and U34350 (N_34350,N_25157,N_25381);
and U34351 (N_34351,N_26856,N_28608);
xnor U34352 (N_34352,N_25193,N_27789);
xnor U34353 (N_34353,N_25929,N_27518);
nand U34354 (N_34354,N_26128,N_26693);
nand U34355 (N_34355,N_28968,N_29546);
nand U34356 (N_34356,N_28436,N_25456);
and U34357 (N_34357,N_27458,N_29161);
nor U34358 (N_34358,N_28952,N_26995);
nand U34359 (N_34359,N_26177,N_29845);
xor U34360 (N_34360,N_27787,N_25072);
or U34361 (N_34361,N_27719,N_29722);
and U34362 (N_34362,N_29480,N_27380);
and U34363 (N_34363,N_28329,N_29507);
xor U34364 (N_34364,N_25249,N_25009);
and U34365 (N_34365,N_25826,N_29496);
or U34366 (N_34366,N_26790,N_26205);
and U34367 (N_34367,N_26326,N_28790);
nand U34368 (N_34368,N_25675,N_26023);
and U34369 (N_34369,N_29692,N_27268);
and U34370 (N_34370,N_29209,N_29247);
xor U34371 (N_34371,N_27095,N_28855);
and U34372 (N_34372,N_29547,N_29717);
nand U34373 (N_34373,N_25294,N_29306);
nand U34374 (N_34374,N_27289,N_26732);
nor U34375 (N_34375,N_25839,N_27957);
xnor U34376 (N_34376,N_26162,N_25820);
nand U34377 (N_34377,N_26414,N_27199);
xor U34378 (N_34378,N_26900,N_27054);
nor U34379 (N_34379,N_27258,N_25061);
nand U34380 (N_34380,N_28039,N_27205);
or U34381 (N_34381,N_26843,N_25994);
or U34382 (N_34382,N_29809,N_28086);
nand U34383 (N_34383,N_28487,N_27887);
nor U34384 (N_34384,N_25174,N_25826);
nand U34385 (N_34385,N_29008,N_25705);
nor U34386 (N_34386,N_29476,N_25651);
or U34387 (N_34387,N_25969,N_29864);
nor U34388 (N_34388,N_26383,N_27120);
nor U34389 (N_34389,N_25108,N_27749);
nand U34390 (N_34390,N_28258,N_25607);
xor U34391 (N_34391,N_28817,N_25120);
and U34392 (N_34392,N_27917,N_26106);
xor U34393 (N_34393,N_26865,N_27497);
xnor U34394 (N_34394,N_29673,N_25231);
nand U34395 (N_34395,N_26292,N_28092);
nor U34396 (N_34396,N_26942,N_29837);
or U34397 (N_34397,N_26121,N_28595);
xnor U34398 (N_34398,N_26536,N_28822);
nor U34399 (N_34399,N_29148,N_29975);
xor U34400 (N_34400,N_28266,N_25030);
nand U34401 (N_34401,N_27272,N_28088);
or U34402 (N_34402,N_28758,N_28379);
nand U34403 (N_34403,N_26072,N_27267);
and U34404 (N_34404,N_25219,N_29435);
or U34405 (N_34405,N_27875,N_29394);
nor U34406 (N_34406,N_28170,N_26660);
xnor U34407 (N_34407,N_27824,N_28460);
nor U34408 (N_34408,N_29210,N_26008);
xor U34409 (N_34409,N_29762,N_27699);
or U34410 (N_34410,N_25195,N_25264);
and U34411 (N_34411,N_25244,N_26531);
xor U34412 (N_34412,N_27730,N_27799);
nor U34413 (N_34413,N_28019,N_27692);
or U34414 (N_34414,N_29054,N_29737);
xnor U34415 (N_34415,N_27157,N_27057);
nand U34416 (N_34416,N_27822,N_28678);
nand U34417 (N_34417,N_29680,N_25991);
or U34418 (N_34418,N_26924,N_26696);
nand U34419 (N_34419,N_28824,N_26273);
and U34420 (N_34420,N_27219,N_28202);
xor U34421 (N_34421,N_28568,N_25432);
xnor U34422 (N_34422,N_28706,N_28951);
nand U34423 (N_34423,N_29457,N_25018);
nand U34424 (N_34424,N_26251,N_25950);
nor U34425 (N_34425,N_27286,N_29710);
nor U34426 (N_34426,N_26389,N_29094);
or U34427 (N_34427,N_26221,N_29644);
nand U34428 (N_34428,N_29688,N_25847);
nor U34429 (N_34429,N_28730,N_26779);
nand U34430 (N_34430,N_25230,N_28630);
or U34431 (N_34431,N_27810,N_25226);
or U34432 (N_34432,N_28960,N_27868);
and U34433 (N_34433,N_29807,N_26629);
nand U34434 (N_34434,N_25051,N_28311);
or U34435 (N_34435,N_26791,N_27769);
or U34436 (N_34436,N_26086,N_28161);
xnor U34437 (N_34437,N_25795,N_25212);
nor U34438 (N_34438,N_28058,N_26231);
nor U34439 (N_34439,N_26825,N_26180);
or U34440 (N_34440,N_28835,N_25099);
xnor U34441 (N_34441,N_27561,N_26505);
nand U34442 (N_34442,N_25962,N_26950);
and U34443 (N_34443,N_27991,N_25198);
xor U34444 (N_34444,N_26707,N_27806);
nor U34445 (N_34445,N_29922,N_26881);
nand U34446 (N_34446,N_28654,N_27521);
or U34447 (N_34447,N_26140,N_26114);
nor U34448 (N_34448,N_29721,N_25020);
or U34449 (N_34449,N_26245,N_25256);
and U34450 (N_34450,N_25860,N_26141);
nor U34451 (N_34451,N_26469,N_27520);
xor U34452 (N_34452,N_28650,N_27300);
and U34453 (N_34453,N_28471,N_27785);
nand U34454 (N_34454,N_29162,N_28917);
xnor U34455 (N_34455,N_29997,N_25277);
xnor U34456 (N_34456,N_26459,N_28439);
and U34457 (N_34457,N_28532,N_28665);
and U34458 (N_34458,N_25433,N_25211);
and U34459 (N_34459,N_29349,N_26688);
or U34460 (N_34460,N_27079,N_27447);
and U34461 (N_34461,N_28445,N_25151);
xor U34462 (N_34462,N_25539,N_27420);
and U34463 (N_34463,N_27216,N_27461);
and U34464 (N_34464,N_29128,N_25568);
nor U34465 (N_34465,N_29032,N_28715);
nand U34466 (N_34466,N_25697,N_28041);
nand U34467 (N_34467,N_27180,N_28636);
nor U34468 (N_34468,N_25776,N_27416);
or U34469 (N_34469,N_27676,N_26006);
xnor U34470 (N_34470,N_25527,N_26880);
and U34471 (N_34471,N_29879,N_25536);
nand U34472 (N_34472,N_26036,N_27095);
and U34473 (N_34473,N_28338,N_26705);
nand U34474 (N_34474,N_25785,N_27360);
and U34475 (N_34475,N_26477,N_26851);
or U34476 (N_34476,N_28899,N_27665);
nor U34477 (N_34477,N_27351,N_27749);
nand U34478 (N_34478,N_26579,N_29690);
nand U34479 (N_34479,N_29566,N_26122);
nor U34480 (N_34480,N_27552,N_29887);
or U34481 (N_34481,N_29279,N_29298);
and U34482 (N_34482,N_29762,N_25083);
nand U34483 (N_34483,N_25149,N_25231);
xnor U34484 (N_34484,N_28565,N_29944);
and U34485 (N_34485,N_29337,N_29839);
and U34486 (N_34486,N_27634,N_25696);
nand U34487 (N_34487,N_25248,N_28212);
nor U34488 (N_34488,N_29506,N_25397);
nand U34489 (N_34489,N_25542,N_27231);
nand U34490 (N_34490,N_28361,N_27719);
or U34491 (N_34491,N_26601,N_26661);
nor U34492 (N_34492,N_26697,N_25239);
xor U34493 (N_34493,N_26919,N_27046);
nand U34494 (N_34494,N_26394,N_29256);
and U34495 (N_34495,N_27335,N_29528);
and U34496 (N_34496,N_29202,N_27941);
and U34497 (N_34497,N_27523,N_27514);
or U34498 (N_34498,N_27213,N_28291);
nand U34499 (N_34499,N_26661,N_29376);
and U34500 (N_34500,N_29611,N_25490);
nor U34501 (N_34501,N_29043,N_29021);
nor U34502 (N_34502,N_29965,N_28925);
nand U34503 (N_34503,N_26744,N_29004);
or U34504 (N_34504,N_29846,N_26838);
or U34505 (N_34505,N_29675,N_27479);
nor U34506 (N_34506,N_25836,N_28302);
nor U34507 (N_34507,N_25785,N_26815);
nor U34508 (N_34508,N_25153,N_28864);
nor U34509 (N_34509,N_26760,N_29530);
xnor U34510 (N_34510,N_29238,N_28874);
nor U34511 (N_34511,N_26527,N_27052);
nand U34512 (N_34512,N_25389,N_28544);
nor U34513 (N_34513,N_29833,N_27759);
and U34514 (N_34514,N_29995,N_26682);
nor U34515 (N_34515,N_27817,N_25878);
or U34516 (N_34516,N_29124,N_26080);
and U34517 (N_34517,N_27124,N_29313);
or U34518 (N_34518,N_29684,N_27641);
xnor U34519 (N_34519,N_27562,N_29506);
or U34520 (N_34520,N_29733,N_26254);
nor U34521 (N_34521,N_25988,N_26506);
xor U34522 (N_34522,N_26991,N_27549);
or U34523 (N_34523,N_27276,N_26928);
nor U34524 (N_34524,N_27665,N_25578);
nand U34525 (N_34525,N_26678,N_28569);
xor U34526 (N_34526,N_26150,N_27999);
xor U34527 (N_34527,N_29349,N_27713);
nand U34528 (N_34528,N_29642,N_27600);
and U34529 (N_34529,N_26948,N_25083);
nand U34530 (N_34530,N_26130,N_29366);
nand U34531 (N_34531,N_29336,N_27358);
xor U34532 (N_34532,N_28241,N_25956);
or U34533 (N_34533,N_28575,N_27890);
nor U34534 (N_34534,N_29974,N_28990);
and U34535 (N_34535,N_27594,N_28369);
and U34536 (N_34536,N_27873,N_26927);
nor U34537 (N_34537,N_26849,N_27958);
nand U34538 (N_34538,N_26644,N_29779);
nor U34539 (N_34539,N_29786,N_29277);
nand U34540 (N_34540,N_28637,N_28824);
nand U34541 (N_34541,N_28640,N_26434);
xor U34542 (N_34542,N_28368,N_26449);
or U34543 (N_34543,N_27218,N_25250);
nor U34544 (N_34544,N_25731,N_28527);
nor U34545 (N_34545,N_29642,N_26270);
or U34546 (N_34546,N_29443,N_27926);
or U34547 (N_34547,N_29277,N_26754);
xnor U34548 (N_34548,N_29893,N_25176);
nand U34549 (N_34549,N_28417,N_27738);
and U34550 (N_34550,N_29852,N_25940);
or U34551 (N_34551,N_25323,N_25237);
xor U34552 (N_34552,N_29446,N_28380);
nor U34553 (N_34553,N_26148,N_28138);
or U34554 (N_34554,N_25491,N_27011);
nor U34555 (N_34555,N_25620,N_29764);
nand U34556 (N_34556,N_26115,N_27086);
and U34557 (N_34557,N_29551,N_25526);
and U34558 (N_34558,N_29192,N_25639);
nor U34559 (N_34559,N_27565,N_26869);
or U34560 (N_34560,N_29581,N_26327);
nand U34561 (N_34561,N_26011,N_26052);
nor U34562 (N_34562,N_29051,N_29744);
nor U34563 (N_34563,N_28482,N_26204);
nor U34564 (N_34564,N_27919,N_27052);
nand U34565 (N_34565,N_28778,N_26117);
and U34566 (N_34566,N_28805,N_25361);
and U34567 (N_34567,N_26544,N_28382);
or U34568 (N_34568,N_26481,N_29827);
nand U34569 (N_34569,N_25581,N_29647);
and U34570 (N_34570,N_28951,N_25378);
xnor U34571 (N_34571,N_29725,N_28564);
nand U34572 (N_34572,N_29715,N_25504);
and U34573 (N_34573,N_26478,N_28278);
and U34574 (N_34574,N_27346,N_29339);
xnor U34575 (N_34575,N_29989,N_27006);
or U34576 (N_34576,N_26686,N_26067);
or U34577 (N_34577,N_28585,N_29242);
or U34578 (N_34578,N_27783,N_29557);
and U34579 (N_34579,N_26045,N_29480);
and U34580 (N_34580,N_29678,N_25367);
xnor U34581 (N_34581,N_29678,N_27917);
nor U34582 (N_34582,N_25700,N_25801);
or U34583 (N_34583,N_28739,N_29072);
nand U34584 (N_34584,N_25908,N_28127);
xnor U34585 (N_34585,N_25615,N_27287);
nor U34586 (N_34586,N_28753,N_28383);
and U34587 (N_34587,N_26412,N_26317);
nor U34588 (N_34588,N_27686,N_26975);
nor U34589 (N_34589,N_27795,N_27288);
nand U34590 (N_34590,N_28908,N_28292);
and U34591 (N_34591,N_28035,N_25317);
or U34592 (N_34592,N_25594,N_28954);
nor U34593 (N_34593,N_25245,N_28140);
and U34594 (N_34594,N_29934,N_29929);
nor U34595 (N_34595,N_25819,N_25069);
or U34596 (N_34596,N_25000,N_25577);
xor U34597 (N_34597,N_27594,N_29563);
xnor U34598 (N_34598,N_28104,N_26417);
xor U34599 (N_34599,N_27746,N_29283);
nor U34600 (N_34600,N_28736,N_28384);
nand U34601 (N_34601,N_28397,N_25750);
or U34602 (N_34602,N_25034,N_26768);
nor U34603 (N_34603,N_25257,N_27563);
nor U34604 (N_34604,N_29947,N_27825);
and U34605 (N_34605,N_29628,N_29705);
and U34606 (N_34606,N_27274,N_28007);
or U34607 (N_34607,N_27805,N_27503);
xnor U34608 (N_34608,N_28418,N_29280);
or U34609 (N_34609,N_25441,N_29477);
or U34610 (N_34610,N_25440,N_29823);
nor U34611 (N_34611,N_28182,N_27723);
or U34612 (N_34612,N_25000,N_29351);
or U34613 (N_34613,N_26514,N_29282);
nand U34614 (N_34614,N_25217,N_26231);
xnor U34615 (N_34615,N_26537,N_28522);
nand U34616 (N_34616,N_29555,N_29281);
or U34617 (N_34617,N_29842,N_26152);
nor U34618 (N_34618,N_29263,N_26282);
and U34619 (N_34619,N_28778,N_25305);
or U34620 (N_34620,N_29529,N_28867);
and U34621 (N_34621,N_25748,N_28117);
xnor U34622 (N_34622,N_25006,N_28521);
nand U34623 (N_34623,N_27658,N_27796);
and U34624 (N_34624,N_29323,N_28461);
nand U34625 (N_34625,N_27988,N_26597);
nor U34626 (N_34626,N_26372,N_25424);
or U34627 (N_34627,N_27381,N_28070);
or U34628 (N_34628,N_25178,N_27148);
nand U34629 (N_34629,N_25735,N_26342);
nand U34630 (N_34630,N_29150,N_25579);
nand U34631 (N_34631,N_28513,N_28845);
xor U34632 (N_34632,N_27657,N_26040);
nor U34633 (N_34633,N_26014,N_29615);
or U34634 (N_34634,N_27471,N_28302);
xor U34635 (N_34635,N_29058,N_26259);
xnor U34636 (N_34636,N_26109,N_27162);
or U34637 (N_34637,N_29586,N_29830);
nand U34638 (N_34638,N_28711,N_27844);
nand U34639 (N_34639,N_27655,N_28668);
or U34640 (N_34640,N_29641,N_27754);
nand U34641 (N_34641,N_26637,N_29141);
xnor U34642 (N_34642,N_28760,N_27730);
xor U34643 (N_34643,N_27734,N_25923);
and U34644 (N_34644,N_25231,N_25625);
xor U34645 (N_34645,N_25002,N_27509);
and U34646 (N_34646,N_29417,N_29831);
nand U34647 (N_34647,N_26370,N_27105);
nand U34648 (N_34648,N_28959,N_28188);
nor U34649 (N_34649,N_27246,N_28754);
xnor U34650 (N_34650,N_29878,N_27851);
and U34651 (N_34651,N_27092,N_27061);
nor U34652 (N_34652,N_29051,N_26981);
or U34653 (N_34653,N_26745,N_25808);
and U34654 (N_34654,N_26426,N_25896);
xor U34655 (N_34655,N_27066,N_28767);
nor U34656 (N_34656,N_27719,N_27956);
and U34657 (N_34657,N_28678,N_25142);
and U34658 (N_34658,N_26392,N_29433);
and U34659 (N_34659,N_27104,N_26538);
and U34660 (N_34660,N_26843,N_26291);
or U34661 (N_34661,N_25142,N_29760);
nand U34662 (N_34662,N_25441,N_28513);
nor U34663 (N_34663,N_29275,N_29791);
and U34664 (N_34664,N_25592,N_26525);
nand U34665 (N_34665,N_28578,N_29427);
xor U34666 (N_34666,N_25971,N_26042);
nand U34667 (N_34667,N_25448,N_28814);
and U34668 (N_34668,N_25407,N_28615);
or U34669 (N_34669,N_26880,N_26999);
nand U34670 (N_34670,N_25646,N_25560);
or U34671 (N_34671,N_25629,N_28794);
or U34672 (N_34672,N_27143,N_26888);
and U34673 (N_34673,N_27311,N_28568);
and U34674 (N_34674,N_25868,N_27270);
xnor U34675 (N_34675,N_28886,N_25675);
and U34676 (N_34676,N_28972,N_26382);
and U34677 (N_34677,N_25287,N_28950);
nor U34678 (N_34678,N_27282,N_27678);
nor U34679 (N_34679,N_25467,N_27162);
and U34680 (N_34680,N_25541,N_25180);
or U34681 (N_34681,N_28439,N_25802);
or U34682 (N_34682,N_26207,N_28762);
or U34683 (N_34683,N_25172,N_28912);
and U34684 (N_34684,N_25719,N_28579);
nor U34685 (N_34685,N_26510,N_28170);
nor U34686 (N_34686,N_25977,N_29830);
and U34687 (N_34687,N_29754,N_29184);
nand U34688 (N_34688,N_28942,N_29229);
and U34689 (N_34689,N_26318,N_26479);
and U34690 (N_34690,N_26673,N_26787);
and U34691 (N_34691,N_27113,N_27685);
and U34692 (N_34692,N_28970,N_25309);
nand U34693 (N_34693,N_28071,N_26028);
nand U34694 (N_34694,N_27545,N_26495);
nor U34695 (N_34695,N_25102,N_27119);
and U34696 (N_34696,N_28368,N_28243);
or U34697 (N_34697,N_28633,N_29268);
nand U34698 (N_34698,N_29918,N_28691);
or U34699 (N_34699,N_26191,N_29329);
nor U34700 (N_34700,N_29777,N_27885);
nor U34701 (N_34701,N_29039,N_28119);
or U34702 (N_34702,N_27394,N_26308);
or U34703 (N_34703,N_27724,N_28999);
nand U34704 (N_34704,N_26177,N_25144);
nor U34705 (N_34705,N_27411,N_25613);
nor U34706 (N_34706,N_25523,N_27946);
and U34707 (N_34707,N_27978,N_26306);
nor U34708 (N_34708,N_27687,N_27466);
nand U34709 (N_34709,N_28813,N_29421);
and U34710 (N_34710,N_26885,N_26104);
and U34711 (N_34711,N_29839,N_27172);
xor U34712 (N_34712,N_27954,N_25000);
and U34713 (N_34713,N_26977,N_25870);
nor U34714 (N_34714,N_26383,N_28263);
and U34715 (N_34715,N_26906,N_26271);
and U34716 (N_34716,N_25865,N_29897);
xor U34717 (N_34717,N_25533,N_25965);
and U34718 (N_34718,N_29109,N_28930);
xnor U34719 (N_34719,N_29246,N_28432);
nor U34720 (N_34720,N_27642,N_28549);
and U34721 (N_34721,N_25217,N_26863);
nor U34722 (N_34722,N_27330,N_26305);
and U34723 (N_34723,N_29116,N_26120);
or U34724 (N_34724,N_25879,N_28170);
nor U34725 (N_34725,N_28230,N_28545);
nor U34726 (N_34726,N_26331,N_27484);
or U34727 (N_34727,N_27260,N_27890);
and U34728 (N_34728,N_26476,N_26751);
nor U34729 (N_34729,N_26888,N_27272);
or U34730 (N_34730,N_28009,N_25347);
xor U34731 (N_34731,N_26538,N_25620);
xor U34732 (N_34732,N_26843,N_27686);
nor U34733 (N_34733,N_28611,N_26612);
nor U34734 (N_34734,N_29262,N_27250);
xor U34735 (N_34735,N_29386,N_29696);
xnor U34736 (N_34736,N_26024,N_25603);
xnor U34737 (N_34737,N_26964,N_28969);
or U34738 (N_34738,N_27681,N_25564);
and U34739 (N_34739,N_29009,N_26064);
or U34740 (N_34740,N_25965,N_27748);
nor U34741 (N_34741,N_28356,N_27185);
nor U34742 (N_34742,N_25777,N_28897);
or U34743 (N_34743,N_28125,N_29005);
nand U34744 (N_34744,N_29241,N_28979);
or U34745 (N_34745,N_29938,N_26084);
or U34746 (N_34746,N_28658,N_28385);
or U34747 (N_34747,N_26177,N_26124);
nand U34748 (N_34748,N_27943,N_29148);
or U34749 (N_34749,N_26216,N_28775);
or U34750 (N_34750,N_26214,N_27581);
xor U34751 (N_34751,N_29192,N_29356);
and U34752 (N_34752,N_25903,N_28995);
nor U34753 (N_34753,N_29792,N_27300);
xor U34754 (N_34754,N_25196,N_26650);
xor U34755 (N_34755,N_29352,N_28811);
or U34756 (N_34756,N_28105,N_26531);
or U34757 (N_34757,N_26587,N_28022);
nor U34758 (N_34758,N_26493,N_29992);
or U34759 (N_34759,N_29052,N_29379);
nor U34760 (N_34760,N_28197,N_26280);
xor U34761 (N_34761,N_25792,N_26209);
nor U34762 (N_34762,N_29992,N_27689);
nor U34763 (N_34763,N_26701,N_27270);
and U34764 (N_34764,N_25992,N_29781);
nand U34765 (N_34765,N_25026,N_29274);
and U34766 (N_34766,N_29355,N_26026);
nand U34767 (N_34767,N_28721,N_25045);
nor U34768 (N_34768,N_28584,N_28217);
and U34769 (N_34769,N_29890,N_25967);
and U34770 (N_34770,N_25488,N_26667);
xnor U34771 (N_34771,N_29128,N_27198);
or U34772 (N_34772,N_25690,N_27192);
nor U34773 (N_34773,N_27993,N_27593);
nor U34774 (N_34774,N_26374,N_27281);
and U34775 (N_34775,N_28648,N_26712);
nand U34776 (N_34776,N_28872,N_26106);
and U34777 (N_34777,N_27536,N_26608);
xor U34778 (N_34778,N_25444,N_25074);
nor U34779 (N_34779,N_28450,N_27022);
or U34780 (N_34780,N_29370,N_25958);
and U34781 (N_34781,N_25232,N_25923);
and U34782 (N_34782,N_26937,N_29024);
nor U34783 (N_34783,N_27870,N_29731);
xnor U34784 (N_34784,N_29575,N_26783);
and U34785 (N_34785,N_29664,N_27870);
nand U34786 (N_34786,N_28145,N_25707);
xor U34787 (N_34787,N_29393,N_29681);
and U34788 (N_34788,N_29518,N_28745);
or U34789 (N_34789,N_26605,N_26520);
nor U34790 (N_34790,N_26528,N_25918);
and U34791 (N_34791,N_28944,N_25217);
or U34792 (N_34792,N_29746,N_29593);
and U34793 (N_34793,N_27529,N_28613);
or U34794 (N_34794,N_28561,N_27277);
and U34795 (N_34795,N_26370,N_27085);
and U34796 (N_34796,N_25256,N_29660);
nor U34797 (N_34797,N_28094,N_27574);
nand U34798 (N_34798,N_29273,N_26193);
nand U34799 (N_34799,N_27083,N_27368);
nand U34800 (N_34800,N_25634,N_25660);
or U34801 (N_34801,N_25542,N_27010);
nand U34802 (N_34802,N_26716,N_28959);
or U34803 (N_34803,N_29779,N_27008);
and U34804 (N_34804,N_29142,N_27998);
nand U34805 (N_34805,N_26648,N_29523);
and U34806 (N_34806,N_28831,N_28690);
or U34807 (N_34807,N_27063,N_29768);
xnor U34808 (N_34808,N_25625,N_25858);
xnor U34809 (N_34809,N_28923,N_26000);
nand U34810 (N_34810,N_26509,N_27405);
and U34811 (N_34811,N_27764,N_28600);
nor U34812 (N_34812,N_26082,N_26254);
or U34813 (N_34813,N_27220,N_29817);
xnor U34814 (N_34814,N_29856,N_27931);
nor U34815 (N_34815,N_25937,N_25564);
and U34816 (N_34816,N_27938,N_26811);
and U34817 (N_34817,N_27358,N_28238);
xor U34818 (N_34818,N_27958,N_25953);
xor U34819 (N_34819,N_27178,N_28499);
or U34820 (N_34820,N_25395,N_28489);
and U34821 (N_34821,N_25555,N_26215);
or U34822 (N_34822,N_26300,N_25625);
and U34823 (N_34823,N_28943,N_26449);
or U34824 (N_34824,N_26013,N_28219);
and U34825 (N_34825,N_26213,N_25804);
nor U34826 (N_34826,N_25755,N_26101);
nor U34827 (N_34827,N_28196,N_26156);
xor U34828 (N_34828,N_27389,N_29141);
nand U34829 (N_34829,N_29506,N_27648);
and U34830 (N_34830,N_28355,N_26447);
xnor U34831 (N_34831,N_29669,N_28328);
nor U34832 (N_34832,N_29211,N_27641);
and U34833 (N_34833,N_25414,N_28429);
or U34834 (N_34834,N_26592,N_25383);
nand U34835 (N_34835,N_27912,N_26283);
nand U34836 (N_34836,N_26700,N_29756);
and U34837 (N_34837,N_25857,N_28255);
nor U34838 (N_34838,N_29568,N_25366);
and U34839 (N_34839,N_26764,N_27351);
and U34840 (N_34840,N_27012,N_27892);
nor U34841 (N_34841,N_27269,N_27984);
xor U34842 (N_34842,N_29398,N_26773);
nand U34843 (N_34843,N_27327,N_26017);
or U34844 (N_34844,N_27676,N_25779);
or U34845 (N_34845,N_26692,N_28135);
nand U34846 (N_34846,N_26734,N_26748);
or U34847 (N_34847,N_27407,N_25473);
xor U34848 (N_34848,N_26840,N_25668);
and U34849 (N_34849,N_25324,N_28858);
xor U34850 (N_34850,N_25683,N_25105);
xor U34851 (N_34851,N_26285,N_27663);
and U34852 (N_34852,N_27163,N_28924);
or U34853 (N_34853,N_27131,N_27725);
or U34854 (N_34854,N_27658,N_28692);
nor U34855 (N_34855,N_26928,N_26783);
nor U34856 (N_34856,N_29922,N_25316);
or U34857 (N_34857,N_27908,N_29576);
and U34858 (N_34858,N_27103,N_29406);
and U34859 (N_34859,N_28635,N_26472);
nor U34860 (N_34860,N_27283,N_26018);
and U34861 (N_34861,N_26742,N_25602);
nand U34862 (N_34862,N_26890,N_25627);
xor U34863 (N_34863,N_27382,N_26075);
nor U34864 (N_34864,N_27488,N_27395);
nor U34865 (N_34865,N_26227,N_28119);
xor U34866 (N_34866,N_26345,N_26248);
and U34867 (N_34867,N_25048,N_26518);
nor U34868 (N_34868,N_27042,N_28054);
nor U34869 (N_34869,N_28390,N_29815);
nor U34870 (N_34870,N_26647,N_25546);
nand U34871 (N_34871,N_25901,N_29539);
nor U34872 (N_34872,N_26744,N_28675);
nand U34873 (N_34873,N_25752,N_28168);
or U34874 (N_34874,N_25701,N_25216);
or U34875 (N_34875,N_25209,N_26345);
nor U34876 (N_34876,N_27141,N_29699);
or U34877 (N_34877,N_25680,N_29752);
or U34878 (N_34878,N_29825,N_28613);
or U34879 (N_34879,N_29186,N_29942);
or U34880 (N_34880,N_27218,N_26133);
nand U34881 (N_34881,N_28093,N_27182);
xor U34882 (N_34882,N_26502,N_25120);
nand U34883 (N_34883,N_28273,N_25690);
nor U34884 (N_34884,N_26323,N_27187);
nand U34885 (N_34885,N_27315,N_27472);
and U34886 (N_34886,N_25912,N_25619);
or U34887 (N_34887,N_25946,N_27214);
or U34888 (N_34888,N_29415,N_26846);
nor U34889 (N_34889,N_25431,N_26811);
or U34890 (N_34890,N_27263,N_27262);
nor U34891 (N_34891,N_25358,N_26208);
xnor U34892 (N_34892,N_26410,N_26126);
nor U34893 (N_34893,N_25507,N_27721);
or U34894 (N_34894,N_29886,N_26247);
nor U34895 (N_34895,N_27516,N_25475);
nand U34896 (N_34896,N_27677,N_28766);
nand U34897 (N_34897,N_29520,N_29181);
and U34898 (N_34898,N_29828,N_27723);
nand U34899 (N_34899,N_29156,N_26072);
or U34900 (N_34900,N_27288,N_26762);
nor U34901 (N_34901,N_27008,N_28783);
nand U34902 (N_34902,N_29259,N_28178);
nand U34903 (N_34903,N_28520,N_29927);
nor U34904 (N_34904,N_25417,N_26324);
nor U34905 (N_34905,N_29080,N_27456);
or U34906 (N_34906,N_25655,N_27270);
or U34907 (N_34907,N_29833,N_26603);
xor U34908 (N_34908,N_26002,N_29955);
xor U34909 (N_34909,N_29424,N_25767);
xnor U34910 (N_34910,N_25389,N_25995);
or U34911 (N_34911,N_29663,N_28023);
and U34912 (N_34912,N_26371,N_28562);
or U34913 (N_34913,N_25194,N_26512);
xor U34914 (N_34914,N_29561,N_26705);
nor U34915 (N_34915,N_29616,N_29771);
nand U34916 (N_34916,N_29913,N_25729);
nor U34917 (N_34917,N_29632,N_27815);
nor U34918 (N_34918,N_27218,N_29802);
xor U34919 (N_34919,N_26126,N_27584);
or U34920 (N_34920,N_28255,N_29094);
and U34921 (N_34921,N_28872,N_29860);
nand U34922 (N_34922,N_27223,N_29642);
xnor U34923 (N_34923,N_27541,N_28994);
nor U34924 (N_34924,N_27747,N_25717);
and U34925 (N_34925,N_29887,N_28228);
nand U34926 (N_34926,N_25588,N_25067);
and U34927 (N_34927,N_26918,N_27160);
nor U34928 (N_34928,N_28922,N_25770);
or U34929 (N_34929,N_29862,N_25472);
nor U34930 (N_34930,N_28280,N_25625);
and U34931 (N_34931,N_29444,N_27733);
or U34932 (N_34932,N_29659,N_25023);
and U34933 (N_34933,N_25030,N_26555);
xor U34934 (N_34934,N_25901,N_28207);
and U34935 (N_34935,N_28729,N_29135);
or U34936 (N_34936,N_28052,N_28720);
nor U34937 (N_34937,N_27939,N_28245);
or U34938 (N_34938,N_28903,N_25099);
nand U34939 (N_34939,N_26954,N_26296);
and U34940 (N_34940,N_26728,N_27996);
xor U34941 (N_34941,N_26386,N_28695);
nor U34942 (N_34942,N_26849,N_28394);
nand U34943 (N_34943,N_27090,N_25681);
nor U34944 (N_34944,N_25992,N_25352);
or U34945 (N_34945,N_29975,N_29169);
nor U34946 (N_34946,N_28428,N_28261);
or U34947 (N_34947,N_28602,N_26256);
nand U34948 (N_34948,N_25011,N_25843);
nand U34949 (N_34949,N_25802,N_28174);
nor U34950 (N_34950,N_28821,N_27138);
or U34951 (N_34951,N_26757,N_29388);
and U34952 (N_34952,N_28073,N_27197);
nand U34953 (N_34953,N_25646,N_28528);
and U34954 (N_34954,N_27538,N_28266);
and U34955 (N_34955,N_27142,N_28365);
xor U34956 (N_34956,N_26313,N_25434);
xnor U34957 (N_34957,N_25316,N_28642);
or U34958 (N_34958,N_29967,N_25747);
xnor U34959 (N_34959,N_26034,N_26479);
nor U34960 (N_34960,N_29365,N_29363);
or U34961 (N_34961,N_26776,N_28327);
xnor U34962 (N_34962,N_29582,N_25854);
nor U34963 (N_34963,N_29484,N_26241);
nor U34964 (N_34964,N_27150,N_25015);
nand U34965 (N_34965,N_29673,N_27083);
xnor U34966 (N_34966,N_26438,N_27258);
nor U34967 (N_34967,N_25175,N_29100);
and U34968 (N_34968,N_28376,N_29824);
xnor U34969 (N_34969,N_29641,N_27476);
and U34970 (N_34970,N_26944,N_25969);
and U34971 (N_34971,N_25861,N_28994);
xor U34972 (N_34972,N_27273,N_27423);
nand U34973 (N_34973,N_25493,N_28339);
xor U34974 (N_34974,N_29576,N_25079);
nor U34975 (N_34975,N_27117,N_25329);
nand U34976 (N_34976,N_27599,N_25045);
and U34977 (N_34977,N_25314,N_28455);
xor U34978 (N_34978,N_26523,N_28867);
nand U34979 (N_34979,N_25580,N_29262);
nand U34980 (N_34980,N_26888,N_29712);
xnor U34981 (N_34981,N_27668,N_25987);
and U34982 (N_34982,N_26566,N_28652);
or U34983 (N_34983,N_27133,N_28401);
nand U34984 (N_34984,N_29728,N_26082);
xor U34985 (N_34985,N_27871,N_26812);
nor U34986 (N_34986,N_25909,N_26537);
and U34987 (N_34987,N_28040,N_28254);
nand U34988 (N_34988,N_28092,N_27910);
nand U34989 (N_34989,N_28799,N_28215);
or U34990 (N_34990,N_26317,N_25210);
xnor U34991 (N_34991,N_26895,N_28785);
nor U34992 (N_34992,N_29672,N_25556);
and U34993 (N_34993,N_29608,N_26862);
and U34994 (N_34994,N_25969,N_27455);
and U34995 (N_34995,N_28600,N_25485);
nand U34996 (N_34996,N_25245,N_27661);
nand U34997 (N_34997,N_26783,N_25675);
xor U34998 (N_34998,N_26479,N_29956);
or U34999 (N_34999,N_29434,N_25701);
nor U35000 (N_35000,N_32466,N_33767);
and U35001 (N_35001,N_33480,N_31194);
or U35002 (N_35002,N_34061,N_33169);
and U35003 (N_35003,N_32288,N_31259);
nor U35004 (N_35004,N_31813,N_30346);
nor U35005 (N_35005,N_34435,N_31827);
and U35006 (N_35006,N_33594,N_34875);
nor U35007 (N_35007,N_32457,N_33593);
nand U35008 (N_35008,N_30405,N_33402);
or U35009 (N_35009,N_31811,N_32300);
xnor U35010 (N_35010,N_34794,N_31446);
nor U35011 (N_35011,N_33483,N_34826);
or U35012 (N_35012,N_34947,N_31286);
nor U35013 (N_35013,N_31250,N_31274);
nand U35014 (N_35014,N_34820,N_30985);
nand U35015 (N_35015,N_33348,N_33874);
nor U35016 (N_35016,N_31472,N_32456);
nand U35017 (N_35017,N_31884,N_34733);
xnor U35018 (N_35018,N_34949,N_34987);
and U35019 (N_35019,N_32929,N_32625);
xor U35020 (N_35020,N_30158,N_34000);
xnor U35021 (N_35021,N_33681,N_31262);
xnor U35022 (N_35022,N_31842,N_31637);
and U35023 (N_35023,N_32594,N_30299);
nand U35024 (N_35024,N_31909,N_33698);
or U35025 (N_35025,N_31414,N_33140);
xor U35026 (N_35026,N_31658,N_30545);
or U35027 (N_35027,N_32276,N_30017);
and U35028 (N_35028,N_32634,N_30982);
or U35029 (N_35029,N_34264,N_34339);
xnor U35030 (N_35030,N_32937,N_33410);
nand U35031 (N_35031,N_32818,N_33122);
and U35032 (N_35032,N_32319,N_30209);
nor U35033 (N_35033,N_30398,N_30802);
xnor U35034 (N_35034,N_34953,N_30778);
or U35035 (N_35035,N_31569,N_31801);
or U35036 (N_35036,N_31240,N_32562);
nand U35037 (N_35037,N_33512,N_33964);
nor U35038 (N_35038,N_34661,N_30311);
or U35039 (N_35039,N_34031,N_32337);
nand U35040 (N_35040,N_30320,N_32142);
xnor U35041 (N_35041,N_33761,N_33923);
nand U35042 (N_35042,N_31885,N_31871);
nor U35043 (N_35043,N_34167,N_34812);
nor U35044 (N_35044,N_32870,N_31398);
nand U35045 (N_35045,N_30335,N_31341);
or U35046 (N_35046,N_33296,N_33183);
nand U35047 (N_35047,N_31180,N_30461);
and U35048 (N_35048,N_33050,N_31897);
nand U35049 (N_35049,N_30304,N_32563);
and U35050 (N_35050,N_31055,N_32965);
and U35051 (N_35051,N_30929,N_34180);
or U35052 (N_35052,N_30309,N_33824);
nand U35053 (N_35053,N_30554,N_31843);
nor U35054 (N_35054,N_30983,N_33559);
xnor U35055 (N_35055,N_32931,N_32406);
nand U35056 (N_35056,N_34950,N_30087);
nor U35057 (N_35057,N_34507,N_32785);
xor U35058 (N_35058,N_34508,N_32877);
nor U35059 (N_35059,N_30762,N_32536);
or U35060 (N_35060,N_34293,N_31866);
or U35061 (N_35061,N_34727,N_30737);
xnor U35062 (N_35062,N_34725,N_30996);
or U35063 (N_35063,N_34647,N_34536);
xnor U35064 (N_35064,N_31605,N_32051);
or U35065 (N_35065,N_31289,N_32685);
or U35066 (N_35066,N_32942,N_30914);
xnor U35067 (N_35067,N_31874,N_34576);
nor U35068 (N_35068,N_31880,N_30843);
xnor U35069 (N_35069,N_31382,N_30500);
or U35070 (N_35070,N_34432,N_34194);
and U35071 (N_35071,N_30485,N_31851);
xnor U35072 (N_35072,N_30056,N_31731);
nor U35073 (N_35073,N_34497,N_31601);
or U35074 (N_35074,N_33668,N_31548);
or U35075 (N_35075,N_34430,N_33872);
or U35076 (N_35076,N_33821,N_30849);
nand U35077 (N_35077,N_32910,N_31780);
or U35078 (N_35078,N_32390,N_31782);
nor U35079 (N_35079,N_32986,N_31957);
nor U35080 (N_35080,N_33830,N_33044);
or U35081 (N_35081,N_32404,N_31052);
or U35082 (N_35082,N_32556,N_33574);
nand U35083 (N_35083,N_34053,N_33445);
and U35084 (N_35084,N_30960,N_33401);
and U35085 (N_35085,N_34713,N_33525);
nand U35086 (N_35086,N_34801,N_33469);
nor U35087 (N_35087,N_32753,N_30492);
nand U35088 (N_35088,N_34858,N_31197);
and U35089 (N_35089,N_30907,N_33712);
nand U35090 (N_35090,N_31012,N_34496);
and U35091 (N_35091,N_33591,N_33231);
xnor U35092 (N_35092,N_33474,N_34296);
nand U35093 (N_35093,N_34521,N_32181);
or U35094 (N_35094,N_31890,N_34433);
xor U35095 (N_35095,N_30959,N_30466);
or U35096 (N_35096,N_31256,N_32991);
or U35097 (N_35097,N_33446,N_34933);
xnor U35098 (N_35098,N_30555,N_33714);
and U35099 (N_35099,N_34093,N_32282);
xnor U35100 (N_35100,N_31931,N_32869);
or U35101 (N_35101,N_30343,N_30046);
nand U35102 (N_35102,N_33451,N_31374);
nand U35103 (N_35103,N_32430,N_32540);
and U35104 (N_35104,N_34232,N_30387);
xor U35105 (N_35105,N_34193,N_34027);
nand U35106 (N_35106,N_31253,N_32264);
and U35107 (N_35107,N_31936,N_30260);
or U35108 (N_35108,N_34550,N_34625);
nor U35109 (N_35109,N_30697,N_33031);
nand U35110 (N_35110,N_34443,N_34611);
or U35111 (N_35111,N_32180,N_33277);
nor U35112 (N_35112,N_33543,N_32628);
nor U35113 (N_35113,N_32972,N_33170);
nand U35114 (N_35114,N_30129,N_30610);
and U35115 (N_35115,N_34566,N_34864);
xor U35116 (N_35116,N_33126,N_30036);
nand U35117 (N_35117,N_33364,N_34237);
nand U35118 (N_35118,N_33936,N_32314);
xnor U35119 (N_35119,N_30077,N_32672);
or U35120 (N_35120,N_31429,N_33938);
and U35121 (N_35121,N_30360,N_33240);
and U35122 (N_35122,N_33785,N_34278);
and U35123 (N_35123,N_33705,N_32623);
nand U35124 (N_35124,N_30862,N_30073);
or U35125 (N_35125,N_31376,N_33590);
xor U35126 (N_35126,N_32567,N_33511);
nor U35127 (N_35127,N_31610,N_30986);
nor U35128 (N_35128,N_32673,N_30663);
or U35129 (N_35129,N_32487,N_32218);
nor U35130 (N_35130,N_30266,N_30037);
nor U35131 (N_35131,N_33003,N_31997);
nor U35132 (N_35132,N_33455,N_32291);
and U35133 (N_35133,N_30772,N_33492);
xor U35134 (N_35134,N_31734,N_32982);
and U35135 (N_35135,N_32738,N_31744);
nand U35136 (N_35136,N_30112,N_34347);
nor U35137 (N_35137,N_30720,N_31098);
xnor U35138 (N_35138,N_33314,N_30809);
nor U35139 (N_35139,N_30845,N_30686);
nor U35140 (N_35140,N_32599,N_34104);
nor U35141 (N_35141,N_33301,N_32071);
nand U35142 (N_35142,N_31748,N_32401);
or U35143 (N_35143,N_32909,N_32076);
or U35144 (N_35144,N_33459,N_33981);
xnor U35145 (N_35145,N_32241,N_34262);
xnor U35146 (N_35146,N_34301,N_32546);
xnor U35147 (N_35147,N_30374,N_32043);
and U35148 (N_35148,N_33198,N_33907);
nand U35149 (N_35149,N_34250,N_32897);
nand U35150 (N_35150,N_33279,N_34165);
nor U35151 (N_35151,N_33333,N_32676);
nor U35152 (N_35152,N_30789,N_34852);
nand U35153 (N_35153,N_31457,N_32526);
and U35154 (N_35154,N_33566,N_34900);
and U35155 (N_35155,N_32169,N_31802);
or U35156 (N_35156,N_34276,N_33935);
nand U35157 (N_35157,N_33069,N_33613);
nand U35158 (N_35158,N_30392,N_31205);
nor U35159 (N_35159,N_30863,N_33097);
nand U35160 (N_35160,N_32829,N_30828);
and U35161 (N_35161,N_32185,N_32094);
nor U35162 (N_35162,N_32863,N_32453);
nand U35163 (N_35163,N_30113,N_31657);
nor U35164 (N_35164,N_32032,N_34789);
xnor U35165 (N_35165,N_31303,N_30380);
nand U35166 (N_35166,N_32149,N_32771);
nand U35167 (N_35167,N_30652,N_33804);
nor U35168 (N_35168,N_33866,N_32615);
xor U35169 (N_35169,N_34998,N_32883);
or U35170 (N_35170,N_31302,N_30830);
nand U35171 (N_35171,N_33528,N_34499);
nand U35172 (N_35172,N_31327,N_32465);
nand U35173 (N_35173,N_31943,N_34537);
xnor U35174 (N_35174,N_31774,N_30117);
xor U35175 (N_35175,N_34174,N_32956);
nor U35176 (N_35176,N_33639,N_32092);
nand U35177 (N_35177,N_32055,N_34094);
xnor U35178 (N_35178,N_31638,N_34436);
nor U35179 (N_35179,N_30462,N_34468);
nand U35180 (N_35180,N_31769,N_34086);
nand U35181 (N_35181,N_31178,N_30124);
and U35182 (N_35182,N_34962,N_34838);
nor U35183 (N_35183,N_31057,N_32793);
and U35184 (N_35184,N_30055,N_32788);
and U35185 (N_35185,N_30518,N_30451);
or U35186 (N_35186,N_32955,N_34187);
xnor U35187 (N_35187,N_32195,N_31913);
nand U35188 (N_35188,N_33690,N_33220);
and U35189 (N_35189,N_31311,N_32919);
and U35190 (N_35190,N_34960,N_34686);
or U35191 (N_35191,N_31528,N_30578);
nor U35192 (N_35192,N_34522,N_30991);
or U35193 (N_35193,N_33181,N_32507);
nor U35194 (N_35194,N_32297,N_32932);
nand U35195 (N_35195,N_30370,N_31070);
nor U35196 (N_35196,N_32455,N_33020);
and U35197 (N_35197,N_34901,N_33890);
xnor U35198 (N_35198,N_34955,N_30365);
nand U35199 (N_35199,N_31187,N_32443);
nor U35200 (N_35200,N_30390,N_33141);
xnor U35201 (N_35201,N_33107,N_33948);
or U35202 (N_35202,N_32702,N_33950);
nand U35203 (N_35203,N_31476,N_30875);
nand U35204 (N_35204,N_30742,N_30459);
or U35205 (N_35205,N_30665,N_34216);
or U35206 (N_35206,N_30759,N_30488);
and U35207 (N_35207,N_32005,N_30101);
xnor U35208 (N_35208,N_32777,N_32378);
and U35209 (N_35209,N_32516,N_32895);
and U35210 (N_35210,N_33070,N_33431);
nand U35211 (N_35211,N_31221,N_33222);
nand U35212 (N_35212,N_33243,N_33699);
or U35213 (N_35213,N_34695,N_32022);
xnor U35214 (N_35214,N_33408,N_32235);
xor U35215 (N_35215,N_32093,N_30035);
xor U35216 (N_35216,N_33532,N_30989);
and U35217 (N_35217,N_31225,N_34416);
and U35218 (N_35218,N_34684,N_33498);
nand U35219 (N_35219,N_34289,N_33683);
or U35220 (N_35220,N_33206,N_31437);
or U35221 (N_35221,N_30972,N_30600);
and U35222 (N_35222,N_32060,N_31352);
nor U35223 (N_35223,N_34030,N_32530);
xnor U35224 (N_35224,N_33368,N_30886);
nand U35225 (N_35225,N_30711,N_31881);
and U35226 (N_35226,N_30619,N_33148);
or U35227 (N_35227,N_34361,N_34452);
nor U35228 (N_35228,N_30753,N_33667);
nor U35229 (N_35229,N_30322,N_32402);
or U35230 (N_35230,N_30700,N_30074);
xor U35231 (N_35231,N_32136,N_34850);
and U35232 (N_35232,N_33197,N_31358);
and U35233 (N_35233,N_33823,N_33766);
or U35234 (N_35234,N_30840,N_30199);
nand U35235 (N_35235,N_32423,N_34798);
nand U35236 (N_35236,N_34085,N_33839);
and U35237 (N_35237,N_32807,N_32340);
xor U35238 (N_35238,N_33173,N_33079);
or U35239 (N_35239,N_34772,N_34151);
or U35240 (N_35240,N_31726,N_32460);
nor U35241 (N_35241,N_34996,N_34195);
xnor U35242 (N_35242,N_33743,N_31073);
or U35243 (N_35243,N_34631,N_30999);
nand U35244 (N_35244,N_33005,N_32105);
nand U35245 (N_35245,N_30443,N_33618);
xnor U35246 (N_35246,N_31222,N_30230);
nand U35247 (N_35247,N_32439,N_31993);
nand U35248 (N_35248,N_30970,N_32368);
nor U35249 (N_35249,N_30687,N_34786);
xnor U35250 (N_35250,N_34424,N_30321);
and U35251 (N_35251,N_30237,N_32718);
or U35252 (N_35252,N_33774,N_34136);
xnor U35253 (N_35253,N_33125,N_30942);
nor U35254 (N_35254,N_32379,N_33340);
nor U35255 (N_35255,N_34905,N_30958);
xor U35256 (N_35256,N_30897,N_31952);
nand U35257 (N_35257,N_31017,N_33685);
xnor U35258 (N_35258,N_33925,N_32486);
or U35259 (N_35259,N_34848,N_33893);
nor U35260 (N_35260,N_33619,N_30210);
nand U35261 (N_35261,N_30010,N_31338);
or U35262 (N_35262,N_30783,N_33799);
or U35263 (N_35263,N_34716,N_31718);
nand U35264 (N_35264,N_31093,N_33916);
and U35265 (N_35265,N_33624,N_31316);
nand U35266 (N_35266,N_30272,N_34284);
xnor U35267 (N_35267,N_30526,N_34616);
xnor U35268 (N_35268,N_31410,N_32707);
or U35269 (N_35269,N_30632,N_30564);
and U35270 (N_35270,N_30421,N_33553);
nor U35271 (N_35271,N_31166,N_31666);
or U35272 (N_35272,N_33878,N_34087);
or U35273 (N_35273,N_31103,N_33424);
xor U35274 (N_35274,N_34454,N_34314);
nor U35275 (N_35275,N_33167,N_30096);
and U35276 (N_35276,N_32867,N_30011);
or U35277 (N_35277,N_33385,N_34170);
and U35278 (N_35278,N_32520,N_33837);
nor U35279 (N_35279,N_30706,N_32735);
nor U35280 (N_35280,N_30995,N_30726);
xor U35281 (N_35281,N_32966,N_33349);
and U35282 (N_35282,N_33626,N_32153);
nor U35283 (N_35283,N_31284,N_32251);
xnor U35284 (N_35284,N_30801,N_34704);
or U35285 (N_35285,N_34349,N_33282);
nand U35286 (N_35286,N_33342,N_32096);
xnor U35287 (N_35287,N_30330,N_31521);
nor U35288 (N_35288,N_32429,N_31143);
xnor U35289 (N_35289,N_31413,N_33165);
nor U35290 (N_35290,N_33276,N_34045);
or U35291 (N_35291,N_32392,N_32683);
nand U35292 (N_35292,N_30356,N_32736);
nor U35293 (N_35293,N_31160,N_31270);
nand U35294 (N_35294,N_34326,N_32138);
nand U35295 (N_35295,N_34805,N_34006);
nor U35296 (N_35296,N_31593,N_30883);
xnor U35297 (N_35297,N_33249,N_30698);
nand U35298 (N_35298,N_31405,N_31743);
or U35299 (N_35299,N_34570,N_34883);
and U35300 (N_35300,N_34897,N_30009);
and U35301 (N_35301,N_34379,N_30739);
or U35302 (N_35302,N_30105,N_33978);
or U35303 (N_35303,N_31814,N_31014);
xnor U35304 (N_35304,N_30550,N_32916);
xnor U35305 (N_35305,N_31648,N_31242);
nand U35306 (N_35306,N_34816,N_34234);
and U35307 (N_35307,N_34723,N_32287);
nand U35308 (N_35308,N_31434,N_33735);
nor U35309 (N_35309,N_33632,N_33177);
and U35310 (N_35310,N_34032,N_33047);
xor U35311 (N_35311,N_34985,N_33739);
nor U35312 (N_35312,N_30206,N_33175);
nand U35313 (N_35313,N_30859,N_30505);
or U35314 (N_35314,N_33753,N_31389);
nand U35315 (N_35315,N_32791,N_30641);
and U35316 (N_35316,N_32190,N_30524);
nor U35317 (N_35317,N_33099,N_34580);
xor U35318 (N_35318,N_30864,N_34881);
nand U35319 (N_35319,N_34307,N_33980);
or U35320 (N_35320,N_31497,N_32508);
and U35321 (N_35321,N_31035,N_31927);
nand U35322 (N_35322,N_32728,N_34068);
nand U35323 (N_35323,N_30024,N_32559);
nand U35324 (N_35324,N_32593,N_34345);
and U35325 (N_35325,N_31230,N_33136);
nor U35326 (N_35326,N_31182,N_33355);
xor U35327 (N_35327,N_33992,N_32754);
or U35328 (N_35328,N_30172,N_33610);
or U35329 (N_35329,N_32463,N_34658);
or U35330 (N_35330,N_30342,N_30084);
and U35331 (N_35331,N_33537,N_33219);
nor U35332 (N_35332,N_32209,N_30803);
and U35333 (N_35333,N_33157,N_31611);
or U35334 (N_35334,N_30140,N_34303);
nand U35335 (N_35335,N_30973,N_32321);
nand U35336 (N_35336,N_32981,N_34977);
nor U35337 (N_35337,N_32131,N_31531);
nand U35338 (N_35338,N_30558,N_33363);
xnor U35339 (N_35339,N_34198,N_32686);
nand U35340 (N_35340,N_34783,N_34331);
or U35341 (N_35341,N_30850,N_32211);
and U35342 (N_35342,N_30193,N_34354);
xor U35343 (N_35343,N_31381,N_32970);
or U35344 (N_35344,N_32663,N_33952);
xor U35345 (N_35345,N_31454,N_32998);
xor U35346 (N_35346,N_32246,N_31479);
nand U35347 (N_35347,N_32033,N_34976);
and U35348 (N_35348,N_33150,N_30549);
xnor U35349 (N_35349,N_33317,N_30598);
nor U35350 (N_35350,N_31527,N_31096);
nor U35351 (N_35351,N_32997,N_31120);
nand U35352 (N_35352,N_34229,N_32644);
and U35353 (N_35353,N_30039,N_33650);
and U35354 (N_35354,N_33841,N_30487);
or U35355 (N_35355,N_30576,N_33082);
and U35356 (N_35356,N_32146,N_34777);
nor U35357 (N_35357,N_34890,N_32284);
and U35358 (N_35358,N_32589,N_34012);
xor U35359 (N_35359,N_32480,N_30650);
xor U35360 (N_35360,N_32098,N_30810);
or U35361 (N_35361,N_32611,N_32317);
nand U35362 (N_35362,N_31043,N_33765);
or U35363 (N_35363,N_30441,N_34598);
or U35364 (N_35364,N_34075,N_33749);
or U35365 (N_35365,N_31373,N_32498);
nor U35366 (N_35366,N_33625,N_32476);
and U35367 (N_35367,N_33404,N_32256);
and U35368 (N_35368,N_32274,N_31272);
nor U35369 (N_35369,N_30302,N_33724);
nand U35370 (N_35370,N_34313,N_33061);
nor U35371 (N_35371,N_34449,N_30314);
or U35372 (N_35372,N_33315,N_33702);
or U35373 (N_35373,N_31757,N_32884);
nand U35374 (N_35374,N_33731,N_34098);
or U35375 (N_35375,N_33584,N_34302);
xnor U35376 (N_35376,N_32836,N_31183);
nor U35377 (N_35377,N_30643,N_33054);
nand U35378 (N_35378,N_34830,N_32003);
nor U35379 (N_35379,N_32565,N_34503);
and U35380 (N_35380,N_30258,N_34400);
nand U35381 (N_35381,N_31059,N_31932);
nand U35382 (N_35382,N_34226,N_31815);
nand U35383 (N_35383,N_33991,N_32677);
or U35384 (N_35384,N_31714,N_32386);
or U35385 (N_35385,N_33599,N_30041);
xnor U35386 (N_35386,N_31760,N_33635);
xor U35387 (N_35387,N_34135,N_31649);
and U35388 (N_35388,N_33782,N_31618);
xor U35389 (N_35389,N_30766,N_33119);
or U35390 (N_35390,N_31267,N_33558);
nand U35391 (N_35391,N_32776,N_32061);
xnor U35392 (N_35392,N_32252,N_33787);
xnor U35393 (N_35393,N_31904,N_32550);
or U35394 (N_35394,N_31204,N_30291);
nor U35395 (N_35395,N_31124,N_30214);
xor U35396 (N_35396,N_31032,N_32715);
nor U35397 (N_35397,N_32268,N_31525);
xnor U35398 (N_35398,N_32583,N_31329);
xnor U35399 (N_35399,N_30563,N_33853);
xnor U35400 (N_35400,N_30635,N_33772);
or U35401 (N_35401,N_30949,N_31717);
nand U35402 (N_35402,N_31285,N_34177);
or U35403 (N_35403,N_34272,N_34806);
and U35404 (N_35404,N_33746,N_33059);
xor U35405 (N_35405,N_34362,N_34802);
nand U35406 (N_35406,N_34385,N_30372);
nor U35407 (N_35407,N_31268,N_33216);
and U35408 (N_35408,N_31438,N_32270);
and U35409 (N_35409,N_30428,N_33186);
nor U35410 (N_35410,N_31603,N_31509);
nand U35411 (N_35411,N_32204,N_33611);
and U35412 (N_35412,N_34002,N_34809);
and U35413 (N_35413,N_32109,N_33678);
and U35414 (N_35414,N_31218,N_31732);
xnor U35415 (N_35415,N_30175,N_32855);
xnor U35416 (N_35416,N_31620,N_34779);
and U35417 (N_35417,N_31107,N_34708);
or U35418 (N_35418,N_30718,N_33638);
xor U35419 (N_35419,N_31201,N_32619);
nor U35420 (N_35420,N_31536,N_33770);
nor U35421 (N_35421,N_31962,N_33018);
nor U35422 (N_35422,N_32134,N_30267);
xnor U35423 (N_35423,N_34642,N_31106);
or U35424 (N_35424,N_31226,N_33211);
and U35425 (N_35425,N_33760,N_32202);
nor U35426 (N_35426,N_33101,N_33922);
or U35427 (N_35427,N_32706,N_31979);
and U35428 (N_35428,N_31565,N_33997);
or U35429 (N_35429,N_31712,N_34102);
xnor U35430 (N_35430,N_31841,N_30353);
and U35431 (N_35431,N_32091,N_31005);
nand U35432 (N_35432,N_34069,N_30283);
nor U35433 (N_35433,N_34399,N_30556);
xor U35434 (N_35434,N_32364,N_31778);
nor U35435 (N_35435,N_33008,N_33245);
xnor U35436 (N_35436,N_33608,N_33264);
nand U35437 (N_35437,N_33396,N_33727);
or U35438 (N_35438,N_34144,N_31383);
or U35439 (N_35439,N_31305,N_31199);
or U35440 (N_35440,N_34579,N_33442);
nand U35441 (N_35441,N_30676,N_30426);
nand U35442 (N_35442,N_32737,N_32415);
xor U35443 (N_35443,N_31704,N_34747);
nand U35444 (N_35444,N_33075,N_34185);
and U35445 (N_35445,N_30577,N_34956);
or U35446 (N_35446,N_30484,N_31858);
xnor U35447 (N_35447,N_31144,N_33795);
xnor U35448 (N_35448,N_30820,N_31313);
nor U35449 (N_35449,N_32219,N_33603);
or U35450 (N_35450,N_32482,N_33247);
or U35451 (N_35451,N_30068,N_30834);
xnor U35452 (N_35452,N_32543,N_31860);
nor U35453 (N_35453,N_31336,N_31956);
and U35454 (N_35454,N_30953,N_31707);
nand U35455 (N_35455,N_30086,N_33902);
xor U35456 (N_35456,N_34348,N_33049);
nand U35457 (N_35457,N_32713,N_34523);
xnor U35458 (N_35458,N_30660,N_32835);
or U35459 (N_35459,N_34231,N_34267);
and U35460 (N_35460,N_34969,N_32808);
or U35461 (N_35461,N_32842,N_32127);
or U35462 (N_35462,N_34610,N_33897);
nand U35463 (N_35463,N_30666,N_34533);
nor U35464 (N_35464,N_34613,N_33343);
or U35465 (N_35465,N_34271,N_32744);
or U35466 (N_35466,N_31485,N_30190);
nor U35467 (N_35467,N_34358,N_32188);
and U35468 (N_35468,N_33002,N_34567);
or U35469 (N_35469,N_32393,N_33291);
or U35470 (N_35470,N_30174,N_32385);
xnor U35471 (N_35471,N_34089,N_33856);
nor U35472 (N_35472,N_31703,N_32339);
nand U35473 (N_35473,N_30444,N_33425);
nand U35474 (N_35474,N_30918,N_32865);
nand U35475 (N_35475,N_33213,N_34336);
nand U35476 (N_35476,N_33094,N_31715);
xor U35477 (N_35477,N_34082,N_34917);
nor U35478 (N_35478,N_33820,N_30509);
xnor U35479 (N_35479,N_33693,N_33691);
and U35480 (N_35480,N_31447,N_30453);
nor U35481 (N_35481,N_34861,N_30623);
xnor U35482 (N_35482,N_34070,N_30054);
xnor U35483 (N_35483,N_33858,N_34126);
or U35484 (N_35484,N_31384,N_32560);
and U35485 (N_35485,N_34880,N_34831);
nand U35486 (N_35486,N_34510,N_33899);
nand U35487 (N_35487,N_32362,N_34311);
xor U35488 (N_35488,N_32436,N_34448);
and U35489 (N_35489,N_30701,N_30908);
nor U35490 (N_35490,N_34051,N_32613);
xor U35491 (N_35491,N_30798,N_30498);
nor U35492 (N_35492,N_33665,N_34207);
nor U35493 (N_35493,N_33748,N_32627);
and U35494 (N_35494,N_33529,N_30228);
or U35495 (N_35495,N_30042,N_32356);
or U35496 (N_35496,N_32758,N_34846);
or U35497 (N_35497,N_30135,N_34241);
and U35498 (N_35498,N_31261,N_30255);
or U35499 (N_35499,N_34124,N_34186);
nor U35500 (N_35500,N_30780,N_34494);
or U35501 (N_35501,N_32725,N_32585);
xnor U35502 (N_35502,N_31089,N_33230);
nand U35503 (N_35503,N_32234,N_33623);
and U35504 (N_35504,N_34819,N_33473);
or U35505 (N_35505,N_32196,N_33738);
xnor U35506 (N_35506,N_33697,N_30544);
nor U35507 (N_35507,N_31248,N_33571);
or U35508 (N_35508,N_34142,N_33888);
and U35509 (N_35509,N_33456,N_32572);
nand U35510 (N_35510,N_34367,N_32154);
and U35511 (N_35511,N_33214,N_34722);
or U35512 (N_35512,N_34991,N_34254);
or U35513 (N_35513,N_33413,N_33440);
xor U35514 (N_35514,N_33199,N_30842);
xnor U35515 (N_35515,N_30889,N_31754);
or U35516 (N_35516,N_30489,N_32524);
nand U35517 (N_35517,N_30419,N_30574);
nand U35518 (N_35518,N_31898,N_33640);
nor U35519 (N_35519,N_30276,N_30377);
xor U35520 (N_35520,N_34659,N_32165);
or U35521 (N_35521,N_31489,N_31543);
or U35522 (N_35522,N_30692,N_34935);
and U35523 (N_35523,N_31153,N_30784);
xor U35524 (N_35524,N_31809,N_30002);
or U35525 (N_35525,N_31797,N_32857);
and U35526 (N_35526,N_33615,N_33526);
nor U35527 (N_35527,N_30601,N_34190);
and U35528 (N_35528,N_33283,N_30250);
nor U35529 (N_35529,N_34355,N_33100);
nand U35530 (N_35530,N_32355,N_33269);
nor U35531 (N_35531,N_32924,N_32258);
or U35532 (N_35532,N_31464,N_31679);
or U35533 (N_35533,N_31944,N_33388);
xor U35534 (N_35534,N_34461,N_31938);
or U35535 (N_35535,N_31783,N_30814);
nand U35536 (N_35536,N_34277,N_30779);
and U35537 (N_35537,N_34426,N_34431);
and U35538 (N_35538,N_33994,N_32509);
nor U35539 (N_35539,N_33205,N_31507);
nand U35540 (N_35540,N_32506,N_34615);
xnor U35541 (N_35541,N_32069,N_31319);
nor U35542 (N_35542,N_31886,N_31711);
or U35543 (N_35543,N_32038,N_31873);
xor U35544 (N_35544,N_34624,N_33998);
nor U35545 (N_35545,N_34769,N_30616);
nand U35546 (N_35546,N_34650,N_32223);
and U35547 (N_35547,N_30310,N_34199);
or U35548 (N_35548,N_33630,N_33676);
nor U35549 (N_35549,N_31539,N_34203);
nand U35550 (N_35550,N_30085,N_33012);
xor U35551 (N_35551,N_34176,N_34775);
nor U35552 (N_35552,N_33692,N_32089);
and U35553 (N_35553,N_33711,N_34560);
nor U35554 (N_35554,N_34915,N_30375);
and U35555 (N_35555,N_31998,N_30713);
or U35556 (N_35556,N_34381,N_31853);
nand U35557 (N_35557,N_34849,N_32958);
nor U35558 (N_35558,N_30729,N_31224);
nand U35559 (N_35559,N_32514,N_33912);
nand U35560 (N_35560,N_32659,N_33793);
nor U35561 (N_35561,N_30648,N_33850);
nor U35562 (N_35562,N_33535,N_30865);
nor U35563 (N_35563,N_30838,N_30404);
nand U35564 (N_35564,N_34405,N_33448);
and U35565 (N_35565,N_34391,N_33827);
xor U35566 (N_35566,N_30690,N_30319);
and U35567 (N_35567,N_33956,N_33908);
nor U35568 (N_35568,N_34395,N_31517);
nand U35569 (N_35569,N_33710,N_30231);
nor U35570 (N_35570,N_31372,N_33185);
and U35571 (N_35571,N_34784,N_31483);
or U35572 (N_35572,N_33664,N_32048);
and U35573 (N_35573,N_33903,N_33089);
nor U35574 (N_35574,N_33726,N_31469);
nand U35575 (N_35575,N_30281,N_30062);
and U35576 (N_35576,N_32407,N_34048);
and U35577 (N_35577,N_32690,N_30307);
xor U35578 (N_35578,N_34079,N_32905);
or U35579 (N_35579,N_32654,N_31254);
and U35580 (N_35580,N_34065,N_31150);
nand U35581 (N_35581,N_33253,N_33707);
nand U35582 (N_35582,N_31347,N_33411);
xor U35583 (N_35583,N_34179,N_30440);
and U35584 (N_35584,N_34466,N_33399);
nand U35585 (N_35585,N_33000,N_30366);
or U35586 (N_35586,N_32653,N_32497);
or U35587 (N_35587,N_30994,N_34058);
and U35588 (N_35588,N_30811,N_34256);
xor U35589 (N_35589,N_30541,N_33251);
nor U35590 (N_35590,N_34832,N_32012);
or U35591 (N_35591,N_34158,N_32176);
nor U35592 (N_35592,N_34230,N_34224);
xnor U35593 (N_35593,N_34040,N_33246);
nor U35594 (N_35594,N_31033,N_33928);
nand U35595 (N_35595,N_30770,N_31257);
and U35596 (N_35596,N_32638,N_32734);
nor U35597 (N_35597,N_33694,N_30933);
nor U35598 (N_35598,N_33255,N_33518);
or U35599 (N_35599,N_33583,N_32382);
nor U35600 (N_35600,N_30717,N_31958);
or U35601 (N_35601,N_30790,N_33300);
and U35602 (N_35602,N_33302,N_32549);
xnor U35603 (N_35603,N_31730,N_33095);
nand U35604 (N_35604,N_32324,N_34333);
or U35605 (N_35605,N_34759,N_34957);
nand U35606 (N_35606,N_33118,N_31680);
nand U35607 (N_35607,N_33900,N_31213);
xnor U35608 (N_35608,N_34252,N_33239);
and U35609 (N_35609,N_33225,N_30877);
xor U35610 (N_35610,N_30282,N_30785);
or U35611 (N_35611,N_31960,N_31038);
xor U35612 (N_35612,N_33262,N_34632);
xnor U35613 (N_35613,N_30008,N_34121);
nor U35614 (N_35614,N_34184,N_30693);
xnor U35615 (N_35615,N_33491,N_33695);
and U35616 (N_35616,N_31579,N_32823);
and U35617 (N_35617,N_31784,N_30955);
xnor U35618 (N_35618,N_30926,N_30527);
and U35619 (N_35619,N_33708,N_34951);
nand U35620 (N_35620,N_31937,N_30013);
and U35621 (N_35621,N_32126,N_34945);
and U35622 (N_35622,N_30724,N_34346);
xor U35623 (N_35623,N_33515,N_31542);
xor U35624 (N_35624,N_34337,N_30497);
and U35625 (N_35625,N_34149,N_30407);
nor U35626 (N_35626,N_34920,N_34371);
nand U35627 (N_35627,N_31693,N_33934);
and U35628 (N_35628,N_30806,N_33716);
and U35629 (N_35629,N_30715,N_34168);
xnor U35630 (N_35630,N_34676,N_34756);
xor U35631 (N_35631,N_32626,N_31522);
xnor U35632 (N_35632,N_33873,N_33836);
and U35633 (N_35633,N_31173,N_33013);
nand U35634 (N_35634,N_33883,N_31888);
xor U35635 (N_35635,N_31360,N_31612);
or U35636 (N_35636,N_34909,N_31959);
nor U35637 (N_35637,N_32846,N_30080);
or U35638 (N_35638,N_33816,N_30341);
and U35639 (N_35639,N_31315,N_31660);
xnor U35640 (N_35640,N_34730,N_32602);
or U35641 (N_35641,N_30797,N_34755);
or U35642 (N_35642,N_30138,N_31696);
xnor U35643 (N_35643,N_31816,N_31039);
or U35644 (N_35644,N_33815,N_30154);
nor U35645 (N_35645,N_30879,N_34043);
or U35646 (N_35646,N_34573,N_33331);
nor U35647 (N_35647,N_31036,N_33132);
nor U35648 (N_35648,N_32002,N_33163);
or U35649 (N_35649,N_30236,N_33152);
or U35650 (N_35650,N_30552,N_32631);
nand U35651 (N_35651,N_33801,N_34088);
or U35652 (N_35652,N_34545,N_34839);
and U35653 (N_35653,N_33461,N_31188);
nor U35654 (N_35654,N_32213,N_34663);
and U35655 (N_35655,N_31061,N_34375);
xnor U35656 (N_35656,N_31145,N_30033);
nand U35657 (N_35657,N_33166,N_30950);
nand U35658 (N_35658,N_33207,N_34984);
nand U35659 (N_35659,N_33530,N_31415);
nand U35660 (N_35660,N_34693,N_31790);
or U35661 (N_35661,N_33880,N_34372);
xnor U35662 (N_35662,N_30916,N_30617);
and U35663 (N_35663,N_30373,N_31951);
or U35664 (N_35664,N_30219,N_34813);
nand U35665 (N_35665,N_31668,N_34130);
and U35666 (N_35666,N_33892,N_31010);
xnor U35667 (N_35667,N_32853,N_33965);
or U35668 (N_35668,N_34164,N_31390);
nand U35669 (N_35669,N_30238,N_33447);
and U35670 (N_35670,N_32017,N_32028);
or U35671 (N_35671,N_32307,N_31823);
and U35672 (N_35672,N_31862,N_33389);
nor U35673 (N_35673,N_34872,N_33248);
xor U35674 (N_35674,N_31629,N_30336);
and U35675 (N_35675,N_33113,N_30539);
xor U35676 (N_35676,N_30430,N_34903);
or U35677 (N_35677,N_30542,N_34703);
nor U35678 (N_35678,N_34473,N_33178);
nor U35679 (N_35679,N_34178,N_32844);
xor U35680 (N_35680,N_33832,N_31641);
nor U35681 (N_35681,N_31020,N_30768);
nor U35682 (N_35682,N_31642,N_34694);
nor U35683 (N_35683,N_30156,N_30516);
or U35684 (N_35684,N_34141,N_32116);
nor U35685 (N_35685,N_30159,N_31872);
nand U35686 (N_35686,N_31487,N_33514);
nand U35687 (N_35687,N_34236,N_30589);
nor U35688 (N_35688,N_32871,N_31596);
and U35689 (N_35689,N_30034,N_31655);
nand U35690 (N_35690,N_34904,N_33781);
nor U35691 (N_35691,N_31661,N_31136);
and U35692 (N_35692,N_30510,N_32575);
nand U35693 (N_35693,N_30218,N_30072);
or U35694 (N_35694,N_30178,N_30202);
xor U35695 (N_35695,N_34936,N_33942);
xor U35696 (N_35696,N_32597,N_31395);
nand U35697 (N_35697,N_33304,N_34474);
nor U35698 (N_35698,N_31283,N_30367);
nand U35699 (N_35699,N_34815,N_31553);
nand U35700 (N_35700,N_33060,N_30247);
xor U35701 (N_35701,N_32889,N_33453);
and U35702 (N_35702,N_34583,N_33562);
nand U35703 (N_35703,N_31086,N_31235);
or U35704 (N_35704,N_30704,N_33226);
nand U35705 (N_35705,N_30653,N_32996);
or U35706 (N_35706,N_31216,N_30425);
nor U35707 (N_35707,N_30109,N_31000);
xor U35708 (N_35708,N_32370,N_32412);
nand U35709 (N_35709,N_31817,N_33808);
or U35710 (N_35710,N_32866,N_31719);
and U35711 (N_35711,N_34442,N_30708);
nand U35712 (N_35712,N_34259,N_31220);
or U35713 (N_35713,N_31549,N_31572);
nor U35714 (N_35714,N_30977,N_33324);
nand U35715 (N_35715,N_32742,N_32113);
xor U35716 (N_35716,N_33962,N_30448);
xnor U35717 (N_35717,N_33421,N_33971);
nor U35718 (N_35718,N_33612,N_33607);
or U35719 (N_35719,N_33454,N_31701);
nor U35720 (N_35720,N_31625,N_32311);
and U35721 (N_35721,N_32547,N_30153);
or U35722 (N_35722,N_34797,N_32416);
or U35723 (N_35723,N_30003,N_31555);
or U35724 (N_35724,N_34290,N_33117);
xnor U35725 (N_35725,N_32338,N_31307);
and U35726 (N_35726,N_32208,N_33768);
xnor U35727 (N_35727,N_31826,N_30151);
nor U35728 (N_35728,N_34974,N_31097);
nand U35729 (N_35729,N_34255,N_33600);
and U35730 (N_35730,N_31628,N_31411);
nor U35731 (N_35731,N_30388,N_33298);
or U35732 (N_35732,N_33966,N_30139);
and U35733 (N_35733,N_34327,N_32112);
nand U35734 (N_35734,N_32377,N_34882);
nand U35735 (N_35735,N_32951,N_34889);
xnor U35736 (N_35736,N_30575,N_33806);
nand U35737 (N_35737,N_30344,N_31626);
nor U35738 (N_35738,N_30031,N_33736);
nand U35739 (N_35739,N_30246,N_31068);
nand U35740 (N_35740,N_31739,N_32175);
or U35741 (N_35741,N_32764,N_34823);
and U35742 (N_35742,N_32148,N_30866);
xnor U35743 (N_35743,N_33550,N_31635);
and U35744 (N_35744,N_33655,N_32703);
nand U35745 (N_35745,N_31264,N_33071);
nand U35746 (N_35746,N_30065,N_34225);
or U35747 (N_35747,N_32391,N_33617);
nand U35748 (N_35748,N_31753,N_31318);
or U35749 (N_35749,N_30878,N_33426);
and U35750 (N_35750,N_34217,N_30021);
nor U35751 (N_35751,N_33990,N_33083);
xor U35752 (N_35752,N_31747,N_34525);
or U35753 (N_35753,N_32226,N_34532);
and U35754 (N_35754,N_31388,N_32147);
and U35755 (N_35755,N_31672,N_34219);
or U35756 (N_35756,N_32034,N_32277);
and U35757 (N_35757,N_32538,N_34999);
or U35758 (N_35758,N_30249,N_34885);
nand U35759 (N_35759,N_33007,N_30682);
or U35760 (N_35760,N_32760,N_34469);
xor U35761 (N_35761,N_34456,N_32124);
nor U35762 (N_35762,N_33894,N_34161);
or U35763 (N_35763,N_31015,N_32962);
or U35764 (N_35764,N_31129,N_30043);
nand U35765 (N_35765,N_34992,N_30393);
nand U35766 (N_35766,N_30473,N_32925);
and U35767 (N_35767,N_33840,N_31157);
or U35768 (N_35768,N_33725,N_33829);
nand U35769 (N_35769,N_33444,N_34778);
or U35770 (N_35770,N_30512,N_34119);
xnor U35771 (N_35771,N_34274,N_31526);
nor U35772 (N_35772,N_32814,N_30122);
nor U35773 (N_35773,N_32166,N_33522);
nor U35774 (N_35774,N_33347,N_30173);
or U35775 (N_35775,N_30741,N_33696);
nand U35776 (N_35776,N_32822,N_34108);
nand U35777 (N_35777,N_31671,N_32856);
nor U35778 (N_35778,N_30007,N_33318);
nor U35779 (N_35779,N_31929,N_31955);
xor U35780 (N_35780,N_31427,N_34026);
and U35781 (N_35781,N_32348,N_30095);
nand U35782 (N_35782,N_31072,N_31768);
and U35783 (N_35783,N_33127,N_34014);
or U35784 (N_35784,N_33642,N_33450);
nand U35785 (N_35785,N_32481,N_32344);
and U35786 (N_35786,N_32031,N_34312);
xor U35787 (N_35787,N_30749,N_33428);
nor U35788 (N_35788,N_34574,N_33917);
and U35789 (N_35789,N_32804,N_33319);
nand U35790 (N_35790,N_34552,N_32930);
nand U35791 (N_35791,N_30411,N_34981);
or U35792 (N_35792,N_32172,N_34506);
xnor U35793 (N_35793,N_31512,N_30167);
and U35794 (N_35794,N_34943,N_34542);
and U35795 (N_35795,N_32900,N_31986);
and U35796 (N_35796,N_33513,N_32074);
and U35797 (N_35797,N_34428,N_31007);
or U35798 (N_35798,N_34540,N_30760);
or U35799 (N_35799,N_33734,N_30015);
nand U35800 (N_35800,N_34873,N_33969);
xor U35801 (N_35801,N_34417,N_31444);
nand U35802 (N_35802,N_31217,N_30507);
nor U35803 (N_35803,N_32396,N_32679);
and U35804 (N_35804,N_34279,N_33275);
nand U35805 (N_35805,N_34979,N_34244);
or U35806 (N_35806,N_34561,N_31420);
nand U35807 (N_35807,N_31477,N_32821);
and U35808 (N_35808,N_32293,N_30964);
and U35809 (N_35809,N_34605,N_34155);
nor U35810 (N_35810,N_33789,N_30800);
nor U35811 (N_35811,N_30470,N_31878);
nand U35812 (N_35812,N_30909,N_34046);
or U35813 (N_35813,N_33763,N_30241);
nor U35814 (N_35814,N_34211,N_32231);
or U35815 (N_35815,N_34389,N_31228);
xor U35816 (N_35816,N_33145,N_32458);
nor U35817 (N_35817,N_33029,N_32341);
xor U35818 (N_35818,N_34227,N_32182);
and U35819 (N_35819,N_32969,N_34870);
and U35820 (N_35820,N_31819,N_30243);
xnor U35821 (N_35821,N_32184,N_31244);
nor U35822 (N_35822,N_34691,N_34868);
and U35823 (N_35823,N_30324,N_33341);
nand U35824 (N_35824,N_31299,N_31128);
or U35825 (N_35825,N_31236,N_33022);
nand U35826 (N_35826,N_30286,N_31558);
xor U35827 (N_35827,N_32987,N_31466);
nor U35828 (N_35828,N_34427,N_34152);
xor U35829 (N_35829,N_30765,N_32792);
xnor U35830 (N_35830,N_30229,N_33621);
nor U35831 (N_35831,N_33987,N_33503);
and U35832 (N_35832,N_32674,N_31354);
nand U35833 (N_35833,N_31847,N_34233);
nand U35834 (N_35834,N_33633,N_30787);
xor U35835 (N_35835,N_34005,N_32301);
nor U35836 (N_35836,N_31399,N_33376);
nand U35837 (N_35837,N_34833,N_31501);
nor U35838 (N_35838,N_33303,N_30721);
xor U35839 (N_35839,N_34134,N_32490);
or U35840 (N_35840,N_30157,N_32114);
xor U35841 (N_35841,N_34591,N_32162);
and U35842 (N_35842,N_32107,N_32192);
nor U35843 (N_35843,N_31833,N_33819);
nor U35844 (N_35844,N_30851,N_30297);
xor U35845 (N_35845,N_32100,N_34029);
and U35846 (N_35846,N_31577,N_30559);
and U35847 (N_35847,N_30227,N_30403);
or U35848 (N_35848,N_33554,N_32203);
nor U35849 (N_35849,N_33737,N_34851);
nand U35850 (N_35850,N_32440,N_33929);
nand U35851 (N_35851,N_32143,N_33723);
xor U35852 (N_35852,N_34724,N_34246);
and U35853 (N_35853,N_33672,N_30184);
or U35854 (N_35854,N_31764,N_31456);
xor U35855 (N_35855,N_34317,N_34123);
or U35856 (N_35856,N_31293,N_31777);
nor U35857 (N_35857,N_33826,N_34821);
xnor U35858 (N_35858,N_31848,N_31462);
nor U35859 (N_35859,N_33006,N_31455);
nor U35860 (N_35860,N_31900,N_32133);
nand U35861 (N_35861,N_31118,N_31834);
nor U35862 (N_35862,N_32058,N_34906);
nor U35863 (N_35863,N_32376,N_30049);
or U35864 (N_35864,N_31066,N_33086);
nand U35865 (N_35865,N_31796,N_33489);
xor U35866 (N_35866,N_33400,N_32775);
xor U35867 (N_35867,N_31386,N_30078);
nor U35868 (N_35868,N_32719,N_32733);
and U35869 (N_35869,N_33084,N_34434);
or U35870 (N_35870,N_33419,N_31850);
or U35871 (N_35871,N_34735,N_31795);
nor U35872 (N_35872,N_34516,N_30680);
nor U35873 (N_35873,N_31300,N_34073);
nor U35874 (N_35874,N_31273,N_34527);
nor U35875 (N_35875,N_33091,N_30903);
xnor U35876 (N_35876,N_34665,N_30147);
nand U35877 (N_35877,N_31925,N_31966);
or U35878 (N_35878,N_30261,N_32533);
or U35879 (N_35879,N_34242,N_32426);
or U35880 (N_35880,N_30481,N_30019);
and U35881 (N_35881,N_33391,N_34218);
or U35882 (N_35882,N_30813,N_30674);
nand U35883 (N_35883,N_30691,N_32479);
or U35884 (N_35884,N_34471,N_34007);
and U35885 (N_35885,N_32085,N_32650);
or U35886 (N_35886,N_34757,N_34639);
nor U35887 (N_35887,N_31899,N_33616);
xnor U35888 (N_35888,N_30100,N_33266);
or U35889 (N_35889,N_30703,N_33974);
or U35890 (N_35890,N_31903,N_33649);
and U35891 (N_35891,N_31911,N_33982);
and U35892 (N_35892,N_32519,N_34781);
xnor U35893 (N_35893,N_31156,N_30082);
nor U35894 (N_35894,N_31298,N_33078);
xnor U35895 (N_35895,N_33561,N_32569);
xnor U35896 (N_35896,N_30896,N_30670);
and U35897 (N_35897,N_34547,N_30044);
and U35898 (N_35898,N_31211,N_32812);
nor U35899 (N_35899,N_32279,N_31785);
xnor U35900 (N_35900,N_30200,N_33328);
and U35901 (N_35901,N_32620,N_30540);
and U35902 (N_35902,N_32123,N_34091);
xor U35903 (N_35903,N_31195,N_33730);
xor U35904 (N_35904,N_33751,N_33414);
xor U35905 (N_35905,N_34145,N_34305);
xor U35906 (N_35906,N_33779,N_32007);
and U35907 (N_35907,N_34095,N_34923);
nand U35908 (N_35908,N_32464,N_33661);
xor U35909 (N_35909,N_33433,N_30306);
xnor U35910 (N_35910,N_31369,N_32995);
nand U35911 (N_35911,N_30683,N_30364);
nor U35912 (N_35912,N_31245,N_34954);
xnor U35913 (N_35913,N_31602,N_34288);
xnor U35914 (N_35914,N_32554,N_30771);
nand U35915 (N_35915,N_34056,N_30782);
nor U35916 (N_35916,N_33677,N_34596);
and U35917 (N_35917,N_32806,N_33352);
nor U35918 (N_35918,N_34332,N_30992);
xnor U35919 (N_35919,N_32724,N_33229);
and U35920 (N_35920,N_32789,N_32903);
nor U35921 (N_35921,N_33783,N_31053);
and U35922 (N_35922,N_31123,N_30571);
nor U35923 (N_35923,N_33943,N_32070);
nand U35924 (N_35924,N_32328,N_33374);
xor U35925 (N_35925,N_34369,N_33156);
xor U35926 (N_35926,N_32387,N_32664);
or U35927 (N_35927,N_31940,N_34097);
nand U35928 (N_35928,N_34578,N_30023);
or U35929 (N_35929,N_33346,N_34114);
xor U35930 (N_35930,N_34702,N_33353);
xnor U35931 (N_35931,N_34090,N_32534);
and U35932 (N_35932,N_31083,N_32437);
and U35933 (N_35933,N_32669,N_33228);
or U35934 (N_35934,N_34673,N_33728);
nor U35935 (N_35935,N_32907,N_32265);
and U35936 (N_35936,N_32187,N_34568);
xnor U35937 (N_35937,N_31639,N_31004);
xnor U35938 (N_35938,N_32827,N_31090);
or U35939 (N_35939,N_32920,N_34692);
or U35940 (N_35940,N_34010,N_32710);
nor U35941 (N_35941,N_30454,N_33221);
or U35942 (N_35942,N_31758,N_31994);
xor U35943 (N_35943,N_30090,N_34698);
xor U35944 (N_35944,N_31614,N_30222);
nor U35945 (N_35945,N_30235,N_34774);
and U35946 (N_35946,N_31541,N_33834);
or U35947 (N_35947,N_30092,N_31237);
and U35948 (N_35948,N_31725,N_30189);
or U35949 (N_35949,N_30273,N_34320);
or U35950 (N_35950,N_30829,N_32886);
and U35951 (N_35951,N_30947,N_33653);
xnor U35952 (N_35952,N_31345,N_31875);
and U35953 (N_35953,N_30566,N_31169);
nand U35954 (N_35954,N_34983,N_33682);
xor U35955 (N_35955,N_31024,N_31088);
xnor U35956 (N_35956,N_32545,N_33509);
nor U35957 (N_35957,N_33915,N_30205);
nor U35958 (N_35958,N_32499,N_32474);
and U35959 (N_35959,N_30906,N_32922);
nor U35960 (N_35960,N_31200,N_32614);
or U35961 (N_35961,N_32833,N_32824);
or U35962 (N_35962,N_31835,N_30477);
nand U35963 (N_35963,N_32261,N_34621);
xor U35964 (N_35964,N_30808,N_31676);
nand U35965 (N_35965,N_30945,N_30871);
and U35966 (N_35966,N_30621,N_32132);
nand U35967 (N_35967,N_34791,N_34677);
xor U35968 (N_35968,N_31771,N_32216);
nor U35969 (N_35969,N_30318,N_33187);
nand U35970 (N_35970,N_33098,N_32398);
nand U35971 (N_35971,N_33754,N_34557);
and U35972 (N_35972,N_31776,N_30893);
or U35973 (N_35973,N_32227,N_30185);
xnor U35974 (N_35974,N_34470,N_32077);
and U35975 (N_35975,N_32603,N_31458);
nor U35976 (N_35976,N_31861,N_31406);
xnor U35977 (N_35977,N_30359,N_31074);
xnor U35978 (N_35978,N_31365,N_31654);
nor U35979 (N_35979,N_31623,N_32874);
and U35980 (N_35980,N_32081,N_31547);
nand U35981 (N_35981,N_34679,N_33555);
and U35982 (N_35982,N_34965,N_33088);
xor U35983 (N_35983,N_34526,N_34620);
and U35984 (N_35984,N_33093,N_33924);
or U35985 (N_35985,N_30186,N_32711);
xnor U35986 (N_35986,N_31845,N_33471);
xnor U35987 (N_35987,N_30384,N_30757);
xnor U35988 (N_35988,N_32882,N_33383);
nand U35989 (N_35989,N_34968,N_30781);
and U35990 (N_35990,N_33267,N_33796);
xor U35991 (N_35991,N_32748,N_30496);
or U35992 (N_35992,N_32933,N_30355);
and U35993 (N_35993,N_32420,N_34640);
nor U35994 (N_35994,N_31181,N_30604);
nor U35995 (N_35995,N_30194,N_34263);
xor U35996 (N_35996,N_33930,N_31567);
xnor U35997 (N_35997,N_30537,N_34483);
nor U35998 (N_35998,N_33196,N_34409);
xnor U35999 (N_35999,N_32944,N_32119);
nor U36000 (N_36000,N_31857,N_34365);
nor U36001 (N_36001,N_31530,N_33323);
nand U36002 (N_36002,N_33945,N_31756);
or U36003 (N_36003,N_31545,N_33927);
and U36004 (N_36004,N_30594,N_32140);
xnor U36005 (N_36005,N_31766,N_34762);
nand U36006 (N_36006,N_30940,N_31067);
and U36007 (N_36007,N_34421,N_30998);
xnor U36008 (N_36008,N_31353,N_33963);
nor U36009 (N_36009,N_34352,N_33954);
xor U36010 (N_36010,N_34490,N_34612);
nor U36011 (N_36011,N_32671,N_34201);
nor U36012 (N_36012,N_33641,N_33752);
xnor U36013 (N_36013,N_31697,N_32639);
or U36014 (N_36014,N_32503,N_31154);
or U36015 (N_36015,N_30980,N_32553);
nand U36016 (N_36016,N_33270,N_30695);
nor U36017 (N_36017,N_33546,N_30557);
nand U36018 (N_36018,N_30130,N_33351);
or U36019 (N_36019,N_32779,N_31924);
and U36020 (N_36020,N_32847,N_34359);
or U36021 (N_36021,N_31839,N_31812);
and U36022 (N_36022,N_33065,N_31115);
nor U36023 (N_36023,N_34300,N_34100);
nor U36024 (N_36024,N_30111,N_33507);
and U36025 (N_36025,N_30793,N_34842);
xor U36026 (N_36026,N_32696,N_31215);
or U36027 (N_36027,N_31695,N_34948);
xnor U36028 (N_36028,N_34140,N_30164);
nand U36029 (N_36029,N_34705,N_30938);
and U36030 (N_36030,N_33622,N_33051);
nor U36031 (N_36031,N_34323,N_33946);
nand U36032 (N_36032,N_32418,N_34924);
or U36033 (N_36033,N_34344,N_33237);
xnor U36034 (N_36034,N_34188,N_30463);
and U36035 (N_36035,N_31735,N_32815);
nand U36036 (N_36036,N_33479,N_30565);
or U36037 (N_36037,N_33438,N_31745);
xnor U36038 (N_36038,N_30352,N_31939);
nand U36039 (N_36039,N_34210,N_33920);
or U36040 (N_36040,N_31830,N_31535);
xor U36041 (N_36041,N_34406,N_33068);
nor U36042 (N_36042,N_34478,N_33485);
or U36043 (N_36043,N_33372,N_33778);
nor U36044 (N_36044,N_34446,N_32365);
and U36045 (N_36045,N_30855,N_34122);
nand U36046 (N_36046,N_34914,N_31251);
nor U36047 (N_36047,N_30170,N_30298);
or U36048 (N_36048,N_30910,N_32852);
or U36049 (N_36049,N_30464,N_30224);
nor U36050 (N_36050,N_30094,N_33953);
xnor U36051 (N_36051,N_32994,N_31189);
and U36052 (N_36052,N_31849,N_31493);
and U36053 (N_36053,N_32830,N_34500);
nand U36054 (N_36054,N_30191,N_34633);
or U36055 (N_36055,N_31287,N_30188);
or U36056 (N_36056,N_31502,N_30409);
and U36057 (N_36057,N_33200,N_30446);
xor U36058 (N_36058,N_31636,N_34143);
and U36059 (N_36059,N_33080,N_30315);
nand U36060 (N_36060,N_32701,N_34773);
nor U36061 (N_36061,N_34117,N_33418);
xor U36062 (N_36062,N_30503,N_34402);
nand U36063 (N_36063,N_32305,N_31575);
nor U36064 (N_36064,N_34459,N_30740);
and U36065 (N_36065,N_30207,N_31294);
nand U36066 (N_36066,N_30502,N_33891);
nor U36067 (N_36067,N_30106,N_34415);
nor U36068 (N_36068,N_30967,N_32750);
xor U36069 (N_36069,N_32768,N_33579);
nand U36070 (N_36070,N_34859,N_30456);
nand U36071 (N_36071,N_31142,N_30719);
nor U36072 (N_36072,N_32767,N_33339);
and U36073 (N_36073,N_33325,N_32729);
or U36074 (N_36074,N_34785,N_33666);
nor U36075 (N_36075,N_32591,N_30066);
and U36076 (N_36076,N_30777,N_31800);
and U36077 (N_36077,N_31583,N_32403);
or U36078 (N_36078,N_34249,N_31824);
xor U36079 (N_36079,N_32101,N_34382);
and U36080 (N_36080,N_33278,N_32151);
nor U36081 (N_36081,N_32141,N_32813);
xor U36082 (N_36082,N_34064,N_33468);
or U36083 (N_36083,N_30880,N_34517);
and U36084 (N_36084,N_31908,N_32963);
or U36085 (N_36085,N_34137,N_34101);
nor U36086 (N_36086,N_31461,N_33863);
xor U36087 (N_36087,N_33215,N_34181);
and U36088 (N_36088,N_33160,N_33877);
or U36089 (N_36089,N_33629,N_34800);
or U36090 (N_36090,N_34397,N_33563);
and U36091 (N_36091,N_31765,N_31278);
or U36092 (N_36092,N_34646,N_31460);
or U36093 (N_36093,N_31837,N_32485);
or U36094 (N_36094,N_32120,N_32315);
or U36095 (N_36095,N_32380,N_31673);
and U36096 (N_36096,N_32961,N_33572);
xnor U36097 (N_36097,N_34113,N_31342);
and U36098 (N_36098,N_31412,N_30647);
and U36099 (N_36099,N_34997,N_31537);
or U36100 (N_36100,N_30350,N_30240);
xor U36101 (N_36101,N_31095,N_34038);
nand U36102 (N_36102,N_32097,N_32483);
nand U36103 (N_36103,N_34856,N_32838);
nand U36104 (N_36104,N_33854,N_31863);
nor U36105 (N_36105,N_31239,N_34202);
xnor U36106 (N_36106,N_32527,N_33259);
or U36107 (N_36107,N_33862,N_31087);
and U36108 (N_36108,N_31500,N_31378);
or U36109 (N_36109,N_30792,N_30248);
or U36110 (N_36110,N_31586,N_33493);
xnor U36111 (N_36111,N_34052,N_34034);
and U36112 (N_36112,N_31060,N_33143);
nand U36113 (N_36113,N_30514,N_33496);
nor U36114 (N_36114,N_31027,N_31775);
xor U36115 (N_36115,N_30091,N_33637);
nor U36116 (N_36116,N_32531,N_32066);
or U36117 (N_36117,N_32008,N_33654);
nor U36118 (N_36118,N_34033,N_31260);
and U36119 (N_36119,N_33487,N_33232);
nand U36120 (N_36120,N_31644,N_33159);
nor U36121 (N_36121,N_33142,N_33112);
nor U36122 (N_36122,N_34196,N_31773);
or U36123 (N_36123,N_31992,N_31355);
or U36124 (N_36124,N_34062,N_30269);
nor U36125 (N_36125,N_34489,N_30988);
xnor U36126 (N_36126,N_32727,N_34763);
xnor U36127 (N_36127,N_31203,N_33972);
nand U36128 (N_36128,N_31402,N_34022);
nor U36129 (N_36129,N_31075,N_33814);
and U36130 (N_36130,N_30957,N_32004);
xor U36131 (N_36131,N_31779,N_32699);
and U36132 (N_36132,N_30076,N_31423);
nor U36133 (N_36133,N_34553,N_33204);
nor U36134 (N_36134,N_30203,N_31667);
nand U36135 (N_36135,N_34304,N_32752);
xnor U36136 (N_36136,N_34297,N_33042);
or U36137 (N_36137,N_31312,N_34511);
and U36138 (N_36138,N_32787,N_30179);
and U36139 (N_36139,N_32419,N_31825);
nand U36140 (N_36140,N_34157,N_30075);
nand U36141 (N_36141,N_33717,N_34594);
or U36142 (N_36142,N_34714,N_30163);
and U36143 (N_36143,N_30317,N_34913);
nor U36144 (N_36144,N_31163,N_31003);
and U36145 (N_36145,N_30922,N_30048);
xnor U36146 (N_36146,N_34047,N_30745);
nor U36147 (N_36147,N_33023,N_32249);
nand U36148 (N_36148,N_32308,N_32952);
nor U36149 (N_36149,N_31631,N_34847);
nor U36150 (N_36150,N_31504,N_32052);
and U36151 (N_36151,N_32875,N_30217);
nor U36152 (N_36152,N_31159,N_31854);
and U36153 (N_36153,N_30279,N_30469);
nand U36154 (N_36154,N_31916,N_33644);
xnor U36155 (N_36155,N_34247,N_33648);
or U36156 (N_36156,N_31116,N_32239);
nor U36157 (N_36157,N_31684,N_32233);
xnor U36158 (N_36158,N_30796,N_34275);
or U36159 (N_36159,N_31685,N_31080);
xor U36160 (N_36160,N_33855,N_34066);
nor U36161 (N_36161,N_32400,N_31574);
or U36162 (N_36162,N_33155,N_30449);
nor U36163 (N_36163,N_30152,N_34701);
nand U36164 (N_36164,N_33462,N_31513);
nor U36165 (N_36165,N_33040,N_32206);
nor U36166 (N_36166,N_34457,N_32271);
and U36167 (N_36167,N_32751,N_34479);
or U36168 (N_36168,N_34963,N_33307);
xnor U36169 (N_36169,N_32641,N_34175);
and U36170 (N_36170,N_33092,N_32890);
xnor U36171 (N_36171,N_34546,N_30979);
nand U36172 (N_36172,N_34298,N_32244);
nand U36173 (N_36173,N_34514,N_31829);
nand U36174 (N_36174,N_32772,N_33662);
xor U36175 (N_36175,N_34827,N_33289);
nor U36176 (N_36176,N_30242,N_32574);
xnor U36177 (N_36177,N_30025,N_32515);
xor U36178 (N_36178,N_30732,N_30032);
xnor U36179 (N_36179,N_33497,N_30491);
and U36180 (N_36180,N_30615,N_33287);
or U36181 (N_36181,N_34081,N_30551);
and U36182 (N_36182,N_31949,N_33564);
or U36183 (N_36183,N_31314,N_31550);
nor U36184 (N_36184,N_31592,N_30974);
nor U36185 (N_36185,N_30396,N_30474);
and U36186 (N_36186,N_34384,N_30221);
nor U36187 (N_36187,N_34501,N_30915);
nand U36188 (N_36188,N_34810,N_32477);
and U36189 (N_36189,N_32243,N_34092);
or U36190 (N_36190,N_32496,N_30234);
xnor U36191 (N_36191,N_31304,N_33123);
xor U36192 (N_36192,N_34515,N_30030);
nand U36193 (N_36193,N_32510,N_34004);
xnor U36194 (N_36194,N_31190,N_30026);
and U36195 (N_36195,N_34376,N_33817);
or U36196 (N_36196,N_31990,N_32280);
xnor U36197 (N_36197,N_34543,N_34390);
or U36198 (N_36198,N_33128,N_32159);
xor U36199 (N_36199,N_33597,N_32904);
nor U36200 (N_36200,N_30746,N_30018);
and U36201 (N_36201,N_30546,N_31025);
and U36202 (N_36202,N_30583,N_32938);
and U36203 (N_36203,N_31049,N_32523);
xor U36204 (N_36204,N_34884,N_33321);
nand U36205 (N_36205,N_34518,N_34462);
or U36206 (N_36206,N_32428,N_31176);
nor U36207 (N_36207,N_32330,N_31869);
xor U36208 (N_36208,N_34378,N_32295);
or U36209 (N_36209,N_31155,N_31632);
or U36210 (N_36210,N_34682,N_34793);
nand U36211 (N_36211,N_30408,N_33847);
and U36212 (N_36212,N_32323,N_31030);
and U36213 (N_36213,N_33423,N_30882);
xor U36214 (N_36214,N_32029,N_30976);
xor U36215 (N_36215,N_33940,N_34706);
nor U36216 (N_36216,N_34392,N_30673);
and U36217 (N_36217,N_32046,N_34549);
nand U36218 (N_36218,N_30612,N_32794);
or U36219 (N_36219,N_32039,N_32898);
and U36220 (N_36220,N_32468,N_30895);
and U36221 (N_36221,N_32913,N_32773);
nand U36222 (N_36222,N_33576,N_34513);
and U36223 (N_36223,N_30284,N_30328);
or U36224 (N_36224,N_32343,N_31792);
xor U36225 (N_36225,N_31576,N_31409);
nand U36226 (N_36226,N_31459,N_34235);
nor U36227 (N_36227,N_33271,N_31026);
or U36228 (N_36228,N_34745,N_34342);
or U36229 (N_36229,N_34750,N_32318);
nor U36230 (N_36230,N_32862,N_32444);
nor U36231 (N_36231,N_31146,N_31379);
and U36232 (N_36232,N_30677,N_33476);
nor U36233 (N_36233,N_31063,N_32595);
and U36234 (N_36234,N_31852,N_34502);
nand U36235 (N_36235,N_30029,N_30431);
or U36236 (N_36236,N_31422,N_32179);
and U36237 (N_36237,N_30755,N_30225);
xnor U36238 (N_36238,N_31321,N_31750);
or U36239 (N_36239,N_33130,N_33236);
xor U36240 (N_36240,N_31737,N_33715);
xor U36241 (N_36241,N_33657,N_33250);
and U36242 (N_36242,N_32015,N_30971);
or U36243 (N_36243,N_32494,N_33660);
xor U36244 (N_36244,N_30457,N_31855);
and U36245 (N_36245,N_34595,N_30961);
xnor U36246 (N_36246,N_32198,N_32943);
or U36247 (N_36247,N_34021,N_30378);
nand U36248 (N_36248,N_30439,N_31568);
and U36249 (N_36249,N_34982,N_34139);
or U36250 (N_36250,N_32647,N_33422);
or U36251 (N_36251,N_31238,N_34569);
xor U36252 (N_36252,N_31243,N_31914);
or U36253 (N_36253,N_30331,N_30819);
or U36254 (N_36254,N_31375,N_33631);
nand U36255 (N_36255,N_32763,N_34308);
xnor U36256 (N_36256,N_32160,N_33254);
or U36257 (N_36257,N_31079,N_32555);
xnor U36258 (N_36258,N_34796,N_33337);
or U36259 (N_36259,N_34752,N_32462);
xnor U36260 (N_36260,N_31691,N_32229);
and U36261 (N_36261,N_34742,N_30602);
nand U36262 (N_36262,N_32762,N_34921);
nor U36263 (N_36263,N_30420,N_31584);
nor U36264 (N_36264,N_33133,N_33238);
xnor U36265 (N_36265,N_34531,N_30831);
xnor U36266 (N_36266,N_32811,N_33208);
nand U36267 (N_36267,N_34804,N_30083);
nor U36268 (N_36268,N_33604,N_30626);
or U36269 (N_36269,N_30171,N_34156);
xnor U36270 (N_36270,N_32139,N_30590);
xor U36271 (N_36271,N_31065,N_30334);
nand U36272 (N_36272,N_32983,N_34529);
nor U36273 (N_36273,N_34111,N_30501);
nand U36274 (N_36274,N_33184,N_34764);
nor U36275 (N_36275,N_30658,N_32059);
xor U36276 (N_36276,N_31818,N_33744);
nor U36277 (N_36277,N_33959,N_32110);
nand U36278 (N_36278,N_31524,N_30401);
nor U36279 (N_36279,N_34874,N_33103);
or U36280 (N_36280,N_32934,N_30925);
and U36281 (N_36281,N_32125,N_32358);
and U36282 (N_36282,N_33429,N_34078);
or U36283 (N_36283,N_30069,N_33620);
or U36284 (N_36284,N_30323,N_34129);
and U36285 (N_36285,N_31865,N_31544);
xnor U36286 (N_36286,N_34383,N_32505);
nor U36287 (N_36287,N_34674,N_33335);
and U36288 (N_36288,N_31767,N_31137);
and U36289 (N_36289,N_34401,N_30969);
or U36290 (N_36290,N_34782,N_34940);
and U36291 (N_36291,N_33598,N_31665);
and U36292 (N_36292,N_31893,N_34711);
xor U36293 (N_36293,N_32006,N_31720);
xor U36294 (N_36294,N_30905,N_31416);
nand U36295 (N_36295,N_31408,N_31580);
nand U36296 (N_36296,N_30131,N_32695);
nand U36297 (N_36297,N_34116,N_30675);
nor U36298 (N_36298,N_31252,N_34544);
nand U36299 (N_36299,N_30050,N_33545);
nor U36300 (N_36300,N_33544,N_31045);
xnor U36301 (N_36301,N_30371,N_34328);
xor U36302 (N_36302,N_30821,N_30585);
or U36303 (N_36303,N_30486,N_31448);
nor U36304 (N_36304,N_34360,N_34584);
xor U36305 (N_36305,N_33309,N_33955);
nand U36306 (N_36306,N_33064,N_32269);
nor U36307 (N_36307,N_30921,N_34978);
or U36308 (N_36308,N_32941,N_33575);
or U36309 (N_36309,N_33901,N_32732);
nand U36310 (N_36310,N_31954,N_34666);
and U36311 (N_36311,N_33999,N_30437);
nor U36312 (N_36312,N_32577,N_33524);
nand U36313 (N_36313,N_32656,N_34888);
and U36314 (N_36314,N_30860,N_31942);
or U36315 (N_36315,N_32199,N_31034);
xnor U36316 (N_36316,N_33392,N_31320);
nor U36317 (N_36317,N_33581,N_30308);
and U36318 (N_36318,N_31984,N_34205);
and U36319 (N_36319,N_30301,N_33380);
nand U36320 (N_36320,N_33977,N_34340);
nor U36321 (N_36321,N_32649,N_34281);
or U36322 (N_36322,N_34648,N_30932);
or U36323 (N_36323,N_31721,N_32469);
xor U36324 (N_36324,N_33876,N_33911);
nor U36325 (N_36325,N_34766,N_30631);
or U36326 (N_36326,N_31523,N_32425);
xor U36327 (N_36327,N_31838,N_33675);
nor U36328 (N_36328,N_33120,N_34683);
xor U36329 (N_36329,N_33290,N_31051);
nor U36330 (N_36330,N_33057,N_31292);
and U36331 (N_36331,N_32289,N_34049);
or U36332 (N_36332,N_33700,N_30622);
and U36333 (N_36333,N_30161,N_32024);
xnor U36334 (N_36334,N_33941,N_31713);
xnor U36335 (N_36335,N_32144,N_31441);
nand U36336 (N_36336,N_32608,N_32405);
and U36337 (N_36337,N_33477,N_30196);
and U36338 (N_36338,N_33944,N_31193);
xor U36339 (N_36339,N_31905,N_34622);
nor U36340 (N_36340,N_33849,N_34321);
nor U36341 (N_36341,N_31983,N_32409);
xnor U36342 (N_36342,N_34477,N_31595);
nor U36343 (N_36343,N_33825,N_34834);
and U36344 (N_36344,N_32161,N_33747);
nand U36345 (N_36345,N_34420,N_30923);
or U36346 (N_36346,N_33852,N_32248);
and U36347 (N_36347,N_31761,N_31656);
and U36348 (N_36348,N_34368,N_32861);
and U36349 (N_36349,N_32021,N_30296);
nor U36350 (N_36350,N_34958,N_34110);
xnor U36351 (N_36351,N_31965,N_30097);
or U36352 (N_36352,N_30628,N_33506);
or U36353 (N_36353,N_34899,N_34324);
nand U36354 (N_36354,N_32099,N_30867);
and U36355 (N_36355,N_31759,N_32947);
or U36356 (N_36356,N_30223,N_33771);
and U36357 (N_36357,N_32128,N_31508);
nand U36358 (N_36358,N_31557,N_32796);
or U36359 (N_36359,N_30052,N_30414);
or U36360 (N_36360,N_32250,N_32237);
and U36361 (N_36361,N_32230,N_33053);
or U36362 (N_36362,N_30022,N_31934);
or U36363 (N_36363,N_34601,N_30442);
nor U36364 (N_36364,N_30278,N_30937);
nand U36365 (N_36365,N_30433,N_30418);
xnor U36366 (N_36366,N_31233,N_31330);
nand U36367 (N_36367,N_31348,N_33914);
nor U36368 (N_36368,N_34841,N_32191);
nand U36369 (N_36369,N_30847,N_32122);
and U36370 (N_36370,N_30735,N_32616);
nand U36371 (N_36371,N_32275,N_32366);
nand U36372 (N_36372,N_32700,N_32607);
nor U36373 (N_36373,N_31168,N_30606);
or U36374 (N_36374,N_33960,N_34476);
or U36375 (N_36375,N_33993,N_30363);
nand U36376 (N_36376,N_33533,N_31482);
and U36377 (N_36377,N_31571,N_33658);
and U36378 (N_36378,N_32215,N_34163);
or U36379 (N_36379,N_30833,N_31492);
and U36380 (N_36380,N_33520,N_33986);
nor U36381 (N_36381,N_34739,N_32049);
xor U36382 (N_36382,N_33534,N_30702);
and U36383 (N_36383,N_30168,N_31891);
nor U36384 (N_36384,N_33595,N_31975);
or U36385 (N_36385,N_30166,N_31570);
xor U36386 (N_36386,N_30927,N_33810);
xnor U36387 (N_36387,N_34520,N_32537);
or U36388 (N_36388,N_32542,N_34172);
nor U36389 (N_36389,N_32984,N_33706);
or U36390 (N_36390,N_30274,N_31474);
and U36391 (N_36391,N_31963,N_31019);
or U36392 (N_36392,N_30904,N_31357);
nor U36393 (N_36393,N_33032,N_33369);
xor U36394 (N_36394,N_34707,N_31084);
and U36395 (N_36395,N_30823,N_33861);
or U36396 (N_36396,N_30593,N_33803);
or U36397 (N_36397,N_34213,N_31417);
nor U36398 (N_36398,N_33995,N_30887);
nand U36399 (N_36399,N_30581,N_30773);
nor U36400 (N_36400,N_34709,N_30733);
and U36401 (N_36401,N_32178,N_33842);
or U36402 (N_36402,N_30689,N_31484);
or U36403 (N_36403,N_31645,N_30638);
nor U36404 (N_36404,N_31326,N_34749);
xnor U36405 (N_36405,N_32286,N_33026);
and U36406 (N_36406,N_34787,N_32473);
and U36407 (N_36407,N_31961,N_32918);
and U36408 (N_36408,N_34715,N_31859);
or U36409 (N_36409,N_31716,N_31119);
or U36410 (N_36410,N_32978,N_34966);
or U36411 (N_36411,N_34316,N_32050);
nor U36412 (N_36412,N_32651,N_32876);
xnor U36413 (N_36413,N_34162,N_33234);
or U36414 (N_36414,N_32717,N_34878);
and U36415 (N_36415,N_32709,N_32640);
xor U36416 (N_36416,N_30911,N_31895);
or U36417 (N_36417,N_32253,N_34386);
or U36418 (N_36418,N_33256,N_33958);
and U36419 (N_36419,N_34484,N_31781);
and U36420 (N_36420,N_33224,N_34696);
nand U36421 (N_36421,N_30450,N_32740);
or U36422 (N_36422,N_32850,N_32692);
nand U36423 (N_36423,N_31451,N_30525);
nor U36424 (N_36424,N_31918,N_33066);
xnor U36425 (N_36425,N_31258,N_31689);
nor U36426 (N_36426,N_33443,N_30963);
or U36427 (N_36427,N_33261,N_33085);
or U36428 (N_36428,N_31491,N_30182);
and U36429 (N_36429,N_34863,N_30888);
or U36430 (N_36430,N_30475,N_33149);
and U36431 (N_36431,N_33371,N_34171);
xnor U36432 (N_36432,N_30562,N_30060);
nor U36433 (N_36433,N_34015,N_32493);
or U36434 (N_36434,N_33412,N_30694);
nor U36435 (N_36435,N_32064,N_31467);
or U36436 (N_36436,N_34425,N_33931);
nand U36437 (N_36437,N_30385,N_32668);
nor U36438 (N_36438,N_31212,N_32964);
and U36439 (N_36439,N_32892,N_34524);
xnor U36440 (N_36440,N_32173,N_30734);
or U36441 (N_36441,N_32121,N_34618);
xor U36442 (N_36442,N_30920,N_32371);
nor U36443 (N_36443,N_33076,N_34555);
or U36444 (N_36444,N_34268,N_34710);
nand U36445 (N_36445,N_32803,N_33144);
xor U36446 (N_36446,N_31752,N_32755);
xnor U36447 (N_36447,N_32157,N_32504);
and U36448 (N_36448,N_31976,N_30137);
nor U36449 (N_36449,N_34394,N_32888);
and U36450 (N_36450,N_31126,N_33592);
nand U36451 (N_36451,N_34495,N_32584);
nand U36452 (N_36452,N_33909,N_30614);
xor U36453 (N_36453,N_30000,N_33976);
nor U36454 (N_36454,N_30480,N_30671);
and U36455 (N_36455,N_34638,N_32027);
and U36456 (N_36456,N_32632,N_32103);
and U36457 (N_36457,N_33063,N_31985);
nand U36458 (N_36458,N_32693,N_33970);
xor U36459 (N_36459,N_32360,N_34076);
and U36460 (N_36460,N_33484,N_31690);
nand U36461 (N_36461,N_31247,N_33025);
nor U36462 (N_36462,N_31029,N_34609);
or U36463 (N_36463,N_32831,N_32600);
nor U36464 (N_36464,N_31351,N_33038);
and U36465 (N_36465,N_31762,N_31789);
xor U36466 (N_36466,N_34212,N_32660);
xor U36467 (N_36467,N_31101,N_34035);
and U36468 (N_36468,N_31424,N_34016);
nor U36469 (N_36469,N_32681,N_32723);
nor U36470 (N_36470,N_34844,N_30934);
nor U36471 (N_36471,N_32072,N_32832);
or U36472 (N_36472,N_34492,N_30254);
nand U36473 (N_36473,N_33776,N_30288);
and U36474 (N_36474,N_33750,N_31361);
xnor U36475 (N_36475,N_32449,N_30607);
or U36476 (N_36476,N_30901,N_30434);
nor U36477 (N_36477,N_31138,N_31394);
xnor U36478 (N_36478,N_34729,N_30495);
xor U36479 (N_36479,N_34488,N_33886);
nor U36480 (N_36480,N_30618,N_30402);
or U36481 (N_36481,N_34617,N_34248);
nor U36482 (N_36482,N_33541,N_33811);
nor U36483 (N_36483,N_33010,N_33124);
and U36484 (N_36484,N_34743,N_31141);
or U36485 (N_36485,N_34505,N_31044);
nor U36486 (N_36486,N_34925,N_33263);
nor U36487 (N_36487,N_31443,N_32353);
xor U36488 (N_36488,N_34699,N_30289);
or U36489 (N_36489,N_34964,N_34651);
and U36490 (N_36490,N_34153,N_32044);
and U36491 (N_36491,N_30445,N_31082);
nor U36492 (N_36492,N_34146,N_34441);
nor U36493 (N_36493,N_33538,N_32194);
and U36494 (N_36494,N_30413,N_33722);
nor U36495 (N_36495,N_34444,N_34438);
or U36496 (N_36496,N_32351,N_33882);
and U36497 (N_36497,N_30180,N_33041);
nand U36498 (N_36498,N_32541,N_31751);
or U36499 (N_36499,N_30339,N_33106);
xor U36500 (N_36500,N_34600,N_34458);
or U36501 (N_36501,N_34877,N_30756);
nor U36502 (N_36502,N_32421,N_34020);
nand U36503 (N_36503,N_33115,N_31185);
nor U36504 (N_36504,N_34282,N_30093);
or U36505 (N_36505,N_30874,N_32484);
and U36506 (N_36506,N_32666,N_31470);
and U36507 (N_36507,N_34318,N_31191);
nand U36508 (N_36508,N_32212,N_30978);
nor U36509 (N_36509,N_32837,N_30192);
nand U36510 (N_36510,N_32000,N_30499);
xnor U36511 (N_36511,N_34619,N_34083);
nand U36512 (N_36512,N_33386,N_32901);
and U36513 (N_36513,N_33096,N_31309);
or U36514 (N_36514,N_31894,N_34761);
nor U36515 (N_36515,N_33432,N_32612);
nand U36516 (N_36516,N_31440,N_34869);
nor U36517 (N_36517,N_33272,N_34989);
and U36518 (N_36518,N_34280,N_32155);
or U36519 (N_36519,N_31646,N_33542);
or U36520 (N_36520,N_34451,N_32988);
and U36521 (N_36521,N_30347,N_33162);
xor U36522 (N_36522,N_30946,N_30966);
or U36523 (N_36523,N_32467,N_32037);
nor U36524 (N_36524,N_30118,N_30685);
nand U36525 (N_36525,N_33373,N_33179);
or U36526 (N_36526,N_30233,N_31368);
and U36527 (N_36527,N_34919,N_31002);
and U36528 (N_36528,N_30567,N_32451);
xor U36529 (N_36529,N_30743,N_32915);
nand U36530 (N_36530,N_32570,N_33194);
nand U36531 (N_36531,N_30530,N_30891);
nand U36532 (N_36532,N_32731,N_32851);
and U36533 (N_36533,N_32435,N_31702);
or U36534 (N_36534,N_32501,N_31425);
or U36535 (N_36535,N_30001,N_34990);
and U36536 (N_36536,N_34562,N_32745);
nand U36537 (N_36537,N_30807,N_30143);
nand U36538 (N_36538,N_32359,N_30852);
nor U36539 (N_36539,N_34023,N_31495);
nor U36540 (N_36540,N_34351,N_30767);
nor U36541 (N_36541,N_33646,N_31478);
nor U36542 (N_36542,N_33557,N_32845);
or U36543 (N_36543,N_30629,N_30187);
and U36544 (N_36544,N_33805,N_32357);
nand U36545 (N_36545,N_34586,N_34009);
or U36546 (N_36546,N_32629,N_30478);
xnor U36547 (N_36547,N_34911,N_34741);
nand U36548 (N_36548,N_32684,N_34753);
nor U36549 (N_36549,N_33652,N_34941);
xnor U36550 (N_36550,N_32352,N_31738);
nand U36551 (N_36551,N_32257,N_34918);
nand U36552 (N_36552,N_33297,N_33192);
nor U36553 (N_36553,N_34445,N_34593);
nor U36554 (N_36554,N_31452,N_31995);
or U36555 (N_36555,N_34751,N_33464);
xnor U36556 (N_36556,N_33024,N_34636);
and U36557 (N_36557,N_31968,N_31078);
or U36558 (N_36558,N_30521,N_31428);
and U36559 (N_36559,N_31442,N_32564);
xor U36560 (N_36560,N_34074,N_34790);
xor U36561 (N_36561,N_30220,N_31552);
or U36562 (N_36562,N_33074,N_30215);
nor U36563 (N_36563,N_33798,N_34912);
nand U36564 (N_36564,N_30268,N_30857);
and U36565 (N_36565,N_32011,N_33452);
nor U36566 (N_36566,N_30824,N_32921);
nand U36567 (N_36567,N_31140,N_34025);
or U36568 (N_36568,N_33720,N_34719);
and U36569 (N_36569,N_31973,N_30651);
nand U36570 (N_36570,N_31563,N_30936);
nor U36571 (N_36571,N_30259,N_33121);
nor U36572 (N_36572,N_32596,N_34214);
nand U36573 (N_36573,N_34191,N_30115);
xor U36574 (N_36574,N_31148,N_34597);
or U36575 (N_36575,N_30799,N_34660);
and U36576 (N_36576,N_31214,N_31788);
or U36577 (N_36577,N_33508,N_32267);
and U36578 (N_36578,N_30522,N_31688);
xor U36579 (N_36579,N_33033,N_31529);
nand U36580 (N_36580,N_31130,N_31708);
nor U36581 (N_36581,N_32304,N_31339);
and U36582 (N_36582,N_33268,N_34922);
nand U36583 (N_36583,N_34286,N_34258);
or U36584 (N_36584,N_33016,N_33460);
nor U36585 (N_36585,N_30774,N_31822);
and U36586 (N_36586,N_34946,N_32273);
and U36587 (N_36587,N_33299,N_33067);
or U36588 (N_36588,N_33949,N_30226);
nand U36589 (N_36589,N_30337,N_34209);
nand U36590 (N_36590,N_32873,N_30912);
xnor U36591 (N_36591,N_31297,N_32939);
nor U36592 (N_36592,N_32658,N_34814);
or U36593 (N_36593,N_33153,N_30053);
xnor U36594 (N_36594,N_33294,N_31099);
nand U36595 (N_36595,N_34538,N_31040);
and U36596 (N_36596,N_30376,N_33741);
or U36597 (N_36597,N_32424,N_30183);
nand U36598 (N_36598,N_31391,N_34447);
nor U36599 (N_36599,N_33895,N_31566);
nand U36600 (N_36600,N_34243,N_34041);
nand U36601 (N_36601,N_30312,N_34315);
or U36602 (N_36602,N_32441,N_32434);
nor U36603 (N_36603,N_30624,N_32539);
or U36604 (N_36604,N_31663,N_34558);
nor U36605 (N_36605,N_31864,N_31023);
or U36606 (N_36606,N_34811,N_31896);
and U36607 (N_36607,N_33887,N_32342);
or U36608 (N_36608,N_30040,N_30608);
nand U36609 (N_36609,N_34986,N_33757);
and U36610 (N_36610,N_30395,N_30533);
xnor U36611 (N_36611,N_30667,N_33244);
or U36612 (N_36612,N_33818,N_31001);
nor U36613 (N_36613,N_30981,N_34534);
or U36614 (N_36614,N_30890,N_32566);
and U36615 (N_36615,N_30295,N_32990);
nor U36616 (N_36616,N_30400,N_31733);
nand U36617 (N_36617,N_30438,N_34829);
nor U36618 (N_36618,N_30634,N_33951);
nand U36619 (N_36619,N_34455,N_30368);
nand U36620 (N_36620,N_31241,N_31117);
xor U36621 (N_36621,N_30884,N_31740);
and U36622 (N_36622,N_34662,N_30669);
and U36623 (N_36623,N_32687,N_32240);
nand U36624 (N_36624,N_32960,N_33688);
or U36625 (N_36625,N_30452,N_34818);
and U36626 (N_36626,N_33202,N_34867);
and U36627 (N_36627,N_33614,N_30016);
nand U36628 (N_36628,N_31449,N_32587);
nand U36629 (N_36629,N_30145,N_30696);
or U36630 (N_36630,N_31149,N_30422);
and U36631 (N_36631,N_34910,N_33295);
nor U36632 (N_36632,N_32117,N_32488);
xnor U36633 (N_36633,N_30876,N_31401);
nand U36634 (N_36634,N_30494,N_31709);
and U36635 (N_36635,N_30257,N_33577);
or U36636 (N_36636,N_32309,N_30553);
xnor U36637 (N_36637,N_31877,N_30479);
and U36638 (N_36638,N_31325,N_31279);
xor U36639 (N_36639,N_33072,N_34688);
xnor U36640 (N_36640,N_32189,N_34824);
nor U36641 (N_36641,N_34902,N_32414);
nor U36642 (N_36642,N_32757,N_31883);
nor U36643 (N_36643,N_30569,N_33146);
nor U36644 (N_36644,N_30716,N_30627);
nand U36645 (N_36645,N_34942,N_34788);
and U36646 (N_36646,N_31371,N_30362);
nor U36647 (N_36647,N_31746,N_30338);
and U36648 (N_36648,N_30596,N_30460);
or U36649 (N_36649,N_31056,N_33686);
xor U36650 (N_36650,N_31430,N_34377);
and U36651 (N_36651,N_33499,N_34024);
or U36652 (N_36652,N_33195,N_34551);
or U36653 (N_36653,N_34855,N_31821);
xnor U36654 (N_36654,N_34338,N_34896);
xor U36655 (N_36655,N_33596,N_30812);
xnor U36656 (N_36656,N_30169,N_33549);
and U36657 (N_36657,N_34626,N_34019);
or U36658 (N_36658,N_34758,N_32292);
xnor U36659 (N_36659,N_31198,N_32217);
xnor U36660 (N_36660,N_32940,N_31439);
nand U36661 (N_36661,N_34629,N_33327);
and U36662 (N_36662,N_31510,N_32336);
xor U36663 (N_36663,N_30586,N_34734);
and U36664 (N_36664,N_33367,N_33087);
xnor U36665 (N_36665,N_30098,N_31608);
nor U36666 (N_36666,N_33039,N_33939);
or U36667 (N_36667,N_30165,N_32512);
nor U36668 (N_36668,N_34554,N_34760);
or U36669 (N_36669,N_32186,N_33961);
or U36670 (N_36670,N_34667,N_31659);
and U36671 (N_36671,N_34204,N_33077);
nor U36672 (N_36672,N_31887,N_32438);
nand U36673 (N_36673,N_34746,N_33495);
nand U36674 (N_36674,N_31634,N_32747);
xor U36675 (N_36675,N_30417,N_34602);
nor U36676 (N_36676,N_33058,N_30684);
nor U36677 (N_36677,N_31806,N_30263);
nand U36678 (N_36678,N_31131,N_33573);
xnor U36679 (N_36679,N_31058,N_33281);
nand U36680 (N_36680,N_33382,N_33988);
xor U36681 (N_36681,N_30655,N_34228);
nor U36682 (N_36682,N_30103,N_32891);
and U36683 (N_36683,N_32661,N_33004);
xor U36684 (N_36684,N_31836,N_32801);
nor U36685 (N_36685,N_30027,N_32225);
and U36686 (N_36686,N_34604,N_32063);
or U36687 (N_36687,N_32137,N_31006);
nor U36688 (N_36688,N_33354,N_34645);
or U36689 (N_36689,N_33344,N_32247);
or U36690 (N_36690,N_32296,N_30197);
nand U36691 (N_36691,N_34482,N_30429);
and U36692 (N_36692,N_30465,N_33833);
and U36693 (N_36693,N_33174,N_33755);
and U36694 (N_36694,N_30786,N_34931);
or U36695 (N_36695,N_32054,N_31223);
and U36696 (N_36696,N_33104,N_32878);
and U36697 (N_36697,N_33338,N_34973);
xnor U36698 (N_36698,N_33516,N_30672);
nand U36699 (N_36699,N_30534,N_32325);
or U36700 (N_36700,N_33280,N_32068);
or U36701 (N_36701,N_31436,N_31651);
nand U36702 (N_36702,N_30047,N_34795);
xor U36703 (N_36703,N_33252,N_30265);
or U36704 (N_36704,N_31037,N_31516);
nor U36705 (N_36705,N_30045,N_34807);
nor U36706 (N_36706,N_32881,N_34898);
xor U36707 (N_36707,N_30568,N_32908);
xnor U36708 (N_36708,N_34285,N_30520);
nand U36709 (N_36709,N_34192,N_30637);
xnor U36710 (N_36710,N_34929,N_33869);
or U36711 (N_36711,N_30788,N_30126);
and U36712 (N_36712,N_33780,N_31147);
nor U36713 (N_36713,N_33233,N_30924);
and U36714 (N_36714,N_34221,N_32704);
and U36715 (N_36715,N_33947,N_31231);
xor U36716 (N_36716,N_30805,N_34050);
nand U36717 (N_36717,N_32492,N_34039);
or U36718 (N_36718,N_31810,N_31334);
xor U36719 (N_36719,N_31064,N_31906);
nor U36720 (N_36720,N_33090,N_30348);
or U36721 (N_36721,N_32313,N_30839);
or U36722 (N_36722,N_32968,N_33475);
nand U36723 (N_36723,N_32025,N_31011);
nor U36724 (N_36724,N_30944,N_31912);
and U36725 (N_36725,N_33427,N_30383);
xnor U36726 (N_36726,N_34836,N_30561);
nor U36727 (N_36727,N_32726,N_32645);
and U36728 (N_36728,N_33457,N_32714);
and U36729 (N_36729,N_33670,N_32422);
or U36730 (N_36730,N_30144,N_30605);
nor U36731 (N_36731,N_30132,N_33329);
nand U36732 (N_36732,N_30776,N_30410);
nor U36733 (N_36733,N_33463,N_33437);
and U36734 (N_36734,N_33802,N_31151);
nand U36735 (N_36735,N_32272,N_34273);
and U36736 (N_36736,N_30873,N_31674);
nand U36737 (N_36737,N_32294,N_32316);
and U36738 (N_36738,N_32053,N_31028);
nand U36739 (N_36739,N_33784,N_32528);
xnor U36740 (N_36740,N_34581,N_31308);
nor U36741 (N_36741,N_32010,N_32263);
nand U36742 (N_36742,N_34036,N_34672);
nand U36743 (N_36743,N_31069,N_33875);
xor U36744 (N_36744,N_31515,N_30455);
or U36745 (N_36745,N_30262,N_33014);
and U36746 (N_36746,N_30201,N_32914);
nor U36747 (N_36747,N_34475,N_34971);
xor U36748 (N_36748,N_31112,N_31889);
nand U36749 (N_36749,N_33560,N_33967);
or U36750 (N_36750,N_30415,N_30057);
or U36751 (N_36751,N_32326,N_34373);
nand U36752 (N_36752,N_33606,N_34067);
and U36753 (N_36753,N_32177,N_31919);
nor U36754 (N_36754,N_31407,N_30099);
nand U36755 (N_36755,N_30020,N_33109);
and U36756 (N_36756,N_33201,N_32408);
nand U36757 (N_36757,N_31280,N_33671);
nor U36758 (N_36758,N_32800,N_30968);
nand U36759 (N_36759,N_30836,N_34393);
nor U36760 (N_36760,N_33056,N_31356);
or U36761 (N_36761,N_31670,N_34208);
xor U36762 (N_36762,N_32369,N_34535);
xor U36763 (N_36763,N_34412,N_30633);
and U36764 (N_36764,N_32040,N_31594);
nor U36765 (N_36765,N_32461,N_32254);
and U36766 (N_36766,N_33504,N_32581);
xnor U36767 (N_36767,N_32500,N_34011);
or U36768 (N_36768,N_32923,N_31219);
nor U36769 (N_36769,N_34291,N_30822);
or U36770 (N_36770,N_33105,N_31786);
and U36771 (N_36771,N_34822,N_34690);
and U36772 (N_36772,N_34737,N_31970);
nand U36773 (N_36773,N_33709,N_30639);
nand U36774 (N_36774,N_30389,N_34150);
and U36775 (N_36775,N_32410,N_32974);
and U36776 (N_36776,N_33265,N_32917);
or U36777 (N_36777,N_31630,N_34845);
xor U36778 (N_36778,N_31271,N_33556);
nand U36779 (N_36779,N_34077,N_31207);
nor U36780 (N_36780,N_34655,N_31310);
and U36781 (N_36781,N_31503,N_30764);
or U36782 (N_36782,N_31031,N_34548);
nor U36783 (N_36783,N_34721,N_32129);
xnor U36784 (N_36784,N_31971,N_32601);
nand U36785 (N_36785,N_34363,N_31418);
xor U36786 (N_36786,N_30931,N_34072);
xnor U36787 (N_36787,N_34589,N_30435);
and U36788 (N_36788,N_32383,N_32016);
or U36789 (N_36789,N_32090,N_31681);
nor U36790 (N_36790,N_33043,N_30204);
or U36791 (N_36791,N_31882,N_32977);
and U36792 (N_36792,N_33889,N_30251);
nand U36793 (N_36793,N_34738,N_33188);
nor U36794 (N_36794,N_31647,N_32936);
and U36795 (N_36795,N_32887,N_34862);
and U36796 (N_36796,N_34952,N_30208);
and U36797 (N_36797,N_34643,N_33394);
nor U36798 (N_36798,N_34967,N_32992);
and U36799 (N_36799,N_34975,N_31615);
and U36800 (N_36800,N_31799,N_31532);
nand U36801 (N_36801,N_34138,N_33800);
nand U36802 (N_36802,N_32104,N_32927);
xor U36803 (N_36803,N_30975,N_32858);
and U36804 (N_36804,N_32065,N_32880);
xor U36805 (N_36805,N_30681,N_30997);
and U36806 (N_36806,N_33996,N_34972);
and U36807 (N_36807,N_30125,N_30656);
xor U36808 (N_36808,N_31989,N_34509);
nand U36809 (N_36809,N_30868,N_32568);
and U36810 (N_36810,N_31465,N_33129);
xor U36811 (N_36811,N_31831,N_33081);
nor U36812 (N_36812,N_32896,N_31184);
nor U36813 (N_36813,N_31337,N_31170);
nand U36814 (N_36814,N_30543,N_33176);
and U36815 (N_36815,N_34112,N_32592);
nor U36816 (N_36816,N_32817,N_31662);
or U36817 (N_36817,N_31917,N_33030);
nor U36818 (N_36818,N_34959,N_31692);
or U36819 (N_36819,N_31820,N_31710);
nand U36820 (N_36820,N_33332,N_34767);
nor U36821 (N_36821,N_32312,N_30595);
xnor U36822 (N_36822,N_30071,N_31581);
nor U36823 (N_36823,N_33313,N_34891);
xnor U36824 (N_36824,N_34222,N_32949);
xor U36825 (N_36825,N_32770,N_33415);
or U36826 (N_36826,N_30705,N_31076);
nand U36827 (N_36827,N_33932,N_33449);
xnor U36828 (N_36828,N_30536,N_34485);
xor U36829 (N_36829,N_34980,N_31102);
nand U36830 (N_36830,N_32579,N_34843);
xnor U36831 (N_36831,N_32078,N_34939);
or U36832 (N_36832,N_33570,N_30841);
xnor U36833 (N_36833,N_30707,N_31514);
nand U36834 (N_36834,N_34147,N_31322);
xor U36835 (N_36835,N_31480,N_31453);
or U36836 (N_36836,N_31996,N_34634);
nor U36837 (N_36837,N_34325,N_34132);
nor U36838 (N_36838,N_32283,N_34387);
and U36839 (N_36839,N_32959,N_30333);
xor U36840 (N_36840,N_34927,N_30028);
nand U36841 (N_36841,N_34419,N_31177);
xnor U36842 (N_36842,N_32993,N_31705);
nor U36843 (N_36843,N_32975,N_34493);
and U36844 (N_36844,N_30993,N_34197);
nand U36845 (N_36845,N_33135,N_30630);
nand U36846 (N_36846,N_34563,N_31135);
and U36847 (N_36847,N_33191,N_34637);
or U36848 (N_36848,N_32026,N_32214);
and U36849 (N_36849,N_30930,N_31486);
nand U36850 (N_36850,N_31621,N_31534);
nand U36851 (N_36851,N_33154,N_31306);
or U36852 (N_36852,N_33390,N_32953);
nor U36853 (N_36853,N_33680,N_34283);
or U36854 (N_36854,N_30943,N_34689);
or U36855 (N_36855,N_33019,N_31463);
xnor U36856 (N_36856,N_31915,N_34559);
nand U36857 (N_36857,N_32281,N_33398);
nor U36858 (N_36858,N_30825,N_32245);
or U36859 (N_36859,N_32989,N_33973);
xor U36860 (N_36860,N_34886,N_33979);
nor U36861 (N_36861,N_32459,N_33359);
nor U36862 (N_36862,N_30313,N_30818);
and U36863 (N_36863,N_34571,N_30714);
nand U36864 (N_36864,N_31202,N_33486);
or U36865 (N_36865,N_33284,N_33759);
and U36866 (N_36866,N_33732,N_33881);
nand U36867 (N_36867,N_30014,N_31121);
or U36868 (N_36868,N_32902,N_31496);
nand U36869 (N_36869,N_33602,N_30869);
or U36870 (N_36870,N_33539,N_34491);
nand U36871 (N_36871,N_32205,N_33242);
and U36872 (N_36872,N_34414,N_33258);
xor U36873 (N_36873,N_30369,N_32712);
nor U36874 (N_36874,N_34422,N_33807);
nor U36875 (N_36875,N_34628,N_32381);
nor U36876 (N_36876,N_34865,N_34206);
nor U36877 (N_36877,N_33036,N_32746);
nand U36878 (N_36878,N_30640,N_30081);
nand U36879 (N_36879,N_33523,N_30902);
or U36880 (N_36880,N_31071,N_33586);
nand U36881 (N_36881,N_32450,N_31678);
nand U36882 (N_36882,N_33536,N_32171);
nand U36883 (N_36883,N_30089,N_30358);
nand U36884 (N_36884,N_32957,N_31400);
xnor U36885 (N_36885,N_34556,N_33790);
or U36886 (N_36886,N_33565,N_31125);
nor U36887 (N_36887,N_33867,N_32716);
xnor U36888 (N_36888,N_32643,N_32475);
or U36889 (N_36889,N_33420,N_32828);
or U36890 (N_36890,N_31598,N_33860);
or U36891 (N_36891,N_34429,N_31127);
nand U36892 (N_36892,N_31403,N_34893);
or U36893 (N_36893,N_30547,N_34063);
and U36894 (N_36894,N_31727,N_34257);
nand U36895 (N_36895,N_32680,N_31481);
nor U36896 (N_36896,N_30738,N_34608);
or U36897 (N_36897,N_31972,N_33885);
and U36898 (N_36898,N_32985,N_31606);
nand U36899 (N_36899,N_32495,N_33788);
xor U36900 (N_36900,N_30587,N_30059);
or U36901 (N_36901,N_34697,N_34853);
or U36902 (N_36902,N_34238,N_33835);
and U36903 (N_36903,N_32491,N_33647);
or U36904 (N_36904,N_31590,N_32167);
or U36905 (N_36905,N_32678,N_33926);
nand U36906 (N_36906,N_31132,N_33257);
nor U36907 (N_36907,N_32697,N_31328);
and U36908 (N_36908,N_31139,N_33326);
nand U36909 (N_36909,N_32306,N_32200);
or U36910 (N_36910,N_32511,N_33792);
nand U36911 (N_36911,N_31269,N_31171);
xor U36912 (N_36912,N_33273,N_34055);
or U36913 (N_36913,N_30005,N_32518);
nand U36914 (N_36914,N_32899,N_32384);
xor U36915 (N_36915,N_34771,N_31229);
nand U36916 (N_36916,N_34866,N_31275);
xor U36917 (N_36917,N_32798,N_31426);
or U36918 (N_36918,N_32893,N_33009);
nor U36919 (N_36919,N_33674,N_31573);
nor U36920 (N_36920,N_33904,N_32682);
xor U36921 (N_36921,N_31227,N_31982);
or U36922 (N_36922,N_31868,N_33227);
nor U36923 (N_36923,N_30211,N_34970);
nor U36924 (N_36924,N_32513,N_30664);
xnor U36925 (N_36925,N_31179,N_33898);
or U36926 (N_36926,N_33046,N_33161);
xnor U36927 (N_36927,N_31387,N_34306);
nand U36928 (N_36928,N_32082,N_33813);
or U36929 (N_36929,N_32335,N_30795);
nor U36930 (N_36930,N_34350,N_32648);
or U36931 (N_36931,N_33527,N_33601);
nand U36932 (N_36932,N_31192,N_32688);
nor U36933 (N_36933,N_30423,N_33718);
nand U36934 (N_36934,N_33288,N_32722);
and U36935 (N_36935,N_31551,N_30198);
nor U36936 (N_36936,N_31016,N_33628);
xnor U36937 (N_36937,N_33578,N_31977);
nand U36938 (N_36938,N_31902,N_30349);
xnor U36939 (N_36939,N_32786,N_31772);
and U36940 (N_36940,N_30128,N_31210);
or U36941 (N_36941,N_33350,N_32606);
xor U36942 (N_36942,N_32327,N_31948);
and U36943 (N_36943,N_32266,N_31018);
xor U36944 (N_36944,N_32667,N_34054);
nor U36945 (N_36945,N_31499,N_31832);
nand U36946 (N_36946,N_32979,N_32108);
or U36947 (N_36947,N_33500,N_31008);
and U36948 (N_36948,N_30775,N_33552);
nor U36949 (N_36949,N_31021,N_33466);
nand U36950 (N_36950,N_31421,N_34299);
nor U36951 (N_36951,N_30951,N_32042);
xor U36952 (N_36952,N_32637,N_32260);
nor U36953 (N_36953,N_31350,N_33517);
xnor U36954 (N_36954,N_34887,N_33330);
nor U36955 (N_36955,N_33168,N_33547);
or U36956 (N_36956,N_30649,N_31803);
nand U36957 (N_36957,N_32586,N_32361);
or U36958 (N_36958,N_32708,N_30962);
or U36959 (N_36959,N_32106,N_32825);
nand U36960 (N_36960,N_31494,N_32790);
and U36961 (N_36961,N_31910,N_30070);
nor U36962 (N_36962,N_31196,N_32395);
and U36963 (N_36963,N_31981,N_30662);
nand U36964 (N_36964,N_30761,N_33409);
and U36965 (N_36965,N_32056,N_33762);
and U36966 (N_36966,N_34240,N_30340);
nor U36967 (N_36967,N_32298,N_34463);
nand U36968 (N_36968,N_32854,N_31133);
and U36969 (N_36969,N_32859,N_33035);
nand U36970 (N_36970,N_33569,N_30948);
nand U36971 (N_36971,N_32950,N_30592);
nor U36972 (N_36972,N_31741,N_30504);
or U36973 (N_36973,N_33110,N_31991);
or U36974 (N_36974,N_31675,N_32346);
and U36975 (N_36975,N_31364,N_34465);
nor U36976 (N_36976,N_34681,N_31538);
xor U36977 (N_36977,N_33436,N_33223);
nand U36978 (N_36978,N_34799,N_32810);
nor U36979 (N_36979,N_33701,N_32826);
nand U36980 (N_36980,N_32578,N_33687);
nand U36981 (N_36981,N_33713,N_34685);
xor U36982 (N_36982,N_31385,N_32730);
xor U36983 (N_36983,N_33721,N_34335);
nand U36984 (N_36984,N_30599,N_31946);
nand U36985 (N_36985,N_31652,N_32220);
and U36986 (N_36986,N_34189,N_33985);
xor U36987 (N_36987,N_30699,N_31564);
and U36988 (N_36988,N_31042,N_32675);
xor U36989 (N_36989,N_32799,N_33306);
xor U36990 (N_36990,N_33189,N_34028);
xor U36991 (N_36991,N_33193,N_30588);
nor U36992 (N_36992,N_30804,N_30332);
and U36993 (N_36993,N_32035,N_34319);
nor U36994 (N_36994,N_33397,N_34776);
nand U36995 (N_36995,N_32670,N_33362);
nand U36996 (N_36996,N_32020,N_30305);
and U36997 (N_36997,N_34329,N_30476);
xnor U36998 (N_36998,N_31999,N_34017);
nand U36999 (N_36999,N_34403,N_31920);
or U37000 (N_37000,N_31804,N_30661);
nand U37001 (N_37001,N_30123,N_33203);
xor U37002 (N_37002,N_30794,N_33235);
nor U37003 (N_37003,N_32945,N_30351);
or U37004 (N_37004,N_30519,N_32971);
nand U37005 (N_37005,N_31396,N_32605);
and U37006 (N_37006,N_33151,N_33048);
nor U37007 (N_37007,N_30939,N_32864);
nor U37008 (N_37008,N_31556,N_30110);
nor U37009 (N_37009,N_33334,N_34481);
nand U37010 (N_37010,N_31588,N_33037);
and U37011 (N_37011,N_30391,N_30064);
nor U37012 (N_37012,N_34590,N_31617);
or U37013 (N_37013,N_31794,N_32954);
or U37014 (N_37014,N_33656,N_31450);
xor U37015 (N_37015,N_33531,N_34396);
xor U37016 (N_37016,N_33286,N_31520);
xor U37017 (N_37017,N_32652,N_34720);
and U37018 (N_37018,N_33458,N_30844);
or U37019 (N_37019,N_30120,N_32417);
nor U37020 (N_37020,N_32073,N_32926);
or U37021 (N_37021,N_30316,N_33589);
nor U37022 (N_37022,N_32164,N_30427);
xnor U37023 (N_37023,N_32047,N_30856);
xnor U37024 (N_37024,N_31980,N_31158);
xor U37025 (N_37025,N_33673,N_33669);
nor U37026 (N_37026,N_33417,N_30827);
or U37027 (N_37027,N_31134,N_34487);
nor U37028 (N_37028,N_30579,N_31787);
xnor U37029 (N_37029,N_34765,N_33831);
xnor U37030 (N_37030,N_33846,N_30861);
or U37031 (N_37031,N_30292,N_32075);
and U37032 (N_37032,N_31597,N_34575);
and U37033 (N_37033,N_33777,N_30816);
nor U37034 (N_37034,N_30644,N_32741);
nor U37035 (N_37035,N_32705,N_31380);
nor U37036 (N_37036,N_32980,N_31370);
or U37037 (N_37037,N_32522,N_32310);
and U37038 (N_37038,N_32636,N_34013);
nor U37039 (N_37039,N_34109,N_32841);
xnor U37040 (N_37040,N_31094,N_33719);
nor U37041 (N_37041,N_32329,N_32095);
and U37042 (N_37042,N_32375,N_32030);
and U37043 (N_37043,N_34565,N_31964);
nor U37044 (N_37044,N_30763,N_30710);
and U37045 (N_37045,N_31290,N_30712);
nand U37046 (N_37046,N_34539,N_30406);
or U37047 (N_37047,N_32642,N_32228);
or U37048 (N_37048,N_30436,N_34057);
xor U37049 (N_37049,N_32749,N_30424);
nand U37050 (N_37050,N_30329,N_34926);
xor U37051 (N_37051,N_34675,N_34018);
or U37052 (N_37052,N_31664,N_32163);
or U37053 (N_37053,N_32819,N_34407);
or U37054 (N_37054,N_31619,N_30659);
nor U37055 (N_37055,N_31600,N_33311);
nand U37056 (N_37056,N_34731,N_33551);
or U37057 (N_37057,N_34907,N_31186);
or U37058 (N_37058,N_32816,N_30591);
or U37059 (N_37059,N_34603,N_32834);
nor U37060 (N_37060,N_31828,N_33312);
and U37061 (N_37061,N_33465,N_30954);
or U37062 (N_37062,N_31921,N_31488);
nand U37063 (N_37063,N_32367,N_32598);
or U37064 (N_37064,N_33488,N_32347);
xor U37065 (N_37065,N_31009,N_32894);
nand U37066 (N_37066,N_33073,N_31749);
nand U37067 (N_37067,N_30361,N_33322);
nor U37068 (N_37068,N_33634,N_31892);
nand U37069 (N_37069,N_32388,N_32839);
nor U37070 (N_37070,N_32079,N_34585);
and U37071 (N_37071,N_30148,N_31650);
nor U37072 (N_37072,N_33116,N_30287);
nand U37073 (N_37073,N_30758,N_33580);
nand U37074 (N_37074,N_30136,N_34934);
nor U37075 (N_37075,N_33361,N_32720);
nand U37076 (N_37076,N_34148,N_30573);
and U37077 (N_37077,N_33643,N_32145);
nand U37078 (N_37078,N_34519,N_33983);
nor U37079 (N_37079,N_30119,N_33651);
nor U37080 (N_37080,N_32778,N_32088);
nor U37081 (N_37081,N_30709,N_33027);
or U37082 (N_37082,N_31947,N_31540);
nand U37083 (N_37083,N_32630,N_30751);
xor U37084 (N_37084,N_34453,N_32333);
nor U37085 (N_37085,N_34712,N_34215);
nand U37086 (N_37086,N_34995,N_32259);
xor U37087 (N_37087,N_33786,N_32221);
or U37088 (N_37088,N_33582,N_32571);
and U37089 (N_37089,N_30256,N_31162);
or U37090 (N_37090,N_34423,N_32848);
or U37091 (N_37091,N_34182,N_30051);
nor U37092 (N_37092,N_33356,N_30548);
nor U37093 (N_37093,N_31091,N_33305);
and U37094 (N_37094,N_33377,N_30736);
nor U37095 (N_37095,N_30511,N_34260);
nor U37096 (N_37096,N_31054,N_32657);
nand U37097 (N_37097,N_34128,N_34908);
nor U37098 (N_37098,N_34120,N_34744);
xnor U37099 (N_37099,N_32238,N_32633);
nand U37100 (N_37100,N_31722,N_33114);
nand U37101 (N_37101,N_32009,N_32018);
nor U37102 (N_37102,N_34728,N_31276);
and U37103 (N_37103,N_30490,N_34644);
and U37104 (N_37104,N_34678,N_33729);
and U37105 (N_37105,N_32470,N_33134);
nor U37106 (N_37106,N_30102,N_30468);
xnor U37107 (N_37107,N_31533,N_34717);
xor U37108 (N_37108,N_32906,N_31346);
and U37109 (N_37109,N_32557,N_33567);
xnor U37110 (N_37110,N_30108,N_31323);
nand U37111 (N_37111,N_30965,N_31870);
nor U37112 (N_37112,N_34071,N_31699);
nand U37113 (N_37113,N_33906,N_30570);
nand U37114 (N_37114,N_33379,N_30107);
or U37115 (N_37115,N_33062,N_32023);
nor U37116 (N_37116,N_34200,N_30290);
and U37117 (N_37117,N_30088,N_30382);
nand U37118 (N_37118,N_31805,N_30162);
nand U37119 (N_37119,N_34808,N_32334);
nor U37120 (N_37120,N_32618,N_32622);
and U37121 (N_37121,N_30181,N_30535);
or U37122 (N_37122,N_32694,N_32489);
or U37123 (N_37123,N_34467,N_32349);
nor U37124 (N_37124,N_34125,N_31359);
and U37125 (N_37125,N_33989,N_33482);
xnor U37126 (N_37126,N_34440,N_30657);
and U37127 (N_37127,N_32168,N_30513);
nand U37128 (N_37128,N_33568,N_31105);
or U37129 (N_37129,N_34127,N_32928);
and U37130 (N_37130,N_31092,N_32809);
and U37131 (N_37131,N_34096,N_32840);
xnor U37132 (N_37132,N_30747,N_32374);
xnor U37133 (N_37133,N_32255,N_32067);
or U37134 (N_37134,N_33218,N_31798);
xor U37135 (N_37135,N_31518,N_33828);
nand U37136 (N_37136,N_31677,N_32087);
or U37137 (N_37137,N_34410,N_33521);
nand U37138 (N_37138,N_34183,N_34292);
and U37139 (N_37139,N_33519,N_33797);
and U37140 (N_37140,N_33844,N_33021);
nor U37141 (N_37141,N_33171,N_31281);
and U37142 (N_37142,N_34504,N_31950);
and U37143 (N_37143,N_31349,N_33791);
xor U37144 (N_37144,N_31969,N_30345);
nor U37145 (N_37145,N_33387,N_33407);
or U37146 (N_37146,N_32086,N_30815);
xor U37147 (N_37147,N_34269,N_32820);
xor U37148 (N_37148,N_34653,N_30642);
and U37149 (N_37149,N_30754,N_34404);
xor U37150 (N_37150,N_31585,N_31393);
nand U37151 (N_37151,N_30303,N_31793);
or U37152 (N_37152,N_31475,N_30531);
and U37153 (N_37153,N_31104,N_31111);
or U37154 (N_37154,N_34357,N_33138);
and U37155 (N_37155,N_34439,N_31505);
or U37156 (N_37156,N_33370,N_32013);
or U37157 (N_37157,N_30853,N_31846);
nor U37158 (N_37158,N_32156,N_33034);
or U37159 (N_37159,N_34131,N_33108);
nand U37160 (N_37160,N_33984,N_31265);
xor U37161 (N_37161,N_34398,N_33308);
nor U37162 (N_37162,N_32320,N_33910);
nand U37163 (N_37163,N_34498,N_32999);
nand U37164 (N_37164,N_30354,N_32797);
nor U37165 (N_37165,N_30956,N_31263);
nor U37166 (N_37166,N_30252,N_30300);
nor U37167 (N_37167,N_31344,N_31935);
xor U37168 (N_37168,N_32350,N_31856);
nand U37169 (N_37169,N_30645,N_33182);
or U37170 (N_37170,N_33975,N_30528);
xnor U37171 (N_37171,N_34408,N_34630);
or U37172 (N_37172,N_31445,N_33851);
nor U37173 (N_37173,N_34437,N_33403);
nand U37174 (N_37174,N_31246,N_32447);
or U37175 (N_37175,N_34380,N_32452);
nand U37176 (N_37176,N_30146,N_32588);
and U37177 (N_37177,N_34160,N_32062);
xnor U37178 (N_37178,N_31622,N_30458);
nand U37179 (N_37179,N_31546,N_32373);
and U37180 (N_37180,N_30280,N_30750);
or U37181 (N_37181,N_30848,N_34541);
xnor U37182 (N_37182,N_30858,N_32394);
xor U37183 (N_37183,N_33689,N_31624);
nand U37184 (N_37184,N_32973,N_31419);
or U37185 (N_37185,N_31687,N_30987);
and U37186 (N_37186,N_31706,N_33937);
and U37187 (N_37187,N_31433,N_31930);
and U37188 (N_37188,N_30846,N_33896);
nand U37189 (N_37189,N_31108,N_30058);
or U37190 (N_37190,N_30325,N_30611);
nand U37191 (N_37191,N_34857,N_31206);
and U37192 (N_37192,N_32911,N_33395);
xnor U37193 (N_37193,N_32472,N_33870);
nor U37194 (N_37194,N_31234,N_31953);
nand U37195 (N_37195,N_30532,N_33740);
and U37196 (N_37196,N_34988,N_33310);
and U37197 (N_37197,N_33742,N_32780);
nor U37198 (N_37198,N_32232,N_32655);
and U37199 (N_37199,N_32322,N_33864);
and U37200 (N_37200,N_34879,N_32442);
nand U37201 (N_37201,N_31174,N_31978);
or U37202 (N_37202,N_33921,N_34623);
nand U37203 (N_37203,N_31808,N_34780);
nand U37204 (N_37204,N_30061,N_32721);
and U37205 (N_37205,N_34592,N_33588);
and U37206 (N_37206,N_33320,N_30412);
nor U37207 (N_37207,N_31616,N_34895);
or U37208 (N_37208,N_34388,N_33809);
nand U37209 (N_37209,N_33733,N_32354);
xor U37210 (N_37210,N_31471,N_32976);
nand U37211 (N_37211,N_34572,N_30728);
xor U37212 (N_37212,N_34413,N_30769);
nand U37213 (N_37213,N_34220,N_32805);
nor U37214 (N_37214,N_33913,N_32558);
nand U37215 (N_37215,N_33490,N_31296);
or U37216 (N_37216,N_33540,N_32665);
or U37217 (N_37217,N_31901,N_34099);
or U37218 (N_37218,N_34876,N_32431);
nand U37219 (N_37219,N_31165,N_32609);
nor U37220 (N_37220,N_34654,N_33345);
nor U37221 (N_37221,N_32521,N_31840);
or U37222 (N_37222,N_32689,N_34223);
nand U37223 (N_37223,N_30679,N_33131);
xnor U37224 (N_37224,N_34582,N_32432);
nand U37225 (N_37225,N_33180,N_34037);
nor U37226 (N_37226,N_32036,N_31928);
xor U37227 (N_37227,N_31643,N_32590);
xnor U37228 (N_37228,N_30899,N_32552);
xor U37229 (N_37229,N_34464,N_34042);
nand U37230 (N_37230,N_31700,N_33111);
and U37231 (N_37231,N_34930,N_34105);
nor U37232 (N_37232,N_34599,N_33663);
or U37233 (N_37233,N_33435,N_31255);
and U37234 (N_37234,N_31723,N_33918);
nand U37235 (N_37235,N_31604,N_30472);
or U37236 (N_37236,N_32525,N_32529);
xor U37237 (N_37237,N_31232,N_31511);
xnor U37238 (N_37238,N_30506,N_34840);
and U37239 (N_37239,N_33758,N_30467);
nand U37240 (N_37240,N_32471,N_32299);
nor U37241 (N_37241,N_32262,N_31633);
or U37242 (N_37242,N_33585,N_30038);
and U37243 (N_37243,N_30006,N_33260);
and U37244 (N_37244,N_33316,N_31807);
xnor U37245 (N_37245,N_30285,N_31682);
xor U37246 (N_37246,N_30381,N_31578);
xor U37247 (N_37247,N_31742,N_33011);
xor U37248 (N_37248,N_31506,N_32331);
or U37249 (N_37249,N_33605,N_31013);
xnor U37250 (N_37250,N_34322,N_34118);
and U37251 (N_37251,N_30508,N_30913);
and U37252 (N_37252,N_31367,N_34450);
nand U37253 (N_37253,N_30678,N_30603);
and U37254 (N_37254,N_34993,N_33968);
xnor U37255 (N_37255,N_34656,N_33794);
nor U37256 (N_37256,N_30752,N_32548);
nor U37257 (N_37257,N_30326,N_31907);
nand U37258 (N_37258,N_33360,N_33028);
xor U37259 (N_37259,N_33505,N_30063);
xor U37260 (N_37260,N_34366,N_34932);
xnor U37261 (N_37261,N_30870,N_31498);
xnor U37262 (N_37262,N_30748,N_30582);
or U37263 (N_37263,N_31770,N_33147);
xnor U37264 (N_37264,N_33933,N_30668);
nor U37265 (N_37265,N_33285,N_32222);
or U37266 (N_37266,N_31763,N_34486);
nor U37267 (N_37267,N_32783,N_33052);
nor U37268 (N_37268,N_30482,N_31333);
xor U37269 (N_37269,N_34133,N_30004);
nand U37270 (N_37270,N_34330,N_31729);
and U37271 (N_37271,N_32573,N_34871);
xor U37272 (N_37272,N_32946,N_31175);
and U37273 (N_37273,N_31109,N_34103);
and U37274 (N_37274,N_31114,N_30900);
nor U37275 (N_37275,N_32332,N_33957);
nor U37276 (N_37276,N_34266,N_31164);
nand U37277 (N_37277,N_34472,N_32478);
nand U37278 (N_37278,N_32765,N_31609);
nand U37279 (N_37279,N_33434,N_32860);
xnor U37280 (N_37280,N_33055,N_30688);
xnor U37281 (N_37281,N_30613,N_30264);
and U37282 (N_37282,N_33017,N_32041);
or U37283 (N_37283,N_33439,N_32290);
and U37284 (N_37284,N_30580,N_32948);
nand U37285 (N_37285,N_34657,N_30142);
nor U37286 (N_37286,N_31291,N_32130);
or U37287 (N_37287,N_32399,N_32345);
nor U37288 (N_37288,N_33745,N_31694);
xnor U37289 (N_37289,N_32201,N_34860);
nor U37290 (N_37290,N_34564,N_33764);
nand U37291 (N_37291,N_30837,N_32759);
xor U37292 (N_37292,N_34364,N_31876);
nor U37293 (N_37293,N_33158,N_31562);
and U37294 (N_37294,N_34287,N_32610);
or U37295 (N_37295,N_32115,N_34084);
or U37296 (N_37296,N_31404,N_31640);
nor U37297 (N_37297,N_34173,N_32242);
and U37298 (N_37298,N_30399,N_34664);
nor U37299 (N_37299,N_32433,N_30141);
nor U37300 (N_37300,N_34854,N_33357);
and U37301 (N_37301,N_31724,N_31048);
xor U37302 (N_37302,N_32084,N_33358);
xnor U37303 (N_37303,N_30990,N_32617);
nand U37304 (N_37304,N_32446,N_30832);
xnor U37305 (N_37305,N_31122,N_30493);
and U37306 (N_37306,N_30127,N_34008);
xor U37307 (N_37307,N_30935,N_32761);
xor U37308 (N_37308,N_31945,N_30941);
xor U37309 (N_37309,N_30232,N_31332);
nor U37310 (N_37310,N_32517,N_33217);
and U37311 (N_37311,N_33645,N_33859);
xor U37312 (N_37312,N_34748,N_31152);
xor U37313 (N_37313,N_33704,N_30133);
nor U37314 (N_37314,N_30239,N_31607);
nand U37315 (N_37315,N_30722,N_34916);
xnor U37316 (N_37316,N_34341,N_32691);
or U37317 (N_37317,N_32302,N_31560);
and U37318 (N_37318,N_33502,N_30791);
nor U37319 (N_37319,N_32057,N_34928);
and U37320 (N_37320,N_33879,N_33838);
nor U37321 (N_37321,N_31288,N_33679);
nor U37322 (N_37322,N_34115,N_32843);
xor U37323 (N_37323,N_34792,N_30572);
and U37324 (N_37324,N_34803,N_33102);
nand U37325 (N_37325,N_33467,N_30885);
or U37326 (N_37326,N_32582,N_32193);
nand U37327 (N_37327,N_32502,N_31172);
and U37328 (N_37328,N_31335,N_33137);
xor U37329 (N_37329,N_32183,N_34370);
or U37330 (N_37330,N_30149,N_32001);
nor U37331 (N_37331,N_30134,N_31208);
and U37332 (N_37332,N_30483,N_32781);
or U37333 (N_37333,N_30386,N_33848);
and U37334 (N_37334,N_31209,N_31249);
xor U37335 (N_37335,N_32935,N_34169);
nand U37336 (N_37336,N_30116,N_32427);
nor U37337 (N_37337,N_34003,N_34669);
and U37338 (N_37338,N_31331,N_33478);
or U37339 (N_37339,N_34374,N_31627);
and U37340 (N_37340,N_34718,N_33441);
nand U37341 (N_37341,N_30625,N_31473);
nor U37342 (N_37342,N_30919,N_30609);
or U37343 (N_37343,N_30293,N_33857);
or U37344 (N_37344,N_32411,N_31077);
nor U37345 (N_37345,N_31582,N_32756);
nor U37346 (N_37346,N_32158,N_30277);
nor U37347 (N_37347,N_34894,N_31343);
and U37348 (N_37348,N_30447,N_33481);
nor U37349 (N_37349,N_34512,N_34245);
or U37350 (N_37350,N_34668,N_34670);
or U37351 (N_37351,N_34356,N_30394);
nand U37352 (N_37352,N_32197,N_31110);
nand U37353 (N_37353,N_31587,N_33381);
or U37354 (N_37354,N_30730,N_31791);
xnor U37355 (N_37355,N_31161,N_31554);
or U37356 (N_37356,N_30538,N_31967);
nand U37357 (N_37357,N_34652,N_30397);
or U37358 (N_37358,N_31317,N_33919);
nand U37359 (N_37359,N_31167,N_32014);
nand U37360 (N_37360,N_33627,N_34253);
and U37361 (N_37361,N_32576,N_31047);
nand U37362 (N_37362,N_33164,N_31941);
and U37363 (N_37363,N_34310,N_30160);
and U37364 (N_37364,N_31397,N_33274);
nor U37365 (N_37365,N_33884,N_32083);
or U37366 (N_37366,N_34261,N_33871);
and U37367 (N_37367,N_33812,N_34740);
or U37368 (N_37368,N_33139,N_33365);
xnor U37369 (N_37369,N_32774,N_34627);
or U37370 (N_37370,N_30928,N_30894);
nor U37371 (N_37371,N_33406,N_30079);
xnor U37372 (N_37372,N_33212,N_31698);
nor U37373 (N_37373,N_33001,N_33822);
and U37374 (N_37374,N_31432,N_32621);
and U37375 (N_37375,N_34944,N_31974);
nor U37376 (N_37376,N_31468,N_30114);
and U37377 (N_37377,N_30517,N_32782);
or U37378 (N_37378,N_33209,N_34938);
xnor U37379 (N_37379,N_33609,N_34828);
xor U37380 (N_37380,N_31926,N_34680);
nor U37381 (N_37381,N_30984,N_33703);
and U37382 (N_37382,N_33510,N_30646);
or U37383 (N_37383,N_31295,N_33501);
or U37384 (N_37384,N_34635,N_31363);
nand U37385 (N_37385,N_34837,N_34817);
xnor U37386 (N_37386,N_30104,N_30245);
or U37387 (N_37387,N_31844,N_32532);
and U37388 (N_37388,N_33756,N_31728);
or U37389 (N_37389,N_33773,N_33865);
xor U37390 (N_37390,N_32210,N_34892);
or U37391 (N_37391,N_32868,N_30294);
xor U37392 (N_37392,N_34961,N_31669);
nor U37393 (N_37393,N_32967,N_34060);
xor U37394 (N_37394,N_34480,N_31282);
or U37395 (N_37395,N_30523,N_32170);
nand U37396 (N_37396,N_33241,N_33366);
nand U37397 (N_37397,N_32739,N_31041);
or U37398 (N_37398,N_30177,N_32879);
or U37399 (N_37399,N_31490,N_30560);
xnor U37400 (N_37400,N_30212,N_33384);
nand U37401 (N_37401,N_31613,N_30620);
and U37402 (N_37402,N_30826,N_30327);
and U37403 (N_37403,N_30744,N_31559);
and U37404 (N_37404,N_33292,N_30253);
xor U37405 (N_37405,N_34825,N_33775);
and U37406 (N_37406,N_31879,N_32372);
nor U37407 (N_37407,N_34700,N_32849);
xor U37408 (N_37408,N_32802,N_31922);
xnor U37409 (N_37409,N_31923,N_30275);
or U37410 (N_37410,N_34754,N_31431);
and U37411 (N_37411,N_32397,N_30067);
nor U37412 (N_37412,N_34768,N_34607);
or U37413 (N_37413,N_34460,N_33472);
or U37414 (N_37414,N_34353,N_34411);
xor U37415 (N_37415,N_33393,N_31933);
nor U37416 (N_37416,N_34671,N_31392);
nand U37417 (N_37417,N_30150,N_34588);
nor U37418 (N_37418,N_34736,N_34528);
nor U37419 (N_37419,N_30723,N_34994);
nor U37420 (N_37420,N_30654,N_34614);
or U37421 (N_37421,N_32445,N_30917);
nor U37422 (N_37422,N_30155,N_33843);
nor U37423 (N_37423,N_32413,N_32743);
and U37424 (N_37424,N_31435,N_32912);
nand U37425 (N_37425,N_32278,N_30271);
and U37426 (N_37426,N_32784,N_31266);
or U37427 (N_37427,N_33636,N_33868);
nand U37428 (N_37428,N_32448,N_32624);
or U37429 (N_37429,N_34239,N_32535);
nor U37430 (N_37430,N_32207,N_31277);
xnor U37431 (N_37431,N_31867,N_30584);
or U37432 (N_37432,N_30213,N_31377);
xnor U37433 (N_37433,N_30270,N_30121);
nor U37434 (N_37434,N_32389,N_30872);
and U37435 (N_37435,N_30515,N_32135);
or U37436 (N_37436,N_34649,N_31085);
nand U37437 (N_37437,N_33470,N_31653);
or U37438 (N_37438,N_34835,N_34265);
nor U37439 (N_37439,N_33172,N_30216);
nor U37440 (N_37440,N_32080,N_30176);
or U37441 (N_37441,N_31599,N_31561);
nor U37442 (N_37442,N_34343,N_32561);
nor U37443 (N_37443,N_34334,N_34166);
or U37444 (N_37444,N_32118,N_31362);
nor U37445 (N_37445,N_33684,N_32544);
nor U37446 (N_37446,N_34732,N_34530);
or U37447 (N_37447,N_33190,N_30731);
nor U37448 (N_37448,N_33015,N_32285);
and U37449 (N_37449,N_32303,N_34726);
nor U37450 (N_37450,N_32045,N_33587);
or U37451 (N_37451,N_33405,N_34606);
nand U37452 (N_37452,N_34770,N_32174);
nor U37453 (N_37453,N_34106,N_30597);
nor U37454 (N_37454,N_34641,N_32872);
nor U37455 (N_37455,N_33494,N_34001);
and U37456 (N_37456,N_33659,N_33293);
xnor U37457 (N_37457,N_31683,N_31987);
and U37458 (N_37458,N_32551,N_31100);
xnor U37459 (N_37459,N_33430,N_33210);
or U37460 (N_37460,N_32604,N_32795);
nor U37461 (N_37461,N_30727,N_31755);
nor U37462 (N_37462,N_31340,N_33416);
xnor U37463 (N_37463,N_30357,N_33375);
nor U37464 (N_37464,N_32662,N_30636);
xor U37465 (N_37465,N_34251,N_31324);
or U37466 (N_37466,N_31988,N_30881);
or U37467 (N_37467,N_34107,N_31591);
or U37468 (N_37468,N_34154,N_30892);
nor U37469 (N_37469,N_34309,N_31050);
and U37470 (N_37470,N_32635,N_32769);
nor U37471 (N_37471,N_32102,N_30012);
or U37472 (N_37472,N_30898,N_32646);
nor U37473 (N_37473,N_30817,N_33045);
nand U37474 (N_37474,N_31686,N_30835);
or U37475 (N_37475,N_30952,N_31301);
nor U37476 (N_37476,N_34059,N_32111);
xor U37477 (N_37477,N_31589,N_34687);
and U37478 (N_37478,N_34294,N_30244);
or U37479 (N_37479,N_34270,N_32698);
nand U37480 (N_37480,N_34937,N_32224);
nor U37481 (N_37481,N_33548,N_32236);
or U37482 (N_37482,N_30432,N_33769);
or U37483 (N_37483,N_34418,N_32580);
xor U37484 (N_37484,N_34159,N_33845);
xor U37485 (N_37485,N_33905,N_34577);
or U37486 (N_37486,N_34080,N_32019);
and U37487 (N_37487,N_31081,N_31736);
and U37488 (N_37488,N_33336,N_32766);
or U37489 (N_37489,N_31519,N_34587);
or U37490 (N_37490,N_31022,N_30416);
nand U37491 (N_37491,N_30471,N_32885);
nand U37492 (N_37492,N_34044,N_33378);
and U37493 (N_37493,N_30529,N_32363);
nor U37494 (N_37494,N_31046,N_30195);
xor U37495 (N_37495,N_32454,N_32150);
nand U37496 (N_37496,N_32152,N_31062);
nand U37497 (N_37497,N_30379,N_31113);
nand U37498 (N_37498,N_30725,N_34295);
nor U37499 (N_37499,N_30854,N_31366);
or U37500 (N_37500,N_34215,N_32845);
nand U37501 (N_37501,N_34385,N_32063);
and U37502 (N_37502,N_31186,N_32622);
and U37503 (N_37503,N_33987,N_34639);
nand U37504 (N_37504,N_31399,N_33964);
and U37505 (N_37505,N_34658,N_33175);
xor U37506 (N_37506,N_34285,N_30091);
or U37507 (N_37507,N_30945,N_33864);
nand U37508 (N_37508,N_32748,N_33562);
nand U37509 (N_37509,N_31181,N_33755);
and U37510 (N_37510,N_30170,N_32166);
xnor U37511 (N_37511,N_32125,N_30635);
nor U37512 (N_37512,N_34281,N_31345);
and U37513 (N_37513,N_34547,N_31939);
nor U37514 (N_37514,N_32061,N_32949);
xnor U37515 (N_37515,N_32113,N_30720);
nand U37516 (N_37516,N_32572,N_33071);
nand U37517 (N_37517,N_31833,N_30906);
or U37518 (N_37518,N_31233,N_32184);
nand U37519 (N_37519,N_31879,N_30652);
xnor U37520 (N_37520,N_32589,N_31518);
nand U37521 (N_37521,N_32404,N_33057);
nand U37522 (N_37522,N_31599,N_33163);
and U37523 (N_37523,N_31051,N_33012);
or U37524 (N_37524,N_31451,N_33590);
or U37525 (N_37525,N_33644,N_33044);
xor U37526 (N_37526,N_34246,N_30321);
xor U37527 (N_37527,N_33974,N_34898);
and U37528 (N_37528,N_34655,N_34972);
or U37529 (N_37529,N_33761,N_31617);
nor U37530 (N_37530,N_32295,N_34090);
nor U37531 (N_37531,N_31480,N_34648);
or U37532 (N_37532,N_31799,N_32519);
xor U37533 (N_37533,N_31116,N_30313);
xnor U37534 (N_37534,N_33263,N_32103);
nand U37535 (N_37535,N_31797,N_32408);
and U37536 (N_37536,N_30335,N_31533);
nor U37537 (N_37537,N_32593,N_32537);
or U37538 (N_37538,N_34579,N_30884);
or U37539 (N_37539,N_33519,N_32272);
nand U37540 (N_37540,N_34308,N_31213);
nand U37541 (N_37541,N_30485,N_34664);
nor U37542 (N_37542,N_32242,N_31876);
xnor U37543 (N_37543,N_34006,N_31297);
and U37544 (N_37544,N_34875,N_34507);
and U37545 (N_37545,N_33942,N_32463);
nor U37546 (N_37546,N_33473,N_31649);
xor U37547 (N_37547,N_32223,N_33524);
and U37548 (N_37548,N_30416,N_31678);
or U37549 (N_37549,N_31871,N_33615);
or U37550 (N_37550,N_34255,N_34625);
and U37551 (N_37551,N_32885,N_31480);
nor U37552 (N_37552,N_30320,N_33768);
nand U37553 (N_37553,N_32923,N_33041);
nand U37554 (N_37554,N_32064,N_30838);
xnor U37555 (N_37555,N_31654,N_34010);
or U37556 (N_37556,N_34694,N_31336);
xnor U37557 (N_37557,N_30794,N_34929);
nor U37558 (N_37558,N_31756,N_31854);
xnor U37559 (N_37559,N_30180,N_31583);
xor U37560 (N_37560,N_31628,N_33916);
or U37561 (N_37561,N_33395,N_32167);
and U37562 (N_37562,N_31327,N_32997);
and U37563 (N_37563,N_33357,N_32564);
xnor U37564 (N_37564,N_31639,N_31173);
and U37565 (N_37565,N_32972,N_31922);
nor U37566 (N_37566,N_34532,N_33303);
xor U37567 (N_37567,N_31093,N_33267);
nor U37568 (N_37568,N_34252,N_32504);
xor U37569 (N_37569,N_34273,N_31682);
xnor U37570 (N_37570,N_32157,N_34244);
xnor U37571 (N_37571,N_31906,N_32121);
xor U37572 (N_37572,N_34794,N_30543);
or U37573 (N_37573,N_30365,N_34209);
or U37574 (N_37574,N_33706,N_34952);
nor U37575 (N_37575,N_32492,N_33878);
or U37576 (N_37576,N_30512,N_34673);
nand U37577 (N_37577,N_33645,N_31739);
nand U37578 (N_37578,N_33457,N_34667);
or U37579 (N_37579,N_33933,N_32530);
xnor U37580 (N_37580,N_34996,N_33080);
nand U37581 (N_37581,N_31783,N_34109);
or U37582 (N_37582,N_33583,N_33351);
or U37583 (N_37583,N_32261,N_33817);
and U37584 (N_37584,N_31748,N_34795);
and U37585 (N_37585,N_30411,N_34438);
xor U37586 (N_37586,N_30707,N_32269);
or U37587 (N_37587,N_34714,N_33561);
and U37588 (N_37588,N_30083,N_33700);
nor U37589 (N_37589,N_31222,N_31545);
nor U37590 (N_37590,N_31485,N_34859);
nor U37591 (N_37591,N_32045,N_34393);
nor U37592 (N_37592,N_34462,N_31329);
nand U37593 (N_37593,N_31551,N_34817);
nand U37594 (N_37594,N_33231,N_31509);
nand U37595 (N_37595,N_31654,N_31040);
nor U37596 (N_37596,N_30393,N_34491);
nand U37597 (N_37597,N_31552,N_31606);
or U37598 (N_37598,N_31951,N_30404);
or U37599 (N_37599,N_33644,N_32743);
nor U37600 (N_37600,N_30115,N_30004);
xnor U37601 (N_37601,N_33938,N_34559);
or U37602 (N_37602,N_34163,N_32948);
xor U37603 (N_37603,N_30026,N_34733);
nor U37604 (N_37604,N_31273,N_30327);
nor U37605 (N_37605,N_32870,N_34255);
xor U37606 (N_37606,N_32451,N_34029);
xnor U37607 (N_37607,N_32373,N_33121);
xor U37608 (N_37608,N_34086,N_33969);
nand U37609 (N_37609,N_30930,N_33116);
nor U37610 (N_37610,N_33586,N_30865);
nand U37611 (N_37611,N_32768,N_33590);
xnor U37612 (N_37612,N_31832,N_30762);
nor U37613 (N_37613,N_31386,N_31892);
or U37614 (N_37614,N_30789,N_31333);
or U37615 (N_37615,N_32150,N_32792);
xnor U37616 (N_37616,N_33902,N_30855);
and U37617 (N_37617,N_33108,N_34972);
xnor U37618 (N_37618,N_32038,N_33246);
xor U37619 (N_37619,N_30848,N_34009);
or U37620 (N_37620,N_34982,N_30003);
or U37621 (N_37621,N_33799,N_31662);
xnor U37622 (N_37622,N_34111,N_33004);
and U37623 (N_37623,N_30203,N_31830);
xnor U37624 (N_37624,N_34811,N_31006);
xor U37625 (N_37625,N_31969,N_31924);
or U37626 (N_37626,N_30742,N_33574);
or U37627 (N_37627,N_31723,N_30442);
and U37628 (N_37628,N_30313,N_31025);
xnor U37629 (N_37629,N_32368,N_34490);
or U37630 (N_37630,N_32579,N_33392);
and U37631 (N_37631,N_33952,N_30978);
xor U37632 (N_37632,N_32464,N_31198);
nand U37633 (N_37633,N_30413,N_33884);
and U37634 (N_37634,N_30706,N_34629);
nand U37635 (N_37635,N_30506,N_31849);
and U37636 (N_37636,N_33110,N_34367);
nor U37637 (N_37637,N_34520,N_30438);
and U37638 (N_37638,N_33025,N_30876);
nand U37639 (N_37639,N_34805,N_32162);
nor U37640 (N_37640,N_32338,N_34778);
xnor U37641 (N_37641,N_34883,N_33693);
or U37642 (N_37642,N_33960,N_33128);
nand U37643 (N_37643,N_30929,N_32375);
or U37644 (N_37644,N_31777,N_33387);
nor U37645 (N_37645,N_33934,N_30739);
and U37646 (N_37646,N_31485,N_34620);
and U37647 (N_37647,N_30768,N_32375);
nand U37648 (N_37648,N_31709,N_34342);
nor U37649 (N_37649,N_34299,N_30991);
nor U37650 (N_37650,N_33793,N_32987);
or U37651 (N_37651,N_33267,N_32206);
and U37652 (N_37652,N_30779,N_34697);
nor U37653 (N_37653,N_33969,N_31822);
nand U37654 (N_37654,N_31580,N_30706);
xor U37655 (N_37655,N_34316,N_34155);
or U37656 (N_37656,N_32259,N_33116);
nand U37657 (N_37657,N_33943,N_31627);
and U37658 (N_37658,N_33018,N_31076);
nor U37659 (N_37659,N_32529,N_32399);
or U37660 (N_37660,N_33639,N_33776);
nand U37661 (N_37661,N_34562,N_32383);
nand U37662 (N_37662,N_31113,N_34462);
nor U37663 (N_37663,N_33018,N_31190);
and U37664 (N_37664,N_31875,N_33924);
xor U37665 (N_37665,N_31497,N_34043);
nor U37666 (N_37666,N_34054,N_30300);
nand U37667 (N_37667,N_34148,N_33584);
nand U37668 (N_37668,N_30469,N_33194);
or U37669 (N_37669,N_33456,N_34568);
or U37670 (N_37670,N_31176,N_33046);
nand U37671 (N_37671,N_34961,N_34685);
xor U37672 (N_37672,N_32915,N_32524);
nand U37673 (N_37673,N_32638,N_32576);
or U37674 (N_37674,N_30346,N_34294);
or U37675 (N_37675,N_33862,N_31648);
xnor U37676 (N_37676,N_33059,N_30089);
and U37677 (N_37677,N_32771,N_32655);
nor U37678 (N_37678,N_30758,N_33219);
or U37679 (N_37679,N_30390,N_32955);
and U37680 (N_37680,N_32507,N_33147);
or U37681 (N_37681,N_34147,N_32388);
and U37682 (N_37682,N_32708,N_31889);
or U37683 (N_37683,N_30756,N_31528);
nor U37684 (N_37684,N_33889,N_34989);
or U37685 (N_37685,N_31470,N_33838);
and U37686 (N_37686,N_30230,N_32768);
nor U37687 (N_37687,N_34385,N_33255);
nand U37688 (N_37688,N_31572,N_34674);
xnor U37689 (N_37689,N_31703,N_33338);
or U37690 (N_37690,N_32758,N_31974);
xor U37691 (N_37691,N_31308,N_34117);
xnor U37692 (N_37692,N_34843,N_32264);
and U37693 (N_37693,N_32891,N_31181);
nor U37694 (N_37694,N_34032,N_30285);
and U37695 (N_37695,N_34190,N_30649);
nand U37696 (N_37696,N_34700,N_34152);
and U37697 (N_37697,N_30161,N_30619);
or U37698 (N_37698,N_30600,N_34770);
or U37699 (N_37699,N_33574,N_31398);
nand U37700 (N_37700,N_34643,N_33778);
nor U37701 (N_37701,N_30414,N_33396);
and U37702 (N_37702,N_31187,N_34202);
and U37703 (N_37703,N_30044,N_32844);
nor U37704 (N_37704,N_34771,N_32074);
and U37705 (N_37705,N_33237,N_31839);
and U37706 (N_37706,N_32941,N_30100);
xor U37707 (N_37707,N_33010,N_30101);
nor U37708 (N_37708,N_33376,N_32830);
or U37709 (N_37709,N_34732,N_34937);
nand U37710 (N_37710,N_32051,N_34606);
nand U37711 (N_37711,N_33665,N_31712);
xnor U37712 (N_37712,N_31264,N_32724);
nand U37713 (N_37713,N_32012,N_31524);
or U37714 (N_37714,N_31821,N_34297);
xor U37715 (N_37715,N_32879,N_34582);
nand U37716 (N_37716,N_32260,N_30429);
xnor U37717 (N_37717,N_34016,N_30206);
or U37718 (N_37718,N_33410,N_34058);
xnor U37719 (N_37719,N_31498,N_31512);
xor U37720 (N_37720,N_33259,N_32315);
nand U37721 (N_37721,N_31263,N_33710);
or U37722 (N_37722,N_34038,N_34148);
xnor U37723 (N_37723,N_30325,N_30943);
and U37724 (N_37724,N_32609,N_30012);
and U37725 (N_37725,N_31757,N_30010);
nor U37726 (N_37726,N_34010,N_32174);
xor U37727 (N_37727,N_34368,N_32331);
and U37728 (N_37728,N_34753,N_31270);
or U37729 (N_37729,N_31845,N_34859);
xor U37730 (N_37730,N_32337,N_31105);
xnor U37731 (N_37731,N_32697,N_32632);
nand U37732 (N_37732,N_32967,N_33946);
nand U37733 (N_37733,N_32772,N_34399);
nor U37734 (N_37734,N_31745,N_30110);
and U37735 (N_37735,N_33197,N_30353);
and U37736 (N_37736,N_30061,N_31463);
or U37737 (N_37737,N_32066,N_32257);
and U37738 (N_37738,N_33843,N_30778);
nor U37739 (N_37739,N_30612,N_33882);
or U37740 (N_37740,N_34471,N_32268);
nor U37741 (N_37741,N_34009,N_34142);
nand U37742 (N_37742,N_31758,N_33311);
nand U37743 (N_37743,N_32494,N_30413);
or U37744 (N_37744,N_33611,N_33729);
or U37745 (N_37745,N_34965,N_32516);
nor U37746 (N_37746,N_34774,N_30867);
xor U37747 (N_37747,N_34088,N_31398);
and U37748 (N_37748,N_30859,N_30670);
xor U37749 (N_37749,N_34325,N_32832);
or U37750 (N_37750,N_30630,N_31044);
and U37751 (N_37751,N_31031,N_34972);
xnor U37752 (N_37752,N_34739,N_32202);
xor U37753 (N_37753,N_32656,N_33511);
or U37754 (N_37754,N_32172,N_30732);
nor U37755 (N_37755,N_34522,N_34793);
xor U37756 (N_37756,N_30484,N_32635);
and U37757 (N_37757,N_30898,N_34164);
nand U37758 (N_37758,N_31712,N_33214);
nand U37759 (N_37759,N_32668,N_33704);
xnor U37760 (N_37760,N_33433,N_32442);
nand U37761 (N_37761,N_33593,N_32722);
nand U37762 (N_37762,N_31406,N_34845);
xor U37763 (N_37763,N_33831,N_30372);
or U37764 (N_37764,N_34623,N_33646);
nor U37765 (N_37765,N_33787,N_33003);
and U37766 (N_37766,N_30325,N_33322);
and U37767 (N_37767,N_31224,N_31784);
xnor U37768 (N_37768,N_32365,N_34104);
nand U37769 (N_37769,N_32091,N_31436);
or U37770 (N_37770,N_32499,N_32537);
xnor U37771 (N_37771,N_31705,N_31868);
or U37772 (N_37772,N_34487,N_31968);
nand U37773 (N_37773,N_34140,N_30720);
and U37774 (N_37774,N_32480,N_34577);
nor U37775 (N_37775,N_31525,N_30716);
and U37776 (N_37776,N_34269,N_32916);
nand U37777 (N_37777,N_32164,N_34116);
or U37778 (N_37778,N_34110,N_34173);
nand U37779 (N_37779,N_34116,N_34210);
nand U37780 (N_37780,N_32365,N_32966);
or U37781 (N_37781,N_31891,N_34094);
or U37782 (N_37782,N_34740,N_33364);
xnor U37783 (N_37783,N_34280,N_31093);
nor U37784 (N_37784,N_30404,N_33840);
or U37785 (N_37785,N_33353,N_33300);
nor U37786 (N_37786,N_33907,N_31691);
xor U37787 (N_37787,N_34762,N_31047);
nand U37788 (N_37788,N_31811,N_31068);
xor U37789 (N_37789,N_34829,N_30707);
or U37790 (N_37790,N_31408,N_32136);
or U37791 (N_37791,N_32609,N_32028);
nor U37792 (N_37792,N_34540,N_31670);
and U37793 (N_37793,N_33750,N_33576);
nor U37794 (N_37794,N_34456,N_33361);
nand U37795 (N_37795,N_32527,N_33907);
and U37796 (N_37796,N_32532,N_32431);
and U37797 (N_37797,N_31407,N_33035);
nand U37798 (N_37798,N_31205,N_33720);
and U37799 (N_37799,N_31251,N_32971);
xor U37800 (N_37800,N_33722,N_31657);
nor U37801 (N_37801,N_30946,N_32970);
or U37802 (N_37802,N_33055,N_33457);
or U37803 (N_37803,N_33690,N_30580);
and U37804 (N_37804,N_33557,N_31120);
nor U37805 (N_37805,N_30853,N_30804);
xor U37806 (N_37806,N_34626,N_31110);
nor U37807 (N_37807,N_32751,N_32717);
nand U37808 (N_37808,N_30129,N_31568);
or U37809 (N_37809,N_31185,N_34458);
nor U37810 (N_37810,N_32357,N_32161);
nand U37811 (N_37811,N_33783,N_31717);
nand U37812 (N_37812,N_33869,N_31873);
or U37813 (N_37813,N_34239,N_33241);
xor U37814 (N_37814,N_30903,N_34926);
nand U37815 (N_37815,N_30868,N_34520);
nand U37816 (N_37816,N_32742,N_33835);
nor U37817 (N_37817,N_31992,N_32350);
xor U37818 (N_37818,N_34277,N_32782);
and U37819 (N_37819,N_31778,N_31443);
nand U37820 (N_37820,N_32962,N_33898);
nand U37821 (N_37821,N_31935,N_34088);
or U37822 (N_37822,N_32373,N_30198);
nor U37823 (N_37823,N_30461,N_32247);
and U37824 (N_37824,N_30264,N_30053);
xor U37825 (N_37825,N_31860,N_30070);
nor U37826 (N_37826,N_33974,N_33728);
nor U37827 (N_37827,N_32960,N_32131);
nor U37828 (N_37828,N_31216,N_32196);
xor U37829 (N_37829,N_34498,N_30522);
nor U37830 (N_37830,N_34911,N_30649);
nand U37831 (N_37831,N_31416,N_30676);
nor U37832 (N_37832,N_34995,N_34158);
and U37833 (N_37833,N_30857,N_32362);
nor U37834 (N_37834,N_34159,N_32786);
nor U37835 (N_37835,N_31704,N_34570);
nor U37836 (N_37836,N_33256,N_32066);
nor U37837 (N_37837,N_33560,N_33670);
nor U37838 (N_37838,N_33153,N_34885);
nor U37839 (N_37839,N_33340,N_30944);
nor U37840 (N_37840,N_33763,N_32530);
and U37841 (N_37841,N_30068,N_34396);
nor U37842 (N_37842,N_33452,N_30114);
nor U37843 (N_37843,N_33427,N_31992);
or U37844 (N_37844,N_34430,N_34272);
nor U37845 (N_37845,N_30073,N_31669);
nand U37846 (N_37846,N_34789,N_30568);
and U37847 (N_37847,N_32250,N_31190);
xnor U37848 (N_37848,N_32169,N_31693);
or U37849 (N_37849,N_31281,N_31821);
nand U37850 (N_37850,N_34394,N_32566);
or U37851 (N_37851,N_31237,N_34625);
xnor U37852 (N_37852,N_33147,N_30051);
or U37853 (N_37853,N_30273,N_34690);
or U37854 (N_37854,N_31757,N_31482);
nand U37855 (N_37855,N_32321,N_33194);
or U37856 (N_37856,N_30764,N_30974);
nand U37857 (N_37857,N_32037,N_33794);
nor U37858 (N_37858,N_34207,N_33208);
xor U37859 (N_37859,N_33845,N_32901);
xor U37860 (N_37860,N_31325,N_30776);
nand U37861 (N_37861,N_30225,N_30304);
xnor U37862 (N_37862,N_31602,N_34989);
nand U37863 (N_37863,N_30007,N_30420);
or U37864 (N_37864,N_33192,N_30768);
or U37865 (N_37865,N_30684,N_34713);
or U37866 (N_37866,N_34442,N_34324);
nor U37867 (N_37867,N_32561,N_30515);
xnor U37868 (N_37868,N_30250,N_30005);
xor U37869 (N_37869,N_33383,N_34479);
or U37870 (N_37870,N_30428,N_31846);
nor U37871 (N_37871,N_31602,N_33731);
and U37872 (N_37872,N_31576,N_30827);
nand U37873 (N_37873,N_31973,N_32321);
nand U37874 (N_37874,N_32277,N_32132);
nand U37875 (N_37875,N_31251,N_34932);
nand U37876 (N_37876,N_32001,N_30562);
xnor U37877 (N_37877,N_34527,N_32259);
nor U37878 (N_37878,N_31536,N_30986);
nand U37879 (N_37879,N_34692,N_34744);
nor U37880 (N_37880,N_31530,N_31677);
nor U37881 (N_37881,N_30363,N_33943);
nor U37882 (N_37882,N_34406,N_30301);
and U37883 (N_37883,N_32815,N_30564);
nor U37884 (N_37884,N_33634,N_33911);
nor U37885 (N_37885,N_34531,N_34983);
and U37886 (N_37886,N_31717,N_34680);
xnor U37887 (N_37887,N_33901,N_33764);
or U37888 (N_37888,N_31419,N_34243);
nor U37889 (N_37889,N_33952,N_33256);
or U37890 (N_37890,N_32861,N_31104);
xnor U37891 (N_37891,N_32372,N_34621);
or U37892 (N_37892,N_34048,N_30188);
and U37893 (N_37893,N_33521,N_32775);
nor U37894 (N_37894,N_33094,N_33285);
or U37895 (N_37895,N_31373,N_34381);
nor U37896 (N_37896,N_34298,N_30328);
xor U37897 (N_37897,N_31213,N_32755);
nand U37898 (N_37898,N_34000,N_32967);
xor U37899 (N_37899,N_34587,N_31330);
xnor U37900 (N_37900,N_34679,N_31048);
and U37901 (N_37901,N_33562,N_33402);
nor U37902 (N_37902,N_32358,N_34542);
or U37903 (N_37903,N_30119,N_31445);
and U37904 (N_37904,N_31888,N_30202);
nor U37905 (N_37905,N_34586,N_33405);
nand U37906 (N_37906,N_34124,N_32612);
and U37907 (N_37907,N_34979,N_30745);
nor U37908 (N_37908,N_32348,N_33767);
or U37909 (N_37909,N_30479,N_33529);
xnor U37910 (N_37910,N_34330,N_30468);
xnor U37911 (N_37911,N_33771,N_31210);
xnor U37912 (N_37912,N_33693,N_32193);
xnor U37913 (N_37913,N_30899,N_32876);
xnor U37914 (N_37914,N_33147,N_32141);
or U37915 (N_37915,N_34922,N_31156);
nor U37916 (N_37916,N_30085,N_34377);
xnor U37917 (N_37917,N_31766,N_32858);
nand U37918 (N_37918,N_33277,N_32705);
and U37919 (N_37919,N_33111,N_31556);
nand U37920 (N_37920,N_30890,N_32133);
or U37921 (N_37921,N_31860,N_31996);
nand U37922 (N_37922,N_34253,N_34663);
and U37923 (N_37923,N_30771,N_34488);
nand U37924 (N_37924,N_30180,N_32553);
xor U37925 (N_37925,N_31479,N_31920);
and U37926 (N_37926,N_31786,N_34009);
nand U37927 (N_37927,N_33640,N_34154);
or U37928 (N_37928,N_31843,N_33679);
or U37929 (N_37929,N_33402,N_30161);
or U37930 (N_37930,N_34225,N_34710);
nor U37931 (N_37931,N_30315,N_31409);
nand U37932 (N_37932,N_32619,N_34631);
and U37933 (N_37933,N_30344,N_32936);
xor U37934 (N_37934,N_33877,N_30518);
nor U37935 (N_37935,N_32734,N_34864);
or U37936 (N_37936,N_32300,N_33967);
nand U37937 (N_37937,N_33181,N_31113);
nor U37938 (N_37938,N_30421,N_32715);
nor U37939 (N_37939,N_34184,N_33253);
or U37940 (N_37940,N_31750,N_32435);
nand U37941 (N_37941,N_32128,N_33924);
and U37942 (N_37942,N_30959,N_32131);
xor U37943 (N_37943,N_31952,N_30484);
nand U37944 (N_37944,N_32907,N_33139);
nor U37945 (N_37945,N_32191,N_33625);
nand U37946 (N_37946,N_33016,N_30411);
or U37947 (N_37947,N_32129,N_30041);
and U37948 (N_37948,N_30261,N_31996);
or U37949 (N_37949,N_30933,N_32287);
nor U37950 (N_37950,N_33822,N_32906);
nor U37951 (N_37951,N_30607,N_33388);
nand U37952 (N_37952,N_32948,N_32212);
nand U37953 (N_37953,N_30299,N_30085);
xor U37954 (N_37954,N_30543,N_31948);
nand U37955 (N_37955,N_30044,N_33209);
nand U37956 (N_37956,N_30989,N_30231);
or U37957 (N_37957,N_31136,N_31143);
or U37958 (N_37958,N_33416,N_31418);
or U37959 (N_37959,N_34012,N_31128);
nand U37960 (N_37960,N_33464,N_32449);
or U37961 (N_37961,N_33895,N_34062);
or U37962 (N_37962,N_32437,N_31977);
and U37963 (N_37963,N_31752,N_30752);
nand U37964 (N_37964,N_30055,N_31706);
and U37965 (N_37965,N_34419,N_30167);
and U37966 (N_37966,N_32839,N_33943);
nor U37967 (N_37967,N_30384,N_31565);
nand U37968 (N_37968,N_32664,N_30360);
or U37969 (N_37969,N_33525,N_32403);
nor U37970 (N_37970,N_33153,N_31931);
or U37971 (N_37971,N_31942,N_32927);
and U37972 (N_37972,N_34335,N_32240);
or U37973 (N_37973,N_31887,N_31048);
nand U37974 (N_37974,N_30600,N_32162);
and U37975 (N_37975,N_31123,N_31039);
nand U37976 (N_37976,N_32818,N_30236);
or U37977 (N_37977,N_31224,N_31891);
nor U37978 (N_37978,N_32148,N_30105);
nand U37979 (N_37979,N_30563,N_30427);
nor U37980 (N_37980,N_31800,N_33944);
and U37981 (N_37981,N_34190,N_30689);
nor U37982 (N_37982,N_32588,N_30462);
or U37983 (N_37983,N_33668,N_33146);
xnor U37984 (N_37984,N_30181,N_33592);
and U37985 (N_37985,N_34111,N_33783);
and U37986 (N_37986,N_31251,N_30981);
xor U37987 (N_37987,N_34606,N_32139);
and U37988 (N_37988,N_33012,N_30639);
or U37989 (N_37989,N_30060,N_34621);
nor U37990 (N_37990,N_30403,N_34065);
and U37991 (N_37991,N_32766,N_30479);
and U37992 (N_37992,N_32799,N_34904);
nor U37993 (N_37993,N_30067,N_34395);
or U37994 (N_37994,N_32839,N_34422);
nor U37995 (N_37995,N_30653,N_30812);
nor U37996 (N_37996,N_33247,N_32874);
xnor U37997 (N_37997,N_33458,N_34464);
nor U37998 (N_37998,N_34606,N_33669);
xnor U37999 (N_37999,N_30723,N_30613);
nand U38000 (N_38000,N_31698,N_31658);
xor U38001 (N_38001,N_34502,N_32183);
and U38002 (N_38002,N_32329,N_34773);
nor U38003 (N_38003,N_34903,N_30653);
nor U38004 (N_38004,N_34465,N_30315);
xor U38005 (N_38005,N_30690,N_32866);
nand U38006 (N_38006,N_30525,N_30626);
and U38007 (N_38007,N_32637,N_33066);
nor U38008 (N_38008,N_34985,N_31842);
and U38009 (N_38009,N_30370,N_33840);
and U38010 (N_38010,N_33610,N_33636);
nand U38011 (N_38011,N_33817,N_30211);
nor U38012 (N_38012,N_31548,N_34573);
and U38013 (N_38013,N_30233,N_34910);
nor U38014 (N_38014,N_33676,N_34876);
nand U38015 (N_38015,N_33157,N_31278);
xor U38016 (N_38016,N_30066,N_34413);
or U38017 (N_38017,N_31738,N_31312);
nand U38018 (N_38018,N_33479,N_34616);
or U38019 (N_38019,N_34691,N_31485);
xor U38020 (N_38020,N_31222,N_34533);
nor U38021 (N_38021,N_30126,N_31013);
or U38022 (N_38022,N_32161,N_34821);
nor U38023 (N_38023,N_34757,N_34055);
nor U38024 (N_38024,N_33165,N_30885);
xnor U38025 (N_38025,N_33990,N_32973);
nand U38026 (N_38026,N_32940,N_34267);
or U38027 (N_38027,N_30481,N_30598);
nand U38028 (N_38028,N_32641,N_32168);
nor U38029 (N_38029,N_34517,N_32504);
xnor U38030 (N_38030,N_32825,N_33739);
or U38031 (N_38031,N_31581,N_30205);
nand U38032 (N_38032,N_30490,N_30951);
nor U38033 (N_38033,N_32665,N_30145);
xnor U38034 (N_38034,N_33917,N_30820);
nand U38035 (N_38035,N_30728,N_30923);
nand U38036 (N_38036,N_31126,N_31428);
xnor U38037 (N_38037,N_33688,N_30802);
nor U38038 (N_38038,N_32619,N_34039);
and U38039 (N_38039,N_34865,N_32191);
nand U38040 (N_38040,N_33216,N_30685);
and U38041 (N_38041,N_30442,N_34745);
xnor U38042 (N_38042,N_33096,N_34306);
nand U38043 (N_38043,N_30069,N_34441);
or U38044 (N_38044,N_34271,N_34724);
and U38045 (N_38045,N_34468,N_30075);
or U38046 (N_38046,N_33126,N_31963);
nor U38047 (N_38047,N_30453,N_31190);
and U38048 (N_38048,N_32475,N_30619);
nor U38049 (N_38049,N_34769,N_31692);
nand U38050 (N_38050,N_33587,N_31529);
or U38051 (N_38051,N_34854,N_30058);
nand U38052 (N_38052,N_33688,N_34314);
or U38053 (N_38053,N_30710,N_30771);
or U38054 (N_38054,N_33439,N_33952);
xnor U38055 (N_38055,N_31349,N_30468);
nand U38056 (N_38056,N_34020,N_32389);
or U38057 (N_38057,N_30818,N_33447);
xnor U38058 (N_38058,N_34194,N_32052);
nor U38059 (N_38059,N_30345,N_33679);
nor U38060 (N_38060,N_30984,N_32461);
nand U38061 (N_38061,N_33400,N_34717);
nand U38062 (N_38062,N_34045,N_32546);
nor U38063 (N_38063,N_30753,N_32015);
nand U38064 (N_38064,N_30685,N_32869);
xor U38065 (N_38065,N_30667,N_32741);
nor U38066 (N_38066,N_31128,N_33650);
nor U38067 (N_38067,N_30010,N_34047);
nand U38068 (N_38068,N_33348,N_30451);
nor U38069 (N_38069,N_31328,N_34862);
nand U38070 (N_38070,N_34365,N_34213);
or U38071 (N_38071,N_31326,N_33987);
and U38072 (N_38072,N_30250,N_33301);
and U38073 (N_38073,N_34788,N_33641);
xnor U38074 (N_38074,N_30152,N_30334);
and U38075 (N_38075,N_32934,N_31631);
and U38076 (N_38076,N_33143,N_34764);
and U38077 (N_38077,N_34746,N_31546);
xnor U38078 (N_38078,N_34028,N_32656);
xnor U38079 (N_38079,N_34371,N_30081);
and U38080 (N_38080,N_30080,N_31465);
or U38081 (N_38081,N_34478,N_30677);
xnor U38082 (N_38082,N_31123,N_34395);
nand U38083 (N_38083,N_34747,N_33427);
or U38084 (N_38084,N_34752,N_30343);
and U38085 (N_38085,N_32353,N_30527);
nor U38086 (N_38086,N_31215,N_34837);
nand U38087 (N_38087,N_32683,N_30100);
nand U38088 (N_38088,N_31181,N_31296);
or U38089 (N_38089,N_31689,N_32254);
xnor U38090 (N_38090,N_32021,N_33592);
nor U38091 (N_38091,N_31472,N_33501);
xor U38092 (N_38092,N_32452,N_31853);
or U38093 (N_38093,N_33012,N_34895);
nor U38094 (N_38094,N_31552,N_32392);
xnor U38095 (N_38095,N_31459,N_31182);
or U38096 (N_38096,N_34855,N_31745);
xor U38097 (N_38097,N_34273,N_32559);
nand U38098 (N_38098,N_34571,N_32083);
and U38099 (N_38099,N_31280,N_33258);
nand U38100 (N_38100,N_31221,N_32200);
and U38101 (N_38101,N_30097,N_31922);
xnor U38102 (N_38102,N_32943,N_34154);
or U38103 (N_38103,N_30629,N_34471);
xor U38104 (N_38104,N_30313,N_32000);
xor U38105 (N_38105,N_34276,N_30843);
nor U38106 (N_38106,N_32175,N_33156);
nor U38107 (N_38107,N_30970,N_34171);
or U38108 (N_38108,N_33751,N_32909);
xnor U38109 (N_38109,N_31663,N_33745);
or U38110 (N_38110,N_34590,N_34400);
xor U38111 (N_38111,N_32342,N_32377);
xor U38112 (N_38112,N_30017,N_31780);
xnor U38113 (N_38113,N_32643,N_32266);
xnor U38114 (N_38114,N_32683,N_34145);
or U38115 (N_38115,N_30503,N_34045);
or U38116 (N_38116,N_34462,N_34087);
or U38117 (N_38117,N_32160,N_30140);
xnor U38118 (N_38118,N_31487,N_31383);
or U38119 (N_38119,N_34476,N_30928);
xnor U38120 (N_38120,N_32188,N_31052);
xnor U38121 (N_38121,N_30382,N_30678);
nand U38122 (N_38122,N_33477,N_30823);
xor U38123 (N_38123,N_30000,N_32733);
nor U38124 (N_38124,N_32238,N_34431);
nand U38125 (N_38125,N_30274,N_30920);
or U38126 (N_38126,N_31100,N_31947);
and U38127 (N_38127,N_32297,N_34414);
and U38128 (N_38128,N_34884,N_33337);
nand U38129 (N_38129,N_30883,N_31825);
nor U38130 (N_38130,N_32294,N_34166);
or U38131 (N_38131,N_32240,N_32118);
nor U38132 (N_38132,N_33903,N_32837);
xor U38133 (N_38133,N_33214,N_32078);
nor U38134 (N_38134,N_32882,N_30852);
or U38135 (N_38135,N_31000,N_30339);
or U38136 (N_38136,N_30837,N_30741);
nand U38137 (N_38137,N_31660,N_31291);
xor U38138 (N_38138,N_34816,N_34175);
xnor U38139 (N_38139,N_32513,N_30251);
or U38140 (N_38140,N_31659,N_32910);
nor U38141 (N_38141,N_32392,N_32546);
or U38142 (N_38142,N_33747,N_32515);
and U38143 (N_38143,N_30304,N_30188);
xnor U38144 (N_38144,N_30139,N_34214);
or U38145 (N_38145,N_33265,N_30212);
nand U38146 (N_38146,N_31346,N_30868);
xnor U38147 (N_38147,N_32446,N_33389);
nor U38148 (N_38148,N_33294,N_30485);
or U38149 (N_38149,N_34560,N_33068);
nor U38150 (N_38150,N_32942,N_31904);
xnor U38151 (N_38151,N_32659,N_30964);
nand U38152 (N_38152,N_31733,N_34150);
xor U38153 (N_38153,N_33642,N_34032);
and U38154 (N_38154,N_34091,N_31841);
nor U38155 (N_38155,N_31204,N_34472);
or U38156 (N_38156,N_31624,N_32102);
nand U38157 (N_38157,N_31759,N_30510);
nand U38158 (N_38158,N_33516,N_33311);
nor U38159 (N_38159,N_32255,N_34810);
xnor U38160 (N_38160,N_31636,N_31017);
or U38161 (N_38161,N_31321,N_30679);
and U38162 (N_38162,N_30332,N_33885);
and U38163 (N_38163,N_30906,N_32073);
xnor U38164 (N_38164,N_32505,N_32933);
or U38165 (N_38165,N_34856,N_32143);
nand U38166 (N_38166,N_30591,N_34067);
xor U38167 (N_38167,N_32708,N_32995);
nand U38168 (N_38168,N_32658,N_33705);
or U38169 (N_38169,N_31423,N_30573);
xnor U38170 (N_38170,N_34521,N_32401);
nor U38171 (N_38171,N_30485,N_34505);
nor U38172 (N_38172,N_31071,N_30235);
and U38173 (N_38173,N_33952,N_31766);
and U38174 (N_38174,N_33007,N_33118);
nor U38175 (N_38175,N_30932,N_30397);
or U38176 (N_38176,N_31482,N_34585);
or U38177 (N_38177,N_32710,N_34914);
nor U38178 (N_38178,N_32859,N_33141);
nand U38179 (N_38179,N_34758,N_33298);
and U38180 (N_38180,N_34675,N_34455);
xnor U38181 (N_38181,N_34384,N_31355);
and U38182 (N_38182,N_34469,N_34330);
and U38183 (N_38183,N_30192,N_33231);
xor U38184 (N_38184,N_33184,N_33633);
xor U38185 (N_38185,N_33644,N_31145);
xnor U38186 (N_38186,N_34992,N_31770);
or U38187 (N_38187,N_30295,N_31772);
or U38188 (N_38188,N_34818,N_34638);
or U38189 (N_38189,N_32853,N_33505);
xnor U38190 (N_38190,N_34074,N_34152);
and U38191 (N_38191,N_33637,N_30080);
and U38192 (N_38192,N_33162,N_31260);
and U38193 (N_38193,N_31811,N_30182);
nand U38194 (N_38194,N_32486,N_30844);
or U38195 (N_38195,N_32970,N_30078);
or U38196 (N_38196,N_34065,N_32760);
nor U38197 (N_38197,N_33100,N_31918);
nor U38198 (N_38198,N_34470,N_31270);
and U38199 (N_38199,N_30876,N_33819);
nor U38200 (N_38200,N_30839,N_32055);
or U38201 (N_38201,N_33180,N_31960);
nand U38202 (N_38202,N_32988,N_31377);
xnor U38203 (N_38203,N_30572,N_34537);
nor U38204 (N_38204,N_34962,N_32869);
or U38205 (N_38205,N_30199,N_31463);
or U38206 (N_38206,N_33415,N_34277);
xnor U38207 (N_38207,N_33412,N_32884);
nand U38208 (N_38208,N_30706,N_32396);
xnor U38209 (N_38209,N_30839,N_33692);
or U38210 (N_38210,N_30923,N_31490);
or U38211 (N_38211,N_33525,N_33150);
nand U38212 (N_38212,N_34454,N_31654);
or U38213 (N_38213,N_32802,N_33592);
and U38214 (N_38214,N_32117,N_30695);
nor U38215 (N_38215,N_34876,N_32778);
xnor U38216 (N_38216,N_30208,N_30124);
nor U38217 (N_38217,N_30548,N_31018);
and U38218 (N_38218,N_30021,N_32754);
xnor U38219 (N_38219,N_34027,N_30140);
nor U38220 (N_38220,N_32543,N_31427);
or U38221 (N_38221,N_34480,N_33428);
or U38222 (N_38222,N_34826,N_33213);
or U38223 (N_38223,N_34925,N_30810);
and U38224 (N_38224,N_31685,N_31359);
nand U38225 (N_38225,N_33702,N_32897);
or U38226 (N_38226,N_34399,N_34581);
and U38227 (N_38227,N_33018,N_31712);
xnor U38228 (N_38228,N_32825,N_34142);
nand U38229 (N_38229,N_31088,N_31663);
xor U38230 (N_38230,N_34675,N_30539);
xnor U38231 (N_38231,N_33699,N_32782);
and U38232 (N_38232,N_33409,N_31595);
and U38233 (N_38233,N_31193,N_31794);
and U38234 (N_38234,N_34654,N_33203);
xnor U38235 (N_38235,N_30001,N_34968);
or U38236 (N_38236,N_34602,N_33850);
or U38237 (N_38237,N_33320,N_32476);
or U38238 (N_38238,N_34507,N_34852);
xor U38239 (N_38239,N_32108,N_30447);
or U38240 (N_38240,N_30134,N_34028);
xnor U38241 (N_38241,N_34252,N_31820);
xnor U38242 (N_38242,N_30898,N_33208);
or U38243 (N_38243,N_33685,N_31256);
or U38244 (N_38244,N_34342,N_32131);
nand U38245 (N_38245,N_32635,N_32365);
nand U38246 (N_38246,N_31493,N_34388);
nor U38247 (N_38247,N_30654,N_31408);
nand U38248 (N_38248,N_33328,N_34653);
or U38249 (N_38249,N_33814,N_30582);
xnor U38250 (N_38250,N_30731,N_30361);
or U38251 (N_38251,N_32753,N_33611);
nor U38252 (N_38252,N_30571,N_33000);
xor U38253 (N_38253,N_30068,N_31362);
nor U38254 (N_38254,N_31263,N_34630);
and U38255 (N_38255,N_32263,N_34322);
and U38256 (N_38256,N_32504,N_32471);
nor U38257 (N_38257,N_34487,N_30686);
nand U38258 (N_38258,N_31621,N_30227);
and U38259 (N_38259,N_33725,N_30908);
xnor U38260 (N_38260,N_34467,N_32273);
xnor U38261 (N_38261,N_34350,N_32901);
nand U38262 (N_38262,N_33633,N_31444);
xor U38263 (N_38263,N_31339,N_30127);
nand U38264 (N_38264,N_30478,N_32420);
nor U38265 (N_38265,N_31431,N_33304);
nand U38266 (N_38266,N_31947,N_32927);
and U38267 (N_38267,N_30383,N_32252);
xnor U38268 (N_38268,N_33243,N_32774);
nand U38269 (N_38269,N_30297,N_34575);
and U38270 (N_38270,N_34096,N_32827);
nor U38271 (N_38271,N_30048,N_31635);
and U38272 (N_38272,N_32055,N_33815);
and U38273 (N_38273,N_31461,N_33641);
or U38274 (N_38274,N_33279,N_32315);
xnor U38275 (N_38275,N_33675,N_31774);
nor U38276 (N_38276,N_31852,N_31609);
xor U38277 (N_38277,N_32222,N_31744);
nand U38278 (N_38278,N_30478,N_33943);
xor U38279 (N_38279,N_30036,N_32519);
xor U38280 (N_38280,N_33003,N_34846);
and U38281 (N_38281,N_31191,N_34589);
nand U38282 (N_38282,N_30899,N_32547);
and U38283 (N_38283,N_34710,N_33399);
nand U38284 (N_38284,N_30625,N_33808);
or U38285 (N_38285,N_30249,N_31543);
nor U38286 (N_38286,N_34905,N_34977);
or U38287 (N_38287,N_31724,N_31229);
xnor U38288 (N_38288,N_34223,N_30166);
nand U38289 (N_38289,N_31895,N_33173);
xor U38290 (N_38290,N_30562,N_34731);
or U38291 (N_38291,N_32142,N_32908);
and U38292 (N_38292,N_30092,N_34185);
nor U38293 (N_38293,N_32357,N_32533);
and U38294 (N_38294,N_34370,N_32348);
and U38295 (N_38295,N_31717,N_30146);
or U38296 (N_38296,N_33386,N_31671);
xor U38297 (N_38297,N_34830,N_34613);
and U38298 (N_38298,N_32622,N_30837);
or U38299 (N_38299,N_31437,N_34879);
nor U38300 (N_38300,N_34099,N_30002);
and U38301 (N_38301,N_33494,N_31043);
nor U38302 (N_38302,N_34901,N_31593);
xor U38303 (N_38303,N_33248,N_33905);
or U38304 (N_38304,N_34798,N_34619);
and U38305 (N_38305,N_32220,N_32720);
nor U38306 (N_38306,N_31821,N_31118);
nand U38307 (N_38307,N_30135,N_31552);
or U38308 (N_38308,N_31956,N_32835);
and U38309 (N_38309,N_31024,N_33991);
nand U38310 (N_38310,N_30438,N_30727);
or U38311 (N_38311,N_34004,N_32316);
and U38312 (N_38312,N_34441,N_32234);
nor U38313 (N_38313,N_34893,N_33468);
or U38314 (N_38314,N_31427,N_30285);
or U38315 (N_38315,N_34150,N_32341);
or U38316 (N_38316,N_31131,N_30275);
and U38317 (N_38317,N_30289,N_33024);
nor U38318 (N_38318,N_32683,N_33188);
nand U38319 (N_38319,N_30398,N_32939);
nand U38320 (N_38320,N_33721,N_34359);
nand U38321 (N_38321,N_32460,N_30016);
and U38322 (N_38322,N_34396,N_32649);
and U38323 (N_38323,N_34475,N_30217);
or U38324 (N_38324,N_32530,N_34878);
nor U38325 (N_38325,N_34362,N_31179);
nor U38326 (N_38326,N_34574,N_30961);
or U38327 (N_38327,N_34433,N_31138);
nor U38328 (N_38328,N_34945,N_30649);
nor U38329 (N_38329,N_32976,N_33339);
and U38330 (N_38330,N_31863,N_33372);
nand U38331 (N_38331,N_34436,N_32815);
and U38332 (N_38332,N_34185,N_34220);
nand U38333 (N_38333,N_31937,N_33882);
or U38334 (N_38334,N_32550,N_31787);
xor U38335 (N_38335,N_32879,N_31912);
nor U38336 (N_38336,N_33284,N_30228);
xor U38337 (N_38337,N_30243,N_34748);
xor U38338 (N_38338,N_32928,N_34174);
nand U38339 (N_38339,N_33992,N_31948);
xnor U38340 (N_38340,N_32199,N_32461);
xnor U38341 (N_38341,N_30389,N_31774);
nor U38342 (N_38342,N_32022,N_31416);
nor U38343 (N_38343,N_31921,N_32567);
nor U38344 (N_38344,N_34236,N_33045);
nor U38345 (N_38345,N_34417,N_32397);
or U38346 (N_38346,N_33211,N_34105);
and U38347 (N_38347,N_31495,N_33747);
or U38348 (N_38348,N_32838,N_32735);
nor U38349 (N_38349,N_34340,N_32887);
nand U38350 (N_38350,N_32956,N_32805);
xor U38351 (N_38351,N_32421,N_33895);
and U38352 (N_38352,N_33350,N_32172);
nor U38353 (N_38353,N_31433,N_34342);
nor U38354 (N_38354,N_31901,N_32017);
or U38355 (N_38355,N_30508,N_34594);
nor U38356 (N_38356,N_30746,N_31177);
nor U38357 (N_38357,N_31801,N_34144);
nand U38358 (N_38358,N_33250,N_34119);
xnor U38359 (N_38359,N_32151,N_31443);
xor U38360 (N_38360,N_32850,N_31241);
or U38361 (N_38361,N_30558,N_31904);
and U38362 (N_38362,N_34385,N_31575);
xor U38363 (N_38363,N_33114,N_33617);
nand U38364 (N_38364,N_30292,N_34592);
or U38365 (N_38365,N_33821,N_32588);
and U38366 (N_38366,N_30947,N_33515);
nor U38367 (N_38367,N_30938,N_34355);
and U38368 (N_38368,N_32817,N_30164);
nand U38369 (N_38369,N_34546,N_34525);
nand U38370 (N_38370,N_33595,N_30078);
and U38371 (N_38371,N_33007,N_34585);
nor U38372 (N_38372,N_34371,N_33165);
nor U38373 (N_38373,N_32217,N_30561);
xnor U38374 (N_38374,N_34068,N_30220);
nand U38375 (N_38375,N_33895,N_30036);
nor U38376 (N_38376,N_34272,N_31498);
xnor U38377 (N_38377,N_32859,N_32201);
nand U38378 (N_38378,N_30420,N_30536);
nand U38379 (N_38379,N_31175,N_34795);
nor U38380 (N_38380,N_30146,N_32328);
nand U38381 (N_38381,N_34125,N_32093);
and U38382 (N_38382,N_32888,N_33389);
and U38383 (N_38383,N_34672,N_33446);
or U38384 (N_38384,N_31191,N_30706);
nor U38385 (N_38385,N_34732,N_30005);
xnor U38386 (N_38386,N_30951,N_32145);
nand U38387 (N_38387,N_30593,N_30598);
nand U38388 (N_38388,N_33958,N_34378);
and U38389 (N_38389,N_32685,N_30277);
and U38390 (N_38390,N_33894,N_34248);
and U38391 (N_38391,N_31921,N_30755);
or U38392 (N_38392,N_33415,N_33500);
xor U38393 (N_38393,N_31786,N_32677);
xor U38394 (N_38394,N_30765,N_34315);
and U38395 (N_38395,N_30332,N_30661);
nand U38396 (N_38396,N_32684,N_30124);
nor U38397 (N_38397,N_33244,N_33203);
and U38398 (N_38398,N_34953,N_33384);
nor U38399 (N_38399,N_34410,N_34834);
or U38400 (N_38400,N_33469,N_31588);
xor U38401 (N_38401,N_30540,N_31343);
and U38402 (N_38402,N_33901,N_30035);
nor U38403 (N_38403,N_32070,N_32584);
or U38404 (N_38404,N_32091,N_32850);
or U38405 (N_38405,N_32730,N_31596);
xnor U38406 (N_38406,N_33423,N_31667);
and U38407 (N_38407,N_31108,N_34119);
nand U38408 (N_38408,N_33617,N_33282);
and U38409 (N_38409,N_32031,N_34215);
nand U38410 (N_38410,N_30686,N_33684);
or U38411 (N_38411,N_30591,N_30998);
nand U38412 (N_38412,N_34090,N_33351);
and U38413 (N_38413,N_34843,N_31875);
nand U38414 (N_38414,N_34366,N_32119);
and U38415 (N_38415,N_30967,N_34292);
and U38416 (N_38416,N_32365,N_30448);
nor U38417 (N_38417,N_32093,N_30361);
and U38418 (N_38418,N_31003,N_34971);
nor U38419 (N_38419,N_30557,N_34061);
or U38420 (N_38420,N_30532,N_30821);
or U38421 (N_38421,N_33185,N_32032);
or U38422 (N_38422,N_32761,N_33499);
and U38423 (N_38423,N_30069,N_30961);
and U38424 (N_38424,N_33443,N_34893);
xnor U38425 (N_38425,N_34430,N_32392);
and U38426 (N_38426,N_33889,N_32526);
nand U38427 (N_38427,N_32884,N_33178);
xor U38428 (N_38428,N_30568,N_34156);
or U38429 (N_38429,N_33039,N_34480);
nand U38430 (N_38430,N_33656,N_30136);
xor U38431 (N_38431,N_31654,N_34591);
or U38432 (N_38432,N_30424,N_32748);
and U38433 (N_38433,N_31874,N_33080);
nand U38434 (N_38434,N_32533,N_34662);
xnor U38435 (N_38435,N_33347,N_30787);
nand U38436 (N_38436,N_33631,N_30240);
nand U38437 (N_38437,N_34807,N_34546);
xnor U38438 (N_38438,N_33661,N_32842);
and U38439 (N_38439,N_31419,N_32781);
or U38440 (N_38440,N_33823,N_33590);
and U38441 (N_38441,N_30901,N_31594);
and U38442 (N_38442,N_32179,N_34977);
nor U38443 (N_38443,N_33880,N_32112);
nor U38444 (N_38444,N_30069,N_34479);
or U38445 (N_38445,N_31987,N_31006);
and U38446 (N_38446,N_31838,N_31463);
and U38447 (N_38447,N_31289,N_34690);
and U38448 (N_38448,N_31252,N_32683);
nor U38449 (N_38449,N_31762,N_33858);
nand U38450 (N_38450,N_30957,N_31561);
and U38451 (N_38451,N_32081,N_32097);
xnor U38452 (N_38452,N_31355,N_30058);
nor U38453 (N_38453,N_34991,N_30890);
nor U38454 (N_38454,N_30011,N_33624);
or U38455 (N_38455,N_32792,N_32598);
and U38456 (N_38456,N_30222,N_32284);
xnor U38457 (N_38457,N_30831,N_34508);
xor U38458 (N_38458,N_30000,N_32594);
and U38459 (N_38459,N_32710,N_34203);
nor U38460 (N_38460,N_32064,N_30448);
or U38461 (N_38461,N_31213,N_32016);
and U38462 (N_38462,N_33826,N_33767);
and U38463 (N_38463,N_30937,N_32802);
xnor U38464 (N_38464,N_30851,N_34120);
nand U38465 (N_38465,N_32287,N_30159);
xnor U38466 (N_38466,N_30912,N_34394);
nor U38467 (N_38467,N_30549,N_31371);
nor U38468 (N_38468,N_30852,N_32563);
nor U38469 (N_38469,N_31625,N_32079);
xnor U38470 (N_38470,N_30447,N_33979);
and U38471 (N_38471,N_30814,N_34261);
or U38472 (N_38472,N_33539,N_32448);
xnor U38473 (N_38473,N_34465,N_32078);
xor U38474 (N_38474,N_31499,N_34117);
xor U38475 (N_38475,N_30552,N_31285);
xnor U38476 (N_38476,N_30350,N_30413);
nand U38477 (N_38477,N_34173,N_30841);
nand U38478 (N_38478,N_33199,N_30774);
nand U38479 (N_38479,N_30612,N_34131);
and U38480 (N_38480,N_30449,N_32524);
nor U38481 (N_38481,N_33521,N_33797);
nor U38482 (N_38482,N_34291,N_33491);
nand U38483 (N_38483,N_31784,N_34479);
xor U38484 (N_38484,N_34000,N_33357);
or U38485 (N_38485,N_33406,N_31117);
nor U38486 (N_38486,N_33813,N_33707);
and U38487 (N_38487,N_31322,N_30492);
and U38488 (N_38488,N_33993,N_33783);
xnor U38489 (N_38489,N_31807,N_33626);
and U38490 (N_38490,N_34539,N_30739);
nor U38491 (N_38491,N_31552,N_30540);
and U38492 (N_38492,N_33465,N_30015);
xnor U38493 (N_38493,N_31188,N_33747);
nor U38494 (N_38494,N_33806,N_34176);
or U38495 (N_38495,N_34569,N_32472);
or U38496 (N_38496,N_32784,N_32857);
nor U38497 (N_38497,N_31705,N_34837);
or U38498 (N_38498,N_33633,N_32947);
nor U38499 (N_38499,N_32137,N_31943);
xor U38500 (N_38500,N_34843,N_32616);
nor U38501 (N_38501,N_30870,N_31886);
and U38502 (N_38502,N_33792,N_32353);
and U38503 (N_38503,N_34042,N_33357);
nand U38504 (N_38504,N_34176,N_30943);
xor U38505 (N_38505,N_31266,N_33637);
xnor U38506 (N_38506,N_31289,N_33099);
or U38507 (N_38507,N_34433,N_34878);
xor U38508 (N_38508,N_32170,N_32724);
and U38509 (N_38509,N_34083,N_33182);
xnor U38510 (N_38510,N_33478,N_30878);
and U38511 (N_38511,N_32185,N_31248);
and U38512 (N_38512,N_34067,N_33868);
xnor U38513 (N_38513,N_32319,N_31462);
nor U38514 (N_38514,N_30877,N_33034);
nor U38515 (N_38515,N_30808,N_30298);
and U38516 (N_38516,N_34619,N_33581);
xor U38517 (N_38517,N_30030,N_34350);
xor U38518 (N_38518,N_32586,N_32537);
xor U38519 (N_38519,N_30060,N_32925);
and U38520 (N_38520,N_30816,N_33842);
or U38521 (N_38521,N_34363,N_32085);
nor U38522 (N_38522,N_34939,N_31883);
nor U38523 (N_38523,N_30975,N_31372);
or U38524 (N_38524,N_34113,N_34833);
nand U38525 (N_38525,N_31394,N_34366);
or U38526 (N_38526,N_34846,N_33021);
xnor U38527 (N_38527,N_31006,N_31061);
and U38528 (N_38528,N_34060,N_31946);
and U38529 (N_38529,N_30320,N_33285);
nand U38530 (N_38530,N_34956,N_31572);
nand U38531 (N_38531,N_30453,N_30295);
nor U38532 (N_38532,N_34398,N_30117);
nor U38533 (N_38533,N_32254,N_34497);
or U38534 (N_38534,N_31932,N_31926);
or U38535 (N_38535,N_34095,N_31389);
nand U38536 (N_38536,N_32290,N_31686);
nand U38537 (N_38537,N_30663,N_32697);
or U38538 (N_38538,N_31279,N_34388);
and U38539 (N_38539,N_33949,N_31876);
or U38540 (N_38540,N_30218,N_32975);
nand U38541 (N_38541,N_30883,N_30741);
nand U38542 (N_38542,N_30374,N_30892);
or U38543 (N_38543,N_30376,N_34653);
nand U38544 (N_38544,N_33631,N_31840);
or U38545 (N_38545,N_33293,N_31402);
and U38546 (N_38546,N_34936,N_30514);
and U38547 (N_38547,N_34816,N_34178);
nor U38548 (N_38548,N_32382,N_33031);
or U38549 (N_38549,N_34437,N_31623);
nor U38550 (N_38550,N_33347,N_31863);
or U38551 (N_38551,N_32506,N_31181);
and U38552 (N_38552,N_33181,N_30162);
or U38553 (N_38553,N_30906,N_34510);
xnor U38554 (N_38554,N_34049,N_31358);
xnor U38555 (N_38555,N_33862,N_33870);
or U38556 (N_38556,N_33616,N_31858);
nand U38557 (N_38557,N_33450,N_34900);
and U38558 (N_38558,N_34638,N_30912);
nand U38559 (N_38559,N_30752,N_34650);
nor U38560 (N_38560,N_34757,N_30064);
nor U38561 (N_38561,N_31147,N_33293);
nand U38562 (N_38562,N_34985,N_30010);
or U38563 (N_38563,N_31416,N_31939);
xor U38564 (N_38564,N_31493,N_33109);
and U38565 (N_38565,N_33691,N_34645);
nand U38566 (N_38566,N_34289,N_30001);
xnor U38567 (N_38567,N_32529,N_32990);
or U38568 (N_38568,N_34848,N_32301);
and U38569 (N_38569,N_30035,N_31540);
nor U38570 (N_38570,N_33256,N_32894);
nand U38571 (N_38571,N_30779,N_30941);
or U38572 (N_38572,N_32675,N_33953);
xor U38573 (N_38573,N_33465,N_34512);
or U38574 (N_38574,N_31160,N_31433);
or U38575 (N_38575,N_33504,N_34696);
xor U38576 (N_38576,N_32422,N_32527);
nand U38577 (N_38577,N_34849,N_33967);
xnor U38578 (N_38578,N_34060,N_31736);
or U38579 (N_38579,N_31920,N_30193);
nor U38580 (N_38580,N_33203,N_30988);
nand U38581 (N_38581,N_33565,N_30525);
nand U38582 (N_38582,N_34236,N_34992);
nand U38583 (N_38583,N_34339,N_33024);
xnor U38584 (N_38584,N_30693,N_30671);
nand U38585 (N_38585,N_32936,N_33196);
nor U38586 (N_38586,N_31415,N_33551);
or U38587 (N_38587,N_31426,N_31721);
or U38588 (N_38588,N_32909,N_32632);
and U38589 (N_38589,N_30691,N_31010);
or U38590 (N_38590,N_33023,N_31301);
and U38591 (N_38591,N_33358,N_31810);
nand U38592 (N_38592,N_32686,N_30879);
or U38593 (N_38593,N_31049,N_32180);
nor U38594 (N_38594,N_34177,N_31270);
or U38595 (N_38595,N_31347,N_31041);
xor U38596 (N_38596,N_34257,N_31119);
xor U38597 (N_38597,N_33984,N_31305);
nand U38598 (N_38598,N_32929,N_31245);
and U38599 (N_38599,N_31381,N_30716);
nor U38600 (N_38600,N_30486,N_30174);
nand U38601 (N_38601,N_30460,N_34039);
and U38602 (N_38602,N_30647,N_33363);
nor U38603 (N_38603,N_34642,N_30191);
nand U38604 (N_38604,N_30043,N_30421);
and U38605 (N_38605,N_30672,N_30150);
nand U38606 (N_38606,N_34031,N_32142);
nand U38607 (N_38607,N_32233,N_31955);
xnor U38608 (N_38608,N_32486,N_30593);
nand U38609 (N_38609,N_31663,N_31125);
nand U38610 (N_38610,N_30195,N_31494);
and U38611 (N_38611,N_33214,N_31947);
nand U38612 (N_38612,N_34758,N_34401);
nand U38613 (N_38613,N_33565,N_34679);
and U38614 (N_38614,N_31860,N_32407);
nor U38615 (N_38615,N_31546,N_33632);
and U38616 (N_38616,N_30073,N_31206);
or U38617 (N_38617,N_34056,N_32567);
nor U38618 (N_38618,N_30990,N_33583);
and U38619 (N_38619,N_34527,N_31524);
and U38620 (N_38620,N_32375,N_30215);
or U38621 (N_38621,N_33965,N_32029);
or U38622 (N_38622,N_30634,N_34886);
and U38623 (N_38623,N_31072,N_31579);
or U38624 (N_38624,N_30996,N_31122);
nor U38625 (N_38625,N_30401,N_31829);
xnor U38626 (N_38626,N_33605,N_32798);
xor U38627 (N_38627,N_31305,N_32399);
nor U38628 (N_38628,N_34499,N_31627);
nor U38629 (N_38629,N_34282,N_34991);
or U38630 (N_38630,N_31597,N_33922);
or U38631 (N_38631,N_32069,N_33374);
nor U38632 (N_38632,N_33297,N_31161);
nor U38633 (N_38633,N_32275,N_31408);
xor U38634 (N_38634,N_30259,N_32549);
xnor U38635 (N_38635,N_32368,N_34985);
xnor U38636 (N_38636,N_33091,N_33333);
nor U38637 (N_38637,N_30718,N_33322);
and U38638 (N_38638,N_31205,N_31701);
nand U38639 (N_38639,N_31011,N_32527);
nand U38640 (N_38640,N_32597,N_30450);
or U38641 (N_38641,N_31122,N_33544);
nand U38642 (N_38642,N_31905,N_34498);
nand U38643 (N_38643,N_32557,N_33965);
nand U38644 (N_38644,N_30929,N_32828);
and U38645 (N_38645,N_30220,N_31083);
nand U38646 (N_38646,N_32431,N_33371);
and U38647 (N_38647,N_30392,N_31143);
xnor U38648 (N_38648,N_32479,N_33760);
or U38649 (N_38649,N_32328,N_34190);
xnor U38650 (N_38650,N_32778,N_33652);
nand U38651 (N_38651,N_30066,N_32599);
nor U38652 (N_38652,N_34015,N_30080);
or U38653 (N_38653,N_32248,N_30861);
nor U38654 (N_38654,N_30441,N_32607);
nor U38655 (N_38655,N_31083,N_30882);
nand U38656 (N_38656,N_32816,N_30468);
xnor U38657 (N_38657,N_33735,N_31527);
and U38658 (N_38658,N_32241,N_31527);
nand U38659 (N_38659,N_33404,N_31705);
nor U38660 (N_38660,N_30312,N_33919);
nand U38661 (N_38661,N_33438,N_33683);
and U38662 (N_38662,N_34731,N_31945);
xnor U38663 (N_38663,N_33560,N_30384);
and U38664 (N_38664,N_30662,N_31307);
nand U38665 (N_38665,N_34399,N_33712);
nand U38666 (N_38666,N_30444,N_32344);
and U38667 (N_38667,N_34335,N_30525);
nor U38668 (N_38668,N_30025,N_30881);
nor U38669 (N_38669,N_31084,N_33790);
nor U38670 (N_38670,N_34925,N_32117);
nand U38671 (N_38671,N_30180,N_34879);
nor U38672 (N_38672,N_34085,N_34443);
nor U38673 (N_38673,N_31686,N_31688);
nand U38674 (N_38674,N_34310,N_31865);
nand U38675 (N_38675,N_31110,N_32720);
and U38676 (N_38676,N_34208,N_31678);
or U38677 (N_38677,N_34426,N_33559);
or U38678 (N_38678,N_34725,N_30354);
or U38679 (N_38679,N_32964,N_30129);
xor U38680 (N_38680,N_33485,N_31849);
nor U38681 (N_38681,N_30262,N_33510);
and U38682 (N_38682,N_32958,N_31199);
nand U38683 (N_38683,N_32741,N_31273);
nor U38684 (N_38684,N_33929,N_32626);
xor U38685 (N_38685,N_30014,N_30425);
or U38686 (N_38686,N_33246,N_32139);
xnor U38687 (N_38687,N_30250,N_34045);
xnor U38688 (N_38688,N_33037,N_34111);
xnor U38689 (N_38689,N_31460,N_30467);
or U38690 (N_38690,N_33072,N_34559);
or U38691 (N_38691,N_34659,N_32061);
xnor U38692 (N_38692,N_31626,N_30336);
nand U38693 (N_38693,N_31556,N_33354);
nand U38694 (N_38694,N_32988,N_32160);
nand U38695 (N_38695,N_30420,N_34647);
and U38696 (N_38696,N_33217,N_34676);
xnor U38697 (N_38697,N_30099,N_32666);
or U38698 (N_38698,N_33733,N_33636);
nor U38699 (N_38699,N_34690,N_34434);
and U38700 (N_38700,N_34274,N_31209);
and U38701 (N_38701,N_30616,N_33687);
xnor U38702 (N_38702,N_34572,N_30980);
nor U38703 (N_38703,N_31455,N_31982);
nor U38704 (N_38704,N_33735,N_34468);
nand U38705 (N_38705,N_31876,N_30609);
or U38706 (N_38706,N_31429,N_30923);
and U38707 (N_38707,N_30137,N_30607);
xor U38708 (N_38708,N_31592,N_33002);
xor U38709 (N_38709,N_33283,N_31558);
nor U38710 (N_38710,N_32457,N_34952);
nand U38711 (N_38711,N_33342,N_33446);
or U38712 (N_38712,N_32848,N_33363);
nand U38713 (N_38713,N_31131,N_31340);
and U38714 (N_38714,N_33612,N_32966);
nor U38715 (N_38715,N_33061,N_33751);
nor U38716 (N_38716,N_30684,N_34470);
xnor U38717 (N_38717,N_34217,N_33431);
nor U38718 (N_38718,N_32676,N_30274);
nand U38719 (N_38719,N_31467,N_32167);
nor U38720 (N_38720,N_31160,N_34659);
nor U38721 (N_38721,N_32133,N_30826);
nand U38722 (N_38722,N_33480,N_31567);
xor U38723 (N_38723,N_31650,N_33304);
nand U38724 (N_38724,N_34696,N_32233);
and U38725 (N_38725,N_34492,N_30866);
nand U38726 (N_38726,N_31311,N_34330);
and U38727 (N_38727,N_31127,N_34411);
nand U38728 (N_38728,N_32858,N_33339);
nand U38729 (N_38729,N_34482,N_31048);
and U38730 (N_38730,N_33530,N_33913);
nand U38731 (N_38731,N_30968,N_30842);
or U38732 (N_38732,N_32660,N_34654);
and U38733 (N_38733,N_31331,N_33027);
xor U38734 (N_38734,N_33231,N_34429);
nor U38735 (N_38735,N_30116,N_30315);
and U38736 (N_38736,N_33531,N_34273);
nand U38737 (N_38737,N_32818,N_31734);
nand U38738 (N_38738,N_34687,N_31727);
and U38739 (N_38739,N_32779,N_33045);
and U38740 (N_38740,N_30550,N_32141);
xnor U38741 (N_38741,N_34149,N_32330);
and U38742 (N_38742,N_33255,N_30649);
xor U38743 (N_38743,N_30629,N_34863);
or U38744 (N_38744,N_31107,N_30736);
xnor U38745 (N_38745,N_32582,N_30652);
xnor U38746 (N_38746,N_31101,N_30446);
or U38747 (N_38747,N_34533,N_33089);
and U38748 (N_38748,N_30208,N_30531);
nand U38749 (N_38749,N_31440,N_30900);
nor U38750 (N_38750,N_32010,N_34637);
nand U38751 (N_38751,N_30809,N_33001);
nor U38752 (N_38752,N_33184,N_33508);
and U38753 (N_38753,N_31876,N_31140);
nand U38754 (N_38754,N_30394,N_33272);
and U38755 (N_38755,N_30067,N_32821);
nor U38756 (N_38756,N_30003,N_30818);
nor U38757 (N_38757,N_32517,N_31247);
or U38758 (N_38758,N_33577,N_30426);
and U38759 (N_38759,N_33235,N_30904);
nor U38760 (N_38760,N_32377,N_31624);
nand U38761 (N_38761,N_31443,N_33731);
nor U38762 (N_38762,N_30807,N_30122);
nor U38763 (N_38763,N_33206,N_30119);
and U38764 (N_38764,N_30247,N_31300);
and U38765 (N_38765,N_30783,N_31240);
or U38766 (N_38766,N_31172,N_32860);
and U38767 (N_38767,N_33533,N_34266);
nor U38768 (N_38768,N_33519,N_32487);
or U38769 (N_38769,N_31930,N_32948);
and U38770 (N_38770,N_30023,N_30546);
and U38771 (N_38771,N_34204,N_33103);
or U38772 (N_38772,N_30286,N_33297);
and U38773 (N_38773,N_32197,N_31862);
or U38774 (N_38774,N_30719,N_30906);
or U38775 (N_38775,N_32076,N_34383);
or U38776 (N_38776,N_32343,N_34161);
nor U38777 (N_38777,N_31496,N_34066);
or U38778 (N_38778,N_34405,N_32021);
or U38779 (N_38779,N_33049,N_33142);
or U38780 (N_38780,N_33660,N_33412);
nand U38781 (N_38781,N_34672,N_31068);
nor U38782 (N_38782,N_34613,N_33952);
xnor U38783 (N_38783,N_34846,N_30410);
nor U38784 (N_38784,N_30945,N_32195);
xnor U38785 (N_38785,N_32698,N_34142);
and U38786 (N_38786,N_34400,N_31676);
nand U38787 (N_38787,N_33653,N_30497);
or U38788 (N_38788,N_33884,N_33545);
xnor U38789 (N_38789,N_30767,N_32293);
nand U38790 (N_38790,N_31375,N_34057);
or U38791 (N_38791,N_34769,N_31425);
nor U38792 (N_38792,N_31020,N_32253);
and U38793 (N_38793,N_33410,N_34297);
nor U38794 (N_38794,N_32898,N_34583);
and U38795 (N_38795,N_32685,N_34663);
or U38796 (N_38796,N_32772,N_31113);
nand U38797 (N_38797,N_31532,N_33989);
or U38798 (N_38798,N_33940,N_33134);
nand U38799 (N_38799,N_34962,N_34093);
nor U38800 (N_38800,N_33736,N_33380);
xnor U38801 (N_38801,N_33102,N_33804);
and U38802 (N_38802,N_31290,N_34318);
nand U38803 (N_38803,N_34130,N_33623);
or U38804 (N_38804,N_30462,N_31400);
or U38805 (N_38805,N_30403,N_33735);
or U38806 (N_38806,N_32945,N_32759);
nand U38807 (N_38807,N_33122,N_32755);
nand U38808 (N_38808,N_30123,N_31129);
and U38809 (N_38809,N_34108,N_30730);
or U38810 (N_38810,N_33960,N_30550);
nand U38811 (N_38811,N_32757,N_33152);
and U38812 (N_38812,N_32427,N_31748);
xnor U38813 (N_38813,N_31930,N_30831);
or U38814 (N_38814,N_33574,N_33851);
xnor U38815 (N_38815,N_31921,N_31710);
nor U38816 (N_38816,N_30936,N_31098);
nor U38817 (N_38817,N_30101,N_32840);
xnor U38818 (N_38818,N_33760,N_32137);
xor U38819 (N_38819,N_31974,N_33710);
or U38820 (N_38820,N_31092,N_31270);
nor U38821 (N_38821,N_30956,N_30203);
xor U38822 (N_38822,N_33139,N_33253);
or U38823 (N_38823,N_32712,N_33754);
or U38824 (N_38824,N_34075,N_30915);
nor U38825 (N_38825,N_33883,N_31880);
xnor U38826 (N_38826,N_34843,N_31561);
xor U38827 (N_38827,N_30726,N_34930);
and U38828 (N_38828,N_33286,N_34692);
or U38829 (N_38829,N_30334,N_32877);
nor U38830 (N_38830,N_31690,N_31797);
and U38831 (N_38831,N_31244,N_33870);
or U38832 (N_38832,N_32150,N_34026);
xor U38833 (N_38833,N_33115,N_30444);
and U38834 (N_38834,N_34796,N_32739);
xor U38835 (N_38835,N_31408,N_31906);
nand U38836 (N_38836,N_34628,N_32511);
xnor U38837 (N_38837,N_30267,N_31874);
and U38838 (N_38838,N_34220,N_33420);
or U38839 (N_38839,N_32526,N_32935);
xnor U38840 (N_38840,N_34341,N_30228);
and U38841 (N_38841,N_34358,N_34320);
and U38842 (N_38842,N_31323,N_34942);
nor U38843 (N_38843,N_30360,N_34302);
xnor U38844 (N_38844,N_33468,N_33167);
xnor U38845 (N_38845,N_31205,N_33343);
or U38846 (N_38846,N_32769,N_31052);
and U38847 (N_38847,N_31476,N_32514);
nand U38848 (N_38848,N_33674,N_32463);
nand U38849 (N_38849,N_34072,N_32253);
nor U38850 (N_38850,N_30895,N_34317);
and U38851 (N_38851,N_30253,N_33092);
nand U38852 (N_38852,N_32238,N_32038);
or U38853 (N_38853,N_34706,N_33757);
nor U38854 (N_38854,N_34022,N_34941);
nand U38855 (N_38855,N_32228,N_30914);
or U38856 (N_38856,N_30117,N_33186);
nor U38857 (N_38857,N_33125,N_32961);
nor U38858 (N_38858,N_34957,N_32396);
xor U38859 (N_38859,N_30986,N_33248);
and U38860 (N_38860,N_31482,N_31365);
xor U38861 (N_38861,N_34576,N_34183);
xnor U38862 (N_38862,N_33661,N_30504);
nor U38863 (N_38863,N_34968,N_30776);
xor U38864 (N_38864,N_33889,N_34663);
nor U38865 (N_38865,N_31733,N_34890);
and U38866 (N_38866,N_34103,N_33114);
nand U38867 (N_38867,N_31335,N_34982);
and U38868 (N_38868,N_32362,N_34351);
nor U38869 (N_38869,N_32397,N_30579);
or U38870 (N_38870,N_30940,N_30810);
nor U38871 (N_38871,N_30886,N_30804);
xor U38872 (N_38872,N_34539,N_34980);
and U38873 (N_38873,N_30206,N_30988);
or U38874 (N_38874,N_33377,N_31802);
nor U38875 (N_38875,N_32738,N_30410);
xor U38876 (N_38876,N_33605,N_32339);
xnor U38877 (N_38877,N_32283,N_32051);
and U38878 (N_38878,N_30159,N_30000);
or U38879 (N_38879,N_34056,N_30132);
nor U38880 (N_38880,N_33008,N_34855);
nor U38881 (N_38881,N_30204,N_30802);
and U38882 (N_38882,N_31075,N_30367);
and U38883 (N_38883,N_32963,N_30065);
nand U38884 (N_38884,N_34967,N_31504);
nor U38885 (N_38885,N_34402,N_31952);
nand U38886 (N_38886,N_34524,N_31071);
xor U38887 (N_38887,N_32026,N_33450);
nor U38888 (N_38888,N_33835,N_32919);
or U38889 (N_38889,N_31642,N_30200);
nand U38890 (N_38890,N_32119,N_30911);
xnor U38891 (N_38891,N_34481,N_31719);
nand U38892 (N_38892,N_31049,N_32111);
nand U38893 (N_38893,N_31185,N_34472);
or U38894 (N_38894,N_31401,N_30147);
nand U38895 (N_38895,N_34680,N_31964);
or U38896 (N_38896,N_34549,N_30942);
nor U38897 (N_38897,N_33136,N_30746);
nand U38898 (N_38898,N_33738,N_32980);
nor U38899 (N_38899,N_32601,N_30222);
nand U38900 (N_38900,N_32235,N_32876);
xor U38901 (N_38901,N_34913,N_34241);
nor U38902 (N_38902,N_34715,N_34409);
nor U38903 (N_38903,N_33520,N_31286);
xnor U38904 (N_38904,N_34804,N_34063);
xnor U38905 (N_38905,N_30965,N_31097);
xor U38906 (N_38906,N_33029,N_30197);
or U38907 (N_38907,N_33723,N_34330);
xnor U38908 (N_38908,N_30128,N_31142);
xor U38909 (N_38909,N_34448,N_32571);
nand U38910 (N_38910,N_31984,N_34364);
and U38911 (N_38911,N_33104,N_32004);
or U38912 (N_38912,N_30075,N_33983);
xnor U38913 (N_38913,N_32773,N_30865);
xor U38914 (N_38914,N_30135,N_31715);
or U38915 (N_38915,N_30804,N_31867);
nor U38916 (N_38916,N_33640,N_31324);
xnor U38917 (N_38917,N_34510,N_34100);
xnor U38918 (N_38918,N_32560,N_32013);
or U38919 (N_38919,N_34007,N_33118);
and U38920 (N_38920,N_34549,N_34208);
or U38921 (N_38921,N_30110,N_32774);
xnor U38922 (N_38922,N_32776,N_33734);
nor U38923 (N_38923,N_32490,N_32730);
nand U38924 (N_38924,N_33682,N_31458);
or U38925 (N_38925,N_34722,N_34501);
and U38926 (N_38926,N_30435,N_32855);
xnor U38927 (N_38927,N_34039,N_34414);
xor U38928 (N_38928,N_33133,N_30392);
and U38929 (N_38929,N_31327,N_32438);
or U38930 (N_38930,N_30883,N_30702);
nand U38931 (N_38931,N_33356,N_32473);
nand U38932 (N_38932,N_31996,N_33346);
xnor U38933 (N_38933,N_30632,N_30950);
and U38934 (N_38934,N_34961,N_30423);
nand U38935 (N_38935,N_32908,N_30954);
nand U38936 (N_38936,N_30394,N_34506);
or U38937 (N_38937,N_32538,N_33884);
nor U38938 (N_38938,N_31578,N_30302);
nand U38939 (N_38939,N_34156,N_32218);
or U38940 (N_38940,N_33952,N_31598);
and U38941 (N_38941,N_33453,N_32096);
nor U38942 (N_38942,N_31350,N_34261);
nor U38943 (N_38943,N_34853,N_31499);
and U38944 (N_38944,N_30900,N_33002);
or U38945 (N_38945,N_32828,N_30447);
or U38946 (N_38946,N_32977,N_31218);
and U38947 (N_38947,N_34406,N_33246);
nand U38948 (N_38948,N_31516,N_33574);
nand U38949 (N_38949,N_30314,N_33274);
and U38950 (N_38950,N_34345,N_34234);
nor U38951 (N_38951,N_30007,N_31958);
nand U38952 (N_38952,N_33022,N_32539);
nand U38953 (N_38953,N_33680,N_31157);
or U38954 (N_38954,N_32003,N_32144);
xor U38955 (N_38955,N_30678,N_31484);
and U38956 (N_38956,N_33058,N_34293);
and U38957 (N_38957,N_32541,N_32438);
and U38958 (N_38958,N_30907,N_34689);
xnor U38959 (N_38959,N_32159,N_32766);
nor U38960 (N_38960,N_30224,N_31375);
and U38961 (N_38961,N_32584,N_33310);
nor U38962 (N_38962,N_31766,N_31425);
nor U38963 (N_38963,N_33849,N_32906);
nor U38964 (N_38964,N_34287,N_32082);
nor U38965 (N_38965,N_34621,N_34834);
xnor U38966 (N_38966,N_33217,N_32019);
and U38967 (N_38967,N_32572,N_31112);
nor U38968 (N_38968,N_30423,N_30822);
or U38969 (N_38969,N_31675,N_31942);
or U38970 (N_38970,N_33138,N_33455);
nor U38971 (N_38971,N_31801,N_32468);
and U38972 (N_38972,N_31024,N_33585);
xnor U38973 (N_38973,N_31540,N_34792);
xnor U38974 (N_38974,N_33158,N_32616);
nor U38975 (N_38975,N_32949,N_34632);
nor U38976 (N_38976,N_32693,N_31518);
nand U38977 (N_38977,N_34395,N_34723);
and U38978 (N_38978,N_33869,N_32197);
or U38979 (N_38979,N_30668,N_31629);
and U38980 (N_38980,N_30391,N_34331);
xnor U38981 (N_38981,N_31645,N_32193);
or U38982 (N_38982,N_34374,N_34500);
nor U38983 (N_38983,N_31779,N_34285);
nand U38984 (N_38984,N_30712,N_30321);
and U38985 (N_38985,N_31265,N_32581);
xor U38986 (N_38986,N_34023,N_30237);
nor U38987 (N_38987,N_33835,N_31234);
and U38988 (N_38988,N_31766,N_33748);
nand U38989 (N_38989,N_33053,N_31253);
xor U38990 (N_38990,N_34491,N_34549);
xnor U38991 (N_38991,N_30797,N_33019);
nor U38992 (N_38992,N_31125,N_34548);
or U38993 (N_38993,N_30886,N_31396);
and U38994 (N_38994,N_31340,N_34054);
nor U38995 (N_38995,N_33868,N_33041);
nand U38996 (N_38996,N_31436,N_31391);
or U38997 (N_38997,N_34364,N_32876);
and U38998 (N_38998,N_32043,N_30430);
and U38999 (N_38999,N_30329,N_30421);
and U39000 (N_39000,N_31483,N_34176);
or U39001 (N_39001,N_34330,N_33484);
xnor U39002 (N_39002,N_31759,N_34410);
xnor U39003 (N_39003,N_30126,N_30970);
or U39004 (N_39004,N_33453,N_34837);
or U39005 (N_39005,N_32911,N_32283);
and U39006 (N_39006,N_33186,N_30202);
xnor U39007 (N_39007,N_32514,N_30761);
nand U39008 (N_39008,N_33726,N_30939);
or U39009 (N_39009,N_31750,N_30456);
nor U39010 (N_39010,N_30736,N_30726);
nand U39011 (N_39011,N_31616,N_31748);
nor U39012 (N_39012,N_34570,N_31444);
nand U39013 (N_39013,N_31946,N_34978);
or U39014 (N_39014,N_32310,N_30345);
and U39015 (N_39015,N_32048,N_32400);
xnor U39016 (N_39016,N_30118,N_33861);
nor U39017 (N_39017,N_32594,N_32760);
xnor U39018 (N_39018,N_34197,N_33008);
or U39019 (N_39019,N_33366,N_32796);
nor U39020 (N_39020,N_31713,N_32172);
or U39021 (N_39021,N_32629,N_30690);
xor U39022 (N_39022,N_32828,N_31788);
nor U39023 (N_39023,N_30687,N_34424);
or U39024 (N_39024,N_33309,N_30144);
xnor U39025 (N_39025,N_30690,N_30256);
and U39026 (N_39026,N_32079,N_30644);
or U39027 (N_39027,N_33838,N_31001);
and U39028 (N_39028,N_30860,N_32848);
nor U39029 (N_39029,N_34705,N_31000);
or U39030 (N_39030,N_33761,N_33258);
nor U39031 (N_39031,N_32809,N_33860);
nor U39032 (N_39032,N_34194,N_34517);
nor U39033 (N_39033,N_30949,N_34261);
or U39034 (N_39034,N_34659,N_31097);
or U39035 (N_39035,N_33413,N_34889);
nand U39036 (N_39036,N_31778,N_30111);
xnor U39037 (N_39037,N_33256,N_31678);
nor U39038 (N_39038,N_31575,N_31657);
or U39039 (N_39039,N_32045,N_34689);
and U39040 (N_39040,N_32773,N_32248);
and U39041 (N_39041,N_31156,N_32761);
xnor U39042 (N_39042,N_34533,N_30820);
or U39043 (N_39043,N_31881,N_34877);
or U39044 (N_39044,N_33156,N_33293);
or U39045 (N_39045,N_33859,N_31499);
nor U39046 (N_39046,N_31549,N_34158);
xnor U39047 (N_39047,N_31132,N_34127);
nor U39048 (N_39048,N_32729,N_31284);
nor U39049 (N_39049,N_30763,N_34980);
nand U39050 (N_39050,N_33265,N_32260);
or U39051 (N_39051,N_30871,N_33822);
and U39052 (N_39052,N_32383,N_32269);
nand U39053 (N_39053,N_32260,N_34833);
xnor U39054 (N_39054,N_33890,N_33244);
nand U39055 (N_39055,N_31617,N_34508);
xnor U39056 (N_39056,N_34172,N_32902);
nor U39057 (N_39057,N_33842,N_33071);
or U39058 (N_39058,N_34006,N_34651);
xor U39059 (N_39059,N_31823,N_33631);
and U39060 (N_39060,N_33171,N_34244);
and U39061 (N_39061,N_32675,N_30243);
nor U39062 (N_39062,N_30433,N_34165);
nand U39063 (N_39063,N_32463,N_32545);
xor U39064 (N_39064,N_31531,N_34521);
and U39065 (N_39065,N_34866,N_30547);
nand U39066 (N_39066,N_34458,N_31966);
or U39067 (N_39067,N_32952,N_33816);
nand U39068 (N_39068,N_32215,N_30728);
nor U39069 (N_39069,N_30677,N_32931);
or U39070 (N_39070,N_30340,N_30977);
or U39071 (N_39071,N_33629,N_32123);
or U39072 (N_39072,N_31033,N_34856);
nor U39073 (N_39073,N_31201,N_31786);
xor U39074 (N_39074,N_31133,N_32865);
xor U39075 (N_39075,N_32504,N_33294);
nand U39076 (N_39076,N_33854,N_33493);
or U39077 (N_39077,N_31274,N_32971);
nor U39078 (N_39078,N_34581,N_30326);
or U39079 (N_39079,N_33601,N_32314);
xor U39080 (N_39080,N_33085,N_33858);
nand U39081 (N_39081,N_30095,N_31033);
and U39082 (N_39082,N_30031,N_31726);
and U39083 (N_39083,N_34664,N_33605);
or U39084 (N_39084,N_30325,N_34777);
and U39085 (N_39085,N_34635,N_31117);
or U39086 (N_39086,N_30576,N_34826);
and U39087 (N_39087,N_34890,N_33680);
nor U39088 (N_39088,N_31729,N_30278);
and U39089 (N_39089,N_32240,N_32464);
and U39090 (N_39090,N_31954,N_31812);
nor U39091 (N_39091,N_30417,N_31729);
nand U39092 (N_39092,N_33983,N_34567);
xnor U39093 (N_39093,N_30456,N_30693);
nor U39094 (N_39094,N_34511,N_34420);
xnor U39095 (N_39095,N_30596,N_30297);
or U39096 (N_39096,N_30723,N_30810);
or U39097 (N_39097,N_30280,N_32935);
nor U39098 (N_39098,N_33553,N_32230);
or U39099 (N_39099,N_33007,N_30068);
xnor U39100 (N_39100,N_32475,N_31927);
or U39101 (N_39101,N_33438,N_30502);
and U39102 (N_39102,N_31979,N_30615);
and U39103 (N_39103,N_34561,N_32364);
and U39104 (N_39104,N_33381,N_32431);
xnor U39105 (N_39105,N_33162,N_34343);
xnor U39106 (N_39106,N_34695,N_34561);
and U39107 (N_39107,N_33207,N_31534);
nand U39108 (N_39108,N_33080,N_33130);
and U39109 (N_39109,N_34951,N_33314);
or U39110 (N_39110,N_32097,N_30140);
and U39111 (N_39111,N_34499,N_32909);
xor U39112 (N_39112,N_34644,N_33441);
nor U39113 (N_39113,N_30741,N_32296);
and U39114 (N_39114,N_32248,N_30233);
or U39115 (N_39115,N_32428,N_30691);
and U39116 (N_39116,N_33744,N_31295);
and U39117 (N_39117,N_32299,N_32544);
and U39118 (N_39118,N_32773,N_30171);
nor U39119 (N_39119,N_30778,N_30834);
nor U39120 (N_39120,N_34460,N_32816);
xnor U39121 (N_39121,N_30124,N_33313);
or U39122 (N_39122,N_32092,N_33870);
xor U39123 (N_39123,N_31530,N_32608);
and U39124 (N_39124,N_30839,N_34666);
and U39125 (N_39125,N_33948,N_34338);
nand U39126 (N_39126,N_30590,N_30163);
or U39127 (N_39127,N_33334,N_33303);
and U39128 (N_39128,N_33659,N_30514);
nor U39129 (N_39129,N_32854,N_30308);
or U39130 (N_39130,N_31420,N_31203);
nand U39131 (N_39131,N_34278,N_32772);
nand U39132 (N_39132,N_30178,N_34797);
or U39133 (N_39133,N_30657,N_34642);
nand U39134 (N_39134,N_31330,N_33094);
or U39135 (N_39135,N_32547,N_34206);
nor U39136 (N_39136,N_34149,N_31811);
xnor U39137 (N_39137,N_30490,N_34472);
or U39138 (N_39138,N_33827,N_33524);
xnor U39139 (N_39139,N_31907,N_31175);
or U39140 (N_39140,N_33218,N_33819);
and U39141 (N_39141,N_33251,N_34990);
or U39142 (N_39142,N_30407,N_30564);
or U39143 (N_39143,N_34048,N_30997);
nand U39144 (N_39144,N_34169,N_30272);
nand U39145 (N_39145,N_30943,N_31730);
or U39146 (N_39146,N_31344,N_32549);
xor U39147 (N_39147,N_32853,N_34332);
nand U39148 (N_39148,N_32686,N_31083);
or U39149 (N_39149,N_30091,N_32602);
or U39150 (N_39150,N_32778,N_34770);
and U39151 (N_39151,N_32139,N_32830);
xnor U39152 (N_39152,N_34405,N_31084);
nor U39153 (N_39153,N_33030,N_31601);
nor U39154 (N_39154,N_31251,N_32990);
and U39155 (N_39155,N_30415,N_34885);
or U39156 (N_39156,N_30289,N_31305);
nor U39157 (N_39157,N_30143,N_34914);
and U39158 (N_39158,N_32117,N_34142);
nand U39159 (N_39159,N_34177,N_33617);
or U39160 (N_39160,N_34511,N_34539);
xnor U39161 (N_39161,N_32976,N_33130);
and U39162 (N_39162,N_32553,N_31563);
xor U39163 (N_39163,N_33629,N_30833);
or U39164 (N_39164,N_33623,N_30214);
and U39165 (N_39165,N_34584,N_31766);
xnor U39166 (N_39166,N_34082,N_33584);
or U39167 (N_39167,N_33617,N_32565);
and U39168 (N_39168,N_31418,N_32930);
and U39169 (N_39169,N_31707,N_32508);
nand U39170 (N_39170,N_32108,N_31950);
or U39171 (N_39171,N_34438,N_34249);
and U39172 (N_39172,N_31174,N_32171);
and U39173 (N_39173,N_33524,N_32587);
or U39174 (N_39174,N_31805,N_34919);
and U39175 (N_39175,N_31526,N_33470);
or U39176 (N_39176,N_32927,N_33581);
nand U39177 (N_39177,N_30884,N_30021);
and U39178 (N_39178,N_31429,N_33147);
nor U39179 (N_39179,N_31351,N_33813);
nand U39180 (N_39180,N_33936,N_33391);
xnor U39181 (N_39181,N_32752,N_31494);
or U39182 (N_39182,N_32546,N_33739);
and U39183 (N_39183,N_32820,N_31010);
and U39184 (N_39184,N_31516,N_34406);
nand U39185 (N_39185,N_33514,N_33981);
xnor U39186 (N_39186,N_31999,N_31031);
and U39187 (N_39187,N_34162,N_30593);
or U39188 (N_39188,N_31728,N_30020);
and U39189 (N_39189,N_31305,N_32771);
nand U39190 (N_39190,N_31902,N_31132);
nand U39191 (N_39191,N_30438,N_31871);
nand U39192 (N_39192,N_31380,N_31471);
nor U39193 (N_39193,N_34327,N_33405);
xor U39194 (N_39194,N_32638,N_33517);
or U39195 (N_39195,N_31071,N_33303);
xnor U39196 (N_39196,N_30542,N_31760);
xnor U39197 (N_39197,N_30554,N_31303);
nor U39198 (N_39198,N_30745,N_30137);
xor U39199 (N_39199,N_33022,N_30384);
xnor U39200 (N_39200,N_34870,N_33067);
and U39201 (N_39201,N_33419,N_31749);
nor U39202 (N_39202,N_33564,N_30345);
or U39203 (N_39203,N_34497,N_31035);
xnor U39204 (N_39204,N_32625,N_32519);
xor U39205 (N_39205,N_33284,N_30001);
or U39206 (N_39206,N_34290,N_32899);
nor U39207 (N_39207,N_32187,N_31215);
nand U39208 (N_39208,N_31720,N_32345);
nand U39209 (N_39209,N_32555,N_31243);
and U39210 (N_39210,N_33827,N_34147);
xor U39211 (N_39211,N_32667,N_34660);
nor U39212 (N_39212,N_31233,N_31227);
and U39213 (N_39213,N_31225,N_31003);
and U39214 (N_39214,N_30787,N_34063);
or U39215 (N_39215,N_31954,N_31343);
or U39216 (N_39216,N_30491,N_33789);
nor U39217 (N_39217,N_31444,N_31949);
or U39218 (N_39218,N_32411,N_33741);
or U39219 (N_39219,N_31965,N_31037);
and U39220 (N_39220,N_32266,N_34808);
nor U39221 (N_39221,N_32518,N_30336);
nor U39222 (N_39222,N_31299,N_34990);
nand U39223 (N_39223,N_33529,N_34934);
or U39224 (N_39224,N_33328,N_34185);
nor U39225 (N_39225,N_33591,N_34545);
nor U39226 (N_39226,N_31922,N_30532);
xnor U39227 (N_39227,N_32839,N_32280);
nor U39228 (N_39228,N_30867,N_33537);
or U39229 (N_39229,N_31031,N_31471);
nand U39230 (N_39230,N_31513,N_30636);
or U39231 (N_39231,N_31418,N_30927);
xor U39232 (N_39232,N_30722,N_30700);
or U39233 (N_39233,N_32512,N_34208);
xor U39234 (N_39234,N_34056,N_34114);
or U39235 (N_39235,N_31615,N_34238);
nor U39236 (N_39236,N_33255,N_32526);
or U39237 (N_39237,N_33379,N_32145);
xnor U39238 (N_39238,N_32373,N_31601);
or U39239 (N_39239,N_33047,N_34774);
and U39240 (N_39240,N_32577,N_34153);
and U39241 (N_39241,N_34933,N_30798);
nand U39242 (N_39242,N_30821,N_30116);
or U39243 (N_39243,N_32818,N_32354);
xor U39244 (N_39244,N_31264,N_32755);
nor U39245 (N_39245,N_33538,N_31551);
xor U39246 (N_39246,N_30024,N_34494);
nor U39247 (N_39247,N_32458,N_31786);
or U39248 (N_39248,N_33250,N_30453);
xor U39249 (N_39249,N_30068,N_32439);
and U39250 (N_39250,N_32975,N_31584);
or U39251 (N_39251,N_34571,N_31243);
nand U39252 (N_39252,N_34614,N_34629);
and U39253 (N_39253,N_34665,N_32263);
or U39254 (N_39254,N_34260,N_33667);
nor U39255 (N_39255,N_33730,N_34679);
or U39256 (N_39256,N_32908,N_31911);
nor U39257 (N_39257,N_30888,N_30755);
nor U39258 (N_39258,N_30934,N_34149);
xor U39259 (N_39259,N_32720,N_33340);
or U39260 (N_39260,N_34737,N_32292);
nor U39261 (N_39261,N_32419,N_30897);
or U39262 (N_39262,N_31497,N_31635);
nand U39263 (N_39263,N_30480,N_30069);
or U39264 (N_39264,N_33248,N_30727);
or U39265 (N_39265,N_32015,N_30212);
and U39266 (N_39266,N_30928,N_34212);
and U39267 (N_39267,N_31315,N_31278);
or U39268 (N_39268,N_31705,N_31222);
and U39269 (N_39269,N_33447,N_32336);
or U39270 (N_39270,N_32494,N_31434);
or U39271 (N_39271,N_31263,N_30554);
or U39272 (N_39272,N_33286,N_32623);
nand U39273 (N_39273,N_31398,N_31663);
nor U39274 (N_39274,N_30193,N_34953);
or U39275 (N_39275,N_33443,N_31123);
nor U39276 (N_39276,N_33318,N_33207);
nand U39277 (N_39277,N_30277,N_30327);
nor U39278 (N_39278,N_31223,N_30070);
nand U39279 (N_39279,N_32911,N_33196);
nand U39280 (N_39280,N_31593,N_31190);
and U39281 (N_39281,N_33298,N_31638);
or U39282 (N_39282,N_31295,N_33121);
or U39283 (N_39283,N_31174,N_34428);
and U39284 (N_39284,N_33663,N_32983);
xnor U39285 (N_39285,N_33016,N_33009);
nor U39286 (N_39286,N_31755,N_34413);
or U39287 (N_39287,N_32224,N_30727);
and U39288 (N_39288,N_34042,N_30054);
nand U39289 (N_39289,N_33255,N_31141);
or U39290 (N_39290,N_33717,N_31255);
nor U39291 (N_39291,N_33069,N_32530);
nor U39292 (N_39292,N_31495,N_33433);
and U39293 (N_39293,N_30890,N_33938);
nand U39294 (N_39294,N_33213,N_32046);
nand U39295 (N_39295,N_31586,N_34119);
xor U39296 (N_39296,N_33681,N_31191);
xnor U39297 (N_39297,N_32508,N_33367);
and U39298 (N_39298,N_33903,N_33795);
or U39299 (N_39299,N_31883,N_33880);
or U39300 (N_39300,N_34201,N_31683);
or U39301 (N_39301,N_34539,N_32076);
or U39302 (N_39302,N_31489,N_32753);
nand U39303 (N_39303,N_31409,N_32478);
or U39304 (N_39304,N_31057,N_34310);
nor U39305 (N_39305,N_32807,N_30599);
nand U39306 (N_39306,N_30347,N_30176);
xnor U39307 (N_39307,N_34960,N_31669);
nor U39308 (N_39308,N_30852,N_34631);
xor U39309 (N_39309,N_34559,N_34271);
or U39310 (N_39310,N_32850,N_31511);
xnor U39311 (N_39311,N_34294,N_32673);
xor U39312 (N_39312,N_31880,N_32292);
nand U39313 (N_39313,N_30042,N_30827);
nor U39314 (N_39314,N_33267,N_32409);
or U39315 (N_39315,N_33273,N_34193);
and U39316 (N_39316,N_32158,N_34102);
and U39317 (N_39317,N_32043,N_31261);
nand U39318 (N_39318,N_30886,N_31280);
or U39319 (N_39319,N_34957,N_33075);
nor U39320 (N_39320,N_32019,N_34753);
nand U39321 (N_39321,N_32093,N_33694);
nand U39322 (N_39322,N_34738,N_32148);
or U39323 (N_39323,N_31519,N_31904);
and U39324 (N_39324,N_34528,N_34450);
nor U39325 (N_39325,N_32667,N_33942);
xor U39326 (N_39326,N_33715,N_32265);
and U39327 (N_39327,N_30824,N_33125);
or U39328 (N_39328,N_31931,N_31773);
nand U39329 (N_39329,N_34416,N_33168);
xor U39330 (N_39330,N_32950,N_34028);
and U39331 (N_39331,N_34945,N_30149);
and U39332 (N_39332,N_34435,N_33869);
xor U39333 (N_39333,N_31545,N_34170);
nor U39334 (N_39334,N_34798,N_34782);
and U39335 (N_39335,N_34225,N_32606);
or U39336 (N_39336,N_33544,N_33860);
and U39337 (N_39337,N_30985,N_31308);
nand U39338 (N_39338,N_33675,N_33023);
and U39339 (N_39339,N_30877,N_31193);
and U39340 (N_39340,N_31734,N_31706);
nand U39341 (N_39341,N_32435,N_30059);
xnor U39342 (N_39342,N_32930,N_32622);
xor U39343 (N_39343,N_30652,N_32203);
xnor U39344 (N_39344,N_30940,N_34518);
nand U39345 (N_39345,N_31545,N_31043);
nor U39346 (N_39346,N_30145,N_30355);
xor U39347 (N_39347,N_33722,N_33974);
nor U39348 (N_39348,N_31973,N_32602);
and U39349 (N_39349,N_32533,N_30528);
nand U39350 (N_39350,N_34052,N_30580);
nand U39351 (N_39351,N_33206,N_33663);
and U39352 (N_39352,N_34005,N_30162);
xnor U39353 (N_39353,N_32776,N_31727);
xnor U39354 (N_39354,N_32485,N_34621);
nand U39355 (N_39355,N_31553,N_31781);
nor U39356 (N_39356,N_30199,N_33816);
xor U39357 (N_39357,N_30956,N_33184);
or U39358 (N_39358,N_32712,N_31524);
and U39359 (N_39359,N_31510,N_31296);
nor U39360 (N_39360,N_33024,N_34596);
and U39361 (N_39361,N_32663,N_32139);
nand U39362 (N_39362,N_34758,N_31495);
nor U39363 (N_39363,N_34450,N_31005);
xnor U39364 (N_39364,N_31756,N_33485);
xnor U39365 (N_39365,N_34400,N_31458);
nor U39366 (N_39366,N_33210,N_33903);
or U39367 (N_39367,N_30004,N_31479);
nand U39368 (N_39368,N_31893,N_33010);
and U39369 (N_39369,N_33521,N_32858);
and U39370 (N_39370,N_30056,N_34056);
and U39371 (N_39371,N_31239,N_33480);
nor U39372 (N_39372,N_30429,N_34009);
or U39373 (N_39373,N_30198,N_31464);
nor U39374 (N_39374,N_32388,N_33006);
xor U39375 (N_39375,N_30136,N_30809);
xnor U39376 (N_39376,N_34250,N_32635);
or U39377 (N_39377,N_33919,N_34185);
nand U39378 (N_39378,N_31028,N_32941);
nor U39379 (N_39379,N_33086,N_30769);
nor U39380 (N_39380,N_33250,N_30130);
or U39381 (N_39381,N_31482,N_31371);
nor U39382 (N_39382,N_34413,N_34324);
and U39383 (N_39383,N_33398,N_33766);
nor U39384 (N_39384,N_32410,N_30161);
and U39385 (N_39385,N_33590,N_32348);
nor U39386 (N_39386,N_33440,N_34964);
nor U39387 (N_39387,N_34313,N_30589);
xnor U39388 (N_39388,N_33786,N_30010);
or U39389 (N_39389,N_33548,N_31552);
or U39390 (N_39390,N_32540,N_32362);
nor U39391 (N_39391,N_31116,N_30694);
or U39392 (N_39392,N_30867,N_31593);
nand U39393 (N_39393,N_30714,N_33480);
nand U39394 (N_39394,N_32753,N_31010);
xor U39395 (N_39395,N_33221,N_31147);
nand U39396 (N_39396,N_31918,N_32780);
nor U39397 (N_39397,N_34628,N_31971);
or U39398 (N_39398,N_34229,N_30707);
or U39399 (N_39399,N_31148,N_32744);
nor U39400 (N_39400,N_31043,N_33000);
or U39401 (N_39401,N_32887,N_33675);
and U39402 (N_39402,N_33889,N_32269);
or U39403 (N_39403,N_30891,N_30030);
and U39404 (N_39404,N_34644,N_34851);
nand U39405 (N_39405,N_32036,N_33994);
and U39406 (N_39406,N_34463,N_34989);
xor U39407 (N_39407,N_31073,N_31400);
nor U39408 (N_39408,N_32839,N_34213);
xor U39409 (N_39409,N_33600,N_30141);
xor U39410 (N_39410,N_30089,N_33868);
xor U39411 (N_39411,N_30430,N_32646);
nor U39412 (N_39412,N_33646,N_32937);
nand U39413 (N_39413,N_34391,N_34385);
xor U39414 (N_39414,N_30956,N_32221);
xor U39415 (N_39415,N_30327,N_34087);
or U39416 (N_39416,N_33911,N_30422);
nand U39417 (N_39417,N_30283,N_33645);
nor U39418 (N_39418,N_32122,N_31426);
or U39419 (N_39419,N_30732,N_32917);
xnor U39420 (N_39420,N_33467,N_31329);
nand U39421 (N_39421,N_31279,N_32970);
xnor U39422 (N_39422,N_34054,N_34487);
xnor U39423 (N_39423,N_34466,N_30548);
xnor U39424 (N_39424,N_30015,N_33021);
or U39425 (N_39425,N_34436,N_32070);
and U39426 (N_39426,N_30664,N_32090);
nor U39427 (N_39427,N_32424,N_32135);
and U39428 (N_39428,N_33961,N_30689);
nand U39429 (N_39429,N_33698,N_34120);
or U39430 (N_39430,N_30295,N_33055);
and U39431 (N_39431,N_30479,N_33955);
xnor U39432 (N_39432,N_34442,N_33347);
nor U39433 (N_39433,N_32662,N_33338);
or U39434 (N_39434,N_34436,N_34618);
xor U39435 (N_39435,N_31208,N_31030);
nor U39436 (N_39436,N_31674,N_32481);
nand U39437 (N_39437,N_30875,N_34430);
or U39438 (N_39438,N_31308,N_32634);
or U39439 (N_39439,N_34728,N_31541);
nor U39440 (N_39440,N_31686,N_34862);
xor U39441 (N_39441,N_34790,N_31114);
nand U39442 (N_39442,N_30097,N_31057);
or U39443 (N_39443,N_31259,N_32639);
xor U39444 (N_39444,N_32969,N_32033);
nor U39445 (N_39445,N_32963,N_34083);
xnor U39446 (N_39446,N_33652,N_32373);
xor U39447 (N_39447,N_31436,N_33666);
and U39448 (N_39448,N_30712,N_33799);
nor U39449 (N_39449,N_34448,N_34504);
xor U39450 (N_39450,N_31448,N_30524);
nor U39451 (N_39451,N_31428,N_30397);
and U39452 (N_39452,N_34699,N_32288);
nor U39453 (N_39453,N_30456,N_34394);
or U39454 (N_39454,N_33425,N_31074);
xnor U39455 (N_39455,N_31414,N_32433);
nand U39456 (N_39456,N_34397,N_32357);
nand U39457 (N_39457,N_34548,N_32629);
xor U39458 (N_39458,N_32781,N_31754);
nand U39459 (N_39459,N_32664,N_30366);
xnor U39460 (N_39460,N_31912,N_32297);
nor U39461 (N_39461,N_32391,N_31473);
xnor U39462 (N_39462,N_34081,N_33901);
nor U39463 (N_39463,N_31249,N_31292);
nor U39464 (N_39464,N_31047,N_33077);
nor U39465 (N_39465,N_30045,N_31503);
nand U39466 (N_39466,N_30722,N_34866);
nor U39467 (N_39467,N_31029,N_32125);
nand U39468 (N_39468,N_30800,N_30335);
xor U39469 (N_39469,N_30995,N_34624);
or U39470 (N_39470,N_32492,N_30788);
xnor U39471 (N_39471,N_32605,N_34385);
or U39472 (N_39472,N_32760,N_30014);
xor U39473 (N_39473,N_30727,N_32465);
nand U39474 (N_39474,N_33695,N_34240);
xnor U39475 (N_39475,N_34371,N_33868);
or U39476 (N_39476,N_31803,N_32072);
xnor U39477 (N_39477,N_34923,N_31214);
nand U39478 (N_39478,N_31734,N_32846);
nor U39479 (N_39479,N_32241,N_32668);
nand U39480 (N_39480,N_32368,N_33672);
nand U39481 (N_39481,N_32505,N_32971);
xnor U39482 (N_39482,N_33567,N_32567);
nand U39483 (N_39483,N_31696,N_31472);
xnor U39484 (N_39484,N_31156,N_33175);
and U39485 (N_39485,N_30169,N_33197);
or U39486 (N_39486,N_33116,N_33851);
xnor U39487 (N_39487,N_33078,N_34767);
nand U39488 (N_39488,N_32368,N_33853);
xnor U39489 (N_39489,N_30438,N_30403);
xor U39490 (N_39490,N_30924,N_31030);
or U39491 (N_39491,N_32174,N_33192);
xnor U39492 (N_39492,N_31725,N_34007);
nor U39493 (N_39493,N_33457,N_32880);
nor U39494 (N_39494,N_33195,N_32883);
or U39495 (N_39495,N_34819,N_31738);
xor U39496 (N_39496,N_32398,N_32183);
and U39497 (N_39497,N_33663,N_33452);
nand U39498 (N_39498,N_32546,N_32139);
and U39499 (N_39499,N_30226,N_33127);
and U39500 (N_39500,N_30356,N_33414);
and U39501 (N_39501,N_34275,N_34277);
xor U39502 (N_39502,N_32509,N_33640);
and U39503 (N_39503,N_32530,N_33946);
nor U39504 (N_39504,N_33636,N_34449);
and U39505 (N_39505,N_32287,N_33336);
xnor U39506 (N_39506,N_33100,N_34061);
or U39507 (N_39507,N_30681,N_31064);
nor U39508 (N_39508,N_33913,N_31478);
or U39509 (N_39509,N_30063,N_34002);
nor U39510 (N_39510,N_30939,N_32613);
and U39511 (N_39511,N_31556,N_31999);
nand U39512 (N_39512,N_34466,N_32856);
nand U39513 (N_39513,N_31971,N_33649);
xnor U39514 (N_39514,N_33657,N_34364);
or U39515 (N_39515,N_31835,N_30575);
and U39516 (N_39516,N_34111,N_30427);
and U39517 (N_39517,N_31828,N_30467);
and U39518 (N_39518,N_30421,N_30412);
nor U39519 (N_39519,N_30046,N_33552);
or U39520 (N_39520,N_30435,N_34953);
or U39521 (N_39521,N_32017,N_31794);
or U39522 (N_39522,N_34076,N_34492);
nand U39523 (N_39523,N_30560,N_33695);
xor U39524 (N_39524,N_33144,N_32508);
and U39525 (N_39525,N_33531,N_33869);
and U39526 (N_39526,N_31190,N_30662);
xnor U39527 (N_39527,N_31975,N_30014);
xor U39528 (N_39528,N_32146,N_30984);
xnor U39529 (N_39529,N_34488,N_34710);
nor U39530 (N_39530,N_33396,N_33952);
and U39531 (N_39531,N_33067,N_34571);
or U39532 (N_39532,N_33445,N_31042);
nand U39533 (N_39533,N_31604,N_34281);
and U39534 (N_39534,N_34027,N_32330);
nor U39535 (N_39535,N_33844,N_33568);
nand U39536 (N_39536,N_30817,N_31552);
nand U39537 (N_39537,N_32550,N_34730);
or U39538 (N_39538,N_31875,N_32129);
and U39539 (N_39539,N_34574,N_31538);
nor U39540 (N_39540,N_32549,N_32598);
and U39541 (N_39541,N_34715,N_31429);
nor U39542 (N_39542,N_34701,N_33128);
and U39543 (N_39543,N_30367,N_32206);
xnor U39544 (N_39544,N_32457,N_30216);
nor U39545 (N_39545,N_33381,N_34161);
and U39546 (N_39546,N_34514,N_30028);
nor U39547 (N_39547,N_32241,N_31930);
nor U39548 (N_39548,N_33200,N_30511);
or U39549 (N_39549,N_34273,N_34838);
xnor U39550 (N_39550,N_31305,N_31752);
and U39551 (N_39551,N_32770,N_30092);
nand U39552 (N_39552,N_34245,N_33388);
or U39553 (N_39553,N_34419,N_33087);
or U39554 (N_39554,N_31350,N_31643);
xor U39555 (N_39555,N_32349,N_30736);
nor U39556 (N_39556,N_33872,N_34605);
and U39557 (N_39557,N_32243,N_33112);
nand U39558 (N_39558,N_34690,N_34165);
xor U39559 (N_39559,N_31749,N_30044);
nor U39560 (N_39560,N_32178,N_34679);
nor U39561 (N_39561,N_30888,N_34926);
or U39562 (N_39562,N_33614,N_31816);
nor U39563 (N_39563,N_33290,N_33748);
nor U39564 (N_39564,N_30363,N_31557);
xor U39565 (N_39565,N_30344,N_32450);
nor U39566 (N_39566,N_33204,N_30439);
or U39567 (N_39567,N_34162,N_31716);
or U39568 (N_39568,N_31904,N_30844);
xor U39569 (N_39569,N_34312,N_33073);
nor U39570 (N_39570,N_33747,N_33758);
xor U39571 (N_39571,N_30412,N_32057);
xnor U39572 (N_39572,N_31455,N_33204);
or U39573 (N_39573,N_30724,N_31248);
nor U39574 (N_39574,N_31097,N_32360);
and U39575 (N_39575,N_34112,N_32159);
nand U39576 (N_39576,N_33432,N_30146);
xnor U39577 (N_39577,N_34015,N_32003);
nor U39578 (N_39578,N_33190,N_33463);
or U39579 (N_39579,N_33669,N_34553);
xor U39580 (N_39580,N_33452,N_31761);
xnor U39581 (N_39581,N_31328,N_32187);
xor U39582 (N_39582,N_32800,N_33471);
xnor U39583 (N_39583,N_30673,N_33025);
nor U39584 (N_39584,N_30235,N_33673);
or U39585 (N_39585,N_34672,N_31232);
and U39586 (N_39586,N_31886,N_34436);
or U39587 (N_39587,N_33227,N_33888);
and U39588 (N_39588,N_33062,N_33458);
nand U39589 (N_39589,N_30458,N_33977);
nor U39590 (N_39590,N_31035,N_33126);
xnor U39591 (N_39591,N_33174,N_32825);
xor U39592 (N_39592,N_30344,N_32331);
or U39593 (N_39593,N_34490,N_33791);
or U39594 (N_39594,N_33463,N_30414);
nor U39595 (N_39595,N_32175,N_34481);
xor U39596 (N_39596,N_31140,N_34370);
and U39597 (N_39597,N_31051,N_32414);
and U39598 (N_39598,N_30487,N_34544);
nor U39599 (N_39599,N_30519,N_34894);
nand U39600 (N_39600,N_31233,N_31157);
or U39601 (N_39601,N_33094,N_31612);
nor U39602 (N_39602,N_33132,N_30855);
or U39603 (N_39603,N_34797,N_32950);
nor U39604 (N_39604,N_34143,N_33863);
nor U39605 (N_39605,N_33833,N_30714);
xnor U39606 (N_39606,N_32007,N_32890);
nor U39607 (N_39607,N_32616,N_31442);
xor U39608 (N_39608,N_33454,N_34206);
xnor U39609 (N_39609,N_34709,N_30929);
or U39610 (N_39610,N_34314,N_31396);
nand U39611 (N_39611,N_33474,N_32969);
nand U39612 (N_39612,N_33178,N_30295);
nor U39613 (N_39613,N_34510,N_32918);
nand U39614 (N_39614,N_34987,N_32550);
nand U39615 (N_39615,N_34839,N_33688);
and U39616 (N_39616,N_34823,N_31240);
or U39617 (N_39617,N_34693,N_32175);
nor U39618 (N_39618,N_33857,N_32468);
nand U39619 (N_39619,N_30065,N_31619);
xnor U39620 (N_39620,N_33817,N_31541);
nand U39621 (N_39621,N_31010,N_31906);
xor U39622 (N_39622,N_30572,N_30840);
xor U39623 (N_39623,N_31122,N_32061);
nor U39624 (N_39624,N_33093,N_32345);
nand U39625 (N_39625,N_30989,N_34972);
xor U39626 (N_39626,N_30486,N_32169);
nor U39627 (N_39627,N_34126,N_33947);
nor U39628 (N_39628,N_30403,N_31088);
xor U39629 (N_39629,N_34352,N_32458);
xnor U39630 (N_39630,N_30172,N_32336);
xor U39631 (N_39631,N_30367,N_31983);
nand U39632 (N_39632,N_34990,N_30901);
and U39633 (N_39633,N_34107,N_32452);
or U39634 (N_39634,N_31084,N_32605);
xnor U39635 (N_39635,N_31905,N_30708);
nor U39636 (N_39636,N_34217,N_32160);
or U39637 (N_39637,N_34101,N_32638);
and U39638 (N_39638,N_30259,N_34426);
xor U39639 (N_39639,N_31405,N_33266);
or U39640 (N_39640,N_33053,N_31182);
nor U39641 (N_39641,N_32632,N_31424);
or U39642 (N_39642,N_34296,N_34003);
nand U39643 (N_39643,N_30440,N_31063);
and U39644 (N_39644,N_32537,N_33009);
nand U39645 (N_39645,N_31948,N_34714);
nor U39646 (N_39646,N_31133,N_34225);
and U39647 (N_39647,N_32539,N_33977);
and U39648 (N_39648,N_33692,N_34999);
or U39649 (N_39649,N_31397,N_31511);
nand U39650 (N_39650,N_31912,N_34793);
and U39651 (N_39651,N_32345,N_30936);
xor U39652 (N_39652,N_34282,N_33249);
and U39653 (N_39653,N_33423,N_33789);
nand U39654 (N_39654,N_33867,N_32594);
nand U39655 (N_39655,N_34583,N_34153);
or U39656 (N_39656,N_31560,N_31175);
xor U39657 (N_39657,N_33243,N_33721);
xor U39658 (N_39658,N_31343,N_30000);
nor U39659 (N_39659,N_33202,N_33483);
nor U39660 (N_39660,N_33477,N_33764);
nor U39661 (N_39661,N_31649,N_31852);
xor U39662 (N_39662,N_33295,N_30516);
and U39663 (N_39663,N_32675,N_31191);
xor U39664 (N_39664,N_33533,N_33531);
nand U39665 (N_39665,N_31800,N_31211);
and U39666 (N_39666,N_32599,N_30800);
and U39667 (N_39667,N_32505,N_34836);
nand U39668 (N_39668,N_32322,N_30640);
or U39669 (N_39669,N_33998,N_34781);
or U39670 (N_39670,N_33162,N_34495);
or U39671 (N_39671,N_33984,N_34315);
nand U39672 (N_39672,N_32072,N_31686);
and U39673 (N_39673,N_33633,N_30482);
or U39674 (N_39674,N_34822,N_31699);
xor U39675 (N_39675,N_33619,N_30859);
xor U39676 (N_39676,N_30640,N_34161);
and U39677 (N_39677,N_32855,N_31384);
or U39678 (N_39678,N_34062,N_34850);
and U39679 (N_39679,N_32949,N_32190);
or U39680 (N_39680,N_33976,N_33666);
nand U39681 (N_39681,N_34668,N_31413);
xnor U39682 (N_39682,N_30733,N_30506);
xor U39683 (N_39683,N_31336,N_34498);
nand U39684 (N_39684,N_33732,N_33158);
and U39685 (N_39685,N_32915,N_30942);
nor U39686 (N_39686,N_30520,N_34351);
nor U39687 (N_39687,N_30396,N_30139);
and U39688 (N_39688,N_32996,N_32927);
nor U39689 (N_39689,N_30965,N_31387);
nor U39690 (N_39690,N_33256,N_33257);
and U39691 (N_39691,N_34536,N_31229);
nand U39692 (N_39692,N_32476,N_34197);
xor U39693 (N_39693,N_34089,N_33992);
or U39694 (N_39694,N_32227,N_32648);
nor U39695 (N_39695,N_34143,N_33937);
xor U39696 (N_39696,N_32626,N_32945);
and U39697 (N_39697,N_32009,N_31872);
or U39698 (N_39698,N_30550,N_34262);
xor U39699 (N_39699,N_34345,N_33960);
or U39700 (N_39700,N_32387,N_31687);
or U39701 (N_39701,N_31395,N_31492);
nor U39702 (N_39702,N_33504,N_30304);
nand U39703 (N_39703,N_31151,N_30234);
and U39704 (N_39704,N_33216,N_33328);
or U39705 (N_39705,N_30741,N_31008);
nand U39706 (N_39706,N_34806,N_31659);
nand U39707 (N_39707,N_31348,N_34967);
and U39708 (N_39708,N_30118,N_31402);
xor U39709 (N_39709,N_31706,N_31602);
or U39710 (N_39710,N_34380,N_33934);
and U39711 (N_39711,N_30747,N_33570);
nand U39712 (N_39712,N_30943,N_32465);
nand U39713 (N_39713,N_30574,N_30232);
xnor U39714 (N_39714,N_31712,N_31679);
or U39715 (N_39715,N_33821,N_30936);
xnor U39716 (N_39716,N_30194,N_32579);
nand U39717 (N_39717,N_34824,N_31295);
nor U39718 (N_39718,N_32972,N_30164);
nor U39719 (N_39719,N_30079,N_32541);
or U39720 (N_39720,N_30873,N_32004);
nor U39721 (N_39721,N_30025,N_32982);
or U39722 (N_39722,N_33467,N_30984);
or U39723 (N_39723,N_34144,N_33130);
xnor U39724 (N_39724,N_32652,N_30806);
xor U39725 (N_39725,N_30726,N_34434);
nor U39726 (N_39726,N_32438,N_32602);
xnor U39727 (N_39727,N_31959,N_30122);
or U39728 (N_39728,N_31743,N_32605);
and U39729 (N_39729,N_30157,N_33321);
and U39730 (N_39730,N_31885,N_31500);
nor U39731 (N_39731,N_30090,N_32121);
or U39732 (N_39732,N_32848,N_33687);
nor U39733 (N_39733,N_34489,N_33086);
and U39734 (N_39734,N_31404,N_34720);
xnor U39735 (N_39735,N_30946,N_33291);
or U39736 (N_39736,N_32021,N_33481);
or U39737 (N_39737,N_32826,N_30211);
nor U39738 (N_39738,N_32058,N_33413);
xor U39739 (N_39739,N_31419,N_33736);
nor U39740 (N_39740,N_30805,N_31550);
nor U39741 (N_39741,N_34005,N_31553);
or U39742 (N_39742,N_33071,N_32074);
xor U39743 (N_39743,N_32671,N_31736);
or U39744 (N_39744,N_34010,N_34647);
nor U39745 (N_39745,N_30500,N_31924);
and U39746 (N_39746,N_31129,N_32296);
and U39747 (N_39747,N_31098,N_32472);
or U39748 (N_39748,N_30159,N_31289);
nand U39749 (N_39749,N_31003,N_33648);
or U39750 (N_39750,N_34999,N_31411);
xor U39751 (N_39751,N_31576,N_32446);
xnor U39752 (N_39752,N_33847,N_30867);
nor U39753 (N_39753,N_33602,N_31699);
nor U39754 (N_39754,N_34753,N_34931);
nand U39755 (N_39755,N_31406,N_30322);
nand U39756 (N_39756,N_31945,N_30642);
nand U39757 (N_39757,N_32259,N_33286);
and U39758 (N_39758,N_31228,N_33715);
and U39759 (N_39759,N_34010,N_31033);
nor U39760 (N_39760,N_30870,N_30135);
nor U39761 (N_39761,N_31931,N_32026);
and U39762 (N_39762,N_33830,N_30355);
nand U39763 (N_39763,N_31301,N_34190);
xor U39764 (N_39764,N_30040,N_32866);
or U39765 (N_39765,N_31236,N_33739);
nor U39766 (N_39766,N_32695,N_30326);
and U39767 (N_39767,N_32800,N_34752);
nor U39768 (N_39768,N_34603,N_32589);
xnor U39769 (N_39769,N_34652,N_31504);
nand U39770 (N_39770,N_33292,N_32802);
and U39771 (N_39771,N_32124,N_33414);
and U39772 (N_39772,N_31923,N_30959);
and U39773 (N_39773,N_33633,N_34120);
nor U39774 (N_39774,N_32909,N_34416);
or U39775 (N_39775,N_30841,N_31172);
or U39776 (N_39776,N_32355,N_31394);
and U39777 (N_39777,N_30862,N_30259);
and U39778 (N_39778,N_32342,N_34242);
and U39779 (N_39779,N_33833,N_34153);
or U39780 (N_39780,N_30971,N_31106);
nor U39781 (N_39781,N_30161,N_34595);
xor U39782 (N_39782,N_33543,N_31267);
nor U39783 (N_39783,N_30574,N_31631);
nand U39784 (N_39784,N_31978,N_34778);
or U39785 (N_39785,N_34363,N_32464);
and U39786 (N_39786,N_30338,N_34117);
xor U39787 (N_39787,N_32731,N_34950);
xor U39788 (N_39788,N_31620,N_33011);
nor U39789 (N_39789,N_30634,N_32610);
and U39790 (N_39790,N_31555,N_31615);
nand U39791 (N_39791,N_31837,N_30326);
and U39792 (N_39792,N_34886,N_31720);
xor U39793 (N_39793,N_31047,N_31668);
xor U39794 (N_39794,N_33031,N_34636);
nand U39795 (N_39795,N_33895,N_34905);
or U39796 (N_39796,N_31721,N_31714);
or U39797 (N_39797,N_30488,N_30674);
nor U39798 (N_39798,N_30067,N_33917);
nor U39799 (N_39799,N_32114,N_33433);
nand U39800 (N_39800,N_34760,N_32457);
nor U39801 (N_39801,N_31714,N_32803);
nand U39802 (N_39802,N_34284,N_32584);
or U39803 (N_39803,N_32621,N_32223);
nand U39804 (N_39804,N_30320,N_34780);
and U39805 (N_39805,N_31855,N_33007);
and U39806 (N_39806,N_31156,N_32358);
and U39807 (N_39807,N_34101,N_32060);
xor U39808 (N_39808,N_32743,N_34013);
nand U39809 (N_39809,N_32504,N_34496);
xor U39810 (N_39810,N_33463,N_30747);
and U39811 (N_39811,N_30392,N_31601);
xnor U39812 (N_39812,N_34161,N_33272);
or U39813 (N_39813,N_34656,N_33813);
nor U39814 (N_39814,N_34021,N_34376);
or U39815 (N_39815,N_30300,N_31161);
or U39816 (N_39816,N_32485,N_32553);
and U39817 (N_39817,N_34446,N_34408);
nand U39818 (N_39818,N_32996,N_32608);
nor U39819 (N_39819,N_30405,N_30978);
nor U39820 (N_39820,N_32061,N_34516);
or U39821 (N_39821,N_33285,N_33334);
nand U39822 (N_39822,N_30592,N_30012);
and U39823 (N_39823,N_34156,N_33426);
or U39824 (N_39824,N_33801,N_32921);
xnor U39825 (N_39825,N_31837,N_34041);
and U39826 (N_39826,N_34089,N_30353);
and U39827 (N_39827,N_30186,N_33082);
nor U39828 (N_39828,N_33288,N_33809);
nand U39829 (N_39829,N_33485,N_33240);
nand U39830 (N_39830,N_30331,N_33567);
and U39831 (N_39831,N_30158,N_31643);
nand U39832 (N_39832,N_32513,N_30408);
and U39833 (N_39833,N_31601,N_33591);
and U39834 (N_39834,N_31913,N_31377);
and U39835 (N_39835,N_33929,N_30173);
xnor U39836 (N_39836,N_33474,N_32785);
or U39837 (N_39837,N_32142,N_34806);
xnor U39838 (N_39838,N_31364,N_32912);
nand U39839 (N_39839,N_31781,N_34091);
and U39840 (N_39840,N_32859,N_33641);
nor U39841 (N_39841,N_32233,N_34807);
and U39842 (N_39842,N_32318,N_32998);
and U39843 (N_39843,N_31991,N_30451);
and U39844 (N_39844,N_30439,N_31762);
nor U39845 (N_39845,N_31685,N_33509);
xor U39846 (N_39846,N_34081,N_30847);
nand U39847 (N_39847,N_31080,N_32252);
or U39848 (N_39848,N_31603,N_33466);
nor U39849 (N_39849,N_33789,N_34848);
nor U39850 (N_39850,N_32566,N_31575);
nor U39851 (N_39851,N_34532,N_32159);
nor U39852 (N_39852,N_32275,N_34903);
nor U39853 (N_39853,N_30665,N_33009);
nand U39854 (N_39854,N_31077,N_33894);
xor U39855 (N_39855,N_31826,N_33959);
and U39856 (N_39856,N_30519,N_32062);
nor U39857 (N_39857,N_31868,N_34937);
or U39858 (N_39858,N_34925,N_33026);
nand U39859 (N_39859,N_30328,N_32754);
nand U39860 (N_39860,N_31367,N_32032);
nand U39861 (N_39861,N_32439,N_31568);
nor U39862 (N_39862,N_33055,N_33573);
nor U39863 (N_39863,N_32922,N_31467);
nor U39864 (N_39864,N_31690,N_30391);
or U39865 (N_39865,N_30978,N_34006);
nor U39866 (N_39866,N_32276,N_34200);
xor U39867 (N_39867,N_32939,N_31970);
and U39868 (N_39868,N_34324,N_31882);
nand U39869 (N_39869,N_31054,N_30268);
xor U39870 (N_39870,N_31188,N_32930);
and U39871 (N_39871,N_31895,N_31115);
and U39872 (N_39872,N_31736,N_34964);
nor U39873 (N_39873,N_31288,N_34353);
and U39874 (N_39874,N_32938,N_32095);
nor U39875 (N_39875,N_34232,N_34994);
or U39876 (N_39876,N_32584,N_33601);
xor U39877 (N_39877,N_34117,N_34347);
or U39878 (N_39878,N_31420,N_32075);
or U39879 (N_39879,N_34131,N_33416);
or U39880 (N_39880,N_33572,N_31884);
nor U39881 (N_39881,N_32766,N_32822);
nand U39882 (N_39882,N_31055,N_33457);
or U39883 (N_39883,N_31422,N_31619);
nand U39884 (N_39884,N_30854,N_34825);
and U39885 (N_39885,N_30822,N_32026);
xnor U39886 (N_39886,N_33044,N_31840);
and U39887 (N_39887,N_34247,N_31602);
or U39888 (N_39888,N_30682,N_33053);
and U39889 (N_39889,N_32257,N_30107);
nor U39890 (N_39890,N_31792,N_30575);
nand U39891 (N_39891,N_34555,N_33201);
nor U39892 (N_39892,N_33969,N_30304);
nor U39893 (N_39893,N_30843,N_33818);
nand U39894 (N_39894,N_30713,N_33049);
xor U39895 (N_39895,N_30200,N_32378);
or U39896 (N_39896,N_33431,N_32913);
or U39897 (N_39897,N_33158,N_32260);
nor U39898 (N_39898,N_33126,N_31207);
xnor U39899 (N_39899,N_33620,N_31366);
xnor U39900 (N_39900,N_31781,N_30104);
nand U39901 (N_39901,N_33213,N_31108);
and U39902 (N_39902,N_34451,N_34502);
nand U39903 (N_39903,N_30725,N_34183);
nand U39904 (N_39904,N_30251,N_33515);
nand U39905 (N_39905,N_32557,N_30391);
nand U39906 (N_39906,N_32232,N_30529);
xor U39907 (N_39907,N_34061,N_30869);
or U39908 (N_39908,N_34902,N_34300);
nand U39909 (N_39909,N_32091,N_31015);
nand U39910 (N_39910,N_32873,N_30788);
and U39911 (N_39911,N_33778,N_34908);
and U39912 (N_39912,N_31141,N_30627);
or U39913 (N_39913,N_30880,N_31377);
and U39914 (N_39914,N_31584,N_33758);
xor U39915 (N_39915,N_30317,N_33008);
nand U39916 (N_39916,N_34420,N_30596);
nor U39917 (N_39917,N_31368,N_33077);
or U39918 (N_39918,N_32920,N_32110);
and U39919 (N_39919,N_31247,N_34002);
or U39920 (N_39920,N_31719,N_34636);
nand U39921 (N_39921,N_33274,N_30907);
xnor U39922 (N_39922,N_31290,N_33361);
nand U39923 (N_39923,N_30928,N_34446);
nor U39924 (N_39924,N_33274,N_32961);
nand U39925 (N_39925,N_32929,N_34509);
or U39926 (N_39926,N_33494,N_33038);
or U39927 (N_39927,N_31266,N_34077);
or U39928 (N_39928,N_34581,N_32844);
and U39929 (N_39929,N_30455,N_34435);
nor U39930 (N_39930,N_32192,N_32324);
nand U39931 (N_39931,N_34181,N_30948);
or U39932 (N_39932,N_30805,N_31263);
nand U39933 (N_39933,N_30002,N_32885);
and U39934 (N_39934,N_32027,N_30434);
nand U39935 (N_39935,N_33610,N_34247);
or U39936 (N_39936,N_31788,N_32936);
and U39937 (N_39937,N_30313,N_33272);
nand U39938 (N_39938,N_34787,N_31699);
or U39939 (N_39939,N_34121,N_32382);
nand U39940 (N_39940,N_32307,N_33520);
xor U39941 (N_39941,N_32240,N_34253);
and U39942 (N_39942,N_30084,N_31972);
or U39943 (N_39943,N_31618,N_30594);
and U39944 (N_39944,N_32466,N_31604);
xnor U39945 (N_39945,N_34164,N_31526);
xor U39946 (N_39946,N_34367,N_34137);
nand U39947 (N_39947,N_31581,N_32958);
and U39948 (N_39948,N_34432,N_33680);
or U39949 (N_39949,N_34452,N_31609);
xor U39950 (N_39950,N_31309,N_32840);
xor U39951 (N_39951,N_33476,N_31781);
and U39952 (N_39952,N_33543,N_34117);
and U39953 (N_39953,N_33520,N_34207);
nor U39954 (N_39954,N_34512,N_31783);
nor U39955 (N_39955,N_31236,N_30740);
xnor U39956 (N_39956,N_31993,N_31941);
nand U39957 (N_39957,N_30386,N_34269);
and U39958 (N_39958,N_31250,N_32607);
or U39959 (N_39959,N_30877,N_34887);
or U39960 (N_39960,N_33558,N_31143);
nor U39961 (N_39961,N_33042,N_34672);
nor U39962 (N_39962,N_31297,N_33921);
nand U39963 (N_39963,N_34963,N_34981);
or U39964 (N_39964,N_34327,N_34003);
nor U39965 (N_39965,N_30952,N_33121);
xnor U39966 (N_39966,N_33957,N_33712);
or U39967 (N_39967,N_33860,N_34099);
nor U39968 (N_39968,N_34243,N_32021);
nor U39969 (N_39969,N_34132,N_30194);
nand U39970 (N_39970,N_33877,N_30299);
nand U39971 (N_39971,N_31539,N_30180);
xor U39972 (N_39972,N_30708,N_34612);
nand U39973 (N_39973,N_33197,N_34144);
or U39974 (N_39974,N_32115,N_32451);
nand U39975 (N_39975,N_32640,N_33345);
and U39976 (N_39976,N_34015,N_31364);
nor U39977 (N_39977,N_34016,N_31435);
nand U39978 (N_39978,N_33397,N_34858);
xor U39979 (N_39979,N_32372,N_30551);
nor U39980 (N_39980,N_30142,N_31460);
nand U39981 (N_39981,N_33477,N_34697);
nor U39982 (N_39982,N_30173,N_32436);
nand U39983 (N_39983,N_33245,N_32469);
nor U39984 (N_39984,N_31774,N_32989);
nand U39985 (N_39985,N_31291,N_34207);
xnor U39986 (N_39986,N_33709,N_34209);
nor U39987 (N_39987,N_30994,N_34739);
nor U39988 (N_39988,N_30549,N_30279);
xor U39989 (N_39989,N_34596,N_32008);
nand U39990 (N_39990,N_34765,N_30316);
nand U39991 (N_39991,N_31246,N_33658);
xor U39992 (N_39992,N_30659,N_33731);
xnor U39993 (N_39993,N_34656,N_30523);
nand U39994 (N_39994,N_32858,N_33682);
or U39995 (N_39995,N_32300,N_30179);
nand U39996 (N_39996,N_33780,N_33709);
nor U39997 (N_39997,N_30366,N_31319);
and U39998 (N_39998,N_30878,N_33545);
xor U39999 (N_39999,N_33287,N_34074);
nand U40000 (N_40000,N_38095,N_38648);
or U40001 (N_40001,N_35111,N_39100);
and U40002 (N_40002,N_38378,N_35462);
nand U40003 (N_40003,N_38860,N_39444);
xnor U40004 (N_40004,N_37988,N_35104);
nand U40005 (N_40005,N_38468,N_36807);
or U40006 (N_40006,N_37983,N_39682);
and U40007 (N_40007,N_38722,N_35426);
nor U40008 (N_40008,N_38526,N_39744);
or U40009 (N_40009,N_35871,N_38653);
nor U40010 (N_40010,N_39732,N_37481);
nand U40011 (N_40011,N_35656,N_37699);
nor U40012 (N_40012,N_37864,N_38743);
and U40013 (N_40013,N_35161,N_36922);
xor U40014 (N_40014,N_35954,N_35296);
xor U40015 (N_40015,N_35942,N_36615);
or U40016 (N_40016,N_35466,N_35067);
nand U40017 (N_40017,N_36951,N_35668);
xor U40018 (N_40018,N_39893,N_38100);
or U40019 (N_40019,N_37692,N_35892);
nand U40020 (N_40020,N_38242,N_37621);
nor U40021 (N_40021,N_35762,N_36860);
and U40022 (N_40022,N_37047,N_38727);
and U40023 (N_40023,N_38372,N_39642);
nand U40024 (N_40024,N_36466,N_37042);
nand U40025 (N_40025,N_38880,N_37541);
nand U40026 (N_40026,N_35253,N_37505);
nand U40027 (N_40027,N_36819,N_39422);
nor U40028 (N_40028,N_39330,N_37099);
nand U40029 (N_40029,N_36436,N_39602);
xor U40030 (N_40030,N_35481,N_35110);
xnor U40031 (N_40031,N_37901,N_39574);
nor U40032 (N_40032,N_36600,N_38348);
and U40033 (N_40033,N_39426,N_35363);
and U40034 (N_40034,N_36825,N_36540);
xor U40035 (N_40035,N_36306,N_37272);
nand U40036 (N_40036,N_38582,N_37343);
nand U40037 (N_40037,N_35168,N_38996);
or U40038 (N_40038,N_35131,N_37204);
nor U40039 (N_40039,N_37706,N_37034);
nor U40040 (N_40040,N_35840,N_37325);
nand U40041 (N_40041,N_35715,N_38855);
xnor U40042 (N_40042,N_39714,N_37708);
nor U40043 (N_40043,N_38199,N_37517);
and U40044 (N_40044,N_36167,N_36550);
and U40045 (N_40045,N_37188,N_35877);
and U40046 (N_40046,N_36791,N_36658);
xor U40047 (N_40047,N_35378,N_37591);
nor U40048 (N_40048,N_38944,N_37021);
nand U40049 (N_40049,N_37165,N_39521);
nand U40050 (N_40050,N_38583,N_37233);
or U40051 (N_40051,N_35555,N_39360);
and U40052 (N_40052,N_37599,N_36004);
nor U40053 (N_40053,N_36773,N_35554);
nand U40054 (N_40054,N_37922,N_37812);
xor U40055 (N_40055,N_35820,N_39763);
nor U40056 (N_40056,N_39498,N_38364);
nand U40057 (N_40057,N_39664,N_38902);
or U40058 (N_40058,N_37886,N_36835);
xor U40059 (N_40059,N_35227,N_36412);
nand U40060 (N_40060,N_35003,N_37435);
and U40061 (N_40061,N_36671,N_38363);
nand U40062 (N_40062,N_36169,N_36303);
and U40063 (N_40063,N_38802,N_38377);
xnor U40064 (N_40064,N_36445,N_36226);
xnor U40065 (N_40065,N_37347,N_37083);
nand U40066 (N_40066,N_36931,N_39910);
xnor U40067 (N_40067,N_37738,N_37202);
nand U40068 (N_40068,N_39186,N_35394);
or U40069 (N_40069,N_38057,N_35205);
nor U40070 (N_40070,N_37556,N_37789);
nor U40071 (N_40071,N_38266,N_37977);
and U40072 (N_40072,N_36644,N_37129);
or U40073 (N_40073,N_38098,N_36850);
nand U40074 (N_40074,N_37829,N_39601);
nor U40075 (N_40075,N_35091,N_39470);
and U40076 (N_40076,N_38233,N_38326);
nand U40077 (N_40077,N_36162,N_39812);
nor U40078 (N_40078,N_37206,N_39449);
or U40079 (N_40079,N_38719,N_39719);
nand U40080 (N_40080,N_35005,N_39181);
xor U40081 (N_40081,N_38573,N_38252);
and U40082 (N_40082,N_36564,N_35603);
nand U40083 (N_40083,N_35976,N_35155);
and U40084 (N_40084,N_37551,N_36417);
or U40085 (N_40085,N_38675,N_38999);
and U40086 (N_40086,N_37164,N_38205);
nand U40087 (N_40087,N_37120,N_39971);
or U40088 (N_40088,N_37746,N_37667);
nand U40089 (N_40089,N_36295,N_35611);
nor U40090 (N_40090,N_36896,N_35445);
and U40091 (N_40091,N_37562,N_38449);
nand U40092 (N_40092,N_37903,N_37716);
xor U40093 (N_40093,N_37795,N_37357);
or U40094 (N_40094,N_38932,N_39215);
or U40095 (N_40095,N_36499,N_39094);
nand U40096 (N_40096,N_38877,N_39972);
nor U40097 (N_40097,N_36752,N_36316);
nand U40098 (N_40098,N_38190,N_38504);
nand U40099 (N_40099,N_36214,N_35927);
nand U40100 (N_40100,N_37130,N_38894);
nand U40101 (N_40101,N_35360,N_35440);
xor U40102 (N_40102,N_37145,N_38460);
nor U40103 (N_40103,N_37902,N_37919);
xnor U40104 (N_40104,N_38056,N_35086);
or U40105 (N_40105,N_35267,N_37463);
xnor U40106 (N_40106,N_39241,N_39064);
nor U40107 (N_40107,N_37192,N_36885);
nor U40108 (N_40108,N_39488,N_37390);
nor U40109 (N_40109,N_38136,N_38714);
xnor U40110 (N_40110,N_37462,N_35053);
nor U40111 (N_40111,N_35446,N_37745);
and U40112 (N_40112,N_36977,N_36753);
or U40113 (N_40113,N_35951,N_36131);
nand U40114 (N_40114,N_37014,N_39684);
and U40115 (N_40115,N_37991,N_38300);
nand U40116 (N_40116,N_35000,N_35128);
nor U40117 (N_40117,N_37909,N_38376);
and U40118 (N_40118,N_39561,N_37679);
or U40119 (N_40119,N_36118,N_39520);
and U40120 (N_40120,N_35536,N_39443);
or U40121 (N_40121,N_38443,N_38997);
nor U40122 (N_40122,N_38030,N_37533);
nor U40123 (N_40123,N_36362,N_38977);
xor U40124 (N_40124,N_37298,N_37867);
nand U40125 (N_40125,N_38751,N_39441);
or U40126 (N_40126,N_38984,N_35088);
and U40127 (N_40127,N_36206,N_38303);
or U40128 (N_40128,N_39138,N_36985);
nor U40129 (N_40129,N_38404,N_39547);
or U40130 (N_40130,N_36231,N_36395);
and U40131 (N_40131,N_39029,N_37781);
nor U40132 (N_40132,N_38122,N_35051);
xnor U40133 (N_40133,N_37008,N_38625);
nor U40134 (N_40134,N_36211,N_37048);
or U40135 (N_40135,N_38606,N_37411);
or U40136 (N_40136,N_37931,N_36660);
nor U40137 (N_40137,N_35211,N_38116);
nand U40138 (N_40138,N_38695,N_38532);
and U40139 (N_40139,N_37531,N_39410);
nor U40140 (N_40140,N_35609,N_35882);
nor U40141 (N_40141,N_38344,N_37324);
nor U40142 (N_40142,N_35369,N_39674);
nor U40143 (N_40143,N_38649,N_38638);
nand U40144 (N_40144,N_35006,N_39324);
and U40145 (N_40145,N_37518,N_35780);
nand U40146 (N_40146,N_35852,N_37964);
or U40147 (N_40147,N_38288,N_36581);
nor U40148 (N_40148,N_36370,N_39124);
and U40149 (N_40149,N_37813,N_39501);
or U40150 (N_40150,N_37539,N_35242);
nor U40151 (N_40151,N_38257,N_38282);
nand U40152 (N_40152,N_39002,N_35746);
or U40153 (N_40153,N_35190,N_39354);
and U40154 (N_40154,N_35027,N_37979);
xnor U40155 (N_40155,N_36607,N_35008);
nand U40156 (N_40156,N_38674,N_38801);
and U40157 (N_40157,N_36763,N_35260);
nor U40158 (N_40158,N_36684,N_36081);
xnor U40159 (N_40159,N_38427,N_35239);
or U40160 (N_40160,N_35799,N_36341);
or U40161 (N_40161,N_36034,N_36256);
or U40162 (N_40162,N_39115,N_37450);
and U40163 (N_40163,N_35574,N_37513);
xnor U40164 (N_40164,N_39127,N_38729);
and U40165 (N_40165,N_37516,N_38644);
nor U40166 (N_40166,N_36947,N_37861);
nor U40167 (N_40167,N_35888,N_37924);
nor U40168 (N_40168,N_39901,N_39711);
and U40169 (N_40169,N_35818,N_38230);
xnor U40170 (N_40170,N_38875,N_37857);
and U40171 (N_40171,N_37117,N_35591);
nor U40172 (N_40172,N_39922,N_35766);
nand U40173 (N_40173,N_37836,N_35560);
xor U40174 (N_40174,N_35614,N_39681);
or U40175 (N_40175,N_36522,N_38898);
and U40176 (N_40176,N_39982,N_39276);
xnor U40177 (N_40177,N_38508,N_36715);
xor U40178 (N_40178,N_37362,N_36203);
nand U40179 (N_40179,N_35066,N_37990);
nor U40180 (N_40180,N_38793,N_36146);
xor U40181 (N_40181,N_36641,N_38487);
xnor U40182 (N_40182,N_36403,N_36862);
nand U40183 (N_40183,N_38628,N_38294);
nor U40184 (N_40184,N_37035,N_36802);
or U40185 (N_40185,N_39069,N_35548);
nand U40186 (N_40186,N_37624,N_36024);
nor U40187 (N_40187,N_37664,N_36806);
nor U40188 (N_40188,N_39286,N_39586);
or U40189 (N_40189,N_37754,N_36039);
nor U40190 (N_40190,N_35136,N_38130);
xnor U40191 (N_40191,N_36317,N_36552);
and U40192 (N_40192,N_35180,N_39183);
or U40193 (N_40193,N_37578,N_35809);
nor U40194 (N_40194,N_36220,N_36419);
nor U40195 (N_40195,N_35203,N_38853);
or U40196 (N_40196,N_36778,N_37189);
and U40197 (N_40197,N_39479,N_35345);
nand U40198 (N_40198,N_39243,N_35596);
xnor U40199 (N_40199,N_36283,N_36032);
nor U40200 (N_40200,N_38187,N_38014);
and U40201 (N_40201,N_36765,N_35215);
or U40202 (N_40202,N_38151,N_35889);
and U40203 (N_40203,N_36863,N_35659);
or U40204 (N_40204,N_37464,N_35350);
nand U40205 (N_40205,N_37452,N_36215);
nand U40206 (N_40206,N_36062,N_38626);
nand U40207 (N_40207,N_39960,N_37474);
and U40208 (N_40208,N_35972,N_35737);
nand U40209 (N_40209,N_36733,N_36265);
nor U40210 (N_40210,N_35404,N_38071);
and U40211 (N_40211,N_35571,N_39679);
xor U40212 (N_40212,N_37495,N_39762);
nand U40213 (N_40213,N_35056,N_36135);
or U40214 (N_40214,N_35226,N_35830);
xnor U40215 (N_40215,N_39340,N_36350);
nor U40216 (N_40216,N_38960,N_39167);
xor U40217 (N_40217,N_36194,N_37548);
xnor U40218 (N_40218,N_39843,N_35077);
xnor U40219 (N_40219,N_38097,N_35802);
nor U40220 (N_40220,N_36614,N_38519);
nor U40221 (N_40221,N_36814,N_35558);
nor U40222 (N_40222,N_35270,N_38935);
and U40223 (N_40223,N_36302,N_37156);
or U40224 (N_40224,N_35773,N_37788);
or U40225 (N_40225,N_37765,N_38995);
or U40226 (N_40226,N_37482,N_37076);
xnor U40227 (N_40227,N_36331,N_39404);
xnor U40228 (N_40228,N_37530,N_37652);
nor U40229 (N_40229,N_38873,N_35549);
xor U40230 (N_40230,N_36795,N_37786);
nor U40231 (N_40231,N_39366,N_35801);
nand U40232 (N_40232,N_36139,N_38211);
nand U40233 (N_40233,N_38076,N_39209);
and U40234 (N_40234,N_37088,N_38170);
or U40235 (N_40235,N_36213,N_36358);
nand U40236 (N_40236,N_39596,N_38134);
nor U40237 (N_40237,N_39423,N_35035);
or U40238 (N_40238,N_37802,N_38567);
nand U40239 (N_40239,N_38384,N_39944);
nor U40240 (N_40240,N_36707,N_35079);
or U40241 (N_40241,N_38911,N_38315);
and U40242 (N_40242,N_37568,N_37693);
nor U40243 (N_40243,N_39841,N_38991);
and U40244 (N_40244,N_36962,N_39567);
xnor U40245 (N_40245,N_36347,N_35414);
nor U40246 (N_40246,N_38424,N_37649);
or U40247 (N_40247,N_38618,N_37115);
xor U40248 (N_40248,N_35425,N_37507);
and U40249 (N_40249,N_36784,N_38948);
and U40250 (N_40250,N_39387,N_35074);
nand U40251 (N_40251,N_37328,N_37808);
xor U40252 (N_40252,N_37413,N_35633);
nand U40253 (N_40253,N_37395,N_36332);
and U40254 (N_40254,N_39385,N_38402);
or U40255 (N_40255,N_35480,N_35777);
and U40256 (N_40256,N_36234,N_39525);
and U40257 (N_40257,N_39578,N_35935);
xor U40258 (N_40258,N_35014,N_36558);
and U40259 (N_40259,N_38311,N_38044);
nand U40260 (N_40260,N_37590,N_36170);
nand U40261 (N_40261,N_37564,N_35418);
nor U40262 (N_40262,N_37195,N_39786);
and U40263 (N_40263,N_37797,N_38631);
nor U40264 (N_40264,N_39053,N_37442);
xor U40265 (N_40265,N_39199,N_37025);
nand U40266 (N_40266,N_35071,N_36230);
or U40267 (N_40267,N_35095,N_36013);
and U40268 (N_40268,N_39870,N_38810);
xnor U40269 (N_40269,N_39620,N_38678);
nand U40270 (N_40270,N_38886,N_37532);
nor U40271 (N_40271,N_38682,N_39236);
nor U40272 (N_40272,N_35070,N_37213);
or U40273 (N_40273,N_35754,N_36424);
nor U40274 (N_40274,N_37234,N_35714);
or U40275 (N_40275,N_37461,N_36526);
nand U40276 (N_40276,N_38803,N_35007);
xor U40277 (N_40277,N_38926,N_36810);
or U40278 (N_40278,N_37028,N_35087);
and U40279 (N_40279,N_38856,N_39861);
or U40280 (N_40280,N_35312,N_35616);
or U40281 (N_40281,N_38261,N_35020);
nor U40282 (N_40282,N_37140,N_37663);
and U40283 (N_40283,N_35415,N_35955);
nor U40284 (N_40284,N_37330,N_36373);
and U40285 (N_40285,N_38456,N_36887);
nand U40286 (N_40286,N_39144,N_35430);
or U40287 (N_40287,N_38223,N_35594);
nor U40288 (N_40288,N_39273,N_39742);
nor U40289 (N_40289,N_39318,N_35285);
nand U40290 (N_40290,N_36340,N_37589);
xor U40291 (N_40291,N_36544,N_36545);
nand U40292 (N_40292,N_38276,N_37739);
xor U40293 (N_40293,N_38409,N_36524);
and U40294 (N_40294,N_37170,N_39553);
xor U40295 (N_40295,N_39457,N_39357);
nand U40296 (N_40296,N_38800,N_37874);
or U40297 (N_40297,N_35678,N_35843);
xnor U40298 (N_40298,N_37199,N_36503);
and U40299 (N_40299,N_37329,N_39832);
or U40300 (N_40300,N_39891,N_39631);
or U40301 (N_40301,N_35405,N_36443);
and U40302 (N_40302,N_35846,N_38435);
nand U40303 (N_40303,N_37185,N_37618);
xor U40304 (N_40304,N_39489,N_36656);
nand U40305 (N_40305,N_35585,N_36553);
nor U40306 (N_40306,N_39780,N_39776);
nor U40307 (N_40307,N_39809,N_39595);
nor U40308 (N_40308,N_37065,N_38467);
nand U40309 (N_40309,N_38844,N_39746);
or U40310 (N_40310,N_37225,N_39311);
nand U40311 (N_40311,N_36228,N_38702);
or U40312 (N_40312,N_37554,N_36255);
xor U40313 (N_40313,N_38167,N_38084);
and U40314 (N_40314,N_37950,N_36668);
xor U40315 (N_40315,N_37023,N_39874);
nand U40316 (N_40316,N_37794,N_38281);
or U40317 (N_40317,N_37602,N_39075);
or U40318 (N_40318,N_38015,N_37080);
nand U40319 (N_40319,N_35520,N_38652);
and U40320 (N_40320,N_35865,N_36601);
or U40321 (N_40321,N_39855,N_36312);
xor U40322 (N_40322,N_38804,N_35826);
nor U40323 (N_40323,N_37038,N_36884);
or U40324 (N_40324,N_35338,N_38848);
nor U40325 (N_40325,N_38368,N_35719);
or U40326 (N_40326,N_36346,N_36045);
nor U40327 (N_40327,N_38365,N_39690);
nor U40328 (N_40328,N_35220,N_35769);
nor U40329 (N_40329,N_36904,N_37559);
or U40330 (N_40330,N_38092,N_38453);
and U40331 (N_40331,N_39698,N_36383);
nand U40332 (N_40332,N_35080,N_38710);
nand U40333 (N_40333,N_39300,N_35717);
nand U40334 (N_40334,N_39765,N_36803);
xnor U40335 (N_40335,N_36879,N_35249);
nand U40336 (N_40336,N_39755,N_36478);
nand U40337 (N_40337,N_37987,N_35283);
xnor U40338 (N_40338,N_39775,N_38045);
or U40339 (N_40339,N_35461,N_37306);
and U40340 (N_40340,N_37388,N_38235);
nor U40341 (N_40341,N_38910,N_36680);
xor U40342 (N_40342,N_35858,N_38597);
nor U40343 (N_40343,N_39701,N_36809);
or U40344 (N_40344,N_37106,N_35647);
nor U40345 (N_40345,N_35109,N_38826);
xor U40346 (N_40346,N_37546,N_38073);
xnor U40347 (N_40347,N_39047,N_39139);
nand U40348 (N_40348,N_35867,N_38983);
or U40349 (N_40349,N_39799,N_37587);
and U40350 (N_40350,N_35417,N_35307);
nand U40351 (N_40351,N_39473,N_35269);
and U40352 (N_40352,N_38185,N_39382);
or U40353 (N_40353,N_39274,N_38025);
xnor U40354 (N_40354,N_36304,N_35512);
or U40355 (N_40355,N_37181,N_37910);
nor U40356 (N_40356,N_35097,N_37301);
nor U40357 (N_40357,N_36177,N_36400);
nand U40358 (N_40358,N_38499,N_36975);
nor U40359 (N_40359,N_36520,N_37792);
nand U40360 (N_40360,N_39331,N_38643);
nor U40361 (N_40361,N_38335,N_36178);
xor U40362 (N_40362,N_38240,N_37271);
and U40363 (N_40363,N_35488,N_37895);
nor U40364 (N_40364,N_36221,N_39436);
nor U40365 (N_40365,N_38473,N_37107);
nor U40366 (N_40366,N_36826,N_36543);
and U40367 (N_40367,N_36834,N_38392);
nor U40368 (N_40368,N_38849,N_38574);
or U40369 (N_40369,N_37240,N_36473);
nand U40370 (N_40370,N_37776,N_37593);
nand U40371 (N_40371,N_37488,N_39081);
nor U40372 (N_40372,N_39579,N_35620);
nand U40373 (N_40373,N_39162,N_38947);
xor U40374 (N_40374,N_35586,N_38740);
and U40375 (N_40375,N_35492,N_35981);
xnor U40376 (N_40376,N_36998,N_39011);
or U40377 (N_40377,N_37498,N_39604);
or U40378 (N_40378,N_36175,N_39234);
or U40379 (N_40379,N_39691,N_37597);
or U40380 (N_40380,N_39953,N_36950);
nor U40381 (N_40381,N_37997,N_37643);
nand U40382 (N_40382,N_38918,N_35043);
nand U40383 (N_40383,N_37421,N_35037);
and U40384 (N_40384,N_37758,N_38807);
xor U40385 (N_40385,N_39367,N_39315);
and U40386 (N_40386,N_37501,N_37611);
xor U40387 (N_40387,N_39233,N_39519);
nor U40388 (N_40388,N_35519,N_37059);
and U40389 (N_40389,N_36248,N_35496);
nor U40390 (N_40390,N_39980,N_39424);
or U40391 (N_40391,N_36467,N_39509);
nor U40392 (N_40392,N_37661,N_39802);
and U40393 (N_40393,N_36409,N_39342);
and U40394 (N_40394,N_38485,N_36264);
and U40395 (N_40395,N_35721,N_38655);
nor U40396 (N_40396,N_39288,N_36730);
or U40397 (N_40397,N_39878,N_35686);
nand U40398 (N_40398,N_35805,N_39463);
xor U40399 (N_40399,N_38283,N_36136);
nor U40400 (N_40400,N_38132,N_39440);
nor U40401 (N_40401,N_36800,N_37926);
xor U40402 (N_40402,N_38731,N_39514);
xnor U40403 (N_40403,N_36128,N_35956);
nand U40404 (N_40404,N_35544,N_39510);
and U40405 (N_40405,N_36687,N_37804);
nor U40406 (N_40406,N_37852,N_36416);
nand U40407 (N_40407,N_37859,N_39425);
xor U40408 (N_40408,N_39790,N_38557);
nor U40409 (N_40409,N_37359,N_36993);
and U40410 (N_40410,N_39591,N_36547);
or U40411 (N_40411,N_37166,N_37102);
nand U40412 (N_40412,N_37223,N_36193);
nand U40413 (N_40413,N_35228,N_38559);
nand U40414 (N_40414,N_39329,N_35120);
xnor U40415 (N_40415,N_37623,N_35989);
and U40416 (N_40416,N_37489,N_37119);
or U40417 (N_40417,N_36508,N_39542);
nor U40418 (N_40418,N_36273,N_39439);
xnor U40419 (N_40419,N_36469,N_35158);
and U40420 (N_40420,N_37446,N_39560);
or U40421 (N_40421,N_38382,N_36134);
xor U40422 (N_40422,N_35062,N_39245);
or U40423 (N_40423,N_35709,N_38397);
xnor U40424 (N_40424,N_35793,N_36593);
nor U40425 (N_40425,N_37002,N_38061);
nor U40426 (N_40426,N_35710,N_36844);
or U40427 (N_40427,N_37383,N_38824);
xnor U40428 (N_40428,N_35085,N_37478);
or U40429 (N_40429,N_35272,N_35996);
xor U40430 (N_40430,N_36669,N_39563);
nand U40431 (N_40431,N_39196,N_36396);
and U40432 (N_40432,N_36461,N_37209);
nand U40433 (N_40433,N_37538,N_36455);
nor U40434 (N_40434,N_36992,N_38884);
nand U40435 (N_40435,N_38159,N_39344);
and U40436 (N_40436,N_39713,N_37892);
xor U40437 (N_40437,N_39941,N_37900);
nor U40438 (N_40438,N_38032,N_36204);
nor U40439 (N_40439,N_36165,N_37999);
and U40440 (N_40440,N_35610,N_35367);
nor U40441 (N_40441,N_39600,N_39702);
or U40442 (N_40442,N_38333,N_37869);
nand U40443 (N_40443,N_37082,N_38328);
xnor U40444 (N_40444,N_39229,N_37976);
and U40445 (N_40445,N_39590,N_37053);
or U40446 (N_40446,N_35978,N_36647);
xor U40447 (N_40447,N_39527,N_36352);
nor U40448 (N_40448,N_39198,N_39882);
nor U40449 (N_40449,N_39013,N_39524);
nor U40450 (N_40450,N_35167,N_38897);
nand U40451 (N_40451,N_39380,N_37437);
xnor U40452 (N_40452,N_38792,N_37515);
xnor U40453 (N_40453,N_35811,N_36238);
xnor U40454 (N_40454,N_37400,N_35564);
nor U40455 (N_40455,N_36421,N_36389);
nand U40456 (N_40456,N_35191,N_37424);
xnor U40457 (N_40457,N_37845,N_38505);
and U40458 (N_40458,N_35624,N_35997);
xnor U40459 (N_40459,N_37607,N_37735);
and U40460 (N_40460,N_36685,N_36190);
and U40461 (N_40461,N_38290,N_35464);
nor U40462 (N_40462,N_39597,N_37617);
nand U40463 (N_40463,N_39195,N_39207);
nor U40464 (N_40464,N_37430,N_38863);
nor U40465 (N_40465,N_36839,N_38296);
nor U40466 (N_40466,N_39237,N_38490);
or U40467 (N_40467,N_39728,N_38815);
or U40468 (N_40468,N_36718,N_38812);
nor U40469 (N_40469,N_38987,N_35510);
or U40470 (N_40470,N_39572,N_35287);
and U40471 (N_40471,N_38500,N_36491);
xnor U40472 (N_40472,N_36571,N_36102);
nand U40473 (N_40473,N_38789,N_37459);
or U40474 (N_40474,N_35775,N_37820);
or U40475 (N_40475,N_39370,N_39408);
nor U40476 (N_40476,N_37094,N_35685);
xnor U40477 (N_40477,N_39582,N_38492);
and U40478 (N_40478,N_38823,N_39883);
and U40479 (N_40479,N_38677,N_35838);
xnor U40480 (N_40480,N_35293,N_37208);
or U40481 (N_40481,N_39628,N_37353);
or U40482 (N_40482,N_39598,N_37963);
or U40483 (N_40483,N_36768,N_39748);
nor U40484 (N_40484,N_35171,N_36980);
or U40485 (N_40485,N_37975,N_38245);
or U40486 (N_40486,N_37441,N_35883);
nand U40487 (N_40487,N_36866,N_37540);
and U40488 (N_40488,N_36319,N_39903);
nand U40489 (N_40489,N_36725,N_38580);
and U40490 (N_40490,N_36551,N_38882);
nor U40491 (N_40491,N_36832,N_37029);
and U40492 (N_40492,N_37402,N_37259);
nor U40493 (N_40493,N_38201,N_39968);
or U40494 (N_40494,N_36723,N_39929);
nor U40495 (N_40495,N_35924,N_38528);
and U40496 (N_40496,N_35410,N_36476);
xnor U40497 (N_40497,N_37855,N_37755);
nand U40498 (N_40498,N_37000,N_37220);
and U40499 (N_40499,N_37332,N_39087);
or U40500 (N_40500,N_36309,N_35371);
nor U40501 (N_40501,N_35295,N_37001);
or U40502 (N_40502,N_36738,N_37238);
xor U40503 (N_40503,N_39751,N_38157);
xor U40504 (N_40504,N_38144,N_37469);
or U40505 (N_40505,N_37672,N_36065);
nor U40506 (N_40506,N_38733,N_35791);
nor U40507 (N_40507,N_38430,N_37937);
and U40508 (N_40508,N_37367,N_37338);
or U40509 (N_40509,N_36908,N_37177);
nor U40510 (N_40510,N_37064,N_38964);
or U40511 (N_40511,N_39617,N_36023);
nand U40512 (N_40512,N_36785,N_38651);
xnor U40513 (N_40513,N_36640,N_38813);
xor U40514 (N_40514,N_37711,N_38482);
or U40515 (N_40515,N_35139,N_37475);
nor U40516 (N_40516,N_37257,N_36981);
and U40517 (N_40517,N_36015,N_36654);
nand U40518 (N_40518,N_37473,N_38149);
xor U40519 (N_40519,N_37282,N_35819);
nand U40520 (N_40520,N_36191,N_37360);
or U40521 (N_40521,N_38093,N_35315);
and U40522 (N_40522,N_36747,N_39869);
nor U40523 (N_40523,N_38118,N_38291);
or U40524 (N_40524,N_37816,N_37876);
xnor U40525 (N_40525,N_39316,N_35500);
or U40526 (N_40526,N_37237,N_35828);
nand U40527 (N_40527,N_37563,N_36114);
xor U40528 (N_40528,N_39848,N_39759);
xor U40529 (N_40529,N_38068,N_39708);
xor U40530 (N_40530,N_38135,N_36902);
and U40531 (N_40531,N_39267,N_39540);
and U40532 (N_40532,N_37550,N_35539);
nor U40533 (N_40533,N_37303,N_38064);
nor U40534 (N_40534,N_37331,N_39170);
nand U40535 (N_40535,N_39113,N_38284);
xnor U40536 (N_40536,N_35320,N_36851);
nor U40537 (N_40537,N_39727,N_39310);
xor U40538 (N_40538,N_39393,N_37992);
or U40539 (N_40539,N_37807,N_36613);
nand U40540 (N_40540,N_38091,N_39208);
or U40541 (N_40541,N_39838,N_36033);
nor U40542 (N_40542,N_37557,N_35870);
xnor U40543 (N_40543,N_35577,N_36000);
xor U40544 (N_40544,N_35025,N_39725);
nor U40545 (N_40545,N_36355,N_36489);
xor U40546 (N_40546,N_38513,N_35973);
or U40547 (N_40547,N_37942,N_35038);
nor U40548 (N_40548,N_35957,N_39830);
or U40549 (N_40549,N_36774,N_36037);
nor U40550 (N_40550,N_37944,N_37255);
nand U40551 (N_40551,N_39337,N_38103);
nor U40552 (N_40552,N_35334,N_38317);
nor U40553 (N_40553,N_39362,N_38830);
nand U40554 (N_40554,N_35116,N_38096);
and U40555 (N_40555,N_39807,N_39866);
nor U40556 (N_40556,N_35650,N_35706);
or U40557 (N_40557,N_37334,N_36123);
xnor U40558 (N_40558,N_37139,N_39017);
xor U40559 (N_40559,N_35324,N_35040);
xnor U40560 (N_40560,N_39289,N_38236);
nor U40561 (N_40561,N_35436,N_36141);
nand U40562 (N_40562,N_39159,N_36789);
or U40563 (N_40563,N_38082,N_36827);
or U40564 (N_40564,N_38186,N_36293);
and U40565 (N_40565,N_38247,N_39834);
nand U40566 (N_40566,N_39492,N_35001);
xor U40567 (N_40567,N_36637,N_36174);
xnor U40568 (N_40568,N_39432,N_38246);
nand U40569 (N_40569,N_37216,N_36188);
nor U40570 (N_40570,N_36260,N_36051);
nor U40571 (N_40571,N_39639,N_38010);
xor U40572 (N_40572,N_35567,N_39296);
nand U40573 (N_40573,N_37239,N_39956);
nand U40574 (N_40574,N_35649,N_36936);
nand U40575 (N_40575,N_38287,N_39394);
and U40576 (N_40576,N_36681,N_35031);
or U40577 (N_40577,N_35969,N_35580);
nand U40578 (N_40578,N_37837,N_39522);
and U40579 (N_40579,N_39794,N_35059);
nand U40580 (N_40580,N_36143,N_35705);
xnor U40581 (N_40581,N_35143,N_39961);
nand U40582 (N_40582,N_39661,N_36115);
nand U40583 (N_40583,N_35789,N_39782);
or U40584 (N_40584,N_38008,N_37198);
or U40585 (N_40585,N_36253,N_39182);
or U40586 (N_40586,N_35076,N_36597);
xor U40587 (N_40587,N_38673,N_37485);
nor U40588 (N_40588,N_39148,N_36793);
nor U40589 (N_40589,N_39784,N_38602);
nand U40590 (N_40590,N_36808,N_35332);
nand U40591 (N_40591,N_37881,N_36963);
or U40592 (N_40592,N_38928,N_37671);
or U40593 (N_40593,N_39907,N_39483);
or U40594 (N_40594,N_38034,N_39833);
nand U40595 (N_40595,N_39309,N_35535);
and U40596 (N_40596,N_38415,N_36129);
and U40597 (N_40597,N_35300,N_39994);
nor U40598 (N_40598,N_35758,N_35049);
nand U40599 (N_40599,N_36072,N_35195);
or U40600 (N_40600,N_38307,N_37251);
xor U40601 (N_40601,N_35508,N_38868);
xor U40602 (N_40602,N_35864,N_38318);
or U40603 (N_40603,N_35640,N_37157);
xor U40604 (N_40604,N_36053,N_35855);
xor U40605 (N_40605,N_37815,N_39263);
nand U40606 (N_40606,N_36001,N_36453);
xor U40607 (N_40607,N_37722,N_39715);
nand U40608 (N_40608,N_39939,N_39254);
xor U40609 (N_40609,N_35911,N_38060);
nor U40610 (N_40610,N_37715,N_39261);
or U40611 (N_40611,N_38414,N_37210);
and U40612 (N_40612,N_39459,N_39168);
nor U40613 (N_40613,N_35385,N_39645);
or U40614 (N_40614,N_39131,N_35256);
and U40615 (N_40615,N_37763,N_35004);
or U40616 (N_40616,N_39825,N_38697);
or U40617 (N_40617,N_39771,N_39652);
nor U40618 (N_40618,N_35975,N_36092);
and U40619 (N_40619,N_35925,N_38587);
nand U40620 (N_40620,N_37730,N_38560);
or U40621 (N_40621,N_39614,N_35831);
nand U40622 (N_40622,N_38152,N_35210);
xor U40623 (N_40623,N_39073,N_38750);
or U40624 (N_40624,N_39141,N_39427);
nand U40625 (N_40625,N_36974,N_35442);
nand U40626 (N_40626,N_35763,N_36515);
nand U40627 (N_40627,N_39246,N_37787);
nand U40628 (N_40628,N_39526,N_37184);
nand U40629 (N_40629,N_35186,N_39202);
or U40630 (N_40630,N_38799,N_38562);
xnor U40631 (N_40631,N_39482,N_36127);
or U40632 (N_40632,N_37118,N_37100);
nand U40633 (N_40633,N_37698,N_37158);
nor U40634 (N_40634,N_38295,N_35380);
nor U40635 (N_40635,N_38065,N_38917);
and U40636 (N_40636,N_38905,N_38747);
xnor U40637 (N_40637,N_38020,N_39230);
xnor U40638 (N_40638,N_37472,N_36661);
or U40639 (N_40639,N_36390,N_39616);
xor U40640 (N_40640,N_35114,N_35305);
nand U40641 (N_40641,N_37772,N_39877);
nand U40642 (N_40642,N_37142,N_36991);
and U40643 (N_40643,N_35931,N_35182);
and U40644 (N_40644,N_35152,N_35246);
nor U40645 (N_40645,N_37358,N_39472);
and U40646 (N_40646,N_38726,N_38538);
and U40647 (N_40647,N_39608,N_36392);
nor U40648 (N_40648,N_38970,N_36030);
and U40649 (N_40649,N_36497,N_37622);
nor U40650 (N_40650,N_38006,N_39722);
nor U40651 (N_40651,N_39648,N_35727);
xnor U40652 (N_40652,N_39466,N_36029);
nand U40653 (N_40653,N_37916,N_35505);
nor U40654 (N_40654,N_36638,N_36439);
xnor U40655 (N_40655,N_39325,N_35393);
and U40656 (N_40656,N_39967,N_39686);
and U40657 (N_40657,N_36828,N_39851);
and U40658 (N_40658,N_36986,N_36454);
xnor U40659 (N_40659,N_38503,N_38314);
or U40660 (N_40660,N_37918,N_35880);
nand U40661 (N_40661,N_36935,N_37480);
and U40662 (N_40662,N_36901,N_39863);
xnor U40663 (N_40663,N_39914,N_36003);
xnor U40664 (N_40664,N_37929,N_36567);
xor U40665 (N_40665,N_35451,N_35331);
xnor U40666 (N_40666,N_35379,N_35692);
or U40667 (N_40667,N_36163,N_38362);
nor U40668 (N_40668,N_35456,N_35083);
nor U40669 (N_40669,N_37971,N_35009);
or U40670 (N_40670,N_38543,N_38260);
and U40671 (N_40671,N_37702,N_37194);
xor U40672 (N_40672,N_37884,N_39688);
nand U40673 (N_40673,N_36915,N_36080);
or U40674 (N_40674,N_36557,N_38229);
nor U40675 (N_40675,N_39532,N_36924);
or U40676 (N_40676,N_36465,N_39411);
nor U40677 (N_40677,N_38209,N_39641);
xnor U40678 (N_40678,N_35604,N_37954);
nor U40679 (N_40679,N_39804,N_37753);
or U40680 (N_40680,N_37570,N_37822);
or U40681 (N_40681,N_35042,N_39098);
nand U40682 (N_40682,N_36195,N_36232);
and U40683 (N_40683,N_38754,N_38581);
xor U40684 (N_40684,N_35660,N_39294);
nor U40685 (N_40685,N_35600,N_38555);
nand U40686 (N_40686,N_37134,N_38146);
and U40687 (N_40687,N_38972,N_39227);
nor U40688 (N_40688,N_36729,N_35184);
and U40689 (N_40689,N_37732,N_37093);
xor U40690 (N_40690,N_37349,N_35546);
and U40691 (N_40691,N_35552,N_35234);
nand U40692 (N_40692,N_39268,N_39632);
xnor U40693 (N_40693,N_37426,N_35221);
and U40694 (N_40694,N_38219,N_36132);
or U40695 (N_40695,N_39353,N_38117);
and U40696 (N_40696,N_35946,N_36611);
and U40697 (N_40697,N_39613,N_35879);
or U40698 (N_40698,N_39811,N_37022);
or U40699 (N_40699,N_36224,N_36327);
xnor U40700 (N_40700,N_36233,N_35169);
xor U40701 (N_40701,N_36181,N_35311);
xnor U40702 (N_40702,N_38204,N_35386);
nand U40703 (N_40703,N_35964,N_37308);
or U40704 (N_40704,N_35903,N_36158);
or U40705 (N_40705,N_36320,N_39206);
xor U40706 (N_40706,N_36939,N_38623);
nor U40707 (N_40707,N_35375,N_39180);
nor U40708 (N_40708,N_37394,N_37734);
and U40709 (N_40709,N_38657,N_35501);
nand U40710 (N_40710,N_37519,N_35034);
nor U40711 (N_40711,N_35096,N_37150);
nor U40712 (N_40712,N_38617,N_38489);
nor U40713 (N_40713,N_37246,N_39927);
nor U40714 (N_40714,N_36954,N_36565);
or U40715 (N_40715,N_38024,N_38746);
nor U40716 (N_40716,N_37736,N_38310);
or U40717 (N_40717,N_37340,N_39248);
nand U40718 (N_40718,N_37377,N_37406);
or U40719 (N_40719,N_35915,N_38831);
nand U40720 (N_40720,N_35225,N_39752);
xor U40721 (N_40721,N_36628,N_38825);
nor U40722 (N_40722,N_35563,N_39951);
nor U40723 (N_40723,N_37467,N_38264);
nand U40724 (N_40724,N_36479,N_37211);
nor U40725 (N_40725,N_38600,N_38193);
or U40726 (N_40726,N_39247,N_36790);
xor U40727 (N_40727,N_38725,N_39815);
nor U40728 (N_40728,N_38051,N_38463);
xor U40729 (N_40729,N_35808,N_39923);
or U40730 (N_40730,N_36812,N_35816);
nand U40731 (N_40731,N_38011,N_35245);
and U40732 (N_40732,N_39039,N_36679);
or U40733 (N_40733,N_36277,N_38820);
nor U40734 (N_40734,N_36599,N_35891);
and U40735 (N_40735,N_37336,N_37063);
or U40736 (N_40736,N_35118,N_36166);
and U40737 (N_40737,N_36662,N_39564);
nor U40738 (N_40738,N_35065,N_37769);
or U40739 (N_40739,N_37883,N_38769);
xor U40740 (N_40740,N_37547,N_39242);
and U40741 (N_40741,N_36815,N_35108);
nor U40742 (N_40742,N_37890,N_39909);
and U40743 (N_40743,N_38676,N_39879);
and U40744 (N_40744,N_37191,N_37161);
or U40745 (N_40745,N_35905,N_37212);
or U40746 (N_40746,N_38270,N_35438);
nand U40747 (N_40747,N_37993,N_35862);
or U40748 (N_40748,N_38141,N_36423);
xnor U40749 (N_40749,N_36608,N_39810);
xnor U40750 (N_40750,N_35458,N_38102);
or U40751 (N_40751,N_38604,N_36509);
and U40752 (N_40752,N_36338,N_39363);
or U40753 (N_40753,N_39853,N_39154);
or U40754 (N_40754,N_39894,N_39846);
nand U40755 (N_40755,N_39624,N_35958);
xor U40756 (N_40756,N_38829,N_39260);
or U40757 (N_40757,N_36659,N_35759);
or U40758 (N_40758,N_39086,N_39312);
or U40759 (N_40759,N_36300,N_36682);
nor U40760 (N_40760,N_37027,N_36425);
nor U40761 (N_40761,N_36442,N_38214);
and U40762 (N_40762,N_38220,N_38795);
or U40763 (N_40763,N_37057,N_37613);
or U40764 (N_40764,N_35707,N_36356);
nand U40765 (N_40765,N_37147,N_39997);
nor U40766 (N_40766,N_35084,N_39554);
and U40767 (N_40767,N_35537,N_39545);
xor U40768 (N_40768,N_38426,N_36208);
or U40769 (N_40769,N_39987,N_38645);
and U40770 (N_40770,N_35630,N_35423);
nand U40771 (N_40771,N_39581,N_36449);
xnor U40772 (N_40772,N_39902,N_36531);
nand U40773 (N_40773,N_39018,N_39056);
and U40774 (N_40774,N_35857,N_37930);
nand U40775 (N_40775,N_38796,N_38255);
and U40776 (N_40776,N_37311,N_36012);
nand U40777 (N_40777,N_36710,N_36794);
xnor U40778 (N_40778,N_37268,N_35992);
nor U40779 (N_40779,N_35204,N_38037);
and U40780 (N_40780,N_36559,N_39981);
and U40781 (N_40781,N_35963,N_36401);
or U40782 (N_40782,N_38111,N_38169);
xnor U40783 (N_40783,N_37847,N_38253);
or U40784 (N_40784,N_35325,N_35934);
and U40785 (N_40785,N_36021,N_35266);
nor U40786 (N_40786,N_38425,N_39249);
xnor U40787 (N_40787,N_37275,N_35839);
xor U40788 (N_40788,N_38713,N_35201);
and U40789 (N_40789,N_35800,N_36414);
nand U40790 (N_40790,N_36971,N_35745);
or U40791 (N_40791,N_36865,N_39670);
or U40792 (N_40792,N_35487,N_38700);
xor U40793 (N_40793,N_36205,N_37814);
nor U40794 (N_40794,N_37015,N_39873);
or U40795 (N_40795,N_38243,N_35122);
xor U40796 (N_40796,N_35471,N_37182);
nand U40797 (N_40797,N_36888,N_36063);
or U40798 (N_40798,N_37375,N_37549);
nand U40799 (N_40799,N_35094,N_38412);
and U40800 (N_40800,N_39166,N_38196);
nand U40801 (N_40801,N_37345,N_35771);
nor U40802 (N_40802,N_35617,N_39349);
nor U40803 (N_40803,N_36125,N_36486);
nor U40804 (N_40804,N_39025,N_36709);
and U40805 (N_40805,N_36574,N_38331);
and U40806 (N_40806,N_38797,N_37870);
and U40807 (N_40807,N_37752,N_36534);
and U40808 (N_40808,N_39699,N_36173);
nor U40809 (N_40809,N_35172,N_39402);
xor U40810 (N_40810,N_37851,N_37719);
and U40811 (N_40811,N_38738,N_39816);
and U40812 (N_40812,N_35966,N_37705);
xnor U40813 (N_40813,N_38846,N_36701);
xor U40814 (N_40814,N_37927,N_37817);
xnor U40815 (N_40815,N_39906,N_36868);
nor U40816 (N_40816,N_37676,N_35388);
and U40817 (N_40817,N_38531,N_35755);
nor U40818 (N_40818,N_39768,N_35506);
xor U40819 (N_40819,N_37962,N_35208);
xor U40820 (N_40820,N_38518,N_35774);
or U40821 (N_40821,N_36967,N_38086);
and U40822 (N_40822,N_35450,N_38522);
nand U40823 (N_40823,N_36148,N_39107);
xnor U40824 (N_40824,N_36106,N_39252);
nand U40825 (N_40825,N_39697,N_39435);
and U40826 (N_40826,N_39172,N_39840);
or U40827 (N_40827,N_37342,N_36572);
nand U40828 (N_40828,N_35277,N_39842);
nand U40829 (N_40829,N_39282,N_35434);
xor U40830 (N_40830,N_35060,N_39764);
nor U40831 (N_40831,N_38446,N_35752);
xnor U40832 (N_40832,N_39570,N_35258);
xnor U40833 (N_40833,N_35304,N_35542);
or U40834 (N_40834,N_39886,N_37773);
and U40835 (N_40835,N_39417,N_37293);
and U40836 (N_40836,N_36618,N_37013);
and U40837 (N_40837,N_35938,N_38063);
nand U40838 (N_40838,N_36589,N_39864);
and U40839 (N_40839,N_37258,N_37190);
and U40840 (N_40840,N_35396,N_39403);
xor U40841 (N_40841,N_38696,N_38593);
nand U40842 (N_40842,N_39609,N_37583);
nand U40843 (N_40843,N_37639,N_39573);
xnor U40844 (N_40844,N_38174,N_37438);
and U40845 (N_40845,N_35424,N_35381);
nor U40846 (N_40846,N_35170,N_38388);
nor U40847 (N_40847,N_35361,N_36301);
or U40848 (N_40848,N_37853,N_36605);
and U40849 (N_40849,N_38441,N_35467);
xnor U40850 (N_40850,N_36430,N_37952);
and U40851 (N_40851,N_38808,N_38990);
nand U40852 (N_40852,N_35112,N_35623);
nand U40853 (N_40853,N_37941,N_38026);
or U40854 (N_40854,N_36299,N_36385);
or U40855 (N_40855,N_35365,N_36912);
nand U40856 (N_40856,N_37327,N_39298);
xor U40857 (N_40857,N_35543,N_36724);
nor U40858 (N_40858,N_39550,N_37068);
xnor U40859 (N_40859,N_38208,N_36997);
or U40860 (N_40860,N_37026,N_39911);
xor U40861 (N_40861,N_38973,N_39082);
nor U40862 (N_40862,N_38711,N_38753);
xnor U40863 (N_40863,N_36702,N_37039);
or U40864 (N_40864,N_39716,N_38872);
nor U40865 (N_40865,N_35248,N_35474);
nor U40866 (N_40866,N_35123,N_39920);
xor U40867 (N_40867,N_35740,N_37688);
and U40868 (N_40868,N_36094,N_37385);
nor U40869 (N_40869,N_36804,N_38530);
nand U40870 (N_40870,N_36359,N_36374);
nand U40871 (N_40871,N_37577,N_36492);
and U40872 (N_40872,N_35884,N_37440);
and U40873 (N_40873,N_37333,N_37090);
xnor U40874 (N_40874,N_39666,N_39214);
and U40875 (N_40875,N_38385,N_36722);
and U40876 (N_40876,N_38694,N_36554);
or U40877 (N_40877,N_37344,N_36562);
and U40878 (N_40878,N_39476,N_36898);
and U40879 (N_40879,N_35893,N_36712);
nor U40880 (N_40880,N_37070,N_38395);
and U40881 (N_40881,N_39529,N_39279);
and U40882 (N_40882,N_35337,N_39190);
and U40883 (N_40883,N_35878,N_38798);
nand U40884 (N_40884,N_39384,N_39950);
nand U40885 (N_40885,N_36969,N_36460);
nand U40886 (N_40886,N_36556,N_36917);
or U40887 (N_40887,N_38755,N_35923);
and U40888 (N_40888,N_38478,N_37299);
xor U40889 (N_40889,N_39556,N_39565);
xor U40890 (N_40890,N_35273,N_37893);
nor U40891 (N_40891,N_36368,N_39723);
xnor U40892 (N_40892,N_39657,N_35635);
nand U40893 (N_40893,N_39240,N_36874);
xnor U40894 (N_40894,N_35937,N_36652);
and U40895 (N_40895,N_38693,N_37865);
and U40896 (N_40896,N_39420,N_35592);
xnor U40897 (N_40897,N_36930,N_36027);
nor U40898 (N_40898,N_37948,N_38379);
nand U40899 (N_40899,N_39192,N_37726);
xor U40900 (N_40900,N_35654,N_39057);
nand U40901 (N_40901,N_38238,N_39562);
xnor U40902 (N_40902,N_36075,N_35223);
and U40903 (N_40903,N_36073,N_38017);
and U40904 (N_40904,N_37315,N_38561);
nand U40905 (N_40905,N_39077,N_38232);
or U40906 (N_40906,N_37172,N_36705);
nand U40907 (N_40907,N_35196,N_37779);
or U40908 (N_40908,N_39313,N_37725);
xnor U40909 (N_40909,N_35901,N_38506);
nand U40910 (N_40910,N_39004,N_36853);
nor U40911 (N_40911,N_36433,N_37775);
xor U40912 (N_40912,N_38915,N_36836);
xnor U40913 (N_40913,N_39091,N_38874);
or U40914 (N_40914,N_36259,N_39157);
and U40915 (N_40915,N_39534,N_35622);
nor U40916 (N_40916,N_36089,N_36315);
nor U40917 (N_40917,N_38345,N_35292);
or U40918 (N_40918,N_38524,N_39475);
nor U40919 (N_40919,N_39275,N_37897);
nor U40920 (N_40920,N_37019,N_35906);
nand U40921 (N_40921,N_35364,N_38542);
or U40922 (N_40922,N_36399,N_38250);
or U40923 (N_40923,N_39533,N_37595);
xor U40924 (N_40924,N_38349,N_37921);
nor U40925 (N_40925,N_37269,N_37036);
nand U40926 (N_40926,N_37245,N_37524);
nand U40927 (N_40927,N_37040,N_35962);
xor U40928 (N_40928,N_37291,N_36257);
nand U40929 (N_40929,N_39948,N_39400);
and U40930 (N_40930,N_38609,N_35720);
xor U40931 (N_40931,N_35724,N_36084);
nor U40932 (N_40932,N_37397,N_37509);
and U40933 (N_40933,N_38540,N_37768);
nor U40934 (N_40934,N_39984,N_38563);
and U40935 (N_40935,N_37263,N_39797);
or U40936 (N_40936,N_39026,N_38131);
xnor U40937 (N_40937,N_38459,N_35885);
nand U40938 (N_40938,N_39888,N_36953);
and U40939 (N_40939,N_37784,N_36642);
nor U40940 (N_40940,N_37419,N_38774);
and U40941 (N_40941,N_38053,N_36946);
nand U40942 (N_40942,N_37416,N_35648);
xnor U40943 (N_40943,N_38050,N_37985);
and U40944 (N_40944,N_38909,N_36824);
xor U40945 (N_40945,N_35713,N_35141);
or U40946 (N_40946,N_38906,N_35744);
or U40947 (N_40947,N_38544,N_39290);
nor U40948 (N_40948,N_35876,N_37573);
or U40949 (N_40949,N_35532,N_38901);
nor U40950 (N_40950,N_38356,N_39068);
nand U40951 (N_40951,N_39036,N_39164);
xnor U40952 (N_40952,N_35943,N_35527);
and U40953 (N_40953,N_35529,N_38683);
and U40954 (N_40954,N_37911,N_36271);
nor U40955 (N_40955,N_39568,N_39978);
nor U40956 (N_40956,N_38007,N_39665);
xnor U40957 (N_40957,N_35750,N_35910);
nor U40958 (N_40958,N_36822,N_39654);
xor U40959 (N_40959,N_38706,N_39111);
or U40960 (N_40960,N_37030,N_35117);
nor U40961 (N_40961,N_38280,N_36870);
nand U40962 (N_40962,N_38773,N_38224);
and U40963 (N_40963,N_39431,N_37687);
xor U40964 (N_40964,N_35493,N_39860);
or U40965 (N_40965,N_38658,N_36767);
xor U40966 (N_40966,N_36335,N_35768);
xnor U40967 (N_40967,N_36664,N_39014);
nand U40968 (N_40968,N_39022,N_35712);
or U40969 (N_40969,N_35142,N_39932);
and U40970 (N_40970,N_37766,N_37984);
xor U40971 (N_40971,N_38878,N_39757);
nand U40972 (N_40972,N_37341,N_37490);
nor U40973 (N_40973,N_36895,N_38454);
and U40974 (N_40974,N_35531,N_36838);
xor U40975 (N_40975,N_38924,N_35482);
xor U40976 (N_40976,N_39090,N_37310);
nor U40977 (N_40977,N_38313,N_35125);
xor U40978 (N_40978,N_39571,N_38432);
nand U40979 (N_40979,N_36482,N_39651);
nand U40980 (N_40980,N_38207,N_37588);
xor U40981 (N_40981,N_35977,N_37171);
and U40982 (N_40982,N_37791,N_37520);
or U40983 (N_40983,N_36052,N_36864);
and U40984 (N_40984,N_39346,N_37376);
nor U40985 (N_40985,N_39912,N_39918);
nand U40986 (N_40986,N_37044,N_36038);
xnor U40987 (N_40987,N_39399,N_37323);
or U40988 (N_40988,N_38137,N_39104);
nor U40989 (N_40989,N_35782,N_37229);
xnor U40990 (N_40990,N_38541,N_37935);
and U40991 (N_40991,N_36846,N_39044);
or U40992 (N_40992,N_35429,N_37141);
and U40993 (N_40993,N_36573,N_38734);
xnor U40994 (N_40994,N_35908,N_35556);
nand U40995 (N_40995,N_38486,N_35047);
nand U40996 (N_40996,N_38048,N_39041);
xor U40997 (N_40997,N_37348,N_39839);
nand U40998 (N_40998,N_39438,N_36966);
nor U40999 (N_40999,N_35217,N_37227);
or U41000 (N_41000,N_37193,N_38126);
nand U41001 (N_41001,N_36192,N_35970);
nor U41002 (N_41002,N_35494,N_35632);
nor U41003 (N_41003,N_35696,N_37078);
and U41004 (N_41004,N_37696,N_35357);
xor U41005 (N_41005,N_35179,N_35784);
xor U41006 (N_41006,N_38021,N_35561);
or U41007 (N_41007,N_37483,N_35023);
or U41008 (N_41008,N_35078,N_38147);
xnor U41009 (N_41009,N_38129,N_39991);
and U41010 (N_41010,N_38386,N_39588);
or U41011 (N_41011,N_38218,N_38373);
nor U41012 (N_41012,N_35033,N_35636);
xnor U41013 (N_41013,N_38124,N_39052);
nor U41014 (N_41014,N_38615,N_37502);
nand U41015 (N_41015,N_37934,N_37873);
xor U41016 (N_41016,N_36201,N_36294);
or U41017 (N_41017,N_38077,N_36249);
or U41018 (N_41018,N_37849,N_37654);
nand U41019 (N_41019,N_39676,N_37243);
nor U41020 (N_41020,N_37432,N_39023);
and U41021 (N_41021,N_38027,N_38716);
and U41022 (N_41022,N_39253,N_39962);
xnor U41023 (N_41023,N_37326,N_35333);
xnor U41024 (N_41024,N_35797,N_35145);
or U41025 (N_41025,N_37095,N_39930);
or U41026 (N_41026,N_39787,N_39012);
or U41027 (N_41027,N_36776,N_38380);
xnor U41028 (N_41028,N_39103,N_39507);
nor U41029 (N_41029,N_39339,N_39610);
nor U41030 (N_41030,N_39003,N_36771);
nand U41031 (N_41031,N_35513,N_36900);
and U41032 (N_41032,N_35872,N_38249);
or U41033 (N_41033,N_36921,N_38776);
xor U41034 (N_41034,N_35914,N_38078);
and U41035 (N_41035,N_38470,N_35194);
or U41036 (N_41036,N_38352,N_38069);
nor U41037 (N_41037,N_36943,N_38494);
or U41038 (N_41038,N_35897,N_38422);
and U41039 (N_41039,N_35069,N_39896);
nand U41040 (N_41040,N_36210,N_38545);
xnor U41041 (N_41041,N_36781,N_36651);
or U41042 (N_41042,N_35298,N_37552);
nand U41043 (N_41043,N_36945,N_39189);
nor U41044 (N_41044,N_39897,N_35579);
nor U41045 (N_41045,N_39378,N_37494);
or U41046 (N_41046,N_36159,N_39693);
xnor U41047 (N_41047,N_35156,N_39733);
xnor U41048 (N_41048,N_35748,N_37121);
nand U41049 (N_41049,N_39785,N_39673);
nor U41050 (N_41050,N_37468,N_35530);
and U41051 (N_41051,N_39783,N_38656);
nand U41052 (N_41052,N_35475,N_38298);
nor U41053 (N_41053,N_38904,N_37834);
xnor U41054 (N_41054,N_35559,N_37097);
or U41055 (N_41055,N_38387,N_36955);
and U41056 (N_41056,N_38822,N_39947);
xnor U41057 (N_41057,N_35741,N_38320);
and U41058 (N_41058,N_37066,N_35538);
or U41059 (N_41059,N_39072,N_39396);
xnor U41060 (N_41060,N_37680,N_36386);
xnor U41061 (N_41061,N_35887,N_39551);
or U41062 (N_41062,N_38510,N_35484);
xor U41063 (N_41063,N_35553,N_35733);
and U41064 (N_41064,N_38838,N_37744);
or U41065 (N_41065,N_35960,N_35254);
or U41066 (N_41066,N_38226,N_39721);
or U41067 (N_41067,N_39224,N_38464);
or U41068 (N_41068,N_36716,N_35667);
and U41069 (N_41069,N_38664,N_39821);
xor U41070 (N_41070,N_35178,N_35174);
nand U41071 (N_41071,N_35399,N_37544);
nor U41072 (N_41072,N_37153,N_38319);
nand U41073 (N_41073,N_37717,N_36458);
xor U41074 (N_41074,N_37961,N_37368);
nand U41075 (N_41075,N_38945,N_39070);
and U41076 (N_41076,N_35138,N_37774);
or U41077 (N_41077,N_39499,N_37405);
xnor U41078 (N_41078,N_36083,N_35804);
xor U41079 (N_41079,N_37923,N_37084);
nand U41080 (N_41080,N_39010,N_38058);
xor U41081 (N_41081,N_38194,N_37644);
and U41082 (N_41082,N_36028,N_38639);
or U41083 (N_41083,N_38782,N_35849);
nand U41084 (N_41084,N_36560,N_36077);
or U41085 (N_41085,N_35829,N_36044);
nand U41086 (N_41086,N_39490,N_39965);
xnor U41087 (N_41087,N_38083,N_39126);
nor U41088 (N_41088,N_36258,N_35541);
and U41089 (N_41089,N_35323,N_35229);
nand U41090 (N_41090,N_39559,N_37109);
nand U41091 (N_41091,N_36889,N_35336);
nor U41092 (N_41092,N_37281,N_38369);
and U41093 (N_41093,N_35874,N_35441);
nor U41094 (N_41094,N_38210,N_36376);
and U41095 (N_41095,N_37364,N_39409);
or U41096 (N_41096,N_35618,N_37543);
and U41097 (N_41097,N_35147,N_38605);
and U41098 (N_41098,N_38930,N_36286);
or U41099 (N_41099,N_38647,N_37968);
or U41100 (N_41100,N_36537,N_35286);
or U41101 (N_41101,N_39791,N_38166);
nor U41102 (N_41102,N_37178,N_36925);
nor U41103 (N_41103,N_35359,N_36561);
or U41104 (N_41104,N_37724,N_37476);
nor U41105 (N_41105,N_36464,N_39270);
or U41106 (N_41106,N_36229,N_36375);
or U41107 (N_41107,N_36820,N_36343);
nand U41108 (N_41108,N_39430,N_39814);
nor U41109 (N_41109,N_36209,N_38553);
or U41110 (N_41110,N_36296,N_39505);
nor U41111 (N_41111,N_37173,N_36782);
nor U41112 (N_41112,N_39589,N_38428);
or U41113 (N_41113,N_37456,N_39649);
or U41114 (N_41114,N_35781,N_37077);
or U41115 (N_41115,N_36532,N_38274);
or U41116 (N_41116,N_36097,N_39019);
nand U41117 (N_41117,N_35965,N_38892);
or U41118 (N_41118,N_39942,N_39200);
or U41119 (N_41119,N_35200,N_37863);
or U41120 (N_41120,N_37631,N_39035);
xnor U41121 (N_41121,N_38662,N_36196);
nand U41122 (N_41122,N_36086,N_38527);
and U41123 (N_41123,N_36287,N_35497);
xnor U41124 (N_41124,N_35675,N_38480);
nor U41125 (N_41125,N_38851,N_36919);
and U41126 (N_41126,N_37089,N_39552);
or U41127 (N_41127,N_35068,N_38267);
and U41128 (N_41128,N_39415,N_38627);
or U41129 (N_41129,N_37825,N_39584);
or U41130 (N_41130,N_38461,N_38636);
and U41131 (N_41131,N_36996,N_35703);
nand U41132 (N_41132,N_36787,N_36495);
nand U41133 (N_41133,N_36586,N_39097);
and U41134 (N_41134,N_36535,N_35589);
and U41135 (N_41135,N_36610,N_36104);
nor U41136 (N_41136,N_39822,N_37894);
or U41137 (N_41137,N_37433,N_38957);
nand U41138 (N_41138,N_38509,N_36427);
xnor U41139 (N_41139,N_37932,N_39447);
nor U41140 (N_41140,N_36500,N_37958);
xnor U41141 (N_41141,N_39859,N_38916);
xnor U41142 (N_41142,N_39277,N_37830);
and U41143 (N_41143,N_39433,N_39767);
and U41144 (N_41144,N_35792,N_36899);
nor U41145 (N_41145,N_35896,N_39908);
nand U41146 (N_41146,N_36956,N_36805);
nor U41147 (N_41147,N_38357,N_35387);
and U41148 (N_41148,N_36410,N_37906);
nand U41149 (N_41149,N_38547,N_36708);
xnor U41150 (N_41150,N_35525,N_37973);
and U41151 (N_41151,N_37241,N_35621);
or U41152 (N_41152,N_38862,N_36617);
nand U41153 (N_41153,N_35933,N_36377);
xor U41154 (N_41154,N_35779,N_35274);
or U41155 (N_41155,N_38074,N_36378);
nor U41156 (N_41156,N_36451,N_38666);
nand U41157 (N_41157,N_39045,N_36578);
and U41158 (N_41158,N_38982,N_37175);
nor U41159 (N_41159,N_35595,N_37565);
and U41160 (N_41160,N_37839,N_38285);
or U41161 (N_41161,N_37833,N_38923);
xnor U41162 (N_41162,N_35157,N_38836);
nor U41163 (N_41163,N_35137,N_37571);
and U41164 (N_41164,N_39283,N_35449);
xor U41165 (N_41165,N_36041,N_39487);
or U41166 (N_41166,N_36329,N_38496);
xor U41167 (N_41167,N_35832,N_39726);
or U41168 (N_41168,N_36575,N_38114);
nand U41169 (N_41169,N_38688,N_39272);
and U41170 (N_41170,N_35310,N_37508);
xor U41171 (N_41171,N_37986,N_38896);
nand U41172 (N_41172,N_37429,N_37648);
nor U41173 (N_41173,N_37743,N_37608);
nor U41174 (N_41174,N_37628,N_37114);
nor U41175 (N_41175,N_37392,N_37527);
nand U41176 (N_41176,N_39477,N_37626);
nand U41177 (N_41177,N_38764,N_39361);
and U41178 (N_41178,N_39040,N_36759);
and U41179 (N_41179,N_35528,N_39695);
nand U41180 (N_41180,N_37905,N_37125);
nor U41181 (N_41181,N_37138,N_39983);
xnor U41182 (N_41182,N_35421,N_39175);
nand U41183 (N_41183,N_35787,N_39437);
nand U41184 (N_41184,N_37778,N_39042);
nand U41185 (N_41185,N_39605,N_39663);
and U41186 (N_41186,N_39049,N_37447);
xnor U41187 (N_41187,N_36689,N_39904);
and U41188 (N_41188,N_37451,N_38632);
or U41189 (N_41189,N_39913,N_37261);
and U41190 (N_41190,N_35634,N_35803);
nor U41191 (N_41191,N_35372,N_35993);
and U41192 (N_41192,N_36602,N_38234);
nor U41193 (N_41193,N_38842,N_35936);
xor U41194 (N_41194,N_39986,N_37297);
xnor U41195 (N_41195,N_38445,N_35247);
or U41196 (N_41196,N_36247,N_35099);
and U41197 (N_41197,N_36727,N_39718);
nand U41198 (N_41198,N_39101,N_35455);
and U41199 (N_41199,N_39650,N_39945);
or U41200 (N_41200,N_36854,N_39223);
and U41201 (N_41201,N_39871,N_38715);
nand U41202 (N_41202,N_37422,N_38297);
nand U41203 (N_41203,N_35400,N_35739);
nand U41204 (N_41204,N_37748,N_36693);
nand U41205 (N_41205,N_39577,N_37799);
and U41206 (N_41206,N_39146,N_37522);
and U41207 (N_41207,N_39379,N_39108);
xor U41208 (N_41208,N_39258,N_38416);
and U41209 (N_41209,N_37939,N_38127);
or U41210 (N_41210,N_38635,N_36883);
nand U41211 (N_41211,N_39741,N_38177);
and U41212 (N_41212,N_35327,N_37374);
and U41213 (N_41213,N_35098,N_36734);
nand U41214 (N_41214,N_37580,N_35376);
xor U41215 (N_41215,N_36714,N_37810);
nor U41216 (N_41216,N_38899,N_38852);
and U41217 (N_41217,N_35601,N_37535);
nor U41218 (N_41218,N_35511,N_36484);
nor U41219 (N_41219,N_38768,N_35662);
xnor U41220 (N_41220,N_35749,N_38168);
xor U41221 (N_41221,N_36519,N_35240);
nand U41222 (N_41222,N_35860,N_35126);
xor U41223 (N_41223,N_36107,N_38650);
or U41224 (N_41224,N_37067,N_35206);
and U41225 (N_41225,N_36186,N_35271);
and U41226 (N_41226,N_38477,N_35002);
and U41227 (N_41227,N_39687,N_35602);
or U41228 (N_41228,N_35358,N_36251);
and U41229 (N_41229,N_37529,N_35279);
nand U41230 (N_41230,N_38978,N_35664);
or U41231 (N_41231,N_39079,N_39080);
and U41232 (N_41232,N_38434,N_38931);
nand U41233 (N_41233,N_37457,N_37436);
and U41234 (N_41234,N_37947,N_36099);
nand U41235 (N_41235,N_35853,N_38869);
or U41236 (N_41236,N_37995,N_37764);
nand U41237 (N_41237,N_36944,N_39317);
nand U41238 (N_41238,N_38718,N_38818);
or U41239 (N_41239,N_36152,N_37041);
nand U41240 (N_41240,N_39169,N_38105);
and U41241 (N_41241,N_35572,N_38708);
nor U41242 (N_41242,N_37630,N_36663);
xor U41243 (N_41243,N_38737,N_35778);
or U41244 (N_41244,N_39881,N_38724);
and U41245 (N_41245,N_36587,N_39429);
xor U41246 (N_41246,N_36700,N_38128);
xnor U41247 (N_41247,N_35565,N_36672);
xor U41248 (N_41248,N_38123,N_35922);
nand U41249 (N_41249,N_38080,N_37226);
or U41250 (N_41250,N_36843,N_35048);
or U41251 (N_41251,N_36292,N_36457);
xor U41252 (N_41252,N_36020,N_36122);
xor U41253 (N_41253,N_36225,N_36933);
nand U41254 (N_41254,N_38444,N_35583);
and U41255 (N_41255,N_39640,N_39321);
xor U41256 (N_41256,N_38590,N_36666);
nor U41257 (N_41257,N_39061,N_37612);
nor U41258 (N_41258,N_39806,N_37448);
nor U41259 (N_41259,N_39659,N_37108);
xnor U41260 (N_41260,N_35146,N_36365);
and U41261 (N_41261,N_35297,N_38005);
or U41262 (N_41262,N_36216,N_35490);
or U41263 (N_41263,N_37891,N_39974);
nand U41264 (N_41264,N_35873,N_35089);
or U41265 (N_41265,N_39265,N_39278);
and U41266 (N_41266,N_38323,N_37678);
or U41267 (N_41267,N_38101,N_39548);
xor U41268 (N_41268,N_35230,N_35015);
xor U41269 (N_41269,N_39543,N_38150);
and U41270 (N_41270,N_37224,N_37994);
xnor U41271 (N_41271,N_38870,N_38338);
or U41272 (N_41272,N_36281,N_37575);
xnor U41273 (N_41273,N_35677,N_38511);
nor U41274 (N_41274,N_37407,N_35121);
or U41275 (N_41275,N_39592,N_35825);
nand U41276 (N_41276,N_39900,N_38429);
xnor U41277 (N_41277,N_38089,N_38633);
or U41278 (N_41278,N_37925,N_39145);
and U41279 (N_41279,N_38599,N_38554);
and U41280 (N_41280,N_38163,N_39391);
nand U41281 (N_41281,N_35503,N_39171);
nor U41282 (N_41282,N_38286,N_36408);
nand U41283 (N_41283,N_35928,N_37443);
nand U41284 (N_41284,N_37154,N_36645);
nor U41285 (N_41285,N_37445,N_39854);
xor U41286 (N_41286,N_39995,N_36227);
and U41287 (N_41287,N_38767,N_35587);
nand U41288 (N_41288,N_35658,N_37913);
nand U41289 (N_41289,N_38550,N_35233);
xor U41290 (N_41290,N_39135,N_38787);
xnor U41291 (N_41291,N_37943,N_37731);
nor U41292 (N_41292,N_38841,N_35354);
or U41293 (N_41293,N_35356,N_38933);
or U41294 (N_41294,N_37981,N_35491);
and U41295 (N_41295,N_38959,N_35166);
nand U41296 (N_41296,N_39789,N_39585);
nand U41297 (N_41297,N_36057,N_37219);
or U41298 (N_41298,N_35930,N_37504);
nand U41299 (N_41299,N_35244,N_37889);
xnor U41300 (N_41300,N_35738,N_39481);
nor U41301 (N_41301,N_39990,N_38621);
and U41302 (N_41302,N_38728,N_39626);
nand U41303 (N_41303,N_39212,N_37179);
or U41304 (N_41304,N_39858,N_38330);
or U41305 (N_41305,N_38466,N_36591);
xnor U41306 (N_41306,N_38723,N_38217);
xnor U41307 (N_41307,N_39256,N_36690);
xor U41308 (N_41308,N_38730,N_36381);
xnor U41309 (N_41309,N_38440,N_37645);
and U41310 (N_41310,N_39000,N_39629);
nand U41311 (N_41311,N_37017,N_38160);
nand U41312 (N_41312,N_37637,N_39193);
nand U41313 (N_41313,N_38889,N_39704);
nand U41314 (N_41314,N_37320,N_36786);
and U41315 (N_41315,N_38900,N_38614);
or U41316 (N_41316,N_39761,N_35833);
nand U41317 (N_41317,N_39979,N_38879);
nor U41318 (N_41318,N_39364,N_35704);
and U41319 (N_41319,N_36088,N_37579);
or U41320 (N_41320,N_35524,N_38472);
and U41321 (N_41321,N_35346,N_36371);
nor U41322 (N_41322,N_35581,N_36470);
nand U41323 (N_41323,N_38989,N_35160);
nor U41324 (N_41324,N_39798,N_36972);
nand U41325 (N_41325,N_39210,N_35368);
or U41326 (N_41326,N_36274,N_38393);
and U41327 (N_41327,N_35409,N_37316);
nand U41328 (N_41328,N_39063,N_37062);
nor U41329 (N_41329,N_37312,N_39793);
xor U41330 (N_41330,N_39085,N_35465);
xnor U41331 (N_41331,N_36120,N_39740);
xor U41332 (N_41332,N_35980,N_38312);
xor U41333 (N_41333,N_38771,N_36501);
xnor U41334 (N_41334,N_38343,N_35788);
nor U41335 (N_41335,N_36290,N_37683);
nand U41336 (N_41336,N_36876,N_39485);
nor U41337 (N_41337,N_39287,N_36250);
nor U41338 (N_41338,N_37681,N_36151);
nand U41339 (N_41339,N_36323,N_39621);
nor U41340 (N_41340,N_39102,N_39480);
xor U41341 (N_41341,N_38502,N_37162);
and U41342 (N_41342,N_35264,N_35149);
nand U41343 (N_41343,N_36629,N_36085);
nand U41344 (N_41344,N_38772,N_38914);
xor U41345 (N_41345,N_35335,N_38413);
nand U41346 (N_41346,N_36616,N_38161);
nor U41347 (N_41347,N_38646,N_36291);
nand U41348 (N_41348,N_37592,N_38408);
xor U41349 (N_41349,N_39468,N_36928);
xor U41350 (N_41350,N_37493,N_35605);
nor U41351 (N_41351,N_36406,N_35827);
or U41352 (N_41352,N_39778,N_36949);
nor U41353 (N_41353,N_37694,N_39739);
xor U41354 (N_41354,N_39594,N_36504);
and U41355 (N_41355,N_37665,N_35627);
nand U41356 (N_41356,N_36894,N_36970);
and U41357 (N_41357,N_38476,N_35606);
and U41358 (N_41358,N_39259,N_39955);
or U41359 (N_41359,N_37252,N_38322);
nand U41360 (N_41360,N_37393,N_37733);
xor U41361 (N_41361,N_36095,N_35576);
and U41362 (N_41362,N_38358,N_36583);
and U41363 (N_41363,N_37843,N_36694);
nor U41364 (N_41364,N_36760,N_38401);
nor U41365 (N_41365,N_38115,N_38481);
and U41366 (N_41366,N_38329,N_35017);
or U41367 (N_41367,N_37640,N_37710);
nand U41368 (N_41368,N_36333,N_37920);
and U41369 (N_41369,N_36434,N_36882);
nand U41370 (N_41370,N_37584,N_39226);
or U41371 (N_41371,N_39857,N_37167);
nand U41372 (N_41372,N_36070,N_39009);
xor U41373 (N_41373,N_39046,N_38022);
nor U41374 (N_41374,N_35590,N_38819);
nor U41375 (N_41375,N_36262,N_37780);
and U41376 (N_41376,N_38104,N_35352);
xnor U41377 (N_41377,N_38955,N_38709);
xor U41378 (N_41378,N_38742,N_38668);
xnor U41379 (N_41379,N_35540,N_36726);
nor U41380 (N_41380,N_35397,N_36325);
or U41381 (N_41381,N_38436,N_36932);
nor U41382 (N_41382,N_38516,N_37371);
xor U41383 (N_41383,N_38687,N_38248);
or U41384 (N_41384,N_37854,N_38539);
and U41385 (N_41385,N_38110,N_39619);
nor U41386 (N_41386,N_35961,N_36837);
nand U41387 (N_41387,N_35308,N_37218);
or U41388 (N_41388,N_38018,N_38548);
and U41389 (N_41389,N_35045,N_39301);
nand U41390 (N_41390,N_35615,N_35044);
nor U41391 (N_41391,N_35443,N_39660);
xnor U41392 (N_41392,N_38939,N_38966);
nand U41393 (N_41393,N_36772,N_35573);
nand U41394 (N_41394,N_35185,N_38942);
nand U41395 (N_41395,N_37888,N_35909);
xnor U41396 (N_41396,N_38748,N_39647);
nand U41397 (N_41397,N_38680,N_37112);
nand U41398 (N_41398,N_35192,N_36112);
and U41399 (N_41399,N_36533,N_37882);
and U41400 (N_41400,N_37525,N_36841);
nand U41401 (N_41401,N_35162,N_37650);
nand U41402 (N_41402,N_38963,N_39618);
nand U41403 (N_41403,N_35953,N_38036);
nand U41404 (N_41404,N_39555,N_36742);
and U41405 (N_41405,N_37832,N_38781);
and U41406 (N_41406,N_36154,N_36066);
and U41407 (N_41407,N_38701,N_35063);
or U41408 (N_41408,N_37684,N_37727);
or U41409 (N_41409,N_37470,N_39219);
nand U41410 (N_41410,N_36755,N_36082);
xnor U41411 (N_41411,N_38465,N_35772);
or U41412 (N_41412,N_38749,N_36817);
xor U41413 (N_41413,N_36698,N_38907);
and U41414 (N_41414,N_35578,N_36017);
nand U41415 (N_41415,N_37620,N_35198);
nor U41416 (N_41416,N_36189,N_36069);
and U41417 (N_41417,N_36670,N_35824);
nand U41418 (N_41418,N_35383,N_35760);
and U41419 (N_41419,N_37287,N_39615);
nor U41420 (N_41420,N_37386,N_39933);
and U41421 (N_41421,N_39165,N_35916);
or U41422 (N_41422,N_39831,N_38951);
xor U41423 (N_41423,N_36798,N_39060);
and U41424 (N_41424,N_36891,N_39865);
nor U41425 (N_41425,N_35377,N_36619);
nand U41426 (N_41426,N_38411,N_36968);
nor U41427 (N_41427,N_35551,N_38679);
xor U41428 (N_41428,N_36372,N_35912);
xnor U41429 (N_41429,N_37144,N_37410);
and U41430 (N_41430,N_39377,N_35913);
nor U41431 (N_41431,N_35398,N_38864);
nor U41432 (N_41432,N_38293,N_36857);
xor U41433 (N_41433,N_36450,N_35948);
and U41434 (N_41434,N_38013,N_35507);
or U41435 (N_41435,N_36124,N_38671);
and U41436 (N_41436,N_37747,N_37656);
or U41437 (N_41437,N_38140,N_39114);
and U41438 (N_41438,N_35700,N_37321);
nor U41439 (N_41439,N_36144,N_36061);
or U41440 (N_41440,N_39406,N_35921);
nand U41441 (N_41441,N_38992,N_37767);
nand U41442 (N_41442,N_38689,N_35757);
xnor U41443 (N_41443,N_35433,N_37439);
and U41444 (N_41444,N_39633,N_35235);
or U41445 (N_41445,N_39110,N_39683);
nor U41446 (N_41446,N_39940,N_38629);
and U41447 (N_41447,N_36415,N_37647);
nor U41448 (N_41448,N_39150,N_39513);
or U41449 (N_41449,N_37720,N_36746);
xnor U41450 (N_41450,N_36126,N_37061);
nor U41451 (N_41451,N_38949,N_36585);
xor U41452 (N_41452,N_35731,N_39043);
and U41453 (N_41453,N_38305,N_39569);
nor U41454 (N_41454,N_35021,N_35373);
or U41455 (N_41455,N_39491,N_35165);
and U41456 (N_41456,N_35898,N_36625);
nand U41457 (N_41457,N_37009,N_37828);
or U41458 (N_41458,N_38471,N_37605);
nor U41459 (N_41459,N_38273,N_36142);
and U41460 (N_41460,N_39129,N_39105);
nor U41461 (N_41461,N_35813,N_37058);
or U41462 (N_41462,N_38732,N_39959);
and U41463 (N_41463,N_37373,N_39801);
xnor U41464 (N_41464,N_38720,N_36040);
nand U41465 (N_41465,N_38263,N_36988);
or U41466 (N_41466,N_36182,N_37811);
or U41467 (N_41467,N_37149,N_38090);
or U41468 (N_41468,N_38254,N_37949);
and U41469 (N_41469,N_36187,N_35945);
nor U41470 (N_41470,N_39034,N_37928);
nor U41471 (N_41471,N_37265,N_38817);
nand U41472 (N_41472,N_36530,N_38221);
nor U41473 (N_41473,N_37037,N_36539);
nor U41474 (N_41474,N_36237,N_36160);
nand U41475 (N_41475,N_35894,N_38431);
xor U41476 (N_41476,N_39703,N_38182);
nand U41477 (N_41477,N_38180,N_36074);
nand U41478 (N_41478,N_38023,N_37598);
xor U41479 (N_41479,N_38351,N_35057);
or U41480 (N_41480,N_35022,N_36978);
or U41481 (N_41481,N_39109,N_35132);
or U41482 (N_41482,N_37856,N_37729);
nand U41483 (N_41483,N_36171,N_39850);
or U41484 (N_41484,N_35081,N_35940);
nand U41485 (N_41485,N_37636,N_37497);
nand U41486 (N_41486,N_36493,N_36703);
nand U41487 (N_41487,N_37503,N_36989);
xnor U41488 (N_41488,N_37414,N_36223);
nor U41489 (N_41489,N_39535,N_37969);
or U41490 (N_41490,N_36179,N_35795);
and U41491 (N_41491,N_39066,N_38596);
or U41492 (N_41492,N_39123,N_39292);
nand U41493 (N_41493,N_37723,N_35679);
and U41494 (N_41494,N_37858,N_38394);
nor U41495 (N_41495,N_35153,N_36036);
nor U41496 (N_41496,N_38227,N_39446);
nand U41497 (N_41497,N_39250,N_36934);
or U41498 (N_41498,N_36010,N_36990);
xor U41499 (N_41499,N_37534,N_35130);
nand U41500 (N_41500,N_38608,N_36858);
or U41501 (N_41501,N_37500,N_39271);
or U41502 (N_41502,N_35684,N_35055);
or U41503 (N_41503,N_38584,N_39319);
and U41504 (N_41504,N_39194,N_35115);
nand U41505 (N_41505,N_39750,N_38192);
nor U41506 (N_41506,N_38469,N_37668);
or U41507 (N_41507,N_39371,N_38231);
xnor U41508 (N_41508,N_39656,N_38641);
and U41509 (N_41509,N_36150,N_37907);
and U41510 (N_41510,N_39998,N_37878);
nor U41511 (N_41511,N_36580,N_36510);
xnor U41512 (N_41512,N_37122,N_35282);
nand U41513 (N_41513,N_38039,N_38857);
or U41514 (N_41514,N_38447,N_35516);
and U41515 (N_41515,N_36475,N_35413);
nor U41516 (N_41516,N_35075,N_37796);
and U41517 (N_41517,N_36632,N_36047);
nor U41518 (N_41518,N_37821,N_37228);
or U41519 (N_41519,N_36905,N_37996);
nand U41520 (N_41520,N_39153,N_35582);
nand U41521 (N_41521,N_36222,N_39508);
nand U41522 (N_41522,N_39341,N_37511);
or U41523 (N_41523,N_37691,N_37110);
and U41524 (N_41524,N_36740,N_39796);
and U41525 (N_41525,N_35257,N_38579);
nor U41526 (N_41526,N_38965,N_35593);
nor U41527 (N_41527,N_38883,N_38558);
or U41528 (N_41528,N_39779,N_35472);
nor U41529 (N_41529,N_37313,N_38033);
nor U41530 (N_41530,N_35676,N_39262);
xnor U41531 (N_41531,N_38941,N_36697);
nor U41532 (N_41532,N_36090,N_37674);
or U41533 (N_41533,N_38845,N_35732);
or U41534 (N_41534,N_35389,N_36391);
and U41535 (N_41535,N_37274,N_37561);
nor U41536 (N_41536,N_35628,N_39369);
and U41537 (N_41537,N_35339,N_37682);
or U41538 (N_41538,N_36655,N_39074);
or U41539 (N_41539,N_35734,N_39088);
nor U41540 (N_41540,N_39928,N_39495);
xor U41541 (N_41541,N_35416,N_38549);
and U41542 (N_41542,N_36568,N_36829);
and U41543 (N_41543,N_38112,N_35326);
nor U41544 (N_41544,N_35899,N_37318);
nor U41545 (N_41545,N_36276,N_37018);
nand U41546 (N_41546,N_36278,N_37292);
nor U41547 (N_41547,N_37180,N_36646);
nor U41548 (N_41548,N_38744,N_35355);
nand U41549 (N_41549,N_36413,N_36031);
nand U41550 (N_41550,N_36732,N_39675);
or U41551 (N_41551,N_37761,N_38766);
or U41552 (N_41552,N_37762,N_35718);
nand U41553 (N_41553,N_35390,N_39464);
nor U41554 (N_41554,N_38837,N_36577);
and U41555 (N_41555,N_36447,N_36180);
nor U41556 (N_41556,N_36110,N_36161);
and U41557 (N_41557,N_38360,N_39225);
and U41558 (N_41558,N_39712,N_38019);
xnor U41559 (N_41559,N_38437,N_39281);
nand U41560 (N_41560,N_36821,N_37635);
nand U41561 (N_41561,N_37279,N_38088);
nand U41562 (N_41562,N_38304,N_37526);
nor U41563 (N_41563,N_38569,N_37123);
or U41564 (N_41564,N_35850,N_38359);
nand U41565 (N_41565,N_38289,N_38811);
or U41566 (N_41566,N_36764,N_36799);
or U41567 (N_41567,N_37959,N_39089);
or U41568 (N_41568,N_36242,N_39517);
nand U41569 (N_41569,N_35224,N_39059);
xnor U41570 (N_41570,N_36488,N_38324);
or U41571 (N_41571,N_36138,N_39328);
nor U41572 (N_41572,N_35252,N_38761);
or U41573 (N_41573,N_39580,N_35309);
and U41574 (N_41574,N_36282,N_38954);
xnor U41575 (N_41575,N_39297,N_39365);
nand U41576 (N_41576,N_37232,N_39685);
nand U41577 (N_41577,N_37838,N_35454);
or U41578 (N_41578,N_38760,N_39772);
nand U41579 (N_41579,N_36916,N_35834);
nand U41580 (N_41580,N_37651,N_38337);
nor U41581 (N_41581,N_37960,N_36269);
nor U41582 (N_41582,N_37972,N_35030);
nand U41583 (N_41583,N_35722,N_39178);
nand U41584 (N_41584,N_39837,N_39112);
xor U41585 (N_41585,N_36926,N_37354);
and U41586 (N_41586,N_37151,N_36334);
xor U41587 (N_41587,N_37603,N_37409);
or U41588 (N_41588,N_39985,N_37454);
nor U41589 (N_41589,N_37236,N_38125);
and U41590 (N_41590,N_37908,N_39322);
and U41591 (N_41591,N_36596,N_36252);
nor U41592 (N_41592,N_39817,N_38834);
and U41593 (N_41593,N_39374,N_35486);
or U41594 (N_41594,N_36404,N_35479);
nand U41595 (N_41595,N_37284,N_37197);
or U41596 (N_41596,N_39820,N_36068);
nor U41597 (N_41597,N_37967,N_36071);
and U41598 (N_41598,N_36485,N_39462);
and U41599 (N_41599,N_37898,N_36650);
and U41600 (N_41600,N_36008,N_38736);
nand U41601 (N_41601,N_36869,N_39054);
or U41602 (N_41602,N_36636,N_39001);
or U41603 (N_41603,N_37060,N_35103);
nand U41604 (N_41604,N_39345,N_37542);
nor U41605 (N_41605,N_38937,N_35990);
xor U41606 (N_41606,N_35521,N_38325);
and U41607 (N_41607,N_37477,N_35941);
or U41608 (N_41608,N_39471,N_39895);
and U41609 (N_41609,N_37196,N_39007);
and U41610 (N_41610,N_38075,N_36745);
nor U41611 (N_41611,N_36272,N_35485);
nor U41612 (N_41612,N_35767,N_36137);
nor U41613 (N_41613,N_35432,N_38961);
xor U41614 (N_41614,N_39849,N_35790);
and U41615 (N_41615,N_38029,N_37980);
nor U41616 (N_41616,N_36108,N_39845);
xor U41617 (N_41617,N_39293,N_37572);
nand U41618 (N_41618,N_39826,N_39302);
or U41619 (N_41619,N_35238,N_35216);
xor U41620 (N_41620,N_39149,N_36713);
or U41621 (N_41621,N_35199,N_35054);
and U41622 (N_41622,N_36677,N_35875);
or U41623 (N_41623,N_36570,N_37111);
xor U41624 (N_41624,N_39327,N_39557);
nor U41625 (N_41625,N_39308,N_37850);
nor U41626 (N_41626,N_38893,N_35688);
nor U41627 (N_41627,N_39173,N_39285);
or U41628 (N_41628,N_38998,N_38968);
or U41629 (N_41629,N_39299,N_37307);
nor U41630 (N_41630,N_36673,N_37113);
nand U41631 (N_41631,N_37560,N_35695);
and U41632 (N_41632,N_36456,N_37365);
and U41633 (N_41633,N_36590,N_37124);
nor U41634 (N_41634,N_35181,N_39008);
or U41635 (N_41635,N_38866,N_38016);
nand U41636 (N_41636,N_36630,N_37615);
nand U41637 (N_41637,N_37826,N_35837);
nor U41638 (N_41638,N_39134,N_35019);
or U41639 (N_41639,N_38828,N_38703);
and U41640 (N_41640,N_38816,N_38462);
or U41641 (N_41641,N_39541,N_39474);
or U41642 (N_41642,N_37479,N_39852);
xor U41643 (N_41643,N_39197,N_38353);
xor U41644 (N_41644,N_37496,N_38070);
or U41645 (N_41645,N_38969,N_38383);
nand U41646 (N_41646,N_39351,N_37276);
and U41647 (N_41647,N_39636,N_37163);
or U41648 (N_41648,N_39381,N_38148);
nor U41649 (N_41649,N_39516,N_38575);
or U41650 (N_41650,N_38859,N_38642);
xor U41651 (N_41651,N_38805,N_39996);
nor U41652 (N_41652,N_35920,N_35652);
or U41653 (N_41653,N_35073,N_37417);
nand U41654 (N_41654,N_35092,N_39453);
nand U41655 (N_41655,N_37737,N_35687);
or U41656 (N_41656,N_39037,N_35401);
nand U41657 (N_41657,N_38962,N_38523);
nor U41658 (N_41658,N_35412,N_38705);
nor U41659 (N_41659,N_36349,N_35469);
nand U41660 (N_41660,N_36792,N_37486);
xnor U41661 (N_41661,N_38452,N_37553);
or U41662 (N_41662,N_39398,N_39383);
or U41663 (N_41663,N_35683,N_39390);
xnor U41664 (N_41664,N_37569,N_35318);
nand U41665 (N_41665,N_37466,N_38881);
nor U41666 (N_41666,N_39095,N_36631);
and U41667 (N_41667,N_36076,N_35694);
nand U41668 (N_41668,N_38890,N_36639);
or U41669 (N_41669,N_38692,N_37594);
nor U41670 (N_41670,N_38143,N_38001);
nor U41671 (N_41671,N_38448,N_37634);
xor U41672 (N_41672,N_36847,N_38049);
nand U41673 (N_41673,N_38336,N_35735);
nor U41674 (N_41674,N_37408,N_35237);
nand U41675 (N_41675,N_38620,N_38099);
xor U41676 (N_41676,N_37689,N_39187);
nor U41677 (N_41677,N_38929,N_37283);
or U41678 (N_41678,N_37230,N_37956);
or U41679 (N_41679,N_36653,N_38612);
and U41680 (N_41680,N_39506,N_36938);
nor U41681 (N_41681,N_36496,N_39067);
xor U41682 (N_41682,N_35028,N_39304);
nand U41683 (N_41683,N_38515,N_39743);
xor U41684 (N_41684,N_36429,N_39899);
nor U41685 (N_41685,N_35032,N_36517);
nand U41686 (N_41686,N_35859,N_35575);
nor U41687 (N_41687,N_39576,N_36913);
nand U41688 (N_41688,N_38835,N_38354);
and U41689 (N_41689,N_37379,N_38043);
nand U41690 (N_41690,N_35666,N_37168);
xor U41691 (N_41691,N_38155,N_35626);
and U41692 (N_41692,N_37521,N_35926);
or U41693 (N_41693,N_37176,N_37638);
nand U41694 (N_41694,N_39416,N_39179);
nor U41695 (N_41695,N_36440,N_36322);
or U41696 (N_41696,N_35847,N_38109);
nand U41697 (N_41697,N_38536,N_38667);
and U41698 (N_41698,N_37842,N_35504);
or U41699 (N_41699,N_36749,N_38839);
or U41700 (N_41700,N_36067,N_35010);
and U41701 (N_41701,N_35968,N_37809);
nor U41702 (N_41702,N_38777,N_35663);
nand U41703 (N_41703,N_38455,N_35817);
nor U41704 (N_41704,N_35289,N_36098);
or U41705 (N_41705,N_37369,N_39736);
or U41706 (N_41706,N_36842,N_38484);
and U41707 (N_41707,N_37256,N_36310);
nor U41708 (N_41708,N_36153,N_35701);
or U41709 (N_41709,N_39946,N_37471);
nor U41710 (N_41710,N_38919,N_39024);
and U41711 (N_41711,N_37896,N_38833);
nand U41712 (N_41712,N_38367,N_35753);
nor U41713 (N_41713,N_37714,N_38195);
nand U41714 (N_41714,N_37205,N_39808);
or U41715 (N_41715,N_36394,N_38659);
or U41716 (N_41716,N_39531,N_37790);
nor U41717 (N_41717,N_39847,N_36736);
nand U41718 (N_41718,N_39926,N_36754);
xnor U41719 (N_41719,N_35154,N_39707);
nor U41720 (N_41720,N_38079,N_38976);
nor U41721 (N_41721,N_35133,N_38783);
or U41722 (N_41722,N_39758,N_37024);
nor U41723 (N_41723,N_36620,N_36490);
or U41724 (N_41724,N_38577,N_36555);
and U41725 (N_41725,N_35729,N_39622);
xnor U41726 (N_41726,N_36009,N_35039);
xnor U41727 (N_41727,N_38534,N_35643);
nor U41728 (N_41728,N_36308,N_39395);
xor U41729 (N_41729,N_37879,N_35761);
nand U41730 (N_41730,N_36079,N_37155);
nor U41731 (N_41731,N_37086,N_37783);
nor U41732 (N_41732,N_35645,N_38986);
xnor U41733 (N_41733,N_38067,N_38809);
nor U41734 (N_41734,N_36529,N_36494);
or U41735 (N_41735,N_38698,N_37528);
nor U41736 (N_41736,N_37697,N_36566);
and U41737 (N_41737,N_37075,N_36521);
nor U41738 (N_41738,N_38438,N_36779);
or U41739 (N_41739,N_37606,N_36923);
nand U41740 (N_41740,N_39419,N_37352);
or U41741 (N_41741,N_39015,N_39128);
and U41742 (N_41742,N_38113,N_39048);
xnor U41743 (N_41743,N_39174,N_39397);
or U41744 (N_41744,N_39307,N_38637);
and U41745 (N_41745,N_39450,N_39925);
or U41746 (N_41746,N_39587,N_38421);
xnor U41747 (N_41747,N_38054,N_35653);
nor U41748 (N_41748,N_35231,N_39106);
nor U41749 (N_41749,N_37302,N_38347);
nand U41750 (N_41750,N_36480,N_38867);
nor U41751 (N_41751,N_38206,N_38162);
or U41752 (N_41752,N_37012,N_39336);
and U41753 (N_41753,N_35671,N_38665);
xnor U41754 (N_41754,N_35680,N_38031);
or U41755 (N_41755,N_38758,N_36011);
and U41756 (N_41756,N_37512,N_36748);
or U41757 (N_41757,N_37785,N_39500);
nor U41758 (N_41758,N_37169,N_36688);
or U41759 (N_41759,N_37186,N_39031);
or U41760 (N_41760,N_37880,N_35148);
xor U41761 (N_41761,N_39434,N_36852);
nand U41762 (N_41762,N_38757,N_37609);
nor U41763 (N_41763,N_39038,N_37351);
and U41764 (N_41764,N_35036,N_36420);
xor U41765 (N_41765,N_38052,N_36692);
nor U41766 (N_41766,N_35236,N_39284);
nand U41767 (N_41767,N_37749,N_37085);
or U41768 (N_41768,N_36624,N_38450);
nor U41769 (N_41769,N_39949,N_35470);
xor U41770 (N_41770,N_35348,N_39392);
xnor U41771 (N_41771,N_39549,N_35262);
nand U41772 (N_41772,N_38576,N_35499);
xnor U41773 (N_41773,N_39418,N_38765);
and U41774 (N_41774,N_39970,N_38398);
nand U41775 (N_41775,N_36266,N_39805);
nand U41776 (N_41776,N_35107,N_38806);
or U41777 (N_41777,N_38850,N_36121);
or U41778 (N_41778,N_37492,N_39694);
or U41779 (N_41779,N_36743,N_38735);
and U41780 (N_41780,N_37866,N_37675);
and U41781 (N_41781,N_36246,N_38272);
nand U41782 (N_41782,N_38681,N_35988);
nor U41783 (N_41783,N_38887,N_35163);
xnor U41784 (N_41784,N_36906,N_38332);
nand U41785 (N_41785,N_38611,N_37798);
xnor U41786 (N_41786,N_39747,N_35796);
and U41787 (N_41787,N_38601,N_38788);
nand U41788 (N_41788,N_35392,N_38684);
nor U41789 (N_41789,N_36665,N_35932);
or U41790 (N_41790,N_39238,N_37877);
nand U41791 (N_41791,N_36022,N_35489);
nand U41792 (N_41792,N_35281,N_39890);
and U41793 (N_41793,N_37304,N_37700);
xor U41794 (N_41794,N_39749,N_37965);
nand U41795 (N_41795,N_38237,N_35987);
and U41796 (N_41796,N_38663,N_39756);
or U41797 (N_41797,N_39643,N_38410);
or U41798 (N_41798,N_37378,N_38669);
and U41799 (N_41799,N_37686,N_36965);
nor U41800 (N_41800,N_39538,N_38950);
nor U41801 (N_41801,N_37487,N_37875);
xnor U41802 (N_41802,N_37955,N_37215);
or U41803 (N_41803,N_39140,N_37536);
nor U41804 (N_41804,N_38790,N_38537);
and U41805 (N_41805,N_38405,N_36823);
xor U41806 (N_41806,N_36483,N_36018);
nand U41807 (N_41807,N_38690,N_36914);
and U41808 (N_41808,N_35904,N_39348);
or U41809 (N_41809,N_39356,N_35918);
nand U41810 (N_41810,N_39781,N_38908);
xnor U41811 (N_41811,N_38239,N_35106);
or U41812 (N_41812,N_38172,N_39188);
nor U41813 (N_41813,N_35313,N_39671);
or U41814 (N_41814,N_38741,N_35144);
nor U41815 (N_41815,N_35384,N_39005);
and U41816 (N_41816,N_39583,N_37289);
nor U41817 (N_41817,N_39218,N_37005);
xor U41818 (N_41818,N_39963,N_36345);
xor U41819 (N_41819,N_39662,N_38913);
nand U41820 (N_41820,N_36388,N_35093);
xor U41821 (N_41821,N_37912,N_35522);
or U41822 (N_41822,N_35711,N_35349);
nor U41823 (N_41823,N_35090,N_37600);
or U41824 (N_41824,N_35646,N_36961);
and U41825 (N_41825,N_39515,N_36241);
or U41826 (N_41826,N_39829,N_39467);
xor U41827 (N_41827,N_37428,N_36487);
nand U41828 (N_41828,N_35175,N_37011);
xnor U41829 (N_41829,N_36588,N_35284);
nand U41830 (N_41830,N_35929,N_38418);
xnor U41831 (N_41831,N_37104,N_37006);
and U41832 (N_41832,N_38038,N_38865);
or U41833 (N_41833,N_39575,N_35984);
or U41834 (N_41834,N_39936,N_36360);
or U41835 (N_41835,N_38081,N_35952);
nor U41836 (N_41836,N_37453,N_38164);
or U41837 (N_41837,N_38181,N_37207);
or U41838 (N_41838,N_38953,N_39083);
or U41839 (N_41839,N_37604,N_37004);
or U41840 (N_41840,N_36739,N_38121);
and U41841 (N_41841,N_36058,N_38888);
nor U41842 (N_41842,N_35670,N_35127);
and U41843 (N_41843,N_37052,N_35013);
xnor U41844 (N_41844,N_36897,N_36831);
nand U41845 (N_41845,N_37658,N_39705);
nor U41846 (N_41846,N_39078,N_37361);
and U41847 (N_41847,N_37235,N_36183);
or U41848 (N_41848,N_38891,N_37957);
nand U41849 (N_41849,N_37126,N_35302);
nand U41850 (N_41850,N_35150,N_36284);
nand U41851 (N_41851,N_39977,N_39731);
nand U41852 (N_41852,N_39885,N_36367);
nor U41853 (N_41853,N_35751,N_39232);
xnor U41854 (N_41854,N_36344,N_37384);
and U41855 (N_41855,N_35637,N_37425);
and U41856 (N_41856,N_35353,N_39975);
and U41857 (N_41857,N_37160,N_39518);
xor U41858 (N_41858,N_38120,N_38396);
nor U41859 (N_41859,N_36678,N_36948);
nand U41860 (N_41860,N_39943,N_35982);
or U41861 (N_41861,N_35730,N_38564);
nand U41862 (N_41862,N_36267,N_36236);
or U41863 (N_41863,N_37091,N_37305);
xnor U41864 (N_41864,N_36428,N_38938);
and U41865 (N_41865,N_38578,N_36321);
nor U41866 (N_41866,N_38974,N_38339);
and U41867 (N_41867,N_38165,N_39469);
nor U41868 (N_41868,N_38943,N_38721);
xnor U41869 (N_41869,N_38832,N_39835);
nand U41870 (N_41870,N_39413,N_35202);
nor U41871 (N_41871,N_35498,N_39352);
and U41872 (N_41872,N_36622,N_35453);
nor U41873 (N_41873,N_37401,N_37073);
and U41874 (N_41874,N_35569,N_35468);
nand U41875 (N_41875,N_39152,N_39966);
nand U41876 (N_41876,N_35986,N_35866);
xor U41877 (N_41877,N_38442,N_36055);
or U41878 (N_41878,N_39544,N_36384);
xnor U41879 (N_41879,N_35619,N_39593);
and U41880 (N_41880,N_37449,N_39773);
or U41881 (N_41881,N_35129,N_39116);
xor U41882 (N_41882,N_36627,N_36130);
xor U41883 (N_41883,N_36579,N_36903);
nor U41884 (N_41884,N_36518,N_35974);
nor U41885 (N_41885,N_35697,N_39222);
nor U41886 (N_41886,N_36527,N_38188);
and U41887 (N_41887,N_39455,N_35263);
or U41888 (N_41888,N_37270,N_35151);
and U41889 (N_41889,N_38158,N_38321);
or U41890 (N_41890,N_38041,N_36471);
or U41891 (N_41891,N_38417,N_38640);
and U41892 (N_41892,N_35278,N_39958);
xnor U41893 (N_41893,N_35597,N_38391);
or U41894 (N_41894,N_38514,N_36731);
nand U41895 (N_41895,N_36091,N_39706);
or U41896 (N_41896,N_37690,N_37685);
and U41897 (N_41897,N_35835,N_37380);
nand U41898 (N_41898,N_39729,N_36207);
or U41899 (N_41899,N_36761,N_36049);
and U41900 (N_41900,N_39205,N_36538);
or U41901 (N_41901,N_35102,N_38497);
xor U41902 (N_41902,N_36348,N_35890);
nor U41903 (N_41903,N_37273,N_37264);
or U41904 (N_41904,N_39828,N_39625);
and U41905 (N_41905,N_37819,N_35406);
nor U41906 (N_41906,N_37159,N_36202);
xor U41907 (N_41907,N_35420,N_36516);
nor U41908 (N_41908,N_37555,N_35351);
nand U41909 (N_41909,N_36326,N_37848);
nor U41910 (N_41910,N_37614,N_37387);
and U41911 (N_41911,N_37831,N_35011);
nand U41912 (N_41912,N_35815,N_36833);
nor U41913 (N_41913,N_35991,N_36983);
nor U41914 (N_41914,N_38108,N_35495);
xnor U41915 (N_41915,N_36239,N_38265);
nand U41916 (N_41916,N_39333,N_39071);
xnor U41917 (N_41917,N_37335,N_36298);
nand U41918 (N_41918,N_39201,N_37818);
xnor U41919 (N_41919,N_36324,N_37936);
and U41920 (N_41920,N_35275,N_39460);
xnor U41921 (N_41921,N_37760,N_36103);
xnor U41922 (N_41922,N_35798,N_35702);
and U41923 (N_41923,N_38847,N_35306);
or U41924 (N_41924,N_36830,N_36751);
nand U41925 (N_41925,N_36893,N_39658);
or U41926 (N_41926,N_38241,N_39669);
xor U41927 (N_41927,N_39770,N_35669);
nand U41928 (N_41928,N_35642,N_39161);
nor U41929 (N_41929,N_36505,N_35756);
and U41930 (N_41930,N_39314,N_36105);
nor U41931 (N_41931,N_37277,N_36872);
and U41932 (N_41932,N_35863,N_35344);
and U41933 (N_41933,N_37366,N_35607);
nand U41934 (N_41934,N_39442,N_39889);
xor U41935 (N_41935,N_36441,N_36911);
nor U41936 (N_41936,N_36477,N_37673);
or U41937 (N_41937,N_37601,N_35250);
nor U41938 (N_41938,N_36958,N_39497);
nor U41939 (N_41939,N_35024,N_38598);
xor U41940 (N_41940,N_38119,N_38501);
or U41941 (N_41941,N_35188,N_39668);
or U41942 (N_41942,N_38571,N_35902);
and U41943 (N_41943,N_38341,N_36472);
nand U41944 (N_41944,N_39627,N_37072);
or U41945 (N_41945,N_36446,N_36261);
xor U41946 (N_41946,N_38145,N_35947);
or U41947 (N_41947,N_39921,N_37092);
nor U41948 (N_41948,N_38775,N_39753);
and U41949 (N_41949,N_39320,N_37757);
nand U41950 (N_41950,N_38009,N_38491);
nor U41951 (N_41951,N_35814,N_36060);
xor U41952 (N_41952,N_35807,N_39347);
xor U41953 (N_41953,N_37132,N_39993);
nand U41954 (N_41954,N_35639,N_36871);
nor U41955 (N_41955,N_37633,N_37423);
nor U41956 (N_41956,N_37782,N_37396);
xor U41957 (N_41957,N_36149,N_35985);
or U41958 (N_41958,N_35402,N_38389);
or U41959 (N_41959,N_38399,N_37146);
nor U41960 (N_41960,N_35681,N_36219);
nand U41961 (N_41961,N_37399,N_36418);
xnor U41962 (N_41962,N_35900,N_39700);
nor U41963 (N_41963,N_36667,N_39969);
nor U41964 (N_41964,N_36275,N_35176);
or U41965 (N_41965,N_35052,N_38198);
and U41966 (N_41966,N_38479,N_35765);
and U41967 (N_41967,N_36623,N_38654);
and U41968 (N_41968,N_35979,N_38556);
xnor U41969 (N_41969,N_36960,N_39235);
xnor U41970 (N_41970,N_37670,N_38971);
and U41971 (N_41971,N_36548,N_35119);
nand U41972 (N_41972,N_39523,N_37152);
nor U41973 (N_41973,N_35895,N_38302);
xor U41974 (N_41974,N_36512,N_35743);
and U41975 (N_41975,N_38371,N_36116);
or U41976 (N_41976,N_37641,N_36101);
or U41977 (N_41977,N_36426,N_37116);
nand U41978 (N_41978,N_39646,N_39745);
and U41979 (N_41979,N_36111,N_38175);
xor U41980 (N_41980,N_39717,N_37294);
and U41981 (N_41981,N_36507,N_36448);
nor U41982 (N_41982,N_39125,N_38212);
nor U41983 (N_41983,N_37200,N_38269);
nor U41984 (N_41984,N_36796,N_39461);
or U41985 (N_41985,N_35995,N_39375);
or U41986 (N_41986,N_36502,N_37629);
xor U41987 (N_41987,N_39076,N_39528);
and U41988 (N_41988,N_35841,N_39769);
nor U41989 (N_41989,N_35545,N_37953);
nor U41990 (N_41990,N_38483,N_39445);
xor U41991 (N_41991,N_37221,N_38355);
xnor U41992 (N_41992,N_39065,N_39502);
and U41993 (N_41993,N_39221,N_39709);
xnor U41994 (N_41994,N_35448,N_35629);
and U41995 (N_41995,N_38309,N_37824);
xor U41996 (N_41996,N_39051,N_36704);
xnor U41997 (N_41997,N_36910,N_36686);
xor U41998 (N_41998,N_37054,N_39231);
xor U41999 (N_41999,N_39931,N_37403);
and U42000 (N_42000,N_37803,N_36297);
and U42001 (N_42001,N_35343,N_38171);
nor U42002 (N_42002,N_38985,N_36046);
and U42003 (N_42003,N_38588,N_36995);
and U42004 (N_42004,N_39973,N_39976);
xor U42005 (N_42005,N_37016,N_35476);
nor U42006 (N_42006,N_36402,N_35588);
nor U42007 (N_42007,N_35783,N_35101);
and U42008 (N_42008,N_36328,N_37653);
or U42009 (N_42009,N_39465,N_36757);
xor U42010 (N_42010,N_37105,N_36305);
nand U42011 (N_42011,N_35725,N_37582);
nand U42012 (N_42012,N_35845,N_35851);
or U42013 (N_42013,N_35566,N_39021);
nor U42014 (N_42014,N_35280,N_37427);
nor U42015 (N_42015,N_36064,N_35362);
nand U42016 (N_42016,N_35437,N_39055);
xor U42017 (N_42017,N_38956,N_35183);
nor U42018 (N_42018,N_39028,N_37703);
and U42019 (N_42019,N_36218,N_35723);
nor U42020 (N_42020,N_37254,N_36342);
xnor U42021 (N_42021,N_37278,N_35187);
nand U42022 (N_42022,N_35082,N_36285);
or U42023 (N_42023,N_39016,N_37742);
xor U42024 (N_42024,N_38139,N_36676);
nor U42025 (N_42025,N_38594,N_36444);
nor U42026 (N_42026,N_38622,N_36783);
and U42027 (N_42027,N_37728,N_38967);
nor U42028 (N_42028,N_39407,N_36973);
nor U42029 (N_42029,N_36280,N_37415);
or U42030 (N_42030,N_36840,N_39603);
xnor U42031 (N_42031,N_35209,N_35881);
nor U42032 (N_42032,N_38191,N_39876);
or U42033 (N_42033,N_39546,N_39964);
nand U42034 (N_42034,N_37046,N_35641);
xnor U42035 (N_42035,N_37982,N_37586);
and U42036 (N_42036,N_38821,N_39813);
xnor U42037 (N_42037,N_39644,N_37309);
nor U42038 (N_42038,N_36674,N_36696);
nor U42039 (N_42039,N_36140,N_36048);
or U42040 (N_42040,N_39156,N_36987);
xor U42041 (N_42041,N_38085,N_37214);
nand U42042 (N_42042,N_39027,N_37222);
nor U42043 (N_42043,N_39667,N_38156);
nor U42044 (N_42044,N_37707,N_36920);
or U42045 (N_42045,N_39844,N_35770);
and U42046 (N_42046,N_38225,N_37998);
nor U42047 (N_42047,N_35534,N_38213);
and U42048 (N_42048,N_39824,N_36780);
and U42049 (N_42049,N_36744,N_37137);
xnor U42050 (N_42050,N_37940,N_38183);
xor U42051 (N_42051,N_39122,N_35665);
or U42052 (N_42052,N_35265,N_36741);
xnor U42053 (N_42053,N_37071,N_37756);
nand U42054 (N_42054,N_37966,N_36849);
or U42055 (N_42055,N_37610,N_36907);
and U42056 (N_42056,N_36422,N_35517);
or U42057 (N_42057,N_36569,N_38474);
and U42058 (N_42058,N_36157,N_37339);
and U42059 (N_42059,N_35625,N_36172);
xor U42060 (N_42060,N_35058,N_36541);
and U42061 (N_42061,N_35674,N_36563);
nor U42062 (N_42062,N_38940,N_36621);
xnor U42063 (N_42063,N_36212,N_37514);
nand U42064 (N_42064,N_39539,N_39421);
and U42065 (N_42065,N_39737,N_36093);
nand U42066 (N_42066,N_36592,N_38002);
xnor U42067 (N_42067,N_37951,N_37404);
or U42068 (N_42068,N_35428,N_39934);
or U42069 (N_42069,N_35261,N_35452);
nor U42070 (N_42070,N_36706,N_38717);
and U42071 (N_42071,N_39332,N_38433);
nor U42072 (N_42072,N_39630,N_37250);
and U42073 (N_42073,N_36523,N_37625);
and U42074 (N_42074,N_36351,N_38572);
nor U42075 (N_42075,N_35950,N_36788);
nand U42076 (N_42076,N_35518,N_36025);
nor U42077 (N_42077,N_37915,N_39655);
nor U42078 (N_42078,N_39884,N_38327);
nor U42079 (N_42079,N_39988,N_35612);
nor U42080 (N_42080,N_35439,N_38568);
or U42081 (N_42081,N_37713,N_35523);
nand U42082 (N_42082,N_37793,N_36200);
nor U42083 (N_42083,N_39130,N_35822);
or U42084 (N_42084,N_39823,N_36721);
nand U42085 (N_42085,N_36164,N_36657);
xnor U42086 (N_42086,N_35255,N_35259);
xnor U42087 (N_42087,N_38439,N_37846);
nand U42088 (N_42088,N_37253,N_35821);
xnor U42089 (N_42089,N_39213,N_36942);
or U42090 (N_42090,N_38592,N_36407);
nand U42091 (N_42091,N_39291,N_37840);
xor U42092 (N_42092,N_38794,N_38613);
xor U42093 (N_42093,N_39151,N_37131);
xnor U42094 (N_42094,N_36719,N_37914);
nor U42095 (N_42095,N_35374,N_36380);
and U42096 (N_42096,N_37288,N_38672);
and U42097 (N_42097,N_37244,N_38607);
or U42098 (N_42098,N_37381,N_35444);
and U42099 (N_42099,N_35317,N_37917);
nand U42100 (N_42100,N_35301,N_38407);
xnor U42101 (N_42101,N_36769,N_36002);
xor U42102 (N_42102,N_36217,N_36432);
and U42103 (N_42103,N_36364,N_38475);
nand U42104 (N_42104,N_39306,N_36604);
nor U42105 (N_42105,N_37444,N_36168);
nor U42106 (N_42106,N_39599,N_35672);
nand U42107 (N_42107,N_38179,N_39117);
xnor U42108 (N_42108,N_35164,N_35998);
nor U42109 (N_42109,N_37098,N_37079);
xnor U42110 (N_42110,N_36254,N_38778);
nor U42111 (N_42111,N_37616,N_37771);
xnor U42112 (N_42112,N_38374,N_39211);
or U42113 (N_42113,N_35243,N_36438);
and U42114 (N_42114,N_37677,N_38876);
nor U42115 (N_42115,N_39388,N_36762);
nand U42116 (N_42116,N_39637,N_36353);
xor U42117 (N_42117,N_36043,N_35463);
nand U42118 (N_42118,N_37431,N_36199);
xnor U42119 (N_42119,N_39634,N_36717);
or U42120 (N_42120,N_38493,N_36927);
nand U42121 (N_42121,N_37491,N_36976);
nor U42122 (N_42122,N_39456,N_36318);
or U42123 (N_42123,N_36606,N_37709);
nand U42124 (N_42124,N_36999,N_35631);
and U42125 (N_42125,N_38507,N_37666);
xnor U42126 (N_42126,N_35691,N_35638);
nand U42127 (N_42127,N_35907,N_38552);
or U42128 (N_42128,N_37391,N_37751);
nand U42129 (N_42129,N_38451,N_36918);
nor U42130 (N_42130,N_35509,N_38133);
nand U42131 (N_42131,N_38262,N_38301);
and U42132 (N_42132,N_36984,N_39458);
nor U42133 (N_42133,N_38551,N_36113);
nand U42134 (N_42134,N_36856,N_36119);
and U42135 (N_42135,N_37183,N_36720);
and U42136 (N_42136,N_37460,N_39537);
or U42137 (N_42137,N_39033,N_37133);
or U42138 (N_42138,N_35061,N_37296);
or U42139 (N_42139,N_37003,N_36880);
and U42140 (N_42140,N_36463,N_37712);
nor U42141 (N_42141,N_35212,N_37627);
xnor U42142 (N_42142,N_36878,N_36354);
or U42143 (N_42143,N_36634,N_39386);
nand U42144 (N_42144,N_35291,N_35716);
and U42145 (N_42145,N_39999,N_37187);
nand U42146 (N_42146,N_35598,N_38403);
nand U42147 (N_42147,N_38630,N_35959);
nor U42148 (N_42148,N_38595,N_35232);
and U42149 (N_42149,N_36877,N_36026);
and U42150 (N_42150,N_37938,N_39957);
nor U42151 (N_42151,N_38759,N_39724);
nor U42152 (N_42152,N_36964,N_37203);
nor U42153 (N_42153,N_38488,N_39696);
nand U42154 (N_42154,N_36511,N_39720);
xor U42155 (N_42155,N_35342,N_37412);
or U42156 (N_42156,N_37267,N_37989);
nor U42157 (N_42157,N_39062,N_35427);
nor U42158 (N_42158,N_37642,N_35613);
and U42159 (N_42159,N_36145,N_38980);
and U42160 (N_42160,N_38047,N_39412);
nor U42161 (N_42161,N_36683,N_37801);
or U42162 (N_42162,N_38936,N_37020);
nor U42163 (N_42163,N_36336,N_39803);
xor U42164 (N_42164,N_35726,N_36307);
or U42165 (N_42165,N_37096,N_39020);
nand U42166 (N_42166,N_35868,N_39244);
and U42167 (N_42167,N_35395,N_39160);
and U42168 (N_42168,N_37974,N_35197);
nand U42169 (N_42169,N_37143,N_35812);
or U42170 (N_42170,N_36546,N_39355);
xor U42171 (N_42171,N_38340,N_37260);
xor U42172 (N_42172,N_39938,N_36728);
nand U42173 (N_42173,N_36016,N_39623);
or U42174 (N_42174,N_37970,N_37946);
nand U42175 (N_42175,N_37280,N_37899);
nand U42176 (N_42176,N_39494,N_37285);
nand U42177 (N_42177,N_35012,N_39917);
or U42178 (N_42178,N_38215,N_37581);
nor U42179 (N_42179,N_35682,N_35316);
xnor U42180 (N_42180,N_35657,N_38780);
or U42181 (N_42181,N_36648,N_35299);
nor U42182 (N_42182,N_38589,N_37007);
nand U42183 (N_42183,N_38390,N_38256);
nand U42184 (N_42184,N_38840,N_36263);
and U42185 (N_42185,N_38495,N_39414);
nand U42186 (N_42186,N_39992,N_39092);
or U42187 (N_42187,N_39448,N_35016);
nor U42188 (N_42188,N_39738,N_37777);
or U42189 (N_42189,N_36528,N_37662);
nor U42190 (N_42190,N_38670,N_35276);
or U42191 (N_42191,N_35919,N_36042);
nand U42192 (N_42192,N_35268,N_36758);
nor U42193 (N_42193,N_35328,N_39359);
xor U42194 (N_42194,N_37718,N_39678);
and U42195 (N_42195,N_39118,N_38791);
and U42196 (N_42196,N_35435,N_36397);
xor U42197 (N_42197,N_37127,N_37049);
and U42198 (N_42198,N_38770,N_39155);
nor U42199 (N_42199,N_36357,N_37510);
nand U42200 (N_42200,N_39800,N_38895);
nand U42201 (N_42201,N_35041,N_39915);
and U42202 (N_42202,N_36379,N_38142);
or U42203 (N_42203,N_36481,N_36584);
or U42204 (N_42204,N_38346,N_37805);
nor U42205 (N_42205,N_37043,N_39266);
or U42206 (N_42206,N_37248,N_37506);
nand U42207 (N_42207,N_37655,N_37574);
nor U42208 (N_42208,N_37010,N_39836);
nand U42209 (N_42209,N_36514,N_38988);
nand U42210 (N_42210,N_39217,N_38762);
xor U42211 (N_42211,N_36867,N_38299);
nor U42212 (N_42212,N_35550,N_39478);
nor U42213 (N_42213,N_36330,N_39239);
nand U42214 (N_42214,N_39137,N_36459);
xor U42215 (N_42215,N_38784,N_37499);
and U42216 (N_42216,N_36603,N_36245);
and U42217 (N_42217,N_35689,N_38739);
or U42218 (N_42218,N_39452,N_38871);
nand U42219 (N_42219,N_36737,N_38570);
or U42220 (N_42220,N_37567,N_39735);
nand U42221 (N_42221,N_37322,N_35844);
or U42222 (N_42222,N_35105,N_38292);
and U42223 (N_42223,N_37031,N_37806);
nand U42224 (N_42224,N_39692,N_35460);
xor U42225 (N_42225,N_38275,N_39606);
nor U42226 (N_42226,N_38691,N_38003);
nor U42227 (N_42227,N_35193,N_37350);
nor U42228 (N_42228,N_37300,N_37800);
and U42229 (N_42229,N_38457,N_37885);
xor U42230 (N_42230,N_37827,N_36056);
and U42231 (N_42231,N_39454,N_36363);
xnor U42232 (N_42232,N_36649,N_36797);
nor U42233 (N_42233,N_36289,N_35064);
nand U42234 (N_42234,N_37128,N_38028);
nor U42235 (N_42235,N_39689,N_38533);
and U42236 (N_42236,N_37174,N_37201);
nor U42237 (N_42237,N_38228,N_35218);
nor U42238 (N_42238,N_35823,N_35177);
and U42239 (N_42239,N_38040,N_39788);
or U42240 (N_42240,N_38520,N_36096);
nand U42241 (N_42241,N_36369,N_36405);
nor U42242 (N_42242,N_38661,N_38004);
or U42243 (N_42243,N_39503,N_35411);
nand U42244 (N_42244,N_36845,N_36735);
nor U42245 (N_42245,N_35382,N_38153);
and U42246 (N_42246,N_36087,N_35408);
xnor U42247 (N_42247,N_37372,N_38704);
nor U42248 (N_42248,N_36506,N_36635);
and U42249 (N_42249,N_38306,N_37458);
xor U42250 (N_42250,N_37242,N_35944);
nor U42251 (N_42251,N_35322,N_39635);
or U42252 (N_42252,N_38035,N_36156);
xor U42253 (N_42253,N_36612,N_37101);
and U42254 (N_42254,N_39264,N_39251);
and U42255 (N_42255,N_39163,N_38334);
and U42256 (N_42256,N_35391,N_38202);
xor U42257 (N_42257,N_35786,N_35290);
nor U42258 (N_42258,N_39451,N_36875);
and U42259 (N_42259,N_35124,N_38603);
and U42260 (N_42260,N_39892,N_38184);
nand U42261 (N_42261,N_38423,N_38350);
or U42262 (N_42262,N_39343,N_39777);
or U42263 (N_42263,N_36054,N_39142);
xnor U42264 (N_42264,N_37659,N_37721);
or U42265 (N_42265,N_35693,N_39730);
nand U42266 (N_42266,N_37249,N_36059);
nor U42267 (N_42267,N_35189,N_35370);
nor U42268 (N_42268,N_35806,N_39368);
nor U42269 (N_42269,N_36941,N_39185);
or U42270 (N_42270,N_35869,N_36393);
nand U42271 (N_42271,N_36979,N_37860);
nand U42272 (N_42272,N_39819,N_37363);
or U42273 (N_42273,N_37523,N_37418);
nor U42274 (N_42274,N_35526,N_38699);
xor U42275 (N_42275,N_37314,N_36957);
or U42276 (N_42276,N_39566,N_38958);
nand U42277 (N_42277,N_38279,N_39818);
and U42278 (N_42278,N_36695,N_35403);
nand U42279 (N_42279,N_37871,N_39766);
nor U42280 (N_42280,N_39050,N_39119);
or U42281 (N_42281,N_36750,N_39358);
nor U42282 (N_42282,N_38921,N_37081);
or U42283 (N_42283,N_37074,N_37346);
xor U42284 (N_42284,N_35477,N_39760);
nor U42285 (N_42285,N_35994,N_39405);
and U42286 (N_42286,N_35848,N_36594);
and U42287 (N_42287,N_38843,N_39680);
and U42288 (N_42288,N_39868,N_37266);
or U42289 (N_42289,N_39376,N_36811);
nor U42290 (N_42290,N_38361,N_35999);
nand U42291 (N_42291,N_39989,N_36498);
nand U42292 (N_42292,N_39612,N_38203);
nand U42293 (N_42293,N_38498,N_38251);
and U42294 (N_42294,N_37835,N_37887);
and U42295 (N_42295,N_37566,N_35046);
nor U42296 (N_42296,N_36014,N_39504);
and U42297 (N_42297,N_39734,N_35514);
nor U42298 (N_42298,N_39935,N_35419);
or U42299 (N_42299,N_39484,N_39486);
or U42300 (N_42300,N_39132,N_35971);
nand U42301 (N_42301,N_38529,N_38420);
xor U42302 (N_42302,N_36019,N_38912);
xnor U42303 (N_42303,N_37231,N_36155);
nand U42304 (N_42304,N_37841,N_39323);
xor U42305 (N_42305,N_39255,N_38042);
or U42306 (N_42306,N_38619,N_38381);
or U42307 (N_42307,N_35939,N_39875);
and U42308 (N_42308,N_38094,N_35557);
xor U42309 (N_42309,N_37032,N_39952);
xnor U42310 (N_42310,N_37537,N_35447);
or U42311 (N_42311,N_35407,N_35728);
nand U42312 (N_42312,N_36387,N_39754);
xor U42313 (N_42313,N_38586,N_38525);
and U42314 (N_42314,N_35794,N_38200);
or U42315 (N_42315,N_35319,N_39924);
xor U42316 (N_42316,N_35502,N_37420);
or U42317 (N_42317,N_38197,N_36176);
nor U42318 (N_42318,N_35599,N_36861);
nor U42319 (N_42319,N_39867,N_37844);
nand U42320 (N_42320,N_35967,N_39880);
xor U42321 (N_42321,N_37247,N_36474);
and U42322 (N_42322,N_36959,N_35213);
nor U42323 (N_42323,N_39334,N_35140);
xor U42324 (N_42324,N_39350,N_37103);
nor U42325 (N_42325,N_35699,N_38952);
or U42326 (N_42326,N_37868,N_38244);
nand U42327 (N_42327,N_39428,N_38258);
nor U42328 (N_42328,N_38271,N_38610);
xnor U42329 (N_42329,N_39792,N_35321);
xnor U42330 (N_42330,N_36777,N_38634);
nor U42331 (N_42331,N_37704,N_39335);
nor U42332 (N_42332,N_35207,N_35341);
nand U42333 (N_42333,N_35842,N_36452);
xnor U42334 (N_42334,N_38934,N_39326);
or U42335 (N_42335,N_37319,N_36691);
or U42336 (N_42336,N_39269,N_36437);
or U42337 (N_42337,N_38585,N_36770);
nand U42338 (N_42338,N_38546,N_39710);
xnor U42339 (N_42339,N_35917,N_39184);
or U42340 (N_42340,N_35459,N_37337);
xor U42341 (N_42341,N_35651,N_39220);
or U42342 (N_42342,N_37069,N_37632);
and U42343 (N_42343,N_35159,N_37355);
or U42344 (N_42344,N_38827,N_36235);
xnor U42345 (N_42345,N_36313,N_38342);
or U42346 (N_42346,N_37669,N_38745);
nor U42347 (N_42347,N_39905,N_38375);
or U42348 (N_42348,N_37904,N_39295);
xnor U42349 (N_42349,N_38178,N_35747);
nand U42350 (N_42350,N_36881,N_38521);
xnor U42351 (N_42351,N_38712,N_36117);
and U42352 (N_42352,N_35222,N_38994);
and U42353 (N_42353,N_39512,N_36699);
xnor U42354 (N_42354,N_39677,N_36536);
xor U42355 (N_42355,N_38176,N_38922);
and U42356 (N_42356,N_36197,N_38946);
and U42357 (N_42357,N_35431,N_37585);
xnor U42358 (N_42358,N_38062,N_36816);
nor U42359 (N_42359,N_35742,N_38565);
or U42360 (N_42360,N_39536,N_37382);
nand U42361 (N_42361,N_38458,N_38686);
nand U42362 (N_42362,N_37148,N_39093);
nand U42363 (N_42363,N_37135,N_38786);
and U42364 (N_42364,N_37389,N_37434);
nand U42365 (N_42365,N_39827,N_38059);
xnor U42366 (N_42366,N_37862,N_35533);
xnor U42367 (N_42367,N_36892,N_36542);
or U42368 (N_42368,N_36007,N_35473);
or U42369 (N_42369,N_35836,N_39401);
and U42370 (N_42370,N_39872,N_35303);
nand U42371 (N_42371,N_36598,N_38000);
or U42372 (N_42372,N_35861,N_39672);
or U42373 (N_42373,N_35219,N_38685);
nand U42374 (N_42374,N_36982,N_36801);
or U42375 (N_42375,N_39916,N_39373);
or U42376 (N_42376,N_38885,N_36109);
and U42377 (N_42377,N_36314,N_36435);
xnor U42378 (N_42378,N_36766,N_36462);
xnor U42379 (N_42379,N_39856,N_39496);
or U42380 (N_42380,N_37945,N_38566);
and U42381 (N_42381,N_37262,N_39389);
and U42382 (N_42382,N_35314,N_37087);
nand U42383 (N_42383,N_38785,N_35100);
or U42384 (N_42384,N_39006,N_35329);
nor U42385 (N_42385,N_37695,N_35785);
and U42386 (N_42386,N_38814,N_37484);
or U42387 (N_42387,N_36240,N_35698);
and U42388 (N_42388,N_36244,N_39176);
nand U42389 (N_42389,N_38854,N_35644);
nand U42390 (N_42390,N_36513,N_36185);
or U42391 (N_42391,N_37596,N_39058);
and U42392 (N_42392,N_39136,N_39954);
or U42393 (N_42393,N_35764,N_39338);
or U42394 (N_42394,N_38925,N_38173);
xor U42395 (N_42395,N_37576,N_37217);
nand U42396 (N_42396,N_38268,N_35134);
nand U42397 (N_42397,N_37051,N_37750);
and U42398 (N_42398,N_36711,N_38106);
and U42399 (N_42399,N_37978,N_35568);
or U42400 (N_42400,N_37823,N_37290);
nand U42401 (N_42401,N_39303,N_38763);
xnor U42402 (N_42402,N_39121,N_35608);
and U42403 (N_42403,N_37741,N_38308);
nor U42404 (N_42404,N_35029,N_38259);
nand U42405 (N_42405,N_38278,N_36133);
and U42406 (N_42406,N_35776,N_35294);
nand U42407 (N_42407,N_39653,N_36268);
or U42408 (N_42408,N_39096,N_38066);
nand U42409 (N_42409,N_39203,N_36633);
nand U42410 (N_42410,N_38107,N_37646);
or U42411 (N_42411,N_37619,N_36279);
xnor U42412 (N_42412,N_36100,N_39099);
or U42413 (N_42413,N_36929,N_36859);
nor U42414 (N_42414,N_36468,N_39228);
xnor U42415 (N_42415,N_39638,N_36937);
xor U42416 (N_42416,N_36813,N_36006);
nand U42417 (N_42417,N_37317,N_39305);
or U42418 (N_42418,N_38072,N_38087);
or U42419 (N_42419,N_38752,N_35347);
nand U42420 (N_42420,N_35655,N_38419);
xor U42421 (N_42421,N_35072,N_39862);
and U42422 (N_42422,N_38222,N_36848);
and U42423 (N_42423,N_36411,N_36147);
and U42424 (N_42424,N_35135,N_36873);
or U42425 (N_42425,N_37657,N_36382);
or U42426 (N_42426,N_36994,N_39147);
nor U42427 (N_42427,N_35547,N_35673);
or U42428 (N_42428,N_36609,N_36775);
xnor U42429 (N_42429,N_38316,N_35018);
nand U42430 (N_42430,N_35810,N_38406);
xnor U42431 (N_42431,N_38861,N_36366);
nand U42432 (N_42432,N_35251,N_35562);
or U42433 (N_42433,N_39493,N_37933);
or U42434 (N_42434,N_37701,N_37286);
or U42435 (N_42435,N_39133,N_35983);
xor U42436 (N_42436,N_39158,N_35854);
nor U42437 (N_42437,N_39084,N_37558);
xor U42438 (N_42438,N_38277,N_39898);
nor U42439 (N_42439,N_38779,N_35422);
nor U42440 (N_42440,N_35478,N_37136);
nor U42441 (N_42441,N_39511,N_37545);
nand U42442 (N_42442,N_36582,N_39919);
or U42443 (N_42443,N_35241,N_38216);
nor U42444 (N_42444,N_39795,N_37740);
or U42445 (N_42445,N_35483,N_38616);
xor U42446 (N_42446,N_35856,N_36675);
and U42447 (N_42447,N_36909,N_36818);
and U42448 (N_42448,N_37455,N_39030);
or U42449 (N_42449,N_36035,N_36050);
xnor U42450 (N_42450,N_36398,N_35288);
and U42451 (N_42451,N_36361,N_35736);
and U42452 (N_42452,N_36890,N_36005);
nor U42453 (N_42453,N_39216,N_38858);
and U42454 (N_42454,N_35584,N_38975);
xnor U42455 (N_42455,N_36270,N_37356);
and U42456 (N_42456,N_36952,N_35457);
or U42457 (N_42457,N_39257,N_36756);
nor U42458 (N_42458,N_38512,N_36431);
xor U42459 (N_42459,N_36339,N_35570);
or U42460 (N_42460,N_35366,N_35690);
or U42461 (N_42461,N_38400,N_37770);
nand U42462 (N_42462,N_36643,N_38012);
nor U42463 (N_42463,N_39204,N_39611);
and U42464 (N_42464,N_38756,N_37056);
xnor U42465 (N_42465,N_35708,N_39191);
and U42466 (N_42466,N_36886,N_37398);
nand U42467 (N_42467,N_35949,N_36595);
xnor U42468 (N_42468,N_36243,N_39558);
nand U42469 (N_42469,N_38517,N_37872);
nand U42470 (N_42470,N_38189,N_39280);
or U42471 (N_42471,N_36198,N_37033);
or U42472 (N_42472,N_36337,N_35173);
xor U42473 (N_42473,N_35661,N_38920);
nand U42474 (N_42474,N_37055,N_36626);
or U42475 (N_42475,N_38624,N_39774);
nor U42476 (N_42476,N_38366,N_35330);
xor U42477 (N_42477,N_35050,N_38981);
nor U42478 (N_42478,N_36855,N_35214);
and U42479 (N_42479,N_38927,N_39372);
or U42480 (N_42480,N_36311,N_39530);
or U42481 (N_42481,N_37045,N_36078);
or U42482 (N_42482,N_36576,N_38979);
nor U42483 (N_42483,N_38055,N_39607);
nor U42484 (N_42484,N_38154,N_38591);
xor U42485 (N_42485,N_39937,N_38046);
xor U42486 (N_42486,N_39032,N_38660);
and U42487 (N_42487,N_37295,N_38993);
xor U42488 (N_42488,N_35113,N_35026);
or U42489 (N_42489,N_38707,N_36288);
nand U42490 (N_42490,N_39120,N_37660);
xor U42491 (N_42491,N_39177,N_37759);
nand U42492 (N_42492,N_37050,N_39143);
or U42493 (N_42493,N_37465,N_38370);
nor U42494 (N_42494,N_38535,N_36525);
nand U42495 (N_42495,N_35886,N_39887);
nor U42496 (N_42496,N_36549,N_35515);
nor U42497 (N_42497,N_36940,N_36184);
nand U42498 (N_42498,N_35340,N_38138);
xnor U42499 (N_42499,N_37370,N_38903);
nor U42500 (N_42500,N_35428,N_38907);
and U42501 (N_42501,N_39759,N_35758);
xnor U42502 (N_42502,N_36767,N_35961);
nor U42503 (N_42503,N_39288,N_39824);
or U42504 (N_42504,N_38318,N_37668);
nor U42505 (N_42505,N_38911,N_37871);
and U42506 (N_42506,N_37277,N_37481);
nand U42507 (N_42507,N_37086,N_38945);
nand U42508 (N_42508,N_39499,N_36682);
or U42509 (N_42509,N_35771,N_35316);
xnor U42510 (N_42510,N_37542,N_39049);
xnor U42511 (N_42511,N_38936,N_38960);
nor U42512 (N_42512,N_39315,N_37639);
nand U42513 (N_42513,N_37105,N_39301);
xor U42514 (N_42514,N_37015,N_39413);
xor U42515 (N_42515,N_39874,N_37061);
or U42516 (N_42516,N_37143,N_35485);
nand U42517 (N_42517,N_38847,N_35150);
nand U42518 (N_42518,N_38852,N_35502);
nand U42519 (N_42519,N_37542,N_37558);
xor U42520 (N_42520,N_38238,N_39042);
and U42521 (N_42521,N_38660,N_38467);
or U42522 (N_42522,N_36320,N_37683);
or U42523 (N_42523,N_36517,N_38013);
nand U42524 (N_42524,N_36475,N_39335);
nand U42525 (N_42525,N_36735,N_36025);
xor U42526 (N_42526,N_35709,N_37472);
nand U42527 (N_42527,N_37432,N_39300);
or U42528 (N_42528,N_37301,N_39297);
nand U42529 (N_42529,N_37080,N_38047);
or U42530 (N_42530,N_39570,N_35460);
xnor U42531 (N_42531,N_36101,N_38978);
or U42532 (N_42532,N_35186,N_37864);
xnor U42533 (N_42533,N_35564,N_37411);
xnor U42534 (N_42534,N_36995,N_39358);
or U42535 (N_42535,N_35579,N_38768);
and U42536 (N_42536,N_39918,N_38794);
or U42537 (N_42537,N_39825,N_35939);
nor U42538 (N_42538,N_37412,N_39433);
or U42539 (N_42539,N_39750,N_37211);
or U42540 (N_42540,N_36611,N_38115);
and U42541 (N_42541,N_38864,N_38651);
or U42542 (N_42542,N_38824,N_35555);
and U42543 (N_42543,N_37004,N_36256);
xnor U42544 (N_42544,N_38355,N_37206);
or U42545 (N_42545,N_38094,N_38582);
and U42546 (N_42546,N_35493,N_35523);
and U42547 (N_42547,N_38230,N_37786);
or U42548 (N_42548,N_37397,N_36952);
or U42549 (N_42549,N_37652,N_37475);
xor U42550 (N_42550,N_35368,N_39991);
xor U42551 (N_42551,N_36533,N_37800);
or U42552 (N_42552,N_36064,N_35461);
nand U42553 (N_42553,N_38296,N_35097);
nor U42554 (N_42554,N_39014,N_35069);
or U42555 (N_42555,N_36682,N_37793);
or U42556 (N_42556,N_35196,N_37152);
and U42557 (N_42557,N_37732,N_36188);
or U42558 (N_42558,N_39040,N_35482);
xor U42559 (N_42559,N_36063,N_35786);
xor U42560 (N_42560,N_37465,N_35747);
and U42561 (N_42561,N_35484,N_38925);
nor U42562 (N_42562,N_38741,N_36435);
nor U42563 (N_42563,N_39118,N_37761);
and U42564 (N_42564,N_36993,N_39621);
nand U42565 (N_42565,N_38389,N_37467);
or U42566 (N_42566,N_36230,N_38816);
and U42567 (N_42567,N_36220,N_35548);
or U42568 (N_42568,N_39206,N_38538);
nor U42569 (N_42569,N_35941,N_36115);
and U42570 (N_42570,N_38140,N_36444);
xnor U42571 (N_42571,N_37287,N_38796);
or U42572 (N_42572,N_37976,N_37263);
or U42573 (N_42573,N_36334,N_37670);
nand U42574 (N_42574,N_35144,N_36635);
nor U42575 (N_42575,N_38211,N_39248);
and U42576 (N_42576,N_38846,N_38410);
nand U42577 (N_42577,N_39611,N_36791);
or U42578 (N_42578,N_35680,N_37468);
or U42579 (N_42579,N_38002,N_36134);
and U42580 (N_42580,N_36151,N_36799);
nand U42581 (N_42581,N_39030,N_37581);
nand U42582 (N_42582,N_35465,N_35224);
nor U42583 (N_42583,N_39144,N_37269);
and U42584 (N_42584,N_38858,N_36677);
xor U42585 (N_42585,N_37313,N_35585);
or U42586 (N_42586,N_39298,N_37130);
and U42587 (N_42587,N_39475,N_38702);
xnor U42588 (N_42588,N_37533,N_39757);
and U42589 (N_42589,N_39279,N_38133);
and U42590 (N_42590,N_36852,N_36927);
xor U42591 (N_42591,N_35265,N_39365);
or U42592 (N_42592,N_37784,N_37578);
and U42593 (N_42593,N_37179,N_36965);
nor U42594 (N_42594,N_38159,N_36397);
or U42595 (N_42595,N_37442,N_38838);
nand U42596 (N_42596,N_39032,N_38797);
nor U42597 (N_42597,N_39660,N_36739);
or U42598 (N_42598,N_37407,N_35512);
or U42599 (N_42599,N_35305,N_37307);
and U42600 (N_42600,N_39909,N_39384);
nor U42601 (N_42601,N_38185,N_38295);
nor U42602 (N_42602,N_38731,N_36992);
xnor U42603 (N_42603,N_36088,N_37957);
and U42604 (N_42604,N_35713,N_38444);
or U42605 (N_42605,N_36213,N_39289);
nand U42606 (N_42606,N_38161,N_36452);
xor U42607 (N_42607,N_35024,N_37111);
and U42608 (N_42608,N_36383,N_37810);
and U42609 (N_42609,N_37242,N_38371);
nand U42610 (N_42610,N_37950,N_37562);
xnor U42611 (N_42611,N_35591,N_39311);
nand U42612 (N_42612,N_38902,N_39123);
or U42613 (N_42613,N_35383,N_39646);
nand U42614 (N_42614,N_35097,N_38537);
or U42615 (N_42615,N_38837,N_37974);
nand U42616 (N_42616,N_37448,N_36436);
nor U42617 (N_42617,N_35831,N_35331);
xnor U42618 (N_42618,N_38471,N_37196);
and U42619 (N_42619,N_37926,N_39280);
xnor U42620 (N_42620,N_35310,N_38206);
nand U42621 (N_42621,N_36594,N_39619);
xnor U42622 (N_42622,N_36212,N_38597);
nand U42623 (N_42623,N_39648,N_39890);
or U42624 (N_42624,N_39142,N_38790);
nor U42625 (N_42625,N_38155,N_36026);
nand U42626 (N_42626,N_37979,N_37703);
nand U42627 (N_42627,N_36531,N_39908);
nand U42628 (N_42628,N_36021,N_35740);
nand U42629 (N_42629,N_37404,N_36315);
nand U42630 (N_42630,N_37549,N_37998);
nor U42631 (N_42631,N_36679,N_36217);
nor U42632 (N_42632,N_38146,N_35080);
xnor U42633 (N_42633,N_38830,N_38325);
xor U42634 (N_42634,N_36260,N_36992);
nor U42635 (N_42635,N_35191,N_37046);
nand U42636 (N_42636,N_38256,N_39462);
xor U42637 (N_42637,N_36657,N_39222);
nor U42638 (N_42638,N_36954,N_38512);
and U42639 (N_42639,N_35458,N_35455);
and U42640 (N_42640,N_37698,N_36232);
or U42641 (N_42641,N_38285,N_37848);
nor U42642 (N_42642,N_35026,N_35023);
or U42643 (N_42643,N_35740,N_35583);
xnor U42644 (N_42644,N_37591,N_35321);
or U42645 (N_42645,N_39609,N_37231);
or U42646 (N_42646,N_37324,N_37011);
nand U42647 (N_42647,N_38667,N_35917);
xor U42648 (N_42648,N_35338,N_38264);
xor U42649 (N_42649,N_39337,N_37311);
xor U42650 (N_42650,N_35990,N_38595);
nand U42651 (N_42651,N_36879,N_38580);
and U42652 (N_42652,N_37154,N_37070);
xor U42653 (N_42653,N_38474,N_39587);
nor U42654 (N_42654,N_35445,N_37646);
nand U42655 (N_42655,N_37429,N_35266);
xnor U42656 (N_42656,N_38442,N_35447);
nor U42657 (N_42657,N_39230,N_39586);
nor U42658 (N_42658,N_37133,N_38526);
nand U42659 (N_42659,N_37795,N_39718);
or U42660 (N_42660,N_37264,N_39022);
or U42661 (N_42661,N_38798,N_39643);
nand U42662 (N_42662,N_39792,N_35814);
nor U42663 (N_42663,N_38716,N_37296);
xnor U42664 (N_42664,N_36402,N_35621);
nand U42665 (N_42665,N_38983,N_36939);
xor U42666 (N_42666,N_38940,N_35815);
and U42667 (N_42667,N_36050,N_35469);
or U42668 (N_42668,N_36742,N_36511);
or U42669 (N_42669,N_37664,N_37544);
or U42670 (N_42670,N_36037,N_36708);
nand U42671 (N_42671,N_38838,N_38244);
nand U42672 (N_42672,N_38270,N_38766);
and U42673 (N_42673,N_38069,N_39506);
xor U42674 (N_42674,N_38969,N_36805);
xor U42675 (N_42675,N_38209,N_38101);
and U42676 (N_42676,N_36514,N_38453);
or U42677 (N_42677,N_37021,N_38347);
nand U42678 (N_42678,N_37994,N_38956);
xor U42679 (N_42679,N_39272,N_38965);
nand U42680 (N_42680,N_39150,N_37776);
xnor U42681 (N_42681,N_36479,N_37497);
xor U42682 (N_42682,N_38865,N_36711);
and U42683 (N_42683,N_37184,N_35466);
nor U42684 (N_42684,N_35488,N_38604);
xnor U42685 (N_42685,N_36593,N_35529);
or U42686 (N_42686,N_36352,N_36253);
nor U42687 (N_42687,N_38315,N_39462);
nand U42688 (N_42688,N_36792,N_36444);
xor U42689 (N_42689,N_38838,N_36298);
nand U42690 (N_42690,N_35602,N_38759);
or U42691 (N_42691,N_37501,N_39986);
or U42692 (N_42692,N_35157,N_38311);
xnor U42693 (N_42693,N_38714,N_38732);
and U42694 (N_42694,N_36553,N_37304);
or U42695 (N_42695,N_39934,N_35989);
nand U42696 (N_42696,N_35670,N_35399);
nor U42697 (N_42697,N_38549,N_38655);
or U42698 (N_42698,N_38623,N_37311);
xor U42699 (N_42699,N_35578,N_36997);
and U42700 (N_42700,N_38993,N_37450);
or U42701 (N_42701,N_39524,N_37215);
and U42702 (N_42702,N_36432,N_38244);
nand U42703 (N_42703,N_37264,N_39124);
or U42704 (N_42704,N_36590,N_39497);
nand U42705 (N_42705,N_35252,N_37291);
xor U42706 (N_42706,N_38780,N_39875);
nand U42707 (N_42707,N_35792,N_36183);
and U42708 (N_42708,N_37553,N_37989);
or U42709 (N_42709,N_36101,N_36061);
or U42710 (N_42710,N_39527,N_35816);
nand U42711 (N_42711,N_35093,N_35149);
xor U42712 (N_42712,N_38956,N_35692);
and U42713 (N_42713,N_38171,N_36825);
or U42714 (N_42714,N_38078,N_38821);
nor U42715 (N_42715,N_36711,N_36028);
and U42716 (N_42716,N_37744,N_39400);
or U42717 (N_42717,N_39044,N_38014);
and U42718 (N_42718,N_39964,N_39106);
nand U42719 (N_42719,N_36744,N_36848);
or U42720 (N_42720,N_36342,N_37634);
xor U42721 (N_42721,N_37024,N_38246);
nand U42722 (N_42722,N_39419,N_37651);
nand U42723 (N_42723,N_37822,N_39175);
nand U42724 (N_42724,N_36456,N_37838);
and U42725 (N_42725,N_38670,N_39012);
nand U42726 (N_42726,N_36291,N_39084);
nor U42727 (N_42727,N_38351,N_35194);
xnor U42728 (N_42728,N_39627,N_37729);
and U42729 (N_42729,N_39097,N_39440);
or U42730 (N_42730,N_35286,N_36128);
xnor U42731 (N_42731,N_38075,N_35099);
and U42732 (N_42732,N_39439,N_36430);
xor U42733 (N_42733,N_35360,N_39146);
nand U42734 (N_42734,N_39009,N_39481);
nor U42735 (N_42735,N_39455,N_37181);
nor U42736 (N_42736,N_36002,N_35109);
nor U42737 (N_42737,N_38647,N_37304);
nand U42738 (N_42738,N_38866,N_37103);
nor U42739 (N_42739,N_37732,N_39361);
or U42740 (N_42740,N_37924,N_36022);
or U42741 (N_42741,N_39338,N_35538);
nand U42742 (N_42742,N_37374,N_36427);
or U42743 (N_42743,N_39777,N_35732);
xnor U42744 (N_42744,N_36147,N_39712);
nand U42745 (N_42745,N_38733,N_35155);
or U42746 (N_42746,N_38010,N_37322);
xnor U42747 (N_42747,N_39773,N_35909);
and U42748 (N_42748,N_37752,N_36006);
or U42749 (N_42749,N_37236,N_37703);
nand U42750 (N_42750,N_37979,N_39917);
and U42751 (N_42751,N_36763,N_38205);
or U42752 (N_42752,N_36676,N_37875);
or U42753 (N_42753,N_38258,N_36705);
nand U42754 (N_42754,N_39569,N_36969);
nand U42755 (N_42755,N_35087,N_38205);
or U42756 (N_42756,N_35685,N_36703);
nand U42757 (N_42757,N_36731,N_37635);
or U42758 (N_42758,N_38494,N_37370);
nor U42759 (N_42759,N_37083,N_36574);
and U42760 (N_42760,N_36941,N_36108);
or U42761 (N_42761,N_38582,N_38125);
or U42762 (N_42762,N_39970,N_38360);
nand U42763 (N_42763,N_36248,N_39709);
nor U42764 (N_42764,N_39665,N_39277);
nor U42765 (N_42765,N_35055,N_38204);
nor U42766 (N_42766,N_35733,N_35051);
and U42767 (N_42767,N_37494,N_37121);
or U42768 (N_42768,N_37447,N_38521);
nand U42769 (N_42769,N_36032,N_39075);
xor U42770 (N_42770,N_39884,N_37395);
xnor U42771 (N_42771,N_39883,N_39043);
and U42772 (N_42772,N_35085,N_35194);
nor U42773 (N_42773,N_39713,N_36778);
xor U42774 (N_42774,N_37272,N_38724);
xnor U42775 (N_42775,N_38010,N_35454);
or U42776 (N_42776,N_39034,N_36299);
and U42777 (N_42777,N_35412,N_39891);
nand U42778 (N_42778,N_35875,N_38671);
xor U42779 (N_42779,N_39689,N_38616);
and U42780 (N_42780,N_36403,N_38462);
or U42781 (N_42781,N_35042,N_38292);
nand U42782 (N_42782,N_35061,N_37181);
nor U42783 (N_42783,N_35204,N_38300);
xor U42784 (N_42784,N_36104,N_35611);
and U42785 (N_42785,N_36847,N_36939);
nand U42786 (N_42786,N_36356,N_39520);
xnor U42787 (N_42787,N_38424,N_39599);
or U42788 (N_42788,N_38308,N_38694);
nor U42789 (N_42789,N_39010,N_38056);
and U42790 (N_42790,N_38839,N_39534);
nor U42791 (N_42791,N_36192,N_38076);
xor U42792 (N_42792,N_37404,N_37178);
or U42793 (N_42793,N_39759,N_37313);
nand U42794 (N_42794,N_37095,N_35378);
and U42795 (N_42795,N_39347,N_38084);
xor U42796 (N_42796,N_36471,N_39592);
xor U42797 (N_42797,N_39966,N_37297);
nor U42798 (N_42798,N_38270,N_39619);
xnor U42799 (N_42799,N_35952,N_37260);
and U42800 (N_42800,N_36430,N_35377);
or U42801 (N_42801,N_38572,N_36564);
and U42802 (N_42802,N_36455,N_37441);
nand U42803 (N_42803,N_37565,N_37299);
xor U42804 (N_42804,N_36100,N_39800);
or U42805 (N_42805,N_37502,N_37051);
nor U42806 (N_42806,N_38864,N_38459);
xnor U42807 (N_42807,N_39510,N_39570);
nor U42808 (N_42808,N_36187,N_39054);
nor U42809 (N_42809,N_38589,N_39152);
xnor U42810 (N_42810,N_38840,N_37231);
and U42811 (N_42811,N_39401,N_37580);
or U42812 (N_42812,N_36133,N_36265);
and U42813 (N_42813,N_36293,N_38089);
or U42814 (N_42814,N_38840,N_37222);
nor U42815 (N_42815,N_35055,N_37031);
xnor U42816 (N_42816,N_36076,N_37270);
or U42817 (N_42817,N_37514,N_35162);
and U42818 (N_42818,N_38185,N_38000);
or U42819 (N_42819,N_38439,N_36101);
nor U42820 (N_42820,N_36775,N_37326);
nand U42821 (N_42821,N_35711,N_38857);
xor U42822 (N_42822,N_38312,N_37218);
and U42823 (N_42823,N_35092,N_36012);
xnor U42824 (N_42824,N_38840,N_39113);
and U42825 (N_42825,N_37925,N_37537);
or U42826 (N_42826,N_36232,N_39265);
nor U42827 (N_42827,N_38126,N_38042);
nor U42828 (N_42828,N_36410,N_37551);
nor U42829 (N_42829,N_37700,N_36792);
nor U42830 (N_42830,N_35234,N_35540);
xor U42831 (N_42831,N_36547,N_36874);
nor U42832 (N_42832,N_38167,N_35058);
nor U42833 (N_42833,N_37305,N_36248);
nor U42834 (N_42834,N_36641,N_39308);
and U42835 (N_42835,N_36829,N_37770);
and U42836 (N_42836,N_35204,N_39430);
nand U42837 (N_42837,N_37871,N_35690);
and U42838 (N_42838,N_38979,N_37743);
or U42839 (N_42839,N_37234,N_39870);
nand U42840 (N_42840,N_35225,N_36345);
and U42841 (N_42841,N_36181,N_39492);
nand U42842 (N_42842,N_37305,N_37745);
or U42843 (N_42843,N_37589,N_39481);
and U42844 (N_42844,N_38795,N_39222);
nor U42845 (N_42845,N_36255,N_36881);
xor U42846 (N_42846,N_38531,N_38352);
or U42847 (N_42847,N_39794,N_39034);
or U42848 (N_42848,N_37951,N_37095);
or U42849 (N_42849,N_38610,N_37352);
nor U42850 (N_42850,N_36076,N_37835);
xnor U42851 (N_42851,N_38885,N_39052);
nand U42852 (N_42852,N_38395,N_36347);
and U42853 (N_42853,N_39262,N_36655);
and U42854 (N_42854,N_35525,N_39727);
nand U42855 (N_42855,N_39063,N_39575);
nor U42856 (N_42856,N_36135,N_37924);
nor U42857 (N_42857,N_35442,N_35713);
xor U42858 (N_42858,N_38403,N_38094);
nor U42859 (N_42859,N_38108,N_36348);
nor U42860 (N_42860,N_35227,N_38477);
nor U42861 (N_42861,N_36428,N_35765);
and U42862 (N_42862,N_37453,N_35948);
or U42863 (N_42863,N_35487,N_37462);
nand U42864 (N_42864,N_38658,N_35734);
nor U42865 (N_42865,N_37657,N_39236);
nand U42866 (N_42866,N_35173,N_38251);
or U42867 (N_42867,N_35659,N_36195);
and U42868 (N_42868,N_37660,N_37424);
and U42869 (N_42869,N_38462,N_39585);
xnor U42870 (N_42870,N_35031,N_37635);
or U42871 (N_42871,N_35789,N_36879);
xor U42872 (N_42872,N_38611,N_35271);
nor U42873 (N_42873,N_37034,N_35128);
nand U42874 (N_42874,N_37755,N_38539);
or U42875 (N_42875,N_39400,N_36452);
or U42876 (N_42876,N_39192,N_35014);
nor U42877 (N_42877,N_39272,N_38874);
xor U42878 (N_42878,N_38382,N_36357);
xnor U42879 (N_42879,N_39654,N_35764);
or U42880 (N_42880,N_35100,N_38609);
or U42881 (N_42881,N_39558,N_38353);
or U42882 (N_42882,N_37982,N_39792);
nor U42883 (N_42883,N_37397,N_38305);
nand U42884 (N_42884,N_37396,N_35944);
nor U42885 (N_42885,N_38379,N_37619);
or U42886 (N_42886,N_36003,N_35800);
xnor U42887 (N_42887,N_36928,N_39340);
or U42888 (N_42888,N_35702,N_37990);
xor U42889 (N_42889,N_38409,N_36135);
or U42890 (N_42890,N_35133,N_37799);
or U42891 (N_42891,N_35923,N_37054);
nor U42892 (N_42892,N_35320,N_35517);
or U42893 (N_42893,N_38232,N_38347);
and U42894 (N_42894,N_35122,N_39775);
or U42895 (N_42895,N_38621,N_39613);
nor U42896 (N_42896,N_35201,N_35670);
and U42897 (N_42897,N_35790,N_36111);
xnor U42898 (N_42898,N_35429,N_37231);
nand U42899 (N_42899,N_39680,N_38426);
nor U42900 (N_42900,N_35907,N_37379);
nor U42901 (N_42901,N_38465,N_38593);
and U42902 (N_42902,N_36525,N_37142);
or U42903 (N_42903,N_37887,N_39430);
or U42904 (N_42904,N_38360,N_35320);
xnor U42905 (N_42905,N_35822,N_37378);
nand U42906 (N_42906,N_36987,N_39267);
or U42907 (N_42907,N_35656,N_35852);
and U42908 (N_42908,N_36324,N_35538);
xor U42909 (N_42909,N_35346,N_37774);
nand U42910 (N_42910,N_38910,N_36204);
and U42911 (N_42911,N_37277,N_38782);
and U42912 (N_42912,N_36936,N_35882);
and U42913 (N_42913,N_37286,N_37934);
and U42914 (N_42914,N_38506,N_37068);
nand U42915 (N_42915,N_35196,N_38880);
xnor U42916 (N_42916,N_39051,N_38706);
and U42917 (N_42917,N_37657,N_36405);
or U42918 (N_42918,N_36707,N_39106);
nor U42919 (N_42919,N_36646,N_36312);
nor U42920 (N_42920,N_35092,N_38226);
xnor U42921 (N_42921,N_38801,N_36096);
and U42922 (N_42922,N_35975,N_35010);
nand U42923 (N_42923,N_35545,N_38246);
nand U42924 (N_42924,N_39022,N_35671);
nand U42925 (N_42925,N_36876,N_36477);
nand U42926 (N_42926,N_38583,N_39224);
and U42927 (N_42927,N_38238,N_37627);
and U42928 (N_42928,N_37324,N_35897);
xor U42929 (N_42929,N_35145,N_37732);
or U42930 (N_42930,N_38732,N_35893);
nor U42931 (N_42931,N_36243,N_39691);
nand U42932 (N_42932,N_37197,N_39711);
or U42933 (N_42933,N_36899,N_38885);
xnor U42934 (N_42934,N_39980,N_38856);
xor U42935 (N_42935,N_36302,N_35157);
xnor U42936 (N_42936,N_38212,N_39377);
or U42937 (N_42937,N_39075,N_39098);
or U42938 (N_42938,N_38818,N_35012);
and U42939 (N_42939,N_37339,N_36831);
and U42940 (N_42940,N_36250,N_36125);
nand U42941 (N_42941,N_37909,N_38764);
and U42942 (N_42942,N_37453,N_38526);
or U42943 (N_42943,N_36314,N_36512);
nand U42944 (N_42944,N_36225,N_38135);
or U42945 (N_42945,N_35791,N_36809);
and U42946 (N_42946,N_36545,N_39216);
or U42947 (N_42947,N_37251,N_39461);
nand U42948 (N_42948,N_36029,N_37194);
nor U42949 (N_42949,N_35727,N_35687);
nand U42950 (N_42950,N_35495,N_38059);
xnor U42951 (N_42951,N_35530,N_36326);
and U42952 (N_42952,N_35656,N_38507);
or U42953 (N_42953,N_38437,N_39231);
nand U42954 (N_42954,N_38900,N_35911);
and U42955 (N_42955,N_37602,N_38789);
and U42956 (N_42956,N_37127,N_38333);
nor U42957 (N_42957,N_36687,N_36201);
or U42958 (N_42958,N_37616,N_39304);
or U42959 (N_42959,N_36929,N_39075);
or U42960 (N_42960,N_36343,N_39573);
or U42961 (N_42961,N_39219,N_39281);
xor U42962 (N_42962,N_37728,N_38409);
nor U42963 (N_42963,N_36475,N_37311);
xor U42964 (N_42964,N_38517,N_37014);
nor U42965 (N_42965,N_35295,N_39982);
nand U42966 (N_42966,N_37701,N_37031);
nor U42967 (N_42967,N_35263,N_35866);
nor U42968 (N_42968,N_35420,N_35437);
nand U42969 (N_42969,N_35345,N_39514);
or U42970 (N_42970,N_38115,N_39085);
or U42971 (N_42971,N_37974,N_38406);
and U42972 (N_42972,N_36241,N_37245);
and U42973 (N_42973,N_37148,N_35560);
or U42974 (N_42974,N_37663,N_37454);
or U42975 (N_42975,N_38894,N_38495);
and U42976 (N_42976,N_37472,N_37762);
or U42977 (N_42977,N_35781,N_37330);
xnor U42978 (N_42978,N_37873,N_37872);
nor U42979 (N_42979,N_38164,N_37378);
nor U42980 (N_42980,N_38421,N_37023);
nor U42981 (N_42981,N_36752,N_38793);
nand U42982 (N_42982,N_39871,N_36624);
nand U42983 (N_42983,N_38078,N_35492);
and U42984 (N_42984,N_36188,N_39696);
nand U42985 (N_42985,N_37162,N_36982);
nand U42986 (N_42986,N_38030,N_37264);
nor U42987 (N_42987,N_37781,N_38374);
or U42988 (N_42988,N_35988,N_37233);
xnor U42989 (N_42989,N_38222,N_39994);
nor U42990 (N_42990,N_39785,N_38953);
and U42991 (N_42991,N_37203,N_38453);
or U42992 (N_42992,N_36600,N_35194);
xnor U42993 (N_42993,N_37347,N_37394);
xnor U42994 (N_42994,N_39125,N_35177);
and U42995 (N_42995,N_39233,N_38176);
nor U42996 (N_42996,N_35675,N_37961);
xnor U42997 (N_42997,N_36387,N_36471);
nor U42998 (N_42998,N_38355,N_37578);
nor U42999 (N_42999,N_38782,N_39082);
xnor U43000 (N_43000,N_36645,N_39658);
and U43001 (N_43001,N_39704,N_39160);
nand U43002 (N_43002,N_36417,N_35086);
xnor U43003 (N_43003,N_38380,N_36387);
nor U43004 (N_43004,N_38362,N_37337);
nand U43005 (N_43005,N_38825,N_36597);
and U43006 (N_43006,N_39760,N_38426);
nor U43007 (N_43007,N_37062,N_37054);
or U43008 (N_43008,N_38744,N_37212);
nor U43009 (N_43009,N_37582,N_35001);
nand U43010 (N_43010,N_38031,N_39545);
and U43011 (N_43011,N_36999,N_35621);
xnor U43012 (N_43012,N_38216,N_39725);
and U43013 (N_43013,N_36690,N_35704);
nor U43014 (N_43014,N_35949,N_38296);
and U43015 (N_43015,N_39111,N_38048);
xor U43016 (N_43016,N_36650,N_37424);
nor U43017 (N_43017,N_38513,N_38402);
nand U43018 (N_43018,N_35571,N_37554);
nand U43019 (N_43019,N_38220,N_37053);
and U43020 (N_43020,N_39252,N_37037);
xor U43021 (N_43021,N_38663,N_35085);
nor U43022 (N_43022,N_38996,N_36049);
nor U43023 (N_43023,N_39922,N_38572);
nand U43024 (N_43024,N_37751,N_36958);
or U43025 (N_43025,N_35735,N_39446);
or U43026 (N_43026,N_37926,N_35701);
or U43027 (N_43027,N_38321,N_35950);
or U43028 (N_43028,N_39732,N_39127);
and U43029 (N_43029,N_37784,N_36343);
or U43030 (N_43030,N_37891,N_38148);
xor U43031 (N_43031,N_35997,N_38149);
nor U43032 (N_43032,N_35610,N_39716);
nor U43033 (N_43033,N_38683,N_38759);
nor U43034 (N_43034,N_39855,N_39259);
and U43035 (N_43035,N_39924,N_37210);
or U43036 (N_43036,N_39693,N_37310);
and U43037 (N_43037,N_35116,N_35688);
nor U43038 (N_43038,N_37594,N_35841);
nor U43039 (N_43039,N_39413,N_39979);
nand U43040 (N_43040,N_38313,N_37642);
and U43041 (N_43041,N_36901,N_37915);
and U43042 (N_43042,N_35894,N_38758);
xnor U43043 (N_43043,N_38378,N_37582);
nor U43044 (N_43044,N_38730,N_35116);
xor U43045 (N_43045,N_37073,N_38283);
nand U43046 (N_43046,N_36469,N_38061);
and U43047 (N_43047,N_39297,N_39234);
and U43048 (N_43048,N_35835,N_37289);
or U43049 (N_43049,N_38214,N_38807);
nand U43050 (N_43050,N_39451,N_35708);
or U43051 (N_43051,N_39922,N_39272);
xor U43052 (N_43052,N_39764,N_35519);
nand U43053 (N_43053,N_36070,N_39280);
and U43054 (N_43054,N_36727,N_35327);
nor U43055 (N_43055,N_39536,N_35610);
nand U43056 (N_43056,N_36103,N_39016);
or U43057 (N_43057,N_35445,N_37121);
and U43058 (N_43058,N_39682,N_38152);
nor U43059 (N_43059,N_38989,N_35162);
nor U43060 (N_43060,N_39646,N_36191);
xor U43061 (N_43061,N_35220,N_35308);
nand U43062 (N_43062,N_39989,N_38898);
and U43063 (N_43063,N_36983,N_36839);
nor U43064 (N_43064,N_36347,N_39490);
nor U43065 (N_43065,N_35517,N_37040);
nor U43066 (N_43066,N_37379,N_37766);
or U43067 (N_43067,N_38262,N_37534);
xnor U43068 (N_43068,N_35637,N_35445);
xnor U43069 (N_43069,N_39170,N_36035);
or U43070 (N_43070,N_38079,N_37885);
nor U43071 (N_43071,N_35919,N_35887);
and U43072 (N_43072,N_36248,N_38905);
xor U43073 (N_43073,N_37274,N_39523);
nor U43074 (N_43074,N_37694,N_39707);
and U43075 (N_43075,N_37013,N_36701);
nor U43076 (N_43076,N_38165,N_38602);
nand U43077 (N_43077,N_36701,N_37345);
nor U43078 (N_43078,N_39075,N_38178);
nor U43079 (N_43079,N_38066,N_35113);
or U43080 (N_43080,N_37682,N_35268);
and U43081 (N_43081,N_36119,N_38430);
xor U43082 (N_43082,N_37688,N_37400);
xnor U43083 (N_43083,N_37801,N_37855);
xnor U43084 (N_43084,N_35949,N_36565);
xnor U43085 (N_43085,N_36140,N_38525);
and U43086 (N_43086,N_35270,N_36258);
xor U43087 (N_43087,N_36866,N_35321);
nor U43088 (N_43088,N_35950,N_39576);
nor U43089 (N_43089,N_37277,N_39489);
nand U43090 (N_43090,N_36564,N_39829);
nand U43091 (N_43091,N_36003,N_35229);
xor U43092 (N_43092,N_38134,N_36154);
nand U43093 (N_43093,N_38213,N_35097);
xnor U43094 (N_43094,N_37467,N_35849);
and U43095 (N_43095,N_38819,N_36980);
nand U43096 (N_43096,N_35494,N_35325);
and U43097 (N_43097,N_37105,N_39073);
nor U43098 (N_43098,N_37371,N_36361);
nand U43099 (N_43099,N_39020,N_38508);
nand U43100 (N_43100,N_38451,N_35950);
and U43101 (N_43101,N_37380,N_37179);
nand U43102 (N_43102,N_36563,N_37803);
nand U43103 (N_43103,N_39283,N_36555);
nand U43104 (N_43104,N_36382,N_39538);
nor U43105 (N_43105,N_35419,N_38820);
nor U43106 (N_43106,N_37166,N_36571);
xor U43107 (N_43107,N_38978,N_39859);
xnor U43108 (N_43108,N_35045,N_36074);
or U43109 (N_43109,N_35404,N_35499);
nand U43110 (N_43110,N_36007,N_37676);
nand U43111 (N_43111,N_39154,N_37039);
or U43112 (N_43112,N_36357,N_37928);
or U43113 (N_43113,N_38656,N_35706);
nor U43114 (N_43114,N_39395,N_36589);
xnor U43115 (N_43115,N_37089,N_36256);
or U43116 (N_43116,N_38466,N_38504);
nand U43117 (N_43117,N_37494,N_39963);
nand U43118 (N_43118,N_37198,N_36326);
or U43119 (N_43119,N_37099,N_38142);
nor U43120 (N_43120,N_39262,N_38921);
and U43121 (N_43121,N_36557,N_35386);
and U43122 (N_43122,N_38614,N_38742);
or U43123 (N_43123,N_39853,N_35766);
and U43124 (N_43124,N_35312,N_38627);
xor U43125 (N_43125,N_38353,N_38671);
or U43126 (N_43126,N_38943,N_39789);
or U43127 (N_43127,N_38718,N_37990);
or U43128 (N_43128,N_37777,N_39703);
xor U43129 (N_43129,N_36714,N_37106);
nor U43130 (N_43130,N_35341,N_35254);
and U43131 (N_43131,N_38434,N_37502);
xor U43132 (N_43132,N_38374,N_39883);
and U43133 (N_43133,N_38962,N_35867);
and U43134 (N_43134,N_38527,N_35748);
or U43135 (N_43135,N_36522,N_36594);
or U43136 (N_43136,N_38657,N_38386);
and U43137 (N_43137,N_36938,N_38284);
xnor U43138 (N_43138,N_35317,N_36828);
and U43139 (N_43139,N_35440,N_39774);
and U43140 (N_43140,N_39325,N_38735);
xor U43141 (N_43141,N_36712,N_36660);
nand U43142 (N_43142,N_39430,N_35500);
nand U43143 (N_43143,N_39111,N_37122);
and U43144 (N_43144,N_35891,N_35899);
or U43145 (N_43145,N_36423,N_38102);
or U43146 (N_43146,N_37390,N_37820);
or U43147 (N_43147,N_39231,N_37997);
nor U43148 (N_43148,N_38891,N_39821);
and U43149 (N_43149,N_36783,N_35761);
nor U43150 (N_43150,N_37964,N_39112);
nand U43151 (N_43151,N_39933,N_38780);
xnor U43152 (N_43152,N_35068,N_37868);
xor U43153 (N_43153,N_37811,N_38274);
and U43154 (N_43154,N_35153,N_39971);
xnor U43155 (N_43155,N_38529,N_36637);
nand U43156 (N_43156,N_36468,N_38233);
or U43157 (N_43157,N_37580,N_39063);
and U43158 (N_43158,N_39240,N_35992);
xor U43159 (N_43159,N_38377,N_35095);
xor U43160 (N_43160,N_39576,N_37442);
or U43161 (N_43161,N_36954,N_36668);
or U43162 (N_43162,N_36760,N_35903);
and U43163 (N_43163,N_38530,N_37695);
nand U43164 (N_43164,N_36869,N_37762);
or U43165 (N_43165,N_35939,N_36812);
nor U43166 (N_43166,N_39496,N_37619);
xnor U43167 (N_43167,N_39168,N_37547);
nor U43168 (N_43168,N_37128,N_35744);
and U43169 (N_43169,N_37864,N_35632);
and U43170 (N_43170,N_36487,N_36872);
nand U43171 (N_43171,N_37219,N_37708);
or U43172 (N_43172,N_36824,N_37931);
and U43173 (N_43173,N_38674,N_38193);
xnor U43174 (N_43174,N_38016,N_38256);
nand U43175 (N_43175,N_37382,N_35650);
xor U43176 (N_43176,N_36371,N_39761);
nand U43177 (N_43177,N_37474,N_36688);
nand U43178 (N_43178,N_39093,N_38844);
nor U43179 (N_43179,N_37909,N_35405);
nor U43180 (N_43180,N_36682,N_36717);
or U43181 (N_43181,N_36472,N_37553);
or U43182 (N_43182,N_36110,N_39530);
or U43183 (N_43183,N_39693,N_37499);
or U43184 (N_43184,N_35952,N_36952);
xor U43185 (N_43185,N_37377,N_36088);
and U43186 (N_43186,N_39987,N_39837);
nor U43187 (N_43187,N_38601,N_35883);
or U43188 (N_43188,N_38712,N_37838);
xor U43189 (N_43189,N_37880,N_37566);
nand U43190 (N_43190,N_36194,N_39696);
xor U43191 (N_43191,N_37443,N_37150);
nand U43192 (N_43192,N_38600,N_39165);
xor U43193 (N_43193,N_35385,N_37428);
nand U43194 (N_43194,N_38305,N_36743);
nor U43195 (N_43195,N_38443,N_36284);
and U43196 (N_43196,N_37889,N_36271);
xnor U43197 (N_43197,N_38803,N_39396);
nand U43198 (N_43198,N_36673,N_35807);
nor U43199 (N_43199,N_38553,N_35041);
xor U43200 (N_43200,N_35873,N_35387);
or U43201 (N_43201,N_36163,N_38194);
and U43202 (N_43202,N_38666,N_35715);
xnor U43203 (N_43203,N_37680,N_35600);
xor U43204 (N_43204,N_36525,N_36603);
and U43205 (N_43205,N_39497,N_39694);
nor U43206 (N_43206,N_39898,N_39355);
nor U43207 (N_43207,N_38350,N_39874);
or U43208 (N_43208,N_39944,N_36555);
nand U43209 (N_43209,N_37962,N_36897);
and U43210 (N_43210,N_37351,N_39037);
nor U43211 (N_43211,N_38093,N_35660);
nand U43212 (N_43212,N_38774,N_39854);
nor U43213 (N_43213,N_38485,N_38433);
or U43214 (N_43214,N_37607,N_35540);
xor U43215 (N_43215,N_38817,N_36418);
or U43216 (N_43216,N_35961,N_36475);
nand U43217 (N_43217,N_38412,N_35995);
and U43218 (N_43218,N_35904,N_37731);
or U43219 (N_43219,N_36552,N_38862);
xnor U43220 (N_43220,N_37454,N_38925);
or U43221 (N_43221,N_39162,N_39309);
xnor U43222 (N_43222,N_37194,N_39182);
or U43223 (N_43223,N_39362,N_38867);
nand U43224 (N_43224,N_37200,N_36551);
xor U43225 (N_43225,N_38338,N_38689);
nand U43226 (N_43226,N_35794,N_36865);
nor U43227 (N_43227,N_35168,N_39482);
nand U43228 (N_43228,N_37869,N_35376);
or U43229 (N_43229,N_37439,N_38738);
and U43230 (N_43230,N_37701,N_39758);
and U43231 (N_43231,N_36578,N_37001);
nor U43232 (N_43232,N_38766,N_38607);
nor U43233 (N_43233,N_37584,N_37521);
or U43234 (N_43234,N_35306,N_38178);
and U43235 (N_43235,N_35389,N_35825);
or U43236 (N_43236,N_37518,N_38639);
nand U43237 (N_43237,N_39580,N_37723);
or U43238 (N_43238,N_35997,N_39396);
nand U43239 (N_43239,N_35858,N_38496);
nand U43240 (N_43240,N_35701,N_38854);
nand U43241 (N_43241,N_38007,N_35057);
xnor U43242 (N_43242,N_35926,N_36388);
and U43243 (N_43243,N_39435,N_38137);
and U43244 (N_43244,N_37952,N_36556);
and U43245 (N_43245,N_37614,N_36520);
nor U43246 (N_43246,N_35781,N_37511);
xor U43247 (N_43247,N_37761,N_37350);
xor U43248 (N_43248,N_35353,N_36407);
and U43249 (N_43249,N_37911,N_37434);
nor U43250 (N_43250,N_39216,N_38347);
and U43251 (N_43251,N_38180,N_37652);
and U43252 (N_43252,N_37198,N_38480);
or U43253 (N_43253,N_35116,N_35739);
nand U43254 (N_43254,N_36451,N_38177);
nand U43255 (N_43255,N_36602,N_37799);
nand U43256 (N_43256,N_37062,N_39539);
and U43257 (N_43257,N_39656,N_35157);
and U43258 (N_43258,N_38078,N_39933);
nand U43259 (N_43259,N_39949,N_36946);
nand U43260 (N_43260,N_39353,N_37905);
and U43261 (N_43261,N_39421,N_36634);
or U43262 (N_43262,N_38759,N_37109);
nor U43263 (N_43263,N_39716,N_37066);
or U43264 (N_43264,N_36405,N_38780);
or U43265 (N_43265,N_38662,N_37586);
nand U43266 (N_43266,N_38415,N_37971);
or U43267 (N_43267,N_39089,N_37562);
nor U43268 (N_43268,N_38293,N_39750);
or U43269 (N_43269,N_35778,N_36896);
or U43270 (N_43270,N_38492,N_35323);
nor U43271 (N_43271,N_36815,N_38613);
nand U43272 (N_43272,N_39464,N_38729);
nand U43273 (N_43273,N_37028,N_35546);
xnor U43274 (N_43274,N_35636,N_36007);
nand U43275 (N_43275,N_36187,N_38002);
xnor U43276 (N_43276,N_36536,N_35903);
xnor U43277 (N_43277,N_39004,N_35568);
nand U43278 (N_43278,N_39972,N_38916);
nor U43279 (N_43279,N_38746,N_39280);
or U43280 (N_43280,N_39125,N_36975);
xnor U43281 (N_43281,N_38503,N_36412);
or U43282 (N_43282,N_38306,N_37385);
and U43283 (N_43283,N_39597,N_37832);
xnor U43284 (N_43284,N_37763,N_38052);
nor U43285 (N_43285,N_35773,N_38593);
nor U43286 (N_43286,N_35940,N_38846);
or U43287 (N_43287,N_37725,N_39379);
or U43288 (N_43288,N_37158,N_38220);
nand U43289 (N_43289,N_35091,N_39437);
nand U43290 (N_43290,N_35189,N_35267);
xor U43291 (N_43291,N_38063,N_38454);
nand U43292 (N_43292,N_39746,N_35448);
nand U43293 (N_43293,N_37140,N_35876);
or U43294 (N_43294,N_37461,N_36834);
nand U43295 (N_43295,N_39826,N_37493);
or U43296 (N_43296,N_35057,N_36893);
or U43297 (N_43297,N_39038,N_38170);
or U43298 (N_43298,N_38714,N_38595);
nand U43299 (N_43299,N_35697,N_37097);
or U43300 (N_43300,N_36504,N_38875);
xor U43301 (N_43301,N_35646,N_37785);
and U43302 (N_43302,N_36335,N_38634);
nor U43303 (N_43303,N_36792,N_38696);
and U43304 (N_43304,N_38480,N_39463);
or U43305 (N_43305,N_36942,N_39792);
or U43306 (N_43306,N_36852,N_39846);
or U43307 (N_43307,N_37185,N_35896);
xor U43308 (N_43308,N_37540,N_37123);
xnor U43309 (N_43309,N_39640,N_37773);
nor U43310 (N_43310,N_36165,N_37391);
nand U43311 (N_43311,N_38350,N_38468);
nor U43312 (N_43312,N_36753,N_36253);
or U43313 (N_43313,N_37377,N_39751);
and U43314 (N_43314,N_37965,N_36681);
or U43315 (N_43315,N_39688,N_38401);
nor U43316 (N_43316,N_35236,N_36890);
nand U43317 (N_43317,N_37459,N_38696);
and U43318 (N_43318,N_37987,N_37752);
or U43319 (N_43319,N_39487,N_36065);
and U43320 (N_43320,N_38995,N_39049);
or U43321 (N_43321,N_36892,N_35819);
or U43322 (N_43322,N_38629,N_37019);
nor U43323 (N_43323,N_39936,N_37694);
or U43324 (N_43324,N_39603,N_37403);
nand U43325 (N_43325,N_39495,N_36882);
or U43326 (N_43326,N_35656,N_39273);
or U43327 (N_43327,N_35333,N_36213);
and U43328 (N_43328,N_36474,N_37539);
nand U43329 (N_43329,N_38693,N_39356);
xor U43330 (N_43330,N_38989,N_38856);
nand U43331 (N_43331,N_38463,N_39704);
nor U43332 (N_43332,N_36821,N_36613);
and U43333 (N_43333,N_35272,N_39578);
or U43334 (N_43334,N_37181,N_39687);
xnor U43335 (N_43335,N_35880,N_37126);
nand U43336 (N_43336,N_37579,N_37763);
nor U43337 (N_43337,N_36773,N_35032);
xnor U43338 (N_43338,N_37636,N_37308);
or U43339 (N_43339,N_37947,N_37752);
nor U43340 (N_43340,N_36956,N_37008);
and U43341 (N_43341,N_36608,N_39175);
and U43342 (N_43342,N_36719,N_39677);
xor U43343 (N_43343,N_39244,N_38269);
nor U43344 (N_43344,N_35430,N_37975);
nor U43345 (N_43345,N_39370,N_36246);
nor U43346 (N_43346,N_37671,N_39077);
nand U43347 (N_43347,N_35054,N_35422);
or U43348 (N_43348,N_39217,N_35143);
xor U43349 (N_43349,N_35507,N_36381);
nor U43350 (N_43350,N_36462,N_38376);
xnor U43351 (N_43351,N_39729,N_36053);
xnor U43352 (N_43352,N_35857,N_38573);
xnor U43353 (N_43353,N_38292,N_35608);
nor U43354 (N_43354,N_36373,N_37604);
nor U43355 (N_43355,N_35928,N_36245);
nand U43356 (N_43356,N_39432,N_35967);
and U43357 (N_43357,N_36271,N_39409);
nand U43358 (N_43358,N_36588,N_38428);
and U43359 (N_43359,N_35368,N_37835);
xnor U43360 (N_43360,N_38652,N_37174);
xor U43361 (N_43361,N_39136,N_38017);
and U43362 (N_43362,N_37656,N_38989);
or U43363 (N_43363,N_38435,N_38961);
and U43364 (N_43364,N_38754,N_39446);
or U43365 (N_43365,N_37282,N_36222);
xor U43366 (N_43366,N_37856,N_37116);
nand U43367 (N_43367,N_35429,N_36149);
or U43368 (N_43368,N_38034,N_39817);
or U43369 (N_43369,N_36421,N_36671);
nor U43370 (N_43370,N_36732,N_35571);
xor U43371 (N_43371,N_38219,N_36407);
nand U43372 (N_43372,N_35321,N_38650);
nor U43373 (N_43373,N_35624,N_35777);
nor U43374 (N_43374,N_39168,N_35582);
or U43375 (N_43375,N_35753,N_37080);
or U43376 (N_43376,N_39214,N_38828);
xor U43377 (N_43377,N_39947,N_38373);
xnor U43378 (N_43378,N_38985,N_35071);
and U43379 (N_43379,N_37574,N_35047);
or U43380 (N_43380,N_37813,N_36844);
and U43381 (N_43381,N_36646,N_39044);
and U43382 (N_43382,N_39391,N_37161);
nand U43383 (N_43383,N_37037,N_37191);
or U43384 (N_43384,N_38788,N_36189);
and U43385 (N_43385,N_39844,N_37204);
and U43386 (N_43386,N_38423,N_35009);
and U43387 (N_43387,N_38669,N_38371);
and U43388 (N_43388,N_36649,N_35300);
nor U43389 (N_43389,N_37026,N_38705);
xor U43390 (N_43390,N_38497,N_38909);
and U43391 (N_43391,N_35595,N_37106);
nand U43392 (N_43392,N_36295,N_39118);
and U43393 (N_43393,N_35334,N_37086);
xnor U43394 (N_43394,N_38810,N_39478);
nand U43395 (N_43395,N_39708,N_37113);
xor U43396 (N_43396,N_37149,N_38479);
and U43397 (N_43397,N_36792,N_37701);
and U43398 (N_43398,N_38549,N_36014);
nor U43399 (N_43399,N_37354,N_36026);
nor U43400 (N_43400,N_36236,N_38708);
xor U43401 (N_43401,N_36415,N_36165);
and U43402 (N_43402,N_36384,N_39558);
xnor U43403 (N_43403,N_36821,N_39088);
nand U43404 (N_43404,N_38404,N_36303);
nand U43405 (N_43405,N_38770,N_39108);
and U43406 (N_43406,N_36423,N_38259);
xor U43407 (N_43407,N_36281,N_37008);
or U43408 (N_43408,N_35457,N_38845);
xor U43409 (N_43409,N_38435,N_39219);
and U43410 (N_43410,N_36966,N_36463);
or U43411 (N_43411,N_36023,N_36175);
nand U43412 (N_43412,N_37107,N_39201);
nor U43413 (N_43413,N_39617,N_39370);
nor U43414 (N_43414,N_38465,N_38696);
nand U43415 (N_43415,N_39115,N_35855);
nand U43416 (N_43416,N_37917,N_39108);
xnor U43417 (N_43417,N_38873,N_36535);
or U43418 (N_43418,N_35885,N_38491);
xor U43419 (N_43419,N_36799,N_37482);
nor U43420 (N_43420,N_37084,N_36049);
nand U43421 (N_43421,N_38721,N_38683);
and U43422 (N_43422,N_37398,N_35278);
nor U43423 (N_43423,N_37397,N_35374);
xor U43424 (N_43424,N_38585,N_37322);
xor U43425 (N_43425,N_38338,N_37837);
nand U43426 (N_43426,N_37106,N_36232);
or U43427 (N_43427,N_37475,N_36692);
xor U43428 (N_43428,N_39422,N_36344);
nor U43429 (N_43429,N_37753,N_37710);
nand U43430 (N_43430,N_35504,N_37237);
and U43431 (N_43431,N_36021,N_35273);
xnor U43432 (N_43432,N_36475,N_37091);
nor U43433 (N_43433,N_36662,N_35613);
nand U43434 (N_43434,N_38044,N_38847);
xor U43435 (N_43435,N_37309,N_36515);
and U43436 (N_43436,N_36060,N_36819);
and U43437 (N_43437,N_38929,N_39152);
and U43438 (N_43438,N_38958,N_39600);
and U43439 (N_43439,N_36086,N_36678);
xnor U43440 (N_43440,N_39431,N_35401);
or U43441 (N_43441,N_39788,N_35868);
nand U43442 (N_43442,N_38107,N_37503);
xnor U43443 (N_43443,N_39670,N_38432);
nand U43444 (N_43444,N_37992,N_35501);
and U43445 (N_43445,N_37373,N_39239);
and U43446 (N_43446,N_37777,N_39453);
and U43447 (N_43447,N_39837,N_39687);
or U43448 (N_43448,N_39648,N_38754);
and U43449 (N_43449,N_37637,N_36334);
nor U43450 (N_43450,N_38396,N_37849);
nand U43451 (N_43451,N_36521,N_35419);
nor U43452 (N_43452,N_36465,N_38317);
nand U43453 (N_43453,N_37395,N_38771);
or U43454 (N_43454,N_37005,N_35909);
xnor U43455 (N_43455,N_38234,N_37225);
nand U43456 (N_43456,N_35731,N_38274);
xnor U43457 (N_43457,N_37362,N_38122);
nand U43458 (N_43458,N_36430,N_38912);
nand U43459 (N_43459,N_37195,N_39190);
xor U43460 (N_43460,N_38896,N_37244);
and U43461 (N_43461,N_39830,N_37160);
nand U43462 (N_43462,N_39083,N_37491);
or U43463 (N_43463,N_36121,N_37036);
xnor U43464 (N_43464,N_38621,N_36275);
or U43465 (N_43465,N_36338,N_35539);
and U43466 (N_43466,N_37769,N_38844);
and U43467 (N_43467,N_35594,N_39190);
xor U43468 (N_43468,N_37748,N_37616);
or U43469 (N_43469,N_39936,N_38397);
xnor U43470 (N_43470,N_37826,N_37454);
xnor U43471 (N_43471,N_38314,N_35545);
and U43472 (N_43472,N_37179,N_37010);
and U43473 (N_43473,N_39660,N_35996);
nand U43474 (N_43474,N_36763,N_38168);
and U43475 (N_43475,N_39350,N_39026);
xnor U43476 (N_43476,N_36603,N_35570);
nand U43477 (N_43477,N_39694,N_39657);
nor U43478 (N_43478,N_35467,N_35980);
nand U43479 (N_43479,N_36473,N_37681);
or U43480 (N_43480,N_39680,N_35486);
or U43481 (N_43481,N_39004,N_35604);
nor U43482 (N_43482,N_37773,N_38450);
nand U43483 (N_43483,N_37761,N_35554);
nand U43484 (N_43484,N_37055,N_38768);
xnor U43485 (N_43485,N_37551,N_38737);
nor U43486 (N_43486,N_35179,N_36586);
nand U43487 (N_43487,N_37714,N_35538);
and U43488 (N_43488,N_38893,N_37482);
xor U43489 (N_43489,N_36721,N_36934);
nand U43490 (N_43490,N_39351,N_38002);
nand U43491 (N_43491,N_39867,N_37808);
nand U43492 (N_43492,N_38901,N_38544);
xor U43493 (N_43493,N_36605,N_39049);
and U43494 (N_43494,N_38492,N_37645);
xor U43495 (N_43495,N_39838,N_35330);
nand U43496 (N_43496,N_39445,N_35421);
xor U43497 (N_43497,N_39619,N_39189);
nor U43498 (N_43498,N_36899,N_36970);
and U43499 (N_43499,N_39935,N_35127);
xnor U43500 (N_43500,N_39072,N_39529);
or U43501 (N_43501,N_38373,N_39740);
or U43502 (N_43502,N_37785,N_37029);
nand U43503 (N_43503,N_39594,N_38040);
and U43504 (N_43504,N_39279,N_38501);
xor U43505 (N_43505,N_38684,N_38519);
nand U43506 (N_43506,N_35559,N_39558);
nand U43507 (N_43507,N_38857,N_36623);
nor U43508 (N_43508,N_37014,N_38493);
nor U43509 (N_43509,N_36828,N_36605);
nand U43510 (N_43510,N_35043,N_35971);
nand U43511 (N_43511,N_37685,N_39524);
nand U43512 (N_43512,N_35348,N_38661);
or U43513 (N_43513,N_38339,N_39619);
nand U43514 (N_43514,N_35038,N_39820);
xor U43515 (N_43515,N_38032,N_35376);
nand U43516 (N_43516,N_38234,N_39633);
nor U43517 (N_43517,N_36098,N_38099);
xor U43518 (N_43518,N_37288,N_35345);
nor U43519 (N_43519,N_37319,N_37218);
nand U43520 (N_43520,N_37113,N_36460);
or U43521 (N_43521,N_35279,N_36794);
nor U43522 (N_43522,N_38918,N_35666);
nor U43523 (N_43523,N_37714,N_37357);
or U43524 (N_43524,N_38843,N_39462);
nand U43525 (N_43525,N_35706,N_39964);
nor U43526 (N_43526,N_36973,N_35054);
nor U43527 (N_43527,N_36571,N_37502);
xnor U43528 (N_43528,N_36383,N_35885);
xnor U43529 (N_43529,N_39722,N_35432);
or U43530 (N_43530,N_37060,N_35156);
nor U43531 (N_43531,N_37071,N_36889);
nor U43532 (N_43532,N_37231,N_35392);
nor U43533 (N_43533,N_35047,N_38655);
or U43534 (N_43534,N_37196,N_35019);
or U43535 (N_43535,N_36057,N_36288);
nand U43536 (N_43536,N_37086,N_36815);
or U43537 (N_43537,N_39528,N_38740);
and U43538 (N_43538,N_35051,N_35307);
or U43539 (N_43539,N_37476,N_39434);
xnor U43540 (N_43540,N_38782,N_38420);
nand U43541 (N_43541,N_36629,N_35192);
nand U43542 (N_43542,N_39485,N_37930);
nand U43543 (N_43543,N_35374,N_37717);
xor U43544 (N_43544,N_35719,N_35912);
or U43545 (N_43545,N_35827,N_37356);
nor U43546 (N_43546,N_37022,N_39641);
or U43547 (N_43547,N_36872,N_36421);
nand U43548 (N_43548,N_37190,N_38089);
and U43549 (N_43549,N_38574,N_37889);
and U43550 (N_43550,N_39842,N_37477);
nand U43551 (N_43551,N_39104,N_36640);
nor U43552 (N_43552,N_37361,N_36586);
and U43553 (N_43553,N_36325,N_36746);
nor U43554 (N_43554,N_35496,N_39049);
and U43555 (N_43555,N_36048,N_36265);
or U43556 (N_43556,N_38662,N_35513);
and U43557 (N_43557,N_35919,N_36705);
or U43558 (N_43558,N_36197,N_35917);
or U43559 (N_43559,N_36884,N_35607);
nand U43560 (N_43560,N_39274,N_36106);
xnor U43561 (N_43561,N_39625,N_37981);
nand U43562 (N_43562,N_37982,N_35362);
nand U43563 (N_43563,N_39306,N_38400);
or U43564 (N_43564,N_36830,N_37461);
or U43565 (N_43565,N_39925,N_37291);
nor U43566 (N_43566,N_37843,N_37141);
and U43567 (N_43567,N_35644,N_39053);
nor U43568 (N_43568,N_36385,N_36631);
nand U43569 (N_43569,N_35667,N_37831);
nor U43570 (N_43570,N_38074,N_35348);
nand U43571 (N_43571,N_36179,N_37947);
nor U43572 (N_43572,N_37630,N_37081);
nand U43573 (N_43573,N_36322,N_37587);
and U43574 (N_43574,N_37606,N_35730);
xnor U43575 (N_43575,N_38380,N_36561);
nor U43576 (N_43576,N_35254,N_39061);
nand U43577 (N_43577,N_36223,N_36884);
xor U43578 (N_43578,N_39737,N_38260);
xor U43579 (N_43579,N_36598,N_35062);
or U43580 (N_43580,N_36622,N_35831);
nor U43581 (N_43581,N_38818,N_37318);
xnor U43582 (N_43582,N_35770,N_39057);
nand U43583 (N_43583,N_38526,N_38547);
or U43584 (N_43584,N_36819,N_39924);
and U43585 (N_43585,N_36260,N_38675);
nand U43586 (N_43586,N_38715,N_37364);
and U43587 (N_43587,N_37244,N_39394);
nor U43588 (N_43588,N_35839,N_37682);
xor U43589 (N_43589,N_37984,N_37197);
and U43590 (N_43590,N_39504,N_39546);
or U43591 (N_43591,N_36479,N_36352);
nand U43592 (N_43592,N_38123,N_39472);
nor U43593 (N_43593,N_39405,N_39422);
nor U43594 (N_43594,N_39387,N_37660);
nor U43595 (N_43595,N_37866,N_39288);
and U43596 (N_43596,N_37132,N_39842);
xnor U43597 (N_43597,N_39730,N_37886);
xor U43598 (N_43598,N_37148,N_37032);
xnor U43599 (N_43599,N_38403,N_37998);
xor U43600 (N_43600,N_36887,N_38771);
xor U43601 (N_43601,N_37323,N_36014);
and U43602 (N_43602,N_39444,N_39973);
and U43603 (N_43603,N_39016,N_38062);
nand U43604 (N_43604,N_35189,N_35646);
nor U43605 (N_43605,N_39831,N_39222);
or U43606 (N_43606,N_37367,N_39796);
nor U43607 (N_43607,N_36135,N_35876);
nand U43608 (N_43608,N_39354,N_35163);
or U43609 (N_43609,N_36051,N_35062);
xor U43610 (N_43610,N_38860,N_36304);
nand U43611 (N_43611,N_36231,N_39773);
nand U43612 (N_43612,N_39863,N_36093);
xor U43613 (N_43613,N_39257,N_35522);
xnor U43614 (N_43614,N_39304,N_39739);
nor U43615 (N_43615,N_38383,N_35451);
nor U43616 (N_43616,N_38476,N_37590);
and U43617 (N_43617,N_39877,N_35016);
or U43618 (N_43618,N_39691,N_35502);
nand U43619 (N_43619,N_35861,N_38495);
nor U43620 (N_43620,N_37861,N_39197);
xor U43621 (N_43621,N_38281,N_37732);
and U43622 (N_43622,N_38655,N_36631);
nor U43623 (N_43623,N_37235,N_36396);
nor U43624 (N_43624,N_35270,N_39015);
xor U43625 (N_43625,N_35906,N_36443);
and U43626 (N_43626,N_37868,N_35613);
xnor U43627 (N_43627,N_35350,N_37056);
xor U43628 (N_43628,N_37607,N_35269);
or U43629 (N_43629,N_39875,N_39853);
or U43630 (N_43630,N_35514,N_38066);
or U43631 (N_43631,N_39249,N_39110);
nor U43632 (N_43632,N_39185,N_38268);
nand U43633 (N_43633,N_39887,N_35375);
or U43634 (N_43634,N_37980,N_36824);
and U43635 (N_43635,N_39426,N_36406);
nand U43636 (N_43636,N_38773,N_36608);
xnor U43637 (N_43637,N_36346,N_37397);
and U43638 (N_43638,N_39198,N_38115);
or U43639 (N_43639,N_35659,N_37704);
nor U43640 (N_43640,N_36086,N_35868);
or U43641 (N_43641,N_38547,N_39589);
or U43642 (N_43642,N_35352,N_37737);
nand U43643 (N_43643,N_38637,N_36991);
xor U43644 (N_43644,N_38136,N_39083);
nand U43645 (N_43645,N_37711,N_39185);
nor U43646 (N_43646,N_36950,N_37803);
nand U43647 (N_43647,N_38577,N_39934);
xnor U43648 (N_43648,N_39097,N_35605);
xnor U43649 (N_43649,N_39430,N_36215);
xnor U43650 (N_43650,N_39834,N_35698);
xnor U43651 (N_43651,N_36632,N_36521);
or U43652 (N_43652,N_39970,N_39234);
nor U43653 (N_43653,N_35039,N_36294);
nand U43654 (N_43654,N_36900,N_36723);
nor U43655 (N_43655,N_35387,N_36827);
and U43656 (N_43656,N_37558,N_38272);
nand U43657 (N_43657,N_39615,N_35004);
nand U43658 (N_43658,N_36874,N_36948);
or U43659 (N_43659,N_36128,N_37611);
or U43660 (N_43660,N_36528,N_35766);
xnor U43661 (N_43661,N_35234,N_38798);
nor U43662 (N_43662,N_37818,N_38002);
and U43663 (N_43663,N_35695,N_36141);
or U43664 (N_43664,N_38000,N_38748);
and U43665 (N_43665,N_37896,N_35455);
xor U43666 (N_43666,N_39462,N_39871);
nand U43667 (N_43667,N_36227,N_37229);
or U43668 (N_43668,N_35634,N_35196);
or U43669 (N_43669,N_39900,N_38778);
nand U43670 (N_43670,N_36932,N_35728);
and U43671 (N_43671,N_37095,N_39658);
nor U43672 (N_43672,N_37821,N_35272);
and U43673 (N_43673,N_37738,N_39916);
or U43674 (N_43674,N_35444,N_37874);
nand U43675 (N_43675,N_35486,N_35942);
nand U43676 (N_43676,N_36321,N_39881);
xnor U43677 (N_43677,N_35892,N_36912);
nor U43678 (N_43678,N_36424,N_35519);
nand U43679 (N_43679,N_36072,N_37803);
xnor U43680 (N_43680,N_35599,N_36027);
and U43681 (N_43681,N_38669,N_37941);
or U43682 (N_43682,N_37401,N_37188);
or U43683 (N_43683,N_39548,N_37170);
or U43684 (N_43684,N_39512,N_36354);
nor U43685 (N_43685,N_38618,N_38314);
or U43686 (N_43686,N_37175,N_38360);
xor U43687 (N_43687,N_39424,N_35648);
or U43688 (N_43688,N_39990,N_37964);
xnor U43689 (N_43689,N_35125,N_37513);
nand U43690 (N_43690,N_39099,N_36489);
and U43691 (N_43691,N_39676,N_38469);
nand U43692 (N_43692,N_37081,N_37263);
xnor U43693 (N_43693,N_38364,N_35756);
xor U43694 (N_43694,N_39384,N_35833);
xor U43695 (N_43695,N_38535,N_36061);
or U43696 (N_43696,N_39928,N_35666);
and U43697 (N_43697,N_35188,N_38497);
xnor U43698 (N_43698,N_35901,N_38720);
nor U43699 (N_43699,N_38260,N_39032);
nand U43700 (N_43700,N_38905,N_38849);
nor U43701 (N_43701,N_39206,N_38761);
xor U43702 (N_43702,N_39550,N_39732);
nor U43703 (N_43703,N_36022,N_38790);
nor U43704 (N_43704,N_39025,N_37445);
xnor U43705 (N_43705,N_37320,N_38411);
and U43706 (N_43706,N_38366,N_38811);
xnor U43707 (N_43707,N_38149,N_38881);
xnor U43708 (N_43708,N_38258,N_36834);
xor U43709 (N_43709,N_36277,N_35303);
nand U43710 (N_43710,N_38556,N_35287);
nand U43711 (N_43711,N_35210,N_35544);
or U43712 (N_43712,N_39018,N_39825);
xnor U43713 (N_43713,N_38702,N_35950);
xnor U43714 (N_43714,N_37939,N_38874);
xnor U43715 (N_43715,N_37793,N_36660);
nor U43716 (N_43716,N_35978,N_39319);
xnor U43717 (N_43717,N_39981,N_38322);
nor U43718 (N_43718,N_36874,N_39455);
or U43719 (N_43719,N_38408,N_37244);
and U43720 (N_43720,N_38863,N_37630);
nor U43721 (N_43721,N_36819,N_39501);
or U43722 (N_43722,N_39731,N_36740);
xnor U43723 (N_43723,N_38191,N_38883);
nor U43724 (N_43724,N_35241,N_36265);
xnor U43725 (N_43725,N_35489,N_39549);
nor U43726 (N_43726,N_35164,N_38853);
nand U43727 (N_43727,N_36185,N_38701);
nand U43728 (N_43728,N_35934,N_37499);
xor U43729 (N_43729,N_38483,N_36080);
xor U43730 (N_43730,N_37921,N_37641);
or U43731 (N_43731,N_38823,N_37600);
nor U43732 (N_43732,N_38187,N_37249);
nor U43733 (N_43733,N_35695,N_36814);
and U43734 (N_43734,N_35401,N_36513);
and U43735 (N_43735,N_36416,N_36047);
nor U43736 (N_43736,N_37577,N_39492);
nor U43737 (N_43737,N_37640,N_36954);
nand U43738 (N_43738,N_39053,N_35870);
nor U43739 (N_43739,N_38571,N_39758);
nor U43740 (N_43740,N_39939,N_37050);
nand U43741 (N_43741,N_36887,N_39258);
or U43742 (N_43742,N_35465,N_36675);
nand U43743 (N_43743,N_35224,N_35890);
and U43744 (N_43744,N_36042,N_38261);
xnor U43745 (N_43745,N_37526,N_38679);
and U43746 (N_43746,N_37073,N_36044);
and U43747 (N_43747,N_37151,N_36477);
nor U43748 (N_43748,N_35830,N_38582);
and U43749 (N_43749,N_39447,N_38542);
or U43750 (N_43750,N_39704,N_37603);
nand U43751 (N_43751,N_38608,N_35631);
xnor U43752 (N_43752,N_39667,N_38495);
xor U43753 (N_43753,N_35050,N_38673);
and U43754 (N_43754,N_35191,N_35275);
nor U43755 (N_43755,N_37729,N_36202);
nor U43756 (N_43756,N_37858,N_38879);
or U43757 (N_43757,N_39295,N_37119);
nand U43758 (N_43758,N_36465,N_38835);
or U43759 (N_43759,N_39245,N_36719);
and U43760 (N_43760,N_39196,N_39630);
and U43761 (N_43761,N_35859,N_36882);
and U43762 (N_43762,N_38688,N_38017);
nor U43763 (N_43763,N_35003,N_38725);
nor U43764 (N_43764,N_37285,N_38929);
and U43765 (N_43765,N_38665,N_39965);
xor U43766 (N_43766,N_37433,N_39532);
nand U43767 (N_43767,N_38834,N_39929);
and U43768 (N_43768,N_35722,N_39650);
nand U43769 (N_43769,N_39504,N_36040);
xnor U43770 (N_43770,N_35095,N_37644);
and U43771 (N_43771,N_35113,N_38467);
nand U43772 (N_43772,N_36872,N_38235);
nor U43773 (N_43773,N_38137,N_37330);
or U43774 (N_43774,N_36596,N_39197);
and U43775 (N_43775,N_36860,N_39605);
nand U43776 (N_43776,N_36620,N_38491);
xor U43777 (N_43777,N_36763,N_36814);
and U43778 (N_43778,N_38284,N_37115);
xnor U43779 (N_43779,N_35058,N_35683);
and U43780 (N_43780,N_39215,N_39570);
nor U43781 (N_43781,N_37979,N_38546);
nand U43782 (N_43782,N_38774,N_35499);
nor U43783 (N_43783,N_35791,N_36705);
nand U43784 (N_43784,N_36810,N_38409);
or U43785 (N_43785,N_38643,N_39367);
or U43786 (N_43786,N_38240,N_39947);
and U43787 (N_43787,N_36198,N_38456);
and U43788 (N_43788,N_35430,N_38806);
and U43789 (N_43789,N_35579,N_37104);
nand U43790 (N_43790,N_38123,N_36762);
and U43791 (N_43791,N_39822,N_36519);
and U43792 (N_43792,N_35412,N_38285);
and U43793 (N_43793,N_38266,N_38691);
and U43794 (N_43794,N_38178,N_36022);
nand U43795 (N_43795,N_36145,N_39663);
nor U43796 (N_43796,N_35142,N_38975);
nand U43797 (N_43797,N_39860,N_38821);
and U43798 (N_43798,N_36991,N_38306);
and U43799 (N_43799,N_38650,N_37853);
nand U43800 (N_43800,N_38527,N_35952);
nor U43801 (N_43801,N_38245,N_36734);
and U43802 (N_43802,N_38918,N_38418);
or U43803 (N_43803,N_38672,N_39444);
and U43804 (N_43804,N_39338,N_37657);
and U43805 (N_43805,N_37401,N_37165);
or U43806 (N_43806,N_38738,N_39316);
nor U43807 (N_43807,N_38486,N_38063);
or U43808 (N_43808,N_38030,N_37683);
xor U43809 (N_43809,N_38386,N_35939);
or U43810 (N_43810,N_39480,N_35478);
xnor U43811 (N_43811,N_36882,N_39779);
and U43812 (N_43812,N_38882,N_39749);
and U43813 (N_43813,N_36400,N_36099);
and U43814 (N_43814,N_38184,N_38593);
and U43815 (N_43815,N_39279,N_37188);
xor U43816 (N_43816,N_37416,N_38184);
xor U43817 (N_43817,N_36676,N_37237);
or U43818 (N_43818,N_35626,N_36773);
xnor U43819 (N_43819,N_38357,N_35712);
xnor U43820 (N_43820,N_39154,N_36163);
or U43821 (N_43821,N_37971,N_36366);
xor U43822 (N_43822,N_35692,N_37273);
and U43823 (N_43823,N_37035,N_39809);
and U43824 (N_43824,N_39317,N_36772);
and U43825 (N_43825,N_36995,N_37968);
or U43826 (N_43826,N_36746,N_39279);
and U43827 (N_43827,N_36065,N_36327);
xor U43828 (N_43828,N_37811,N_36122);
and U43829 (N_43829,N_36458,N_37713);
and U43830 (N_43830,N_39848,N_37362);
nor U43831 (N_43831,N_38594,N_35067);
xnor U43832 (N_43832,N_38924,N_38128);
and U43833 (N_43833,N_36072,N_35092);
xnor U43834 (N_43834,N_39408,N_36111);
xnor U43835 (N_43835,N_36004,N_39971);
or U43836 (N_43836,N_39521,N_38172);
or U43837 (N_43837,N_39114,N_36487);
xnor U43838 (N_43838,N_36808,N_35625);
nor U43839 (N_43839,N_38405,N_37562);
and U43840 (N_43840,N_38299,N_38433);
nor U43841 (N_43841,N_39878,N_39952);
nor U43842 (N_43842,N_37455,N_36117);
nor U43843 (N_43843,N_39728,N_37571);
nor U43844 (N_43844,N_36265,N_37125);
nand U43845 (N_43845,N_36071,N_39717);
and U43846 (N_43846,N_37364,N_37046);
nor U43847 (N_43847,N_35843,N_37747);
or U43848 (N_43848,N_39074,N_39517);
and U43849 (N_43849,N_38880,N_38695);
or U43850 (N_43850,N_37270,N_37053);
nor U43851 (N_43851,N_36043,N_35840);
or U43852 (N_43852,N_37853,N_37589);
xnor U43853 (N_43853,N_36119,N_35644);
nor U43854 (N_43854,N_36255,N_35087);
xor U43855 (N_43855,N_38025,N_35031);
and U43856 (N_43856,N_39467,N_37939);
nand U43857 (N_43857,N_38876,N_37569);
xor U43858 (N_43858,N_37105,N_37373);
nand U43859 (N_43859,N_37962,N_37038);
nor U43860 (N_43860,N_39098,N_38739);
nor U43861 (N_43861,N_39743,N_35592);
nand U43862 (N_43862,N_39656,N_39026);
or U43863 (N_43863,N_35664,N_37601);
and U43864 (N_43864,N_35733,N_38748);
nand U43865 (N_43865,N_37646,N_36874);
xor U43866 (N_43866,N_36189,N_35432);
nand U43867 (N_43867,N_36210,N_37548);
nand U43868 (N_43868,N_36488,N_39386);
or U43869 (N_43869,N_37765,N_36525);
nand U43870 (N_43870,N_36888,N_35539);
or U43871 (N_43871,N_37570,N_39245);
nor U43872 (N_43872,N_38758,N_37312);
nor U43873 (N_43873,N_37092,N_39203);
xnor U43874 (N_43874,N_35756,N_36012);
nor U43875 (N_43875,N_35796,N_39601);
nor U43876 (N_43876,N_37369,N_36833);
and U43877 (N_43877,N_38157,N_35067);
and U43878 (N_43878,N_36836,N_38610);
or U43879 (N_43879,N_35531,N_36621);
and U43880 (N_43880,N_38757,N_38523);
xnor U43881 (N_43881,N_37917,N_39269);
and U43882 (N_43882,N_38760,N_36810);
or U43883 (N_43883,N_38892,N_39894);
or U43884 (N_43884,N_37715,N_39971);
and U43885 (N_43885,N_36141,N_39929);
and U43886 (N_43886,N_37139,N_36696);
and U43887 (N_43887,N_36066,N_36063);
and U43888 (N_43888,N_38036,N_38208);
and U43889 (N_43889,N_36362,N_36595);
xor U43890 (N_43890,N_38349,N_35246);
or U43891 (N_43891,N_37577,N_39514);
xor U43892 (N_43892,N_39815,N_39784);
or U43893 (N_43893,N_37954,N_36193);
nand U43894 (N_43894,N_35254,N_38592);
nand U43895 (N_43895,N_39589,N_37372);
nor U43896 (N_43896,N_39980,N_36300);
nand U43897 (N_43897,N_35985,N_35095);
xor U43898 (N_43898,N_36788,N_37882);
and U43899 (N_43899,N_38029,N_36192);
nor U43900 (N_43900,N_37627,N_37952);
and U43901 (N_43901,N_36227,N_39859);
and U43902 (N_43902,N_37865,N_38103);
xor U43903 (N_43903,N_36580,N_35234);
xnor U43904 (N_43904,N_38777,N_35537);
and U43905 (N_43905,N_37086,N_38759);
xnor U43906 (N_43906,N_39360,N_37180);
nand U43907 (N_43907,N_38759,N_35780);
xnor U43908 (N_43908,N_37062,N_35049);
nand U43909 (N_43909,N_36807,N_39247);
xnor U43910 (N_43910,N_35679,N_39946);
or U43911 (N_43911,N_37915,N_39306);
nand U43912 (N_43912,N_36118,N_37499);
nor U43913 (N_43913,N_38696,N_35422);
and U43914 (N_43914,N_39964,N_39196);
and U43915 (N_43915,N_38747,N_38265);
xor U43916 (N_43916,N_36714,N_37221);
or U43917 (N_43917,N_36597,N_39271);
nor U43918 (N_43918,N_37955,N_38273);
nand U43919 (N_43919,N_38796,N_38439);
nor U43920 (N_43920,N_38580,N_38107);
nor U43921 (N_43921,N_39271,N_39379);
xnor U43922 (N_43922,N_36047,N_37524);
or U43923 (N_43923,N_39605,N_38985);
and U43924 (N_43924,N_35658,N_38981);
nor U43925 (N_43925,N_39528,N_36971);
nor U43926 (N_43926,N_39739,N_39451);
xnor U43927 (N_43927,N_36130,N_39993);
or U43928 (N_43928,N_35751,N_38779);
nor U43929 (N_43929,N_35351,N_39275);
xnor U43930 (N_43930,N_35388,N_36052);
xor U43931 (N_43931,N_35270,N_36848);
nor U43932 (N_43932,N_36058,N_36190);
xor U43933 (N_43933,N_38490,N_36025);
xor U43934 (N_43934,N_39016,N_39399);
and U43935 (N_43935,N_37615,N_35636);
nor U43936 (N_43936,N_38480,N_38738);
and U43937 (N_43937,N_37744,N_39501);
or U43938 (N_43938,N_37377,N_36697);
nand U43939 (N_43939,N_35260,N_35348);
nor U43940 (N_43940,N_38130,N_37013);
xnor U43941 (N_43941,N_39436,N_36141);
nand U43942 (N_43942,N_36417,N_39371);
nand U43943 (N_43943,N_35132,N_36932);
or U43944 (N_43944,N_38686,N_39084);
nor U43945 (N_43945,N_38985,N_38848);
xnor U43946 (N_43946,N_38156,N_35121);
nor U43947 (N_43947,N_39415,N_38185);
or U43948 (N_43948,N_36121,N_38208);
nor U43949 (N_43949,N_39037,N_37392);
xor U43950 (N_43950,N_37803,N_36298);
or U43951 (N_43951,N_38635,N_36917);
and U43952 (N_43952,N_35530,N_39148);
and U43953 (N_43953,N_38830,N_38985);
or U43954 (N_43954,N_38912,N_39968);
nor U43955 (N_43955,N_36267,N_37587);
nand U43956 (N_43956,N_39810,N_38236);
and U43957 (N_43957,N_38647,N_35842);
nand U43958 (N_43958,N_39884,N_36798);
and U43959 (N_43959,N_38096,N_36813);
and U43960 (N_43960,N_37933,N_35003);
xnor U43961 (N_43961,N_39553,N_37594);
nor U43962 (N_43962,N_36058,N_36590);
nor U43963 (N_43963,N_39472,N_39501);
and U43964 (N_43964,N_38859,N_39466);
nor U43965 (N_43965,N_38093,N_35142);
nor U43966 (N_43966,N_36037,N_38973);
nor U43967 (N_43967,N_39676,N_35241);
xor U43968 (N_43968,N_36084,N_39601);
nand U43969 (N_43969,N_35444,N_39677);
xor U43970 (N_43970,N_38714,N_36365);
xor U43971 (N_43971,N_37480,N_39253);
and U43972 (N_43972,N_37224,N_35389);
or U43973 (N_43973,N_35361,N_37650);
or U43974 (N_43974,N_35814,N_36010);
or U43975 (N_43975,N_39409,N_37599);
and U43976 (N_43976,N_38272,N_36394);
or U43977 (N_43977,N_36433,N_37643);
and U43978 (N_43978,N_35304,N_38406);
and U43979 (N_43979,N_36233,N_36940);
nand U43980 (N_43980,N_36486,N_35741);
nand U43981 (N_43981,N_38871,N_39585);
xnor U43982 (N_43982,N_39708,N_38951);
and U43983 (N_43983,N_39421,N_39217);
xor U43984 (N_43984,N_35934,N_36586);
and U43985 (N_43985,N_39936,N_39654);
nand U43986 (N_43986,N_37048,N_39386);
and U43987 (N_43987,N_38584,N_37127);
or U43988 (N_43988,N_39124,N_39953);
or U43989 (N_43989,N_39064,N_36277);
or U43990 (N_43990,N_36625,N_37852);
nand U43991 (N_43991,N_35949,N_39890);
nand U43992 (N_43992,N_38873,N_38425);
and U43993 (N_43993,N_38259,N_38358);
xnor U43994 (N_43994,N_35193,N_37481);
or U43995 (N_43995,N_38253,N_37737);
and U43996 (N_43996,N_35810,N_37831);
or U43997 (N_43997,N_36238,N_36260);
nand U43998 (N_43998,N_39443,N_37907);
xor U43999 (N_43999,N_39062,N_35189);
nor U44000 (N_44000,N_36671,N_39120);
nand U44001 (N_44001,N_36423,N_35887);
nand U44002 (N_44002,N_37336,N_39755);
or U44003 (N_44003,N_36320,N_39820);
xnor U44004 (N_44004,N_37573,N_39945);
nand U44005 (N_44005,N_38637,N_37056);
xor U44006 (N_44006,N_35807,N_37116);
xnor U44007 (N_44007,N_39086,N_37489);
xor U44008 (N_44008,N_35283,N_38605);
xnor U44009 (N_44009,N_38802,N_39711);
nand U44010 (N_44010,N_36653,N_36523);
or U44011 (N_44011,N_36914,N_38771);
or U44012 (N_44012,N_38082,N_35110);
nand U44013 (N_44013,N_39218,N_37623);
xor U44014 (N_44014,N_38021,N_39326);
nand U44015 (N_44015,N_35872,N_38974);
nand U44016 (N_44016,N_39507,N_35353);
nand U44017 (N_44017,N_35759,N_38738);
or U44018 (N_44018,N_36504,N_37653);
or U44019 (N_44019,N_39034,N_35995);
nand U44020 (N_44020,N_37088,N_39216);
and U44021 (N_44021,N_37841,N_35613);
nand U44022 (N_44022,N_35524,N_38534);
nand U44023 (N_44023,N_36838,N_35004);
and U44024 (N_44024,N_35199,N_35162);
nor U44025 (N_44025,N_36933,N_38742);
xnor U44026 (N_44026,N_36070,N_37539);
nand U44027 (N_44027,N_35949,N_35199);
or U44028 (N_44028,N_35175,N_36075);
nor U44029 (N_44029,N_39412,N_37094);
nor U44030 (N_44030,N_36543,N_38817);
nand U44031 (N_44031,N_38932,N_36612);
nor U44032 (N_44032,N_38059,N_37881);
xnor U44033 (N_44033,N_37130,N_39508);
or U44034 (N_44034,N_35522,N_39554);
xor U44035 (N_44035,N_39394,N_35422);
or U44036 (N_44036,N_39301,N_39659);
or U44037 (N_44037,N_38135,N_36380);
and U44038 (N_44038,N_37629,N_39500);
xor U44039 (N_44039,N_38202,N_38207);
or U44040 (N_44040,N_39280,N_38012);
xnor U44041 (N_44041,N_35081,N_38268);
xnor U44042 (N_44042,N_35657,N_35980);
or U44043 (N_44043,N_36008,N_36259);
nand U44044 (N_44044,N_36199,N_38525);
xnor U44045 (N_44045,N_37335,N_36041);
and U44046 (N_44046,N_39870,N_35298);
and U44047 (N_44047,N_39358,N_36014);
nand U44048 (N_44048,N_37063,N_39048);
or U44049 (N_44049,N_36258,N_36658);
or U44050 (N_44050,N_37227,N_37153);
or U44051 (N_44051,N_35595,N_35648);
and U44052 (N_44052,N_39966,N_37684);
or U44053 (N_44053,N_39171,N_39371);
xor U44054 (N_44054,N_39750,N_35947);
nor U44055 (N_44055,N_36047,N_36588);
xnor U44056 (N_44056,N_36562,N_39511);
nor U44057 (N_44057,N_36304,N_36287);
or U44058 (N_44058,N_37255,N_36665);
and U44059 (N_44059,N_38608,N_38763);
or U44060 (N_44060,N_37600,N_36382);
and U44061 (N_44061,N_35967,N_37012);
nor U44062 (N_44062,N_37339,N_37950);
and U44063 (N_44063,N_35573,N_39632);
nor U44064 (N_44064,N_36941,N_38404);
nand U44065 (N_44065,N_37224,N_35131);
and U44066 (N_44066,N_36954,N_38588);
or U44067 (N_44067,N_37274,N_35903);
xnor U44068 (N_44068,N_37706,N_36815);
nand U44069 (N_44069,N_36595,N_36026);
or U44070 (N_44070,N_36485,N_38632);
nand U44071 (N_44071,N_39988,N_35373);
nor U44072 (N_44072,N_39408,N_39620);
xnor U44073 (N_44073,N_37725,N_35395);
or U44074 (N_44074,N_37127,N_38612);
xnor U44075 (N_44075,N_35672,N_39800);
and U44076 (N_44076,N_35461,N_39586);
and U44077 (N_44077,N_36110,N_39280);
or U44078 (N_44078,N_36632,N_39515);
and U44079 (N_44079,N_36421,N_38449);
and U44080 (N_44080,N_37802,N_37589);
or U44081 (N_44081,N_35721,N_36597);
nor U44082 (N_44082,N_39134,N_38927);
xor U44083 (N_44083,N_36749,N_35317);
nor U44084 (N_44084,N_36480,N_36897);
nand U44085 (N_44085,N_35135,N_35438);
xor U44086 (N_44086,N_38214,N_38038);
nand U44087 (N_44087,N_39790,N_35120);
or U44088 (N_44088,N_36603,N_37371);
or U44089 (N_44089,N_36143,N_37051);
nand U44090 (N_44090,N_39523,N_36649);
xor U44091 (N_44091,N_39028,N_38632);
and U44092 (N_44092,N_37518,N_36591);
nor U44093 (N_44093,N_38468,N_38598);
and U44094 (N_44094,N_38211,N_38264);
nand U44095 (N_44095,N_37439,N_38472);
nand U44096 (N_44096,N_35470,N_39660);
nor U44097 (N_44097,N_37579,N_36293);
nor U44098 (N_44098,N_37167,N_37493);
and U44099 (N_44099,N_35822,N_35366);
nor U44100 (N_44100,N_35437,N_38974);
nor U44101 (N_44101,N_38516,N_38445);
nor U44102 (N_44102,N_35208,N_36680);
nor U44103 (N_44103,N_38741,N_38599);
xnor U44104 (N_44104,N_38286,N_38543);
or U44105 (N_44105,N_39439,N_37452);
or U44106 (N_44106,N_37113,N_39409);
nor U44107 (N_44107,N_38245,N_37715);
and U44108 (N_44108,N_35588,N_36263);
or U44109 (N_44109,N_35060,N_36171);
xnor U44110 (N_44110,N_36298,N_39185);
nor U44111 (N_44111,N_35102,N_39012);
and U44112 (N_44112,N_38739,N_36969);
or U44113 (N_44113,N_38167,N_38696);
nand U44114 (N_44114,N_35010,N_37970);
nor U44115 (N_44115,N_35377,N_36205);
nor U44116 (N_44116,N_38802,N_36955);
and U44117 (N_44117,N_35309,N_39659);
nor U44118 (N_44118,N_37692,N_35197);
xor U44119 (N_44119,N_38126,N_39126);
nor U44120 (N_44120,N_38043,N_38122);
and U44121 (N_44121,N_36000,N_38130);
or U44122 (N_44122,N_38135,N_36859);
nand U44123 (N_44123,N_38663,N_36318);
nand U44124 (N_44124,N_39109,N_37846);
or U44125 (N_44125,N_38787,N_39687);
nand U44126 (N_44126,N_38443,N_39296);
and U44127 (N_44127,N_38841,N_39912);
xnor U44128 (N_44128,N_38080,N_39842);
and U44129 (N_44129,N_35693,N_38177);
nand U44130 (N_44130,N_36863,N_39905);
or U44131 (N_44131,N_39340,N_37546);
and U44132 (N_44132,N_36844,N_39234);
nand U44133 (N_44133,N_37050,N_36471);
and U44134 (N_44134,N_39808,N_35070);
and U44135 (N_44135,N_38770,N_35797);
or U44136 (N_44136,N_38802,N_35875);
nand U44137 (N_44137,N_38581,N_38501);
and U44138 (N_44138,N_39526,N_37886);
or U44139 (N_44139,N_38192,N_36648);
nor U44140 (N_44140,N_35836,N_39836);
or U44141 (N_44141,N_37579,N_39368);
nand U44142 (N_44142,N_38657,N_36299);
xnor U44143 (N_44143,N_36778,N_35763);
nor U44144 (N_44144,N_36410,N_38791);
xor U44145 (N_44145,N_39837,N_39705);
and U44146 (N_44146,N_39605,N_39932);
and U44147 (N_44147,N_35900,N_36116);
nor U44148 (N_44148,N_36392,N_39146);
or U44149 (N_44149,N_39559,N_36961);
nor U44150 (N_44150,N_39029,N_38034);
and U44151 (N_44151,N_36529,N_35523);
or U44152 (N_44152,N_38426,N_37684);
and U44153 (N_44153,N_35090,N_37922);
and U44154 (N_44154,N_39447,N_35775);
nor U44155 (N_44155,N_35121,N_37907);
xor U44156 (N_44156,N_37063,N_37725);
nand U44157 (N_44157,N_36389,N_38768);
and U44158 (N_44158,N_36687,N_37147);
nand U44159 (N_44159,N_37453,N_36585);
nor U44160 (N_44160,N_36774,N_39189);
and U44161 (N_44161,N_35971,N_37379);
and U44162 (N_44162,N_38550,N_39624);
xnor U44163 (N_44163,N_39849,N_38353);
xnor U44164 (N_44164,N_39414,N_37888);
nor U44165 (N_44165,N_39230,N_38967);
nor U44166 (N_44166,N_39443,N_37811);
or U44167 (N_44167,N_39099,N_38090);
and U44168 (N_44168,N_37379,N_36469);
xnor U44169 (N_44169,N_36107,N_38778);
or U44170 (N_44170,N_35744,N_36611);
xor U44171 (N_44171,N_38531,N_37533);
nand U44172 (N_44172,N_38505,N_35634);
xor U44173 (N_44173,N_39411,N_37941);
nand U44174 (N_44174,N_35790,N_39450);
nor U44175 (N_44175,N_37500,N_36409);
xor U44176 (N_44176,N_36828,N_35417);
nor U44177 (N_44177,N_37331,N_35424);
nor U44178 (N_44178,N_38425,N_36245);
xnor U44179 (N_44179,N_37652,N_37816);
xnor U44180 (N_44180,N_35174,N_35577);
xnor U44181 (N_44181,N_37025,N_39804);
or U44182 (N_44182,N_36665,N_36309);
or U44183 (N_44183,N_39557,N_37695);
or U44184 (N_44184,N_36511,N_39090);
xor U44185 (N_44185,N_35705,N_36976);
and U44186 (N_44186,N_39002,N_38239);
nor U44187 (N_44187,N_39319,N_36916);
and U44188 (N_44188,N_36520,N_37206);
xnor U44189 (N_44189,N_39933,N_37063);
nand U44190 (N_44190,N_39631,N_39600);
nand U44191 (N_44191,N_37589,N_35566);
and U44192 (N_44192,N_38417,N_35620);
nor U44193 (N_44193,N_39826,N_37217);
nand U44194 (N_44194,N_35237,N_39711);
and U44195 (N_44195,N_36696,N_39385);
nand U44196 (N_44196,N_37949,N_36848);
nor U44197 (N_44197,N_38963,N_36110);
nor U44198 (N_44198,N_36079,N_39481);
or U44199 (N_44199,N_39339,N_39752);
xnor U44200 (N_44200,N_39516,N_35836);
nor U44201 (N_44201,N_38559,N_37384);
or U44202 (N_44202,N_37441,N_36768);
or U44203 (N_44203,N_39603,N_35173);
nand U44204 (N_44204,N_39111,N_37239);
xnor U44205 (N_44205,N_38827,N_38845);
nand U44206 (N_44206,N_37353,N_38865);
or U44207 (N_44207,N_37611,N_38523);
xor U44208 (N_44208,N_39339,N_39228);
nand U44209 (N_44209,N_39185,N_39339);
xnor U44210 (N_44210,N_35374,N_39757);
or U44211 (N_44211,N_39712,N_36811);
and U44212 (N_44212,N_35150,N_37772);
or U44213 (N_44213,N_38876,N_38854);
or U44214 (N_44214,N_37472,N_39673);
or U44215 (N_44215,N_35561,N_39204);
xnor U44216 (N_44216,N_39671,N_36371);
nand U44217 (N_44217,N_35463,N_36628);
or U44218 (N_44218,N_35926,N_39675);
or U44219 (N_44219,N_39001,N_38590);
xnor U44220 (N_44220,N_36745,N_39093);
nand U44221 (N_44221,N_35273,N_39780);
nor U44222 (N_44222,N_37107,N_35014);
and U44223 (N_44223,N_37350,N_36259);
nor U44224 (N_44224,N_37170,N_36019);
nand U44225 (N_44225,N_39595,N_35707);
nand U44226 (N_44226,N_37761,N_35382);
and U44227 (N_44227,N_35175,N_37433);
nor U44228 (N_44228,N_36618,N_38667);
xnor U44229 (N_44229,N_37522,N_38561);
or U44230 (N_44230,N_35711,N_38940);
nor U44231 (N_44231,N_35700,N_38723);
nor U44232 (N_44232,N_37681,N_37323);
or U44233 (N_44233,N_35926,N_39715);
and U44234 (N_44234,N_35217,N_39209);
nand U44235 (N_44235,N_39642,N_38424);
nor U44236 (N_44236,N_39667,N_35221);
or U44237 (N_44237,N_36949,N_36419);
nand U44238 (N_44238,N_37464,N_36143);
or U44239 (N_44239,N_38947,N_39057);
and U44240 (N_44240,N_37822,N_39596);
nand U44241 (N_44241,N_38867,N_36860);
or U44242 (N_44242,N_37096,N_37778);
xor U44243 (N_44243,N_37788,N_37167);
xnor U44244 (N_44244,N_36623,N_38970);
nor U44245 (N_44245,N_38283,N_37462);
nand U44246 (N_44246,N_38121,N_39694);
xor U44247 (N_44247,N_38687,N_37391);
xor U44248 (N_44248,N_37742,N_37930);
xnor U44249 (N_44249,N_37208,N_36466);
or U44250 (N_44250,N_35018,N_38324);
and U44251 (N_44251,N_36263,N_38796);
and U44252 (N_44252,N_38374,N_36173);
or U44253 (N_44253,N_35777,N_36513);
and U44254 (N_44254,N_35334,N_37670);
nand U44255 (N_44255,N_37227,N_35771);
nand U44256 (N_44256,N_39739,N_36937);
nor U44257 (N_44257,N_37172,N_38667);
or U44258 (N_44258,N_35453,N_37907);
nor U44259 (N_44259,N_35822,N_38758);
nand U44260 (N_44260,N_38931,N_38526);
xor U44261 (N_44261,N_38137,N_37564);
nor U44262 (N_44262,N_37131,N_38496);
or U44263 (N_44263,N_37803,N_37289);
nand U44264 (N_44264,N_35259,N_39021);
nor U44265 (N_44265,N_36099,N_39774);
nand U44266 (N_44266,N_37824,N_38142);
xor U44267 (N_44267,N_37692,N_37520);
nor U44268 (N_44268,N_36471,N_39065);
and U44269 (N_44269,N_37691,N_35287);
or U44270 (N_44270,N_38910,N_37416);
nor U44271 (N_44271,N_36561,N_35194);
nand U44272 (N_44272,N_39778,N_35005);
or U44273 (N_44273,N_39610,N_38345);
and U44274 (N_44274,N_36502,N_37783);
xnor U44275 (N_44275,N_38886,N_39703);
nor U44276 (N_44276,N_38398,N_37656);
xnor U44277 (N_44277,N_35073,N_35651);
nor U44278 (N_44278,N_39427,N_37703);
nor U44279 (N_44279,N_39988,N_37357);
or U44280 (N_44280,N_37171,N_35871);
and U44281 (N_44281,N_39767,N_38514);
nor U44282 (N_44282,N_38797,N_38600);
xor U44283 (N_44283,N_38207,N_35366);
or U44284 (N_44284,N_36570,N_39784);
nand U44285 (N_44285,N_39319,N_37155);
nor U44286 (N_44286,N_35275,N_37854);
xor U44287 (N_44287,N_37851,N_36371);
xnor U44288 (N_44288,N_38156,N_35007);
or U44289 (N_44289,N_38733,N_36092);
xor U44290 (N_44290,N_38861,N_39544);
or U44291 (N_44291,N_39980,N_38419);
xor U44292 (N_44292,N_37486,N_36443);
xor U44293 (N_44293,N_39636,N_36194);
xor U44294 (N_44294,N_35304,N_36575);
nor U44295 (N_44295,N_37142,N_35185);
nor U44296 (N_44296,N_37364,N_35089);
or U44297 (N_44297,N_35642,N_37049);
nand U44298 (N_44298,N_36596,N_35930);
or U44299 (N_44299,N_35190,N_39534);
and U44300 (N_44300,N_36070,N_38195);
nand U44301 (N_44301,N_37451,N_38305);
or U44302 (N_44302,N_35622,N_39024);
nor U44303 (N_44303,N_35561,N_39646);
or U44304 (N_44304,N_37481,N_39136);
xor U44305 (N_44305,N_38824,N_39848);
xor U44306 (N_44306,N_38627,N_37449);
xor U44307 (N_44307,N_37241,N_36832);
nor U44308 (N_44308,N_36514,N_38840);
and U44309 (N_44309,N_38260,N_39188);
nand U44310 (N_44310,N_37618,N_36218);
nand U44311 (N_44311,N_38622,N_39702);
nand U44312 (N_44312,N_36545,N_37412);
xnor U44313 (N_44313,N_36287,N_37889);
or U44314 (N_44314,N_35075,N_38518);
nor U44315 (N_44315,N_38477,N_37056);
or U44316 (N_44316,N_35757,N_35264);
xnor U44317 (N_44317,N_39963,N_36301);
xor U44318 (N_44318,N_37572,N_39787);
xnor U44319 (N_44319,N_37656,N_37632);
or U44320 (N_44320,N_37070,N_39009);
nor U44321 (N_44321,N_38748,N_39273);
xor U44322 (N_44322,N_36245,N_39573);
or U44323 (N_44323,N_36874,N_37920);
nor U44324 (N_44324,N_35279,N_38410);
nor U44325 (N_44325,N_38107,N_36375);
and U44326 (N_44326,N_39540,N_35718);
xor U44327 (N_44327,N_35156,N_39572);
nand U44328 (N_44328,N_38032,N_36206);
or U44329 (N_44329,N_36842,N_37415);
xnor U44330 (N_44330,N_36150,N_37109);
and U44331 (N_44331,N_39785,N_37337);
or U44332 (N_44332,N_36418,N_38781);
nand U44333 (N_44333,N_37335,N_39098);
nand U44334 (N_44334,N_36697,N_36472);
nand U44335 (N_44335,N_36090,N_37344);
or U44336 (N_44336,N_38168,N_35326);
or U44337 (N_44337,N_36568,N_35137);
and U44338 (N_44338,N_39299,N_36006);
nand U44339 (N_44339,N_39937,N_38256);
and U44340 (N_44340,N_39540,N_38546);
xor U44341 (N_44341,N_37909,N_37308);
and U44342 (N_44342,N_39664,N_38919);
nor U44343 (N_44343,N_39883,N_37185);
and U44344 (N_44344,N_38778,N_37870);
xor U44345 (N_44345,N_36498,N_35694);
xor U44346 (N_44346,N_36346,N_38622);
nor U44347 (N_44347,N_38734,N_37052);
nor U44348 (N_44348,N_36961,N_39981);
xor U44349 (N_44349,N_37759,N_35716);
or U44350 (N_44350,N_36664,N_35257);
or U44351 (N_44351,N_35902,N_39246);
xnor U44352 (N_44352,N_35712,N_38401);
xnor U44353 (N_44353,N_37646,N_35466);
nor U44354 (N_44354,N_36259,N_39088);
or U44355 (N_44355,N_38759,N_39705);
nand U44356 (N_44356,N_39134,N_36722);
and U44357 (N_44357,N_36005,N_36504);
nand U44358 (N_44358,N_36761,N_39633);
or U44359 (N_44359,N_37865,N_36876);
nor U44360 (N_44360,N_35521,N_36182);
nor U44361 (N_44361,N_39111,N_37799);
nor U44362 (N_44362,N_39755,N_35212);
nor U44363 (N_44363,N_39173,N_35996);
nor U44364 (N_44364,N_37944,N_36834);
nor U44365 (N_44365,N_36673,N_36594);
and U44366 (N_44366,N_38866,N_37317);
or U44367 (N_44367,N_35237,N_38146);
nor U44368 (N_44368,N_37044,N_38653);
or U44369 (N_44369,N_37198,N_35329);
or U44370 (N_44370,N_37302,N_36202);
nor U44371 (N_44371,N_38841,N_39030);
xor U44372 (N_44372,N_39331,N_36410);
or U44373 (N_44373,N_37756,N_39629);
and U44374 (N_44374,N_39349,N_37133);
xor U44375 (N_44375,N_37034,N_38240);
nand U44376 (N_44376,N_38888,N_39948);
nand U44377 (N_44377,N_37594,N_36517);
xnor U44378 (N_44378,N_37657,N_36435);
nor U44379 (N_44379,N_39889,N_36090);
nor U44380 (N_44380,N_35866,N_37118);
xor U44381 (N_44381,N_35222,N_36052);
or U44382 (N_44382,N_38878,N_39608);
and U44383 (N_44383,N_39025,N_37867);
nor U44384 (N_44384,N_35695,N_39860);
or U44385 (N_44385,N_36180,N_38408);
nor U44386 (N_44386,N_37383,N_36652);
nor U44387 (N_44387,N_39661,N_38633);
nor U44388 (N_44388,N_38769,N_38523);
or U44389 (N_44389,N_35139,N_35779);
and U44390 (N_44390,N_36694,N_35909);
or U44391 (N_44391,N_39636,N_35925);
or U44392 (N_44392,N_39122,N_38135);
nor U44393 (N_44393,N_38630,N_37966);
nor U44394 (N_44394,N_38302,N_38766);
nor U44395 (N_44395,N_39491,N_35213);
and U44396 (N_44396,N_36233,N_36777);
nand U44397 (N_44397,N_37246,N_36831);
nor U44398 (N_44398,N_35966,N_37699);
or U44399 (N_44399,N_39529,N_38644);
nand U44400 (N_44400,N_38635,N_38164);
xor U44401 (N_44401,N_35361,N_39753);
nand U44402 (N_44402,N_39608,N_38846);
xnor U44403 (N_44403,N_39454,N_36204);
xor U44404 (N_44404,N_38253,N_36140);
nor U44405 (N_44405,N_35802,N_39401);
and U44406 (N_44406,N_36239,N_38348);
nand U44407 (N_44407,N_38119,N_35843);
nand U44408 (N_44408,N_37768,N_39897);
or U44409 (N_44409,N_37321,N_37070);
nand U44410 (N_44410,N_35255,N_39282);
and U44411 (N_44411,N_39782,N_36721);
or U44412 (N_44412,N_39442,N_35766);
nor U44413 (N_44413,N_35677,N_36085);
nand U44414 (N_44414,N_39930,N_37224);
and U44415 (N_44415,N_39915,N_35269);
xor U44416 (N_44416,N_38720,N_38532);
xnor U44417 (N_44417,N_35693,N_36990);
xor U44418 (N_44418,N_36366,N_39755);
xnor U44419 (N_44419,N_36621,N_35117);
and U44420 (N_44420,N_38524,N_38319);
and U44421 (N_44421,N_36332,N_35990);
nand U44422 (N_44422,N_39778,N_36263);
and U44423 (N_44423,N_38089,N_35161);
or U44424 (N_44424,N_38223,N_37097);
xor U44425 (N_44425,N_39530,N_38997);
or U44426 (N_44426,N_39563,N_39557);
or U44427 (N_44427,N_39604,N_35574);
xnor U44428 (N_44428,N_35433,N_38738);
xor U44429 (N_44429,N_38971,N_36161);
nand U44430 (N_44430,N_39804,N_37467);
and U44431 (N_44431,N_38481,N_38853);
nor U44432 (N_44432,N_36229,N_36312);
or U44433 (N_44433,N_35731,N_37723);
or U44434 (N_44434,N_36703,N_38194);
nand U44435 (N_44435,N_39015,N_36852);
xor U44436 (N_44436,N_37831,N_37217);
or U44437 (N_44437,N_36400,N_38198);
and U44438 (N_44438,N_38122,N_36282);
nor U44439 (N_44439,N_39722,N_39550);
xor U44440 (N_44440,N_36303,N_38114);
and U44441 (N_44441,N_38123,N_39536);
xor U44442 (N_44442,N_38802,N_38906);
xor U44443 (N_44443,N_36267,N_38606);
and U44444 (N_44444,N_35116,N_39954);
and U44445 (N_44445,N_36358,N_39084);
nand U44446 (N_44446,N_38726,N_37845);
or U44447 (N_44447,N_35255,N_35287);
or U44448 (N_44448,N_36714,N_36547);
nand U44449 (N_44449,N_37494,N_38690);
and U44450 (N_44450,N_38185,N_38784);
xor U44451 (N_44451,N_39183,N_37997);
nand U44452 (N_44452,N_39381,N_35601);
and U44453 (N_44453,N_38842,N_35675);
and U44454 (N_44454,N_38403,N_39931);
and U44455 (N_44455,N_39324,N_35230);
or U44456 (N_44456,N_37047,N_37942);
or U44457 (N_44457,N_38845,N_36337);
xnor U44458 (N_44458,N_38368,N_38716);
or U44459 (N_44459,N_36144,N_38250);
or U44460 (N_44460,N_39633,N_37674);
and U44461 (N_44461,N_36439,N_35993);
nor U44462 (N_44462,N_37766,N_35198);
nand U44463 (N_44463,N_39529,N_37905);
or U44464 (N_44464,N_36249,N_39333);
nand U44465 (N_44465,N_36529,N_37685);
xnor U44466 (N_44466,N_38591,N_36558);
xor U44467 (N_44467,N_38191,N_39857);
xor U44468 (N_44468,N_39161,N_36466);
nor U44469 (N_44469,N_37284,N_38104);
or U44470 (N_44470,N_39543,N_35105);
nand U44471 (N_44471,N_39031,N_37168);
or U44472 (N_44472,N_35418,N_38986);
or U44473 (N_44473,N_35440,N_37110);
nand U44474 (N_44474,N_35870,N_36601);
xnor U44475 (N_44475,N_37727,N_38041);
and U44476 (N_44476,N_36773,N_36850);
or U44477 (N_44477,N_37374,N_36637);
nand U44478 (N_44478,N_35686,N_35560);
or U44479 (N_44479,N_38133,N_39382);
or U44480 (N_44480,N_35437,N_39042);
and U44481 (N_44481,N_38193,N_37769);
xor U44482 (N_44482,N_38471,N_37125);
or U44483 (N_44483,N_37931,N_39863);
xnor U44484 (N_44484,N_38818,N_37150);
or U44485 (N_44485,N_35758,N_38254);
and U44486 (N_44486,N_38926,N_37651);
and U44487 (N_44487,N_38694,N_36081);
nand U44488 (N_44488,N_38683,N_38221);
nor U44489 (N_44489,N_38373,N_37418);
xor U44490 (N_44490,N_36868,N_37630);
and U44491 (N_44491,N_36232,N_35553);
or U44492 (N_44492,N_39633,N_38439);
or U44493 (N_44493,N_35965,N_35051);
or U44494 (N_44494,N_38945,N_38624);
and U44495 (N_44495,N_35856,N_37120);
or U44496 (N_44496,N_36032,N_37758);
or U44497 (N_44497,N_36440,N_36657);
nand U44498 (N_44498,N_39573,N_35776);
nor U44499 (N_44499,N_39756,N_38318);
xnor U44500 (N_44500,N_35788,N_37368);
nand U44501 (N_44501,N_39237,N_36233);
nor U44502 (N_44502,N_36536,N_39933);
xor U44503 (N_44503,N_35705,N_38830);
nor U44504 (N_44504,N_36840,N_36217);
nor U44505 (N_44505,N_35572,N_38458);
xor U44506 (N_44506,N_38115,N_35178);
xnor U44507 (N_44507,N_35682,N_36440);
nand U44508 (N_44508,N_36093,N_37483);
or U44509 (N_44509,N_36670,N_37169);
xnor U44510 (N_44510,N_35853,N_38540);
xnor U44511 (N_44511,N_36561,N_35843);
nand U44512 (N_44512,N_38106,N_38160);
and U44513 (N_44513,N_39861,N_37869);
and U44514 (N_44514,N_39748,N_39270);
or U44515 (N_44515,N_37084,N_35174);
and U44516 (N_44516,N_38155,N_39910);
or U44517 (N_44517,N_38604,N_36856);
and U44518 (N_44518,N_39055,N_37465);
nand U44519 (N_44519,N_38360,N_36672);
nor U44520 (N_44520,N_37442,N_36102);
nor U44521 (N_44521,N_36301,N_35460);
nand U44522 (N_44522,N_37990,N_38598);
nand U44523 (N_44523,N_39875,N_39175);
and U44524 (N_44524,N_36528,N_39328);
nand U44525 (N_44525,N_39580,N_36495);
and U44526 (N_44526,N_35954,N_38809);
or U44527 (N_44527,N_35641,N_35000);
or U44528 (N_44528,N_39708,N_36998);
nand U44529 (N_44529,N_37022,N_35867);
nor U44530 (N_44530,N_36463,N_37539);
and U44531 (N_44531,N_37301,N_39653);
and U44532 (N_44532,N_37240,N_39572);
or U44533 (N_44533,N_38547,N_39453);
or U44534 (N_44534,N_35019,N_37825);
and U44535 (N_44535,N_36855,N_36447);
nand U44536 (N_44536,N_36034,N_36088);
nor U44537 (N_44537,N_35112,N_35823);
nand U44538 (N_44538,N_39711,N_37602);
nor U44539 (N_44539,N_37603,N_35816);
nor U44540 (N_44540,N_35935,N_36015);
or U44541 (N_44541,N_36175,N_39727);
xnor U44542 (N_44542,N_36858,N_36135);
nor U44543 (N_44543,N_35549,N_37262);
nor U44544 (N_44544,N_36967,N_39524);
and U44545 (N_44545,N_37820,N_38056);
or U44546 (N_44546,N_38581,N_36474);
or U44547 (N_44547,N_35030,N_39056);
and U44548 (N_44548,N_36359,N_36798);
nor U44549 (N_44549,N_36082,N_39567);
or U44550 (N_44550,N_37296,N_39408);
xnor U44551 (N_44551,N_36702,N_36413);
or U44552 (N_44552,N_37621,N_36541);
nand U44553 (N_44553,N_37541,N_35416);
or U44554 (N_44554,N_37830,N_38542);
or U44555 (N_44555,N_36725,N_38729);
or U44556 (N_44556,N_37371,N_35658);
xor U44557 (N_44557,N_37093,N_35028);
nand U44558 (N_44558,N_35979,N_35668);
nand U44559 (N_44559,N_39102,N_39083);
or U44560 (N_44560,N_37633,N_35125);
xor U44561 (N_44561,N_39805,N_39167);
nor U44562 (N_44562,N_38243,N_36112);
and U44563 (N_44563,N_35173,N_36124);
xnor U44564 (N_44564,N_38247,N_35586);
xor U44565 (N_44565,N_37426,N_35193);
and U44566 (N_44566,N_39435,N_39965);
nand U44567 (N_44567,N_38400,N_38615);
nor U44568 (N_44568,N_38749,N_37267);
nor U44569 (N_44569,N_38796,N_37636);
and U44570 (N_44570,N_36249,N_38965);
nor U44571 (N_44571,N_39936,N_35757);
nor U44572 (N_44572,N_36832,N_36431);
or U44573 (N_44573,N_36239,N_35446);
nor U44574 (N_44574,N_35797,N_35988);
nor U44575 (N_44575,N_36914,N_38204);
and U44576 (N_44576,N_35939,N_35993);
or U44577 (N_44577,N_39356,N_39877);
xor U44578 (N_44578,N_35941,N_35271);
and U44579 (N_44579,N_39472,N_39383);
and U44580 (N_44580,N_36172,N_39082);
xor U44581 (N_44581,N_38823,N_36353);
or U44582 (N_44582,N_37178,N_36632);
nor U44583 (N_44583,N_39961,N_35715);
xor U44584 (N_44584,N_36616,N_38596);
nor U44585 (N_44585,N_35733,N_38765);
nand U44586 (N_44586,N_37704,N_36077);
nor U44587 (N_44587,N_35161,N_37643);
xnor U44588 (N_44588,N_35618,N_38738);
nor U44589 (N_44589,N_37746,N_39599);
or U44590 (N_44590,N_35343,N_35117);
nor U44591 (N_44591,N_39233,N_38648);
nor U44592 (N_44592,N_35481,N_39350);
nand U44593 (N_44593,N_39765,N_39478);
xnor U44594 (N_44594,N_35213,N_39903);
nand U44595 (N_44595,N_35149,N_39167);
nor U44596 (N_44596,N_37193,N_39553);
nand U44597 (N_44597,N_37923,N_36254);
or U44598 (N_44598,N_35526,N_36606);
nand U44599 (N_44599,N_36912,N_37866);
and U44600 (N_44600,N_36932,N_35747);
nand U44601 (N_44601,N_38405,N_36874);
nor U44602 (N_44602,N_39165,N_37291);
and U44603 (N_44603,N_37860,N_37035);
and U44604 (N_44604,N_35578,N_35136);
xor U44605 (N_44605,N_37203,N_39458);
xnor U44606 (N_44606,N_39981,N_35340);
nor U44607 (N_44607,N_39945,N_37456);
nand U44608 (N_44608,N_36326,N_35045);
and U44609 (N_44609,N_37094,N_35523);
nor U44610 (N_44610,N_38664,N_36318);
xor U44611 (N_44611,N_39920,N_38455);
xnor U44612 (N_44612,N_37090,N_39815);
or U44613 (N_44613,N_38620,N_37472);
and U44614 (N_44614,N_39331,N_38712);
and U44615 (N_44615,N_38634,N_37527);
xnor U44616 (N_44616,N_36404,N_38584);
and U44617 (N_44617,N_38375,N_39843);
and U44618 (N_44618,N_36687,N_35768);
nor U44619 (N_44619,N_35896,N_37441);
and U44620 (N_44620,N_35025,N_35511);
nand U44621 (N_44621,N_37086,N_38144);
nor U44622 (N_44622,N_36551,N_39290);
nand U44623 (N_44623,N_36012,N_37834);
nor U44624 (N_44624,N_36111,N_39268);
or U44625 (N_44625,N_37859,N_35569);
nand U44626 (N_44626,N_38489,N_37246);
nand U44627 (N_44627,N_39678,N_36598);
nor U44628 (N_44628,N_35507,N_37097);
or U44629 (N_44629,N_39580,N_35412);
nand U44630 (N_44630,N_38326,N_39011);
xor U44631 (N_44631,N_37214,N_39087);
nor U44632 (N_44632,N_37409,N_39976);
or U44633 (N_44633,N_38663,N_37023);
or U44634 (N_44634,N_39215,N_37992);
nor U44635 (N_44635,N_39275,N_35396);
or U44636 (N_44636,N_36691,N_36413);
nor U44637 (N_44637,N_36413,N_35097);
xnor U44638 (N_44638,N_37238,N_36600);
or U44639 (N_44639,N_36853,N_36645);
and U44640 (N_44640,N_36826,N_39922);
xor U44641 (N_44641,N_38898,N_37909);
nand U44642 (N_44642,N_35792,N_37370);
and U44643 (N_44643,N_37111,N_39554);
nor U44644 (N_44644,N_36282,N_39240);
or U44645 (N_44645,N_35906,N_39299);
nor U44646 (N_44646,N_36707,N_36134);
nand U44647 (N_44647,N_37516,N_35828);
xor U44648 (N_44648,N_39800,N_38844);
nor U44649 (N_44649,N_36414,N_37553);
and U44650 (N_44650,N_39268,N_37834);
xnor U44651 (N_44651,N_36422,N_38630);
xor U44652 (N_44652,N_38407,N_36490);
and U44653 (N_44653,N_38372,N_37017);
nand U44654 (N_44654,N_38655,N_35830);
nand U44655 (N_44655,N_37114,N_38044);
and U44656 (N_44656,N_37276,N_39282);
nor U44657 (N_44657,N_39576,N_36261);
nand U44658 (N_44658,N_39634,N_38396);
nor U44659 (N_44659,N_39414,N_37786);
nor U44660 (N_44660,N_37582,N_38158);
xnor U44661 (N_44661,N_39985,N_38635);
and U44662 (N_44662,N_38502,N_37486);
xnor U44663 (N_44663,N_39650,N_38768);
and U44664 (N_44664,N_37777,N_37197);
nor U44665 (N_44665,N_37940,N_36226);
or U44666 (N_44666,N_37231,N_35461);
nor U44667 (N_44667,N_39178,N_35633);
or U44668 (N_44668,N_35460,N_36354);
nand U44669 (N_44669,N_36363,N_39566);
nor U44670 (N_44670,N_38942,N_36444);
nor U44671 (N_44671,N_36028,N_36924);
nand U44672 (N_44672,N_36956,N_35284);
nand U44673 (N_44673,N_37247,N_38853);
nor U44674 (N_44674,N_35847,N_38078);
nand U44675 (N_44675,N_39806,N_35368);
nor U44676 (N_44676,N_35708,N_35185);
nor U44677 (N_44677,N_35919,N_39390);
nand U44678 (N_44678,N_39345,N_36655);
xor U44679 (N_44679,N_39574,N_36311);
and U44680 (N_44680,N_38281,N_35595);
xnor U44681 (N_44681,N_39681,N_38805);
xnor U44682 (N_44682,N_38186,N_36612);
and U44683 (N_44683,N_38666,N_37850);
xor U44684 (N_44684,N_35336,N_37761);
nor U44685 (N_44685,N_39160,N_37091);
or U44686 (N_44686,N_35044,N_35431);
nand U44687 (N_44687,N_37260,N_36193);
nand U44688 (N_44688,N_36985,N_37089);
nand U44689 (N_44689,N_35530,N_35251);
or U44690 (N_44690,N_37020,N_38984);
nand U44691 (N_44691,N_39466,N_36146);
or U44692 (N_44692,N_39782,N_37017);
nor U44693 (N_44693,N_36204,N_38726);
or U44694 (N_44694,N_35794,N_36742);
and U44695 (N_44695,N_39483,N_36325);
or U44696 (N_44696,N_39417,N_35006);
nor U44697 (N_44697,N_39566,N_35047);
or U44698 (N_44698,N_36289,N_37656);
or U44699 (N_44699,N_36030,N_39997);
and U44700 (N_44700,N_36721,N_38990);
xor U44701 (N_44701,N_37787,N_36494);
and U44702 (N_44702,N_38484,N_35064);
nor U44703 (N_44703,N_36661,N_35639);
nand U44704 (N_44704,N_37518,N_36342);
nor U44705 (N_44705,N_35636,N_39465);
and U44706 (N_44706,N_38828,N_37787);
nor U44707 (N_44707,N_36328,N_39207);
and U44708 (N_44708,N_39125,N_37664);
nand U44709 (N_44709,N_35147,N_38894);
xnor U44710 (N_44710,N_36743,N_37483);
nand U44711 (N_44711,N_35175,N_35129);
nand U44712 (N_44712,N_35899,N_38792);
xnor U44713 (N_44713,N_39033,N_35683);
nor U44714 (N_44714,N_38959,N_35407);
nor U44715 (N_44715,N_36974,N_35170);
nor U44716 (N_44716,N_36375,N_38095);
nand U44717 (N_44717,N_37180,N_35602);
nand U44718 (N_44718,N_38135,N_37978);
xor U44719 (N_44719,N_36736,N_38355);
nor U44720 (N_44720,N_37497,N_39147);
or U44721 (N_44721,N_35333,N_36873);
nor U44722 (N_44722,N_36460,N_35600);
xor U44723 (N_44723,N_38829,N_37552);
or U44724 (N_44724,N_39169,N_37641);
or U44725 (N_44725,N_38306,N_37137);
and U44726 (N_44726,N_35103,N_36240);
xor U44727 (N_44727,N_39174,N_39139);
and U44728 (N_44728,N_39084,N_38000);
nor U44729 (N_44729,N_38696,N_36931);
nand U44730 (N_44730,N_36388,N_37368);
nor U44731 (N_44731,N_39307,N_37196);
xnor U44732 (N_44732,N_38904,N_37950);
nand U44733 (N_44733,N_38608,N_35717);
nor U44734 (N_44734,N_36476,N_36537);
nand U44735 (N_44735,N_35928,N_38052);
nor U44736 (N_44736,N_39111,N_35622);
nand U44737 (N_44737,N_37657,N_38467);
nor U44738 (N_44738,N_39609,N_39278);
and U44739 (N_44739,N_36627,N_36476);
xnor U44740 (N_44740,N_35441,N_38566);
xnor U44741 (N_44741,N_39644,N_39111);
and U44742 (N_44742,N_39812,N_37823);
nor U44743 (N_44743,N_35459,N_38781);
xor U44744 (N_44744,N_36475,N_36516);
and U44745 (N_44745,N_36222,N_36503);
or U44746 (N_44746,N_38200,N_37450);
xnor U44747 (N_44747,N_35382,N_36066);
xnor U44748 (N_44748,N_35623,N_35062);
or U44749 (N_44749,N_37751,N_36334);
xor U44750 (N_44750,N_36238,N_36356);
xor U44751 (N_44751,N_38982,N_35803);
nor U44752 (N_44752,N_36400,N_36891);
nor U44753 (N_44753,N_35937,N_36666);
nand U44754 (N_44754,N_39403,N_38874);
nand U44755 (N_44755,N_35125,N_36258);
nor U44756 (N_44756,N_37372,N_38486);
nand U44757 (N_44757,N_38464,N_38155);
xnor U44758 (N_44758,N_35841,N_39779);
or U44759 (N_44759,N_36804,N_35391);
nand U44760 (N_44760,N_38226,N_35410);
nor U44761 (N_44761,N_35457,N_36531);
nand U44762 (N_44762,N_35443,N_36251);
nand U44763 (N_44763,N_35528,N_35997);
and U44764 (N_44764,N_39032,N_35524);
and U44765 (N_44765,N_39026,N_38003);
or U44766 (N_44766,N_35908,N_38477);
and U44767 (N_44767,N_39768,N_38598);
nor U44768 (N_44768,N_39898,N_36041);
nand U44769 (N_44769,N_39816,N_39473);
and U44770 (N_44770,N_39901,N_38679);
or U44771 (N_44771,N_39870,N_38402);
nand U44772 (N_44772,N_37006,N_39756);
or U44773 (N_44773,N_39419,N_36043);
and U44774 (N_44774,N_36165,N_36693);
xnor U44775 (N_44775,N_36929,N_37480);
and U44776 (N_44776,N_38898,N_39596);
nor U44777 (N_44777,N_39359,N_35445);
nand U44778 (N_44778,N_37057,N_36986);
or U44779 (N_44779,N_37115,N_35398);
nand U44780 (N_44780,N_38382,N_36168);
and U44781 (N_44781,N_38272,N_35082);
nand U44782 (N_44782,N_35159,N_39124);
or U44783 (N_44783,N_35967,N_36965);
nand U44784 (N_44784,N_39443,N_37106);
or U44785 (N_44785,N_37844,N_35938);
nand U44786 (N_44786,N_38238,N_35813);
and U44787 (N_44787,N_37731,N_38263);
or U44788 (N_44788,N_39352,N_37805);
nand U44789 (N_44789,N_39595,N_37640);
nor U44790 (N_44790,N_38233,N_37966);
and U44791 (N_44791,N_36457,N_39269);
and U44792 (N_44792,N_39558,N_38301);
and U44793 (N_44793,N_38132,N_35824);
nor U44794 (N_44794,N_39032,N_38985);
or U44795 (N_44795,N_35073,N_38068);
nand U44796 (N_44796,N_37650,N_36157);
nand U44797 (N_44797,N_35138,N_36263);
nand U44798 (N_44798,N_38931,N_37868);
nor U44799 (N_44799,N_39566,N_35523);
nand U44800 (N_44800,N_37672,N_37551);
nand U44801 (N_44801,N_36854,N_38595);
or U44802 (N_44802,N_39805,N_38874);
xnor U44803 (N_44803,N_35099,N_39158);
and U44804 (N_44804,N_38318,N_35117);
or U44805 (N_44805,N_39778,N_39830);
nor U44806 (N_44806,N_38459,N_36890);
nand U44807 (N_44807,N_37573,N_38361);
and U44808 (N_44808,N_35354,N_39275);
and U44809 (N_44809,N_35558,N_35660);
xor U44810 (N_44810,N_36020,N_39244);
nor U44811 (N_44811,N_38796,N_37672);
nand U44812 (N_44812,N_39065,N_36207);
nand U44813 (N_44813,N_38635,N_37309);
nor U44814 (N_44814,N_36580,N_35828);
xor U44815 (N_44815,N_35942,N_39016);
or U44816 (N_44816,N_38684,N_39922);
nand U44817 (N_44817,N_39237,N_39796);
and U44818 (N_44818,N_37086,N_36503);
nand U44819 (N_44819,N_38109,N_35471);
or U44820 (N_44820,N_35620,N_37660);
xor U44821 (N_44821,N_38384,N_36066);
or U44822 (N_44822,N_35698,N_36776);
nor U44823 (N_44823,N_38776,N_38304);
or U44824 (N_44824,N_36343,N_35593);
xor U44825 (N_44825,N_35665,N_38458);
or U44826 (N_44826,N_38267,N_38671);
nand U44827 (N_44827,N_36956,N_38020);
nor U44828 (N_44828,N_36187,N_35408);
or U44829 (N_44829,N_37537,N_38270);
and U44830 (N_44830,N_35923,N_36112);
and U44831 (N_44831,N_37562,N_38508);
xor U44832 (N_44832,N_38489,N_38299);
xnor U44833 (N_44833,N_36942,N_37699);
xor U44834 (N_44834,N_37384,N_35009);
nand U44835 (N_44835,N_36166,N_36735);
or U44836 (N_44836,N_38706,N_39530);
nor U44837 (N_44837,N_36738,N_38565);
nor U44838 (N_44838,N_35946,N_35748);
nor U44839 (N_44839,N_38215,N_35328);
nand U44840 (N_44840,N_35903,N_37229);
xnor U44841 (N_44841,N_36228,N_39278);
or U44842 (N_44842,N_36147,N_38397);
and U44843 (N_44843,N_35004,N_38807);
nor U44844 (N_44844,N_36981,N_37752);
nor U44845 (N_44845,N_35797,N_37330);
or U44846 (N_44846,N_35776,N_36983);
and U44847 (N_44847,N_36763,N_36448);
or U44848 (N_44848,N_38839,N_37196);
xor U44849 (N_44849,N_37709,N_38410);
xor U44850 (N_44850,N_39714,N_36813);
xor U44851 (N_44851,N_37923,N_38630);
and U44852 (N_44852,N_38058,N_38626);
or U44853 (N_44853,N_39508,N_35220);
or U44854 (N_44854,N_39390,N_36043);
xor U44855 (N_44855,N_39725,N_35724);
or U44856 (N_44856,N_38852,N_38316);
and U44857 (N_44857,N_38906,N_36832);
nand U44858 (N_44858,N_35798,N_38065);
xnor U44859 (N_44859,N_39222,N_36658);
nand U44860 (N_44860,N_36938,N_35795);
nand U44861 (N_44861,N_38120,N_37591);
xnor U44862 (N_44862,N_36750,N_36220);
or U44863 (N_44863,N_37092,N_37321);
or U44864 (N_44864,N_38238,N_37194);
and U44865 (N_44865,N_37326,N_38383);
and U44866 (N_44866,N_36401,N_37035);
or U44867 (N_44867,N_39809,N_39390);
or U44868 (N_44868,N_37401,N_35620);
and U44869 (N_44869,N_38228,N_39767);
or U44870 (N_44870,N_39726,N_38164);
nor U44871 (N_44871,N_38239,N_35749);
nand U44872 (N_44872,N_39344,N_35765);
and U44873 (N_44873,N_39630,N_38580);
nor U44874 (N_44874,N_35468,N_36117);
nand U44875 (N_44875,N_39247,N_36810);
xnor U44876 (N_44876,N_35092,N_37260);
or U44877 (N_44877,N_37655,N_35251);
or U44878 (N_44878,N_38621,N_39047);
nand U44879 (N_44879,N_37385,N_35030);
or U44880 (N_44880,N_39607,N_37070);
or U44881 (N_44881,N_38993,N_36802);
xnor U44882 (N_44882,N_36601,N_38636);
nor U44883 (N_44883,N_35584,N_35105);
xor U44884 (N_44884,N_37766,N_35147);
or U44885 (N_44885,N_38811,N_35103);
nand U44886 (N_44886,N_36571,N_39188);
nor U44887 (N_44887,N_39199,N_36146);
xnor U44888 (N_44888,N_35021,N_38666);
xor U44889 (N_44889,N_38680,N_36269);
xnor U44890 (N_44890,N_38642,N_39474);
nand U44891 (N_44891,N_35494,N_37401);
and U44892 (N_44892,N_37661,N_35447);
xor U44893 (N_44893,N_38843,N_38248);
nor U44894 (N_44894,N_37551,N_37129);
nand U44895 (N_44895,N_36413,N_39457);
nand U44896 (N_44896,N_36715,N_37030);
or U44897 (N_44897,N_38663,N_35417);
nand U44898 (N_44898,N_36199,N_38837);
nand U44899 (N_44899,N_37530,N_38659);
nand U44900 (N_44900,N_35368,N_37492);
xor U44901 (N_44901,N_36070,N_39864);
xor U44902 (N_44902,N_39502,N_39986);
xnor U44903 (N_44903,N_38818,N_38904);
or U44904 (N_44904,N_38504,N_35068);
and U44905 (N_44905,N_37454,N_37780);
nand U44906 (N_44906,N_39482,N_39992);
nor U44907 (N_44907,N_35049,N_38619);
nand U44908 (N_44908,N_36113,N_36187);
or U44909 (N_44909,N_35122,N_38526);
and U44910 (N_44910,N_38446,N_38210);
and U44911 (N_44911,N_38497,N_35137);
nand U44912 (N_44912,N_38064,N_36454);
xor U44913 (N_44913,N_36583,N_37812);
or U44914 (N_44914,N_35696,N_37541);
nor U44915 (N_44915,N_36238,N_35008);
nand U44916 (N_44916,N_39061,N_36920);
xor U44917 (N_44917,N_37714,N_39512);
nand U44918 (N_44918,N_36139,N_38259);
and U44919 (N_44919,N_37146,N_35675);
nor U44920 (N_44920,N_38586,N_35441);
xor U44921 (N_44921,N_38101,N_36150);
xor U44922 (N_44922,N_39145,N_37299);
or U44923 (N_44923,N_36130,N_36773);
nor U44924 (N_44924,N_38149,N_35503);
nand U44925 (N_44925,N_36075,N_35539);
and U44926 (N_44926,N_35539,N_37670);
nand U44927 (N_44927,N_39328,N_35437);
or U44928 (N_44928,N_36866,N_38922);
nand U44929 (N_44929,N_36266,N_37129);
nor U44930 (N_44930,N_35681,N_38776);
nor U44931 (N_44931,N_39088,N_36179);
xor U44932 (N_44932,N_39940,N_35513);
or U44933 (N_44933,N_37855,N_37221);
nor U44934 (N_44934,N_38571,N_37534);
nand U44935 (N_44935,N_39610,N_35431);
xnor U44936 (N_44936,N_39959,N_35333);
or U44937 (N_44937,N_39094,N_35345);
nor U44938 (N_44938,N_38460,N_38840);
nand U44939 (N_44939,N_35070,N_38540);
nor U44940 (N_44940,N_39031,N_39577);
or U44941 (N_44941,N_37352,N_37106);
and U44942 (N_44942,N_35509,N_36264);
nor U44943 (N_44943,N_36769,N_35657);
or U44944 (N_44944,N_38248,N_37626);
nor U44945 (N_44945,N_35828,N_35587);
nor U44946 (N_44946,N_37863,N_38757);
xor U44947 (N_44947,N_38767,N_36181);
xor U44948 (N_44948,N_38849,N_35980);
or U44949 (N_44949,N_36762,N_37878);
xnor U44950 (N_44950,N_38728,N_38847);
or U44951 (N_44951,N_39609,N_38003);
and U44952 (N_44952,N_36169,N_36176);
and U44953 (N_44953,N_39772,N_35370);
or U44954 (N_44954,N_35759,N_37510);
and U44955 (N_44955,N_37123,N_36094);
or U44956 (N_44956,N_39940,N_38002);
nor U44957 (N_44957,N_36761,N_39784);
or U44958 (N_44958,N_38251,N_38419);
nand U44959 (N_44959,N_38318,N_39087);
or U44960 (N_44960,N_38117,N_35121);
or U44961 (N_44961,N_35511,N_38908);
and U44962 (N_44962,N_37756,N_38102);
nor U44963 (N_44963,N_38626,N_35796);
xnor U44964 (N_44964,N_35546,N_35915);
or U44965 (N_44965,N_38101,N_35338);
or U44966 (N_44966,N_36073,N_38235);
xor U44967 (N_44967,N_39229,N_39365);
xor U44968 (N_44968,N_39822,N_39960);
and U44969 (N_44969,N_35262,N_38965);
xor U44970 (N_44970,N_35184,N_35117);
nand U44971 (N_44971,N_36274,N_36213);
or U44972 (N_44972,N_35064,N_38984);
xor U44973 (N_44973,N_39747,N_35694);
and U44974 (N_44974,N_38648,N_37308);
or U44975 (N_44975,N_36244,N_37162);
nor U44976 (N_44976,N_37568,N_38519);
nand U44977 (N_44977,N_36435,N_37105);
or U44978 (N_44978,N_36274,N_38573);
nor U44979 (N_44979,N_39792,N_38208);
or U44980 (N_44980,N_36820,N_37647);
nor U44981 (N_44981,N_38881,N_36794);
xnor U44982 (N_44982,N_36514,N_35259);
nor U44983 (N_44983,N_37709,N_37111);
nor U44984 (N_44984,N_39444,N_39290);
nor U44985 (N_44985,N_35388,N_39102);
nand U44986 (N_44986,N_38686,N_37563);
nand U44987 (N_44987,N_39651,N_36132);
xnor U44988 (N_44988,N_39695,N_37582);
nand U44989 (N_44989,N_35326,N_38325);
nor U44990 (N_44990,N_38087,N_36978);
nand U44991 (N_44991,N_38972,N_35280);
nor U44992 (N_44992,N_35450,N_36099);
nand U44993 (N_44993,N_35499,N_38040);
xor U44994 (N_44994,N_38125,N_37071);
xnor U44995 (N_44995,N_35489,N_39551);
or U44996 (N_44996,N_39623,N_37199);
nor U44997 (N_44997,N_39239,N_35164);
nor U44998 (N_44998,N_35345,N_39359);
and U44999 (N_44999,N_35891,N_36816);
nor U45000 (N_45000,N_44447,N_43886);
or U45001 (N_45001,N_43375,N_42938);
xnor U45002 (N_45002,N_41169,N_41270);
nor U45003 (N_45003,N_44863,N_41294);
xnor U45004 (N_45004,N_42273,N_42757);
xnor U45005 (N_45005,N_41666,N_44595);
nand U45006 (N_45006,N_44933,N_41899);
and U45007 (N_45007,N_43645,N_42627);
and U45008 (N_45008,N_40608,N_42105);
nand U45009 (N_45009,N_42220,N_41988);
xnor U45010 (N_45010,N_40165,N_42911);
xnor U45011 (N_45011,N_43474,N_41587);
and U45012 (N_45012,N_42169,N_40888);
xnor U45013 (N_45013,N_44841,N_42988);
or U45014 (N_45014,N_43608,N_42849);
and U45015 (N_45015,N_42855,N_44230);
or U45016 (N_45016,N_42181,N_42623);
and U45017 (N_45017,N_44766,N_44343);
or U45018 (N_45018,N_43925,N_43594);
or U45019 (N_45019,N_40521,N_43577);
xnor U45020 (N_45020,N_41365,N_43634);
nor U45021 (N_45021,N_44453,N_40249);
nor U45022 (N_45022,N_43847,N_41547);
xnor U45023 (N_45023,N_40176,N_44337);
or U45024 (N_45024,N_43076,N_40857);
and U45025 (N_45025,N_41132,N_40152);
nand U45026 (N_45026,N_42585,N_40821);
nor U45027 (N_45027,N_44003,N_42355);
nor U45028 (N_45028,N_42636,N_42526);
nor U45029 (N_45029,N_44523,N_41558);
or U45030 (N_45030,N_40491,N_44200);
and U45031 (N_45031,N_43765,N_40131);
and U45032 (N_45032,N_42511,N_43566);
or U45033 (N_45033,N_41212,N_42590);
nand U45034 (N_45034,N_42824,N_44035);
xnor U45035 (N_45035,N_41425,N_43141);
nor U45036 (N_45036,N_42396,N_42516);
nand U45037 (N_45037,N_43912,N_44616);
or U45038 (N_45038,N_44549,N_43398);
nor U45039 (N_45039,N_44111,N_40171);
xor U45040 (N_45040,N_44402,N_40289);
nor U45041 (N_45041,N_44556,N_40590);
nor U45042 (N_45042,N_44936,N_41143);
nand U45043 (N_45043,N_44949,N_41936);
nand U45044 (N_45044,N_44182,N_41252);
and U45045 (N_45045,N_42972,N_40230);
and U45046 (N_45046,N_44735,N_42225);
nand U45047 (N_45047,N_43845,N_43533);
or U45048 (N_45048,N_40890,N_44350);
and U45049 (N_45049,N_44618,N_42012);
or U45050 (N_45050,N_44123,N_44012);
nand U45051 (N_45051,N_40819,N_41522);
nor U45052 (N_45052,N_41594,N_41351);
or U45053 (N_45053,N_42010,N_41675);
nand U45054 (N_45054,N_42711,N_40808);
or U45055 (N_45055,N_43130,N_42200);
and U45056 (N_45056,N_43035,N_43491);
or U45057 (N_45057,N_40045,N_43430);
nor U45058 (N_45058,N_40381,N_41827);
nor U45059 (N_45059,N_44341,N_43642);
xnor U45060 (N_45060,N_44292,N_42352);
or U45061 (N_45061,N_43609,N_43325);
nor U45062 (N_45062,N_41766,N_44531);
nand U45063 (N_45063,N_40112,N_40475);
xor U45064 (N_45064,N_41427,N_43259);
nor U45065 (N_45065,N_42118,N_40244);
and U45066 (N_45066,N_41886,N_42996);
and U45067 (N_45067,N_42382,N_43535);
and U45068 (N_45068,N_42197,N_41526);
or U45069 (N_45069,N_40267,N_42532);
or U45070 (N_45070,N_41388,N_43589);
nand U45071 (N_45071,N_40101,N_44696);
and U45072 (N_45072,N_44829,N_44150);
nand U45073 (N_45073,N_40735,N_43767);
or U45074 (N_45074,N_41997,N_44855);
nor U45075 (N_45075,N_40726,N_40777);
or U45076 (N_45076,N_40837,N_44299);
nor U45077 (N_45077,N_44922,N_43882);
or U45078 (N_45078,N_40552,N_40030);
nand U45079 (N_45079,N_44613,N_43809);
nand U45080 (N_45080,N_41055,N_41011);
nand U45081 (N_45081,N_44653,N_42402);
and U45082 (N_45082,N_41314,N_43667);
xnor U45083 (N_45083,N_42359,N_42536);
xor U45084 (N_45084,N_44026,N_40015);
nor U45085 (N_45085,N_42228,N_41811);
xor U45086 (N_45086,N_41721,N_42686);
xor U45087 (N_45087,N_40425,N_40712);
nand U45088 (N_45088,N_43274,N_40778);
and U45089 (N_45089,N_41367,N_44311);
and U45090 (N_45090,N_43394,N_40620);
xnor U45091 (N_45091,N_43741,N_43607);
nand U45092 (N_45092,N_43873,N_40321);
nor U45093 (N_45093,N_42769,N_42347);
or U45094 (N_45094,N_44039,N_40013);
nand U45095 (N_45095,N_44471,N_41507);
nor U45096 (N_45096,N_42896,N_44421);
or U45097 (N_45097,N_43071,N_40632);
or U45098 (N_45098,N_44663,N_42377);
and U45099 (N_45099,N_42159,N_43486);
xor U45100 (N_45100,N_43321,N_42109);
nand U45101 (N_45101,N_41433,N_43456);
nor U45102 (N_45102,N_40347,N_44574);
and U45103 (N_45103,N_40629,N_40391);
and U45104 (N_45104,N_42276,N_43461);
or U45105 (N_45105,N_43303,N_41250);
nor U45106 (N_45106,N_40594,N_40037);
nor U45107 (N_45107,N_40515,N_41329);
nor U45108 (N_45108,N_43754,N_40755);
nor U45109 (N_45109,N_40569,N_44697);
nand U45110 (N_45110,N_42662,N_43143);
or U45111 (N_45111,N_40811,N_43763);
xor U45112 (N_45112,N_43999,N_44216);
xor U45113 (N_45113,N_40469,N_41895);
xnor U45114 (N_45114,N_41893,N_40105);
xnor U45115 (N_45115,N_43580,N_43188);
xnor U45116 (N_45116,N_40779,N_41605);
nor U45117 (N_45117,N_42665,N_41945);
xor U45118 (N_45118,N_40287,N_43702);
nor U45119 (N_45119,N_42663,N_44361);
nand U45120 (N_45120,N_40799,N_42306);
nand U45121 (N_45121,N_43406,N_44891);
nand U45122 (N_45122,N_42784,N_41646);
xor U45123 (N_45123,N_44450,N_42198);
xnor U45124 (N_45124,N_40433,N_42263);
nor U45125 (N_45125,N_40946,N_41154);
nor U45126 (N_45126,N_44334,N_44083);
xnor U45127 (N_45127,N_40402,N_42016);
nand U45128 (N_45128,N_42839,N_41468);
and U45129 (N_45129,N_42944,N_44995);
nand U45130 (N_45130,N_41649,N_40276);
nor U45131 (N_45131,N_40256,N_41905);
nand U45132 (N_45132,N_44161,N_44590);
nand U45133 (N_45133,N_42270,N_43373);
and U45134 (N_45134,N_44062,N_41943);
or U45135 (N_45135,N_41268,N_43689);
or U45136 (N_45136,N_41242,N_44907);
nor U45137 (N_45137,N_42042,N_43412);
xor U45138 (N_45138,N_43981,N_40965);
and U45139 (N_45139,N_42094,N_40748);
nor U45140 (N_45140,N_42316,N_40702);
and U45141 (N_45141,N_43249,N_40758);
xor U45142 (N_45142,N_40541,N_42930);
or U45143 (N_45143,N_43938,N_40762);
nor U45144 (N_45144,N_41034,N_40605);
and U45145 (N_45145,N_42956,N_41295);
nand U45146 (N_45146,N_43048,N_40047);
xor U45147 (N_45147,N_43330,N_42335);
xor U45148 (N_45148,N_41640,N_41165);
xnor U45149 (N_45149,N_43895,N_42780);
or U45150 (N_45150,N_42542,N_41681);
xnor U45151 (N_45151,N_43152,N_41138);
nor U45152 (N_45152,N_41341,N_42976);
and U45153 (N_45153,N_42218,N_40102);
xor U45154 (N_45154,N_40023,N_40745);
nor U45155 (N_45155,N_40470,N_42737);
nand U45156 (N_45156,N_40722,N_43069);
or U45157 (N_45157,N_43990,N_40931);
nor U45158 (N_45158,N_40048,N_44815);
or U45159 (N_45159,N_40424,N_44888);
xnor U45160 (N_45160,N_41107,N_42458);
nor U45161 (N_45161,N_44024,N_40178);
xnor U45162 (N_45162,N_40797,N_42264);
nand U45163 (N_45163,N_41791,N_40246);
or U45164 (N_45164,N_41103,N_41933);
or U45165 (N_45165,N_42692,N_40853);
or U45166 (N_45166,N_40365,N_44484);
xnor U45167 (N_45167,N_44319,N_40816);
nor U45168 (N_45168,N_44828,N_42670);
nor U45169 (N_45169,N_44281,N_44972);
and U45170 (N_45170,N_40099,N_44767);
nor U45171 (N_45171,N_42926,N_43180);
or U45172 (N_45172,N_40460,N_44004);
or U45173 (N_45173,N_42986,N_42281);
nand U45174 (N_45174,N_44937,N_40896);
nand U45175 (N_45175,N_42762,N_42096);
or U45176 (N_45176,N_43902,N_40235);
xnor U45177 (N_45177,N_40512,N_40969);
and U45178 (N_45178,N_40690,N_40125);
or U45179 (N_45179,N_44699,N_40567);
xor U45180 (N_45180,N_44301,N_44592);
nor U45181 (N_45181,N_42861,N_42998);
nand U45182 (N_45182,N_44273,N_40883);
and U45183 (N_45183,N_42252,N_40094);
or U45184 (N_45184,N_40867,N_42332);
and U45185 (N_45185,N_44383,N_41908);
xor U45186 (N_45186,N_44969,N_43993);
or U45187 (N_45187,N_43386,N_44858);
or U45188 (N_45188,N_42069,N_43875);
xor U45189 (N_45189,N_44073,N_41368);
or U45190 (N_45190,N_41742,N_41043);
nand U45191 (N_45191,N_41773,N_42560);
or U45192 (N_45192,N_40150,N_42447);
xor U45193 (N_45193,N_44877,N_43883);
xnor U45194 (N_45194,N_44967,N_42357);
and U45195 (N_45195,N_40742,N_44483);
or U45196 (N_45196,N_41027,N_41751);
nand U45197 (N_45197,N_41870,N_40610);
or U45198 (N_45198,N_43813,N_42315);
or U45199 (N_45199,N_42773,N_44805);
xnor U45200 (N_45200,N_40411,N_43155);
xnor U45201 (N_45201,N_41115,N_40582);
nand U45202 (N_45202,N_41450,N_43764);
or U45203 (N_45203,N_43221,N_41041);
and U45204 (N_45204,N_41105,N_40472);
xor U45205 (N_45205,N_40053,N_44948);
nor U45206 (N_45206,N_40953,N_43448);
xor U45207 (N_45207,N_42760,N_43779);
nor U45208 (N_45208,N_44776,N_42939);
or U45209 (N_45209,N_44602,N_40824);
and U45210 (N_45210,N_41150,N_44700);
or U45211 (N_45211,N_41039,N_44676);
nor U45212 (N_45212,N_44226,N_41982);
nand U45213 (N_45213,N_43851,N_44196);
or U45214 (N_45214,N_43279,N_40790);
nand U45215 (N_45215,N_43670,N_41475);
nor U45216 (N_45216,N_41566,N_43294);
and U45217 (N_45217,N_41865,N_42249);
or U45218 (N_45218,N_42707,N_42968);
nand U45219 (N_45219,N_44757,N_40040);
xor U45220 (N_45220,N_42660,N_41494);
nand U45221 (N_45221,N_41922,N_41562);
nand U45222 (N_45222,N_40507,N_41848);
nand U45223 (N_45223,N_42768,N_42212);
nand U45224 (N_45224,N_42024,N_41202);
xnor U45225 (N_45225,N_44156,N_41528);
xor U45226 (N_45226,N_42958,N_43418);
or U45227 (N_45227,N_42597,N_44306);
nand U45228 (N_45228,N_43821,N_40447);
nor U45229 (N_45229,N_41434,N_40630);
or U45230 (N_45230,N_43433,N_40041);
or U45231 (N_45231,N_42476,N_41812);
xnor U45232 (N_45232,N_42605,N_44109);
nor U45233 (N_45233,N_42201,N_41800);
xor U45234 (N_45234,N_41794,N_40090);
or U45235 (N_45235,N_41923,N_44737);
nand U45236 (N_45236,N_44474,N_44218);
nand U45237 (N_45237,N_43811,N_42090);
xor U45238 (N_45238,N_44647,N_40323);
and U45239 (N_45239,N_43653,N_41621);
and U45240 (N_45240,N_43151,N_41354);
xor U45241 (N_45241,N_41338,N_42833);
and U45242 (N_45242,N_44621,N_43116);
or U45243 (N_45243,N_44606,N_42606);
xnor U45244 (N_45244,N_42124,N_44923);
nor U45245 (N_45245,N_44790,N_44690);
nand U45246 (N_45246,N_43336,N_43929);
xnor U45247 (N_45247,N_41819,N_44310);
xnor U45248 (N_45248,N_40951,N_42832);
or U45249 (N_45249,N_44581,N_42565);
nor U45250 (N_45250,N_41086,N_44393);
nor U45251 (N_45251,N_40604,N_41406);
or U45252 (N_45252,N_42406,N_43047);
nor U45253 (N_45253,N_42884,N_42555);
nand U45254 (N_45254,N_42953,N_43078);
and U45255 (N_45255,N_40038,N_42369);
or U45256 (N_45256,N_41009,N_41611);
or U45257 (N_45257,N_41133,N_42806);
xnor U45258 (N_45258,N_43040,N_40028);
xor U45259 (N_45259,N_42550,N_44118);
nand U45260 (N_45260,N_43407,N_43000);
xnor U45261 (N_45261,N_40075,N_41629);
nand U45262 (N_45262,N_43157,N_41961);
xor U45263 (N_45263,N_42966,N_42664);
nand U45264 (N_45264,N_40719,N_43499);
and U45265 (N_45265,N_41173,N_40432);
nand U45266 (N_45266,N_43296,N_42060);
and U45267 (N_45267,N_43198,N_41387);
or U45268 (N_45268,N_42150,N_44479);
or U45269 (N_45269,N_42018,N_44679);
xor U45270 (N_45270,N_44518,N_44555);
xnor U45271 (N_45271,N_42436,N_41733);
and U45272 (N_45272,N_43257,N_40376);
nand U45273 (N_45273,N_42653,N_43013);
nor U45274 (N_45274,N_41277,N_40255);
or U45275 (N_45275,N_42815,N_42876);
and U45276 (N_45276,N_43361,N_40410);
or U45277 (N_45277,N_43639,N_40653);
nand U45278 (N_45278,N_42701,N_42479);
nand U45279 (N_45279,N_42233,N_44803);
and U45280 (N_45280,N_44373,N_44053);
xor U45281 (N_45281,N_42795,N_44030);
nor U45282 (N_45282,N_43314,N_40396);
xor U45283 (N_45283,N_43231,N_41648);
and U45284 (N_45284,N_42433,N_41977);
or U45285 (N_45285,N_43242,N_40714);
and U45286 (N_45286,N_40282,N_42743);
nand U45287 (N_45287,N_40835,N_43260);
nand U45288 (N_45288,N_44353,N_43675);
nand U45289 (N_45289,N_41140,N_40813);
and U45290 (N_45290,N_43001,N_43285);
nand U45291 (N_45291,N_43972,N_44975);
nor U45292 (N_45292,N_43822,N_43072);
nor U45293 (N_45293,N_40976,N_42363);
nand U45294 (N_45294,N_40337,N_41904);
or U45295 (N_45295,N_43804,N_42850);
nor U45296 (N_45296,N_44515,N_41509);
xor U45297 (N_45297,N_44599,N_44104);
or U45298 (N_45298,N_44362,N_41604);
or U45299 (N_45299,N_44138,N_44762);
or U45300 (N_45300,N_41471,N_44066);
xor U45301 (N_45301,N_41006,N_41940);
or U45302 (N_45302,N_40736,N_41631);
nor U45303 (N_45303,N_44856,N_42298);
or U45304 (N_45304,N_41343,N_43464);
xor U45305 (N_45305,N_42652,N_41797);
nor U45306 (N_45306,N_41962,N_41525);
nor U45307 (N_45307,N_41290,N_41069);
or U45308 (N_45308,N_44022,N_44628);
or U45309 (N_45309,N_42919,N_41410);
nor U45310 (N_45310,N_44594,N_41535);
nand U45311 (N_45311,N_42008,N_41803);
or U45312 (N_45312,N_41686,N_41430);
xor U45313 (N_45313,N_43842,N_44905);
and U45314 (N_45314,N_40830,N_44055);
nor U45315 (N_45315,N_40467,N_43651);
nor U45316 (N_45316,N_44386,N_42381);
and U45317 (N_45317,N_43916,N_41466);
nand U45318 (N_45318,N_42822,N_41722);
and U45319 (N_45319,N_41839,N_43050);
xor U45320 (N_45320,N_43801,N_42717);
nand U45321 (N_45321,N_44651,N_44020);
nor U45322 (N_45322,N_40670,N_40263);
and U45323 (N_45323,N_41578,N_41260);
and U45324 (N_45324,N_44149,N_41696);
nand U45325 (N_45325,N_41705,N_41213);
nand U45326 (N_45326,N_44970,N_44296);
xnor U45327 (N_45327,N_44680,N_42860);
or U45328 (N_45328,N_44668,N_41872);
and U45329 (N_45329,N_44826,N_40596);
or U45330 (N_45330,N_40727,N_40860);
xnor U45331 (N_45331,N_44516,N_42716);
xor U45332 (N_45332,N_44333,N_42140);
nand U45333 (N_45333,N_44755,N_42267);
and U45334 (N_45334,N_42778,N_40335);
and U45335 (N_45335,N_43233,N_40279);
nor U45336 (N_45336,N_41040,N_42398);
nor U45337 (N_45337,N_44251,N_40389);
or U45338 (N_45338,N_44712,N_40084);
nor U45339 (N_45339,N_44081,N_42354);
and U45340 (N_45340,N_42487,N_43496);
nor U45341 (N_45341,N_43219,N_41155);
nor U45342 (N_45342,N_44322,N_42823);
or U45343 (N_45343,N_40415,N_40757);
xnor U45344 (N_45344,N_44238,N_41170);
and U45345 (N_45345,N_40925,N_43908);
xnor U45346 (N_45346,N_44040,N_43232);
and U45347 (N_45347,N_41100,N_41072);
or U45348 (N_45348,N_43202,N_42037);
and U45349 (N_45349,N_44874,N_42821);
nor U45350 (N_45350,N_42260,N_44247);
xnor U45351 (N_45351,N_40196,N_44683);
xnor U45352 (N_45352,N_41375,N_40899);
xor U45353 (N_45353,N_43748,N_42954);
xnor U45354 (N_45354,N_42314,N_40769);
nor U45355 (N_45355,N_41673,N_44256);
nand U45356 (N_45356,N_43278,N_41359);
nand U45357 (N_45357,N_40593,N_41552);
xor U45358 (N_45358,N_41110,N_40082);
nand U45359 (N_45359,N_41036,N_43138);
nor U45360 (N_45360,N_40967,N_42345);
and U45361 (N_45361,N_40238,N_43137);
xnor U45362 (N_45362,N_42852,N_40584);
and U45363 (N_45363,N_41976,N_44794);
and U45364 (N_45364,N_42842,N_44637);
or U45365 (N_45365,N_41442,N_42982);
and U45366 (N_45366,N_40897,N_43522);
xor U45367 (N_45367,N_43518,N_42222);
xor U45368 (N_45368,N_42782,N_42294);
nor U45369 (N_45369,N_44538,N_40937);
or U45370 (N_45370,N_41261,N_44655);
or U45371 (N_45371,N_44906,N_42794);
xnor U45372 (N_45372,N_43131,N_40104);
nand U45373 (N_45373,N_42865,N_43490);
and U45374 (N_45374,N_44242,N_41398);
nand U45375 (N_45375,N_40741,N_43719);
and U45376 (N_45376,N_42937,N_44792);
or U45377 (N_45377,N_42735,N_44265);
nor U45378 (N_45378,N_40640,N_40501);
xor U45379 (N_45379,N_43015,N_42759);
and U45380 (N_45380,N_42622,N_42787);
nand U45381 (N_45381,N_42291,N_44671);
xnor U45382 (N_45382,N_43098,N_43211);
or U45383 (N_45383,N_44189,N_44572);
nor U45384 (N_45384,N_40145,N_43696);
nor U45385 (N_45385,N_40909,N_44286);
nor U45386 (N_45386,N_42157,N_43094);
nor U45387 (N_45387,N_43478,N_40342);
nor U45388 (N_45388,N_41088,N_40801);
nand U45389 (N_45389,N_41996,N_41330);
or U45390 (N_45390,N_42631,N_44389);
nor U45391 (N_45391,N_44861,N_44028);
nor U45392 (N_45392,N_40798,N_44406);
nand U45393 (N_45393,N_43403,N_42546);
or U45394 (N_45394,N_42963,N_41855);
nor U45395 (N_45395,N_42728,N_44331);
or U45396 (N_45396,N_41697,N_43065);
xor U45397 (N_45397,N_42380,N_41163);
xor U45398 (N_45398,N_40681,N_44199);
nor U45399 (N_45399,N_40351,N_40483);
xnor U45400 (N_45400,N_40049,N_41930);
xnor U45401 (N_45401,N_44711,N_40587);
or U45402 (N_45402,N_40122,N_42494);
nand U45403 (N_45403,N_40868,N_41775);
nor U45404 (N_45404,N_43305,N_43789);
nor U45405 (N_45405,N_42830,N_44379);
xor U45406 (N_45406,N_43646,N_44088);
nand U45407 (N_45407,N_40181,N_43721);
xor U45408 (N_45408,N_42223,N_41714);
nor U45409 (N_45409,N_43234,N_40905);
xnor U45410 (N_45410,N_40710,N_43251);
nor U45411 (N_45411,N_42709,N_43898);
nor U45412 (N_45412,N_43544,N_42095);
nand U45413 (N_45413,N_40217,N_43364);
or U45414 (N_45414,N_42870,N_44057);
and U45415 (N_45415,N_44287,N_43376);
xor U45416 (N_45416,N_40912,N_41393);
or U45417 (N_45417,N_44879,N_41752);
nor U45418 (N_45418,N_40961,N_44023);
or U45419 (N_45419,N_44662,N_40536);
or U45420 (N_45420,N_40051,N_40197);
and U45421 (N_45421,N_41370,N_40812);
or U45422 (N_45422,N_41449,N_42286);
or U45423 (N_45423,N_44520,N_41804);
and U45424 (N_45424,N_43725,N_43759);
or U45425 (N_45425,N_40394,N_43149);
nand U45426 (N_45426,N_41125,N_40556);
or U45427 (N_45427,N_41498,N_42819);
nor U45428 (N_45428,N_40307,N_41869);
and U45429 (N_45429,N_40142,N_43162);
nor U45430 (N_45430,N_40699,N_41274);
or U45431 (N_45431,N_40124,N_40110);
nor U45432 (N_45432,N_40206,N_43429);
nand U45433 (N_45433,N_41857,N_41576);
and U45434 (N_45434,N_44997,N_44076);
or U45435 (N_45435,N_41090,N_41517);
and U45436 (N_45436,N_43674,N_41291);
and U45437 (N_45437,N_44367,N_40724);
and U45438 (N_45438,N_42324,N_41946);
nand U45439 (N_45439,N_44812,N_41824);
nand U45440 (N_45440,N_42521,N_41642);
and U45441 (N_45441,N_43465,N_44754);
nand U45442 (N_45442,N_40810,N_43027);
and U45443 (N_45443,N_44627,N_44467);
xnor U45444 (N_45444,N_43275,N_41735);
or U45445 (N_45445,N_43846,N_41207);
and U45446 (N_45446,N_44045,N_42858);
xor U45447 (N_45447,N_40825,N_41748);
nand U45448 (N_45448,N_41137,N_42007);
and U45449 (N_45449,N_44043,N_42552);
nor U45450 (N_45450,N_44597,N_44047);
or U45451 (N_45451,N_44845,N_43632);
and U45452 (N_45452,N_41707,N_40527);
or U45453 (N_45453,N_41674,N_44102);
nand U45454 (N_45454,N_44405,N_41716);
xor U45455 (N_45455,N_44171,N_40850);
nand U45456 (N_45456,N_42828,N_44115);
and U45457 (N_45457,N_42610,N_44259);
or U45458 (N_45458,N_40439,N_41241);
nor U45459 (N_45459,N_41198,N_40317);
or U45460 (N_45460,N_43442,N_40578);
xnor U45461 (N_45461,N_41188,N_44571);
nand U45462 (N_45462,N_44782,N_43785);
or U45463 (N_45463,N_41283,N_43192);
or U45464 (N_45464,N_42322,N_41316);
xor U45465 (N_45465,N_44175,N_42840);
and U45466 (N_45466,N_41740,N_42329);
nor U45467 (N_45467,N_44151,N_40295);
nand U45468 (N_45468,N_42505,N_41938);
or U45469 (N_45469,N_44868,N_40129);
xnor U45470 (N_45470,N_41743,N_41537);
xnor U45471 (N_45471,N_40019,N_43382);
and U45472 (N_45472,N_42426,N_44025);
nor U45473 (N_45473,N_42818,N_40676);
nand U45474 (N_45474,N_41149,N_41285);
nor U45475 (N_45475,N_41369,N_41120);
xnor U45476 (N_45476,N_43387,N_40504);
nand U45477 (N_45477,N_41840,N_40212);
nand U45478 (N_45478,N_43392,N_44212);
nand U45479 (N_45479,N_43968,N_40761);
and U45480 (N_45480,N_43264,N_42992);
or U45481 (N_45481,N_40729,N_42459);
and U45482 (N_45482,N_41142,N_41774);
nor U45483 (N_45483,N_41560,N_41779);
or U45484 (N_45484,N_43550,N_44810);
and U45485 (N_45485,N_42601,N_43046);
and U45486 (N_45486,N_43585,N_42211);
or U45487 (N_45487,N_40173,N_44110);
and U45488 (N_45488,N_42006,N_43659);
and U45489 (N_45489,N_44381,N_43985);
and U45490 (N_45490,N_43541,N_43358);
nand U45491 (N_45491,N_40087,N_40623);
or U45492 (N_45492,N_40682,N_41789);
or U45493 (N_45493,N_42507,N_40526);
or U45494 (N_45494,N_40121,N_44527);
nor U45495 (N_45495,N_41297,N_41238);
nor U45496 (N_45496,N_43663,N_42644);
xor U45497 (N_45497,N_42234,N_44748);
and U45498 (N_45498,N_40468,N_44477);
xnor U45499 (N_45499,N_44021,N_41364);
or U45500 (N_45500,N_44390,N_40166);
xor U45501 (N_45501,N_43841,N_43469);
and U45502 (N_45502,N_43459,N_41529);
or U45503 (N_45503,N_40877,N_44596);
and U45504 (N_45504,N_43800,N_41303);
nor U45505 (N_45505,N_42414,N_40453);
nand U45506 (N_45506,N_41873,N_43983);
or U45507 (N_45507,N_40650,N_41201);
nand U45508 (N_45508,N_41879,N_40773);
xnor U45509 (N_45509,N_41969,N_40399);
nand U45510 (N_45510,N_40941,N_42825);
nor U45511 (N_45511,N_43362,N_44716);
nor U45512 (N_45512,N_40560,N_40502);
nor U45513 (N_45513,N_41296,N_41454);
nand U45514 (N_45514,N_44244,N_41031);
nand U45515 (N_45515,N_41921,N_41047);
xnor U45516 (N_45516,N_40619,N_42661);
nor U45517 (N_45517,N_43085,N_42688);
xor U45518 (N_45518,N_41676,N_40747);
nand U45519 (N_45519,N_42537,N_42366);
or U45520 (N_45520,N_44961,N_44747);
nand U45521 (N_45521,N_42812,N_44116);
nand U45522 (N_45522,N_41711,N_42607);
nand U45523 (N_45523,N_44183,N_41342);
xnor U45524 (N_45524,N_44636,N_43636);
xor U45525 (N_45525,N_44665,N_42204);
nor U45526 (N_45526,N_44087,N_41402);
or U45527 (N_45527,N_44872,N_40219);
xor U45528 (N_45528,N_42632,N_41776);
nor U45529 (N_45529,N_41460,N_41978);
nand U45530 (N_45530,N_42541,N_43187);
xnor U45531 (N_45531,N_41606,N_43984);
xnor U45532 (N_45532,N_40846,N_42905);
nand U45533 (N_45533,N_44441,N_44530);
and U45534 (N_45534,N_44860,N_43783);
xor U45535 (N_45535,N_40806,N_42145);
and U45536 (N_45536,N_43506,N_44136);
xnor U45537 (N_45537,N_43352,N_43308);
or U45538 (N_45538,N_42547,N_42873);
nor U45539 (N_45539,N_41651,N_44061);
and U45540 (N_45540,N_42493,N_40434);
nor U45541 (N_45541,N_43795,N_43128);
nand U45542 (N_45542,N_42650,N_42562);
xnor U45543 (N_45543,N_41963,N_41279);
and U45544 (N_45544,N_43782,N_40649);
and U45545 (N_45545,N_41148,N_44233);
and U45546 (N_45546,N_41372,N_42671);
or U45547 (N_45547,N_40442,N_43927);
nand U45548 (N_45548,N_41632,N_40700);
or U45549 (N_45549,N_43976,N_44512);
nor U45550 (N_45550,N_44126,N_42903);
and U45551 (N_45551,N_44634,N_41128);
nand U45552 (N_45552,N_42971,N_44267);
xor U45553 (N_45553,N_41796,N_40393);
nor U45554 (N_45554,N_42564,N_44262);
nand U45555 (N_45555,N_42789,N_44044);
nand U45556 (N_45556,N_44209,N_40203);
or U45557 (N_45557,N_43084,N_41436);
or U45558 (N_45558,N_44809,N_40942);
nand U45559 (N_45559,N_44525,N_43980);
nand U45560 (N_45560,N_42902,N_40261);
xnor U45561 (N_45561,N_42021,N_43318);
or U45562 (N_45562,N_44279,N_41264);
and U45563 (N_45563,N_43705,N_43239);
or U45564 (N_45564,N_41805,N_41320);
and U45565 (N_45565,N_40576,N_44698);
nand U45566 (N_45566,N_40281,N_43716);
nor U45567 (N_45567,N_44469,N_42764);
and U45568 (N_45568,N_43488,N_43790);
or U45569 (N_45569,N_43957,N_40539);
nand U45570 (N_45570,N_41834,N_43183);
xor U45571 (N_45571,N_41346,N_40116);
nand U45572 (N_45572,N_42640,N_43482);
and U45573 (N_45573,N_40898,N_40754);
nand U45574 (N_45574,N_43868,N_41392);
nand U45575 (N_45575,N_41864,N_44506);
nor U45576 (N_45576,N_42698,N_44190);
xnor U45577 (N_45577,N_43631,N_42442);
and U45578 (N_45578,N_41438,N_41323);
nand U45579 (N_45579,N_43028,N_41122);
xor U45580 (N_45580,N_44852,N_40913);
or U45581 (N_45581,N_40070,N_44382);
and U45582 (N_45582,N_44305,N_43444);
xnor U45583 (N_45583,N_43400,N_42765);
nand U45584 (N_45584,N_43252,N_41421);
and U45585 (N_45585,N_41911,N_43276);
and U45586 (N_45586,N_43717,N_44823);
nor U45587 (N_45587,N_40987,N_41456);
xor U45588 (N_45588,N_44865,N_43007);
nor U45589 (N_45589,N_42501,N_42128);
or U45590 (N_45590,N_44650,N_40654);
nor U45591 (N_45591,N_42615,N_43320);
xor U45592 (N_45592,N_41089,N_43335);
nor U45593 (N_45593,N_41058,N_40471);
xor U45594 (N_45594,N_44140,N_43960);
nor U45595 (N_45595,N_43843,N_43599);
nor U45596 (N_45596,N_43905,N_41081);
or U45597 (N_45597,N_40656,N_41687);
and U45598 (N_45598,N_41248,N_44910);
and U45599 (N_45599,N_43447,N_42964);
nor U45600 (N_45600,N_43893,N_44481);
nor U45601 (N_45601,N_40072,N_40147);
xor U45602 (N_45602,N_43353,N_44519);
or U45603 (N_45603,N_44774,N_40005);
and U45604 (N_45604,N_43189,N_40275);
and U45605 (N_45605,N_40164,N_40663);
nand U45606 (N_45606,N_40167,N_44232);
nand U45607 (N_45607,N_41302,N_44913);
or U45608 (N_45608,N_40952,N_43840);
or U45609 (N_45609,N_40143,N_42053);
and U45610 (N_45610,N_43026,N_43937);
and U45611 (N_45611,N_40269,N_44981);
nor U45612 (N_45612,N_44015,N_40960);
and U45613 (N_45613,N_41702,N_41068);
nand U45614 (N_45614,N_40988,N_42126);
xor U45615 (N_45615,N_44883,N_44130);
nand U45616 (N_45616,N_40201,N_40055);
xnor U45617 (N_45617,N_43136,N_42066);
or U45618 (N_45618,N_44324,N_40153);
nor U45619 (N_45619,N_40908,N_43958);
nand U45620 (N_45620,N_42629,N_44180);
xor U45621 (N_45621,N_41278,N_40111);
nand U45622 (N_45622,N_44449,N_43787);
or U45623 (N_45623,N_42675,N_42296);
xnor U45624 (N_45624,N_40103,N_41030);
nand U45625 (N_45625,N_42438,N_44376);
nor U45626 (N_45626,N_43322,N_42890);
or U45627 (N_45627,N_40346,N_41215);
and U45628 (N_45628,N_40180,N_43552);
nor U45629 (N_45629,N_40170,N_40357);
xnor U45630 (N_45630,N_44313,N_44664);
xor U45631 (N_45631,N_40551,N_44723);
and U45632 (N_45632,N_44709,N_43802);
xnor U45633 (N_45633,N_43956,N_41024);
xor U45634 (N_45634,N_44085,N_41083);
xor U45635 (N_45635,N_43457,N_42859);
or U45636 (N_45636,N_44391,N_42983);
nand U45637 (N_45637,N_40862,N_40371);
and U45638 (N_45638,N_43756,N_42445);
nor U45639 (N_45639,N_41255,N_41478);
xnor U45640 (N_45640,N_42706,N_43413);
or U45641 (N_45641,N_42277,N_40086);
or U45642 (N_45642,N_43647,N_43487);
xnor U45643 (N_45643,N_42637,N_40288);
or U45644 (N_45644,N_43810,N_44094);
or U45645 (N_45645,N_42036,N_43238);
or U45646 (N_45646,N_44365,N_44342);
nor U45647 (N_45647,N_40241,N_44942);
xnor U45648 (N_45648,N_41289,N_40208);
xor U45649 (N_45649,N_44903,N_43752);
or U45650 (N_45650,N_43560,N_41422);
nor U45651 (N_45651,N_43343,N_42950);
and U45652 (N_45652,N_43708,N_41947);
and U45653 (N_45653,N_40689,N_40211);
nor U45654 (N_45654,N_43658,N_40766);
or U45655 (N_45655,N_43263,N_40859);
nand U45656 (N_45656,N_44625,N_43122);
xor U45657 (N_45657,N_41544,N_43132);
or U45658 (N_45658,N_43170,N_42386);
xor U45659 (N_45659,N_41231,N_41902);
or U45660 (N_45660,N_44056,N_42231);
and U45661 (N_45661,N_41756,N_44048);
xor U45662 (N_45662,N_41028,N_43918);
or U45663 (N_45663,N_42563,N_40236);
nor U45664 (N_45664,N_41670,N_40531);
nand U45665 (N_45665,N_42463,N_42935);
xor U45666 (N_45666,N_43606,N_44229);
and U45667 (N_45667,N_44357,N_43870);
and U45668 (N_45668,N_43684,N_44645);
xnor U45669 (N_45669,N_44008,N_44097);
or U45670 (N_45670,N_44925,N_41428);
xor U45671 (N_45671,N_43145,N_43163);
nor U45672 (N_45672,N_43859,N_40216);
nor U45673 (N_45673,N_44601,N_43520);
or U45674 (N_45674,N_43042,N_43220);
or U45675 (N_45675,N_41897,N_43755);
and U45676 (N_45676,N_44882,N_42558);
or U45677 (N_45677,N_42300,N_42658);
nor U45678 (N_45678,N_40059,N_44973);
or U45679 (N_45679,N_43724,N_41304);
xnor U45680 (N_45680,N_44052,N_43952);
or U45681 (N_45681,N_42410,N_41563);
or U45682 (N_45682,N_41108,N_44300);
nor U45683 (N_45683,N_40481,N_43692);
nand U45684 (N_45684,N_44559,N_42942);
or U45685 (N_45685,N_43615,N_43959);
or U45686 (N_45686,N_41357,N_41554);
xor U45687 (N_45687,N_43743,N_40488);
nand U45688 (N_45688,N_42156,N_42538);
nand U45689 (N_45689,N_42718,N_41386);
nor U45690 (N_45690,N_42239,N_41726);
and U45691 (N_45691,N_40844,N_43428);
and U45692 (N_45692,N_44661,N_41135);
and U45693 (N_45693,N_40343,N_40783);
xnor U45694 (N_45694,N_40444,N_44423);
nor U45695 (N_45695,N_40678,N_44468);
or U45696 (N_45696,N_42046,N_44522);
xor U45697 (N_45697,N_43992,N_43638);
and U45698 (N_45698,N_42647,N_43582);
nand U45699 (N_45699,N_41033,N_40832);
and U45700 (N_45700,N_41005,N_42400);
xnor U45701 (N_45701,N_42957,N_42307);
nor U45702 (N_45702,N_44163,N_43023);
and U45703 (N_45703,N_41311,N_43293);
xor U45704 (N_45704,N_42180,N_40550);
xor U45705 (N_45705,N_43848,N_40749);
and U45706 (N_45706,N_43301,N_40452);
and U45707 (N_45707,N_40694,N_41409);
nand U45708 (N_45708,N_42897,N_40971);
xor U45709 (N_45709,N_40009,N_44691);
nand U45710 (N_45710,N_43012,N_44167);
nor U45711 (N_45711,N_43435,N_41195);
xor U45712 (N_45712,N_43171,N_44857);
nand U45713 (N_45713,N_44419,N_44713);
or U45714 (N_45714,N_42739,N_44929);
nor U45715 (N_45715,N_40901,N_42990);
nor U45716 (N_45716,N_42695,N_44626);
and U45717 (N_45717,N_41085,N_42337);
and U45718 (N_45718,N_44535,N_42639);
nand U45719 (N_45719,N_40254,N_41121);
nor U45720 (N_45720,N_40266,N_44263);
and U45721 (N_45721,N_41762,N_41934);
or U45722 (N_45722,N_42747,N_40546);
and U45723 (N_45723,N_44593,N_43182);
xnor U45724 (N_45724,N_42383,N_41919);
or U45725 (N_45725,N_44188,N_44103);
nor U45726 (N_45726,N_44016,N_40114);
nor U45727 (N_45727,N_41975,N_42981);
and U45728 (N_45728,N_42719,N_43889);
or U45729 (N_45729,N_41815,N_43110);
nand U45730 (N_45730,N_40572,N_40044);
and U45731 (N_45731,N_40756,N_40591);
and U45732 (N_45732,N_44955,N_40703);
or U45733 (N_45733,N_42067,N_43850);
xnor U45734 (N_45734,N_40855,N_42253);
xor U45735 (N_45735,N_43517,N_42177);
or U45736 (N_45736,N_42304,N_42261);
nand U45737 (N_45737,N_40631,N_44743);
nor U45738 (N_45738,N_44529,N_42881);
or U45739 (N_45739,N_41746,N_42133);
or U45740 (N_45740,N_41620,N_42510);
and U45741 (N_45741,N_44176,N_43377);
and U45742 (N_45742,N_42365,N_40992);
xor U45743 (N_45743,N_43907,N_42151);
and U45744 (N_45744,N_41095,N_43297);
nand U45745 (N_45745,N_41907,N_40248);
or U45746 (N_45746,N_42172,N_43753);
xnor U45747 (N_45747,N_41602,N_40278);
or U45748 (N_45748,N_42677,N_44046);
nor U45749 (N_45749,N_44672,N_40401);
or U45750 (N_45750,N_40284,N_44317);
xnor U45751 (N_45751,N_43123,N_41583);
xor U45752 (N_45752,N_43510,N_43363);
nand U45753 (N_45753,N_41785,N_42474);
and U45754 (N_45754,N_41860,N_44228);
nor U45755 (N_45755,N_41399,N_42594);
and U45756 (N_45756,N_44220,N_44507);
nand U45757 (N_45757,N_42111,N_42928);
or U45758 (N_45758,N_40555,N_44192);
nor U45759 (N_45759,N_40660,N_44253);
or U45760 (N_45760,N_40935,N_40078);
or U45761 (N_45761,N_43286,N_43020);
nor U45762 (N_45762,N_44753,N_42049);
or U45763 (N_45763,N_40760,N_41116);
nand U45764 (N_45764,N_44833,N_41615);
or U45765 (N_45765,N_41144,N_40559);
nand U45766 (N_45766,N_42625,N_40294);
xor U45767 (N_45767,N_43776,N_43484);
xor U45768 (N_45768,N_42123,N_43426);
or U45769 (N_45769,N_40997,N_40795);
xor U45770 (N_45770,N_41506,N_40940);
or U45771 (N_45771,N_42137,N_44924);
nand U45772 (N_45772,N_42014,N_41455);
or U45773 (N_45773,N_41071,N_41597);
and U45774 (N_45774,N_44793,N_42005);
nor U45775 (N_45775,N_42168,N_43344);
nand U45776 (N_45776,N_43267,N_40882);
xnor U45777 (N_45777,N_40511,N_44384);
or U45778 (N_45778,N_41881,N_43529);
nor U45779 (N_45779,N_42465,N_41467);
xnor U45780 (N_45780,N_43281,N_44965);
nand U45781 (N_45781,N_40326,N_44042);
nor U45782 (N_45782,N_41221,N_41580);
nand U45783 (N_45783,N_43223,N_42588);
nand U45784 (N_45784,N_40450,N_43751);
nor U45785 (N_45785,N_44557,N_44940);
xor U45786 (N_45786,N_41968,N_43673);
nand U45787 (N_45787,N_40348,N_41608);
nand U45788 (N_45788,N_43302,N_42672);
or U45789 (N_45789,N_41541,N_41281);
xnor U45790 (N_45790,N_44201,N_44101);
and U45791 (N_45791,N_44508,N_40964);
xor U45792 (N_45792,N_42917,N_44392);
and U45793 (N_45793,N_41501,N_44893);
and U45794 (N_45794,N_40794,N_40891);
nand U45795 (N_45795,N_41187,N_44996);
and U45796 (N_45796,N_42685,N_40646);
and U45797 (N_45797,N_40677,N_43839);
nand U45798 (N_45798,N_42110,N_41240);
or U45799 (N_45799,N_43146,N_42327);
xnor U45800 (N_45800,N_44688,N_40510);
or U45801 (N_45801,N_40637,N_43371);
nor U45802 (N_45802,N_41266,N_42667);
nand U45803 (N_45803,N_44358,N_44813);
nand U45804 (N_45804,N_44444,N_43666);
and U45805 (N_45805,N_40893,N_42279);
nor U45806 (N_45806,N_44902,N_44407);
nor U45807 (N_45807,N_44563,N_40600);
xor U45808 (N_45808,N_41585,N_40588);
nand U45809 (N_45809,N_41591,N_41444);
nor U45810 (N_45810,N_44580,N_42448);
xnor U45811 (N_45811,N_43698,N_42482);
or U45812 (N_45812,N_40318,N_40264);
and U45813 (N_45813,N_41727,N_41010);
and U45814 (N_45814,N_43551,N_42834);
nand U45815 (N_45815,N_42213,N_44460);
nor U45816 (N_45816,N_40829,N_44819);
nor U45817 (N_45817,N_42409,N_40409);
or U45818 (N_45818,N_42004,N_43266);
xnor U45819 (N_45819,N_40385,N_44091);
nor U45820 (N_45820,N_41657,N_44480);
and U45821 (N_45821,N_42075,N_44659);
and U45822 (N_45822,N_40002,N_44831);
xnor U45823 (N_45823,N_43008,N_40304);
and U45824 (N_45824,N_44974,N_43682);
xor U45825 (N_45825,N_41325,N_40107);
xnor U45826 (N_45826,N_44014,N_41767);
or U45827 (N_45827,N_44573,N_42057);
xnor U45828 (N_45828,N_41061,N_44285);
xor U45829 (N_45829,N_42045,N_40627);
nor U45830 (N_45830,N_42086,N_43677);
nand U45831 (N_45831,N_41457,N_44649);
and U45832 (N_45832,N_42492,N_42694);
and U45833 (N_45833,N_42175,N_42235);
nand U45834 (N_45834,N_40330,N_40934);
xor U45835 (N_45835,N_41292,N_44120);
xnor U45836 (N_45836,N_40058,N_41829);
nor U45837 (N_45837,N_41644,N_41397);
nor U45838 (N_45838,N_44497,N_41048);
or U45839 (N_45839,N_40126,N_44796);
or U45840 (N_45840,N_41814,N_41616);
nand U45841 (N_45841,N_42299,N_40352);
xnor U45842 (N_45842,N_43919,N_44837);
and U45843 (N_45843,N_43034,N_43936);
and U45844 (N_45844,N_40183,N_44074);
xnor U45845 (N_45845,N_40329,N_43153);
nor U45846 (N_45846,N_42104,N_44817);
or U45847 (N_45847,N_40902,N_40585);
nor U45848 (N_45848,N_40268,N_44019);
nor U45849 (N_45849,N_43860,N_44610);
nor U45850 (N_45850,N_41035,N_43440);
nand U45851 (N_45851,N_40870,N_43528);
or U45852 (N_45852,N_41161,N_44205);
nand U45853 (N_45853,N_43656,N_43479);
nand U45854 (N_45854,N_42136,N_43081);
or U45855 (N_45855,N_40487,N_42545);
nand U45856 (N_45856,N_43148,N_40975);
nand U45857 (N_45857,N_43063,N_41710);
xor U45858 (N_45858,N_41307,N_43661);
xnor U45859 (N_45859,N_42577,N_40359);
nor U45860 (N_45860,N_41337,N_40390);
xor U45861 (N_45861,N_44612,N_41956);
nor U45862 (N_45862,N_44105,N_41413);
and U45863 (N_45863,N_41385,N_41074);
nor U45864 (N_45864,N_43489,N_42977);
nand U45865 (N_45865,N_43397,N_40592);
nand U45866 (N_45866,N_41565,N_43002);
and U45867 (N_45867,N_40387,N_43420);
or U45868 (N_45868,N_44824,N_41171);
xnor U45869 (N_45869,N_41344,N_40377);
nand U45870 (N_45870,N_42682,N_40057);
nand U45871 (N_45871,N_43032,N_41093);
xor U45872 (N_45872,N_44678,N_43806);
xor U45873 (N_45873,N_40568,N_40869);
xnor U45874 (N_45874,N_44080,N_44408);
or U45875 (N_45875,N_40713,N_43901);
nand U45876 (N_45876,N_43443,N_40449);
and U45877 (N_45877,N_40537,N_41846);
nor U45878 (N_45878,N_40188,N_41808);
or U45879 (N_45879,N_42097,N_42720);
xnor U45880 (N_45880,N_40980,N_40863);
or U45881 (N_45881,N_41920,N_41298);
xnor U45882 (N_45882,N_42373,N_43041);
xnor U45883 (N_45883,N_42624,N_43395);
xnor U45884 (N_45884,N_42602,N_44912);
or U45885 (N_45885,N_43664,N_44966);
nor U45886 (N_45886,N_40373,N_43016);
nor U45887 (N_45887,N_44168,N_43468);
nand U45888 (N_45888,N_41136,N_43612);
nor U45889 (N_45889,N_41753,N_42478);
xor U45890 (N_45890,N_44001,N_40369);
nand U45891 (N_45891,N_40516,N_42952);
nor U45892 (N_45892,N_40615,N_44802);
xor U45893 (N_45893,N_40172,N_42617);
nand U45894 (N_45894,N_44462,N_43581);
nor U45895 (N_45895,N_43794,N_40419);
and U45896 (N_45896,N_44122,N_41216);
xor U45897 (N_45897,N_43928,N_43455);
xnor U45898 (N_45898,N_43161,N_43926);
or U45899 (N_45899,N_42247,N_44202);
nand U45900 (N_45900,N_43003,N_42578);
or U45901 (N_45901,N_40344,N_41200);
or U45902 (N_45902,N_43844,N_44037);
xor U45903 (N_45903,N_40362,N_40895);
or U45904 (N_45904,N_44714,N_43620);
nor U45905 (N_45905,N_43060,N_41654);
nand U45906 (N_45906,N_43565,N_44108);
nand U45907 (N_45907,N_43115,N_43949);
and U45908 (N_45908,N_43525,N_43174);
and U45909 (N_45909,N_40074,N_43521);
nor U45910 (N_45910,N_43900,N_43562);
or U45911 (N_45911,N_41618,N_44881);
nand U45912 (N_45912,N_42912,N_44461);
xnor U45913 (N_45913,N_40448,N_41633);
and U45914 (N_45914,N_41064,N_43497);
or U45915 (N_45915,N_44717,N_44908);
and U45916 (N_45916,N_44050,N_44068);
nand U45917 (N_45917,N_40429,N_42392);
or U45918 (N_45918,N_44112,N_41394);
xnor U45919 (N_45919,N_40876,N_42495);
or U45920 (N_45920,N_42131,N_44598);
or U45921 (N_45921,N_44000,N_40851);
xnor U45922 (N_45922,N_40954,N_42480);
or U45923 (N_45923,N_42877,N_43460);
nand U45924 (N_45924,N_41801,N_44501);
and U45925 (N_45925,N_41439,N_40880);
or U45926 (N_45926,N_41513,N_41464);
nand U45927 (N_45927,N_42761,N_44217);
nand U45928 (N_45928,N_40297,N_42488);
xnor U45929 (N_45929,N_40253,N_44801);
nand U45930 (N_45930,N_43946,N_40213);
xor U45931 (N_45931,N_43829,N_40692);
nor U45932 (N_45932,N_43476,N_44894);
and U45933 (N_45933,N_44673,N_41724);
xor U45934 (N_45934,N_42141,N_42339);
nand U45935 (N_45935,N_41614,N_44106);
or U45936 (N_45936,N_42424,N_43637);
or U45937 (N_45937,N_42378,N_42633);
xor U45938 (N_45938,N_43818,N_42372);
xor U45939 (N_45939,N_42205,N_44685);
or U45940 (N_45940,N_44749,N_41790);
or U45941 (N_45941,N_41786,N_42027);
nand U45942 (N_45942,N_43247,N_41553);
or U45943 (N_45943,N_43688,N_41117);
nand U45944 (N_45944,N_40479,N_42754);
or U45945 (N_45945,N_44137,N_41915);
and U45946 (N_45946,N_43450,N_42353);
nand U45947 (N_45947,N_40014,N_41712);
nand U45948 (N_45948,N_43597,N_40464);
xnor U45949 (N_45949,N_41469,N_40007);
and U45950 (N_45950,N_40715,N_41955);
nor U45951 (N_45951,N_40001,N_43548);
or U45952 (N_45952,N_42869,N_40407);
or U45953 (N_45953,N_41180,N_44250);
nor U45954 (N_45954,N_44960,N_40624);
or U45955 (N_45955,N_44172,N_41795);
nand U45956 (N_45956,N_44198,N_42413);
xnor U45957 (N_45957,N_42248,N_44899);
or U45958 (N_45958,N_43979,N_44584);
nor U45959 (N_45959,N_44901,N_42599);
nor U45960 (N_45960,N_42164,N_40973);
nand U45961 (N_45961,N_42395,N_41405);
and U45962 (N_45962,N_42829,N_41568);
nor U45963 (N_45963,N_41206,N_41493);
xnor U45964 (N_45964,N_44980,N_41097);
xnor U45965 (N_45965,N_40315,N_40370);
or U45966 (N_45966,N_44269,N_41999);
nor U45967 (N_45967,N_42303,N_40336);
or U45968 (N_45968,N_41592,N_42419);
nor U45969 (N_45969,N_41203,N_42216);
nand U45970 (N_45970,N_43648,N_44095);
and U45971 (N_45971,N_44864,N_40643);
xor U45972 (N_45972,N_42457,N_42791);
or U45973 (N_45973,N_42626,N_41607);
and U45974 (N_45974,N_42453,N_40333);
nor U45975 (N_45975,N_42237,N_41448);
and U45976 (N_45976,N_43256,N_40083);
and U45977 (N_45977,N_44656,N_41838);
nand U45978 (N_45978,N_41065,N_44036);
xor U45979 (N_45979,N_43492,N_42427);
or U45980 (N_45980,N_43410,N_41536);
nor U45981 (N_45981,N_41828,N_44174);
and U45982 (N_45982,N_44204,N_41571);
xor U45983 (N_45983,N_43511,N_44511);
xor U45984 (N_45984,N_44318,N_43831);
or U45985 (N_45985,N_43554,N_43619);
nor U45986 (N_45986,N_42817,N_44548);
nand U45987 (N_45987,N_41935,N_40113);
or U45988 (N_45988,N_42098,N_42551);
or U45989 (N_45989,N_40822,N_44089);
nor U45990 (N_45990,N_41485,N_41957);
nand U45991 (N_45991,N_42055,N_41451);
or U45992 (N_45992,N_42721,N_43629);
or U45993 (N_45993,N_44093,N_41787);
nor U45994 (N_45994,N_40791,N_41152);
or U45995 (N_45995,N_42002,N_40701);
xor U45996 (N_45996,N_43989,N_40477);
nor U45997 (N_45997,N_40012,N_41931);
nand U45998 (N_45998,N_44862,N_41051);
or U45999 (N_45999,N_40476,N_44327);
nor U46000 (N_46000,N_43378,N_43217);
or U46001 (N_46001,N_43775,N_40517);
nor U46002 (N_46002,N_42796,N_42149);
or U46003 (N_46003,N_41432,N_43618);
and U46004 (N_46004,N_44338,N_44443);
nor U46005 (N_46005,N_44326,N_42961);
nor U46006 (N_46006,N_43073,N_43935);
and U46007 (N_46007,N_42936,N_40006);
nor U46008 (N_46008,N_41854,N_40651);
or U46009 (N_46009,N_42404,N_43113);
and U46010 (N_46010,N_41151,N_43380);
xor U46011 (N_46011,N_42256,N_40231);
xor U46012 (N_46012,N_41927,N_43411);
nand U46013 (N_46013,N_43280,N_40852);
xor U46014 (N_46014,N_41091,N_44427);
nand U46015 (N_46015,N_44603,N_40349);
and U46016 (N_46016,N_42949,N_43964);
nor U46017 (N_46017,N_44495,N_41888);
xnor U46018 (N_46018,N_41480,N_40174);
or U46019 (N_46019,N_44500,N_41653);
nor U46020 (N_46020,N_41599,N_43707);
or U46021 (N_46021,N_41896,N_40970);
nor U46022 (N_46022,N_40305,N_41521);
or U46023 (N_46023,N_42323,N_40655);
nand U46024 (N_46024,N_44909,N_42290);
and U46025 (N_46025,N_43224,N_41193);
nand U46026 (N_46026,N_40565,N_44554);
or U46027 (N_46027,N_44547,N_44832);
nor U46028 (N_46028,N_42975,N_40273);
nor U46029 (N_46029,N_41465,N_41214);
xnor U46030 (N_46030,N_44144,N_43349);
nand U46031 (N_46031,N_43826,N_42062);
and U46032 (N_46032,N_42001,N_42421);
xor U46033 (N_46033,N_44448,N_41418);
and U46034 (N_46034,N_40428,N_42678);
and U46035 (N_46035,N_40232,N_43805);
and U46036 (N_46036,N_43295,N_40793);
nor U46037 (N_46037,N_44179,N_43678);
nand U46038 (N_46038,N_40823,N_40589);
nand U46039 (N_46039,N_41251,N_41917);
and U46040 (N_46040,N_41026,N_42052);
or U46041 (N_46041,N_41672,N_42461);
xnor U46042 (N_46042,N_44814,N_40000);
or U46043 (N_46043,N_44513,N_41807);
nand U46044 (N_46044,N_41228,N_44885);
nor U46045 (N_46045,N_43075,N_44687);
and U46046 (N_46046,N_41458,N_40207);
nor U46047 (N_46047,N_41851,N_41689);
xor U46048 (N_46048,N_43011,N_44835);
xnor U46049 (N_46049,N_42257,N_40763);
or U46050 (N_46050,N_43434,N_44489);
nand U46051 (N_46051,N_42351,N_43546);
and U46052 (N_46052,N_44884,N_44859);
or U46053 (N_46053,N_42613,N_42989);
xor U46054 (N_46054,N_42927,N_41550);
nand U46055 (N_46055,N_41784,N_41482);
or U46056 (N_46056,N_43304,N_42025);
and U46057 (N_46057,N_43307,N_44387);
or U46058 (N_46058,N_44807,N_40280);
nand U46059 (N_46059,N_44991,N_43208);
nor U46060 (N_46060,N_44433,N_44297);
nand U46061 (N_46061,N_41222,N_43924);
nor U46062 (N_46062,N_43458,N_40948);
or U46063 (N_46063,N_43685,N_41239);
xnor U46064 (N_46064,N_40120,N_44356);
and U46065 (N_46065,N_43021,N_41617);
nor U46066 (N_46066,N_40621,N_44738);
and U46067 (N_46067,N_40881,N_44583);
or U46068 (N_46068,N_44346,N_44096);
nor U46069 (N_46069,N_40356,N_41636);
nor U46070 (N_46070,N_43033,N_41964);
nor U46071 (N_46071,N_41054,N_44207);
nor U46072 (N_46072,N_41709,N_43970);
nor U46073 (N_46073,N_41273,N_44374);
or U46074 (N_46074,N_43205,N_42030);
nor U46075 (N_46075,N_42350,N_44726);
xnor U46076 (N_46076,N_40802,N_40309);
nor U46077 (N_46077,N_41548,N_41013);
or U46078 (N_46078,N_40717,N_42142);
nor U46079 (N_46079,N_40291,N_41515);
or U46080 (N_46080,N_40986,N_40209);
and U46081 (N_46081,N_42003,N_44938);
nand U46082 (N_46082,N_42816,N_41974);
nor U46083 (N_46083,N_40540,N_40836);
nand U46084 (N_46084,N_40158,N_44629);
and U46085 (N_46085,N_40117,N_41538);
xor U46086 (N_46086,N_40628,N_41502);
nand U46087 (N_46087,N_43947,N_42513);
xnor U46088 (N_46088,N_40239,N_44067);
or U46089 (N_46089,N_42925,N_44224);
and U46090 (N_46090,N_42388,N_42040);
and U46091 (N_46091,N_41667,N_41424);
xor U46092 (N_46092,N_42666,N_43053);
nor U46093 (N_46093,N_40134,N_40495);
xnor U46094 (N_46094,N_42673,N_42539);
xor U46095 (N_46095,N_44304,N_40892);
or U46096 (N_46096,N_44082,N_42399);
and U46097 (N_46097,N_42609,N_43298);
or U46098 (N_46098,N_43409,N_41293);
or U46099 (N_46099,N_41704,N_41741);
xor U46100 (N_46100,N_44132,N_44932);
nand U46101 (N_46101,N_43771,N_41249);
xor U46102 (N_46102,N_42485,N_40421);
nor U46103 (N_46103,N_44939,N_41384);
nor U46104 (N_46104,N_44998,N_44706);
nor U46105 (N_46105,N_43526,N_41516);
and U46106 (N_46106,N_42125,N_44765);
xnor U46107 (N_46107,N_41965,N_43381);
nor U46108 (N_46108,N_43693,N_40564);
and U46109 (N_46109,N_43555,N_44260);
or U46110 (N_46110,N_42848,N_42924);
nor U46111 (N_46111,N_42836,N_41750);
and U46112 (N_46112,N_40169,N_40149);
or U46113 (N_46113,N_43817,N_40451);
or U46114 (N_46114,N_44791,N_41299);
or U46115 (N_46115,N_41389,N_43874);
or U46116 (N_46116,N_42195,N_41114);
nor U46117 (N_46117,N_42520,N_42697);
or U46118 (N_46118,N_44954,N_43543);
nand U46119 (N_46119,N_43832,N_42724);
nand U46120 (N_46120,N_41745,N_43014);
nor U46121 (N_46121,N_44141,N_42408);
nand U46122 (N_46122,N_40018,N_40680);
nand U46123 (N_46123,N_43351,N_43777);
or U46124 (N_46124,N_41339,N_41998);
nand U46125 (N_46125,N_43250,N_41634);
nand U46126 (N_46126,N_42119,N_43225);
and U46127 (N_46127,N_41584,N_40731);
and U46128 (N_46128,N_43258,N_43849);
nand U46129 (N_46129,N_41256,N_41845);
xor U46130 (N_46130,N_40561,N_44771);
nor U46131 (N_46131,N_44215,N_40223);
and U46132 (N_46132,N_44946,N_40067);
or U46133 (N_46133,N_44643,N_41669);
nor U46134 (N_46134,N_42862,N_42984);
nor U46135 (N_46135,N_42309,N_40688);
and U46136 (N_46136,N_41701,N_40194);
and U46137 (N_46137,N_41219,N_40991);
xor U46138 (N_46138,N_43737,N_41546);
or U46139 (N_46139,N_40215,N_40438);
or U46140 (N_46140,N_44565,N_44919);
and U46141 (N_46141,N_44355,N_44746);
xnor U46142 (N_46142,N_43124,N_44475);
nor U46143 (N_46143,N_43963,N_40077);
xnor U46144 (N_46144,N_40245,N_42082);
and U46145 (N_46145,N_43037,N_40296);
nor U46146 (N_46146,N_41868,N_40242);
nor U46147 (N_46147,N_42651,N_42108);
nand U46148 (N_46148,N_43055,N_41520);
or U46149 (N_46149,N_43749,N_41462);
or U46150 (N_46150,N_44611,N_42061);
nand U46151 (N_46151,N_42648,N_42187);
nor U46152 (N_46152,N_40226,N_42065);
and U46153 (N_46153,N_43337,N_44034);
or U46154 (N_46154,N_43089,N_44875);
and U46155 (N_46155,N_42693,N_43559);
and U46156 (N_46156,N_43017,N_40190);
or U46157 (N_46157,N_44957,N_41272);
nor U46158 (N_46158,N_41898,N_41390);
and U46159 (N_46159,N_40478,N_43334);
nor U46160 (N_46160,N_42593,N_44838);
and U46161 (N_46161,N_43494,N_43006);
xor U46162 (N_46162,N_40865,N_41757);
and U46163 (N_46163,N_43039,N_42531);
and U46164 (N_46164,N_42356,N_41719);
or U46165 (N_46165,N_41332,N_41596);
nor U46166 (N_46166,N_43018,N_40413);
nand U46167 (N_46167,N_42553,N_43834);
or U46168 (N_46168,N_42029,N_40738);
nor U46169 (N_46169,N_40179,N_41335);
or U46170 (N_46170,N_42544,N_40465);
and U46171 (N_46171,N_42170,N_40894);
nor U46172 (N_46172,N_44897,N_42430);
xor U46173 (N_46173,N_40679,N_42068);
nor U46174 (N_46174,N_43214,N_40849);
nor U46175 (N_46175,N_43892,N_40350);
nand U46176 (N_46176,N_44869,N_43417);
or U46177 (N_46177,N_43178,N_40932);
nor U46178 (N_46178,N_43401,N_43762);
nor U46179 (N_46179,N_42477,N_42687);
and U46180 (N_46180,N_42158,N_44759);
nand U46181 (N_46181,N_43333,N_41863);
nand U46182 (N_46182,N_42620,N_43087);
nor U46183 (N_46183,N_42973,N_44934);
or U46184 (N_46184,N_44375,N_42047);
xor U46185 (N_46185,N_44482,N_40856);
and U46186 (N_46186,N_43483,N_44947);
and U46187 (N_46187,N_43140,N_42814);
and U46188 (N_46188,N_43169,N_40115);
nand U46189 (N_46189,N_42674,N_44666);
or U46190 (N_46190,N_41754,N_43758);
nand U46191 (N_46191,N_43568,N_40725);
and U46192 (N_46192,N_42454,N_41880);
nor U46193 (N_46193,N_44340,N_40944);
nor U46194 (N_46194,N_42063,N_42699);
nand U46195 (N_46195,N_42084,N_44847);
or U46196 (N_46196,N_44437,N_40595);
nand U46197 (N_46197,N_40100,N_42116);
nor U46198 (N_46198,N_41210,N_43603);
nor U46199 (N_46199,N_41913,N_40290);
or U46200 (N_46200,N_43542,N_41628);
and U46201 (N_46201,N_43004,N_40418);
xnor U46202 (N_46202,N_41044,N_40069);
and U46203 (N_46203,N_40032,N_41328);
or U46204 (N_46204,N_42995,N_44347);
nand U46205 (N_46205,N_44693,N_43090);
or U46206 (N_46206,N_40744,N_43819);
or U46207 (N_46207,N_42529,N_41050);
and U46208 (N_46208,N_41798,N_41519);
nand U46209 (N_46209,N_40807,N_43742);
or U46210 (N_46210,N_41638,N_42034);
and U46211 (N_46211,N_41446,N_44177);
nand U46212 (N_46212,N_41022,N_43495);
and U46213 (N_46213,N_41685,N_42077);
xor U46214 (N_46214,N_44638,N_43044);
xor U46215 (N_46215,N_42729,N_44870);
nor U46216 (N_46216,N_40518,N_42093);
nor U46217 (N_46217,N_40917,N_44541);
and U46218 (N_46218,N_44360,N_44125);
xnor U46219 (N_46219,N_41053,N_43516);
or U46220 (N_46220,N_40959,N_44013);
nor U46221 (N_46221,N_44993,N_42955);
nand U46222 (N_46222,N_41408,N_41123);
xnor U46223 (N_46223,N_42863,N_43588);
nand U46224 (N_46224,N_43616,N_42502);
nor U46225 (N_46225,N_43650,N_41698);
or U46226 (N_46226,N_41038,N_44941);
and U46227 (N_46227,N_44078,N_42940);
xor U46228 (N_46228,N_42155,N_43896);
nand U46229 (N_46229,N_42033,N_43372);
xnor U46230 (N_46230,N_40723,N_41842);
xnor U46231 (N_46231,N_44657,N_40577);
nor U46232 (N_46232,N_43405,N_41612);
and U46233 (N_46233,N_43158,N_42790);
xor U46234 (N_46234,N_44619,N_44166);
and U46235 (N_46235,N_42411,N_41288);
nor U46236 (N_46236,N_43399,N_44667);
or U46237 (N_46237,N_41265,N_41452);
nand U46238 (N_46238,N_41483,N_40312);
and U46239 (N_46239,N_42203,N_43287);
nor U46240 (N_46240,N_42035,N_42910);
and U46241 (N_46241,N_41882,N_44491);
nor U46242 (N_46242,N_43058,N_42591);
nor U46243 (N_46243,N_43346,N_40497);
nor U46244 (N_46244,N_42847,N_42807);
nor U46245 (N_46245,N_41948,N_40473);
and U46246 (N_46246,N_41512,N_41909);
xnor U46247 (N_46247,N_43481,N_42916);
nor U46248 (N_46248,N_42878,N_43355);
nand U46249 (N_46249,N_41186,N_40071);
or U46250 (N_46250,N_41435,N_41833);
nor U46251 (N_46251,N_40974,N_43701);
xnor U46252 (N_46252,N_43897,N_40195);
or U46253 (N_46253,N_44579,N_42243);
or U46254 (N_46254,N_41130,N_43070);
nor U46255 (N_46255,N_44551,N_44890);
or U46256 (N_46256,N_44154,N_43604);
xor U46257 (N_46257,N_40025,N_44148);
nor U46258 (N_46258,N_40184,N_41300);
nand U46259 (N_46259,N_41542,N_42302);
or U46260 (N_46260,N_43049,N_41723);
nor U46261 (N_46261,N_42793,N_44780);
nor U46262 (N_46262,N_40586,N_41312);
or U46263 (N_46263,N_43359,N_43660);
and U46264 (N_46264,N_43611,N_42943);
xor U46265 (N_46265,N_43662,N_40845);
and U46266 (N_46266,N_42527,N_44086);
or U46267 (N_46267,N_41910,N_44694);
nor U46268 (N_46268,N_43100,N_42504);
nor U46269 (N_46269,N_41246,N_41334);
xnor U46270 (N_46270,N_43671,N_41156);
or U46271 (N_46271,N_41007,N_40573);
or U46272 (N_46272,N_44002,N_44320);
or U46273 (N_46273,N_42464,N_41567);
xor U46274 (N_46274,N_42429,N_42727);
nor U46275 (N_46275,N_41486,N_43168);
nor U46276 (N_46276,N_43931,N_40989);
nand U46277 (N_46277,N_41015,N_44397);
nand U46278 (N_46278,N_40698,N_42194);
and U46279 (N_46279,N_41229,N_40683);
and U46280 (N_46280,N_40332,N_40017);
nor U46281 (N_46281,N_44432,N_42236);
nor U46282 (N_46282,N_44622,N_42766);
and U46283 (N_46283,N_44732,N_43711);
nor U46284 (N_46284,N_44051,N_42630);
and U46285 (N_46285,N_42153,N_43593);
and U46286 (N_46286,N_43437,N_40635);
xor U46287 (N_46287,N_44731,N_40462);
nand U46288 (N_46288,N_42549,N_40096);
nor U46289 (N_46289,N_43613,N_43788);
nand U46290 (N_46290,N_43485,N_40666);
or U46291 (N_46291,N_44090,N_40490);
nand U46292 (N_46292,N_42330,N_44237);
nand U46293 (N_46293,N_41683,N_42643);
nor U46294 (N_46294,N_41056,N_43920);
or U46295 (N_46295,N_43570,N_41504);
and U46296 (N_46296,N_40089,N_44992);
nand U46297 (N_46297,N_40910,N_41102);
nor U46298 (N_46298,N_44445,N_44487);
nor U46299 (N_46299,N_44631,N_42443);
and U46300 (N_46300,N_42813,N_42523);
xnor U46301 (N_46301,N_44240,N_40430);
or U46302 (N_46302,N_41308,N_42566);
or U46303 (N_46303,N_42753,N_42081);
and U46304 (N_46304,N_44438,N_41508);
nor U46305 (N_46305,N_41382,N_43477);
nand U46306 (N_46306,N_42331,N_41496);
or U46307 (N_46307,N_42767,N_44366);
xor U46308 (N_46308,N_43370,N_41781);
and U46309 (N_46309,N_40923,N_43243);
or U46310 (N_46310,N_40872,N_44129);
or U46311 (N_46311,N_41682,N_41813);
and U46312 (N_46312,N_43971,N_40708);
nor U46313 (N_46313,N_40459,N_40325);
or U46314 (N_46314,N_40386,N_44811);
xor U46315 (N_46315,N_41564,N_42612);
and U46316 (N_46316,N_40065,N_44768);
nand U46317 (N_46317,N_41937,N_43427);
and U46318 (N_46318,N_40534,N_43720);
or U46319 (N_46319,N_41361,N_43676);
xor U46320 (N_46320,N_41700,N_43808);
nand U46321 (N_46321,N_43774,N_44553);
nor U46322 (N_46322,N_42262,N_41986);
xnor U46323 (N_46323,N_42358,N_40618);
nor U46324 (N_46324,N_41049,N_41177);
nor U46325 (N_46325,N_43067,N_40458);
and U46326 (N_46326,N_44575,N_41205);
xor U46327 (N_46327,N_41983,N_40088);
nand U46328 (N_46328,N_41645,N_44968);
and U46329 (N_46329,N_44725,N_41472);
xor U46330 (N_46330,N_41914,N_41098);
nor U46331 (N_46331,N_42856,N_41280);
xor U46332 (N_46332,N_44155,N_43503);
xnor U46333 (N_46333,N_40382,N_41853);
nor U46334 (N_46334,N_44145,N_41324);
xor U46335 (N_46335,N_43147,N_42393);
or U46336 (N_46336,N_41373,N_44364);
nor U46337 (N_46337,N_41225,N_43454);
nor U46338 (N_46338,N_43861,N_41014);
or U46339 (N_46339,N_40064,N_40854);
nand U46340 (N_46340,N_42962,N_40123);
xor U46341 (N_46341,N_41843,N_44290);
or U46342 (N_46342,N_42376,N_44359);
and U46343 (N_46343,N_41755,N_44669);
nand U46344 (N_46344,N_42026,N_44844);
xnor U46345 (N_46345,N_44424,N_42446);
nor U46346 (N_46346,N_43531,N_41734);
nand U46347 (N_46347,N_40392,N_43374);
xor U46348 (N_46348,N_42417,N_40374);
xor U46349 (N_46349,N_42079,N_44476);
or U46350 (N_46350,N_41087,N_40139);
nor U46351 (N_46351,N_42420,N_44345);
xor U46352 (N_46352,N_44867,N_41363);
xor U46353 (N_46353,N_40871,N_43986);
nor U46354 (N_46354,N_40691,N_43338);
nor U46355 (N_46355,N_42746,N_42107);
and U46356 (N_46356,N_41759,N_41404);
nor U46357 (N_46357,N_44904,N_43173);
or U46358 (N_46358,N_41688,N_41990);
or U46359 (N_46359,N_44770,N_44722);
nor U46360 (N_46360,N_44143,N_44380);
and U46361 (N_46361,N_43289,N_42618);
nand U46362 (N_46362,N_40026,N_44309);
or U46363 (N_46363,N_40547,N_42312);
and U46364 (N_46364,N_41861,N_43814);
nor U46365 (N_46365,N_44646,N_42740);
nand U46366 (N_46366,N_43967,N_41175);
nand U46367 (N_46367,N_41021,N_43558);
nand U46368 (N_46368,N_41352,N_44915);
nor U46369 (N_46369,N_44065,N_44272);
nor U46370 (N_46370,N_42645,N_44455);
or U46371 (N_46371,N_41362,N_42749);
or U46372 (N_46372,N_44234,N_43944);
nor U46373 (N_46373,N_44070,N_41317);
nor U46374 (N_46374,N_44197,N_42343);
or U46375 (N_46375,N_40607,N_44614);
or U46376 (N_46376,N_44416,N_41823);
nor U46377 (N_46377,N_44395,N_40818);
xnor U46378 (N_46378,N_43523,N_41331);
nor U46379 (N_46379,N_42092,N_42422);
or U46380 (N_46380,N_40311,N_44605);
nor U46381 (N_46381,N_41661,N_43421);
and U46382 (N_46382,N_42777,N_42880);
xnor U46383 (N_46383,N_43922,N_40093);
nor U46384 (N_46384,N_42894,N_42361);
nor U46385 (N_46385,N_40063,N_40999);
nand U46386 (N_46386,N_41572,N_41693);
xnor U46387 (N_46387,N_40384,N_42397);
nand U46388 (N_46388,N_43665,N_43652);
xnor U46389 (N_46389,N_40157,N_40728);
and U46390 (N_46390,N_40233,N_40234);
or U46391 (N_46391,N_42684,N_43757);
xnor U46392 (N_46392,N_42708,N_42868);
nor U46393 (N_46393,N_42102,N_42031);
or U46394 (N_46394,N_41731,N_43856);
or U46395 (N_46395,N_41932,N_43126);
xor U46396 (N_46396,N_40920,N_42557);
or U46397 (N_46397,N_44818,N_43894);
and U46398 (N_46398,N_44733,N_41162);
nand U46399 (N_46399,N_42483,N_44509);
xor U46400 (N_46400,N_41518,N_43681);
nand U46401 (N_46401,N_42742,N_41577);
nand U46402 (N_46402,N_41008,N_41159);
nand U46403 (N_46403,N_40695,N_41333);
nand U46404 (N_46404,N_43244,N_41497);
nor U46405 (N_46405,N_40667,N_43200);
or U46406 (N_46406,N_43948,N_40950);
and U46407 (N_46407,N_42722,N_41305);
nor U46408 (N_46408,N_44223,N_42425);
or U46409 (N_46409,N_42826,N_43164);
nand U46410 (N_46410,N_44436,N_42999);
or U46411 (N_46411,N_43690,N_43125);
xor U46412 (N_46412,N_44783,N_42914);
nor U46413 (N_46413,N_41189,N_40685);
nor U46414 (N_46414,N_42736,N_44999);
nor U46415 (N_46415,N_43291,N_42401);
or U46416 (N_46416,N_44414,N_44564);
nand U46417 (N_46417,N_41003,N_42348);
and U46418 (N_46418,N_44258,N_44295);
or U46419 (N_46419,N_40668,N_42132);
or U46420 (N_46420,N_41590,N_44463);
nand U46421 (N_46421,N_41534,N_40542);
xnor U46422 (N_46422,N_41366,N_41856);
or U46423 (N_46423,N_42657,N_41588);
xnor U46424 (N_46424,N_41806,N_44536);
nand U46425 (N_46425,N_43229,N_43977);
nand U46426 (N_46426,N_40579,N_44568);
and U46427 (N_46427,N_43852,N_44898);
nor U46428 (N_46428,N_41082,N_43837);
xor U46429 (N_46429,N_43277,N_44544);
or U46430 (N_46430,N_42530,N_42843);
or U46431 (N_46431,N_43236,N_44887);
and U46432 (N_46432,N_43215,N_41662);
or U46433 (N_46433,N_41403,N_44072);
nand U46434 (N_46434,N_40265,N_40228);
nand U46435 (N_46435,N_41104,N_40764);
nand U46436 (N_46436,N_42751,N_42515);
nand U46437 (N_46437,N_43317,N_42490);
and U46438 (N_46438,N_43536,N_43502);
nor U46439 (N_46439,N_43863,N_42466);
nor U46440 (N_46440,N_44871,N_40334);
or U46441 (N_46441,N_44403,N_41906);
or U46442 (N_46442,N_41111,N_40405);
nand U46443 (N_46443,N_44303,N_41876);
and U46444 (N_46444,N_41981,N_43578);
xor U46445 (N_46445,N_43712,N_42705);
and U46446 (N_46446,N_40156,N_40533);
nor U46447 (N_46447,N_42319,N_43300);
and U46448 (N_46448,N_44478,N_42841);
and U46449 (N_46449,N_44977,N_44778);
or U46450 (N_46450,N_41258,N_40274);
xnor U46451 (N_46451,N_42771,N_43591);
xor U46452 (N_46452,N_40673,N_42367);
or U46453 (N_46453,N_44719,N_43331);
nor U46454 (N_46454,N_43191,N_41016);
and U46455 (N_46455,N_42641,N_44585);
or U46456 (N_46456,N_43199,N_42208);
xor U46457 (N_46457,N_40148,N_43556);
or U46458 (N_46458,N_40146,N_44927);
xor U46459 (N_46459,N_41655,N_42167);
xnor U46460 (N_46460,N_40474,N_43833);
or U46461 (N_46461,N_44429,N_41164);
xor U46462 (N_46462,N_40205,N_44944);
and U46463 (N_46463,N_44494,N_44763);
xor U46464 (N_46464,N_43853,N_42113);
nor U46465 (N_46465,N_40788,N_40505);
nand U46466 (N_46466,N_41953,N_42845);
nor U46467 (N_46467,N_44988,N_43865);
xor U46468 (N_46468,N_42579,N_43909);
xor U46469 (N_46469,N_43105,N_41336);
xnor U46470 (N_46470,N_42715,N_44009);
nand U46471 (N_46471,N_43054,N_41928);
or U46472 (N_46472,N_42245,N_42655);
nand U46473 (N_46473,N_42668,N_41301);
nor U46474 (N_46474,N_41176,N_40661);
or U46475 (N_46475,N_43254,N_41663);
and U46476 (N_46476,N_40583,N_40532);
nor U46477 (N_46477,N_41887,N_42921);
or U46478 (N_46478,N_42186,N_43747);
nor U46479 (N_46479,N_42292,N_40638);
and U46480 (N_46480,N_44849,N_43466);
nor U46481 (N_46481,N_40803,N_43513);
xnor U46482 (N_46482,N_40981,N_44986);
or U46483 (N_46483,N_43998,N_41420);
xnor U46484 (N_46484,N_40106,N_44162);
or U46485 (N_46485,N_44587,N_43557);
or U46486 (N_46486,N_41046,N_41971);
nand U46487 (N_46487,N_44225,N_43836);
and U46488 (N_46488,N_40780,N_40322);
xor U46489 (N_46489,N_43547,N_44214);
and U46490 (N_46490,N_40499,N_41017);
xnor U46491 (N_46491,N_40707,N_42827);
nor U46492 (N_46492,N_41012,N_43997);
nor U46493 (N_46493,N_43475,N_44851);
nand U46494 (N_46494,N_43283,N_43365);
and U46495 (N_46495,N_41459,N_43095);
xnor U46496 (N_46496,N_40840,N_43025);
and U46497 (N_46497,N_44266,N_40066);
and U46498 (N_46498,N_42028,N_43104);
or U46499 (N_46499,N_43686,N_41890);
nand U46500 (N_46500,N_42514,N_41023);
nor U46501 (N_46501,N_40994,N_41603);
nor U46502 (N_46502,N_41821,N_41991);
nor U46503 (N_46503,N_40659,N_44010);
nor U46504 (N_46504,N_44411,N_40383);
nor U46505 (N_46505,N_40509,N_40022);
and U46506 (N_46506,N_41778,N_41635);
or U46507 (N_46507,N_44822,N_41569);
nand U46508 (N_46508,N_40647,N_44786);
xor U46509 (N_46509,N_40616,N_42456);
nor U46510 (N_46510,N_43961,N_43598);
nand U46511 (N_46511,N_44127,N_40466);
xnor U46512 (N_46512,N_40657,N_43614);
nor U46513 (N_46513,N_42265,N_40674);
xnor U46514 (N_46514,N_41967,N_44658);
and U46515 (N_46515,N_40492,N_42838);
or U46516 (N_46516,N_40016,N_41788);
and U46517 (N_46517,N_43872,N_42130);
and U46518 (N_46518,N_41112,N_41080);
xnor U46519 (N_46519,N_40068,N_44979);
nor U46520 (N_46520,N_43563,N_43453);
nor U46521 (N_46521,N_42559,N_40805);
and U46522 (N_46522,N_44958,N_43184);
or U46523 (N_46523,N_42154,N_42196);
or U46524 (N_46524,N_43939,N_41601);
nor U46525 (N_46525,N_41287,N_42748);
nand U46526 (N_46526,N_43416,N_43446);
nor U46527 (N_46527,N_42432,N_44158);
nor U46528 (N_46528,N_41172,N_42342);
or U46529 (N_46529,N_42775,N_42076);
or U46530 (N_46530,N_43366,N_44434);
and U46531 (N_46531,N_44950,N_43657);
xor U46532 (N_46532,N_40500,N_44503);
nand U46533 (N_46533,N_41613,N_43988);
and U46534 (N_46534,N_43207,N_41429);
xnor U46535 (N_46535,N_43167,N_43431);
nand U46536 (N_46536,N_41668,N_44600);
xnor U46537 (N_46537,N_41549,N_43082);
nand U46538 (N_46538,N_40549,N_40796);
or U46539 (N_46539,N_40354,N_43798);
or U46540 (N_46540,N_40995,N_43010);
or U46541 (N_46541,N_43114,N_42472);
xor U46542 (N_46542,N_41959,N_43884);
and U46543 (N_46543,N_43248,N_44329);
xor U46544 (N_46544,N_42891,N_44648);
xor U46545 (N_46545,N_44280,N_43093);
nor U46546 (N_46546,N_44836,N_40557);
xnor U46547 (N_46547,N_43210,N_41348);
nand U46548 (N_46548,N_44769,N_40709);
xnor U46549 (N_46549,N_43190,N_42517);
nor U46550 (N_46550,N_43480,N_43206);
and U46551 (N_46551,N_40108,N_42452);
or U46552 (N_46552,N_40814,N_40052);
nand U46553 (N_46553,N_40292,N_42313);
or U46554 (N_46554,N_41783,N_42980);
xor U46555 (N_46555,N_42540,N_41412);
or U46556 (N_46556,N_40397,N_40684);
or U46557 (N_46557,N_41575,N_41484);
nor U46558 (N_46558,N_41555,N_44398);
nand U46559 (N_46559,N_41182,N_44962);
nor U46560 (N_46560,N_43500,N_42091);
or U46561 (N_46561,N_41677,N_43975);
or U46562 (N_46562,N_43119,N_40221);
or U46563 (N_46563,N_41656,N_43553);
and U46564 (N_46564,N_41063,N_42628);
nand U46565 (N_46565,N_40119,N_43313);
xnor U46566 (N_46566,N_40412,N_43714);
nor U46567 (N_46567,N_44146,N_44834);
xor U46568 (N_46568,N_44582,N_44426);
nand U46569 (N_46569,N_44098,N_41223);
or U46570 (N_46570,N_42611,N_43186);
and U46571 (N_46571,N_40878,N_40903);
nand U46572 (N_46572,N_42887,N_42714);
nand U46573 (N_46573,N_43622,N_43576);
and U46574 (N_46574,N_40340,N_40358);
nand U46575 (N_46575,N_40431,N_41768);
or U46576 (N_46576,N_42080,N_43389);
and U46577 (N_46577,N_42522,N_42923);
nand U46578 (N_46578,N_42965,N_40388);
and U46579 (N_46579,N_40062,N_42258);
or U46580 (N_46580,N_41598,N_42835);
nand U46581 (N_46581,N_41415,N_43978);
or U46582 (N_46582,N_44252,N_41411);
and U46583 (N_46583,N_43121,N_44916);
nand U46584 (N_46584,N_43733,N_43319);
and U46585 (N_46585,N_44173,N_43310);
xnor U46586 (N_46586,N_43974,N_41664);
nor U46587 (N_46587,N_40603,N_40224);
or U46588 (N_46588,N_41500,N_40957);
or U46589 (N_46589,N_44633,N_42207);
xor U46590 (N_46590,N_44264,N_40599);
nor U46591 (N_46591,N_43828,N_43471);
nand U46592 (N_46592,N_43111,N_43727);
and U46593 (N_46593,N_43425,N_42772);
and U46594 (N_46594,N_43052,N_42321);
nor U46595 (N_46595,N_41625,N_44114);
or U46596 (N_46596,N_44485,N_42506);
nand U46597 (N_46597,N_40993,N_41885);
or U46598 (N_46598,N_40283,N_41736);
xor U46599 (N_46599,N_40947,N_42450);
or U46600 (N_46600,N_42349,N_43118);
and U46601 (N_46601,N_41505,N_42394);
nand U46602 (N_46602,N_40634,N_40494);
nor U46603 (N_46603,N_43419,N_42710);
xor U46604 (N_46604,N_43195,N_42785);
nand U46605 (N_46605,N_44550,N_42250);
and U46606 (N_46606,N_41315,N_40008);
or U46607 (N_46607,N_41423,N_41191);
or U46608 (N_46608,N_43706,N_43268);
nand U46609 (N_46609,N_42576,N_41717);
nand U46610 (N_46610,N_41737,N_44758);
nor U46611 (N_46611,N_42468,N_41358);
xnor U46612 (N_46612,N_43786,N_44134);
nand U46613 (N_46613,N_42251,N_42301);
nand U46614 (N_46614,N_42899,N_41259);
nand U46615 (N_46615,N_41029,N_42269);
nand U46616 (N_46616,N_43738,N_42152);
nand U46617 (N_46617,N_40360,N_40933);
and U46618 (N_46618,N_44417,N_44608);
xnor U46619 (N_46619,N_40519,N_42013);
and U46620 (N_46620,N_42586,N_40739);
or U46621 (N_46621,N_44533,N_40081);
xnor U46622 (N_46622,N_43246,N_43537);
xnor U46623 (N_46623,N_42289,N_43945);
and U46624 (N_46624,N_41849,N_41593);
nand U46625 (N_46625,N_42621,N_43781);
or U46626 (N_46626,N_41037,N_40601);
nor U46627 (N_46627,N_41972,N_43101);
xnor U46628 (N_46628,N_44473,N_42932);
nor U46629 (N_46629,N_40884,N_42166);
nor U46630 (N_46630,N_43009,N_40076);
nor U46631 (N_46631,N_41489,N_42499);
nand U46632 (N_46632,N_40523,N_42587);
and U46633 (N_46633,N_44892,N_40436);
xor U46634 (N_46634,N_43383,N_41684);
nor U46635 (N_46635,N_44543,N_41582);
xor U46636 (N_46636,N_44060,N_42439);
and U46637 (N_46637,N_41491,N_44422);
xnor U46638 (N_46638,N_44775,N_44577);
nor U46639 (N_46639,N_40118,N_43791);
and U46640 (N_46640,N_40740,N_43467);
xnor U46641 (N_46641,N_41556,N_44552);
xnor U46642 (N_46642,N_42193,N_41488);
nor U46643 (N_46643,N_41837,N_42883);
nor U46644 (N_46644,N_44642,N_44412);
nor U46645 (N_46645,N_40672,N_41729);
xor U46646 (N_46646,N_44328,N_44418);
or U46647 (N_46647,N_40562,N_40496);
nor U46648 (N_46648,N_42489,N_43061);
nor U46649 (N_46649,N_44569,N_43857);
and U46650 (N_46650,N_42189,N_42866);
xnor U46651 (N_46651,N_41817,N_40457);
nor U46652 (N_46652,N_44325,N_44751);
nand U46653 (N_46653,N_44674,N_41070);
xor U46654 (N_46654,N_43038,N_42960);
and U46655 (N_46655,N_43910,N_42888);
xnor U46656 (N_46656,N_41158,N_43586);
or U46657 (N_46657,N_43723,N_41060);
nor U46658 (N_46658,N_40306,N_44532);
or U46659 (N_46659,N_42901,N_40368);
and U46660 (N_46660,N_40782,N_43327);
nor U46661 (N_46661,N_41730,N_40319);
or U46662 (N_46662,N_44952,N_40033);
nor U46663 (N_46663,N_43253,N_42209);
and U46664 (N_46664,N_43379,N_44113);
and U46665 (N_46665,N_40916,N_42571);
or U46666 (N_46666,N_43423,N_44064);
xnor U46667 (N_46667,N_42455,N_44041);
nand U46668 (N_46668,N_42147,N_42978);
nand U46669 (N_46669,N_42646,N_40753);
and U46670 (N_46670,N_44617,N_42368);
xnor U46671 (N_46671,N_41660,N_41841);
and U46672 (N_46672,N_40313,N_42143);
nor U46673 (N_46673,N_43129,N_41545);
nand U46674 (N_46674,N_44926,N_40786);
and U46675 (N_46675,N_40144,N_44917);
xor U46676 (N_46676,N_44092,N_43342);
nand U46677 (N_46677,N_41499,N_42920);
xor U46678 (N_46678,N_44261,N_42039);
and U46679 (N_46679,N_43201,N_41139);
xnor U46680 (N_46680,N_41417,N_42449);
or U46681 (N_46681,N_41994,N_42089);
and U46682 (N_46682,N_42215,N_42820);
nand U46683 (N_46683,N_40644,N_40575);
nor U46684 (N_46684,N_42246,N_43356);
nor U46685 (N_46685,N_43414,N_41884);
and U46686 (N_46686,N_41178,N_41637);
xnor U46687 (N_46687,N_42334,N_44609);
or U46688 (N_46688,N_44987,N_43108);
nor U46689 (N_46689,N_42308,N_41377);
and U46690 (N_46690,N_44566,N_43445);
or U46691 (N_46691,N_41253,N_42583);
or U46692 (N_46692,N_41220,N_44918);
and U46693 (N_46693,N_44956,N_44744);
nor U46694 (N_46694,N_42524,N_43312);
nor U46695 (N_46695,N_43504,N_42403);
nand U46696 (N_46696,N_43994,N_41770);
nand U46697 (N_46697,N_43185,N_41878);
xnor U46698 (N_46698,N_44268,N_44363);
nand U46699 (N_46699,N_40979,N_44591);
or U46700 (N_46700,N_42183,N_41573);
nand U46701 (N_46701,N_41912,N_41257);
nor U46702 (N_46702,N_40664,N_42214);
nand U46703 (N_46703,N_42528,N_42786);
or U46704 (N_46704,N_43654,N_44739);
xor U46705 (N_46705,N_44005,N_41799);
or U46706 (N_46706,N_42423,N_43324);
or U46707 (N_46707,N_41995,N_44615);
and U46708 (N_46708,N_44307,N_41099);
or U46709 (N_46709,N_41918,N_42043);
or U46710 (N_46710,N_40734,N_41659);
nor U46711 (N_46711,N_43621,N_44084);
xor U46712 (N_46712,N_43855,N_41708);
or U46713 (N_46713,N_43602,N_44728);
nand U46714 (N_46714,N_41474,N_40978);
nand U46715 (N_46715,N_44208,N_41145);
or U46716 (N_46716,N_44119,N_43881);
and U46717 (N_46717,N_40260,N_43056);
nor U46718 (N_46718,N_42238,N_42099);
xnor U46719 (N_46719,N_43770,N_43703);
nor U46720 (N_46720,N_42853,N_44873);
and U46721 (N_46721,N_40372,N_40406);
and U46722 (N_46722,N_43534,N_41510);
and U46723 (N_46723,N_42732,N_40597);
or U46724 (N_46724,N_44291,N_44493);
and U46725 (N_46725,N_42050,N_40486);
and U46726 (N_46726,N_41345,N_42895);
and U46727 (N_46727,N_40243,N_42997);
xnor U46728 (N_46728,N_40886,N_44734);
and U46729 (N_46729,N_41199,N_40506);
and U46730 (N_46730,N_42974,N_43142);
or U46731 (N_46731,N_44248,N_43019);
nand U46732 (N_46732,N_42776,N_44785);
nor U46733 (N_46733,N_43704,N_44399);
nand U46734 (N_46734,N_42725,N_42202);
nor U46735 (N_46735,N_41503,N_41738);
xnor U46736 (N_46736,N_42554,N_41077);
nand U46737 (N_46737,N_40277,N_44724);
and U46738 (N_46738,N_42991,N_43193);
nand U46739 (N_46739,N_40963,N_41720);
and U46740 (N_46740,N_43735,N_44740);
nor U46741 (N_46741,N_44670,N_40956);
and U46742 (N_46742,N_41728,N_43966);
nand U46743 (N_46743,N_42681,N_41441);
nor U46744 (N_46744,N_44930,N_44853);
or U46745 (N_46745,N_40622,N_42226);
nor U46746 (N_46746,N_42941,N_40338);
nor U46747 (N_46747,N_44157,N_40784);
xor U46748 (N_46748,N_40693,N_41286);
or U46749 (N_46749,N_43731,N_42070);
or U46750 (N_46750,N_40633,N_42679);
nand U46751 (N_46751,N_42951,N_43871);
nand U46752 (N_46752,N_43572,N_43436);
nor U46753 (N_46753,N_42274,N_43051);
and U46754 (N_46754,N_41574,N_41079);
or U46755 (N_46755,N_41236,N_40508);
nor U46756 (N_46756,N_44213,N_42370);
nor U46757 (N_46757,N_44953,N_44243);
nand U46758 (N_46758,N_42121,N_44459);
or U46759 (N_46759,N_44660,N_40455);
xor U46760 (N_46760,N_44038,N_40911);
nand U46761 (N_46761,N_41126,N_44677);
or U46762 (N_46762,N_40998,N_43273);
nand U46763 (N_46763,N_44560,N_41092);
nor U46764 (N_46764,N_40887,N_42272);
xnor U46765 (N_46765,N_42738,N_40423);
xor U46766 (N_46766,N_43024,N_40566);
or U46767 (N_46767,N_44316,N_43934);
and U46768 (N_46768,N_42467,N_40968);
nor U46769 (N_46769,N_43354,N_43820);
nand U46770 (N_46770,N_40091,N_42011);
nand U46771 (N_46771,N_44854,N_43083);
or U46772 (N_46772,N_40598,N_44896);
nand U46773 (N_46773,N_42811,N_41168);
and U46774 (N_46774,N_43573,N_41327);
or U46775 (N_46775,N_42802,N_42831);
xnor U46776 (N_46776,N_42804,N_42569);
nand U46777 (N_46777,N_41929,N_43729);
and U46778 (N_46778,N_40815,N_40367);
nand U46779 (N_46779,N_42174,N_43600);
or U46780 (N_46780,N_43390,N_42412);
and U46781 (N_46781,N_42230,N_43472);
or U46782 (N_46782,N_40073,N_43713);
or U46783 (N_46783,N_44011,N_42712);
or U46784 (N_46784,N_42875,N_41235);
nor U46785 (N_46785,N_40900,N_42750);
and U46786 (N_46786,N_44772,N_41379);
and U46787 (N_46787,N_42221,N_42690);
or U46788 (N_46788,N_44718,N_40938);
nor U46789 (N_46789,N_42434,N_40639);
nor U46790 (N_46790,N_43730,N_43127);
nand U46791 (N_46791,N_42106,N_44534);
nand U46792 (N_46792,N_43913,N_44288);
nor U46793 (N_46793,N_43203,N_40366);
or U46794 (N_46794,N_42134,N_43630);
xor U46795 (N_46795,N_41725,N_42229);
nor U46796 (N_46796,N_40641,N_43498);
xnor U46797 (N_46797,N_41539,N_41619);
nor U46798 (N_46798,N_43583,N_40697);
nor U46799 (N_46799,N_44496,N_43402);
and U46800 (N_46800,N_42072,N_44246);
and U46801 (N_46801,N_42909,N_44827);
nand U46802 (N_46802,N_41586,N_44159);
nor U46803 (N_46803,N_44830,N_42676);
nand U46804 (N_46804,N_41226,N_44135);
xor U46805 (N_46805,N_44007,N_43360);
xnor U46806 (N_46806,N_43367,N_44635);
xor U46807 (N_46807,N_40154,N_43815);
nor U46808 (N_46808,N_42654,N_40827);
xor U46809 (N_46809,N_42023,N_44777);
and U46810 (N_46810,N_40403,N_43515);
xor U46811 (N_46811,N_42642,N_43736);
xnor U46812 (N_46812,N_44800,N_42584);
nand U46813 (N_46813,N_41903,N_44249);
nor U46814 (N_46814,N_44760,N_43728);
nor U46815 (N_46815,N_43422,N_42469);
nand U46816 (N_46816,N_40310,N_41793);
or U46817 (N_46817,N_41650,N_43527);
xnor U46818 (N_46818,N_42241,N_43951);
and U46819 (N_46819,N_42889,N_40658);
xor U46820 (N_46820,N_42683,N_44131);
nand U46821 (N_46821,N_41694,N_44959);
xnor U46822 (N_46822,N_41057,N_42763);
or U46823 (N_46823,N_40625,N_43005);
or U46824 (N_46824,N_44721,N_41321);
xnor U46825 (N_46825,N_40990,N_43154);
or U46826 (N_46826,N_40395,N_44797);
and U46827 (N_46827,N_42379,N_41461);
nand U46828 (N_46828,N_40027,N_44219);
xnor U46829 (N_46829,N_42311,N_40705);
nand U46830 (N_46830,N_41862,N_40776);
and U46831 (N_46831,N_43987,N_40772);
or U46832 (N_46832,N_42148,N_42689);
nor U46833 (N_46833,N_41826,N_40446);
or U46834 (N_46834,N_44846,N_40775);
or U46835 (N_46835,N_41889,N_43628);
nor U46836 (N_46836,N_41440,N_42182);
xor U46837 (N_46837,N_44077,N_42444);
and U46838 (N_46838,N_40612,N_42659);
xnor U46839 (N_46839,N_41247,N_44689);
and U46840 (N_46840,N_41218,N_41692);
nor U46841 (N_46841,N_42893,N_42101);
nor U46842 (N_46842,N_44567,N_44275);
nor U46843 (N_46843,N_42570,N_40949);
xnor U46844 (N_46844,N_41160,N_42948);
xor U46845 (N_46845,N_44681,N_44654);
nand U46846 (N_46846,N_43415,N_40198);
nor U46847 (N_46847,N_42115,N_44029);
nor U46848 (N_46848,N_44293,N_41245);
and U46849 (N_46849,N_44312,N_40316);
and U46850 (N_46850,N_40982,N_44984);
nand U46851 (N_46851,N_43683,N_44369);
xor U46852 (N_46852,N_42907,N_42731);
nor U46853 (N_46853,N_41243,N_42931);
xor U46854 (N_46854,N_43080,N_41094);
and U46855 (N_46855,N_43732,N_41141);
or U46856 (N_46856,N_43539,N_42947);
xor U46857 (N_46857,N_41523,N_43680);
xnor U46858 (N_46858,N_43272,N_40972);
and U46859 (N_46859,N_43933,N_40301);
and U46860 (N_46860,N_43079,N_40327);
nor U46861 (N_46861,N_42160,N_40686);
and U46862 (N_46862,N_42371,N_44193);
nor U46863 (N_46863,N_40530,N_40456);
or U46864 (N_46864,N_40443,N_43739);
nand U46865 (N_46865,N_40258,N_44842);
or U46866 (N_46866,N_44561,N_41835);
xnor U46867 (N_46867,N_41630,N_41533);
xnor U46868 (N_46868,N_40861,N_42589);
xnor U46869 (N_46869,N_44704,N_43610);
nand U46870 (N_46870,N_44586,N_42851);
or U46871 (N_46871,N_43059,N_42512);
nor U46872 (N_46872,N_40189,N_41109);
and U46873 (N_46873,N_42192,N_41153);
xnor U46874 (N_46874,N_42462,N_40482);
nor U46875 (N_46875,N_41900,N_44524);
xnor U46876 (N_46876,N_40128,N_43404);
nand U46877 (N_46877,N_44589,N_43540);
and U46878 (N_46878,N_44570,N_43877);
nand U46879 (N_46879,N_42882,N_40308);
or U46880 (N_46880,N_44308,N_40789);
nand U46881 (N_46881,N_44187,N_42700);
and U46882 (N_46882,N_42534,N_40996);
or U46883 (N_46883,N_41476,N_40545);
nor U46884 (N_46884,N_43584,N_40004);
nand U46885 (N_46885,N_42041,N_44194);
and U46886 (N_46886,N_40378,N_40240);
xnor U46887 (N_46887,N_42305,N_42481);
xnor U46888 (N_46888,N_41980,N_43799);
and U46889 (N_46889,N_42184,N_43212);
and U46890 (N_46890,N_43165,N_43626);
xnor U46891 (N_46891,N_41254,N_41479);
nand U46892 (N_46892,N_40270,N_43282);
nand U46893 (N_46893,N_41032,N_44931);
nand U46894 (N_46894,N_42054,N_41000);
or U46895 (N_46895,N_43858,N_43965);
xor U46896 (N_46896,N_41850,N_43388);
and U46897 (N_46897,N_42285,N_44378);
or U46898 (N_46898,N_43509,N_44349);
and U46899 (N_46899,N_43156,N_44221);
nand U46900 (N_46900,N_42451,N_43326);
nor U46901 (N_46901,N_43306,N_41761);
nor U46902 (N_46902,N_41134,N_44964);
xor U46903 (N_46903,N_43096,N_44488);
or U46904 (N_46904,N_44271,N_40138);
nor U46905 (N_46905,N_42723,N_44695);
or U46906 (N_46906,N_41780,N_43036);
or U46907 (N_46907,N_40817,N_44049);
xor U46908 (N_46908,N_40498,N_40563);
xnor U46909 (N_46909,N_42500,N_43687);
nor U46910 (N_46910,N_40746,N_44302);
xnor U46911 (N_46911,N_41652,N_42805);
or U46912 (N_46912,N_40414,N_41647);
or U46913 (N_46913,N_43204,N_42360);
nor U46914 (N_46914,N_41690,N_42781);
xor U46915 (N_46915,N_44588,N_44006);
or U46916 (N_46916,N_41349,N_41679);
or U46917 (N_46917,N_40636,N_44169);
and U46918 (N_46918,N_40328,N_43029);
nand U46919 (N_46919,N_41949,N_41894);
nor U46920 (N_46920,N_44639,N_40417);
and U46921 (N_46921,N_43031,N_40520);
or U46922 (N_46922,N_44499,N_40461);
or U46923 (N_46923,N_43878,N_43643);
or U46924 (N_46924,N_43601,N_42297);
nand U46925 (N_46925,N_41984,N_41706);
nor U46926 (N_46926,N_42792,N_42078);
nand U46927 (N_46927,N_40966,N_40842);
nand U46928 (N_46928,N_41492,N_42146);
or U46929 (N_46929,N_40222,N_40918);
nand U46930 (N_46930,N_41950,N_40163);
nand U46931 (N_46931,N_44492,N_41941);
and U46932 (N_46932,N_40809,N_43350);
nor U46933 (N_46933,N_44315,N_41641);
nor U46934 (N_46934,N_42803,N_43903);
and U46935 (N_46935,N_41263,N_41527);
nor U46936 (N_46936,N_42915,N_40130);
or U46937 (N_46937,N_44983,N_43462);
nor U46938 (N_46938,N_43715,N_40375);
nor U46939 (N_46939,N_44943,N_40671);
and U46940 (N_46940,N_44558,N_43323);
or U46941 (N_46941,N_43885,N_42318);
nor U46942 (N_46942,N_42874,N_42190);
nor U46943 (N_46943,N_43932,N_44976);
or U46944 (N_46944,N_41665,N_43134);
nor U46945 (N_46945,N_43507,N_44442);
or U46946 (N_46946,N_42946,N_42886);
or U46947 (N_46947,N_42188,N_40642);
nor U46948 (N_46948,N_42779,N_43514);
or U46949 (N_46949,N_43773,N_44420);
or U46950 (N_46950,N_44708,N_43265);
nor U46951 (N_46951,N_43699,N_41062);
xor U46952 (N_46952,N_41356,N_43066);
xnor U46953 (N_46953,N_42733,N_41119);
xnor U46954 (N_46954,N_43954,N_41262);
nand U46955 (N_46955,N_44351,N_41822);
or U46956 (N_46956,N_41118,N_41765);
or U46957 (N_46957,N_43237,N_42574);
or U46958 (N_46958,N_44745,N_43109);
nand U46959 (N_46959,N_43172,N_43332);
xor U46960 (N_46960,N_43769,N_42435);
or U46961 (N_46961,N_43596,N_41194);
nor U46962 (N_46962,N_43803,N_43102);
nand U46963 (N_46963,N_40345,N_42922);
xor U46964 (N_46964,N_40906,N_41019);
xor U46965 (N_46965,N_40645,N_40285);
or U46966 (N_46966,N_41166,N_41275);
and U46967 (N_46967,N_43816,N_43655);
xnor U46968 (N_46968,N_42227,N_41831);
and U46969 (N_46969,N_41224,N_42317);
and U46970 (N_46970,N_43879,N_42328);
xnor U46971 (N_46971,N_41284,N_44921);
nand U46972 (N_46972,N_41059,N_42608);
xnor U46973 (N_46973,N_41076,N_42333);
xnor U46974 (N_46974,N_41866,N_42431);
or U46975 (N_46975,N_40732,N_40151);
nand U46976 (N_46976,N_42929,N_42185);
nor U46977 (N_46977,N_43159,N_40380);
xnor U46978 (N_46978,N_44186,N_42120);
nand U46979 (N_46979,N_44033,N_40298);
and U46980 (N_46980,N_44504,N_41600);
or U46981 (N_46981,N_43973,N_42295);
xor U46982 (N_46982,N_42730,N_42259);
xor U46983 (N_46983,N_41204,N_40463);
xor U46984 (N_46984,N_42242,N_40838);
nor U46985 (N_46985,N_40202,N_40648);
xor U46986 (N_46986,N_41237,N_44452);
or U46987 (N_46987,N_41514,N_42808);
xor U46988 (N_46988,N_41217,N_43133);
nand U46989 (N_46989,N_40907,N_43345);
xnor U46990 (N_46990,N_41313,N_42088);
nand U46991 (N_46991,N_40050,N_44843);
or U46992 (N_46992,N_40914,N_43668);
and U46993 (N_46993,N_40250,N_40787);
or U46994 (N_46994,N_44339,N_42179);
nand U46995 (N_46995,N_40400,N_42696);
xor U46996 (N_46996,N_42970,N_40804);
nor U46997 (N_46997,N_40199,N_44502);
xor U46998 (N_46998,N_40135,N_43194);
nor U46999 (N_46999,N_41610,N_42649);
xor U47000 (N_47000,N_40765,N_40548);
nor U47001 (N_47001,N_41966,N_40042);
xor U47002 (N_47002,N_43441,N_43887);
or U47003 (N_47003,N_44675,N_40984);
nand U47004 (N_47004,N_40085,N_41511);
nor U47005 (N_47005,N_43396,N_43288);
or U47006 (N_47006,N_44164,N_42240);
and U47007 (N_47007,N_43625,N_41747);
and U47008 (N_47008,N_42440,N_40848);
or U47009 (N_47009,N_44848,N_41771);
xnor U47010 (N_47010,N_44684,N_43772);
nand U47011 (N_47011,N_41901,N_42518);
nand U47012 (N_47012,N_41769,N_44283);
xor U47013 (N_47013,N_43530,N_44472);
nand U47014 (N_47014,N_44372,N_40420);
nor U47015 (N_47015,N_44682,N_41282);
nand U47016 (N_47016,N_44348,N_41973);
nor U47017 (N_47017,N_43545,N_42898);
nor U47018 (N_47018,N_41309,N_44458);
nor U47019 (N_47019,N_41810,N_43120);
xor U47020 (N_47020,N_43150,N_41543);
nor U47021 (N_47021,N_43240,N_43617);
and U47022 (N_47022,N_40247,N_43451);
or U47023 (N_47023,N_40602,N_44486);
nor U47024 (N_47024,N_41559,N_44139);
xor U47025 (N_47025,N_42219,N_44707);
nor U47026 (N_47026,N_42275,N_40926);
nand U47027 (N_47027,N_44323,N_42162);
nand U47028 (N_47028,N_42638,N_43635);
xor U47029 (N_47029,N_43940,N_44289);
or U47030 (N_47030,N_42389,N_43835);
xor U47031 (N_47031,N_42112,N_40943);
nor U47032 (N_47032,N_40866,N_42364);
and U47033 (N_47033,N_44235,N_42244);
or U47034 (N_47034,N_43679,N_41758);
xor U47035 (N_47035,N_44750,N_43181);
xnor U47036 (N_47036,N_41892,N_41739);
nand U47037 (N_47037,N_43177,N_41883);
or U47038 (N_47038,N_44239,N_41380);
xor U47039 (N_47039,N_41487,N_40983);
xor U47040 (N_47040,N_43627,N_42484);
xnor U47041 (N_47041,N_42100,N_40720);
or U47042 (N_47042,N_41551,N_41749);
nand U47043 (N_47043,N_40011,N_40435);
nand U47044 (N_47044,N_40767,N_42017);
nor U47045 (N_47045,N_42000,N_41579);
nor U47046 (N_47046,N_40958,N_41993);
or U47047 (N_47047,N_44742,N_43222);
or U47048 (N_47048,N_43328,N_42755);
or U47049 (N_47049,N_42809,N_44715);
xnor U47050 (N_47050,N_43508,N_42799);
nand U47051 (N_47051,N_44720,N_40272);
or U47052 (N_47052,N_43432,N_42741);
or U47053 (N_47053,N_41360,N_44075);
nand U47054 (N_47054,N_43564,N_42969);
or U47055 (N_47055,N_41871,N_41113);
and U47056 (N_47056,N_41197,N_41891);
and U47057 (N_47057,N_43097,N_42117);
and U47058 (N_47058,N_40454,N_40141);
xnor U47059 (N_47059,N_40493,N_44562);
nor U47060 (N_47060,N_44866,N_40445);
nand U47061 (N_47061,N_43995,N_44344);
xor U47062 (N_47062,N_43385,N_40514);
nand U47063 (N_47063,N_44781,N_43574);
nand U47064 (N_47064,N_40915,N_43501);
and U47065 (N_47065,N_40828,N_42497);
nor U47066 (N_47066,N_44705,N_42362);
xor U47067 (N_47067,N_43942,N_44840);
or U47068 (N_47068,N_44761,N_40718);
and U47069 (N_47069,N_41146,N_40168);
nor U47070 (N_47070,N_43950,N_40843);
or U47071 (N_47071,N_41426,N_41622);
nand U47072 (N_47072,N_42486,N_44703);
or U47073 (N_47073,N_40252,N_43309);
nand U47074 (N_47074,N_40160,N_41045);
nand U47075 (N_47075,N_41269,N_44294);
or U47076 (N_47076,N_40800,N_44701);
nand U47077 (N_47077,N_42713,N_43197);
xnor U47078 (N_47078,N_44440,N_43064);
and U47079 (N_47079,N_40921,N_42344);
nand U47080 (N_47080,N_44370,N_41561);
xor U47081 (N_47081,N_41954,N_42473);
and U47082 (N_47082,N_44470,N_41174);
nand U47083 (N_47083,N_41052,N_41951);
xnor U47084 (N_47084,N_43921,N_44799);
and U47085 (N_47085,N_40904,N_40161);
nor U47086 (N_47086,N_41096,N_44276);
xor U47087 (N_47087,N_44231,N_44505);
xor U47088 (N_47088,N_41183,N_44354);
nor U47089 (N_47089,N_44644,N_42341);
nand U47090 (N_47090,N_43393,N_42879);
nand U47091 (N_47091,N_42543,N_41234);
xor U47092 (N_47092,N_44054,N_43718);
and U47093 (N_47093,N_44314,N_44816);
or U47094 (N_47094,N_43823,N_44652);
and U47095 (N_47095,N_42232,N_42756);
or U47096 (N_47096,N_40293,N_44804);
or U47097 (N_47097,N_40841,N_42758);
and U47098 (N_47098,N_44385,N_42022);
and U47099 (N_47099,N_44377,N_40704);
nand U47100 (N_47100,N_42867,N_41732);
and U47101 (N_47101,N_40962,N_44542);
nand U47102 (N_47102,N_44032,N_42083);
and U47103 (N_47103,N_42384,N_42744);
nand U47104 (N_47104,N_40538,N_43103);
xnor U47105 (N_47105,N_44409,N_44107);
xor U47106 (N_47106,N_42864,N_40341);
nand U47107 (N_47107,N_42634,N_42788);
or U47108 (N_47108,N_44184,N_42519);
nor U47109 (N_47109,N_42581,N_44400);
xnor U47110 (N_47110,N_41190,N_43368);
nor U47111 (N_47111,N_44454,N_43838);
xnor U47112 (N_47112,N_43807,N_43099);
and U47113 (N_47113,N_41830,N_43092);
nor U47114 (N_47114,N_40669,N_42635);
nand U47115 (N_47115,N_43672,N_41782);
and U47116 (N_47116,N_42338,N_40977);
nand U47117 (N_47117,N_40752,N_40733);
nand U47118 (N_47118,N_44195,N_43866);
or U47119 (N_47119,N_43176,N_43911);
xor U47120 (N_47120,N_41431,N_43218);
xnor U47121 (N_47121,N_43043,N_41490);
nand U47122 (N_47122,N_40227,N_44876);
and U47123 (N_47123,N_42122,N_44521);
nand U47124 (N_47124,N_41383,N_44456);
nand U47125 (N_47125,N_40826,N_44978);
and U47126 (N_47126,N_43230,N_41820);
nor U47127 (N_47127,N_43567,N_41147);
nor U47128 (N_47128,N_41844,N_41481);
xnor U47129 (N_47129,N_40525,N_43347);
xor U47130 (N_47130,N_41419,N_44756);
xnor U47131 (N_47131,N_41101,N_43904);
nor U47132 (N_47132,N_44410,N_41453);
or U47133 (N_47133,N_42287,N_44607);
nor U47134 (N_47134,N_42048,N_40617);
xnor U47135 (N_47135,N_42604,N_40097);
nand U47136 (N_47136,N_43292,N_40833);
or U47137 (N_47137,N_40109,N_42374);
or U47138 (N_47138,N_42282,N_44540);
nor U47139 (N_47139,N_43463,N_43030);
or U47140 (N_47140,N_44133,N_42703);
nand U47141 (N_47141,N_42798,N_43969);
xor U47142 (N_47142,N_40929,N_44147);
nor U47143 (N_47143,N_44510,N_43792);
nand U47144 (N_47144,N_44465,N_40320);
and U47145 (N_47145,N_43891,N_40730);
xnor U47146 (N_47146,N_40484,N_40060);
or U47147 (N_47147,N_40792,N_41858);
nand U47148 (N_47148,N_40889,N_43740);
nor U47149 (N_47149,N_43139,N_41131);
xnor U47150 (N_47150,N_44526,N_42019);
nor U47151 (N_47151,N_44920,N_41540);
xnor U47152 (N_47152,N_41777,N_40528);
and U47153 (N_47153,N_43512,N_40021);
nor U47154 (N_47154,N_43867,N_43962);
or U47155 (N_47155,N_44788,N_40580);
nand U47156 (N_47156,N_41319,N_42288);
nand U47157 (N_47157,N_44710,N_44971);
nor U47158 (N_47158,N_42071,N_40331);
xor U47159 (N_47159,N_43700,N_44514);
nand U47160 (N_47160,N_44165,N_42278);
or U47161 (N_47161,N_40220,N_44914);
or U47162 (N_47162,N_40079,N_42680);
nand U47163 (N_47163,N_44490,N_42199);
nand U47164 (N_47164,N_41623,N_43780);
nor U47165 (N_47165,N_44886,N_40834);
nor U47166 (N_47166,N_44435,N_41942);
xor U47167 (N_47167,N_43906,N_42600);
nor U47168 (N_47168,N_40039,N_40524);
and U47169 (N_47169,N_40061,N_41792);
and U47170 (N_47170,N_40300,N_43538);
nand U47171 (N_47171,N_43644,N_42254);
nor U47172 (N_47172,N_40031,N_40544);
xor U47173 (N_47173,N_44539,N_44752);
and U47174 (N_47174,N_42592,N_40864);
and U47175 (N_47175,N_42509,N_44702);
nand U47176 (N_47176,N_41989,N_44170);
nand U47177 (N_47177,N_41570,N_43255);
and U47178 (N_47178,N_41066,N_40858);
xnor U47179 (N_47179,N_40706,N_42854);
nand U47180 (N_47180,N_40182,N_43633);
nor U47181 (N_47181,N_43057,N_44185);
nor U47182 (N_47182,N_42900,N_44298);
and U47183 (N_47183,N_43561,N_43899);
nor U47184 (N_47184,N_42503,N_40192);
nand U47185 (N_47185,N_40441,N_43746);
and U47186 (N_47186,N_44191,N_44528);
nand U47187 (N_47187,N_40919,N_43955);
and U47188 (N_47188,N_42475,N_40489);
and U47189 (N_47189,N_42752,N_41395);
and U47190 (N_47190,N_41371,N_42020);
or U47191 (N_47191,N_40675,N_41004);
and U47192 (N_47192,N_40928,N_44321);
nand U47193 (N_47193,N_43854,N_44124);
or U47194 (N_47194,N_40136,N_41018);
or U47195 (N_47195,N_41347,N_42206);
and U47196 (N_47196,N_44911,N_41470);
nand U47197 (N_47197,N_43213,N_42934);
xnor U47198 (N_47198,N_43812,N_42471);
nor U47199 (N_47199,N_43227,N_42533);
and U47200 (N_47200,N_40737,N_42598);
or U47201 (N_47201,N_44982,N_41680);
and U47202 (N_47202,N_40200,N_40137);
nor U47203 (N_47203,N_44415,N_42191);
nand U47204 (N_47204,N_40010,N_40426);
nand U47205 (N_47205,N_43827,N_43106);
nand U47206 (N_47206,N_43241,N_40422);
or U47207 (N_47207,N_42580,N_42556);
or U47208 (N_47208,N_44951,N_43869);
nor U47209 (N_47209,N_40696,N_43575);
nor U47210 (N_47210,N_40404,N_41443);
xor U47211 (N_47211,N_40271,N_44203);
nand U47212 (N_47212,N_43216,N_41192);
xnor U47213 (N_47213,N_40339,N_44900);
or U47214 (N_47214,N_44428,N_41271);
or U47215 (N_47215,N_40553,N_42074);
or U47216 (N_47216,N_41185,N_44257);
and U47217 (N_47217,N_43135,N_43797);
nand U47218 (N_47218,N_42596,N_41002);
and U47219 (N_47219,N_41232,N_42567);
or U47220 (N_47220,N_42985,N_42726);
xnor U47221 (N_47221,N_41699,N_44686);
nand U47222 (N_47222,N_40503,N_43760);
and U47223 (N_47223,N_43917,N_41581);
nand U47224 (N_47224,N_42161,N_44152);
and U47225 (N_47225,N_41944,N_42945);
or U47226 (N_47226,N_44806,N_40535);
and U47227 (N_47227,N_43088,N_42415);
and U47228 (N_47228,N_40036,N_41626);
xor U47229 (N_47229,N_44990,N_44878);
and U47230 (N_47230,N_42375,N_43709);
and U47231 (N_47231,N_40614,N_44576);
and U47232 (N_47232,N_43166,N_41939);
xor U47233 (N_47233,N_41124,N_40770);
and U47234 (N_47234,N_42616,N_41916);
or U47235 (N_47235,N_41227,N_44779);
nand U47236 (N_47236,N_44017,N_41695);
or U47237 (N_47237,N_43077,N_44241);
xor U47238 (N_47238,N_44451,N_43271);
and U47239 (N_47239,N_40570,N_44517);
nor U47240 (N_47240,N_42691,N_44439);
xnor U47241 (N_47241,N_44446,N_44784);
nand U47242 (N_47242,N_44624,N_40711);
nand U47243 (N_47243,N_41267,N_42498);
and U47244 (N_47244,N_41209,N_43519);
or U47245 (N_47245,N_44839,N_40185);
or U47246 (N_47246,N_41847,N_42127);
and U47247 (N_47247,N_41713,N_44787);
or U47248 (N_47248,N_40259,N_41400);
or U47249 (N_47249,N_40175,N_43144);
and U47250 (N_47250,N_44121,N_40785);
nand U47251 (N_47251,N_41867,N_40095);
xor U47252 (N_47252,N_43864,N_41958);
and U47253 (N_47253,N_42575,N_40571);
nor U47254 (N_47254,N_43595,N_44994);
xor U47255 (N_47255,N_40873,N_43590);
nand U47256 (N_47256,N_42416,N_41463);
and U47257 (N_47257,N_44332,N_44466);
nand U47258 (N_47258,N_44396,N_44206);
xnor U47259 (N_47259,N_44945,N_40985);
or U47260 (N_47260,N_44210,N_41609);
xor U47261 (N_47261,N_40874,N_41859);
nor U47262 (N_47262,N_41078,N_41671);
xor U47263 (N_47263,N_43235,N_44254);
nand U47264 (N_47264,N_41196,N_44789);
nor U47265 (N_47265,N_40513,N_41992);
and U47266 (N_47266,N_44464,N_40924);
nor U47267 (N_47267,N_40303,N_40229);
nand U47268 (N_47268,N_43761,N_41073);
and U47269 (N_47269,N_44985,N_43086);
and U47270 (N_47270,N_40939,N_43824);
nand U47271 (N_47271,N_41353,N_44764);
or U47272 (N_47272,N_42135,N_44736);
or U47273 (N_47273,N_43091,N_42064);
nor U47274 (N_47274,N_41184,N_44128);
nand U47275 (N_47275,N_40936,N_42603);
and U47276 (N_47276,N_43196,N_41987);
or U47277 (N_47277,N_40127,N_44236);
nand U47278 (N_47278,N_40665,N_41764);
nor U47279 (N_47279,N_43439,N_43505);
and U47280 (N_47280,N_43493,N_41852);
or U47281 (N_47281,N_41042,N_40140);
and U47282 (N_47282,N_40416,N_44284);
or U47283 (N_47283,N_40771,N_42129);
nand U47284 (N_47284,N_44795,N_41230);
and U47285 (N_47285,N_42582,N_43449);
nor U47286 (N_47286,N_40204,N_41318);
or U47287 (N_47287,N_42139,N_41925);
and U47288 (N_47288,N_41414,N_44178);
or U47289 (N_47289,N_42009,N_43299);
or U47290 (N_47290,N_44578,N_44211);
and U47291 (N_47291,N_43744,N_43691);
nand U47292 (N_47292,N_40155,N_41924);
or U47293 (N_47293,N_40626,N_41744);
xor U47294 (N_47294,N_41350,N_42391);
xor U47295 (N_47295,N_44142,N_44640);
or U47296 (N_47296,N_43341,N_42051);
and U47297 (N_47297,N_42525,N_44027);
xnor U47298 (N_47298,N_42266,N_42336);
nor U47299 (N_47299,N_43695,N_43391);
and U47300 (N_47300,N_41532,N_42908);
and U47301 (N_47301,N_40193,N_40133);
or U47302 (N_47302,N_40831,N_41020);
nand U47303 (N_47303,N_43734,N_41127);
xnor U47304 (N_47304,N_41157,N_43876);
or U47305 (N_47305,N_40132,N_44425);
nor U47306 (N_47306,N_43340,N_43569);
and U47307 (N_47307,N_42656,N_41624);
and U47308 (N_47308,N_44058,N_44277);
nand U47309 (N_47309,N_43316,N_42176);
nand U47310 (N_47310,N_41381,N_44825);
nand U47311 (N_47311,N_44430,N_42800);
and U47312 (N_47312,N_41211,N_44371);
nor U47313 (N_47313,N_44245,N_40379);
nor U47314 (N_47314,N_41244,N_44880);
nand U47315 (N_47315,N_40662,N_43112);
nand U47316 (N_47316,N_42087,N_42326);
nand U47317 (N_47317,N_43228,N_43357);
nor U47318 (N_47318,N_41001,N_44741);
nand U47319 (N_47319,N_42979,N_40879);
and U47320 (N_47320,N_41179,N_41208);
xor U47321 (N_47321,N_41378,N_44730);
nand U47322 (N_47322,N_43532,N_43269);
or U47323 (N_47323,N_40162,N_43587);
and U47324 (N_47324,N_44498,N_44099);
nor U47325 (N_47325,N_44620,N_43914);
nand U47326 (N_47326,N_42704,N_43784);
nand U47327 (N_47327,N_41473,N_43778);
or U47328 (N_47328,N_42774,N_40922);
xor U47329 (N_47329,N_42846,N_41809);
and U47330 (N_47330,N_44278,N_41836);
or U47331 (N_47331,N_41401,N_44989);
nand U47332 (N_47332,N_41877,N_43329);
nor U47333 (N_47333,N_41181,N_40186);
or U47334 (N_47334,N_43880,N_40177);
or U47335 (N_47335,N_40687,N_40187);
or U47336 (N_47336,N_44330,N_42044);
and U47337 (N_47337,N_43284,N_40652);
nand U47338 (N_47338,N_42210,N_43262);
or U47339 (N_47339,N_43915,N_42535);
xnor U47340 (N_47340,N_40774,N_42224);
or U47341 (N_47341,N_43438,N_42114);
xnor U47342 (N_47342,N_40485,N_41407);
xor U47343 (N_47343,N_40262,N_41960);
xor U47344 (N_47344,N_42407,N_42508);
nor U47345 (N_47345,N_42293,N_42280);
xor U47346 (N_47346,N_44388,N_44069);
nand U47347 (N_47347,N_44117,N_40875);
or U47348 (N_47348,N_43750,N_42103);
xnor U47349 (N_47349,N_41715,N_42255);
nor U47350 (N_47350,N_40302,N_44071);
nor U47351 (N_47351,N_41557,N_43226);
nor U47352 (N_47352,N_43579,N_43022);
nand U47353 (N_47353,N_43941,N_43862);
or U47354 (N_47354,N_42073,N_40361);
nand U47355 (N_47355,N_44895,N_43796);
and U47356 (N_47356,N_43592,N_41477);
nand U47357 (N_47357,N_42993,N_42340);
nand U47358 (N_47358,N_42595,N_44808);
nor U47359 (N_47359,N_41391,N_43209);
nor U47360 (N_47360,N_40257,N_40606);
nand U47361 (N_47361,N_43369,N_40398);
nand U47362 (N_47362,N_40043,N_43270);
xnor U47363 (N_47363,N_42496,N_41025);
or U47364 (N_47364,N_41084,N_42987);
nor U47365 (N_47365,N_44546,N_42283);
and U47366 (N_47366,N_44692,N_44335);
or U47367 (N_47367,N_41326,N_41396);
nor U47368 (N_47368,N_44336,N_41322);
nand U47369 (N_47369,N_43160,N_40098);
or U47370 (N_47370,N_40324,N_43745);
nand U47371 (N_47371,N_41818,N_42959);
or U47372 (N_47372,N_41531,N_41376);
nor U47373 (N_47373,N_44270,N_40035);
and U47374 (N_47374,N_44457,N_42437);
xnor U47375 (N_47375,N_42173,N_42346);
nand U47376 (N_47376,N_40558,N_42144);
nor U47377 (N_47377,N_41524,N_44063);
and U47378 (N_47378,N_41772,N_42918);
or U47379 (N_47379,N_40543,N_42797);
nor U47380 (N_47380,N_43768,N_42770);
or U47381 (N_47381,N_40314,N_41816);
or U47382 (N_47382,N_41832,N_42271);
or U47383 (N_47383,N_44773,N_42325);
and U47384 (N_47384,N_42428,N_42783);
or U47385 (N_47385,N_41530,N_43315);
and U47386 (N_47386,N_41595,N_44018);
xnor U47387 (N_47387,N_42933,N_44160);
xnor U47388 (N_47388,N_42913,N_43641);
and U47389 (N_47389,N_44227,N_42801);
and U47390 (N_47390,N_40751,N_44394);
nor U47391 (N_47391,N_43623,N_43571);
nand U47392 (N_47392,N_41643,N_41703);
nor U47393 (N_47393,N_44928,N_43722);
nand U47394 (N_47394,N_42320,N_44274);
or U47395 (N_47395,N_43424,N_41416);
and U47396 (N_47396,N_43452,N_40522);
nor U47397 (N_47397,N_43549,N_44368);
nand U47398 (N_47398,N_42745,N_44850);
or U47399 (N_47399,N_41306,N_43311);
xor U47400 (N_47400,N_40020,N_42491);
xor U47401 (N_47401,N_40930,N_43982);
and U47402 (N_47402,N_42614,N_43890);
xor U47403 (N_47403,N_40820,N_41340);
or U47404 (N_47404,N_44821,N_42548);
and U47405 (N_47405,N_41926,N_44889);
nand U47406 (N_47406,N_43830,N_41437);
or U47407 (N_47407,N_44401,N_44729);
or U47408 (N_47408,N_42460,N_42994);
nand U47409 (N_47409,N_41589,N_43245);
nand U47410 (N_47410,N_40363,N_43953);
nand U47411 (N_47411,N_40408,N_41874);
and U47412 (N_47412,N_44282,N_43649);
xnor U47413 (N_47413,N_40046,N_41355);
nor U47414 (N_47414,N_42138,N_43408);
xor U47415 (N_47415,N_44413,N_43888);
nor U47416 (N_47416,N_40768,N_43710);
nand U47417 (N_47417,N_40927,N_43669);
nand U47418 (N_47418,N_41167,N_41067);
nand U47419 (N_47419,N_43261,N_44727);
nand U47420 (N_47420,N_41825,N_41802);
or U47421 (N_47421,N_42268,N_40480);
nor U47422 (N_47422,N_44079,N_40945);
and U47423 (N_47423,N_42390,N_44545);
xor U47424 (N_47424,N_43179,N_42284);
and U47425 (N_47425,N_40251,N_40440);
and U47426 (N_47426,N_40716,N_41760);
nor U47427 (N_47427,N_43825,N_41718);
nor U47428 (N_47428,N_40054,N_40839);
xnor U47429 (N_47429,N_42418,N_42702);
xnor U47430 (N_47430,N_41447,N_42568);
nor U47431 (N_47431,N_43793,N_44031);
xnor U47432 (N_47432,N_40003,N_44604);
nor U47433 (N_47433,N_42810,N_40743);
and U47434 (N_47434,N_40024,N_42038);
nor U47435 (N_47435,N_43943,N_42734);
nand U47436 (N_47436,N_41985,N_42669);
and U47437 (N_47437,N_44181,N_42470);
nand U47438 (N_47438,N_41763,N_40159);
xor U47439 (N_47439,N_44537,N_42885);
and U47440 (N_47440,N_41374,N_40092);
and U47441 (N_47441,N_42904,N_44404);
nand U47442 (N_47442,N_42857,N_43348);
xnor U47443 (N_47443,N_41445,N_40214);
or U47444 (N_47444,N_40759,N_43062);
or U47445 (N_47445,N_43766,N_40056);
or U47446 (N_47446,N_42385,N_41276);
nand U47447 (N_47447,N_41310,N_42573);
nor U47448 (N_47448,N_40355,N_42059);
and U47449 (N_47449,N_44431,N_44059);
nor U47450 (N_47450,N_44100,N_44222);
xor U47451 (N_47451,N_42619,N_43473);
or U47452 (N_47452,N_42085,N_42217);
xor U47453 (N_47453,N_43923,N_41979);
nor U47454 (N_47454,N_44820,N_43117);
nand U47455 (N_47455,N_42165,N_42871);
nor U47456 (N_47456,N_40080,N_44630);
nand U47457 (N_47457,N_42178,N_41129);
nand U47458 (N_47458,N_40581,N_43930);
or U47459 (N_47459,N_44641,N_40750);
nor U47460 (N_47460,N_41233,N_44255);
and U47461 (N_47461,N_43290,N_40554);
or U47462 (N_47462,N_40437,N_40955);
nor U47463 (N_47463,N_40237,N_44623);
and U47464 (N_47464,N_43175,N_42837);
nor U47465 (N_47465,N_43470,N_40574);
nor U47466 (N_47466,N_42906,N_40299);
nand U47467 (N_47467,N_40210,N_40721);
xor U47468 (N_47468,N_44632,N_43697);
xor U47469 (N_47469,N_42171,N_43996);
nand U47470 (N_47470,N_41639,N_43694);
nand U47471 (N_47471,N_40353,N_41627);
nand U47472 (N_47472,N_43068,N_40781);
or U47473 (N_47473,N_41970,N_42058);
or U47474 (N_47474,N_43991,N_40286);
and U47475 (N_47475,N_40218,N_40847);
nand U47476 (N_47476,N_42163,N_40034);
nor U47477 (N_47477,N_42310,N_42967);
xor U47478 (N_47478,N_41678,N_41952);
nand U47479 (N_47479,N_41658,N_40885);
xnor U47480 (N_47480,N_42032,N_40611);
and U47481 (N_47481,N_43384,N_43074);
and U47482 (N_47482,N_43726,N_42844);
nand U47483 (N_47483,N_40225,N_44798);
or U47484 (N_47484,N_42441,N_42872);
xor U47485 (N_47485,N_42892,N_41691);
nor U47486 (N_47486,N_41495,N_44352);
or U47487 (N_47487,N_43107,N_41075);
or U47488 (N_47488,N_41106,N_40191);
xor U47489 (N_47489,N_43524,N_42572);
nand U47490 (N_47490,N_43339,N_41875);
and U47491 (N_47491,N_42405,N_44935);
or U47492 (N_47492,N_43624,N_43045);
xor U47493 (N_47493,N_44153,N_40364);
or U47494 (N_47494,N_43640,N_40029);
xor U47495 (N_47495,N_40427,N_42015);
xor U47496 (N_47496,N_42387,N_40609);
and U47497 (N_47497,N_44963,N_42561);
xnor U47498 (N_47498,N_40613,N_43605);
or U47499 (N_47499,N_42056,N_40529);
nor U47500 (N_47500,N_41545,N_42822);
nand U47501 (N_47501,N_42556,N_44290);
xnor U47502 (N_47502,N_41541,N_41881);
xnor U47503 (N_47503,N_43620,N_42248);
and U47504 (N_47504,N_40819,N_44271);
and U47505 (N_47505,N_40191,N_42529);
or U47506 (N_47506,N_42899,N_44504);
nand U47507 (N_47507,N_40949,N_40146);
nor U47508 (N_47508,N_43802,N_41850);
nor U47509 (N_47509,N_42198,N_41464);
or U47510 (N_47510,N_43886,N_40873);
and U47511 (N_47511,N_42983,N_43960);
nor U47512 (N_47512,N_42425,N_42978);
nand U47513 (N_47513,N_42646,N_44858);
xor U47514 (N_47514,N_40725,N_42837);
nor U47515 (N_47515,N_41541,N_41809);
xnor U47516 (N_47516,N_41209,N_42343);
nand U47517 (N_47517,N_40819,N_42325);
nor U47518 (N_47518,N_44815,N_43311);
nor U47519 (N_47519,N_42446,N_40343);
nor U47520 (N_47520,N_40354,N_40501);
nor U47521 (N_47521,N_43256,N_44802);
nor U47522 (N_47522,N_43219,N_43765);
nor U47523 (N_47523,N_40295,N_40345);
xnor U47524 (N_47524,N_43061,N_40473);
nor U47525 (N_47525,N_43300,N_42841);
nor U47526 (N_47526,N_42688,N_43864);
nand U47527 (N_47527,N_40706,N_42732);
and U47528 (N_47528,N_42985,N_40895);
and U47529 (N_47529,N_41899,N_41875);
nor U47530 (N_47530,N_41710,N_44528);
nand U47531 (N_47531,N_44912,N_42380);
nor U47532 (N_47532,N_43654,N_42846);
nand U47533 (N_47533,N_44635,N_40275);
nand U47534 (N_47534,N_42316,N_44190);
or U47535 (N_47535,N_44627,N_44275);
nor U47536 (N_47536,N_41500,N_40139);
xnor U47537 (N_47537,N_41650,N_42256);
xor U47538 (N_47538,N_42999,N_43652);
xnor U47539 (N_47539,N_41906,N_41976);
or U47540 (N_47540,N_40507,N_42357);
and U47541 (N_47541,N_40335,N_40856);
and U47542 (N_47542,N_44121,N_41170);
nand U47543 (N_47543,N_41372,N_42161);
nor U47544 (N_47544,N_42511,N_42973);
and U47545 (N_47545,N_44936,N_44006);
nor U47546 (N_47546,N_44497,N_44526);
or U47547 (N_47547,N_41840,N_40245);
xor U47548 (N_47548,N_41605,N_43751);
nand U47549 (N_47549,N_42339,N_43015);
xnor U47550 (N_47550,N_41482,N_42627);
or U47551 (N_47551,N_44400,N_40325);
nand U47552 (N_47552,N_43563,N_40496);
and U47553 (N_47553,N_43312,N_41164);
nor U47554 (N_47554,N_40905,N_42050);
or U47555 (N_47555,N_41667,N_42256);
nor U47556 (N_47556,N_40962,N_43652);
nor U47557 (N_47557,N_42701,N_44379);
nand U47558 (N_47558,N_40357,N_44677);
and U47559 (N_47559,N_44319,N_42175);
and U47560 (N_47560,N_44350,N_43409);
nor U47561 (N_47561,N_41033,N_43209);
nor U47562 (N_47562,N_42557,N_43825);
or U47563 (N_47563,N_44728,N_41021);
or U47564 (N_47564,N_40094,N_41124);
xor U47565 (N_47565,N_42809,N_40701);
nor U47566 (N_47566,N_44306,N_40070);
or U47567 (N_47567,N_40685,N_41750);
or U47568 (N_47568,N_44575,N_40101);
nand U47569 (N_47569,N_44273,N_44826);
and U47570 (N_47570,N_44255,N_40382);
xor U47571 (N_47571,N_44264,N_41765);
xor U47572 (N_47572,N_41458,N_40514);
nor U47573 (N_47573,N_40808,N_41426);
xor U47574 (N_47574,N_44048,N_43470);
and U47575 (N_47575,N_40958,N_43347);
xnor U47576 (N_47576,N_40186,N_43262);
and U47577 (N_47577,N_44357,N_40663);
nand U47578 (N_47578,N_42768,N_43173);
xor U47579 (N_47579,N_41182,N_42432);
and U47580 (N_47580,N_40834,N_44146);
nor U47581 (N_47581,N_41837,N_41269);
or U47582 (N_47582,N_43107,N_42585);
nor U47583 (N_47583,N_43324,N_42171);
or U47584 (N_47584,N_41010,N_44556);
xor U47585 (N_47585,N_41494,N_43691);
nand U47586 (N_47586,N_42781,N_44886);
nand U47587 (N_47587,N_40489,N_44649);
nor U47588 (N_47588,N_40041,N_41282);
or U47589 (N_47589,N_40950,N_42282);
nor U47590 (N_47590,N_41038,N_41192);
nor U47591 (N_47591,N_43756,N_40888);
or U47592 (N_47592,N_41656,N_42581);
xnor U47593 (N_47593,N_40317,N_42148);
or U47594 (N_47594,N_42306,N_41772);
nor U47595 (N_47595,N_42952,N_40180);
nor U47596 (N_47596,N_40397,N_41411);
or U47597 (N_47597,N_43858,N_42855);
or U47598 (N_47598,N_44797,N_41456);
nor U47599 (N_47599,N_40156,N_41856);
xor U47600 (N_47600,N_42778,N_40666);
nand U47601 (N_47601,N_41002,N_43131);
xor U47602 (N_47602,N_44431,N_43659);
or U47603 (N_47603,N_41617,N_41793);
and U47604 (N_47604,N_41747,N_43459);
and U47605 (N_47605,N_44197,N_42078);
nor U47606 (N_47606,N_40415,N_41190);
xnor U47607 (N_47607,N_40066,N_40049);
and U47608 (N_47608,N_41563,N_43330);
xnor U47609 (N_47609,N_41144,N_43589);
and U47610 (N_47610,N_40040,N_40440);
and U47611 (N_47611,N_44954,N_43803);
and U47612 (N_47612,N_42586,N_41155);
or U47613 (N_47613,N_41918,N_40033);
nor U47614 (N_47614,N_43946,N_43603);
or U47615 (N_47615,N_40976,N_44372);
or U47616 (N_47616,N_43411,N_40882);
or U47617 (N_47617,N_40373,N_43510);
nand U47618 (N_47618,N_42309,N_40613);
nand U47619 (N_47619,N_41629,N_41726);
and U47620 (N_47620,N_43736,N_41658);
nor U47621 (N_47621,N_43641,N_44694);
and U47622 (N_47622,N_40151,N_44563);
and U47623 (N_47623,N_44194,N_42802);
nand U47624 (N_47624,N_41977,N_41159);
nand U47625 (N_47625,N_44696,N_43040);
and U47626 (N_47626,N_41006,N_40296);
xor U47627 (N_47627,N_44494,N_44539);
and U47628 (N_47628,N_41513,N_42388);
nand U47629 (N_47629,N_41811,N_44774);
xnor U47630 (N_47630,N_40614,N_40836);
or U47631 (N_47631,N_42796,N_43260);
nand U47632 (N_47632,N_40143,N_44315);
nand U47633 (N_47633,N_41635,N_44568);
nand U47634 (N_47634,N_41224,N_40088);
or U47635 (N_47635,N_43060,N_44960);
and U47636 (N_47636,N_41160,N_41061);
nor U47637 (N_47637,N_40399,N_41510);
nand U47638 (N_47638,N_40965,N_40276);
nor U47639 (N_47639,N_42104,N_40327);
nor U47640 (N_47640,N_40409,N_43698);
nor U47641 (N_47641,N_40002,N_44450);
nor U47642 (N_47642,N_43129,N_42971);
or U47643 (N_47643,N_42218,N_43239);
xor U47644 (N_47644,N_43650,N_41537);
and U47645 (N_47645,N_40909,N_42874);
and U47646 (N_47646,N_42087,N_40826);
nand U47647 (N_47647,N_43052,N_40084);
nor U47648 (N_47648,N_40481,N_40603);
nand U47649 (N_47649,N_44892,N_40578);
and U47650 (N_47650,N_42583,N_41959);
nand U47651 (N_47651,N_42620,N_41268);
xor U47652 (N_47652,N_44207,N_40301);
or U47653 (N_47653,N_40163,N_43848);
xnor U47654 (N_47654,N_41937,N_44859);
nand U47655 (N_47655,N_40511,N_42794);
and U47656 (N_47656,N_41462,N_41217);
and U47657 (N_47657,N_44975,N_42932);
nand U47658 (N_47658,N_44844,N_41867);
nor U47659 (N_47659,N_44578,N_40679);
and U47660 (N_47660,N_42483,N_42702);
xnor U47661 (N_47661,N_44374,N_43221);
xor U47662 (N_47662,N_44542,N_41990);
xnor U47663 (N_47663,N_41972,N_41678);
nand U47664 (N_47664,N_44022,N_42453);
xor U47665 (N_47665,N_44439,N_44851);
nor U47666 (N_47666,N_43176,N_44089);
and U47667 (N_47667,N_42378,N_40760);
xor U47668 (N_47668,N_40828,N_41906);
xnor U47669 (N_47669,N_44450,N_40516);
and U47670 (N_47670,N_41509,N_42055);
and U47671 (N_47671,N_41352,N_40374);
nand U47672 (N_47672,N_41131,N_44527);
nand U47673 (N_47673,N_44194,N_42426);
xnor U47674 (N_47674,N_44043,N_42268);
xor U47675 (N_47675,N_43597,N_40693);
nor U47676 (N_47676,N_42914,N_41364);
xnor U47677 (N_47677,N_40113,N_42445);
nand U47678 (N_47678,N_42840,N_43274);
or U47679 (N_47679,N_40017,N_41969);
and U47680 (N_47680,N_40963,N_40562);
xor U47681 (N_47681,N_40041,N_41252);
nand U47682 (N_47682,N_40819,N_43683);
nand U47683 (N_47683,N_42558,N_40876);
xnor U47684 (N_47684,N_41509,N_44786);
nor U47685 (N_47685,N_44602,N_43316);
xor U47686 (N_47686,N_44610,N_40503);
and U47687 (N_47687,N_43749,N_44322);
xnor U47688 (N_47688,N_43351,N_44894);
nand U47689 (N_47689,N_40955,N_43069);
nand U47690 (N_47690,N_41379,N_41933);
nor U47691 (N_47691,N_44247,N_41458);
nor U47692 (N_47692,N_40591,N_42939);
or U47693 (N_47693,N_42844,N_44579);
and U47694 (N_47694,N_40094,N_42263);
or U47695 (N_47695,N_44479,N_42832);
nand U47696 (N_47696,N_42517,N_40534);
nor U47697 (N_47697,N_44541,N_43812);
nor U47698 (N_47698,N_43681,N_41403);
nand U47699 (N_47699,N_44222,N_41556);
nand U47700 (N_47700,N_40582,N_40503);
nand U47701 (N_47701,N_43035,N_44857);
and U47702 (N_47702,N_43030,N_44452);
or U47703 (N_47703,N_44862,N_40286);
or U47704 (N_47704,N_40580,N_40051);
nand U47705 (N_47705,N_41017,N_44410);
nand U47706 (N_47706,N_41530,N_40952);
nand U47707 (N_47707,N_44261,N_44465);
nor U47708 (N_47708,N_41505,N_44704);
and U47709 (N_47709,N_43311,N_42224);
and U47710 (N_47710,N_41267,N_41673);
nand U47711 (N_47711,N_44041,N_40896);
xnor U47712 (N_47712,N_40207,N_41415);
nand U47713 (N_47713,N_41140,N_42685);
or U47714 (N_47714,N_44721,N_42846);
xnor U47715 (N_47715,N_44720,N_43206);
or U47716 (N_47716,N_41622,N_41156);
nand U47717 (N_47717,N_41561,N_41119);
nor U47718 (N_47718,N_41378,N_41438);
nand U47719 (N_47719,N_40800,N_42027);
and U47720 (N_47720,N_44470,N_44606);
xor U47721 (N_47721,N_40701,N_43480);
nor U47722 (N_47722,N_41961,N_44425);
nor U47723 (N_47723,N_44585,N_43394);
and U47724 (N_47724,N_42068,N_42986);
and U47725 (N_47725,N_42214,N_41340);
xor U47726 (N_47726,N_40512,N_40211);
or U47727 (N_47727,N_44439,N_41846);
nand U47728 (N_47728,N_44195,N_42574);
xnor U47729 (N_47729,N_43548,N_42915);
nand U47730 (N_47730,N_40175,N_41014);
nor U47731 (N_47731,N_43275,N_43020);
nor U47732 (N_47732,N_41302,N_43164);
nand U47733 (N_47733,N_40385,N_43055);
nand U47734 (N_47734,N_42973,N_42175);
xor U47735 (N_47735,N_42178,N_40479);
or U47736 (N_47736,N_43540,N_44804);
and U47737 (N_47737,N_43710,N_43184);
nor U47738 (N_47738,N_43124,N_41330);
xor U47739 (N_47739,N_41546,N_41675);
nor U47740 (N_47740,N_41796,N_44862);
and U47741 (N_47741,N_41135,N_44291);
and U47742 (N_47742,N_41296,N_43268);
nand U47743 (N_47743,N_43604,N_41485);
xor U47744 (N_47744,N_44632,N_44599);
and U47745 (N_47745,N_44168,N_43748);
nor U47746 (N_47746,N_41054,N_44808);
and U47747 (N_47747,N_43605,N_42602);
nor U47748 (N_47748,N_40675,N_42199);
and U47749 (N_47749,N_44886,N_43094);
xor U47750 (N_47750,N_42204,N_43780);
nor U47751 (N_47751,N_40205,N_41814);
xnor U47752 (N_47752,N_44520,N_40525);
nor U47753 (N_47753,N_40539,N_42550);
nor U47754 (N_47754,N_41221,N_40177);
nor U47755 (N_47755,N_44468,N_44651);
or U47756 (N_47756,N_41606,N_40034);
or U47757 (N_47757,N_41977,N_43360);
and U47758 (N_47758,N_44578,N_43156);
or U47759 (N_47759,N_41019,N_43582);
nor U47760 (N_47760,N_42444,N_44601);
nor U47761 (N_47761,N_41435,N_41533);
and U47762 (N_47762,N_41060,N_43142);
and U47763 (N_47763,N_40004,N_43298);
or U47764 (N_47764,N_41871,N_41622);
xnor U47765 (N_47765,N_42631,N_40513);
or U47766 (N_47766,N_44441,N_43731);
or U47767 (N_47767,N_44801,N_43836);
or U47768 (N_47768,N_42775,N_43118);
nor U47769 (N_47769,N_43913,N_41292);
and U47770 (N_47770,N_40695,N_42004);
nand U47771 (N_47771,N_41718,N_44521);
nor U47772 (N_47772,N_43101,N_43670);
and U47773 (N_47773,N_40457,N_42606);
or U47774 (N_47774,N_44924,N_41884);
nand U47775 (N_47775,N_43555,N_42553);
xnor U47776 (N_47776,N_44462,N_44722);
and U47777 (N_47777,N_44771,N_44841);
xnor U47778 (N_47778,N_41170,N_41754);
or U47779 (N_47779,N_40675,N_44534);
xor U47780 (N_47780,N_43538,N_43784);
nor U47781 (N_47781,N_43800,N_40206);
nor U47782 (N_47782,N_44833,N_41952);
or U47783 (N_47783,N_43247,N_40046);
and U47784 (N_47784,N_42644,N_44144);
nand U47785 (N_47785,N_43259,N_42239);
nor U47786 (N_47786,N_42896,N_43152);
and U47787 (N_47787,N_41077,N_42164);
or U47788 (N_47788,N_43430,N_44726);
nand U47789 (N_47789,N_40807,N_40818);
nor U47790 (N_47790,N_44257,N_40247);
and U47791 (N_47791,N_43069,N_41193);
and U47792 (N_47792,N_44772,N_44500);
nand U47793 (N_47793,N_40542,N_40469);
nor U47794 (N_47794,N_40854,N_41314);
and U47795 (N_47795,N_42469,N_42319);
or U47796 (N_47796,N_43214,N_43096);
nand U47797 (N_47797,N_44595,N_40715);
and U47798 (N_47798,N_40649,N_42823);
nand U47799 (N_47799,N_41114,N_43026);
nand U47800 (N_47800,N_41280,N_42848);
and U47801 (N_47801,N_43266,N_43825);
nor U47802 (N_47802,N_44317,N_43527);
or U47803 (N_47803,N_40300,N_42228);
and U47804 (N_47804,N_43577,N_41437);
nand U47805 (N_47805,N_43224,N_40948);
nand U47806 (N_47806,N_44490,N_41886);
or U47807 (N_47807,N_41986,N_43000);
and U47808 (N_47808,N_40621,N_41064);
nand U47809 (N_47809,N_40204,N_42055);
nor U47810 (N_47810,N_44510,N_41885);
and U47811 (N_47811,N_43160,N_43467);
nor U47812 (N_47812,N_44477,N_41449);
and U47813 (N_47813,N_44771,N_42072);
and U47814 (N_47814,N_42827,N_43978);
nor U47815 (N_47815,N_42228,N_41651);
nand U47816 (N_47816,N_42725,N_41865);
xnor U47817 (N_47817,N_40743,N_41045);
nand U47818 (N_47818,N_44818,N_44684);
nor U47819 (N_47819,N_43959,N_43007);
or U47820 (N_47820,N_44278,N_40105);
nand U47821 (N_47821,N_43436,N_43353);
and U47822 (N_47822,N_40365,N_44048);
nand U47823 (N_47823,N_40624,N_40741);
or U47824 (N_47824,N_41995,N_43259);
xor U47825 (N_47825,N_43577,N_42294);
and U47826 (N_47826,N_41906,N_40920);
and U47827 (N_47827,N_44534,N_40589);
or U47828 (N_47828,N_43985,N_44954);
and U47829 (N_47829,N_44520,N_44488);
and U47830 (N_47830,N_42267,N_42495);
nor U47831 (N_47831,N_42133,N_41571);
nor U47832 (N_47832,N_43468,N_41553);
xnor U47833 (N_47833,N_40296,N_43576);
nand U47834 (N_47834,N_43142,N_44756);
or U47835 (N_47835,N_43066,N_40545);
nand U47836 (N_47836,N_40798,N_44092);
nor U47837 (N_47837,N_41884,N_40963);
xor U47838 (N_47838,N_44304,N_40738);
xnor U47839 (N_47839,N_44916,N_43329);
nand U47840 (N_47840,N_43720,N_42526);
nand U47841 (N_47841,N_43739,N_40765);
or U47842 (N_47842,N_43604,N_42636);
or U47843 (N_47843,N_42205,N_44147);
xnor U47844 (N_47844,N_44394,N_40024);
nor U47845 (N_47845,N_42742,N_40582);
nor U47846 (N_47846,N_44359,N_44695);
nand U47847 (N_47847,N_41438,N_41737);
or U47848 (N_47848,N_44021,N_40550);
and U47849 (N_47849,N_41855,N_41471);
and U47850 (N_47850,N_40753,N_44958);
nor U47851 (N_47851,N_42814,N_41408);
nand U47852 (N_47852,N_40816,N_40679);
xnor U47853 (N_47853,N_43803,N_41487);
nor U47854 (N_47854,N_42424,N_40364);
nand U47855 (N_47855,N_40150,N_40295);
nor U47856 (N_47856,N_43367,N_41013);
or U47857 (N_47857,N_41343,N_41951);
nand U47858 (N_47858,N_41240,N_43440);
or U47859 (N_47859,N_43103,N_44718);
nand U47860 (N_47860,N_40915,N_41952);
xnor U47861 (N_47861,N_42991,N_42445);
or U47862 (N_47862,N_44683,N_42278);
nand U47863 (N_47863,N_42043,N_44667);
nand U47864 (N_47864,N_44943,N_44589);
and U47865 (N_47865,N_40501,N_42894);
xnor U47866 (N_47866,N_41675,N_43097);
nand U47867 (N_47867,N_41879,N_43640);
and U47868 (N_47868,N_42914,N_40725);
or U47869 (N_47869,N_44708,N_43012);
and U47870 (N_47870,N_41772,N_44287);
nor U47871 (N_47871,N_40670,N_42528);
nor U47872 (N_47872,N_43606,N_44338);
and U47873 (N_47873,N_44273,N_41233);
nand U47874 (N_47874,N_43802,N_42412);
nand U47875 (N_47875,N_44891,N_41345);
nor U47876 (N_47876,N_42897,N_41534);
nand U47877 (N_47877,N_43707,N_43427);
or U47878 (N_47878,N_43163,N_42184);
nand U47879 (N_47879,N_44413,N_44816);
or U47880 (N_47880,N_43006,N_43308);
nand U47881 (N_47881,N_41540,N_41946);
or U47882 (N_47882,N_44381,N_40754);
or U47883 (N_47883,N_43474,N_42153);
nand U47884 (N_47884,N_40489,N_44547);
nor U47885 (N_47885,N_43048,N_43878);
xnor U47886 (N_47886,N_44357,N_40161);
xor U47887 (N_47887,N_43156,N_40464);
xnor U47888 (N_47888,N_40880,N_41779);
nor U47889 (N_47889,N_41009,N_44152);
nor U47890 (N_47890,N_40746,N_40177);
and U47891 (N_47891,N_44652,N_41395);
xor U47892 (N_47892,N_40952,N_41236);
nand U47893 (N_47893,N_42404,N_42193);
xnor U47894 (N_47894,N_41438,N_41946);
nor U47895 (N_47895,N_42749,N_42888);
xor U47896 (N_47896,N_42290,N_41523);
xor U47897 (N_47897,N_43087,N_42911);
or U47898 (N_47898,N_40888,N_44099);
and U47899 (N_47899,N_40346,N_41134);
nor U47900 (N_47900,N_40235,N_40660);
nor U47901 (N_47901,N_42859,N_42410);
and U47902 (N_47902,N_44061,N_40602);
xnor U47903 (N_47903,N_44810,N_42382);
nor U47904 (N_47904,N_42534,N_40909);
nand U47905 (N_47905,N_41806,N_40241);
nand U47906 (N_47906,N_43992,N_42803);
nand U47907 (N_47907,N_43253,N_41237);
nand U47908 (N_47908,N_44309,N_44968);
nand U47909 (N_47909,N_42942,N_40285);
xor U47910 (N_47910,N_44846,N_43045);
nor U47911 (N_47911,N_40776,N_42323);
or U47912 (N_47912,N_43295,N_42311);
nand U47913 (N_47913,N_40727,N_42264);
xor U47914 (N_47914,N_43779,N_42013);
nor U47915 (N_47915,N_42578,N_44354);
xnor U47916 (N_47916,N_40364,N_43100);
or U47917 (N_47917,N_40585,N_43092);
or U47918 (N_47918,N_43919,N_43120);
and U47919 (N_47919,N_42161,N_40093);
and U47920 (N_47920,N_40749,N_43956);
or U47921 (N_47921,N_43801,N_41938);
xnor U47922 (N_47922,N_42699,N_42269);
nor U47923 (N_47923,N_40675,N_42194);
xnor U47924 (N_47924,N_43694,N_42907);
nand U47925 (N_47925,N_42115,N_44922);
and U47926 (N_47926,N_44195,N_40738);
nand U47927 (N_47927,N_43101,N_43931);
xor U47928 (N_47928,N_44398,N_42521);
or U47929 (N_47929,N_42487,N_44099);
or U47930 (N_47930,N_41072,N_44454);
and U47931 (N_47931,N_41072,N_43926);
and U47932 (N_47932,N_44132,N_40324);
and U47933 (N_47933,N_44786,N_43821);
xnor U47934 (N_47934,N_44974,N_44896);
nand U47935 (N_47935,N_40123,N_41778);
and U47936 (N_47936,N_43457,N_44208);
or U47937 (N_47937,N_41467,N_43231);
and U47938 (N_47938,N_40490,N_40901);
and U47939 (N_47939,N_42234,N_40085);
or U47940 (N_47940,N_44313,N_43676);
or U47941 (N_47941,N_44541,N_42021);
or U47942 (N_47942,N_44405,N_42786);
xnor U47943 (N_47943,N_44498,N_42715);
and U47944 (N_47944,N_41157,N_43599);
nor U47945 (N_47945,N_44582,N_41638);
xnor U47946 (N_47946,N_44651,N_41007);
and U47947 (N_47947,N_44815,N_42803);
nor U47948 (N_47948,N_42734,N_44833);
xor U47949 (N_47949,N_41483,N_44377);
nor U47950 (N_47950,N_43314,N_43329);
or U47951 (N_47951,N_41824,N_40319);
or U47952 (N_47952,N_44473,N_44289);
nand U47953 (N_47953,N_44784,N_41290);
nor U47954 (N_47954,N_43141,N_43994);
nand U47955 (N_47955,N_42098,N_42401);
xor U47956 (N_47956,N_41285,N_41501);
nand U47957 (N_47957,N_44594,N_43306);
nor U47958 (N_47958,N_41370,N_42863);
or U47959 (N_47959,N_42085,N_43050);
xor U47960 (N_47960,N_42888,N_40967);
xor U47961 (N_47961,N_43760,N_42181);
and U47962 (N_47962,N_44318,N_41512);
nor U47963 (N_47963,N_40567,N_41714);
nand U47964 (N_47964,N_43586,N_43095);
and U47965 (N_47965,N_44240,N_43837);
and U47966 (N_47966,N_40545,N_43985);
nor U47967 (N_47967,N_44764,N_44415);
or U47968 (N_47968,N_42783,N_44037);
nor U47969 (N_47969,N_43980,N_43244);
nor U47970 (N_47970,N_43080,N_42323);
or U47971 (N_47971,N_42180,N_42995);
xnor U47972 (N_47972,N_40080,N_41066);
or U47973 (N_47973,N_42529,N_44316);
or U47974 (N_47974,N_44472,N_43676);
and U47975 (N_47975,N_43677,N_44255);
and U47976 (N_47976,N_43222,N_41534);
and U47977 (N_47977,N_43686,N_40177);
nor U47978 (N_47978,N_43830,N_42344);
and U47979 (N_47979,N_42298,N_40755);
or U47980 (N_47980,N_42897,N_43076);
xor U47981 (N_47981,N_41621,N_42432);
or U47982 (N_47982,N_44914,N_40057);
xor U47983 (N_47983,N_42364,N_41818);
nor U47984 (N_47984,N_44649,N_41916);
nand U47985 (N_47985,N_42077,N_40603);
nand U47986 (N_47986,N_41722,N_42530);
nand U47987 (N_47987,N_42972,N_40619);
and U47988 (N_47988,N_43216,N_44547);
nor U47989 (N_47989,N_40578,N_40438);
nand U47990 (N_47990,N_40354,N_40782);
nor U47991 (N_47991,N_41626,N_42966);
and U47992 (N_47992,N_41714,N_40436);
xor U47993 (N_47993,N_40072,N_43215);
or U47994 (N_47994,N_43309,N_44135);
nand U47995 (N_47995,N_40893,N_42619);
or U47996 (N_47996,N_41041,N_44629);
or U47997 (N_47997,N_41507,N_40877);
and U47998 (N_47998,N_41690,N_43856);
nor U47999 (N_47999,N_43735,N_44025);
or U48000 (N_48000,N_40068,N_41061);
or U48001 (N_48001,N_40521,N_40088);
nand U48002 (N_48002,N_40460,N_42316);
nand U48003 (N_48003,N_44280,N_44868);
or U48004 (N_48004,N_42179,N_42954);
and U48005 (N_48005,N_44332,N_40282);
nor U48006 (N_48006,N_43532,N_40782);
and U48007 (N_48007,N_42795,N_40249);
or U48008 (N_48008,N_43509,N_40110);
and U48009 (N_48009,N_42792,N_40285);
xor U48010 (N_48010,N_40546,N_42087);
xor U48011 (N_48011,N_42459,N_41689);
or U48012 (N_48012,N_40662,N_41431);
nand U48013 (N_48013,N_40333,N_43991);
nand U48014 (N_48014,N_40359,N_43175);
nand U48015 (N_48015,N_43488,N_43718);
and U48016 (N_48016,N_40546,N_44671);
nand U48017 (N_48017,N_44100,N_44822);
or U48018 (N_48018,N_42055,N_40033);
or U48019 (N_48019,N_44083,N_40180);
or U48020 (N_48020,N_40517,N_40208);
or U48021 (N_48021,N_43723,N_41667);
nand U48022 (N_48022,N_40183,N_41682);
or U48023 (N_48023,N_41994,N_41119);
or U48024 (N_48024,N_41256,N_43511);
and U48025 (N_48025,N_42700,N_41804);
nand U48026 (N_48026,N_40094,N_40863);
or U48027 (N_48027,N_40829,N_42815);
nor U48028 (N_48028,N_42972,N_42010);
nor U48029 (N_48029,N_41994,N_43220);
nand U48030 (N_48030,N_44438,N_40542);
and U48031 (N_48031,N_42608,N_43528);
xor U48032 (N_48032,N_40230,N_42089);
or U48033 (N_48033,N_43101,N_40018);
and U48034 (N_48034,N_40591,N_44491);
or U48035 (N_48035,N_42302,N_43226);
nand U48036 (N_48036,N_40842,N_42143);
nor U48037 (N_48037,N_43571,N_41235);
and U48038 (N_48038,N_41742,N_40736);
and U48039 (N_48039,N_42778,N_42652);
nand U48040 (N_48040,N_44380,N_43385);
or U48041 (N_48041,N_42155,N_44084);
nand U48042 (N_48042,N_43437,N_44591);
and U48043 (N_48043,N_41968,N_42091);
or U48044 (N_48044,N_40225,N_42150);
and U48045 (N_48045,N_40305,N_41724);
nand U48046 (N_48046,N_40213,N_41381);
nor U48047 (N_48047,N_41181,N_40790);
and U48048 (N_48048,N_41468,N_42016);
or U48049 (N_48049,N_43759,N_42044);
or U48050 (N_48050,N_41509,N_40648);
xor U48051 (N_48051,N_41364,N_40222);
nor U48052 (N_48052,N_41127,N_43505);
xor U48053 (N_48053,N_41413,N_44052);
and U48054 (N_48054,N_40836,N_44454);
or U48055 (N_48055,N_42249,N_40014);
nand U48056 (N_48056,N_40303,N_42329);
xnor U48057 (N_48057,N_40362,N_42851);
and U48058 (N_48058,N_40492,N_43162);
nor U48059 (N_48059,N_40856,N_44516);
or U48060 (N_48060,N_40420,N_42914);
and U48061 (N_48061,N_42451,N_44371);
and U48062 (N_48062,N_40109,N_43298);
xnor U48063 (N_48063,N_43863,N_40018);
nor U48064 (N_48064,N_41454,N_43963);
and U48065 (N_48065,N_41870,N_43968);
nand U48066 (N_48066,N_43918,N_43366);
nand U48067 (N_48067,N_43992,N_41620);
nand U48068 (N_48068,N_41741,N_44770);
nand U48069 (N_48069,N_44921,N_41345);
xor U48070 (N_48070,N_42643,N_43528);
nand U48071 (N_48071,N_43229,N_40948);
and U48072 (N_48072,N_41461,N_42142);
xnor U48073 (N_48073,N_41115,N_43233);
or U48074 (N_48074,N_41543,N_42099);
or U48075 (N_48075,N_43216,N_42367);
xor U48076 (N_48076,N_40795,N_44092);
and U48077 (N_48077,N_40612,N_44953);
and U48078 (N_48078,N_44920,N_42946);
or U48079 (N_48079,N_42896,N_44646);
nand U48080 (N_48080,N_40882,N_43123);
nor U48081 (N_48081,N_40584,N_42992);
and U48082 (N_48082,N_41679,N_44609);
xor U48083 (N_48083,N_42221,N_43339);
or U48084 (N_48084,N_42765,N_43771);
or U48085 (N_48085,N_43548,N_43303);
nor U48086 (N_48086,N_40688,N_44318);
and U48087 (N_48087,N_41347,N_40530);
nor U48088 (N_48088,N_41679,N_41677);
and U48089 (N_48089,N_42254,N_40031);
or U48090 (N_48090,N_44825,N_42844);
and U48091 (N_48091,N_41529,N_42818);
and U48092 (N_48092,N_41770,N_40641);
and U48093 (N_48093,N_41972,N_41970);
xor U48094 (N_48094,N_41511,N_44300);
nand U48095 (N_48095,N_44198,N_40274);
nand U48096 (N_48096,N_41938,N_40540);
nand U48097 (N_48097,N_43893,N_40412);
nor U48098 (N_48098,N_40152,N_43785);
nand U48099 (N_48099,N_43799,N_43916);
and U48100 (N_48100,N_43979,N_41826);
or U48101 (N_48101,N_41412,N_44137);
or U48102 (N_48102,N_42418,N_41868);
xnor U48103 (N_48103,N_42777,N_43318);
xor U48104 (N_48104,N_42829,N_43910);
and U48105 (N_48105,N_42804,N_40145);
nor U48106 (N_48106,N_42875,N_44693);
xnor U48107 (N_48107,N_44789,N_42088);
or U48108 (N_48108,N_41568,N_41105);
xor U48109 (N_48109,N_41948,N_42330);
and U48110 (N_48110,N_44842,N_41807);
or U48111 (N_48111,N_41932,N_44979);
and U48112 (N_48112,N_41039,N_41417);
nor U48113 (N_48113,N_44406,N_41369);
xnor U48114 (N_48114,N_43332,N_44662);
nor U48115 (N_48115,N_43735,N_42193);
xnor U48116 (N_48116,N_41464,N_41280);
and U48117 (N_48117,N_42399,N_43350);
or U48118 (N_48118,N_41741,N_40639);
and U48119 (N_48119,N_41997,N_42377);
or U48120 (N_48120,N_41736,N_44550);
nor U48121 (N_48121,N_42256,N_40363);
or U48122 (N_48122,N_44585,N_40978);
nor U48123 (N_48123,N_42165,N_42228);
xnor U48124 (N_48124,N_43874,N_44627);
nand U48125 (N_48125,N_41901,N_40335);
xor U48126 (N_48126,N_42629,N_40312);
xnor U48127 (N_48127,N_43580,N_42169);
nand U48128 (N_48128,N_40094,N_44282);
and U48129 (N_48129,N_41758,N_44538);
nor U48130 (N_48130,N_42701,N_43079);
xor U48131 (N_48131,N_40125,N_40064);
nand U48132 (N_48132,N_42208,N_40543);
nand U48133 (N_48133,N_44436,N_42263);
nand U48134 (N_48134,N_42002,N_41681);
and U48135 (N_48135,N_44571,N_40800);
and U48136 (N_48136,N_41243,N_41859);
or U48137 (N_48137,N_43506,N_41030);
or U48138 (N_48138,N_40342,N_44146);
xnor U48139 (N_48139,N_42514,N_43461);
or U48140 (N_48140,N_44358,N_41724);
or U48141 (N_48141,N_44917,N_43908);
or U48142 (N_48142,N_43554,N_44228);
xnor U48143 (N_48143,N_40727,N_43583);
and U48144 (N_48144,N_40029,N_41547);
nand U48145 (N_48145,N_41647,N_43093);
nand U48146 (N_48146,N_44476,N_44963);
nor U48147 (N_48147,N_43352,N_41730);
or U48148 (N_48148,N_41458,N_41830);
nor U48149 (N_48149,N_42852,N_42828);
and U48150 (N_48150,N_44605,N_42970);
xnor U48151 (N_48151,N_42205,N_42008);
nand U48152 (N_48152,N_43881,N_43991);
or U48153 (N_48153,N_41953,N_41710);
nor U48154 (N_48154,N_44686,N_44847);
xor U48155 (N_48155,N_44294,N_42154);
xor U48156 (N_48156,N_41754,N_40372);
xnor U48157 (N_48157,N_43811,N_43395);
and U48158 (N_48158,N_42548,N_44382);
nor U48159 (N_48159,N_43321,N_40174);
or U48160 (N_48160,N_41176,N_40942);
or U48161 (N_48161,N_40659,N_42903);
nand U48162 (N_48162,N_44247,N_43148);
nand U48163 (N_48163,N_40609,N_40971);
and U48164 (N_48164,N_41667,N_44595);
nand U48165 (N_48165,N_43398,N_40023);
xnor U48166 (N_48166,N_40806,N_43620);
nor U48167 (N_48167,N_44766,N_40525);
nand U48168 (N_48168,N_41076,N_40867);
and U48169 (N_48169,N_40346,N_42022);
or U48170 (N_48170,N_42908,N_41855);
nor U48171 (N_48171,N_40060,N_43197);
or U48172 (N_48172,N_44089,N_42187);
and U48173 (N_48173,N_44848,N_43335);
and U48174 (N_48174,N_41922,N_41015);
xor U48175 (N_48175,N_40816,N_42975);
xor U48176 (N_48176,N_44349,N_41304);
nor U48177 (N_48177,N_42274,N_43597);
and U48178 (N_48178,N_41445,N_42917);
nor U48179 (N_48179,N_42718,N_43112);
nand U48180 (N_48180,N_43585,N_43627);
nor U48181 (N_48181,N_41935,N_40084);
nor U48182 (N_48182,N_44196,N_42987);
nor U48183 (N_48183,N_42996,N_41542);
and U48184 (N_48184,N_40916,N_44558);
nor U48185 (N_48185,N_42005,N_42418);
nor U48186 (N_48186,N_44659,N_44026);
xor U48187 (N_48187,N_41698,N_41240);
nor U48188 (N_48188,N_44620,N_42681);
and U48189 (N_48189,N_42003,N_42498);
or U48190 (N_48190,N_41964,N_40166);
xor U48191 (N_48191,N_40995,N_41862);
and U48192 (N_48192,N_44697,N_42597);
nor U48193 (N_48193,N_41687,N_42348);
or U48194 (N_48194,N_42657,N_43615);
or U48195 (N_48195,N_42686,N_41724);
xnor U48196 (N_48196,N_42145,N_42392);
xnor U48197 (N_48197,N_43143,N_43962);
or U48198 (N_48198,N_40571,N_42989);
and U48199 (N_48199,N_42542,N_40433);
nor U48200 (N_48200,N_41491,N_43067);
nand U48201 (N_48201,N_43580,N_44562);
xor U48202 (N_48202,N_41948,N_43658);
nor U48203 (N_48203,N_41387,N_41126);
and U48204 (N_48204,N_44818,N_42920);
and U48205 (N_48205,N_41668,N_44233);
or U48206 (N_48206,N_43162,N_44978);
or U48207 (N_48207,N_42113,N_43995);
or U48208 (N_48208,N_41741,N_40578);
and U48209 (N_48209,N_43151,N_41627);
xor U48210 (N_48210,N_41912,N_42606);
nand U48211 (N_48211,N_43229,N_40337);
xor U48212 (N_48212,N_42118,N_41486);
and U48213 (N_48213,N_41622,N_40645);
and U48214 (N_48214,N_43263,N_42113);
nor U48215 (N_48215,N_43521,N_43105);
or U48216 (N_48216,N_43201,N_43348);
nor U48217 (N_48217,N_41473,N_40443);
and U48218 (N_48218,N_42519,N_41765);
or U48219 (N_48219,N_43174,N_40092);
nand U48220 (N_48220,N_42545,N_41278);
xor U48221 (N_48221,N_44459,N_43322);
or U48222 (N_48222,N_43885,N_42645);
nand U48223 (N_48223,N_43391,N_42748);
xor U48224 (N_48224,N_42746,N_42634);
or U48225 (N_48225,N_43296,N_41622);
or U48226 (N_48226,N_44069,N_41099);
or U48227 (N_48227,N_44746,N_44887);
nand U48228 (N_48228,N_44377,N_43788);
or U48229 (N_48229,N_43712,N_42936);
nand U48230 (N_48230,N_43824,N_42299);
xnor U48231 (N_48231,N_43161,N_42477);
or U48232 (N_48232,N_42979,N_42457);
or U48233 (N_48233,N_44152,N_43158);
and U48234 (N_48234,N_43284,N_41641);
or U48235 (N_48235,N_40440,N_41413);
and U48236 (N_48236,N_43118,N_40262);
xnor U48237 (N_48237,N_41713,N_40169);
xor U48238 (N_48238,N_44468,N_43398);
or U48239 (N_48239,N_42358,N_42606);
or U48240 (N_48240,N_41624,N_44814);
nor U48241 (N_48241,N_41500,N_43019);
nand U48242 (N_48242,N_43796,N_42832);
nand U48243 (N_48243,N_44632,N_41019);
nand U48244 (N_48244,N_42363,N_43320);
or U48245 (N_48245,N_44472,N_43739);
and U48246 (N_48246,N_41622,N_40609);
nand U48247 (N_48247,N_43048,N_44680);
or U48248 (N_48248,N_43718,N_43402);
nand U48249 (N_48249,N_42892,N_41120);
or U48250 (N_48250,N_43281,N_40867);
or U48251 (N_48251,N_41947,N_41159);
and U48252 (N_48252,N_41443,N_40705);
nor U48253 (N_48253,N_41528,N_44596);
xor U48254 (N_48254,N_43682,N_41875);
xnor U48255 (N_48255,N_42137,N_44734);
nor U48256 (N_48256,N_43206,N_42956);
or U48257 (N_48257,N_44821,N_42159);
or U48258 (N_48258,N_40066,N_43128);
xnor U48259 (N_48259,N_44278,N_43989);
nand U48260 (N_48260,N_44092,N_40321);
nor U48261 (N_48261,N_42201,N_43853);
nor U48262 (N_48262,N_42570,N_40447);
or U48263 (N_48263,N_41755,N_43498);
or U48264 (N_48264,N_43270,N_43420);
and U48265 (N_48265,N_43561,N_44643);
and U48266 (N_48266,N_41493,N_41548);
and U48267 (N_48267,N_41237,N_44438);
and U48268 (N_48268,N_41161,N_42808);
xnor U48269 (N_48269,N_44124,N_43124);
and U48270 (N_48270,N_44911,N_41173);
xnor U48271 (N_48271,N_44977,N_43487);
nor U48272 (N_48272,N_44820,N_41804);
xor U48273 (N_48273,N_42157,N_43014);
nor U48274 (N_48274,N_43884,N_41623);
and U48275 (N_48275,N_44171,N_44425);
nand U48276 (N_48276,N_42852,N_40151);
and U48277 (N_48277,N_40580,N_44586);
xnor U48278 (N_48278,N_42175,N_40120);
nand U48279 (N_48279,N_41423,N_44262);
or U48280 (N_48280,N_42391,N_41805);
or U48281 (N_48281,N_41043,N_43781);
nand U48282 (N_48282,N_40110,N_42110);
or U48283 (N_48283,N_42332,N_42623);
xnor U48284 (N_48284,N_42210,N_41621);
nand U48285 (N_48285,N_40254,N_42819);
and U48286 (N_48286,N_40467,N_41755);
or U48287 (N_48287,N_41201,N_44304);
or U48288 (N_48288,N_41087,N_43363);
xnor U48289 (N_48289,N_43553,N_43618);
xor U48290 (N_48290,N_44827,N_40733);
nand U48291 (N_48291,N_40451,N_44101);
nand U48292 (N_48292,N_40947,N_43459);
or U48293 (N_48293,N_43536,N_40357);
and U48294 (N_48294,N_41479,N_43045);
or U48295 (N_48295,N_41525,N_41725);
xnor U48296 (N_48296,N_44881,N_40665);
or U48297 (N_48297,N_43183,N_40182);
or U48298 (N_48298,N_42536,N_41673);
and U48299 (N_48299,N_43006,N_44929);
nor U48300 (N_48300,N_40875,N_41827);
nand U48301 (N_48301,N_43771,N_44129);
xor U48302 (N_48302,N_43503,N_41213);
or U48303 (N_48303,N_43133,N_40970);
and U48304 (N_48304,N_40103,N_42183);
nand U48305 (N_48305,N_44454,N_41696);
xor U48306 (N_48306,N_44463,N_44198);
xor U48307 (N_48307,N_40807,N_43913);
nor U48308 (N_48308,N_44653,N_40671);
nand U48309 (N_48309,N_43857,N_42699);
or U48310 (N_48310,N_44919,N_40670);
nor U48311 (N_48311,N_40289,N_41184);
nand U48312 (N_48312,N_41570,N_44907);
or U48313 (N_48313,N_41964,N_44011);
xnor U48314 (N_48314,N_43933,N_42559);
or U48315 (N_48315,N_42696,N_42143);
nor U48316 (N_48316,N_41961,N_44114);
xnor U48317 (N_48317,N_41521,N_42517);
xnor U48318 (N_48318,N_43077,N_40876);
nand U48319 (N_48319,N_42220,N_42764);
or U48320 (N_48320,N_42013,N_41229);
nor U48321 (N_48321,N_41076,N_44920);
nand U48322 (N_48322,N_44726,N_42339);
nand U48323 (N_48323,N_42359,N_44733);
and U48324 (N_48324,N_41585,N_41276);
nand U48325 (N_48325,N_41237,N_43437);
nor U48326 (N_48326,N_40075,N_43844);
and U48327 (N_48327,N_42552,N_43950);
nor U48328 (N_48328,N_43450,N_42162);
or U48329 (N_48329,N_44568,N_40549);
or U48330 (N_48330,N_43548,N_40148);
or U48331 (N_48331,N_42132,N_44933);
and U48332 (N_48332,N_44556,N_43754);
or U48333 (N_48333,N_44058,N_42573);
or U48334 (N_48334,N_42954,N_43261);
and U48335 (N_48335,N_40780,N_40159);
nor U48336 (N_48336,N_42785,N_41521);
nor U48337 (N_48337,N_40940,N_42384);
and U48338 (N_48338,N_42504,N_42824);
and U48339 (N_48339,N_41706,N_41431);
or U48340 (N_48340,N_41476,N_42988);
or U48341 (N_48341,N_40421,N_40899);
or U48342 (N_48342,N_41564,N_44485);
xor U48343 (N_48343,N_43155,N_41990);
and U48344 (N_48344,N_44049,N_44213);
xnor U48345 (N_48345,N_40497,N_43583);
nor U48346 (N_48346,N_40013,N_44170);
xnor U48347 (N_48347,N_41170,N_42350);
or U48348 (N_48348,N_42775,N_43500);
nand U48349 (N_48349,N_40350,N_43224);
nand U48350 (N_48350,N_44862,N_44095);
nor U48351 (N_48351,N_42437,N_41729);
and U48352 (N_48352,N_44429,N_42034);
or U48353 (N_48353,N_42298,N_41642);
xnor U48354 (N_48354,N_44857,N_40648);
xor U48355 (N_48355,N_43933,N_40261);
and U48356 (N_48356,N_42783,N_43294);
nor U48357 (N_48357,N_42331,N_40861);
and U48358 (N_48358,N_41361,N_42938);
or U48359 (N_48359,N_44183,N_43225);
xor U48360 (N_48360,N_44080,N_40927);
nand U48361 (N_48361,N_42595,N_40294);
nand U48362 (N_48362,N_44132,N_40547);
nand U48363 (N_48363,N_44973,N_44249);
xnor U48364 (N_48364,N_40294,N_41548);
xor U48365 (N_48365,N_40218,N_44592);
and U48366 (N_48366,N_43697,N_41470);
or U48367 (N_48367,N_41488,N_42272);
nand U48368 (N_48368,N_42306,N_42018);
nand U48369 (N_48369,N_40456,N_42257);
nor U48370 (N_48370,N_43506,N_41141);
nor U48371 (N_48371,N_44634,N_42531);
nor U48372 (N_48372,N_44892,N_42857);
xnor U48373 (N_48373,N_40372,N_41095);
and U48374 (N_48374,N_41813,N_43292);
nand U48375 (N_48375,N_44155,N_43379);
nand U48376 (N_48376,N_40587,N_41927);
and U48377 (N_48377,N_44798,N_42888);
xnor U48378 (N_48378,N_43913,N_42427);
or U48379 (N_48379,N_44830,N_41350);
and U48380 (N_48380,N_42677,N_40074);
nor U48381 (N_48381,N_41195,N_44453);
nor U48382 (N_48382,N_44592,N_42735);
xor U48383 (N_48383,N_43035,N_42820);
nand U48384 (N_48384,N_44032,N_42504);
nand U48385 (N_48385,N_44143,N_41088);
nor U48386 (N_48386,N_43515,N_44648);
and U48387 (N_48387,N_43165,N_41342);
nand U48388 (N_48388,N_43458,N_43927);
or U48389 (N_48389,N_43729,N_44200);
or U48390 (N_48390,N_41559,N_43961);
nand U48391 (N_48391,N_41262,N_40490);
or U48392 (N_48392,N_43095,N_40285);
nor U48393 (N_48393,N_40973,N_40113);
nand U48394 (N_48394,N_41957,N_42464);
xnor U48395 (N_48395,N_40039,N_41067);
or U48396 (N_48396,N_44743,N_44683);
nand U48397 (N_48397,N_40332,N_41239);
or U48398 (N_48398,N_40840,N_41555);
nand U48399 (N_48399,N_42139,N_44370);
xor U48400 (N_48400,N_41539,N_40927);
xor U48401 (N_48401,N_44249,N_43822);
and U48402 (N_48402,N_43737,N_40754);
nor U48403 (N_48403,N_42981,N_40808);
xor U48404 (N_48404,N_41526,N_43050);
and U48405 (N_48405,N_44984,N_42302);
nor U48406 (N_48406,N_42007,N_42454);
or U48407 (N_48407,N_43528,N_41189);
xnor U48408 (N_48408,N_41432,N_42739);
and U48409 (N_48409,N_41506,N_44351);
and U48410 (N_48410,N_40008,N_41292);
nor U48411 (N_48411,N_43256,N_42786);
and U48412 (N_48412,N_43772,N_42883);
nand U48413 (N_48413,N_42892,N_44593);
nor U48414 (N_48414,N_41223,N_44678);
or U48415 (N_48415,N_44937,N_43782);
or U48416 (N_48416,N_43236,N_41000);
and U48417 (N_48417,N_42552,N_42651);
xor U48418 (N_48418,N_40694,N_43794);
and U48419 (N_48419,N_43077,N_41185);
or U48420 (N_48420,N_40066,N_43955);
nand U48421 (N_48421,N_40270,N_44422);
nand U48422 (N_48422,N_42240,N_40121);
and U48423 (N_48423,N_44949,N_40580);
or U48424 (N_48424,N_41221,N_43840);
nor U48425 (N_48425,N_44396,N_43057);
nand U48426 (N_48426,N_42762,N_42554);
xnor U48427 (N_48427,N_43765,N_44913);
nand U48428 (N_48428,N_44067,N_42711);
nand U48429 (N_48429,N_43691,N_44378);
and U48430 (N_48430,N_40903,N_42443);
and U48431 (N_48431,N_44404,N_44968);
xnor U48432 (N_48432,N_41003,N_40488);
or U48433 (N_48433,N_41186,N_41086);
nand U48434 (N_48434,N_44698,N_44139);
nand U48435 (N_48435,N_40108,N_41936);
or U48436 (N_48436,N_43086,N_44657);
and U48437 (N_48437,N_41905,N_42141);
and U48438 (N_48438,N_44546,N_42323);
nor U48439 (N_48439,N_44081,N_41189);
nand U48440 (N_48440,N_43805,N_40143);
nand U48441 (N_48441,N_41163,N_40828);
and U48442 (N_48442,N_43354,N_44388);
nor U48443 (N_48443,N_41487,N_42940);
and U48444 (N_48444,N_42708,N_41232);
or U48445 (N_48445,N_42882,N_42898);
or U48446 (N_48446,N_44190,N_43538);
xor U48447 (N_48447,N_41582,N_43951);
and U48448 (N_48448,N_41195,N_42583);
nand U48449 (N_48449,N_44713,N_41638);
and U48450 (N_48450,N_43544,N_43048);
nand U48451 (N_48451,N_40498,N_44878);
xnor U48452 (N_48452,N_41803,N_42797);
nor U48453 (N_48453,N_41101,N_42555);
and U48454 (N_48454,N_42333,N_42275);
xnor U48455 (N_48455,N_44808,N_44818);
and U48456 (N_48456,N_41471,N_41132);
or U48457 (N_48457,N_42728,N_42117);
and U48458 (N_48458,N_44628,N_44493);
nor U48459 (N_48459,N_43859,N_43490);
nand U48460 (N_48460,N_41156,N_44734);
and U48461 (N_48461,N_43102,N_40450);
or U48462 (N_48462,N_44851,N_43885);
xor U48463 (N_48463,N_40550,N_42977);
and U48464 (N_48464,N_43751,N_40511);
nor U48465 (N_48465,N_40847,N_44093);
nand U48466 (N_48466,N_42370,N_42096);
nand U48467 (N_48467,N_43112,N_41387);
or U48468 (N_48468,N_41280,N_43388);
xnor U48469 (N_48469,N_41633,N_41806);
and U48470 (N_48470,N_42976,N_42972);
nor U48471 (N_48471,N_40468,N_43942);
or U48472 (N_48472,N_42741,N_40484);
or U48473 (N_48473,N_41140,N_40729);
and U48474 (N_48474,N_43465,N_42959);
nor U48475 (N_48475,N_42022,N_44767);
or U48476 (N_48476,N_44642,N_41447);
nand U48477 (N_48477,N_40664,N_41748);
nor U48478 (N_48478,N_44918,N_41148);
nor U48479 (N_48479,N_40401,N_44209);
and U48480 (N_48480,N_44460,N_40617);
xor U48481 (N_48481,N_43498,N_40021);
and U48482 (N_48482,N_40038,N_44574);
or U48483 (N_48483,N_44168,N_41936);
xor U48484 (N_48484,N_40655,N_43407);
or U48485 (N_48485,N_41966,N_42722);
nand U48486 (N_48486,N_44915,N_43148);
and U48487 (N_48487,N_43821,N_41609);
and U48488 (N_48488,N_42228,N_43713);
and U48489 (N_48489,N_44770,N_40291);
or U48490 (N_48490,N_41349,N_41399);
nand U48491 (N_48491,N_44957,N_43487);
nand U48492 (N_48492,N_42596,N_43377);
and U48493 (N_48493,N_43434,N_44274);
or U48494 (N_48494,N_42628,N_41914);
nand U48495 (N_48495,N_42288,N_44624);
xor U48496 (N_48496,N_40576,N_44576);
or U48497 (N_48497,N_42132,N_40188);
or U48498 (N_48498,N_42413,N_41745);
and U48499 (N_48499,N_41411,N_43011);
and U48500 (N_48500,N_44561,N_40723);
xor U48501 (N_48501,N_44931,N_43266);
xor U48502 (N_48502,N_41486,N_41792);
or U48503 (N_48503,N_43755,N_40501);
xor U48504 (N_48504,N_44826,N_43851);
nand U48505 (N_48505,N_43808,N_43530);
and U48506 (N_48506,N_41911,N_44127);
or U48507 (N_48507,N_44931,N_41725);
or U48508 (N_48508,N_40945,N_43536);
nor U48509 (N_48509,N_41971,N_42921);
nand U48510 (N_48510,N_40506,N_44632);
nor U48511 (N_48511,N_43104,N_40864);
nand U48512 (N_48512,N_40326,N_44567);
and U48513 (N_48513,N_42748,N_42929);
or U48514 (N_48514,N_44944,N_43606);
nand U48515 (N_48515,N_42115,N_40650);
nor U48516 (N_48516,N_40220,N_40707);
and U48517 (N_48517,N_44218,N_40127);
nand U48518 (N_48518,N_41199,N_44174);
nor U48519 (N_48519,N_44805,N_43044);
and U48520 (N_48520,N_40388,N_42363);
and U48521 (N_48521,N_44538,N_42318);
nor U48522 (N_48522,N_42349,N_40423);
nor U48523 (N_48523,N_40758,N_43282);
xnor U48524 (N_48524,N_40427,N_41146);
and U48525 (N_48525,N_41439,N_41576);
and U48526 (N_48526,N_41189,N_44692);
nand U48527 (N_48527,N_41438,N_42593);
nand U48528 (N_48528,N_41205,N_42967);
nand U48529 (N_48529,N_43415,N_44959);
nand U48530 (N_48530,N_40869,N_43176);
xnor U48531 (N_48531,N_41411,N_43286);
or U48532 (N_48532,N_41030,N_43111);
nor U48533 (N_48533,N_40549,N_40032);
or U48534 (N_48534,N_41966,N_41977);
xor U48535 (N_48535,N_44874,N_44277);
or U48536 (N_48536,N_42139,N_43365);
and U48537 (N_48537,N_40356,N_40084);
nor U48538 (N_48538,N_41435,N_43899);
and U48539 (N_48539,N_41019,N_40562);
or U48540 (N_48540,N_43469,N_42650);
nand U48541 (N_48541,N_43481,N_40038);
or U48542 (N_48542,N_40525,N_42452);
xnor U48543 (N_48543,N_44220,N_44150);
and U48544 (N_48544,N_43059,N_40467);
xnor U48545 (N_48545,N_43267,N_44601);
nand U48546 (N_48546,N_43953,N_43207);
nor U48547 (N_48547,N_40506,N_41845);
xor U48548 (N_48548,N_43242,N_40643);
or U48549 (N_48549,N_44862,N_44490);
and U48550 (N_48550,N_40280,N_41697);
xnor U48551 (N_48551,N_44585,N_43832);
and U48552 (N_48552,N_41387,N_40106);
nand U48553 (N_48553,N_43413,N_43050);
or U48554 (N_48554,N_43187,N_40978);
and U48555 (N_48555,N_41495,N_40291);
and U48556 (N_48556,N_43104,N_42765);
nand U48557 (N_48557,N_42612,N_44652);
nand U48558 (N_48558,N_43491,N_40641);
xnor U48559 (N_48559,N_43258,N_40792);
xnor U48560 (N_48560,N_40958,N_43702);
or U48561 (N_48561,N_41640,N_41588);
xnor U48562 (N_48562,N_43956,N_41260);
nor U48563 (N_48563,N_40326,N_41336);
nand U48564 (N_48564,N_41595,N_44304);
nor U48565 (N_48565,N_42574,N_40156);
xnor U48566 (N_48566,N_43229,N_44350);
xnor U48567 (N_48567,N_43617,N_43678);
or U48568 (N_48568,N_43687,N_42136);
nor U48569 (N_48569,N_41575,N_41394);
and U48570 (N_48570,N_42415,N_41049);
or U48571 (N_48571,N_41534,N_40142);
and U48572 (N_48572,N_41339,N_44254);
nand U48573 (N_48573,N_44559,N_40524);
or U48574 (N_48574,N_42876,N_40614);
or U48575 (N_48575,N_40994,N_43416);
xor U48576 (N_48576,N_41111,N_43475);
and U48577 (N_48577,N_43696,N_41016);
nand U48578 (N_48578,N_40454,N_43248);
xor U48579 (N_48579,N_41196,N_42020);
nor U48580 (N_48580,N_43855,N_40965);
nor U48581 (N_48581,N_42298,N_41086);
nor U48582 (N_48582,N_42492,N_42166);
nand U48583 (N_48583,N_44225,N_41659);
nor U48584 (N_48584,N_44438,N_43777);
nor U48585 (N_48585,N_42224,N_44023);
and U48586 (N_48586,N_40948,N_44819);
and U48587 (N_48587,N_42758,N_40081);
and U48588 (N_48588,N_40213,N_42514);
nor U48589 (N_48589,N_43610,N_42272);
xnor U48590 (N_48590,N_43998,N_40800);
or U48591 (N_48591,N_42333,N_41693);
or U48592 (N_48592,N_43006,N_40045);
nand U48593 (N_48593,N_41788,N_40573);
and U48594 (N_48594,N_41041,N_43465);
and U48595 (N_48595,N_40484,N_43644);
and U48596 (N_48596,N_42175,N_40383);
or U48597 (N_48597,N_40435,N_44211);
and U48598 (N_48598,N_44884,N_40861);
and U48599 (N_48599,N_41945,N_40632);
or U48600 (N_48600,N_43640,N_43916);
nor U48601 (N_48601,N_42897,N_40688);
nand U48602 (N_48602,N_43288,N_43310);
xor U48603 (N_48603,N_43198,N_42525);
nand U48604 (N_48604,N_43374,N_42688);
xor U48605 (N_48605,N_44849,N_44328);
nor U48606 (N_48606,N_41801,N_42551);
nand U48607 (N_48607,N_43414,N_40747);
xnor U48608 (N_48608,N_42493,N_41731);
or U48609 (N_48609,N_41528,N_43777);
and U48610 (N_48610,N_40110,N_43526);
nand U48611 (N_48611,N_44422,N_43501);
nor U48612 (N_48612,N_43349,N_44857);
nand U48613 (N_48613,N_40313,N_41825);
or U48614 (N_48614,N_44600,N_41475);
xnor U48615 (N_48615,N_44766,N_43186);
nand U48616 (N_48616,N_41800,N_43414);
nor U48617 (N_48617,N_41407,N_41256);
nand U48618 (N_48618,N_40926,N_43833);
nand U48619 (N_48619,N_43149,N_40656);
nor U48620 (N_48620,N_42563,N_43661);
nand U48621 (N_48621,N_44554,N_44644);
nor U48622 (N_48622,N_41323,N_41046);
nand U48623 (N_48623,N_42450,N_41806);
and U48624 (N_48624,N_40023,N_42427);
or U48625 (N_48625,N_41797,N_40522);
nand U48626 (N_48626,N_44256,N_40606);
or U48627 (N_48627,N_41075,N_43872);
nor U48628 (N_48628,N_42164,N_41618);
nor U48629 (N_48629,N_42688,N_42537);
nand U48630 (N_48630,N_40565,N_44161);
or U48631 (N_48631,N_41105,N_40607);
nand U48632 (N_48632,N_43971,N_42483);
nand U48633 (N_48633,N_43488,N_41195);
or U48634 (N_48634,N_44475,N_43538);
or U48635 (N_48635,N_42658,N_44937);
or U48636 (N_48636,N_42173,N_40350);
xnor U48637 (N_48637,N_42742,N_43037);
xnor U48638 (N_48638,N_43801,N_44323);
and U48639 (N_48639,N_42951,N_41340);
and U48640 (N_48640,N_40969,N_44630);
and U48641 (N_48641,N_41803,N_42366);
xnor U48642 (N_48642,N_42814,N_43244);
or U48643 (N_48643,N_40829,N_44836);
nor U48644 (N_48644,N_40679,N_44995);
and U48645 (N_48645,N_42155,N_41232);
nand U48646 (N_48646,N_44979,N_44931);
nand U48647 (N_48647,N_42529,N_42596);
nand U48648 (N_48648,N_43975,N_42338);
or U48649 (N_48649,N_44832,N_43745);
or U48650 (N_48650,N_41326,N_42499);
and U48651 (N_48651,N_42027,N_42256);
xor U48652 (N_48652,N_40560,N_41885);
nand U48653 (N_48653,N_43744,N_40856);
or U48654 (N_48654,N_44720,N_41382);
xnor U48655 (N_48655,N_40659,N_40770);
xnor U48656 (N_48656,N_40781,N_42539);
xnor U48657 (N_48657,N_44589,N_41560);
nand U48658 (N_48658,N_42587,N_43985);
or U48659 (N_48659,N_41344,N_43860);
or U48660 (N_48660,N_41505,N_43831);
and U48661 (N_48661,N_43164,N_44444);
or U48662 (N_48662,N_42956,N_40185);
xnor U48663 (N_48663,N_42620,N_44237);
or U48664 (N_48664,N_42653,N_44217);
nand U48665 (N_48665,N_41581,N_44319);
and U48666 (N_48666,N_43214,N_44728);
nor U48667 (N_48667,N_40288,N_44877);
xnor U48668 (N_48668,N_44785,N_42320);
or U48669 (N_48669,N_40226,N_43560);
xor U48670 (N_48670,N_43641,N_40989);
nor U48671 (N_48671,N_42908,N_43582);
nand U48672 (N_48672,N_41722,N_42127);
or U48673 (N_48673,N_42359,N_44622);
xor U48674 (N_48674,N_44367,N_40340);
nand U48675 (N_48675,N_43801,N_41865);
nor U48676 (N_48676,N_43237,N_43239);
and U48677 (N_48677,N_40816,N_44323);
nand U48678 (N_48678,N_43636,N_40100);
or U48679 (N_48679,N_42266,N_44370);
or U48680 (N_48680,N_41765,N_40081);
and U48681 (N_48681,N_42191,N_40335);
or U48682 (N_48682,N_40221,N_44587);
nand U48683 (N_48683,N_43529,N_43231);
or U48684 (N_48684,N_44427,N_43604);
nand U48685 (N_48685,N_40825,N_42018);
and U48686 (N_48686,N_40330,N_44476);
nand U48687 (N_48687,N_42156,N_42363);
and U48688 (N_48688,N_40651,N_44496);
xnor U48689 (N_48689,N_41245,N_42504);
xor U48690 (N_48690,N_42888,N_44204);
nand U48691 (N_48691,N_42273,N_43637);
nand U48692 (N_48692,N_40248,N_42359);
or U48693 (N_48693,N_44940,N_41953);
and U48694 (N_48694,N_41272,N_44025);
or U48695 (N_48695,N_42900,N_43070);
or U48696 (N_48696,N_40345,N_40657);
nand U48697 (N_48697,N_44821,N_44848);
nand U48698 (N_48698,N_41529,N_44700);
and U48699 (N_48699,N_40146,N_44904);
nand U48700 (N_48700,N_43751,N_41125);
xor U48701 (N_48701,N_40418,N_41803);
or U48702 (N_48702,N_40475,N_43492);
and U48703 (N_48703,N_44627,N_43415);
nor U48704 (N_48704,N_41408,N_40920);
xor U48705 (N_48705,N_44661,N_43895);
and U48706 (N_48706,N_43789,N_44671);
xor U48707 (N_48707,N_43231,N_40936);
or U48708 (N_48708,N_42384,N_40665);
nor U48709 (N_48709,N_43588,N_44765);
xnor U48710 (N_48710,N_40890,N_43433);
or U48711 (N_48711,N_42149,N_44515);
xnor U48712 (N_48712,N_43967,N_43146);
nor U48713 (N_48713,N_42195,N_44008);
xor U48714 (N_48714,N_40621,N_42558);
or U48715 (N_48715,N_44071,N_40749);
nor U48716 (N_48716,N_42312,N_41421);
nor U48717 (N_48717,N_41160,N_42741);
nor U48718 (N_48718,N_41144,N_43029);
or U48719 (N_48719,N_42373,N_42953);
nor U48720 (N_48720,N_41992,N_42704);
xnor U48721 (N_48721,N_44891,N_41358);
nor U48722 (N_48722,N_44302,N_42503);
xor U48723 (N_48723,N_40440,N_40030);
nor U48724 (N_48724,N_44100,N_43715);
or U48725 (N_48725,N_42371,N_43209);
and U48726 (N_48726,N_44859,N_40982);
nand U48727 (N_48727,N_42040,N_41430);
xor U48728 (N_48728,N_40644,N_40058);
nand U48729 (N_48729,N_43760,N_42294);
nand U48730 (N_48730,N_44568,N_40181);
and U48731 (N_48731,N_43910,N_44360);
nand U48732 (N_48732,N_44782,N_42019);
xor U48733 (N_48733,N_43797,N_42092);
xor U48734 (N_48734,N_43899,N_43030);
xor U48735 (N_48735,N_43757,N_44851);
nor U48736 (N_48736,N_44543,N_44767);
nand U48737 (N_48737,N_40653,N_42309);
xor U48738 (N_48738,N_42950,N_41801);
xor U48739 (N_48739,N_41702,N_43797);
or U48740 (N_48740,N_40058,N_41805);
nand U48741 (N_48741,N_41555,N_40624);
and U48742 (N_48742,N_42013,N_44529);
or U48743 (N_48743,N_43926,N_41088);
and U48744 (N_48744,N_42668,N_40728);
or U48745 (N_48745,N_44580,N_42623);
xnor U48746 (N_48746,N_40148,N_42036);
nand U48747 (N_48747,N_40201,N_44552);
or U48748 (N_48748,N_43394,N_41659);
xnor U48749 (N_48749,N_44719,N_41207);
nand U48750 (N_48750,N_42958,N_40009);
or U48751 (N_48751,N_42789,N_44695);
or U48752 (N_48752,N_43119,N_40442);
and U48753 (N_48753,N_41819,N_43027);
nand U48754 (N_48754,N_44164,N_42612);
nor U48755 (N_48755,N_44435,N_43893);
xor U48756 (N_48756,N_44360,N_41924);
xor U48757 (N_48757,N_42064,N_41352);
nor U48758 (N_48758,N_42832,N_42283);
and U48759 (N_48759,N_40922,N_41739);
or U48760 (N_48760,N_41772,N_40171);
nor U48761 (N_48761,N_41784,N_44136);
nor U48762 (N_48762,N_40203,N_42735);
xor U48763 (N_48763,N_43417,N_42379);
and U48764 (N_48764,N_40509,N_40652);
nand U48765 (N_48765,N_40517,N_41683);
and U48766 (N_48766,N_43261,N_42570);
xnor U48767 (N_48767,N_44290,N_41570);
and U48768 (N_48768,N_41691,N_43991);
or U48769 (N_48769,N_43516,N_41527);
or U48770 (N_48770,N_40104,N_42634);
nand U48771 (N_48771,N_42088,N_41914);
or U48772 (N_48772,N_40850,N_42274);
nor U48773 (N_48773,N_41616,N_41940);
nand U48774 (N_48774,N_44812,N_42052);
nor U48775 (N_48775,N_41077,N_41641);
nor U48776 (N_48776,N_44139,N_43035);
and U48777 (N_48777,N_43481,N_42510);
nand U48778 (N_48778,N_41601,N_42294);
or U48779 (N_48779,N_40091,N_41835);
nor U48780 (N_48780,N_43444,N_44255);
xor U48781 (N_48781,N_42464,N_44640);
and U48782 (N_48782,N_42897,N_44765);
xnor U48783 (N_48783,N_43603,N_44552);
xor U48784 (N_48784,N_43703,N_40980);
xor U48785 (N_48785,N_40082,N_42341);
nand U48786 (N_48786,N_43482,N_41412);
and U48787 (N_48787,N_40649,N_44391);
or U48788 (N_48788,N_44884,N_43813);
nand U48789 (N_48789,N_40427,N_43222);
nand U48790 (N_48790,N_43390,N_42627);
or U48791 (N_48791,N_44082,N_44822);
and U48792 (N_48792,N_40725,N_40839);
xnor U48793 (N_48793,N_40964,N_40007);
or U48794 (N_48794,N_44912,N_44157);
xnor U48795 (N_48795,N_40762,N_43268);
or U48796 (N_48796,N_40226,N_40862);
nor U48797 (N_48797,N_43393,N_42422);
xnor U48798 (N_48798,N_41559,N_40087);
xor U48799 (N_48799,N_43648,N_40275);
or U48800 (N_48800,N_44712,N_41122);
or U48801 (N_48801,N_40035,N_42860);
and U48802 (N_48802,N_40377,N_44213);
nand U48803 (N_48803,N_42731,N_43218);
nor U48804 (N_48804,N_43774,N_43110);
or U48805 (N_48805,N_40769,N_41909);
nand U48806 (N_48806,N_40849,N_44290);
nand U48807 (N_48807,N_43252,N_43857);
nor U48808 (N_48808,N_40525,N_42049);
or U48809 (N_48809,N_41374,N_41006);
and U48810 (N_48810,N_42477,N_40965);
and U48811 (N_48811,N_43034,N_43989);
or U48812 (N_48812,N_40769,N_42061);
or U48813 (N_48813,N_40638,N_43260);
nand U48814 (N_48814,N_41590,N_44531);
nand U48815 (N_48815,N_44712,N_41956);
nor U48816 (N_48816,N_41563,N_43849);
or U48817 (N_48817,N_40949,N_41613);
and U48818 (N_48818,N_43789,N_41110);
or U48819 (N_48819,N_42050,N_41758);
nand U48820 (N_48820,N_44622,N_41582);
nand U48821 (N_48821,N_42544,N_44529);
nand U48822 (N_48822,N_44882,N_43812);
nand U48823 (N_48823,N_42768,N_40080);
xnor U48824 (N_48824,N_44979,N_40843);
nand U48825 (N_48825,N_42248,N_41452);
xor U48826 (N_48826,N_43882,N_41548);
or U48827 (N_48827,N_40577,N_41621);
xnor U48828 (N_48828,N_43096,N_41637);
xnor U48829 (N_48829,N_44763,N_44636);
nor U48830 (N_48830,N_40512,N_44766);
and U48831 (N_48831,N_44216,N_41296);
xor U48832 (N_48832,N_42098,N_44232);
xnor U48833 (N_48833,N_41387,N_43083);
and U48834 (N_48834,N_43188,N_41693);
and U48835 (N_48835,N_42054,N_42885);
and U48836 (N_48836,N_43466,N_40201);
nor U48837 (N_48837,N_44414,N_44748);
and U48838 (N_48838,N_42545,N_42882);
or U48839 (N_48839,N_42185,N_41819);
nand U48840 (N_48840,N_40103,N_40329);
xor U48841 (N_48841,N_43396,N_41123);
and U48842 (N_48842,N_41879,N_44451);
nor U48843 (N_48843,N_42881,N_44785);
nand U48844 (N_48844,N_41639,N_41119);
and U48845 (N_48845,N_42319,N_43084);
xnor U48846 (N_48846,N_40792,N_42569);
and U48847 (N_48847,N_40704,N_41640);
or U48848 (N_48848,N_44597,N_42933);
or U48849 (N_48849,N_43635,N_41717);
and U48850 (N_48850,N_43554,N_43794);
or U48851 (N_48851,N_40133,N_42315);
and U48852 (N_48852,N_42060,N_42805);
nor U48853 (N_48853,N_42595,N_44431);
nor U48854 (N_48854,N_41861,N_41546);
xor U48855 (N_48855,N_41997,N_40554);
nand U48856 (N_48856,N_42556,N_42886);
xor U48857 (N_48857,N_44145,N_43363);
nor U48858 (N_48858,N_41404,N_40905);
xor U48859 (N_48859,N_43768,N_42076);
and U48860 (N_48860,N_43798,N_41360);
xnor U48861 (N_48861,N_43367,N_41477);
and U48862 (N_48862,N_41499,N_44580);
xnor U48863 (N_48863,N_42363,N_42909);
nor U48864 (N_48864,N_43054,N_43654);
and U48865 (N_48865,N_40767,N_42621);
nor U48866 (N_48866,N_40725,N_42316);
xnor U48867 (N_48867,N_42438,N_43138);
xor U48868 (N_48868,N_42298,N_42008);
and U48869 (N_48869,N_41714,N_44663);
nand U48870 (N_48870,N_41334,N_40761);
or U48871 (N_48871,N_42356,N_43138);
nand U48872 (N_48872,N_40923,N_43217);
or U48873 (N_48873,N_40964,N_44643);
nand U48874 (N_48874,N_42460,N_43483);
xnor U48875 (N_48875,N_41161,N_41727);
nand U48876 (N_48876,N_43022,N_42341);
nor U48877 (N_48877,N_43934,N_42466);
xnor U48878 (N_48878,N_40600,N_42095);
and U48879 (N_48879,N_43598,N_44982);
and U48880 (N_48880,N_43969,N_42154);
nor U48881 (N_48881,N_43964,N_41045);
or U48882 (N_48882,N_41511,N_42487);
nand U48883 (N_48883,N_42060,N_43027);
or U48884 (N_48884,N_41739,N_41785);
or U48885 (N_48885,N_40752,N_41742);
xor U48886 (N_48886,N_42630,N_42053);
or U48887 (N_48887,N_42780,N_42483);
xnor U48888 (N_48888,N_43375,N_43408);
or U48889 (N_48889,N_41254,N_41913);
or U48890 (N_48890,N_44867,N_41689);
and U48891 (N_48891,N_42235,N_42543);
or U48892 (N_48892,N_40842,N_42609);
nor U48893 (N_48893,N_44811,N_43893);
nand U48894 (N_48894,N_42765,N_43163);
or U48895 (N_48895,N_41279,N_42811);
or U48896 (N_48896,N_42696,N_44418);
xnor U48897 (N_48897,N_43143,N_43738);
or U48898 (N_48898,N_43327,N_42180);
and U48899 (N_48899,N_43377,N_42928);
and U48900 (N_48900,N_44578,N_42902);
nor U48901 (N_48901,N_42149,N_41491);
nand U48902 (N_48902,N_44701,N_41442);
and U48903 (N_48903,N_42678,N_43675);
nor U48904 (N_48904,N_44637,N_43722);
nor U48905 (N_48905,N_43160,N_41024);
or U48906 (N_48906,N_44987,N_43824);
nand U48907 (N_48907,N_40721,N_40762);
or U48908 (N_48908,N_40331,N_40570);
or U48909 (N_48909,N_41019,N_41163);
and U48910 (N_48910,N_44850,N_41711);
nand U48911 (N_48911,N_43609,N_43716);
xor U48912 (N_48912,N_41969,N_43405);
xnor U48913 (N_48913,N_44031,N_43488);
nor U48914 (N_48914,N_43834,N_41438);
nand U48915 (N_48915,N_42491,N_40844);
xnor U48916 (N_48916,N_41012,N_44954);
and U48917 (N_48917,N_40740,N_42587);
and U48918 (N_48918,N_43571,N_40324);
xor U48919 (N_48919,N_44149,N_42338);
nand U48920 (N_48920,N_43229,N_42482);
nor U48921 (N_48921,N_40024,N_40557);
nor U48922 (N_48922,N_42966,N_43388);
nand U48923 (N_48923,N_43355,N_44518);
nor U48924 (N_48924,N_40722,N_43615);
and U48925 (N_48925,N_43056,N_42961);
xnor U48926 (N_48926,N_44908,N_41406);
nor U48927 (N_48927,N_42415,N_43938);
and U48928 (N_48928,N_42419,N_44138);
nand U48929 (N_48929,N_41256,N_41424);
and U48930 (N_48930,N_44466,N_43060);
or U48931 (N_48931,N_42753,N_41897);
xor U48932 (N_48932,N_42572,N_41821);
and U48933 (N_48933,N_44366,N_43408);
xnor U48934 (N_48934,N_41204,N_44622);
or U48935 (N_48935,N_44867,N_42978);
nand U48936 (N_48936,N_44099,N_41304);
and U48937 (N_48937,N_41820,N_41242);
or U48938 (N_48938,N_43338,N_43597);
nor U48939 (N_48939,N_42888,N_41448);
xor U48940 (N_48940,N_41925,N_43079);
xnor U48941 (N_48941,N_42784,N_40653);
and U48942 (N_48942,N_42552,N_43888);
xor U48943 (N_48943,N_41949,N_42063);
or U48944 (N_48944,N_44575,N_40045);
xor U48945 (N_48945,N_43898,N_42077);
and U48946 (N_48946,N_40610,N_40961);
nand U48947 (N_48947,N_40656,N_43018);
or U48948 (N_48948,N_44412,N_43072);
and U48949 (N_48949,N_40891,N_42231);
or U48950 (N_48950,N_40369,N_40064);
nand U48951 (N_48951,N_44283,N_43882);
nand U48952 (N_48952,N_43954,N_42663);
and U48953 (N_48953,N_40970,N_41083);
xor U48954 (N_48954,N_41461,N_40848);
xnor U48955 (N_48955,N_44007,N_44217);
or U48956 (N_48956,N_44705,N_44058);
nand U48957 (N_48957,N_44213,N_43582);
nor U48958 (N_48958,N_43325,N_42996);
and U48959 (N_48959,N_41396,N_40197);
and U48960 (N_48960,N_44428,N_40776);
nor U48961 (N_48961,N_42229,N_43300);
nor U48962 (N_48962,N_43152,N_42057);
nor U48963 (N_48963,N_41406,N_40077);
and U48964 (N_48964,N_42330,N_41262);
nor U48965 (N_48965,N_43963,N_40536);
xnor U48966 (N_48966,N_43623,N_42400);
nand U48967 (N_48967,N_42551,N_42347);
nor U48968 (N_48968,N_43502,N_43151);
xnor U48969 (N_48969,N_44658,N_42155);
nor U48970 (N_48970,N_44235,N_43548);
xnor U48971 (N_48971,N_41475,N_40167);
nor U48972 (N_48972,N_42075,N_42125);
nor U48973 (N_48973,N_44951,N_44426);
xor U48974 (N_48974,N_42377,N_42548);
and U48975 (N_48975,N_40963,N_43764);
nor U48976 (N_48976,N_43951,N_42598);
xor U48977 (N_48977,N_41538,N_40713);
xnor U48978 (N_48978,N_41359,N_43198);
or U48979 (N_48979,N_42083,N_44030);
or U48980 (N_48980,N_42487,N_40035);
nor U48981 (N_48981,N_41857,N_40561);
nand U48982 (N_48982,N_41265,N_43186);
nor U48983 (N_48983,N_41965,N_42376);
or U48984 (N_48984,N_40696,N_42049);
nor U48985 (N_48985,N_41110,N_42759);
and U48986 (N_48986,N_40686,N_41966);
nor U48987 (N_48987,N_40229,N_42639);
nor U48988 (N_48988,N_43627,N_41192);
nand U48989 (N_48989,N_40909,N_41298);
xor U48990 (N_48990,N_41356,N_42877);
and U48991 (N_48991,N_43347,N_42815);
and U48992 (N_48992,N_41618,N_40697);
and U48993 (N_48993,N_42647,N_43565);
and U48994 (N_48994,N_44458,N_43303);
nor U48995 (N_48995,N_43863,N_42406);
and U48996 (N_48996,N_42541,N_41588);
xnor U48997 (N_48997,N_44029,N_43746);
and U48998 (N_48998,N_41652,N_41446);
nand U48999 (N_48999,N_42912,N_42849);
nand U49000 (N_49000,N_42114,N_43234);
xor U49001 (N_49001,N_41669,N_42252);
or U49002 (N_49002,N_42362,N_42128);
or U49003 (N_49003,N_44427,N_43412);
nor U49004 (N_49004,N_40452,N_40725);
or U49005 (N_49005,N_43530,N_41085);
nor U49006 (N_49006,N_42494,N_44294);
xnor U49007 (N_49007,N_44925,N_41378);
or U49008 (N_49008,N_42915,N_43358);
xor U49009 (N_49009,N_40443,N_42399);
and U49010 (N_49010,N_43053,N_42852);
and U49011 (N_49011,N_42251,N_41202);
nor U49012 (N_49012,N_41359,N_44448);
nor U49013 (N_49013,N_41569,N_43832);
xor U49014 (N_49014,N_42690,N_40702);
nand U49015 (N_49015,N_42613,N_40791);
xnor U49016 (N_49016,N_44178,N_42856);
or U49017 (N_49017,N_42113,N_40897);
nor U49018 (N_49018,N_42976,N_42136);
or U49019 (N_49019,N_44855,N_41899);
xnor U49020 (N_49020,N_44181,N_41760);
xor U49021 (N_49021,N_44224,N_44449);
xor U49022 (N_49022,N_43492,N_42258);
nand U49023 (N_49023,N_42869,N_41239);
and U49024 (N_49024,N_44657,N_42678);
nand U49025 (N_49025,N_40695,N_42255);
or U49026 (N_49026,N_43256,N_41828);
and U49027 (N_49027,N_44884,N_41723);
or U49028 (N_49028,N_44900,N_44268);
or U49029 (N_49029,N_40590,N_42111);
xnor U49030 (N_49030,N_40724,N_41349);
nor U49031 (N_49031,N_40948,N_44640);
nor U49032 (N_49032,N_44531,N_43659);
nand U49033 (N_49033,N_43490,N_42774);
nand U49034 (N_49034,N_43007,N_43477);
nor U49035 (N_49035,N_41934,N_40073);
nand U49036 (N_49036,N_44455,N_43459);
and U49037 (N_49037,N_41169,N_43826);
and U49038 (N_49038,N_43492,N_41087);
nor U49039 (N_49039,N_44304,N_43651);
nor U49040 (N_49040,N_43391,N_40664);
or U49041 (N_49041,N_40142,N_41441);
or U49042 (N_49042,N_40076,N_41773);
or U49043 (N_49043,N_44218,N_41907);
or U49044 (N_49044,N_43776,N_41832);
or U49045 (N_49045,N_43840,N_44912);
nor U49046 (N_49046,N_41475,N_44664);
xor U49047 (N_49047,N_44500,N_44472);
nor U49048 (N_49048,N_40897,N_41157);
xor U49049 (N_49049,N_40198,N_42207);
and U49050 (N_49050,N_44660,N_43206);
nor U49051 (N_49051,N_42829,N_42700);
xnor U49052 (N_49052,N_44024,N_40502);
xnor U49053 (N_49053,N_43388,N_43082);
nand U49054 (N_49054,N_43472,N_43821);
nor U49055 (N_49055,N_42550,N_44878);
xnor U49056 (N_49056,N_41173,N_41667);
nor U49057 (N_49057,N_42516,N_44151);
nand U49058 (N_49058,N_41447,N_40162);
and U49059 (N_49059,N_43465,N_43249);
xor U49060 (N_49060,N_41914,N_43815);
and U49061 (N_49061,N_43006,N_44169);
nor U49062 (N_49062,N_41016,N_41746);
or U49063 (N_49063,N_43889,N_41606);
nor U49064 (N_49064,N_41434,N_43102);
nand U49065 (N_49065,N_40090,N_43228);
and U49066 (N_49066,N_44588,N_40594);
or U49067 (N_49067,N_43391,N_40329);
and U49068 (N_49068,N_40528,N_40680);
nand U49069 (N_49069,N_44102,N_40358);
xnor U49070 (N_49070,N_44119,N_40388);
and U49071 (N_49071,N_40820,N_43992);
and U49072 (N_49072,N_40617,N_41391);
or U49073 (N_49073,N_42267,N_42178);
xor U49074 (N_49074,N_44062,N_43517);
xnor U49075 (N_49075,N_44913,N_42617);
xor U49076 (N_49076,N_40197,N_42843);
or U49077 (N_49077,N_42218,N_43542);
nand U49078 (N_49078,N_41478,N_42298);
and U49079 (N_49079,N_41813,N_41876);
nor U49080 (N_49080,N_40781,N_40350);
nor U49081 (N_49081,N_44649,N_43847);
nand U49082 (N_49082,N_40986,N_42711);
nor U49083 (N_49083,N_44929,N_41317);
or U49084 (N_49084,N_41622,N_40386);
nand U49085 (N_49085,N_42696,N_43046);
nor U49086 (N_49086,N_41703,N_42644);
nand U49087 (N_49087,N_43791,N_44697);
or U49088 (N_49088,N_43681,N_40152);
xor U49089 (N_49089,N_41167,N_42201);
nand U49090 (N_49090,N_41662,N_43198);
nor U49091 (N_49091,N_41890,N_40590);
xor U49092 (N_49092,N_42984,N_42548);
xor U49093 (N_49093,N_42383,N_40177);
xnor U49094 (N_49094,N_43246,N_41982);
xnor U49095 (N_49095,N_42377,N_40063);
nor U49096 (N_49096,N_40305,N_42942);
xnor U49097 (N_49097,N_43707,N_41385);
nor U49098 (N_49098,N_42879,N_44981);
xor U49099 (N_49099,N_41385,N_43372);
and U49100 (N_49100,N_43219,N_40466);
xor U49101 (N_49101,N_44929,N_44639);
nor U49102 (N_49102,N_44282,N_42948);
and U49103 (N_49103,N_42125,N_42204);
nand U49104 (N_49104,N_40962,N_41273);
and U49105 (N_49105,N_40272,N_40219);
xnor U49106 (N_49106,N_43313,N_41097);
and U49107 (N_49107,N_40142,N_40955);
or U49108 (N_49108,N_40042,N_42468);
xnor U49109 (N_49109,N_40164,N_41081);
xnor U49110 (N_49110,N_43880,N_42511);
or U49111 (N_49111,N_44775,N_40242);
and U49112 (N_49112,N_41779,N_42102);
xnor U49113 (N_49113,N_43155,N_44659);
nand U49114 (N_49114,N_44373,N_42669);
xnor U49115 (N_49115,N_44547,N_44783);
nand U49116 (N_49116,N_41008,N_44843);
nor U49117 (N_49117,N_43539,N_43642);
and U49118 (N_49118,N_41663,N_43863);
xnor U49119 (N_49119,N_42680,N_43801);
nand U49120 (N_49120,N_43582,N_40517);
nand U49121 (N_49121,N_40038,N_43513);
or U49122 (N_49122,N_40657,N_44801);
nor U49123 (N_49123,N_43126,N_41346);
or U49124 (N_49124,N_44600,N_41278);
and U49125 (N_49125,N_40060,N_42499);
xor U49126 (N_49126,N_44688,N_40485);
xor U49127 (N_49127,N_43021,N_44620);
and U49128 (N_49128,N_43335,N_41341);
xor U49129 (N_49129,N_44802,N_43093);
and U49130 (N_49130,N_43248,N_40324);
or U49131 (N_49131,N_44538,N_41643);
xor U49132 (N_49132,N_40956,N_44005);
nor U49133 (N_49133,N_43944,N_42579);
xnor U49134 (N_49134,N_42041,N_40744);
nand U49135 (N_49135,N_40625,N_41827);
and U49136 (N_49136,N_41083,N_44326);
nor U49137 (N_49137,N_43255,N_43312);
xor U49138 (N_49138,N_44868,N_44537);
xor U49139 (N_49139,N_44123,N_43764);
or U49140 (N_49140,N_43243,N_41569);
or U49141 (N_49141,N_43243,N_41158);
nand U49142 (N_49142,N_41509,N_40696);
or U49143 (N_49143,N_44576,N_41636);
and U49144 (N_49144,N_44644,N_44476);
and U49145 (N_49145,N_44337,N_43765);
nand U49146 (N_49146,N_40467,N_41573);
nor U49147 (N_49147,N_42831,N_44090);
xnor U49148 (N_49148,N_43183,N_43497);
or U49149 (N_49149,N_41245,N_41260);
and U49150 (N_49150,N_43617,N_40290);
xor U49151 (N_49151,N_43680,N_41059);
xnor U49152 (N_49152,N_41243,N_44128);
nor U49153 (N_49153,N_42546,N_42210);
nor U49154 (N_49154,N_44493,N_42015);
or U49155 (N_49155,N_41818,N_42632);
xor U49156 (N_49156,N_42242,N_43533);
and U49157 (N_49157,N_43690,N_41419);
xnor U49158 (N_49158,N_42927,N_42526);
xnor U49159 (N_49159,N_42333,N_42673);
nand U49160 (N_49160,N_44276,N_41695);
nand U49161 (N_49161,N_44390,N_41128);
nand U49162 (N_49162,N_41145,N_44452);
and U49163 (N_49163,N_41361,N_41056);
nor U49164 (N_49164,N_40580,N_41251);
and U49165 (N_49165,N_43312,N_44568);
and U49166 (N_49166,N_40585,N_44894);
nand U49167 (N_49167,N_42209,N_43899);
nor U49168 (N_49168,N_41880,N_44819);
nand U49169 (N_49169,N_40792,N_42014);
and U49170 (N_49170,N_41306,N_44491);
nor U49171 (N_49171,N_41988,N_42915);
nand U49172 (N_49172,N_40654,N_41338);
or U49173 (N_49173,N_40849,N_41607);
xor U49174 (N_49174,N_41609,N_42076);
xnor U49175 (N_49175,N_43898,N_42042);
xnor U49176 (N_49176,N_41304,N_44191);
nand U49177 (N_49177,N_43479,N_43044);
nand U49178 (N_49178,N_42371,N_41489);
nand U49179 (N_49179,N_40060,N_41765);
or U49180 (N_49180,N_43782,N_43879);
nand U49181 (N_49181,N_44223,N_42201);
xnor U49182 (N_49182,N_43437,N_42705);
xor U49183 (N_49183,N_43845,N_41174);
nand U49184 (N_49184,N_44479,N_42848);
nor U49185 (N_49185,N_41399,N_44217);
xnor U49186 (N_49186,N_42775,N_42721);
and U49187 (N_49187,N_43449,N_43157);
xnor U49188 (N_49188,N_40250,N_40709);
xor U49189 (N_49189,N_41514,N_41921);
and U49190 (N_49190,N_42856,N_44054);
nor U49191 (N_49191,N_41421,N_40470);
nor U49192 (N_49192,N_44246,N_41239);
nor U49193 (N_49193,N_43165,N_42235);
or U49194 (N_49194,N_41406,N_42859);
or U49195 (N_49195,N_44859,N_43022);
nand U49196 (N_49196,N_42319,N_40938);
xnor U49197 (N_49197,N_40283,N_41583);
nand U49198 (N_49198,N_44903,N_42790);
or U49199 (N_49199,N_42149,N_41720);
and U49200 (N_49200,N_40820,N_43016);
and U49201 (N_49201,N_41718,N_43946);
nand U49202 (N_49202,N_43772,N_43668);
or U49203 (N_49203,N_40495,N_41457);
nand U49204 (N_49204,N_44954,N_41923);
and U49205 (N_49205,N_40063,N_41786);
nor U49206 (N_49206,N_42980,N_42422);
xor U49207 (N_49207,N_44116,N_40441);
xor U49208 (N_49208,N_43860,N_42918);
xor U49209 (N_49209,N_43489,N_42406);
nor U49210 (N_49210,N_40869,N_42218);
xor U49211 (N_49211,N_43671,N_42443);
nor U49212 (N_49212,N_41445,N_42213);
nor U49213 (N_49213,N_40813,N_41956);
or U49214 (N_49214,N_43062,N_42429);
and U49215 (N_49215,N_40885,N_42997);
xor U49216 (N_49216,N_41258,N_44293);
xor U49217 (N_49217,N_44533,N_44725);
or U49218 (N_49218,N_41570,N_40252);
xor U49219 (N_49219,N_41204,N_44243);
nand U49220 (N_49220,N_42165,N_43472);
or U49221 (N_49221,N_42250,N_40011);
nor U49222 (N_49222,N_44151,N_41592);
nand U49223 (N_49223,N_44593,N_40812);
or U49224 (N_49224,N_42590,N_41720);
nand U49225 (N_49225,N_41333,N_41291);
and U49226 (N_49226,N_40746,N_41295);
nand U49227 (N_49227,N_44287,N_41047);
xnor U49228 (N_49228,N_44487,N_40036);
or U49229 (N_49229,N_40783,N_41891);
and U49230 (N_49230,N_41105,N_44624);
nand U49231 (N_49231,N_43102,N_44942);
or U49232 (N_49232,N_40332,N_43799);
nand U49233 (N_49233,N_43218,N_44839);
nand U49234 (N_49234,N_43693,N_44369);
nand U49235 (N_49235,N_43068,N_43127);
nor U49236 (N_49236,N_43577,N_43930);
nand U49237 (N_49237,N_44544,N_42947);
nor U49238 (N_49238,N_43190,N_41522);
nand U49239 (N_49239,N_41380,N_40840);
nand U49240 (N_49240,N_40037,N_40248);
nand U49241 (N_49241,N_42000,N_42269);
xor U49242 (N_49242,N_42431,N_41096);
or U49243 (N_49243,N_43351,N_44578);
xnor U49244 (N_49244,N_40953,N_43057);
and U49245 (N_49245,N_43038,N_40534);
nand U49246 (N_49246,N_42862,N_42168);
nand U49247 (N_49247,N_44742,N_43343);
xor U49248 (N_49248,N_41059,N_42076);
and U49249 (N_49249,N_43790,N_43112);
nor U49250 (N_49250,N_42553,N_43383);
and U49251 (N_49251,N_40841,N_40607);
or U49252 (N_49252,N_41400,N_41888);
nand U49253 (N_49253,N_41711,N_42385);
nor U49254 (N_49254,N_41169,N_44499);
xor U49255 (N_49255,N_41895,N_44538);
xnor U49256 (N_49256,N_42750,N_40859);
xor U49257 (N_49257,N_40784,N_41719);
and U49258 (N_49258,N_41461,N_42230);
nand U49259 (N_49259,N_43634,N_44715);
and U49260 (N_49260,N_42399,N_40550);
nand U49261 (N_49261,N_40762,N_41493);
and U49262 (N_49262,N_40831,N_42456);
or U49263 (N_49263,N_44160,N_40294);
nor U49264 (N_49264,N_40111,N_42369);
or U49265 (N_49265,N_43242,N_40559);
nand U49266 (N_49266,N_44833,N_40606);
or U49267 (N_49267,N_41786,N_42866);
xnor U49268 (N_49268,N_43438,N_44841);
xnor U49269 (N_49269,N_41741,N_44772);
and U49270 (N_49270,N_42723,N_41983);
nand U49271 (N_49271,N_40676,N_41472);
and U49272 (N_49272,N_42324,N_41888);
nor U49273 (N_49273,N_40990,N_41868);
or U49274 (N_49274,N_40627,N_40711);
nor U49275 (N_49275,N_44117,N_40245);
and U49276 (N_49276,N_44542,N_42066);
and U49277 (N_49277,N_43591,N_42105);
or U49278 (N_49278,N_43347,N_42314);
xor U49279 (N_49279,N_43469,N_43914);
xnor U49280 (N_49280,N_42156,N_41517);
nor U49281 (N_49281,N_43227,N_40580);
and U49282 (N_49282,N_42496,N_40357);
or U49283 (N_49283,N_43838,N_41032);
or U49284 (N_49284,N_40201,N_44184);
xor U49285 (N_49285,N_43987,N_43589);
or U49286 (N_49286,N_42682,N_42478);
and U49287 (N_49287,N_44511,N_44800);
and U49288 (N_49288,N_43581,N_40751);
or U49289 (N_49289,N_40547,N_41655);
xor U49290 (N_49290,N_42556,N_41268);
nor U49291 (N_49291,N_42202,N_42778);
xor U49292 (N_49292,N_41677,N_44588);
nor U49293 (N_49293,N_43164,N_41845);
nand U49294 (N_49294,N_44914,N_44116);
and U49295 (N_49295,N_44650,N_42928);
xor U49296 (N_49296,N_42047,N_40577);
and U49297 (N_49297,N_40366,N_43656);
and U49298 (N_49298,N_44040,N_43199);
or U49299 (N_49299,N_43734,N_42005);
nand U49300 (N_49300,N_42938,N_43424);
and U49301 (N_49301,N_41722,N_41742);
and U49302 (N_49302,N_43069,N_40494);
nor U49303 (N_49303,N_44720,N_42486);
or U49304 (N_49304,N_41812,N_43698);
or U49305 (N_49305,N_40077,N_41792);
nand U49306 (N_49306,N_40766,N_41183);
nor U49307 (N_49307,N_40831,N_43890);
or U49308 (N_49308,N_43572,N_41273);
or U49309 (N_49309,N_44136,N_42455);
nand U49310 (N_49310,N_40528,N_41962);
nand U49311 (N_49311,N_40384,N_43541);
xnor U49312 (N_49312,N_42552,N_42116);
and U49313 (N_49313,N_40847,N_44688);
and U49314 (N_49314,N_44366,N_41854);
or U49315 (N_49315,N_43360,N_41559);
or U49316 (N_49316,N_41873,N_41844);
nor U49317 (N_49317,N_40023,N_44623);
xnor U49318 (N_49318,N_42213,N_40276);
nand U49319 (N_49319,N_41907,N_44911);
and U49320 (N_49320,N_43656,N_40720);
and U49321 (N_49321,N_44019,N_40184);
and U49322 (N_49322,N_41569,N_42025);
or U49323 (N_49323,N_40618,N_42323);
and U49324 (N_49324,N_41242,N_40629);
or U49325 (N_49325,N_42535,N_44825);
or U49326 (N_49326,N_40733,N_44215);
nor U49327 (N_49327,N_44619,N_43429);
and U49328 (N_49328,N_43694,N_40367);
nand U49329 (N_49329,N_41635,N_41670);
nand U49330 (N_49330,N_40716,N_42594);
or U49331 (N_49331,N_43727,N_42349);
nor U49332 (N_49332,N_43365,N_42967);
xnor U49333 (N_49333,N_43316,N_40554);
nand U49334 (N_49334,N_42867,N_41281);
nor U49335 (N_49335,N_40464,N_43010);
or U49336 (N_49336,N_40108,N_44263);
or U49337 (N_49337,N_43441,N_43863);
xnor U49338 (N_49338,N_41060,N_43280);
or U49339 (N_49339,N_43741,N_41762);
nor U49340 (N_49340,N_44332,N_42798);
nor U49341 (N_49341,N_41330,N_43914);
and U49342 (N_49342,N_42732,N_41763);
and U49343 (N_49343,N_44013,N_41220);
and U49344 (N_49344,N_42900,N_41615);
nand U49345 (N_49345,N_43103,N_44812);
or U49346 (N_49346,N_40351,N_44193);
or U49347 (N_49347,N_41387,N_44058);
nand U49348 (N_49348,N_44245,N_41290);
or U49349 (N_49349,N_43015,N_44914);
and U49350 (N_49350,N_41470,N_40744);
or U49351 (N_49351,N_42885,N_44606);
or U49352 (N_49352,N_42601,N_42502);
nand U49353 (N_49353,N_43292,N_41141);
xnor U49354 (N_49354,N_44561,N_41980);
nor U49355 (N_49355,N_40047,N_41121);
nor U49356 (N_49356,N_42686,N_42217);
and U49357 (N_49357,N_42908,N_41715);
nand U49358 (N_49358,N_41760,N_44897);
nand U49359 (N_49359,N_41346,N_44039);
nor U49360 (N_49360,N_42872,N_41232);
xor U49361 (N_49361,N_44187,N_43154);
xor U49362 (N_49362,N_41322,N_41546);
or U49363 (N_49363,N_44923,N_40250);
nand U49364 (N_49364,N_40756,N_41046);
nor U49365 (N_49365,N_44692,N_42231);
nor U49366 (N_49366,N_44085,N_43089);
nand U49367 (N_49367,N_40093,N_44436);
xor U49368 (N_49368,N_42534,N_41220);
nor U49369 (N_49369,N_42065,N_43806);
nor U49370 (N_49370,N_40832,N_43181);
nand U49371 (N_49371,N_41164,N_42148);
xor U49372 (N_49372,N_44251,N_44419);
or U49373 (N_49373,N_40169,N_43914);
xor U49374 (N_49374,N_41808,N_42815);
xnor U49375 (N_49375,N_40228,N_43206);
or U49376 (N_49376,N_44223,N_43887);
nor U49377 (N_49377,N_41231,N_44919);
xor U49378 (N_49378,N_42063,N_44763);
or U49379 (N_49379,N_41932,N_40242);
nor U49380 (N_49380,N_42982,N_41624);
nand U49381 (N_49381,N_42492,N_40836);
xor U49382 (N_49382,N_40858,N_41866);
xnor U49383 (N_49383,N_41015,N_42389);
and U49384 (N_49384,N_41146,N_43893);
or U49385 (N_49385,N_44226,N_40101);
nand U49386 (N_49386,N_43301,N_44209);
nand U49387 (N_49387,N_41506,N_43600);
xor U49388 (N_49388,N_42624,N_42079);
xor U49389 (N_49389,N_43481,N_40070);
and U49390 (N_49390,N_44411,N_43684);
nand U49391 (N_49391,N_44867,N_43720);
or U49392 (N_49392,N_43137,N_40828);
xor U49393 (N_49393,N_44226,N_43941);
or U49394 (N_49394,N_42034,N_44359);
nand U49395 (N_49395,N_42275,N_42687);
nor U49396 (N_49396,N_42358,N_44535);
or U49397 (N_49397,N_43087,N_40260);
or U49398 (N_49398,N_42066,N_44508);
nor U49399 (N_49399,N_42885,N_44137);
xnor U49400 (N_49400,N_44251,N_42005);
xor U49401 (N_49401,N_40409,N_41160);
and U49402 (N_49402,N_40371,N_41978);
or U49403 (N_49403,N_42315,N_43937);
nand U49404 (N_49404,N_42018,N_41304);
nand U49405 (N_49405,N_40984,N_41609);
nor U49406 (N_49406,N_44197,N_41431);
xor U49407 (N_49407,N_42462,N_43285);
nand U49408 (N_49408,N_40383,N_42073);
and U49409 (N_49409,N_44968,N_43198);
xor U49410 (N_49410,N_42357,N_41322);
nor U49411 (N_49411,N_44642,N_43177);
nand U49412 (N_49412,N_41269,N_41411);
or U49413 (N_49413,N_41631,N_41292);
xor U49414 (N_49414,N_41367,N_41031);
xor U49415 (N_49415,N_41817,N_41183);
and U49416 (N_49416,N_40737,N_42788);
nor U49417 (N_49417,N_44075,N_40492);
xor U49418 (N_49418,N_42557,N_42843);
or U49419 (N_49419,N_44495,N_42673);
and U49420 (N_49420,N_40896,N_43617);
nand U49421 (N_49421,N_42580,N_44598);
or U49422 (N_49422,N_44007,N_41051);
nor U49423 (N_49423,N_43165,N_44945);
or U49424 (N_49424,N_40755,N_44589);
or U49425 (N_49425,N_41560,N_43772);
or U49426 (N_49426,N_44624,N_40185);
and U49427 (N_49427,N_42805,N_43450);
xnor U49428 (N_49428,N_42870,N_40705);
xor U49429 (N_49429,N_41981,N_43357);
xor U49430 (N_49430,N_43164,N_44942);
nand U49431 (N_49431,N_42253,N_43796);
nand U49432 (N_49432,N_44416,N_41365);
and U49433 (N_49433,N_40138,N_42720);
nand U49434 (N_49434,N_44416,N_44031);
and U49435 (N_49435,N_40377,N_43526);
xor U49436 (N_49436,N_43018,N_43615);
nor U49437 (N_49437,N_44989,N_41145);
nand U49438 (N_49438,N_41500,N_42921);
xnor U49439 (N_49439,N_40408,N_41398);
xor U49440 (N_49440,N_44837,N_41444);
and U49441 (N_49441,N_44022,N_42709);
nor U49442 (N_49442,N_43219,N_42101);
and U49443 (N_49443,N_42256,N_41293);
nor U49444 (N_49444,N_40191,N_40629);
xnor U49445 (N_49445,N_41113,N_40502);
nand U49446 (N_49446,N_44185,N_43771);
or U49447 (N_49447,N_43458,N_40524);
xnor U49448 (N_49448,N_40441,N_44742);
nor U49449 (N_49449,N_44792,N_43265);
or U49450 (N_49450,N_42548,N_44816);
nor U49451 (N_49451,N_40562,N_43480);
nand U49452 (N_49452,N_44221,N_40188);
nor U49453 (N_49453,N_40358,N_44442);
xnor U49454 (N_49454,N_42322,N_40430);
xnor U49455 (N_49455,N_44900,N_40459);
or U49456 (N_49456,N_41384,N_40555);
nor U49457 (N_49457,N_42772,N_41711);
or U49458 (N_49458,N_43394,N_41002);
xnor U49459 (N_49459,N_42302,N_43031);
or U49460 (N_49460,N_42077,N_41225);
or U49461 (N_49461,N_40323,N_41031);
and U49462 (N_49462,N_43066,N_43196);
or U49463 (N_49463,N_42711,N_44409);
or U49464 (N_49464,N_40188,N_41868);
and U49465 (N_49465,N_43478,N_41493);
xor U49466 (N_49466,N_42154,N_43756);
nor U49467 (N_49467,N_43786,N_43224);
or U49468 (N_49468,N_40006,N_40209);
nand U49469 (N_49469,N_41408,N_44656);
and U49470 (N_49470,N_41798,N_42523);
nand U49471 (N_49471,N_42880,N_44073);
xor U49472 (N_49472,N_41742,N_44652);
xnor U49473 (N_49473,N_44731,N_42095);
and U49474 (N_49474,N_43746,N_41163);
or U49475 (N_49475,N_41487,N_42563);
nand U49476 (N_49476,N_41839,N_41787);
or U49477 (N_49477,N_40262,N_43700);
and U49478 (N_49478,N_43058,N_42435);
nand U49479 (N_49479,N_40494,N_42687);
xnor U49480 (N_49480,N_44985,N_43490);
or U49481 (N_49481,N_44384,N_40384);
and U49482 (N_49482,N_43923,N_41339);
and U49483 (N_49483,N_41735,N_41540);
nand U49484 (N_49484,N_42598,N_42833);
nor U49485 (N_49485,N_41184,N_44366);
or U49486 (N_49486,N_44130,N_42422);
nor U49487 (N_49487,N_41729,N_41343);
and U49488 (N_49488,N_42648,N_41416);
or U49489 (N_49489,N_42195,N_41095);
nand U49490 (N_49490,N_40819,N_44408);
nor U49491 (N_49491,N_44652,N_40850);
nor U49492 (N_49492,N_41428,N_44118);
nor U49493 (N_49493,N_41554,N_42070);
or U49494 (N_49494,N_40401,N_44419);
xnor U49495 (N_49495,N_44360,N_40826);
xnor U49496 (N_49496,N_41948,N_43918);
nand U49497 (N_49497,N_40771,N_42873);
or U49498 (N_49498,N_42896,N_43815);
nand U49499 (N_49499,N_41559,N_42368);
or U49500 (N_49500,N_42946,N_42943);
and U49501 (N_49501,N_44758,N_41081);
or U49502 (N_49502,N_41351,N_40896);
nor U49503 (N_49503,N_42045,N_40732);
or U49504 (N_49504,N_42530,N_44843);
xor U49505 (N_49505,N_44038,N_42329);
nand U49506 (N_49506,N_42270,N_42285);
or U49507 (N_49507,N_44146,N_43077);
nor U49508 (N_49508,N_40298,N_40573);
xnor U49509 (N_49509,N_41092,N_42156);
and U49510 (N_49510,N_44434,N_42063);
nor U49511 (N_49511,N_44080,N_43342);
nand U49512 (N_49512,N_42988,N_40586);
nand U49513 (N_49513,N_40392,N_42648);
and U49514 (N_49514,N_41444,N_41093);
nand U49515 (N_49515,N_41586,N_41561);
or U49516 (N_49516,N_43519,N_44940);
xor U49517 (N_49517,N_41825,N_43828);
or U49518 (N_49518,N_43897,N_40457);
or U49519 (N_49519,N_42096,N_44214);
nor U49520 (N_49520,N_40181,N_40451);
nor U49521 (N_49521,N_40053,N_43165);
and U49522 (N_49522,N_40592,N_40947);
xor U49523 (N_49523,N_43851,N_43326);
nor U49524 (N_49524,N_42152,N_41678);
xnor U49525 (N_49525,N_42779,N_40152);
nor U49526 (N_49526,N_43031,N_44856);
xnor U49527 (N_49527,N_44124,N_41728);
xnor U49528 (N_49528,N_44415,N_41623);
nor U49529 (N_49529,N_41593,N_43188);
or U49530 (N_49530,N_42085,N_44038);
or U49531 (N_49531,N_40118,N_40513);
or U49532 (N_49532,N_43237,N_44111);
xor U49533 (N_49533,N_42108,N_42325);
nor U49534 (N_49534,N_41185,N_40778);
nor U49535 (N_49535,N_41538,N_44234);
nor U49536 (N_49536,N_42769,N_40179);
nor U49537 (N_49537,N_40401,N_41221);
xor U49538 (N_49538,N_40403,N_40801);
and U49539 (N_49539,N_40038,N_43312);
nand U49540 (N_49540,N_42627,N_42479);
nand U49541 (N_49541,N_43003,N_40625);
and U49542 (N_49542,N_42146,N_42156);
nand U49543 (N_49543,N_40507,N_43989);
nand U49544 (N_49544,N_42405,N_43106);
nand U49545 (N_49545,N_42969,N_44805);
xor U49546 (N_49546,N_43343,N_44852);
and U49547 (N_49547,N_42933,N_41810);
and U49548 (N_49548,N_44626,N_44835);
nand U49549 (N_49549,N_44123,N_42662);
and U49550 (N_49550,N_41959,N_41584);
and U49551 (N_49551,N_41364,N_40768);
xnor U49552 (N_49552,N_42824,N_41303);
and U49553 (N_49553,N_43034,N_44035);
nand U49554 (N_49554,N_41421,N_43204);
nor U49555 (N_49555,N_43815,N_41825);
or U49556 (N_49556,N_40127,N_42392);
nor U49557 (N_49557,N_41571,N_44949);
xnor U49558 (N_49558,N_42422,N_42784);
or U49559 (N_49559,N_41989,N_42555);
nor U49560 (N_49560,N_41745,N_41370);
and U49561 (N_49561,N_44773,N_41943);
nand U49562 (N_49562,N_41861,N_43394);
xnor U49563 (N_49563,N_40928,N_43511);
or U49564 (N_49564,N_41311,N_40085);
nand U49565 (N_49565,N_44942,N_42067);
nand U49566 (N_49566,N_41854,N_41257);
xor U49567 (N_49567,N_43813,N_41008);
nor U49568 (N_49568,N_44132,N_42467);
or U49569 (N_49569,N_42380,N_43343);
nand U49570 (N_49570,N_43379,N_42232);
nor U49571 (N_49571,N_42115,N_44177);
or U49572 (N_49572,N_41855,N_41184);
and U49573 (N_49573,N_40654,N_42907);
nor U49574 (N_49574,N_44233,N_43738);
or U49575 (N_49575,N_42148,N_41337);
xor U49576 (N_49576,N_43011,N_40133);
nor U49577 (N_49577,N_44540,N_43084);
nand U49578 (N_49578,N_41516,N_43027);
xor U49579 (N_49579,N_44289,N_44254);
or U49580 (N_49580,N_40669,N_40689);
or U49581 (N_49581,N_44017,N_42354);
xnor U49582 (N_49582,N_44166,N_41230);
xnor U49583 (N_49583,N_44346,N_40789);
and U49584 (N_49584,N_43976,N_44072);
and U49585 (N_49585,N_44598,N_43459);
nand U49586 (N_49586,N_41093,N_41947);
nor U49587 (N_49587,N_40228,N_42202);
or U49588 (N_49588,N_40353,N_40041);
xor U49589 (N_49589,N_43206,N_41204);
nand U49590 (N_49590,N_40449,N_44008);
nor U49591 (N_49591,N_44180,N_43294);
nor U49592 (N_49592,N_40728,N_43536);
xnor U49593 (N_49593,N_44841,N_41737);
and U49594 (N_49594,N_40852,N_42255);
or U49595 (N_49595,N_41213,N_42030);
nor U49596 (N_49596,N_41603,N_44290);
nand U49597 (N_49597,N_44694,N_42411);
and U49598 (N_49598,N_41009,N_41299);
nor U49599 (N_49599,N_42600,N_43092);
or U49600 (N_49600,N_41562,N_43889);
xnor U49601 (N_49601,N_41292,N_44119);
or U49602 (N_49602,N_44221,N_41933);
xor U49603 (N_49603,N_41154,N_44432);
nand U49604 (N_49604,N_42575,N_43571);
nor U49605 (N_49605,N_40810,N_42298);
and U49606 (N_49606,N_44585,N_40782);
nor U49607 (N_49607,N_43531,N_41949);
xor U49608 (N_49608,N_42552,N_40951);
or U49609 (N_49609,N_43082,N_40012);
nand U49610 (N_49610,N_44802,N_43408);
nand U49611 (N_49611,N_41085,N_43522);
nand U49612 (N_49612,N_40546,N_40982);
nor U49613 (N_49613,N_40639,N_43305);
nor U49614 (N_49614,N_40133,N_40425);
nand U49615 (N_49615,N_40571,N_43516);
nand U49616 (N_49616,N_42403,N_43766);
xor U49617 (N_49617,N_42647,N_43751);
xor U49618 (N_49618,N_41760,N_43167);
nor U49619 (N_49619,N_41255,N_42190);
xor U49620 (N_49620,N_40447,N_42624);
nor U49621 (N_49621,N_41330,N_42589);
xor U49622 (N_49622,N_40436,N_42310);
nor U49623 (N_49623,N_42568,N_44426);
xnor U49624 (N_49624,N_44032,N_41807);
xor U49625 (N_49625,N_43931,N_42233);
and U49626 (N_49626,N_41870,N_42024);
nand U49627 (N_49627,N_42498,N_44107);
xor U49628 (N_49628,N_43079,N_40123);
xor U49629 (N_49629,N_41813,N_42052);
nand U49630 (N_49630,N_43635,N_44413);
nor U49631 (N_49631,N_40767,N_41954);
nor U49632 (N_49632,N_42572,N_44763);
or U49633 (N_49633,N_43271,N_41812);
and U49634 (N_49634,N_44734,N_43958);
xnor U49635 (N_49635,N_42374,N_44949);
nand U49636 (N_49636,N_41715,N_44120);
or U49637 (N_49637,N_43430,N_40997);
nor U49638 (N_49638,N_41574,N_43866);
xnor U49639 (N_49639,N_40791,N_43556);
or U49640 (N_49640,N_42891,N_42149);
nand U49641 (N_49641,N_43164,N_43257);
nand U49642 (N_49642,N_40234,N_41389);
nand U49643 (N_49643,N_43878,N_40749);
and U49644 (N_49644,N_40561,N_40014);
or U49645 (N_49645,N_43342,N_44865);
nand U49646 (N_49646,N_41390,N_43382);
and U49647 (N_49647,N_44818,N_44196);
xnor U49648 (N_49648,N_40271,N_42433);
nor U49649 (N_49649,N_44117,N_42312);
xor U49650 (N_49650,N_44528,N_43438);
nor U49651 (N_49651,N_43778,N_43598);
or U49652 (N_49652,N_44641,N_44226);
nand U49653 (N_49653,N_41067,N_40652);
xor U49654 (N_49654,N_44294,N_44983);
nand U49655 (N_49655,N_40702,N_41771);
and U49656 (N_49656,N_40816,N_40856);
xnor U49657 (N_49657,N_40321,N_40731);
xor U49658 (N_49658,N_40439,N_43200);
or U49659 (N_49659,N_41307,N_42083);
or U49660 (N_49660,N_41235,N_40662);
or U49661 (N_49661,N_41855,N_44970);
nand U49662 (N_49662,N_44618,N_40519);
or U49663 (N_49663,N_41765,N_43509);
xnor U49664 (N_49664,N_43862,N_40031);
and U49665 (N_49665,N_44726,N_41958);
or U49666 (N_49666,N_42377,N_40937);
and U49667 (N_49667,N_44332,N_44033);
nand U49668 (N_49668,N_43368,N_44481);
nor U49669 (N_49669,N_41749,N_41653);
and U49670 (N_49670,N_40872,N_41290);
xor U49671 (N_49671,N_41478,N_42253);
xor U49672 (N_49672,N_43245,N_41888);
nand U49673 (N_49673,N_42091,N_40292);
xor U49674 (N_49674,N_40379,N_41366);
and U49675 (N_49675,N_42267,N_42304);
and U49676 (N_49676,N_44472,N_42982);
nor U49677 (N_49677,N_41177,N_43242);
nand U49678 (N_49678,N_41892,N_44682);
or U49679 (N_49679,N_43979,N_42849);
nand U49680 (N_49680,N_43928,N_43286);
nand U49681 (N_49681,N_40509,N_41895);
and U49682 (N_49682,N_42320,N_41928);
nor U49683 (N_49683,N_44304,N_40905);
and U49684 (N_49684,N_41457,N_41591);
or U49685 (N_49685,N_41113,N_44206);
nor U49686 (N_49686,N_41352,N_40113);
nor U49687 (N_49687,N_41493,N_44837);
and U49688 (N_49688,N_40998,N_42633);
and U49689 (N_49689,N_40175,N_44707);
xor U49690 (N_49690,N_44894,N_41318);
xor U49691 (N_49691,N_40158,N_41795);
xor U49692 (N_49692,N_43736,N_42693);
or U49693 (N_49693,N_44336,N_44548);
or U49694 (N_49694,N_43320,N_43490);
or U49695 (N_49695,N_42687,N_43199);
xnor U49696 (N_49696,N_43757,N_42102);
xnor U49697 (N_49697,N_41736,N_40138);
nor U49698 (N_49698,N_40381,N_40094);
nor U49699 (N_49699,N_41319,N_43672);
xnor U49700 (N_49700,N_44982,N_41191);
and U49701 (N_49701,N_43256,N_44635);
xor U49702 (N_49702,N_41576,N_42201);
nand U49703 (N_49703,N_43677,N_44876);
and U49704 (N_49704,N_41247,N_41808);
or U49705 (N_49705,N_44074,N_44001);
xor U49706 (N_49706,N_43120,N_42182);
or U49707 (N_49707,N_41590,N_44633);
xnor U49708 (N_49708,N_41864,N_42663);
xor U49709 (N_49709,N_41481,N_44455);
xnor U49710 (N_49710,N_40495,N_40058);
and U49711 (N_49711,N_44787,N_41451);
xor U49712 (N_49712,N_41320,N_42779);
xor U49713 (N_49713,N_40336,N_43581);
nand U49714 (N_49714,N_42969,N_44151);
and U49715 (N_49715,N_42089,N_43365);
nor U49716 (N_49716,N_43938,N_41259);
nor U49717 (N_49717,N_43880,N_41730);
xor U49718 (N_49718,N_43592,N_44389);
or U49719 (N_49719,N_42299,N_41821);
nand U49720 (N_49720,N_42917,N_44003);
xnor U49721 (N_49721,N_41352,N_40603);
nand U49722 (N_49722,N_43561,N_43299);
or U49723 (N_49723,N_44954,N_40473);
or U49724 (N_49724,N_42924,N_43488);
nor U49725 (N_49725,N_40060,N_42813);
xnor U49726 (N_49726,N_41378,N_41465);
nor U49727 (N_49727,N_42637,N_42532);
and U49728 (N_49728,N_42728,N_40566);
xnor U49729 (N_49729,N_44126,N_44444);
xnor U49730 (N_49730,N_42569,N_40348);
xnor U49731 (N_49731,N_43441,N_43613);
or U49732 (N_49732,N_40424,N_43882);
nor U49733 (N_49733,N_42230,N_44507);
xnor U49734 (N_49734,N_41940,N_44121);
nor U49735 (N_49735,N_40807,N_40427);
nor U49736 (N_49736,N_40082,N_41200);
nor U49737 (N_49737,N_41799,N_43033);
or U49738 (N_49738,N_44241,N_41130);
xor U49739 (N_49739,N_41523,N_43906);
xnor U49740 (N_49740,N_43586,N_43407);
nor U49741 (N_49741,N_40099,N_44848);
xnor U49742 (N_49742,N_43228,N_41017);
xor U49743 (N_49743,N_42241,N_44331);
nor U49744 (N_49744,N_40685,N_40759);
or U49745 (N_49745,N_41404,N_42331);
xor U49746 (N_49746,N_42448,N_42847);
or U49747 (N_49747,N_40774,N_43922);
and U49748 (N_49748,N_40347,N_43763);
or U49749 (N_49749,N_43412,N_42659);
nand U49750 (N_49750,N_43977,N_41524);
nor U49751 (N_49751,N_43403,N_42456);
or U49752 (N_49752,N_41443,N_43064);
nor U49753 (N_49753,N_42262,N_42337);
xor U49754 (N_49754,N_42808,N_43342);
and U49755 (N_49755,N_42131,N_44134);
and U49756 (N_49756,N_44523,N_44436);
nor U49757 (N_49757,N_43179,N_42245);
nand U49758 (N_49758,N_41674,N_42989);
or U49759 (N_49759,N_44003,N_44897);
and U49760 (N_49760,N_40539,N_42052);
or U49761 (N_49761,N_40145,N_43030);
and U49762 (N_49762,N_42323,N_42422);
nor U49763 (N_49763,N_40268,N_40210);
xnor U49764 (N_49764,N_41458,N_43241);
and U49765 (N_49765,N_40970,N_41193);
or U49766 (N_49766,N_42303,N_44044);
nand U49767 (N_49767,N_43661,N_44855);
nand U49768 (N_49768,N_40245,N_41361);
nand U49769 (N_49769,N_44171,N_41402);
nand U49770 (N_49770,N_43369,N_40287);
nand U49771 (N_49771,N_43215,N_44717);
nand U49772 (N_49772,N_43510,N_43014);
nand U49773 (N_49773,N_42976,N_41699);
nor U49774 (N_49774,N_42374,N_44861);
nand U49775 (N_49775,N_44747,N_40180);
xnor U49776 (N_49776,N_44746,N_42060);
and U49777 (N_49777,N_41602,N_43389);
nand U49778 (N_49778,N_44888,N_43147);
nand U49779 (N_49779,N_42658,N_43237);
or U49780 (N_49780,N_40088,N_40738);
or U49781 (N_49781,N_41134,N_43582);
or U49782 (N_49782,N_44792,N_40792);
xor U49783 (N_49783,N_41904,N_41557);
nand U49784 (N_49784,N_43680,N_41981);
and U49785 (N_49785,N_43276,N_44422);
or U49786 (N_49786,N_42950,N_43424);
nand U49787 (N_49787,N_42652,N_44625);
nor U49788 (N_49788,N_41405,N_40683);
or U49789 (N_49789,N_43489,N_42111);
or U49790 (N_49790,N_44112,N_42037);
xnor U49791 (N_49791,N_42726,N_40500);
nor U49792 (N_49792,N_41740,N_43927);
nor U49793 (N_49793,N_40792,N_44120);
nand U49794 (N_49794,N_41923,N_43156);
xor U49795 (N_49795,N_42515,N_40387);
nand U49796 (N_49796,N_44125,N_43265);
and U49797 (N_49797,N_41386,N_44594);
nand U49798 (N_49798,N_42745,N_42628);
and U49799 (N_49799,N_44844,N_44051);
nand U49800 (N_49800,N_43532,N_40434);
or U49801 (N_49801,N_44568,N_44613);
xnor U49802 (N_49802,N_42990,N_42218);
nor U49803 (N_49803,N_40495,N_42939);
nand U49804 (N_49804,N_42447,N_44810);
xor U49805 (N_49805,N_42951,N_41064);
xor U49806 (N_49806,N_44704,N_44787);
nand U49807 (N_49807,N_42802,N_40953);
and U49808 (N_49808,N_44312,N_42122);
or U49809 (N_49809,N_44705,N_41993);
nand U49810 (N_49810,N_40626,N_41790);
or U49811 (N_49811,N_43646,N_42032);
or U49812 (N_49812,N_40784,N_44804);
and U49813 (N_49813,N_43432,N_41013);
and U49814 (N_49814,N_42667,N_44641);
and U49815 (N_49815,N_43160,N_41708);
nand U49816 (N_49816,N_43995,N_42196);
nand U49817 (N_49817,N_41137,N_40873);
xnor U49818 (N_49818,N_43861,N_44935);
or U49819 (N_49819,N_44761,N_40092);
nor U49820 (N_49820,N_40175,N_42831);
nor U49821 (N_49821,N_44412,N_43106);
nand U49822 (N_49822,N_43958,N_40269);
nand U49823 (N_49823,N_43293,N_42814);
or U49824 (N_49824,N_41948,N_40550);
nor U49825 (N_49825,N_44812,N_44292);
nor U49826 (N_49826,N_42092,N_43241);
or U49827 (N_49827,N_43624,N_44029);
and U49828 (N_49828,N_43410,N_40544);
nand U49829 (N_49829,N_40546,N_41574);
xor U49830 (N_49830,N_42996,N_44932);
and U49831 (N_49831,N_42893,N_40678);
or U49832 (N_49832,N_42062,N_40150);
nand U49833 (N_49833,N_44184,N_42026);
nand U49834 (N_49834,N_44718,N_43775);
xnor U49835 (N_49835,N_42784,N_41352);
nor U49836 (N_49836,N_44917,N_41910);
or U49837 (N_49837,N_40967,N_41191);
or U49838 (N_49838,N_40972,N_44582);
nor U49839 (N_49839,N_40769,N_44039);
nor U49840 (N_49840,N_43107,N_42414);
xor U49841 (N_49841,N_40840,N_42631);
or U49842 (N_49842,N_43370,N_43415);
nand U49843 (N_49843,N_40654,N_42111);
xnor U49844 (N_49844,N_41341,N_43227);
or U49845 (N_49845,N_42210,N_42433);
and U49846 (N_49846,N_41663,N_44626);
or U49847 (N_49847,N_43996,N_40092);
and U49848 (N_49848,N_40756,N_40042);
and U49849 (N_49849,N_43214,N_44122);
or U49850 (N_49850,N_42070,N_43201);
nor U49851 (N_49851,N_41260,N_42237);
and U49852 (N_49852,N_42137,N_41146);
xor U49853 (N_49853,N_43760,N_40551);
xor U49854 (N_49854,N_41180,N_43630);
xor U49855 (N_49855,N_41363,N_42464);
nand U49856 (N_49856,N_44658,N_40178);
and U49857 (N_49857,N_41072,N_41493);
nor U49858 (N_49858,N_41646,N_43421);
or U49859 (N_49859,N_43297,N_40712);
xor U49860 (N_49860,N_41438,N_44819);
xor U49861 (N_49861,N_43654,N_44833);
nand U49862 (N_49862,N_43779,N_41740);
or U49863 (N_49863,N_42450,N_42366);
nor U49864 (N_49864,N_44978,N_43435);
and U49865 (N_49865,N_41829,N_44787);
xor U49866 (N_49866,N_43179,N_42253);
nor U49867 (N_49867,N_42835,N_41512);
xnor U49868 (N_49868,N_41372,N_43713);
or U49869 (N_49869,N_40256,N_43292);
nand U49870 (N_49870,N_44710,N_41177);
nor U49871 (N_49871,N_41564,N_44166);
and U49872 (N_49872,N_43646,N_42468);
or U49873 (N_49873,N_42767,N_43632);
nor U49874 (N_49874,N_44814,N_41872);
nand U49875 (N_49875,N_41446,N_44863);
nor U49876 (N_49876,N_41213,N_42573);
nand U49877 (N_49877,N_40201,N_40435);
xnor U49878 (N_49878,N_42540,N_40714);
and U49879 (N_49879,N_44489,N_40198);
nand U49880 (N_49880,N_43680,N_44125);
nor U49881 (N_49881,N_40404,N_44697);
and U49882 (N_49882,N_40187,N_41756);
nor U49883 (N_49883,N_40617,N_41729);
xnor U49884 (N_49884,N_43566,N_43641);
or U49885 (N_49885,N_40147,N_43740);
nor U49886 (N_49886,N_40850,N_41912);
nor U49887 (N_49887,N_42483,N_41177);
nor U49888 (N_49888,N_43689,N_42551);
nor U49889 (N_49889,N_41965,N_43014);
and U49890 (N_49890,N_41336,N_40986);
xor U49891 (N_49891,N_43333,N_40356);
and U49892 (N_49892,N_43426,N_41131);
xnor U49893 (N_49893,N_40380,N_41493);
xor U49894 (N_49894,N_42019,N_40463);
nor U49895 (N_49895,N_40338,N_41817);
and U49896 (N_49896,N_41678,N_42104);
and U49897 (N_49897,N_40737,N_43796);
and U49898 (N_49898,N_42786,N_42990);
xnor U49899 (N_49899,N_44618,N_42588);
xnor U49900 (N_49900,N_43894,N_44592);
xnor U49901 (N_49901,N_44366,N_44828);
nand U49902 (N_49902,N_41516,N_44222);
nor U49903 (N_49903,N_41768,N_41055);
and U49904 (N_49904,N_43865,N_40754);
xor U49905 (N_49905,N_43896,N_43443);
nand U49906 (N_49906,N_43657,N_40324);
and U49907 (N_49907,N_44611,N_44896);
and U49908 (N_49908,N_43930,N_41534);
xor U49909 (N_49909,N_40652,N_43736);
or U49910 (N_49910,N_41641,N_43492);
and U49911 (N_49911,N_43848,N_41967);
or U49912 (N_49912,N_40229,N_42594);
xnor U49913 (N_49913,N_41164,N_40502);
xor U49914 (N_49914,N_44834,N_44846);
nor U49915 (N_49915,N_43416,N_42195);
or U49916 (N_49916,N_40947,N_42670);
xnor U49917 (N_49917,N_41679,N_42453);
nor U49918 (N_49918,N_43461,N_44406);
or U49919 (N_49919,N_43872,N_42765);
nand U49920 (N_49920,N_40841,N_44790);
nand U49921 (N_49921,N_42344,N_42784);
or U49922 (N_49922,N_43730,N_44890);
or U49923 (N_49923,N_41174,N_43134);
xnor U49924 (N_49924,N_41077,N_40786);
and U49925 (N_49925,N_43413,N_41693);
nand U49926 (N_49926,N_44532,N_41645);
or U49927 (N_49927,N_42083,N_40573);
nor U49928 (N_49928,N_44479,N_42662);
and U49929 (N_49929,N_42109,N_43397);
nor U49930 (N_49930,N_43530,N_43995);
xnor U49931 (N_49931,N_42939,N_41300);
nor U49932 (N_49932,N_41770,N_44342);
nand U49933 (N_49933,N_44098,N_42843);
or U49934 (N_49934,N_41301,N_41298);
nor U49935 (N_49935,N_41946,N_43860);
nor U49936 (N_49936,N_41192,N_40053);
or U49937 (N_49937,N_44579,N_42881);
or U49938 (N_49938,N_43059,N_44661);
nand U49939 (N_49939,N_41487,N_43849);
and U49940 (N_49940,N_40419,N_43390);
or U49941 (N_49941,N_41199,N_40481);
and U49942 (N_49942,N_41406,N_44324);
xor U49943 (N_49943,N_40551,N_40264);
and U49944 (N_49944,N_41195,N_44671);
nand U49945 (N_49945,N_40601,N_44494);
xor U49946 (N_49946,N_44181,N_42526);
nor U49947 (N_49947,N_40001,N_42276);
or U49948 (N_49948,N_44417,N_42216);
nand U49949 (N_49949,N_40506,N_41066);
or U49950 (N_49950,N_41846,N_44110);
and U49951 (N_49951,N_41614,N_41442);
nand U49952 (N_49952,N_41547,N_40284);
nor U49953 (N_49953,N_40775,N_42075);
or U49954 (N_49954,N_40158,N_43111);
nor U49955 (N_49955,N_43075,N_43325);
and U49956 (N_49956,N_44630,N_43711);
nand U49957 (N_49957,N_44539,N_41611);
nor U49958 (N_49958,N_43975,N_40341);
and U49959 (N_49959,N_43082,N_40111);
xnor U49960 (N_49960,N_44940,N_43364);
or U49961 (N_49961,N_43489,N_43371);
nor U49962 (N_49962,N_43173,N_40065);
xor U49963 (N_49963,N_40127,N_43737);
nand U49964 (N_49964,N_41338,N_41996);
and U49965 (N_49965,N_43297,N_44963);
nor U49966 (N_49966,N_40091,N_43924);
nand U49967 (N_49967,N_40369,N_43036);
xor U49968 (N_49968,N_40211,N_40306);
or U49969 (N_49969,N_43004,N_43143);
and U49970 (N_49970,N_42897,N_40725);
nor U49971 (N_49971,N_42868,N_44761);
xor U49972 (N_49972,N_42902,N_41630);
xor U49973 (N_49973,N_43569,N_43910);
and U49974 (N_49974,N_41827,N_40243);
or U49975 (N_49975,N_41912,N_43519);
xor U49976 (N_49976,N_41135,N_41065);
nand U49977 (N_49977,N_40386,N_42142);
and U49978 (N_49978,N_43631,N_40783);
nor U49979 (N_49979,N_40026,N_40803);
and U49980 (N_49980,N_43216,N_41006);
nor U49981 (N_49981,N_43387,N_42921);
xnor U49982 (N_49982,N_43014,N_40773);
xnor U49983 (N_49983,N_41495,N_44215);
and U49984 (N_49984,N_43545,N_44921);
nand U49985 (N_49985,N_42773,N_41483);
nand U49986 (N_49986,N_44068,N_43465);
or U49987 (N_49987,N_43120,N_41643);
xor U49988 (N_49988,N_43836,N_44326);
nor U49989 (N_49989,N_44703,N_42322);
nor U49990 (N_49990,N_40530,N_43889);
and U49991 (N_49991,N_43592,N_42879);
nand U49992 (N_49992,N_40924,N_44373);
nand U49993 (N_49993,N_40971,N_41436);
nor U49994 (N_49994,N_43813,N_40416);
and U49995 (N_49995,N_42562,N_43531);
nand U49996 (N_49996,N_41570,N_42896);
xnor U49997 (N_49997,N_43078,N_41054);
nor U49998 (N_49998,N_44686,N_40531);
nand U49999 (N_49999,N_41886,N_41602);
nor UO_0 (O_0,N_45324,N_49415);
xnor UO_1 (O_1,N_45836,N_49822);
or UO_2 (O_2,N_46921,N_48165);
nor UO_3 (O_3,N_45080,N_47679);
nor UO_4 (O_4,N_49425,N_45464);
nor UO_5 (O_5,N_46635,N_46844);
nor UO_6 (O_6,N_47092,N_46122);
or UO_7 (O_7,N_48066,N_46015);
xor UO_8 (O_8,N_47993,N_47295);
and UO_9 (O_9,N_45921,N_46202);
nor UO_10 (O_10,N_48446,N_49774);
and UO_11 (O_11,N_46566,N_46454);
xor UO_12 (O_12,N_47763,N_46753);
or UO_13 (O_13,N_46175,N_46574);
nor UO_14 (O_14,N_49768,N_49860);
xor UO_15 (O_15,N_45598,N_47545);
xor UO_16 (O_16,N_46857,N_48440);
xor UO_17 (O_17,N_45752,N_47903);
or UO_18 (O_18,N_48501,N_49913);
nand UO_19 (O_19,N_45911,N_45115);
xor UO_20 (O_20,N_48202,N_47417);
or UO_21 (O_21,N_46422,N_47929);
and UO_22 (O_22,N_45570,N_46694);
nor UO_23 (O_23,N_49057,N_48568);
or UO_24 (O_24,N_45391,N_46971);
or UO_25 (O_25,N_48227,N_47100);
and UO_26 (O_26,N_48330,N_47951);
nor UO_27 (O_27,N_46813,N_45443);
nand UO_28 (O_28,N_49445,N_45771);
nand UO_29 (O_29,N_46907,N_45841);
xnor UO_30 (O_30,N_49460,N_47387);
xor UO_31 (O_31,N_46763,N_49322);
xor UO_32 (O_32,N_46960,N_49631);
nand UO_33 (O_33,N_46332,N_49030);
and UO_34 (O_34,N_45957,N_48619);
nand UO_35 (O_35,N_46353,N_49624);
and UO_36 (O_36,N_45631,N_47234);
and UO_37 (O_37,N_46046,N_46897);
or UO_38 (O_38,N_45090,N_48098);
or UO_39 (O_39,N_46182,N_49907);
and UO_40 (O_40,N_48693,N_47254);
nor UO_41 (O_41,N_47850,N_46708);
or UO_42 (O_42,N_46311,N_47406);
nand UO_43 (O_43,N_49305,N_48081);
or UO_44 (O_44,N_49837,N_49280);
and UO_45 (O_45,N_46679,N_47625);
or UO_46 (O_46,N_48731,N_47331);
nor UO_47 (O_47,N_46052,N_48069);
xor UO_48 (O_48,N_48076,N_49095);
or UO_49 (O_49,N_49335,N_49553);
nand UO_50 (O_50,N_46469,N_45747);
nor UO_51 (O_51,N_49005,N_47674);
nand UO_52 (O_52,N_49015,N_48567);
and UO_53 (O_53,N_45769,N_48423);
nand UO_54 (O_54,N_48083,N_45894);
nor UO_55 (O_55,N_45927,N_48875);
nor UO_56 (O_56,N_46888,N_48054);
xor UO_57 (O_57,N_49481,N_48253);
nor UO_58 (O_58,N_45823,N_45509);
xor UO_59 (O_59,N_45202,N_49465);
nor UO_60 (O_60,N_46992,N_46630);
nand UO_61 (O_61,N_45863,N_48488);
or UO_62 (O_62,N_47968,N_48761);
or UO_63 (O_63,N_47544,N_48649);
nor UO_64 (O_64,N_45756,N_49055);
xor UO_65 (O_65,N_45359,N_48286);
nor UO_66 (O_66,N_49854,N_48965);
xor UO_67 (O_67,N_48267,N_45337);
nor UO_68 (O_68,N_45540,N_46425);
and UO_69 (O_69,N_45037,N_49618);
or UO_70 (O_70,N_46489,N_49378);
nand UO_71 (O_71,N_49056,N_49111);
nand UO_72 (O_72,N_49935,N_49524);
nand UO_73 (O_73,N_46395,N_48362);
xnor UO_74 (O_74,N_49975,N_45260);
nand UO_75 (O_75,N_48166,N_48425);
or UO_76 (O_76,N_46245,N_46538);
nor UO_77 (O_77,N_49488,N_45355);
nor UO_78 (O_78,N_47312,N_47120);
xnor UO_79 (O_79,N_46858,N_45958);
or UO_80 (O_80,N_45347,N_45288);
xnor UO_81 (O_81,N_46016,N_45567);
and UO_82 (O_82,N_48201,N_45263);
nor UO_83 (O_83,N_49579,N_48867);
or UO_84 (O_84,N_49973,N_45620);
xnor UO_85 (O_85,N_48670,N_49274);
xor UO_86 (O_86,N_47680,N_49841);
or UO_87 (O_87,N_46322,N_49316);
nand UO_88 (O_88,N_46393,N_48575);
nand UO_89 (O_89,N_49431,N_45238);
nor UO_90 (O_90,N_45107,N_48845);
xor UO_91 (O_91,N_48515,N_49674);
nor UO_92 (O_92,N_46204,N_47858);
xor UO_93 (O_93,N_49344,N_47525);
or UO_94 (O_94,N_45221,N_46411);
nor UO_95 (O_95,N_48245,N_47608);
xor UO_96 (O_96,N_47069,N_47512);
nor UO_97 (O_97,N_46354,N_46624);
and UO_98 (O_98,N_46100,N_46220);
xor UO_99 (O_99,N_47440,N_47986);
nor UO_100 (O_100,N_45924,N_45502);
or UO_101 (O_101,N_48973,N_45280);
nor UO_102 (O_102,N_45462,N_45690);
xnor UO_103 (O_103,N_47268,N_46303);
nand UO_104 (O_104,N_48605,N_45009);
xor UO_105 (O_105,N_47155,N_49952);
or UO_106 (O_106,N_45973,N_47463);
nor UO_107 (O_107,N_47731,N_49520);
nor UO_108 (O_108,N_46985,N_45835);
nor UO_109 (O_109,N_46307,N_46607);
and UO_110 (O_110,N_49257,N_49147);
nand UO_111 (O_111,N_49085,N_48294);
or UO_112 (O_112,N_48555,N_49389);
nand UO_113 (O_113,N_45132,N_49444);
or UO_114 (O_114,N_47513,N_46484);
xor UO_115 (O_115,N_47304,N_45493);
nor UO_116 (O_116,N_47727,N_49546);
xor UO_117 (O_117,N_45310,N_47124);
or UO_118 (O_118,N_48114,N_49468);
xor UO_119 (O_119,N_47506,N_46537);
xor UO_120 (O_120,N_46089,N_45980);
nor UO_121 (O_121,N_48410,N_49241);
nor UO_122 (O_122,N_49486,N_47292);
nand UO_123 (O_123,N_49547,N_48496);
and UO_124 (O_124,N_49614,N_48802);
or UO_125 (O_125,N_45802,N_49719);
or UO_126 (O_126,N_45413,N_49130);
or UO_127 (O_127,N_46587,N_46686);
nand UO_128 (O_128,N_48773,N_45209);
nor UO_129 (O_129,N_49778,N_47985);
xor UO_130 (O_130,N_45365,N_45194);
or UO_131 (O_131,N_46993,N_46691);
xnor UO_132 (O_132,N_46285,N_49454);
nor UO_133 (O_133,N_48301,N_45759);
and UO_134 (O_134,N_49590,N_48408);
and UO_135 (O_135,N_46170,N_48335);
nand UO_136 (O_136,N_48836,N_45576);
or UO_137 (O_137,N_48207,N_47219);
and UO_138 (O_138,N_46671,N_47413);
nand UO_139 (O_139,N_45767,N_49027);
nor UO_140 (O_140,N_49140,N_48134);
nor UO_141 (O_141,N_49009,N_49041);
nor UO_142 (O_142,N_49320,N_49174);
or UO_143 (O_143,N_49953,N_48017);
or UO_144 (O_144,N_46756,N_45719);
or UO_145 (O_145,N_45297,N_48378);
nor UO_146 (O_146,N_45490,N_47770);
xor UO_147 (O_147,N_46040,N_49687);
and UO_148 (O_148,N_48130,N_47690);
nor UO_149 (O_149,N_47764,N_46480);
nor UO_150 (O_150,N_45314,N_46515);
and UO_151 (O_151,N_49072,N_46849);
nor UO_152 (O_152,N_47759,N_49155);
and UO_153 (O_153,N_45106,N_48784);
nor UO_154 (O_154,N_45092,N_48862);
or UO_155 (O_155,N_48517,N_48769);
nor UO_156 (O_156,N_45820,N_49177);
nor UO_157 (O_157,N_48226,N_45643);
nand UO_158 (O_158,N_45232,N_48082);
nand UO_159 (O_159,N_48152,N_45308);
nand UO_160 (O_160,N_48285,N_46104);
nand UO_161 (O_161,N_45936,N_49722);
or UO_162 (O_162,N_49353,N_45472);
or UO_163 (O_163,N_48053,N_45654);
or UO_164 (O_164,N_48529,N_45442);
xor UO_165 (O_165,N_47215,N_45910);
xnor UO_166 (O_166,N_49090,N_48158);
or UO_167 (O_167,N_48609,N_49228);
nand UO_168 (O_168,N_46304,N_47734);
and UO_169 (O_169,N_46194,N_47840);
xor UO_170 (O_170,N_45996,N_48903);
nand UO_171 (O_171,N_46447,N_48722);
or UO_172 (O_172,N_49340,N_45041);
nor UO_173 (O_173,N_46051,N_49648);
nand UO_174 (O_174,N_49971,N_48937);
or UO_175 (O_175,N_48975,N_46569);
nor UO_176 (O_176,N_47263,N_45926);
and UO_177 (O_177,N_45094,N_46531);
xnor UO_178 (O_178,N_47516,N_48712);
xor UO_179 (O_179,N_47281,N_48727);
xor UO_180 (O_180,N_47979,N_48871);
and UO_181 (O_181,N_47361,N_45792);
xnor UO_182 (O_182,N_47706,N_49067);
or UO_183 (O_183,N_46092,N_47347);
xor UO_184 (O_184,N_45519,N_47306);
xnor UO_185 (O_185,N_48848,N_48508);
and UO_186 (O_186,N_48827,N_46096);
and UO_187 (O_187,N_46155,N_47446);
xor UO_188 (O_188,N_48264,N_46798);
nor UO_189 (O_189,N_46127,N_48509);
or UO_190 (O_190,N_47602,N_48442);
nor UO_191 (O_191,N_46115,N_46449);
nor UO_192 (O_192,N_47476,N_49360);
or UO_193 (O_193,N_46341,N_46939);
nor UO_194 (O_194,N_46989,N_46709);
or UO_195 (O_195,N_46168,N_46419);
or UO_196 (O_196,N_48469,N_45249);
and UO_197 (O_197,N_49826,N_45180);
and UO_198 (O_198,N_45409,N_45815);
or UO_199 (O_199,N_47536,N_49512);
or UO_200 (O_200,N_48393,N_46034);
nor UO_201 (O_201,N_47345,N_46945);
and UO_202 (O_202,N_46282,N_45342);
nand UO_203 (O_203,N_47225,N_46214);
nand UO_204 (O_204,N_45923,N_49104);
nand UO_205 (O_205,N_46103,N_47125);
xor UO_206 (O_206,N_48334,N_46606);
xnor UO_207 (O_207,N_48870,N_47644);
nor UO_208 (O_208,N_46442,N_47707);
nand UO_209 (O_209,N_49933,N_47747);
or UO_210 (O_210,N_46900,N_48902);
nand UO_211 (O_211,N_48878,N_49004);
nand UO_212 (O_212,N_48172,N_48774);
nor UO_213 (O_213,N_49705,N_45783);
and UO_214 (O_214,N_48224,N_45289);
nor UO_215 (O_215,N_46905,N_47947);
nand UO_216 (O_216,N_47118,N_45373);
and UO_217 (O_217,N_49802,N_47401);
xor UO_218 (O_218,N_48220,N_47587);
and UO_219 (O_219,N_45991,N_45352);
or UO_220 (O_220,N_45328,N_48794);
or UO_221 (O_221,N_49788,N_46856);
and UO_222 (O_222,N_45914,N_47480);
nor UO_223 (O_223,N_48324,N_49379);
nand UO_224 (O_224,N_45676,N_49108);
or UO_225 (O_225,N_48918,N_45210);
or UO_226 (O_226,N_49441,N_45015);
nand UO_227 (O_227,N_47246,N_48126);
or UO_228 (O_228,N_46505,N_47514);
nor UO_229 (O_229,N_46121,N_46359);
and UO_230 (O_230,N_45864,N_47403);
xnor UO_231 (O_231,N_48279,N_49134);
nand UO_232 (O_232,N_48636,N_47896);
nand UO_233 (O_233,N_46731,N_45515);
xor UO_234 (O_234,N_46189,N_47481);
and UO_235 (O_235,N_45514,N_48491);
and UO_236 (O_236,N_47081,N_49219);
nor UO_237 (O_237,N_48830,N_47064);
nor UO_238 (O_238,N_46741,N_49660);
and UO_239 (O_239,N_48854,N_46584);
and UO_240 (O_240,N_49864,N_49411);
and UO_241 (O_241,N_47005,N_48588);
xnor UO_242 (O_242,N_47455,N_47059);
and UO_243 (O_243,N_49079,N_48963);
xnor UO_244 (O_244,N_46809,N_47132);
and UO_245 (O_245,N_49226,N_45197);
xnor UO_246 (O_246,N_46118,N_49630);
or UO_247 (O_247,N_49821,N_45689);
xnor UO_248 (O_248,N_46807,N_48898);
nor UO_249 (O_249,N_46621,N_47523);
or UO_250 (O_250,N_49021,N_46722);
xor UO_251 (O_251,N_49075,N_47335);
and UO_252 (O_252,N_45852,N_48771);
nor UO_253 (O_253,N_46748,N_45492);
xor UO_254 (O_254,N_47569,N_46716);
and UO_255 (O_255,N_49791,N_46467);
or UO_256 (O_256,N_46106,N_48556);
and UO_257 (O_257,N_47846,N_49715);
and UO_258 (O_258,N_49049,N_49811);
xnor UO_259 (O_259,N_46612,N_45089);
xnor UO_260 (O_260,N_47957,N_46755);
or UO_261 (O_261,N_49750,N_49242);
or UO_262 (O_262,N_46056,N_47546);
and UO_263 (O_263,N_47910,N_48648);
nor UO_264 (O_264,N_48317,N_49695);
xor UO_265 (O_265,N_45295,N_48930);
and UO_266 (O_266,N_46319,N_49263);
or UO_267 (O_267,N_49961,N_49686);
or UO_268 (O_268,N_46654,N_49000);
and UO_269 (O_269,N_45206,N_45834);
xnor UO_270 (O_270,N_45292,N_47251);
nand UO_271 (O_271,N_45044,N_48710);
and UO_272 (O_272,N_45954,N_46850);
or UO_273 (O_273,N_48586,N_45406);
or UO_274 (O_274,N_46384,N_46776);
and UO_275 (O_275,N_49679,N_47623);
nand UO_276 (O_276,N_48068,N_48630);
or UO_277 (O_277,N_47435,N_49724);
or UO_278 (O_278,N_45388,N_48949);
or UO_279 (O_279,N_48415,N_45657);
nand UO_280 (O_280,N_45507,N_46737);
nor UO_281 (O_281,N_47857,N_48543);
or UO_282 (O_282,N_45410,N_47889);
nor UO_283 (O_283,N_49135,N_49849);
and UO_284 (O_284,N_47216,N_46605);
xnor UO_285 (O_285,N_48355,N_48671);
and UO_286 (O_286,N_46541,N_45611);
xor UO_287 (O_287,N_46441,N_49487);
and UO_288 (O_288,N_45964,N_45738);
nor UO_289 (O_289,N_47811,N_48487);
nand UO_290 (O_290,N_48148,N_48432);
nor UO_291 (O_291,N_48592,N_48721);
xnor UO_292 (O_292,N_48262,N_48709);
nor UO_293 (O_293,N_49118,N_49582);
and UO_294 (O_294,N_47785,N_49985);
and UO_295 (O_295,N_45001,N_46634);
nand UO_296 (O_296,N_49278,N_45587);
nand UO_297 (O_297,N_47818,N_45699);
or UO_298 (O_298,N_45556,N_48178);
nand UO_299 (O_299,N_46998,N_48382);
or UO_300 (O_300,N_46388,N_48541);
or UO_301 (O_301,N_45018,N_46752);
nor UO_302 (O_302,N_49187,N_46301);
nand UO_303 (O_303,N_48177,N_47130);
nor UO_304 (O_304,N_48512,N_47629);
or UO_305 (O_305,N_49102,N_48979);
xor UO_306 (O_306,N_46642,N_49105);
and UO_307 (O_307,N_45561,N_47470);
or UO_308 (O_308,N_47830,N_47599);
nor UO_309 (O_309,N_49205,N_45329);
or UO_310 (O_310,N_46680,N_46561);
nor UO_311 (O_311,N_45484,N_45166);
and UO_312 (O_312,N_46042,N_46678);
and UO_313 (O_313,N_48683,N_49183);
or UO_314 (O_314,N_46487,N_45368);
nor UO_315 (O_315,N_46500,N_48103);
or UO_316 (O_316,N_48577,N_45239);
and UO_317 (O_317,N_47065,N_45825);
xnor UO_318 (O_318,N_49870,N_48628);
or UO_319 (O_319,N_48367,N_45947);
nor UO_320 (O_320,N_47321,N_48010);
xor UO_321 (O_321,N_47126,N_49188);
xor UO_322 (O_322,N_45114,N_45751);
xnor UO_323 (O_323,N_47802,N_48223);
or UO_324 (O_324,N_45878,N_45582);
and UO_325 (O_325,N_47888,N_45224);
and UO_326 (O_326,N_49645,N_48174);
nand UO_327 (O_327,N_47843,N_46269);
and UO_328 (O_328,N_47672,N_47582);
nand UO_329 (O_329,N_48677,N_49681);
and UO_330 (O_330,N_48782,N_45647);
xor UO_331 (O_331,N_45322,N_46747);
and UO_332 (O_332,N_48591,N_49309);
nand UO_333 (O_333,N_46502,N_49659);
nand UO_334 (O_334,N_47253,N_46173);
xor UO_335 (O_335,N_45457,N_48468);
nand UO_336 (O_336,N_48225,N_47277);
and UO_337 (O_337,N_45816,N_47479);
xor UO_338 (O_338,N_48957,N_49561);
nor UO_339 (O_339,N_48841,N_47036);
and UO_340 (O_340,N_48879,N_49293);
nor UO_341 (O_341,N_48531,N_45574);
nand UO_342 (O_342,N_46069,N_47095);
xnor UO_343 (O_343,N_46184,N_48730);
and UO_344 (O_344,N_47160,N_46721);
or UO_345 (O_345,N_46382,N_45215);
and UO_346 (O_346,N_49338,N_48277);
or UO_347 (O_347,N_48208,N_45504);
nand UO_348 (O_348,N_45299,N_45959);
xor UO_349 (O_349,N_46822,N_49048);
xor UO_350 (O_350,N_46576,N_47927);
nand UO_351 (O_351,N_46032,N_45301);
xnor UO_352 (O_352,N_49051,N_49213);
and UO_353 (O_353,N_46358,N_48091);
nand UO_354 (O_354,N_49697,N_47498);
or UO_355 (O_355,N_49404,N_45380);
nand UO_356 (O_356,N_49221,N_47280);
nor UO_357 (O_357,N_49414,N_45165);
xnor UO_358 (O_358,N_49651,N_46275);
nand UO_359 (O_359,N_49717,N_45169);
nor UO_360 (O_360,N_45192,N_47574);
xor UO_361 (O_361,N_47336,N_47920);
nand UO_362 (O_362,N_46315,N_47886);
nand UO_363 (O_363,N_46966,N_45715);
xor UO_364 (O_364,N_48028,N_46810);
xnor UO_365 (O_365,N_48717,N_49457);
or UO_366 (O_366,N_45278,N_48019);
nand UO_367 (O_367,N_48800,N_48711);
xnor UO_368 (O_368,N_46475,N_47839);
and UO_369 (O_369,N_46037,N_49026);
or UO_370 (O_370,N_49838,N_47354);
nor UO_371 (O_371,N_45590,N_46392);
nand UO_372 (O_372,N_48922,N_47318);
xor UO_373 (O_373,N_46224,N_48893);
or UO_374 (O_374,N_48087,N_48074);
nor UO_375 (O_375,N_47040,N_49673);
or UO_376 (O_376,N_49859,N_47757);
or UO_377 (O_377,N_47908,N_46645);
or UO_378 (O_378,N_48198,N_46720);
xnor UO_379 (O_379,N_45849,N_45644);
and UO_380 (O_380,N_47067,N_49356);
xor UO_381 (O_381,N_47398,N_47866);
or UO_382 (O_382,N_46120,N_48624);
and UO_383 (O_383,N_46216,N_48292);
nor UO_384 (O_384,N_49807,N_45437);
or UO_385 (O_385,N_45276,N_45273);
nand UO_386 (O_386,N_46145,N_46899);
and UO_387 (O_387,N_48196,N_47038);
xnor UO_388 (O_388,N_48329,N_45633);
nor UO_389 (O_389,N_45714,N_45813);
xor UO_390 (O_390,N_47449,N_48389);
nand UO_391 (O_391,N_49270,N_47157);
nor UO_392 (O_392,N_47087,N_48558);
nor UO_393 (O_393,N_48889,N_46166);
xor UO_394 (O_394,N_45832,N_48337);
and UO_395 (O_395,N_47877,N_45744);
xnor UO_396 (O_396,N_45396,N_49620);
or UO_397 (O_397,N_49543,N_49412);
or UO_398 (O_398,N_47752,N_46430);
nor UO_399 (O_399,N_45589,N_45100);
or UO_400 (O_400,N_45242,N_45253);
nor UO_401 (O_401,N_46336,N_47510);
or UO_402 (O_402,N_48559,N_46713);
and UO_403 (O_403,N_45571,N_47116);
or UO_404 (O_404,N_45307,N_48016);
and UO_405 (O_405,N_48175,N_49997);
nand UO_406 (O_406,N_48812,N_48544);
xor UO_407 (O_407,N_47250,N_48779);
xnor UO_408 (O_408,N_47664,N_45489);
nand UO_409 (O_409,N_46935,N_46928);
nand UO_410 (O_410,N_45271,N_47796);
nand UO_411 (O_411,N_49189,N_46906);
or UO_412 (O_412,N_47056,N_46948);
and UO_413 (O_413,N_46625,N_48713);
nor UO_414 (O_414,N_47353,N_46550);
and UO_415 (O_415,N_45763,N_49927);
xor UO_416 (O_416,N_48427,N_48056);
xor UO_417 (O_417,N_47878,N_45984);
nand UO_418 (O_418,N_49564,N_46178);
and UO_419 (O_419,N_45471,N_46828);
nor UO_420 (O_420,N_49967,N_46433);
or UO_421 (O_421,N_48617,N_46055);
nor UO_422 (O_422,N_46924,N_45087);
xnor UO_423 (O_423,N_47020,N_45211);
or UO_424 (O_424,N_48113,N_48001);
nand UO_425 (O_425,N_49502,N_46650);
nand UO_426 (O_426,N_46261,N_49801);
nor UO_427 (O_427,N_47887,N_47483);
and UO_428 (O_428,N_48892,N_48039);
nor UO_429 (O_429,N_47333,N_48006);
nor UO_430 (O_430,N_45588,N_49992);
and UO_431 (O_431,N_45098,N_45151);
nand UO_432 (O_432,N_49753,N_48170);
nand UO_433 (O_433,N_48829,N_49554);
nor UO_434 (O_434,N_48537,N_46931);
xor UO_435 (O_435,N_47824,N_48161);
xor UO_436 (O_436,N_46227,N_46564);
and UO_437 (O_437,N_47776,N_48897);
nor UO_438 (O_438,N_45725,N_47176);
xor UO_439 (O_439,N_48365,N_45701);
xnor UO_440 (O_440,N_46647,N_48764);
xor UO_441 (O_441,N_48043,N_45052);
xor UO_442 (O_442,N_49795,N_45045);
nor UO_443 (O_443,N_48877,N_47152);
xnor UO_444 (O_444,N_48536,N_48633);
nand UO_445 (O_445,N_49331,N_49597);
xor UO_446 (O_446,N_48735,N_47496);
nand UO_447 (O_447,N_46872,N_47870);
xnor UO_448 (O_448,N_45040,N_48302);
xor UO_449 (O_449,N_46386,N_49038);
nor UO_450 (O_450,N_49450,N_47196);
and UO_451 (O_451,N_48562,N_47459);
or UO_452 (O_452,N_45174,N_49399);
and UO_453 (O_453,N_48011,N_47505);
or UO_454 (O_454,N_49946,N_49097);
nand UO_455 (O_455,N_49919,N_47825);
and UO_456 (O_456,N_46101,N_48287);
or UO_457 (O_457,N_49248,N_49970);
and UO_458 (O_458,N_48886,N_45754);
xor UO_459 (O_459,N_48195,N_45277);
and UO_460 (O_460,N_47677,N_46710);
nand UO_461 (O_461,N_45503,N_47025);
and UO_462 (O_462,N_48611,N_47844);
or UO_463 (O_463,N_48806,N_47342);
xor UO_464 (O_464,N_49043,N_47831);
nor UO_465 (O_465,N_45522,N_48243);
nand UO_466 (O_466,N_46081,N_46583);
nor UO_467 (O_467,N_45645,N_48590);
xor UO_468 (O_468,N_49965,N_49976);
xor UO_469 (O_469,N_45648,N_49856);
nor UO_470 (O_470,N_49334,N_47454);
and UO_471 (O_471,N_48763,N_45776);
nand UO_472 (O_472,N_49006,N_49556);
or UO_473 (O_473,N_45007,N_46958);
nand UO_474 (O_474,N_48781,N_49466);
and UO_475 (O_475,N_47188,N_45216);
and UO_476 (O_476,N_46950,N_45086);
nor UO_477 (O_477,N_47329,N_45060);
and UO_478 (O_478,N_49814,N_48869);
or UO_479 (O_479,N_47079,N_48796);
and UO_480 (O_480,N_48641,N_49467);
xnor UO_481 (O_481,N_45703,N_48993);
nor UO_482 (O_482,N_46327,N_48691);
nor UO_483 (O_483,N_48116,N_46623);
nand UO_484 (O_484,N_47928,N_45500);
or UO_485 (O_485,N_49577,N_45270);
xnor UO_486 (O_486,N_45061,N_45895);
nor UO_487 (O_487,N_46592,N_48849);
nand UO_488 (O_488,N_48720,N_47341);
or UO_489 (O_489,N_46513,N_48911);
nor UO_490 (O_490,N_45120,N_47583);
xor UO_491 (O_491,N_45780,N_45420);
nor UO_492 (O_492,N_48197,N_45880);
nand UO_493 (O_493,N_45485,N_46862);
nor UO_494 (O_494,N_47217,N_47052);
and UO_495 (O_495,N_49082,N_47085);
and UO_496 (O_496,N_49698,N_49716);
and UO_497 (O_497,N_46575,N_48485);
and UO_498 (O_498,N_48739,N_46961);
nor UO_499 (O_499,N_49958,N_48353);
nand UO_500 (O_500,N_47183,N_45887);
or UO_501 (O_501,N_48992,N_46539);
nand UO_502 (O_502,N_46219,N_47613);
nand UO_503 (O_503,N_48191,N_47099);
nand UO_504 (O_504,N_47600,N_46344);
xor UO_505 (O_505,N_47478,N_48050);
xor UO_506 (O_506,N_45967,N_47499);
and UO_507 (O_507,N_46853,N_46059);
or UO_508 (O_508,N_45951,N_45794);
nor UO_509 (O_509,N_46190,N_47482);
or UO_510 (O_510,N_45234,N_48390);
nand UO_511 (O_511,N_48308,N_45416);
xnor UO_512 (O_512,N_46452,N_45161);
or UO_513 (O_513,N_49763,N_48809);
or UO_514 (O_514,N_45740,N_46668);
nand UO_515 (O_515,N_47101,N_47173);
nor UO_516 (O_516,N_47634,N_49116);
nand UO_517 (O_517,N_49480,N_48885);
or UO_518 (O_518,N_45491,N_47091);
or UO_519 (O_519,N_47795,N_47148);
or UO_520 (O_520,N_49192,N_49195);
nand UO_521 (O_521,N_47592,N_45712);
nand UO_522 (O_522,N_48109,N_48860);
or UO_523 (O_523,N_47465,N_49253);
xnor UO_524 (O_524,N_48151,N_47862);
or UO_525 (O_525,N_48049,N_46617);
nand UO_526 (O_526,N_47698,N_49771);
nor UO_527 (O_527,N_47307,N_47639);
nand UO_528 (O_528,N_45547,N_47635);
and UO_529 (O_529,N_45865,N_48718);
nand UO_530 (O_530,N_45266,N_49685);
xnor UO_531 (O_531,N_47990,N_47998);
xnor UO_532 (O_532,N_46664,N_47232);
xor UO_533 (O_533,N_48579,N_49164);
or UO_534 (O_534,N_48951,N_47464);
xnor UO_535 (O_535,N_48634,N_45077);
and UO_536 (O_536,N_48916,N_47458);
xnor UO_537 (O_537,N_49664,N_47800);
and UO_538 (O_538,N_46990,N_49789);
and UO_539 (O_539,N_47875,N_45117);
or UO_540 (O_540,N_45520,N_46434);
nand UO_541 (O_541,N_49034,N_45709);
nand UO_542 (O_542,N_47520,N_45551);
or UO_543 (O_543,N_48667,N_49417);
and UO_544 (O_544,N_49922,N_47045);
nand UO_545 (O_545,N_46514,N_49428);
or UO_546 (O_546,N_46929,N_46481);
nand UO_547 (O_547,N_49315,N_45111);
nor UO_548 (O_548,N_48563,N_46889);
nand UO_549 (O_549,N_45640,N_45392);
nand UO_550 (O_550,N_45411,N_49084);
nor UO_551 (O_551,N_49497,N_46496);
nand UO_552 (O_552,N_47647,N_46544);
xor UO_553 (O_553,N_48123,N_46495);
nand UO_554 (O_554,N_48850,N_45608);
xnor UO_555 (O_555,N_49052,N_46771);
xnor UO_556 (O_556,N_45772,N_48940);
or UO_557 (O_557,N_48465,N_45839);
nand UO_558 (O_558,N_45178,N_48080);
nor UO_559 (O_559,N_48414,N_46815);
or UO_560 (O_560,N_46373,N_47290);
nand UO_561 (O_561,N_48012,N_47589);
nor UO_562 (O_562,N_48745,N_46946);
xnor UO_563 (O_563,N_48413,N_49224);
or UO_564 (O_564,N_49522,N_46860);
nor UO_565 (O_565,N_46074,N_48982);
nand UO_566 (O_566,N_49616,N_45679);
or UO_567 (O_567,N_49405,N_47323);
nor UO_568 (O_568,N_46455,N_48637);
or UO_569 (O_569,N_45904,N_48246);
and UO_570 (O_570,N_49277,N_48919);
nand UO_571 (O_571,N_49496,N_49167);
nor UO_572 (O_572,N_46868,N_49375);
nor UO_573 (O_573,N_48306,N_45981);
nand UO_574 (O_574,N_47687,N_49963);
xor UO_575 (O_575,N_46526,N_48618);
nand UO_576 (O_576,N_46991,N_48612);
xnor UO_577 (O_577,N_45163,N_45623);
and UO_578 (O_578,N_48770,N_49987);
xor UO_579 (O_579,N_46254,N_45692);
xnor UO_580 (O_580,N_46791,N_49308);
and UO_581 (O_581,N_46767,N_46593);
nand UO_582 (O_582,N_45312,N_47213);
or UO_583 (O_583,N_49898,N_47055);
xor UO_584 (O_584,N_47247,N_48737);
or UO_585 (O_585,N_46260,N_49218);
xnor UO_586 (O_586,N_46372,N_46404);
nor UO_587 (O_587,N_49016,N_46920);
xor UO_588 (O_588,N_48994,N_48658);
xor UO_589 (O_589,N_49710,N_45173);
and UO_590 (O_590,N_47725,N_45554);
xor UO_591 (O_591,N_47882,N_48995);
xor UO_592 (O_592,N_48765,N_49678);
nand UO_593 (O_593,N_46417,N_49602);
xor UO_594 (O_594,N_46504,N_45626);
and UO_595 (O_595,N_46786,N_49670);
and UO_596 (O_596,N_47293,N_48791);
and UO_597 (O_597,N_45466,N_46073);
and UO_598 (O_598,N_46728,N_46762);
xor UO_599 (O_599,N_48342,N_48906);
nand UO_600 (O_600,N_46049,N_49784);
and UO_601 (O_601,N_49121,N_47201);
xnor UO_602 (O_602,N_49730,N_48639);
or UO_603 (O_603,N_45350,N_47129);
and UO_604 (O_604,N_45838,N_45313);
and UO_605 (O_605,N_49667,N_45562);
and UO_606 (O_606,N_48626,N_47616);
or UO_607 (O_607,N_46764,N_46806);
nand UO_608 (O_608,N_46845,N_48278);
and UO_609 (O_609,N_48097,N_49509);
nand UO_610 (O_610,N_48265,N_46488);
nand UO_611 (O_611,N_45482,N_45367);
or UO_612 (O_612,N_46482,N_47489);
or UO_613 (O_613,N_47901,N_45872);
nor UO_614 (O_614,N_47174,N_49540);
and UO_615 (O_615,N_49657,N_49809);
xor UO_616 (O_616,N_45176,N_46761);
and UO_617 (O_617,N_45427,N_48874);
or UO_618 (O_618,N_49066,N_46299);
and UO_619 (O_619,N_49769,N_46067);
xor UO_620 (O_620,N_45377,N_49387);
nand UO_621 (O_621,N_46128,N_49729);
nor UO_622 (O_622,N_49508,N_49294);
nand UO_623 (O_623,N_47026,N_45004);
or UO_624 (O_624,N_48176,N_47428);
nand UO_625 (O_625,N_45050,N_47349);
xnor UO_626 (O_626,N_48462,N_48998);
xor UO_627 (O_627,N_47442,N_45140);
nand UO_628 (O_628,N_48106,N_45137);
xor UO_629 (O_629,N_48140,N_47841);
xor UO_630 (O_630,N_46714,N_49993);
or UO_631 (O_631,N_49877,N_45903);
nand UO_632 (O_632,N_47504,N_49880);
nand UO_633 (O_633,N_48861,N_48218);
or UO_634 (O_634,N_49394,N_47953);
and UO_635 (O_635,N_49060,N_47343);
xor UO_636 (O_636,N_45303,N_48955);
nand UO_637 (O_637,N_48147,N_49605);
or UO_638 (O_638,N_47285,N_48018);
nand UO_639 (O_639,N_45230,N_45375);
nand UO_640 (O_640,N_45937,N_46098);
nor UO_641 (O_641,N_45706,N_47715);
nor UO_642 (O_642,N_45828,N_46926);
nor UO_643 (O_643,N_46019,N_49846);
nand UO_644 (O_644,N_49536,N_46797);
nand UO_645 (O_645,N_48689,N_46665);
xor UO_646 (O_646,N_46555,N_45800);
or UO_647 (O_647,N_45804,N_45203);
xor UO_648 (O_648,N_48171,N_47938);
and UO_649 (O_649,N_47827,N_47089);
and UO_650 (O_650,N_49892,N_49541);
nand UO_651 (O_651,N_45634,N_46632);
nand UO_652 (O_652,N_47788,N_45167);
nand UO_653 (O_653,N_47322,N_48817);
and UO_654 (O_654,N_48552,N_45778);
or UO_655 (O_655,N_45943,N_49077);
nand UO_656 (O_656,N_46943,N_48646);
nor UO_657 (O_657,N_48048,N_49435);
nand UO_658 (O_658,N_47115,N_47683);
nor UO_659 (O_659,N_45177,N_45304);
xor UO_660 (O_660,N_48467,N_45073);
nand UO_661 (O_661,N_45722,N_46622);
or UO_662 (O_662,N_47303,N_46639);
xnor UO_663 (O_663,N_49995,N_49748);
nor UO_664 (O_664,N_45755,N_45387);
nand UO_665 (O_665,N_45993,N_47708);
or UO_666 (O_666,N_47653,N_48969);
nor UO_667 (O_667,N_47328,N_45378);
nor UO_668 (O_668,N_48325,N_49511);
xnor UO_669 (O_669,N_47240,N_48051);
or UO_670 (O_670,N_45011,N_49348);
and UO_671 (O_671,N_45453,N_48275);
xor UO_672 (O_672,N_48348,N_46697);
nor UO_673 (O_673,N_46394,N_47579);
and UO_674 (O_674,N_47809,N_48811);
nand UO_675 (O_675,N_48479,N_47249);
nor UO_676 (O_676,N_49949,N_49575);
nand UO_677 (O_677,N_47904,N_47302);
and UO_678 (O_678,N_46258,N_46277);
xnor UO_679 (O_679,N_47378,N_47169);
and UO_680 (O_680,N_45764,N_47703);
nor UO_681 (O_681,N_49830,N_45907);
or UO_682 (O_682,N_49545,N_47450);
and UO_683 (O_683,N_47379,N_46944);
nand UO_684 (O_684,N_47697,N_47070);
nor UO_685 (O_685,N_48684,N_46540);
and UO_686 (O_686,N_47351,N_49260);
nor UO_687 (O_687,N_46355,N_46843);
nor UO_688 (O_688,N_49054,N_47184);
xor UO_689 (O_689,N_46896,N_47050);
xor UO_690 (O_690,N_49010,N_45225);
nor UO_691 (O_691,N_46804,N_49182);
xor UO_692 (O_692,N_48792,N_45624);
nand UO_693 (O_693,N_45385,N_46369);
nand UO_694 (O_694,N_46543,N_48987);
or UO_695 (O_695,N_45425,N_49947);
nand UO_696 (O_696,N_47190,N_48844);
xor UO_697 (O_697,N_45463,N_49112);
or UO_698 (O_698,N_49327,N_48890);
and UO_699 (O_699,N_45035,N_46877);
or UO_700 (O_700,N_48585,N_49349);
xnor UO_701 (O_701,N_49558,N_49693);
nand UO_702 (O_702,N_47109,N_46754);
or UO_703 (O_703,N_48535,N_48748);
or UO_704 (O_704,N_48888,N_45429);
or UO_705 (O_705,N_46271,N_49843);
and UO_706 (O_706,N_46171,N_45527);
nor UO_707 (O_707,N_49361,N_45049);
nand UO_708 (O_708,N_45495,N_46789);
xor UO_709 (O_709,N_48293,N_48866);
nand UO_710 (O_710,N_49598,N_45293);
or UO_711 (O_711,N_48435,N_46140);
nor UO_712 (O_712,N_47907,N_47559);
nand UO_713 (O_713,N_45379,N_48094);
xor UO_714 (O_714,N_49490,N_45580);
xnor UO_715 (O_715,N_47735,N_46468);
and UO_716 (O_716,N_49580,N_47621);
nand UO_717 (O_717,N_46159,N_48305);
nor UO_718 (O_718,N_47041,N_45698);
or UO_719 (O_719,N_46692,N_47670);
or UO_720 (O_720,N_47076,N_48157);
nand UO_721 (O_721,N_49125,N_46235);
nor UO_722 (O_722,N_46221,N_48984);
or UO_723 (O_723,N_47086,N_46796);
xor UO_724 (O_724,N_46745,N_49096);
nor UO_725 (O_725,N_49471,N_47352);
and UO_726 (O_726,N_46719,N_47944);
and UO_727 (O_727,N_45994,N_46739);
and UO_728 (O_728,N_48359,N_47962);
nand UO_729 (O_729,N_45309,N_46878);
or UO_730 (O_730,N_46983,N_49144);
and UO_731 (O_731,N_48754,N_48117);
or UO_732 (O_732,N_49966,N_48729);
or UO_733 (O_733,N_46342,N_48498);
nand UO_734 (O_734,N_48451,N_45047);
nand UO_735 (O_735,N_46429,N_46876);
nor UO_736 (O_736,N_46859,N_49766);
nor UO_737 (O_737,N_49609,N_45074);
and UO_738 (O_738,N_45327,N_49646);
xor UO_739 (O_739,N_47699,N_47638);
xor UO_740 (O_740,N_48584,N_45432);
nand UO_741 (O_741,N_47595,N_46875);
or UO_742 (O_742,N_47756,N_49560);
and UO_743 (O_743,N_46023,N_49266);
nand UO_744 (O_744,N_47248,N_46399);
nand UO_745 (O_745,N_47395,N_46673);
xor UO_746 (O_746,N_46117,N_45449);
nor UO_747 (O_747,N_48600,N_49593);
or UO_748 (O_748,N_47704,N_48595);
nand UO_749 (O_749,N_46025,N_47917);
nor UO_750 (O_750,N_46278,N_47106);
or UO_751 (O_751,N_45441,N_48694);
xnor UO_752 (O_752,N_45897,N_47650);
nand UO_753 (O_753,N_47586,N_48128);
or UO_754 (O_754,N_48623,N_48412);
xor UO_755 (O_755,N_47799,N_46071);
nor UO_756 (O_756,N_46693,N_49373);
and UO_757 (O_757,N_46781,N_47468);
xnor UO_758 (O_758,N_47049,N_49243);
nand UO_759 (O_759,N_49956,N_49489);
or UO_760 (O_760,N_46450,N_49114);
xnor UO_761 (O_761,N_45122,N_45281);
nor UO_762 (O_762,N_45247,N_47339);
and UO_763 (O_763,N_49374,N_49767);
and UO_764 (O_764,N_48331,N_47705);
and UO_765 (O_765,N_45599,N_48946);
and UO_766 (O_766,N_48826,N_45256);
nand UO_767 (O_767,N_45535,N_49333);
and UO_768 (O_768,N_48503,N_45405);
nor UO_769 (O_769,N_49549,N_46535);
nand UO_770 (O_770,N_45187,N_49915);
xnor UO_771 (O_771,N_46599,N_48474);
xor UO_772 (O_772,N_45474,N_49638);
and UO_773 (O_773,N_46314,N_48996);
xnor UO_774 (O_774,N_48863,N_46840);
and UO_775 (O_775,N_45812,N_49875);
nor UO_776 (O_776,N_47658,N_48349);
or UO_777 (O_777,N_47429,N_47911);
nand UO_778 (O_778,N_46579,N_49855);
nor UO_779 (O_779,N_46396,N_48938);
xnor UO_780 (O_780,N_47867,N_45065);
and UO_781 (O_781,N_48805,N_48120);
or UO_782 (O_782,N_46956,N_46863);
xnor UO_783 (O_783,N_47954,N_46274);
nor UO_784 (O_784,N_47235,N_49706);
nand UO_785 (O_785,N_49262,N_48482);
nand UO_786 (O_786,N_48828,N_45128);
or UO_787 (O_787,N_47367,N_46557);
xnor UO_788 (O_788,N_48760,N_47135);
xor UO_789 (O_789,N_47034,N_45116);
nor UO_790 (O_790,N_49525,N_47641);
nor UO_791 (O_791,N_46952,N_49008);
nor UO_792 (O_792,N_47614,N_46478);
nor UO_793 (O_793,N_47700,N_46811);
and UO_794 (O_794,N_47952,N_47243);
xnor UO_795 (O_795,N_45916,N_48645);
and UO_796 (O_796,N_49410,N_47750);
nor UO_797 (O_797,N_45750,N_45233);
nor UO_798 (O_798,N_48787,N_46018);
or UO_799 (O_799,N_46567,N_46510);
nand UO_800 (O_800,N_48030,N_48603);
nand UO_801 (O_801,N_47414,N_49815);
xnor UO_802 (O_802,N_46398,N_46165);
or UO_803 (O_803,N_49046,N_46244);
nor UO_804 (O_804,N_47880,N_45129);
and UO_805 (O_805,N_48540,N_47684);
or UO_806 (O_806,N_49282,N_46782);
or UO_807 (O_807,N_45516,N_49944);
xnor UO_808 (O_808,N_46066,N_47786);
nor UO_809 (O_809,N_48230,N_49663);
and UO_810 (O_810,N_49865,N_47334);
nor UO_811 (O_811,N_46263,N_47488);
nor UO_812 (O_812,N_45325,N_48352);
nand UO_813 (O_813,N_46832,N_46553);
nor UO_814 (O_814,N_49749,N_46440);
xnor UO_815 (O_815,N_48814,N_45478);
xnor UO_816 (O_816,N_45435,N_48598);
xnor UO_817 (O_817,N_47035,N_48808);
nand UO_818 (O_818,N_47416,N_45583);
xor UO_819 (O_819,N_45008,N_46865);
or UO_820 (O_820,N_45663,N_49025);
and UO_821 (O_821,N_45672,N_48644);
or UO_822 (O_822,N_49606,N_45056);
nand UO_823 (O_823,N_48855,N_45848);
xor UO_824 (O_824,N_49810,N_49505);
nor UO_825 (O_825,N_47231,N_49214);
or UO_826 (O_826,N_45777,N_47711);
nand UO_827 (O_827,N_49451,N_48092);
or UO_828 (O_828,N_46302,N_45982);
and UO_829 (O_829,N_45473,N_47633);
nand UO_830 (O_830,N_47147,N_46111);
or UO_831 (O_831,N_48187,N_46438);
nor UO_832 (O_832,N_49040,N_49146);
xor UO_833 (O_833,N_48941,N_47973);
nor UO_834 (O_834,N_47814,N_45606);
nand UO_835 (O_835,N_46738,N_49197);
or UO_836 (O_836,N_49429,N_47298);
nor UO_837 (O_837,N_46167,N_46914);
nand UO_838 (O_838,N_49957,N_45513);
nor UO_839 (O_839,N_45637,N_48338);
and UO_840 (O_840,N_47409,N_46385);
nor UO_841 (O_841,N_49161,N_48714);
nor UO_842 (O_842,N_49920,N_49318);
or UO_843 (O_843,N_46803,N_48686);
and UO_844 (O_844,N_48179,N_47732);
nand UO_845 (O_845,N_45021,N_48656);
xnor UO_846 (O_846,N_48818,N_49238);
and UO_847 (O_847,N_47837,N_46852);
nand UO_848 (O_848,N_45511,N_49382);
or UO_849 (O_849,N_48723,N_45434);
and UO_850 (O_850,N_47017,N_49840);
and UO_851 (O_851,N_45666,N_45083);
nor UO_852 (O_852,N_48822,N_47948);
or UO_853 (O_853,N_47965,N_46371);
or UO_854 (O_854,N_47792,N_49751);
nand UO_855 (O_855,N_48460,N_46135);
nand UO_856 (O_856,N_49281,N_48627);
or UO_857 (O_857,N_45439,N_48138);
nor UO_858 (O_858,N_46228,N_47469);
nand UO_859 (O_859,N_49493,N_47452);
nor UO_860 (O_860,N_47593,N_47645);
xnor UO_861 (O_861,N_46594,N_45707);
and UO_862 (O_862,N_45510,N_46231);
xnor UO_863 (O_863,N_47782,N_45093);
nand UO_864 (O_864,N_49701,N_47177);
or UO_865 (O_865,N_49064,N_47812);
nand UO_866 (O_866,N_49127,N_47905);
xor UO_867 (O_867,N_48601,N_46125);
nor UO_868 (O_868,N_46188,N_46830);
xor UO_869 (O_869,N_47581,N_47975);
xor UO_870 (O_870,N_46742,N_48502);
xnor UO_871 (O_871,N_49426,N_49252);
nor UO_872 (O_872,N_46637,N_45622);
and UO_873 (O_873,N_45970,N_45625);
xnor UO_874 (O_874,N_48744,N_45909);
nor UO_875 (O_875,N_47879,N_48304);
nand UO_876 (O_876,N_49903,N_49159);
nand UO_877 (O_877,N_45022,N_45265);
nand UO_878 (O_878,N_49080,N_47738);
nor UO_879 (O_879,N_45227,N_46094);
or UO_880 (O_880,N_46597,N_46308);
xnor UO_881 (O_881,N_48813,N_47992);
or UO_882 (O_882,N_46133,N_45869);
nor UO_883 (O_883,N_47466,N_45941);
xnor UO_884 (O_884,N_47185,N_46816);
nor UO_885 (O_885,N_45196,N_48756);
nor UO_886 (O_886,N_48665,N_49813);
and UO_887 (O_887,N_46949,N_45826);
and UO_888 (O_888,N_48783,N_45005);
nand UO_889 (O_889,N_46364,N_46402);
nor UO_890 (O_890,N_46827,N_49708);
or UO_891 (O_891,N_46346,N_47774);
or UO_892 (O_892,N_47537,N_48392);
or UO_893 (O_893,N_49235,N_49700);
or UO_894 (O_894,N_45038,N_45054);
or UO_895 (O_895,N_48801,N_45660);
xnor UO_896 (O_896,N_46033,N_49756);
nor UO_897 (O_897,N_47158,N_46022);
xor UO_898 (O_898,N_45847,N_45871);
or UO_899 (O_899,N_47111,N_47995);
nand UO_900 (O_900,N_47448,N_45433);
or UO_901 (O_901,N_48314,N_49904);
nand UO_902 (O_902,N_49727,N_46884);
or UO_903 (O_903,N_47541,N_47940);
or UO_904 (O_904,N_45319,N_46735);
nor UO_905 (O_905,N_46711,N_47266);
and UO_906 (O_906,N_46972,N_47094);
or UO_907 (O_907,N_45938,N_45066);
and UO_908 (O_908,N_49544,N_49534);
nor UO_909 (O_909,N_48798,N_46788);
xnor UO_910 (O_910,N_49420,N_48929);
or UO_911 (O_911,N_48507,N_46012);
and UO_912 (O_912,N_45099,N_47771);
and UO_913 (O_913,N_48431,N_49977);
nand UO_914 (O_914,N_45724,N_48666);
nand UO_915 (O_915,N_49983,N_45361);
or UO_916 (O_916,N_49306,N_46941);
and UO_917 (O_917,N_45990,N_48316);
xor UO_918 (O_918,N_46836,N_45741);
xor UO_919 (O_919,N_47212,N_48206);
or UO_920 (O_920,N_48883,N_45758);
nand UO_921 (O_921,N_46523,N_49494);
xnor UO_922 (O_922,N_47384,N_49816);
nor UO_923 (O_923,N_46413,N_49419);
nand UO_924 (O_924,N_45033,N_47337);
xnor UO_925 (O_925,N_45333,N_47720);
nand UO_926 (O_926,N_46727,N_48222);
or UO_927 (O_927,N_46787,N_49217);
nand UO_928 (O_928,N_45614,N_49779);
xor UO_929 (O_929,N_45728,N_48323);
and UO_930 (O_930,N_45091,N_49007);
or UO_931 (O_931,N_46802,N_48741);
and UO_932 (O_932,N_45684,N_49828);
xor UO_933 (O_933,N_48759,N_45678);
xnor UO_934 (O_934,N_46982,N_48239);
or UO_935 (O_935,N_46814,N_46082);
and UO_936 (O_936,N_49357,N_49297);
xnor UO_937 (O_937,N_49584,N_47678);
xor UO_938 (O_938,N_47753,N_46582);
xnor UO_939 (O_939,N_49139,N_45850);
and UO_940 (O_940,N_48956,N_47804);
nand UO_941 (O_941,N_47370,N_46078);
nand UO_942 (O_942,N_48027,N_46288);
xor UO_943 (O_943,N_45096,N_47543);
xor UO_944 (O_944,N_47956,N_45986);
and UO_945 (O_945,N_45857,N_47567);
xor UO_946 (O_946,N_49829,N_48311);
and UO_947 (O_947,N_46026,N_48058);
xor UO_948 (O_948,N_46134,N_46116);
and UO_949 (O_949,N_45059,N_48981);
and UO_950 (O_950,N_47913,N_49694);
and UO_951 (O_951,N_48075,N_47503);
and UO_952 (O_952,N_49350,N_45332);
nand UO_953 (O_953,N_46222,N_46192);
or UO_954 (O_954,N_49733,N_49176);
xor UO_955 (O_955,N_48443,N_46525);
and UO_956 (O_956,N_46108,N_48669);
and UO_957 (O_957,N_48966,N_46628);
xor UO_958 (O_958,N_45559,N_45718);
or UO_959 (O_959,N_49106,N_49636);
nand UO_960 (O_960,N_46670,N_46238);
or UO_961 (O_961,N_47988,N_48159);
nand UO_962 (O_962,N_47591,N_47006);
nor UO_963 (O_963,N_47722,N_46004);
nor UO_964 (O_964,N_48602,N_49623);
and UO_965 (O_965,N_46279,N_47320);
or UO_966 (O_966,N_48040,N_47551);
nor UO_967 (O_967,N_48663,N_48958);
and UO_968 (O_968,N_46962,N_47836);
and UO_969 (O_969,N_46784,N_47047);
or UO_970 (O_970,N_48528,N_48690);
xor UO_971 (O_971,N_48788,N_45272);
nand UO_972 (O_972,N_49622,N_46444);
nor UO_973 (O_973,N_48129,N_48868);
and UO_974 (O_974,N_49755,N_45788);
or UO_975 (O_975,N_49137,N_49033);
nand UO_976 (O_976,N_49982,N_47991);
xor UO_977 (O_977,N_47178,N_47806);
or UO_978 (O_978,N_49271,N_48939);
xor UO_979 (O_979,N_45592,N_47755);
xor UO_980 (O_980,N_45568,N_49070);
or UO_981 (O_981,N_49478,N_48751);
nor UO_982 (O_982,N_45153,N_47733);
or UO_983 (O_983,N_47381,N_45193);
nor UO_984 (O_984,N_45635,N_48404);
and UO_985 (O_985,N_45686,N_45757);
nor UO_986 (O_986,N_48386,N_45269);
nor UO_987 (O_987,N_48360,N_49256);
and UO_988 (O_988,N_49787,N_45840);
nor UO_989 (O_989,N_47172,N_48820);
nand UO_990 (O_990,N_45415,N_46769);
or UO_991 (O_991,N_47371,N_45944);
nor UO_992 (O_992,N_46942,N_48882);
xor UO_993 (O_993,N_46295,N_47028);
or UO_994 (O_994,N_48375,N_47456);
nor UO_995 (O_995,N_45252,N_49268);
xnor UO_996 (O_996,N_49453,N_47745);
and UO_997 (O_997,N_47532,N_47575);
nand UO_998 (O_998,N_49390,N_48989);
xnor UO_999 (O_999,N_46881,N_47919);
and UO_1000 (O_1000,N_45960,N_46400);
or UO_1001 (O_1001,N_46297,N_45564);
or UO_1002 (O_1002,N_45824,N_46109);
nand UO_1003 (O_1003,N_47637,N_49874);
and UO_1004 (O_1004,N_46126,N_45182);
nor UO_1005 (O_1005,N_46397,N_45533);
or UO_1006 (O_1006,N_46556,N_49603);
xor UO_1007 (O_1007,N_46778,N_48962);
xnor UO_1008 (O_1008,N_48767,N_49819);
xnor UO_1009 (O_1009,N_49200,N_47787);
xor UO_1010 (O_1010,N_49103,N_49504);
nand UO_1011 (O_1011,N_46223,N_46201);
nor UO_1012 (O_1012,N_46197,N_48102);
and UO_1013 (O_1013,N_47407,N_48185);
or UO_1014 (O_1014,N_47659,N_47003);
and UO_1015 (O_1015,N_48539,N_47224);
or UO_1016 (O_1016,N_49442,N_47749);
or UO_1017 (O_1017,N_46119,N_45112);
nor UO_1018 (O_1018,N_46215,N_46061);
xor UO_1019 (O_1019,N_49567,N_46659);
nand UO_1020 (O_1020,N_49731,N_47218);
and UO_1021 (O_1021,N_48122,N_45217);
xor UO_1022 (O_1022,N_49615,N_47271);
nand UO_1023 (O_1023,N_49637,N_47955);
nand UO_1024 (O_1024,N_47396,N_46977);
xor UO_1025 (O_1025,N_48221,N_48169);
nor UO_1026 (O_1026,N_47618,N_49943);
nor UO_1027 (O_1027,N_48250,N_48499);
or UO_1028 (O_1028,N_49692,N_48212);
nor UO_1029 (O_1029,N_47773,N_48099);
or UO_1030 (O_1030,N_45386,N_45627);
or UO_1031 (O_1031,N_45732,N_49955);
nor UO_1032 (O_1032,N_47491,N_48834);
or UO_1033 (O_1033,N_46927,N_49721);
xor UO_1034 (O_1034,N_49459,N_47646);
nor UO_1035 (O_1035,N_49974,N_46957);
or UO_1036 (O_1036,N_47326,N_47359);
nor UO_1037 (O_1037,N_47256,N_46963);
xor UO_1038 (O_1038,N_45735,N_46768);
xor UO_1039 (O_1039,N_49916,N_46913);
nor UO_1040 (O_1040,N_46210,N_46916);
nand UO_1041 (O_1041,N_48284,N_45358);
and UO_1042 (O_1042,N_49573,N_47128);
xnor UO_1043 (O_1043,N_47855,N_45298);
nand UO_1044 (O_1044,N_49911,N_46110);
nor UO_1045 (O_1045,N_47060,N_45791);
nand UO_1046 (O_1046,N_48405,N_49363);
and UO_1047 (O_1047,N_49661,N_46013);
or UO_1048 (O_1048,N_46629,N_45734);
xor UO_1049 (O_1049,N_48550,N_48742);
nand UO_1050 (O_1050,N_45600,N_48090);
or UO_1051 (O_1051,N_48971,N_46267);
nor UO_1052 (O_1052,N_46616,N_46162);
and UO_1053 (O_1053,N_47573,N_49433);
nand UO_1054 (O_1054,N_47344,N_45407);
xor UO_1055 (O_1055,N_48915,N_49833);
nand UO_1056 (O_1056,N_45451,N_48042);
or UO_1057 (O_1057,N_46255,N_46079);
xnor UO_1058 (O_1058,N_46829,N_47467);
nand UO_1059 (O_1059,N_45919,N_46652);
and UO_1060 (O_1060,N_49539,N_48478);
xnor UO_1061 (O_1061,N_46825,N_45855);
nor UO_1062 (O_1062,N_48824,N_47902);
nand UO_1063 (O_1063,N_45745,N_49934);
xnor UO_1064 (O_1064,N_47667,N_47267);
nor UO_1065 (O_1065,N_47167,N_49124);
or UO_1066 (O_1066,N_49960,N_49325);
or UO_1067 (O_1067,N_48160,N_46027);
xor UO_1068 (O_1068,N_45896,N_48307);
and UO_1069 (O_1069,N_46653,N_46241);
nor UO_1070 (O_1070,N_46922,N_45236);
xnor UO_1071 (O_1071,N_45526,N_45983);
or UO_1072 (O_1072,N_49012,N_46305);
xor UO_1073 (O_1073,N_47518,N_45597);
or UO_1074 (O_1074,N_49276,N_48700);
and UO_1075 (O_1075,N_46833,N_45766);
or UO_1076 (O_1076,N_46439,N_47391);
and UO_1077 (O_1077,N_46289,N_48419);
nor UO_1078 (O_1078,N_47815,N_49393);
nand UO_1079 (O_1079,N_45874,N_49470);
nor UO_1080 (O_1080,N_49062,N_46867);
or UO_1081 (O_1081,N_47657,N_45157);
nand UO_1082 (O_1082,N_45691,N_46527);
and UO_1083 (O_1083,N_45284,N_47767);
nand UO_1084 (O_1084,N_47999,N_46234);
and UO_1085 (O_1085,N_45501,N_49587);
nor UO_1086 (O_1086,N_48687,N_48107);
and UO_1087 (O_1087,N_49530,N_46129);
nor UO_1088 (O_1088,N_46619,N_47390);
xnor UO_1089 (O_1089,N_46208,N_48273);
nand UO_1090 (O_1090,N_45398,N_49800);
nor UO_1091 (O_1091,N_45064,N_47014);
xor UO_1092 (O_1092,N_46270,N_46045);
and UO_1093 (O_1093,N_46890,N_46682);
nand UO_1094 (O_1094,N_49476,N_49853);
and UO_1095 (O_1095,N_46418,N_46141);
and UO_1096 (O_1096,N_49022,N_49013);
nand UO_1097 (O_1097,N_48258,N_45397);
nor UO_1098 (O_1098,N_49869,N_47288);
nor UO_1099 (O_1099,N_45667,N_45431);
or UO_1100 (O_1100,N_45036,N_46461);
or UO_1101 (O_1101,N_49063,N_49772);
nand UO_1102 (O_1102,N_47264,N_49817);
nand UO_1103 (O_1103,N_45336,N_45147);
and UO_1104 (O_1104,N_45596,N_48920);
and UO_1105 (O_1105,N_48186,N_46485);
and UO_1106 (O_1106,N_49888,N_47001);
and UO_1107 (O_1107,N_49643,N_48917);
nor UO_1108 (O_1108,N_46967,N_46060);
nor UO_1109 (O_1109,N_46997,N_49002);
and UO_1110 (O_1110,N_49912,N_45048);
nand UO_1111 (O_1111,N_45346,N_47197);
or UO_1112 (O_1112,N_46770,N_49086);
and UO_1113 (O_1113,N_45287,N_45821);
xor UO_1114 (O_1114,N_46486,N_45020);
or UO_1115 (O_1115,N_47071,N_47585);
or UO_1116 (O_1116,N_49732,N_45078);
xnor UO_1117 (O_1117,N_49484,N_49918);
nand UO_1118 (O_1118,N_48073,N_47166);
or UO_1119 (O_1119,N_45421,N_48978);
nor UO_1120 (O_1120,N_48597,N_48835);
nand UO_1121 (O_1121,N_48772,N_48506);
nand UO_1122 (O_1122,N_45616,N_46839);
nand UO_1123 (O_1123,N_47611,N_46381);
and UO_1124 (O_1124,N_48927,N_46934);
xnor UO_1125 (O_1125,N_49599,N_46565);
nor UO_1126 (O_1126,N_45971,N_49519);
or UO_1127 (O_1127,N_45426,N_45097);
nand UO_1128 (O_1128,N_47590,N_46759);
or UO_1129 (O_1129,N_45879,N_48310);
xnor UO_1130 (O_1130,N_47419,N_45300);
nor UO_1131 (O_1131,N_46407,N_47997);
and UO_1132 (O_1132,N_45962,N_45891);
nor UO_1133 (O_1133,N_48007,N_48318);
and UO_1134 (O_1134,N_49818,N_47408);
and UO_1135 (O_1135,N_46729,N_47807);
or UO_1136 (O_1136,N_49439,N_47175);
nand UO_1137 (O_1137,N_47709,N_48980);
nand UO_1138 (O_1138,N_46826,N_49527);
nand UO_1139 (O_1139,N_47330,N_47555);
nand UO_1140 (O_1140,N_46420,N_47584);
or UO_1141 (O_1141,N_46218,N_45063);
nor UO_1142 (O_1142,N_46063,N_49044);
or UO_1143 (O_1143,N_49709,N_49384);
xnor UO_1144 (O_1144,N_49068,N_46391);
xnor UO_1145 (O_1145,N_49206,N_45118);
xor UO_1146 (O_1146,N_46048,N_45170);
or UO_1147 (O_1147,N_45105,N_49120);
xnor UO_1148 (O_1148,N_45331,N_49634);
and UO_1149 (O_1149,N_48456,N_45458);
and UO_1150 (O_1150,N_47793,N_45408);
nor UO_1151 (O_1151,N_46424,N_46007);
nor UO_1152 (O_1152,N_48746,N_49273);
nor UO_1153 (O_1153,N_47978,N_46161);
nand UO_1154 (O_1154,N_45185,N_47922);
xnor UO_1155 (O_1155,N_48972,N_46472);
nand UO_1156 (O_1156,N_46799,N_47685);
nor UO_1157 (O_1157,N_45785,N_45031);
nand UO_1158 (O_1158,N_47163,N_49368);
or UO_1159 (O_1159,N_46084,N_47832);
xor UO_1160 (O_1160,N_47058,N_47899);
and UO_1161 (O_1161,N_49332,N_49740);
or UO_1162 (O_1162,N_48880,N_48652);
and UO_1163 (O_1163,N_49909,N_49211);
and UO_1164 (O_1164,N_49764,N_49078);
nand UO_1165 (O_1165,N_46666,N_48490);
xor UO_1166 (O_1166,N_46959,N_49370);
and UO_1167 (O_1167,N_49020,N_47854);
nand UO_1168 (O_1168,N_47193,N_46252);
xnor UO_1169 (O_1169,N_48842,N_48856);
or UO_1170 (O_1170,N_47565,N_45067);
nand UO_1171 (O_1171,N_46151,N_49447);
and UO_1172 (O_1172,N_49594,N_49275);
nand UO_1173 (O_1173,N_47299,N_45906);
nand UO_1174 (O_1174,N_45603,N_45900);
nor UO_1175 (O_1175,N_46740,N_47062);
xnor UO_1176 (O_1176,N_47019,N_47325);
or UO_1177 (O_1177,N_47313,N_47024);
nand UO_1178 (O_1178,N_47817,N_45291);
or UO_1179 (O_1179,N_48023,N_47936);
xor UO_1180 (O_1180,N_47921,N_45214);
or UO_1181 (O_1181,N_47939,N_47457);
nor UO_1182 (O_1182,N_47082,N_48803);
nor UO_1183 (O_1183,N_49239,N_48300);
xnor UO_1184 (O_1184,N_45023,N_47430);
and UO_1185 (O_1185,N_49676,N_47933);
and UO_1186 (O_1186,N_47598,N_49352);
and UO_1187 (O_1187,N_46494,N_47168);
nand UO_1188 (O_1188,N_47374,N_46265);
nand UO_1189 (O_1189,N_47208,N_48067);
nor UO_1190 (O_1190,N_46520,N_46627);
or UO_1191 (O_1191,N_48928,N_45150);
and UO_1192 (O_1192,N_48986,N_49092);
nand UO_1193 (O_1193,N_48977,N_47553);
or UO_1194 (O_1194,N_46846,N_47373);
or UO_1195 (O_1195,N_46999,N_47202);
nor UO_1196 (O_1196,N_48925,N_48213);
nor UO_1197 (O_1197,N_45638,N_47945);
and UO_1198 (O_1198,N_45805,N_45781);
nor UO_1199 (O_1199,N_45591,N_45470);
nand UO_1200 (O_1200,N_48452,N_45664);
nand UO_1201 (O_1201,N_49018,N_46953);
xor UO_1202 (O_1202,N_49984,N_46361);
nand UO_1203 (O_1203,N_48298,N_49247);
or UO_1204 (O_1204,N_47434,N_47451);
nor UO_1205 (O_1205,N_49723,N_49576);
or UO_1206 (O_1206,N_47200,N_45968);
nand UO_1207 (O_1207,N_48086,N_46087);
or UO_1208 (O_1208,N_45279,N_48581);
and UO_1209 (O_1209,N_45774,N_47652);
or UO_1210 (O_1210,N_45404,N_47460);
or UO_1211 (O_1211,N_45019,N_46685);
nor UO_1212 (O_1212,N_46038,N_47607);
nor UO_1213 (O_1213,N_49672,N_49449);
xnor UO_1214 (O_1214,N_45138,N_47397);
or UO_1215 (O_1215,N_49720,N_48421);
nor UO_1216 (O_1216,N_47778,N_45988);
nand UO_1217 (O_1217,N_47009,N_49142);
nor UO_1218 (O_1218,N_46507,N_46640);
nand UO_1219 (O_1219,N_48740,N_45162);
nand UO_1220 (O_1220,N_48181,N_49613);
xor UO_1221 (O_1221,N_49792,N_45549);
nor UO_1222 (O_1222,N_45655,N_47977);
nand UO_1223 (O_1223,N_46465,N_45550);
and UO_1224 (O_1224,N_45888,N_47316);
xnor UO_1225 (O_1225,N_45340,N_46448);
and UO_1226 (O_1226,N_45168,N_48548);
xnor UO_1227 (O_1227,N_47884,N_46187);
or UO_1228 (O_1228,N_47580,N_45207);
xnor UO_1229 (O_1229,N_45141,N_47260);
or UO_1230 (O_1230,N_45809,N_45949);
nand UO_1231 (O_1231,N_46610,N_45139);
nor UO_1232 (O_1232,N_46476,N_48557);
xor UO_1233 (O_1233,N_46601,N_45399);
xor UO_1234 (O_1234,N_45051,N_47477);
nand UO_1235 (O_1235,N_49842,N_48320);
nand UO_1236 (O_1236,N_49406,N_46581);
nand UO_1237 (O_1237,N_47849,N_46611);
and UO_1238 (O_1238,N_47713,N_49808);
nor UO_1239 (O_1239,N_49230,N_47164);
nor UO_1240 (O_1240,N_47358,N_49169);
and UO_1241 (O_1241,N_45181,N_48000);
nor UO_1242 (O_1242,N_46203,N_47004);
or UO_1243 (O_1243,N_48753,N_49954);
or UO_1244 (O_1244,N_48276,N_45579);
nand UO_1245 (O_1245,N_49099,N_47721);
and UO_1246 (O_1246,N_47900,N_45531);
xnor UO_1247 (O_1247,N_48819,N_45542);
nand UO_1248 (O_1248,N_47030,N_47632);
xnor UO_1249 (O_1249,N_47080,N_48795);
or UO_1250 (O_1250,N_48096,N_45870);
xor UO_1251 (O_1251,N_48031,N_47930);
nand UO_1252 (O_1252,N_49600,N_45330);
and UO_1253 (O_1253,N_46675,N_46124);
nand UO_1254 (O_1254,N_47833,N_46548);
xor UO_1255 (O_1255,N_48381,N_46462);
xnor UO_1256 (O_1256,N_48974,N_46571);
nor UO_1257 (O_1257,N_45422,N_46456);
or UO_1258 (O_1258,N_48234,N_47471);
or UO_1259 (O_1259,N_46870,N_46150);
or UO_1260 (O_1260,N_46054,N_47960);
nand UO_1261 (O_1261,N_47860,N_48733);
xor UO_1262 (O_1262,N_49883,N_45267);
or UO_1263 (O_1263,N_48013,N_45246);
xnor UO_1264 (O_1264,N_45779,N_45240);
nor UO_1265 (O_1265,N_46681,N_47426);
xnor UO_1266 (O_1266,N_47668,N_47976);
nor UO_1267 (O_1267,N_47143,N_45341);
and UO_1268 (O_1268,N_46064,N_49190);
nor UO_1269 (O_1269,N_49199,N_46528);
xnor UO_1270 (O_1270,N_47522,N_49491);
xor UO_1271 (O_1271,N_45282,N_47744);
xor UO_1272 (O_1272,N_49145,N_47624);
xor UO_1273 (O_1273,N_48333,N_45861);
nor UO_1274 (O_1274,N_46517,N_48015);
or UO_1275 (O_1275,N_48534,N_45512);
and UO_1276 (O_1276,N_46636,N_48838);
or UO_1277 (O_1277,N_48999,N_45739);
and UO_1278 (O_1278,N_46690,N_47823);
or UO_1279 (O_1279,N_46698,N_45746);
nor UO_1280 (O_1280,N_46268,N_46009);
nand UO_1281 (O_1281,N_47609,N_45862);
nand UO_1282 (O_1282,N_48290,N_45275);
nand UO_1283 (O_1283,N_49728,N_45126);
nand UO_1284 (O_1284,N_49683,N_47211);
nand UO_1285 (O_1285,N_49781,N_47162);
xor UO_1286 (O_1286,N_45814,N_48675);
or UO_1287 (O_1287,N_48511,N_49862);
or UO_1288 (O_1288,N_47205,N_45915);
nor UO_1289 (O_1289,N_49601,N_48145);
nor UO_1290 (O_1290,N_47576,N_46595);
xor UO_1291 (O_1291,N_49851,N_48313);
nor UO_1292 (O_1292,N_48853,N_49942);
nand UO_1293 (O_1293,N_46898,N_48524);
nand UO_1294 (O_1294,N_49902,N_46644);
nor UO_1295 (O_1295,N_48321,N_45528);
nor UO_1296 (O_1296,N_49658,N_46805);
or UO_1297 (O_1297,N_48505,N_48400);
xnor UO_1298 (O_1298,N_47136,N_49133);
or UO_1299 (O_1299,N_45268,N_46792);
xnor UO_1300 (O_1300,N_47615,N_47909);
nor UO_1301 (O_1301,N_46684,N_46035);
nor UO_1302 (O_1302,N_49836,N_45933);
xor UO_1303 (O_1303,N_45102,N_45134);
xor UO_1304 (O_1304,N_49220,N_47425);
nand UO_1305 (O_1305,N_47443,N_49141);
nor UO_1306 (O_1306,N_46097,N_46766);
and UO_1307 (O_1307,N_48385,N_48734);
xor UO_1308 (O_1308,N_46401,N_45885);
or UO_1309 (O_1309,N_46416,N_47279);
or UO_1310 (O_1310,N_45335,N_46348);
and UO_1311 (O_1311,N_45787,N_46077);
and UO_1312 (O_1312,N_45121,N_45058);
or UO_1313 (O_1313,N_49024,N_48894);
and UO_1314 (O_1314,N_47820,N_45069);
nor UO_1315 (O_1315,N_47926,N_49735);
nor UO_1316 (O_1316,N_45143,N_46772);
and UO_1317 (O_1317,N_49979,N_46718);
xor UO_1318 (O_1318,N_46378,N_45966);
nand UO_1319 (O_1319,N_46657,N_45659);
nand UO_1320 (O_1320,N_45125,N_46794);
and UO_1321 (O_1321,N_48326,N_45110);
nand UO_1322 (O_1322,N_47851,N_45913);
or UO_1323 (O_1323,N_45969,N_45713);
xnor UO_1324 (O_1324,N_49249,N_46602);
or UO_1325 (O_1325,N_48775,N_49931);
nor UO_1326 (O_1326,N_48789,N_47380);
nor UO_1327 (O_1327,N_49639,N_49381);
or UO_1328 (O_1328,N_48574,N_46050);
and UO_1329 (O_1329,N_45486,N_48272);
nand UO_1330 (O_1330,N_45191,N_49844);
nand UO_1331 (O_1331,N_46474,N_46955);
nand UO_1332 (O_1332,N_48758,N_49671);
nor UO_1333 (O_1333,N_48459,N_48194);
nor UO_1334 (O_1334,N_49366,N_48203);
and UO_1335 (O_1335,N_48233,N_49418);
nor UO_1336 (O_1336,N_47365,N_47724);
nand UO_1337 (O_1337,N_48699,N_47194);
or UO_1338 (O_1338,N_48576,N_48480);
and UO_1339 (O_1339,N_46984,N_47423);
and UO_1340 (O_1340,N_47604,N_49655);
nand UO_1341 (O_1341,N_48692,N_47394);
nor UO_1342 (O_1342,N_47865,N_47554);
or UO_1343 (O_1343,N_46179,N_49702);
or UO_1344 (O_1344,N_46701,N_47182);
xor UO_1345 (O_1345,N_45183,N_47324);
nand UO_1346 (O_1346,N_46335,N_45158);
xor UO_1347 (O_1347,N_45650,N_45071);
xnor UO_1348 (O_1348,N_49291,N_48358);
or UO_1349 (O_1349,N_49882,N_47932);
or UO_1350 (O_1350,N_49485,N_48560);
nor UO_1351 (O_1351,N_45264,N_49413);
and UO_1352 (O_1352,N_46213,N_47507);
nor UO_1353 (O_1353,N_49894,N_48997);
nand UO_1354 (O_1354,N_48417,N_46696);
nor UO_1355 (O_1355,N_46375,N_48168);
nand UO_1356 (O_1356,N_47206,N_48256);
and UO_1357 (O_1357,N_48923,N_46186);
nor UO_1358 (O_1358,N_48422,N_45079);
or UO_1359 (O_1359,N_46176,N_46492);
or UO_1360 (O_1360,N_49398,N_45553);
nor UO_1361 (O_1361,N_48363,N_46232);
nand UO_1362 (O_1362,N_46272,N_49924);
xnor UO_1363 (O_1363,N_48564,N_47226);
nor UO_1364 (O_1364,N_47898,N_49901);
nand UO_1365 (O_1365,N_48445,N_45438);
and UO_1366 (O_1366,N_48061,N_45286);
and UO_1367 (O_1367,N_49641,N_48606);
or UO_1368 (O_1368,N_47572,N_47061);
nand UO_1369 (O_1369,N_45419,N_48521);
and UO_1370 (O_1370,N_47605,N_49876);
xnor UO_1371 (O_1371,N_48280,N_47783);
nor UO_1372 (O_1372,N_46436,N_48398);
or UO_1373 (O_1373,N_47078,N_47692);
xor UO_1374 (O_1374,N_46251,N_49940);
nor UO_1375 (O_1375,N_46153,N_49388);
nand UO_1376 (O_1376,N_48901,N_46874);
nor UO_1377 (O_1377,N_46851,N_47835);
xor UO_1378 (O_1378,N_49408,N_45859);
nand UO_1379 (O_1379,N_49588,N_45043);
nand UO_1380 (O_1380,N_49158,N_47437);
or UO_1381 (O_1381,N_47596,N_45136);
nand UO_1382 (O_1382,N_46506,N_47287);
nand UO_1383 (O_1383,N_47861,N_45376);
nor UO_1384 (O_1384,N_45155,N_46453);
nand UO_1385 (O_1385,N_46298,N_45363);
nand UO_1386 (O_1386,N_47368,N_47023);
nor UO_1387 (O_1387,N_49783,N_45978);
nand UO_1388 (O_1388,N_46591,N_45302);
and UO_1389 (O_1389,N_48388,N_46532);
nor UO_1390 (O_1390,N_46163,N_45062);
xnor UO_1391 (O_1391,N_47577,N_45860);
and UO_1392 (O_1392,N_46549,N_49094);
or UO_1393 (O_1393,N_49978,N_49402);
or UO_1394 (O_1394,N_49759,N_48241);
nand UO_1395 (O_1395,N_48127,N_47717);
and UO_1396 (O_1396,N_49500,N_49448);
xor UO_1397 (O_1397,N_48240,N_45205);
and UO_1398 (O_1398,N_48484,N_49156);
or UO_1399 (O_1399,N_48406,N_49285);
or UO_1400 (O_1400,N_49422,N_48188);
and UO_1401 (O_1401,N_45867,N_45918);
xnor UO_1402 (O_1402,N_49151,N_46158);
nand UO_1403 (O_1403,N_47404,N_45716);
nor UO_1404 (O_1404,N_49884,N_47931);
nor UO_1405 (O_1405,N_47032,N_45818);
xnor UO_1406 (O_1406,N_47971,N_45685);
nor UO_1407 (O_1407,N_45630,N_48799);
and UO_1408 (O_1408,N_45032,N_46988);
nand UO_1409 (O_1409,N_48616,N_45499);
or UO_1410 (O_1410,N_48680,N_47220);
or UO_1411 (O_1411,N_48629,N_48156);
nand UO_1412 (O_1412,N_45704,N_47914);
or UO_1413 (O_1413,N_49653,N_49204);
xnor UO_1414 (O_1414,N_45222,N_49928);
xor UO_1415 (O_1415,N_46356,N_47980);
or UO_1416 (O_1416,N_46421,N_47156);
or UO_1417 (O_1417,N_48570,N_48340);
nor UO_1418 (O_1418,N_46410,N_49170);
and UO_1419 (O_1419,N_46293,N_46596);
and UO_1420 (O_1420,N_49430,N_47742);
nor UO_1421 (O_1421,N_46031,N_46873);
xor UO_1422 (O_1422,N_46903,N_49117);
xnor UO_1423 (O_1423,N_48659,N_47950);
nand UO_1424 (O_1424,N_47571,N_48615);
xnor UO_1425 (O_1425,N_47236,N_47561);
nor UO_1426 (O_1426,N_48447,N_49824);
and UO_1427 (O_1427,N_49202,N_46318);
and UO_1428 (O_1428,N_49825,N_46700);
and UO_1429 (O_1429,N_49299,N_45784);
xnor UO_1430 (O_1430,N_48526,N_47230);
or UO_1431 (O_1431,N_46521,N_48288);
or UO_1432 (O_1432,N_47526,N_49395);
or UO_1433 (O_1433,N_46524,N_45465);
or UO_1434 (O_1434,N_45487,N_46352);
xnor UO_1435 (O_1435,N_49307,N_49747);
and UO_1436 (O_1436,N_48372,N_47842);
xnor UO_1437 (O_1437,N_46801,N_45873);
xnor UO_1438 (O_1438,N_48057,N_48522);
and UO_1439 (O_1439,N_49001,N_49803);
or UO_1440 (O_1440,N_48900,N_47484);
and UO_1441 (O_1441,N_47276,N_49123);
xnor UO_1442 (O_1442,N_46834,N_48476);
or UO_1443 (O_1443,N_47262,N_49482);
nor UO_1444 (O_1444,N_46047,N_46529);
xor UO_1445 (O_1445,N_45360,N_48115);
nand UO_1446 (O_1446,N_47871,N_48047);
nor UO_1447 (O_1447,N_45095,N_49999);
nand UO_1448 (O_1448,N_49574,N_45070);
or UO_1449 (O_1449,N_46144,N_48865);
or UO_1450 (O_1450,N_45833,N_48747);
or UO_1451 (O_1451,N_45965,N_45710);
nand UO_1452 (O_1452,N_45323,N_46533);
xor UO_1453 (O_1453,N_49762,N_46445);
or UO_1454 (O_1454,N_45952,N_49790);
or UO_1455 (O_1455,N_45517,N_48399);
nand UO_1456 (O_1456,N_47497,N_45123);
nand UO_1457 (O_1457,N_49538,N_47789);
nand UO_1458 (O_1458,N_48614,N_46316);
nand UO_1459 (O_1459,N_47037,N_47989);
nand UO_1460 (O_1460,N_48924,N_49463);
and UO_1461 (O_1461,N_47415,N_48254);
xor UO_1462 (O_1462,N_47073,N_49936);
nor UO_1463 (O_1463,N_45975,N_45932);
and UO_1464 (O_1464,N_47088,N_45680);
and UO_1465 (O_1465,N_49893,N_46824);
or UO_1466 (O_1466,N_48108,N_45743);
or UO_1467 (O_1467,N_45629,N_49529);
xnor UO_1468 (O_1468,N_49930,N_49770);
xnor UO_1469 (O_1469,N_49059,N_47165);
xor UO_1470 (O_1470,N_45084,N_49680);
xnor UO_1471 (O_1471,N_46534,N_49972);
and UO_1472 (O_1472,N_46466,N_46730);
or UO_1473 (O_1473,N_48216,N_45524);
nand UO_1474 (O_1474,N_48896,N_48766);
nor UO_1475 (O_1475,N_47794,N_49396);
and UO_1476 (O_1476,N_49236,N_47890);
or UO_1477 (O_1477,N_49938,N_49959);
xor UO_1478 (O_1478,N_47405,N_49265);
nor UO_1479 (O_1479,N_45003,N_49621);
and UO_1480 (O_1480,N_45034,N_46283);
nor UO_1481 (O_1481,N_48599,N_47892);
nand UO_1482 (O_1482,N_48184,N_45617);
nand UO_1483 (O_1483,N_49595,N_48449);
or UO_1484 (O_1484,N_48571,N_48205);
and UO_1485 (O_1485,N_46368,N_46044);
xnor UO_1486 (O_1486,N_47021,N_48934);
nand UO_1487 (O_1487,N_49510,N_49845);
xnor UO_1488 (O_1488,N_46546,N_47741);
and UO_1489 (O_1489,N_45649,N_48604);
or UO_1490 (O_1490,N_49516,N_49031);
nand UO_1491 (O_1491,N_46325,N_47916);
nor UO_1492 (O_1492,N_46463,N_47265);
and UO_1493 (O_1493,N_49269,N_45720);
and UO_1494 (O_1494,N_45807,N_45950);
or UO_1495 (O_1495,N_49392,N_45558);
nand UO_1496 (O_1496,N_46357,N_49945);
nor UO_1497 (O_1497,N_47377,N_45628);
or UO_1498 (O_1498,N_47578,N_46641);
or UO_1499 (O_1499,N_45285,N_49039);
nor UO_1500 (O_1500,N_46412,N_49531);
nor UO_1501 (O_1501,N_49858,N_45400);
nor UO_1502 (O_1502,N_47119,N_48135);
nor UO_1503 (O_1503,N_49181,N_47282);
or UO_1504 (O_1504,N_46136,N_48533);
nor UO_1505 (O_1505,N_46426,N_46734);
nor UO_1506 (O_1506,N_47688,N_48936);
nor UO_1507 (O_1507,N_45886,N_46183);
or UO_1508 (O_1508,N_49244,N_48755);
nand UO_1509 (O_1509,N_45076,N_48566);
and UO_1510 (O_1510,N_45619,N_45372);
nor UO_1511 (O_1511,N_46493,N_45610);
xor UO_1512 (O_1512,N_49583,N_48736);
nor UO_1513 (O_1513,N_47730,N_45452);
and UO_1514 (O_1514,N_49209,N_47258);
or UO_1515 (O_1515,N_48470,N_48943);
and UO_1516 (O_1516,N_47195,N_45742);
xnor UO_1517 (O_1517,N_48518,N_46780);
or UO_1518 (O_1518,N_47372,N_49537);
nor UO_1519 (O_1519,N_49981,N_47517);
nand UO_1520 (O_1520,N_47441,N_47660);
xnor UO_1521 (O_1521,N_48407,N_49612);
xor UO_1522 (O_1522,N_48777,N_46715);
nor UO_1523 (O_1523,N_46938,N_48037);
nand UO_1524 (O_1524,N_48910,N_45428);
nand UO_1525 (O_1525,N_47746,N_48685);
xor UO_1526 (O_1526,N_48538,N_46891);
nor UO_1527 (O_1527,N_47102,N_48257);
nand UO_1528 (O_1528,N_47834,N_49290);
nand UO_1529 (O_1529,N_46995,N_45219);
or UO_1530 (O_1530,N_47601,N_49499);
or UO_1531 (O_1531,N_46473,N_49896);
and UO_1532 (O_1532,N_45989,N_49831);
nand UO_1533 (O_1533,N_47048,N_45557);
nor UO_1534 (O_1534,N_45109,N_48840);
nand UO_1535 (O_1535,N_45208,N_48237);
nor UO_1536 (O_1536,N_48274,N_48881);
xor UO_1537 (O_1537,N_47227,N_46350);
xnor UO_1538 (O_1538,N_49088,N_46712);
xor UO_1539 (O_1539,N_45401,N_46655);
nand UO_1540 (O_1540,N_46883,N_45693);
nor UO_1541 (O_1541,N_46205,N_46835);
nand UO_1542 (O_1542,N_46847,N_45736);
nor UO_1543 (O_1543,N_48136,N_49157);
or UO_1544 (O_1544,N_47906,N_49298);
nor UO_1545 (O_1545,N_48580,N_49565);
nor UO_1546 (O_1546,N_48908,N_48621);
and UO_1547 (O_1547,N_45651,N_45418);
nor UO_1548 (O_1548,N_49254,N_47473);
nand UO_1549 (O_1549,N_45796,N_45765);
nand UO_1550 (O_1550,N_45354,N_45537);
or UO_1551 (O_1551,N_49736,N_48357);
nor UO_1552 (O_1552,N_45283,N_45940);
nand UO_1553 (O_1553,N_48072,N_46259);
xnor UO_1554 (O_1554,N_47063,N_45057);
nor UO_1555 (O_1555,N_47346,N_45976);
and UO_1556 (O_1556,N_47701,N_45072);
or UO_1557 (O_1557,N_49391,N_49675);
nand UO_1558 (O_1558,N_48493,N_47981);
nand UO_1559 (O_1559,N_45665,N_45445);
nor UO_1560 (O_1560,N_46423,N_46143);
and UO_1561 (O_1561,N_47676,N_46864);
xnor UO_1562 (O_1562,N_46790,N_46114);
xnor UO_1563 (O_1563,N_48726,N_48312);
or UO_1564 (O_1564,N_47533,N_47283);
nor UO_1565 (O_1565,N_48244,N_48839);
nand UO_1566 (O_1566,N_49863,N_47819);
xnor UO_1567 (O_1567,N_46102,N_48105);
nand UO_1568 (O_1568,N_46608,N_45827);
xnor UO_1569 (O_1569,N_49848,N_48356);
nand UO_1570 (O_1570,N_48345,N_49172);
or UO_1571 (O_1571,N_45877,N_47159);
nor UO_1572 (O_1572,N_47508,N_46408);
xnor UO_1573 (O_1573,N_49726,N_48411);
xor UO_1574 (O_1574,N_47563,N_45179);
and UO_1575 (O_1575,N_46917,N_49339);
or UO_1576 (O_1576,N_46131,N_46470);
nand UO_1577 (O_1577,N_46968,N_46248);
or UO_1578 (O_1578,N_45817,N_46638);
or UO_1579 (O_1579,N_45113,N_46387);
nand UO_1580 (O_1580,N_49115,N_49372);
nor UO_1581 (O_1581,N_47538,N_46660);
nand UO_1582 (O_1582,N_46249,N_49311);
nor UO_1583 (O_1583,N_46818,N_48688);
and UO_1584 (O_1584,N_46431,N_45053);
nor UO_1585 (O_1585,N_49432,N_47661);
and UO_1586 (O_1586,N_49175,N_46823);
and UO_1587 (O_1587,N_49409,N_46380);
nor UO_1588 (O_1588,N_48453,N_46779);
and UO_1589 (O_1589,N_45899,N_47987);
nor UO_1590 (O_1590,N_47191,N_45229);
nor UO_1591 (O_1591,N_47366,N_49812);
xnor UO_1592 (O_1592,N_45254,N_48263);
nor UO_1593 (O_1593,N_48698,N_47803);
or UO_1594 (O_1594,N_47393,N_45189);
or UO_1595 (O_1595,N_47011,N_48804);
or UO_1596 (O_1596,N_46290,N_46879);
nor UO_1597 (O_1597,N_45669,N_46003);
nand UO_1598 (O_1598,N_48519,N_49083);
nor UO_1599 (O_1599,N_47022,N_47719);
nand UO_1600 (O_1600,N_48785,N_45808);
nand UO_1601 (O_1601,N_45262,N_49528);
and UO_1602 (O_1602,N_49237,N_49150);
nor UO_1603 (O_1603,N_46560,N_47015);
nand UO_1604 (O_1604,N_46212,N_48380);
and UO_1605 (O_1605,N_47665,N_46904);
or UO_1606 (O_1606,N_49210,N_46491);
or UO_1607 (O_1607,N_49279,N_45681);
and UO_1608 (O_1608,N_49314,N_47856);
and UO_1609 (O_1609,N_45159,N_48651);
nand UO_1610 (O_1610,N_48295,N_48189);
and UO_1611 (O_1611,N_49607,N_47438);
or UO_1612 (O_1612,N_45985,N_45972);
nand UO_1613 (O_1613,N_49364,N_46008);
xnor UO_1614 (O_1614,N_45467,N_47726);
and UO_1615 (O_1615,N_47149,N_46366);
nor UO_1616 (O_1616,N_45831,N_45374);
xnor UO_1617 (O_1617,N_48823,N_46777);
or UO_1618 (O_1618,N_48948,N_46053);
and UO_1619 (O_1619,N_49129,N_49136);
or UO_1620 (O_1620,N_49076,N_45245);
or UO_1621 (O_1621,N_45602,N_45006);
or UO_1622 (O_1622,N_47606,N_46620);
and UO_1623 (O_1623,N_45199,N_46147);
or UO_1624 (O_1624,N_46775,N_47500);
and UO_1625 (O_1625,N_49514,N_49264);
and UO_1626 (O_1626,N_45068,N_48005);
and UO_1627 (O_1627,N_45682,N_49948);
nand UO_1628 (O_1628,N_48876,N_45402);
or UO_1629 (O_1629,N_46437,N_45697);
and UO_1630 (O_1630,N_45694,N_49775);
nor UO_1631 (O_1631,N_46080,N_45883);
xnor UO_1632 (O_1632,N_47447,N_49328);
nor UO_1633 (O_1633,N_46723,N_48719);
and UO_1634 (O_1634,N_48985,N_47338);
and UO_1635 (O_1635,N_46284,N_49354);
and UO_1636 (O_1636,N_48968,N_49906);
nand UO_1637 (O_1637,N_45987,N_49212);
nor UO_1638 (O_1638,N_49718,N_45127);
or UO_1639 (O_1639,N_48281,N_49712);
and UO_1640 (O_1640,N_49286,N_45017);
and UO_1641 (O_1641,N_49923,N_48416);
nor UO_1642 (O_1642,N_46320,N_45046);
nand UO_1643 (O_1643,N_48891,N_49937);
nand UO_1644 (O_1644,N_48022,N_49113);
nor UO_1645 (O_1645,N_48339,N_45175);
xnor UO_1646 (O_1646,N_47663,N_46207);
xnor UO_1647 (O_1647,N_49535,N_46152);
nor UO_1648 (O_1648,N_46105,N_47628);
and UO_1649 (O_1649,N_45461,N_46443);
or UO_1650 (O_1650,N_45618,N_46459);
xnor UO_1651 (O_1651,N_45294,N_46542);
and UO_1652 (O_1652,N_47775,N_45251);
nor UO_1653 (O_1653,N_48020,N_45768);
nand UO_1654 (O_1654,N_48327,N_46588);
nor UO_1655 (O_1655,N_48705,N_48752);
and UO_1656 (O_1656,N_48034,N_45148);
or UO_1657 (O_1657,N_48403,N_46331);
nand UO_1658 (O_1658,N_46736,N_45974);
nor UO_1659 (O_1659,N_49780,N_47462);
nand UO_1660 (O_1660,N_49310,N_46172);
nand UO_1661 (O_1661,N_47848,N_47694);
nor UO_1662 (O_1662,N_47493,N_49873);
nor UO_1663 (O_1663,N_48728,N_48481);
nor UO_1664 (O_1664,N_48026,N_47117);
or UO_1665 (O_1665,N_49991,N_49796);
or UO_1666 (O_1666,N_47630,N_46773);
and UO_1667 (O_1667,N_47671,N_45195);
xor UO_1668 (O_1668,N_45390,N_49872);
and UO_1669 (O_1669,N_45345,N_49255);
and UO_1670 (O_1670,N_47666,N_47643);
and UO_1671 (O_1671,N_49473,N_47568);
xor UO_1672 (O_1672,N_47693,N_48964);
xor UO_1673 (O_1673,N_47883,N_45801);
xnor UO_1674 (O_1674,N_49861,N_45454);
nor UO_1675 (O_1675,N_47181,N_46154);
and UO_1676 (O_1676,N_49611,N_46083);
and UO_1677 (O_1677,N_46765,N_49168);
nor UO_1678 (O_1678,N_47486,N_45135);
nand UO_1679 (O_1679,N_46286,N_48483);
or UO_1680 (O_1680,N_48303,N_48214);
nand UO_1681 (O_1681,N_45893,N_46362);
xnor UO_1682 (O_1682,N_47150,N_49245);
xor UO_1683 (O_1683,N_45963,N_47655);
xor UO_1684 (O_1684,N_49797,N_49053);
nor UO_1685 (O_1685,N_48366,N_46427);
nor UO_1686 (O_1686,N_46969,N_48112);
nand UO_1687 (O_1687,N_49045,N_47284);
nand UO_1688 (O_1688,N_49515,N_49194);
xor UO_1689 (O_1689,N_46820,N_48121);
and UO_1690 (O_1690,N_48454,N_45723);
xnor UO_1691 (O_1691,N_45488,N_45523);
nor UO_1692 (O_1692,N_47214,N_49153);
nor UO_1693 (O_1693,N_45555,N_47748);
xor UO_1694 (O_1694,N_47974,N_46545);
nand UO_1695 (O_1695,N_45688,N_48815);
and UO_1696 (O_1696,N_47418,N_48024);
nor UO_1697 (O_1697,N_45349,N_47090);
nor UO_1698 (O_1698,N_48464,N_49288);
nand UO_1699 (O_1699,N_46328,N_49589);
or UO_1700 (O_1700,N_45220,N_49581);
nor UO_1701 (O_1701,N_47074,N_45505);
xnor UO_1702 (O_1702,N_46403,N_49559);
and UO_1703 (O_1703,N_46547,N_45882);
nor UO_1704 (O_1704,N_49627,N_49047);
nand UO_1705 (O_1705,N_47925,N_49619);
nand UO_1706 (O_1706,N_47134,N_46414);
and UO_1707 (O_1707,N_45424,N_48228);
or UO_1708 (O_1708,N_48620,N_47315);
nand UO_1709 (O_1709,N_48858,N_46160);
nor UO_1710 (O_1710,N_48428,N_46821);
and UO_1711 (O_1711,N_48921,N_45483);
nand UO_1712 (O_1712,N_45468,N_48430);
nor UO_1713 (O_1713,N_45339,N_45658);
nor UO_1714 (O_1714,N_49707,N_46751);
and UO_1715 (O_1715,N_46580,N_46257);
and UO_1716 (O_1716,N_49061,N_48270);
xnor UO_1717 (O_1717,N_45946,N_49019);
nand UO_1718 (O_1718,N_48610,N_47765);
or UO_1719 (O_1719,N_48696,N_45029);
or UO_1720 (O_1720,N_48527,N_49347);
or UO_1721 (O_1721,N_45822,N_48931);
and UO_1722 (O_1722,N_49229,N_46812);
nor UO_1723 (O_1723,N_47790,N_45395);
and UO_1724 (O_1724,N_48494,N_47485);
nor UO_1725 (O_1725,N_47261,N_45382);
nor UO_1726 (O_1726,N_45417,N_46276);
nand UO_1727 (O_1727,N_48361,N_46406);
or UO_1728 (O_1728,N_48724,N_47669);
nor UO_1729 (O_1729,N_47696,N_48153);
nand UO_1730 (O_1730,N_49479,N_46933);
nor UO_1731 (O_1731,N_46689,N_46477);
nand UO_1732 (O_1732,N_46651,N_49677);
nor UO_1733 (O_1733,N_46086,N_47000);
nand UO_1734 (O_1734,N_49737,N_46130);
and UO_1735 (O_1735,N_46065,N_45370);
and UO_1736 (O_1736,N_49586,N_45956);
or UO_1737 (O_1737,N_49878,N_47529);
and UO_1738 (O_1738,N_49760,N_47695);
nor UO_1739 (O_1739,N_46011,N_47728);
nor UO_1740 (O_1740,N_48289,N_47689);
nor UO_1741 (O_1741,N_47552,N_46932);
xor UO_1742 (O_1742,N_49542,N_45014);
and UO_1743 (O_1743,N_49914,N_47994);
nand UO_1744 (O_1744,N_45459,N_48708);
xor UO_1745 (O_1745,N_46028,N_48143);
nor UO_1746 (O_1746,N_49635,N_45671);
xnor UO_1747 (O_1747,N_47829,N_49777);
and UO_1748 (O_1748,N_47961,N_49351);
xnor UO_1749 (O_1749,N_47310,N_45366);
nand UO_1750 (O_1750,N_47360,N_48248);
xnor UO_1751 (O_1751,N_45999,N_49744);
or UO_1752 (O_1752,N_48100,N_46885);
nor UO_1753 (O_1753,N_46246,N_47673);
nor UO_1754 (O_1754,N_49551,N_49569);
or UO_1755 (O_1755,N_47242,N_45250);
or UO_1756 (O_1756,N_48551,N_48268);
xor UO_1757 (O_1757,N_47400,N_49345);
and UO_1758 (O_1758,N_46389,N_47494);
and UO_1759 (O_1759,N_47984,N_48944);
xnor UO_1760 (O_1760,N_49152,N_45979);
nand UO_1761 (O_1761,N_45912,N_49501);
nor UO_1762 (O_1762,N_46088,N_48231);
xnor UO_1763 (O_1763,N_45101,N_47885);
and UO_1764 (O_1764,N_45171,N_46871);
nor UO_1765 (O_1765,N_46345,N_47612);
or UO_1766 (O_1766,N_48583,N_45371);
and UO_1767 (O_1767,N_46598,N_45414);
nor UO_1768 (O_1768,N_48473,N_45119);
xor UO_1769 (O_1769,N_48060,N_47297);
xor UO_1770 (O_1770,N_47104,N_47141);
or UO_1771 (O_1771,N_47798,N_48070);
nand UO_1772 (O_1772,N_49885,N_48434);
or UO_1773 (O_1773,N_45026,N_47872);
and UO_1774 (O_1774,N_45235,N_49517);
nand UO_1775 (O_1775,N_49065,N_48970);
nand UO_1776 (O_1776,N_49042,N_48150);
or UO_1777 (O_1777,N_47501,N_47204);
and UO_1778 (O_1778,N_46522,N_49806);
or UO_1779 (O_1779,N_46006,N_49578);
xnor UO_1780 (O_1780,N_46536,N_49452);
xor UO_1781 (O_1781,N_46978,N_45726);
nand UO_1782 (O_1782,N_49608,N_46195);
xor UO_1783 (O_1783,N_48350,N_49110);
xnor UO_1784 (O_1784,N_49223,N_48988);
nor UO_1785 (O_1785,N_48757,N_48297);
xor UO_1786 (O_1786,N_48935,N_48247);
nand UO_1787 (O_1787,N_49773,N_47619);
nand UO_1788 (O_1788,N_46374,N_49741);
or UO_1789 (O_1789,N_45819,N_47969);
or UO_1790 (O_1790,N_46974,N_46211);
nand UO_1791 (O_1791,N_46174,N_48554);
nand UO_1792 (O_1792,N_46029,N_46068);
and UO_1793 (O_1793,N_47228,N_46503);
and UO_1794 (O_1794,N_47278,N_45731);
nor UO_1795 (O_1795,N_45334,N_49319);
or UO_1796 (O_1796,N_49292,N_45673);
xnor UO_1797 (O_1797,N_48913,N_46340);
nand UO_1798 (O_1798,N_46041,N_47557);
and UO_1799 (O_1799,N_47876,N_48401);
xnor UO_1800 (O_1800,N_49336,N_46349);
nand UO_1801 (O_1801,N_46236,N_47332);
nand UO_1802 (O_1802,N_48545,N_45889);
and UO_1803 (O_1803,N_49570,N_45088);
nor UO_1804 (O_1804,N_46973,N_45922);
nor UO_1805 (O_1805,N_49518,N_48776);
nand UO_1806 (O_1806,N_49087,N_48674);
and UO_1807 (O_1807,N_46573,N_45103);
nor UO_1808 (O_1808,N_45775,N_45727);
or UO_1809 (O_1809,N_48374,N_46996);
nand UO_1810 (O_1810,N_47075,N_47291);
and UO_1811 (O_1811,N_45931,N_48235);
or UO_1812 (O_1812,N_46965,N_48332);
nand UO_1813 (O_1813,N_45393,N_46446);
and UO_1814 (O_1814,N_49805,N_48163);
xor UO_1815 (O_1815,N_48383,N_46577);
nand UO_1816 (O_1816,N_46893,N_45595);
nor UO_1817 (O_1817,N_49632,N_48847);
nand UO_1818 (O_1818,N_48055,N_47558);
and UO_1819 (O_1819,N_48192,N_49434);
xnor UO_1820 (O_1820,N_49462,N_49857);
nor UO_1821 (O_1821,N_45525,N_49179);
nor UO_1822 (O_1822,N_45357,N_46148);
and UO_1823 (O_1823,N_47813,N_48002);
and UO_1824 (O_1824,N_47610,N_48071);
and UO_1825 (O_1825,N_47626,N_45212);
nand UO_1826 (O_1826,N_49215,N_49101);
and UO_1827 (O_1827,N_45577,N_47539);
xnor UO_1828 (O_1828,N_48887,N_46062);
or UO_1829 (O_1829,N_45998,N_47515);
xnor UO_1830 (O_1830,N_49572,N_46057);
nor UO_1831 (O_1831,N_48146,N_49017);
xnor UO_1832 (O_1832,N_47640,N_45585);
xor UO_1833 (O_1833,N_48133,N_48797);
nand UO_1834 (O_1834,N_45055,N_48864);
or UO_1835 (O_1835,N_48041,N_49939);
or UO_1836 (O_1836,N_47138,N_45394);
or UO_1837 (O_1837,N_47527,N_49312);
xor UO_1838 (O_1838,N_45646,N_45027);
or UO_1839 (O_1839,N_49160,N_45530);
or UO_1840 (O_1840,N_48492,N_45383);
nand UO_1841 (O_1841,N_46667,N_49765);
and UO_1842 (O_1842,N_47300,N_49754);
nand UO_1843 (O_1843,N_47008,N_45446);
nand UO_1844 (O_1844,N_45496,N_48119);
and UO_1845 (O_1845,N_48991,N_47296);
nand UO_1846 (O_1846,N_49032,N_45318);
xnor UO_1847 (O_1847,N_46724,N_45902);
and UO_1848 (O_1848,N_46688,N_47642);
or UO_1849 (O_1849,N_48516,N_47620);
nor UO_1850 (O_1850,N_49650,N_45705);
and UO_1851 (O_1851,N_48780,N_49891);
or UO_1852 (O_1852,N_45529,N_45961);
and UO_1853 (O_1853,N_49023,N_45799);
nand UO_1854 (O_1854,N_48947,N_48315);
or UO_1855 (O_1855,N_49550,N_48394);
nor UO_1856 (O_1856,N_49014,N_46717);
or UO_1857 (O_1857,N_45255,N_46253);
or UO_1858 (O_1858,N_47002,N_49989);
or UO_1859 (O_1859,N_49996,N_49383);
nor UO_1860 (O_1860,N_49225,N_46707);
nor UO_1861 (O_1861,N_45920,N_49571);
nand UO_1862 (O_1862,N_46264,N_48183);
xnor UO_1863 (O_1863,N_49617,N_45866);
or UO_1864 (O_1864,N_49342,N_48608);
xor UO_1865 (O_1865,N_47207,N_48582);
and UO_1866 (O_1866,N_49058,N_45593);
nor UO_1867 (O_1867,N_45613,N_46947);
nor UO_1868 (O_1868,N_49071,N_46281);
or UO_1869 (O_1869,N_49665,N_46981);
nand UO_1870 (O_1870,N_49163,N_49986);
xnor UO_1871 (O_1871,N_46758,N_47691);
xor UO_1872 (O_1872,N_46618,N_49203);
xnor UO_1873 (O_1873,N_45670,N_49850);
nand UO_1874 (O_1874,N_49794,N_45025);
nor UO_1875 (O_1875,N_48500,N_46376);
nor UO_1876 (O_1876,N_45930,N_49440);
nor UO_1877 (O_1877,N_45843,N_45085);
and UO_1878 (O_1878,N_45708,N_49699);
xor UO_1879 (O_1879,N_48370,N_46887);
and UO_1880 (O_1880,N_45450,N_47570);
and UO_1881 (O_1881,N_48950,N_47942);
xor UO_1882 (O_1882,N_49879,N_46923);
nor UO_1883 (O_1883,N_46808,N_47891);
nor UO_1884 (O_1884,N_47934,N_46987);
and UO_1885 (O_1885,N_46243,N_47845);
xnor UO_1886 (O_1886,N_47996,N_49477);
nor UO_1887 (O_1887,N_47781,N_48807);
or UO_1888 (O_1888,N_45565,N_48907);
and UO_1889 (O_1889,N_49343,N_45476);
nor UO_1890 (O_1890,N_47153,N_49557);
xor UO_1891 (O_1891,N_45356,N_49401);
or UO_1892 (O_1892,N_47348,N_45244);
or UO_1893 (O_1893,N_48679,N_48111);
xor UO_1894 (O_1894,N_49385,N_45296);
and UO_1895 (O_1895,N_46306,N_48215);
nand UO_1896 (O_1896,N_48668,N_48438);
xor UO_1897 (O_1897,N_45641,N_49852);
or UO_1898 (O_1898,N_47314,N_48790);
xnor UO_1899 (O_1899,N_46795,N_46198);
and UO_1900 (O_1900,N_49296,N_48959);
nand UO_1901 (O_1901,N_49839,N_47410);
and UO_1902 (O_1902,N_48530,N_49362);
or UO_1903 (O_1903,N_46563,N_49227);
nor UO_1904 (O_1904,N_48872,N_47421);
nand UO_1905 (O_1905,N_47431,N_46687);
nand UO_1906 (O_1906,N_49951,N_47131);
and UO_1907 (O_1907,N_46930,N_45479);
nand UO_1908 (O_1908,N_47142,N_48132);
nand UO_1909 (O_1909,N_49185,N_48778);
or UO_1910 (O_1910,N_49358,N_47007);
xor UO_1911 (O_1911,N_46262,N_47145);
and UO_1912 (O_1912,N_49786,N_46831);
and UO_1913 (O_1913,N_48004,N_45797);
or UO_1914 (O_1914,N_46321,N_46072);
or UO_1915 (O_1915,N_49346,N_47791);
and UO_1916 (O_1916,N_49691,N_45436);
xor UO_1917 (O_1917,N_46390,N_48391);
nand UO_1918 (O_1918,N_45642,N_45733);
nand UO_1919 (O_1919,N_46002,N_48703);
and UO_1920 (O_1920,N_45560,N_48444);
or UO_1921 (O_1921,N_48437,N_48344);
xor UO_1922 (O_1922,N_48613,N_47528);
nand UO_1923 (O_1923,N_49222,N_48420);
nand UO_1924 (O_1924,N_49483,N_49887);
nand UO_1925 (O_1925,N_47133,N_49035);
xor UO_1926 (O_1926,N_48635,N_47385);
or UO_1927 (O_1927,N_47737,N_46379);
nand UO_1928 (O_1928,N_47238,N_45575);
and UO_1929 (O_1929,N_47718,N_49969);
nand UO_1930 (O_1930,N_46347,N_46351);
nand UO_1931 (O_1931,N_49758,N_47309);
nand UO_1932 (O_1932,N_49592,N_46338);
nand UO_1933 (O_1933,N_46405,N_47852);
xnor UO_1934 (O_1934,N_47893,N_47255);
nor UO_1935 (O_1935,N_45652,N_48983);
nand UO_1936 (O_1936,N_47743,N_47077);
nor UO_1937 (O_1937,N_45749,N_48525);
nor UO_1938 (O_1938,N_48569,N_45995);
nor UO_1939 (O_1939,N_46894,N_47151);
nand UO_1940 (O_1940,N_45928,N_48371);
nor UO_1941 (O_1941,N_47729,N_46848);
and UO_1942 (O_1942,N_47686,N_48032);
and UO_1943 (O_1943,N_47389,N_47114);
nor UO_1944 (O_1944,N_49591,N_49037);
xor UO_1945 (O_1945,N_49628,N_49171);
nor UO_1946 (O_1946,N_48514,N_46703);
nor UO_1947 (O_1947,N_46674,N_45448);
xor UO_1948 (O_1948,N_48059,N_49889);
nand UO_1949 (O_1949,N_46287,N_49355);
nand UO_1950 (O_1950,N_47386,N_46800);
and UO_1951 (O_1951,N_48852,N_47170);
or UO_1952 (O_1952,N_49261,N_45639);
and UO_1953 (O_1953,N_47186,N_49905);
nor UO_1954 (O_1954,N_49523,N_46370);
and UO_1955 (O_1955,N_49259,N_49173);
xor UO_1956 (O_1956,N_46669,N_49585);
and UO_1957 (O_1957,N_49337,N_49696);
or UO_1958 (O_1958,N_47550,N_45444);
or UO_1959 (O_1959,N_49742,N_47502);
xor UO_1960 (O_1960,N_46886,N_48251);
and UO_1961 (O_1961,N_49475,N_47826);
nor UO_1962 (O_1962,N_48439,N_46726);
xor UO_1963 (O_1963,N_48139,N_47305);
or UO_1964 (O_1964,N_45762,N_45892);
nor UO_1965 (O_1965,N_48523,N_49871);
or UO_1966 (O_1966,N_46646,N_49503);
or UO_1967 (O_1967,N_49424,N_45842);
nand UO_1968 (O_1968,N_45497,N_47937);
and UO_1969 (O_1969,N_46980,N_49455);
and UO_1970 (O_1970,N_47289,N_46123);
xnor UO_1971 (O_1971,N_49131,N_45594);
or UO_1972 (O_1972,N_47816,N_46367);
and UO_1973 (O_1973,N_49649,N_48932);
xnor UO_1974 (O_1974,N_48014,N_48282);
and UO_1975 (O_1975,N_45536,N_47018);
and UO_1976 (O_1976,N_48409,N_45455);
nor UO_1977 (O_1977,N_45793,N_46250);
and UO_1978 (O_1978,N_47766,N_45935);
and UO_1979 (O_1979,N_48167,N_47548);
or UO_1980 (O_1980,N_46312,N_47199);
nand UO_1981 (O_1981,N_47762,N_46191);
nand UO_1982 (O_1982,N_47915,N_49036);
and UO_1983 (O_1983,N_47355,N_45104);
and UO_1984 (O_1984,N_49469,N_45475);
or UO_1985 (O_1985,N_49533,N_49492);
and UO_1986 (O_1986,N_49437,N_48967);
and UO_1987 (O_1987,N_45024,N_49604);
and UO_1988 (O_1988,N_49029,N_49917);
xor UO_1989 (O_1989,N_45992,N_45584);
nand UO_1990 (O_1990,N_48351,N_48343);
nand UO_1991 (O_1991,N_47784,N_48573);
nand UO_1992 (O_1992,N_49456,N_48904);
nand UO_1993 (O_1993,N_45311,N_46233);
nand UO_1994 (O_1994,N_49427,N_49642);
xor UO_1995 (O_1995,N_45683,N_47588);
or UO_1996 (O_1996,N_48319,N_46180);
or UO_1997 (O_1997,N_46793,N_49371);
xor UO_1998 (O_1998,N_48025,N_49154);
xnor UO_1999 (O_1999,N_48455,N_49377);
nor UO_2000 (O_2000,N_45789,N_46643);
nor UO_2001 (O_2001,N_49397,N_46383);
nor UO_2002 (O_2002,N_47054,N_46273);
or UO_2003 (O_2003,N_46309,N_46334);
and UO_2004 (O_2004,N_45218,N_48125);
xnor UO_2005 (O_2005,N_48873,N_46936);
nand UO_2006 (O_2006,N_46377,N_48232);
nor UO_2007 (O_2007,N_49908,N_45351);
and UO_2008 (O_2008,N_49688,N_45013);
or UO_2009 (O_2009,N_46333,N_49566);
and UO_2010 (O_2010,N_47656,N_48542);
and UO_2011 (O_2011,N_49743,N_47140);
xor UO_2012 (O_2012,N_49782,N_45711);
xor UO_2013 (O_2013,N_47257,N_49713);
and UO_2014 (O_2014,N_46861,N_45082);
nand UO_2015 (O_2015,N_48162,N_49929);
and UO_2016 (O_2016,N_48044,N_48368);
nor UO_2017 (O_2017,N_47245,N_47357);
nand UO_2018 (O_2018,N_45696,N_49640);
xnor UO_2019 (O_2019,N_45830,N_46915);
nor UO_2020 (O_2020,N_45898,N_47051);
or UO_2021 (O_2021,N_49568,N_49804);
nand UO_2022 (O_2022,N_47949,N_49191);
and UO_2023 (O_2023,N_45154,N_46841);
nand UO_2024 (O_2024,N_46744,N_47029);
nor UO_2025 (O_2025,N_47241,N_49267);
nand UO_2026 (O_2026,N_48347,N_48657);
or UO_2027 (O_2027,N_45362,N_47105);
xnor UO_2028 (O_2028,N_48144,N_45851);
nor UO_2029 (O_2029,N_49050,N_49776);
nand UO_2030 (O_2030,N_47356,N_45890);
nor UO_2031 (O_2031,N_47675,N_48149);
xor UO_2032 (O_2032,N_47098,N_49329);
and UO_2033 (O_2033,N_47127,N_48768);
or UO_2034 (O_2034,N_45369,N_49941);
nor UO_2035 (O_2035,N_49498,N_46589);
and UO_2036 (O_2036,N_45274,N_45917);
or UO_2037 (O_2037,N_45605,N_49184);
nand UO_2038 (O_2038,N_47881,N_47252);
xor UO_2039 (O_2039,N_46185,N_45607);
xor UO_2040 (O_2040,N_46043,N_46107);
and UO_2041 (O_2041,N_45534,N_49656);
nor UO_2042 (O_2042,N_48750,N_47924);
nand UO_2043 (O_2043,N_47524,N_48260);
xor UO_2044 (O_2044,N_49761,N_45858);
xnor UO_2045 (O_2045,N_47648,N_48259);
and UO_2046 (O_2046,N_45447,N_45477);
nand UO_2047 (O_2047,N_45440,N_49654);
nand UO_2048 (O_2048,N_47535,N_48336);
xnor UO_2049 (O_2049,N_46895,N_49011);
nor UO_2050 (O_2050,N_45258,N_49119);
or UO_2051 (O_2051,N_48899,N_46479);
nand UO_2052 (O_2052,N_47869,N_48546);
nand UO_2053 (O_2053,N_45795,N_46585);
and UO_2054 (O_2054,N_47946,N_48291);
and UO_2055 (O_2055,N_46256,N_45955);
and UO_2056 (O_2056,N_46000,N_48209);
xor UO_2057 (O_2057,N_48632,N_49994);
nor UO_2058 (O_2058,N_47474,N_47244);
or UO_2059 (O_2059,N_49093,N_46132);
and UO_2060 (O_2060,N_46869,N_49793);
and UO_2061 (O_2061,N_49074,N_48078);
or UO_2062 (O_2062,N_49251,N_49166);
and UO_2063 (O_2063,N_48346,N_47012);
nor UO_2064 (O_2064,N_45204,N_47594);
and UO_2065 (O_2065,N_47308,N_46451);
or UO_2066 (O_2066,N_48762,N_47388);
xor UO_2067 (O_2067,N_49073,N_46075);
nor UO_2068 (O_2068,N_45226,N_48520);
or UO_2069 (O_2069,N_45612,N_47863);
nand UO_2070 (O_2070,N_46552,N_45945);
xnor UO_2071 (O_2071,N_48211,N_47039);
or UO_2072 (O_2072,N_48395,N_45939);
and UO_2073 (O_2073,N_48118,N_46783);
nor UO_2074 (O_2074,N_47531,N_48085);
xnor UO_2075 (O_2075,N_49149,N_49689);
nor UO_2076 (O_2076,N_49313,N_45925);
or UO_2077 (O_2077,N_47805,N_49128);
nand UO_2078 (O_2078,N_47972,N_46146);
or UO_2079 (O_2079,N_46001,N_47121);
nor UO_2080 (O_2080,N_46892,N_47171);
nor UO_2081 (O_2081,N_48707,N_49495);
and UO_2082 (O_2082,N_47970,N_49910);
nand UO_2083 (O_2083,N_47239,N_45677);
nand UO_2084 (O_2084,N_49109,N_47031);
nand UO_2085 (O_2085,N_47801,N_47432);
nor UO_2086 (O_2086,N_48961,N_47198);
nor UO_2087 (O_2087,N_46919,N_48101);
nand UO_2088 (O_2088,N_45761,N_49231);
nor UO_2089 (O_2089,N_48513,N_45259);
nor UO_2090 (O_2090,N_47066,N_47847);
or UO_2091 (O_2091,N_46229,N_46976);
and UO_2092 (O_2092,N_48062,N_46169);
and UO_2093 (O_2093,N_47631,N_47636);
or UO_2094 (O_2094,N_45934,N_48269);
xnor UO_2095 (O_2095,N_49326,N_47112);
and UO_2096 (O_2096,N_48857,N_48647);
or UO_2097 (O_2097,N_49666,N_46855);
and UO_2098 (O_2098,N_47382,N_48594);
nor UO_2099 (O_2099,N_45544,N_49555);
nor UO_2100 (O_2100,N_48681,N_47461);
or UO_2101 (O_2101,N_47180,N_49233);
or UO_2102 (O_2102,N_48510,N_48833);
nand UO_2103 (O_2103,N_46662,N_48217);
or UO_2104 (O_2104,N_49464,N_48976);
and UO_2105 (O_2105,N_49752,N_48706);
nand UO_2106 (O_2106,N_46658,N_48786);
or UO_2107 (O_2107,N_46137,N_46217);
nand UO_2108 (O_2108,N_46732,N_46343);
nand UO_2109 (O_2109,N_48749,N_45317);
or UO_2110 (O_2110,N_45942,N_47033);
and UO_2111 (O_2111,N_45532,N_47107);
nand UO_2112 (O_2112,N_49208,N_47103);
or UO_2113 (O_2113,N_45662,N_46428);
xnor UO_2114 (O_2114,N_48486,N_49652);
xor UO_2115 (O_2115,N_45430,N_48960);
nand UO_2116 (O_2116,N_47810,N_45569);
and UO_2117 (O_2117,N_47327,N_46409);
nand UO_2118 (O_2118,N_48561,N_47161);
xor UO_2119 (O_2119,N_49507,N_45845);
nor UO_2120 (O_2120,N_45081,N_47016);
xor UO_2121 (O_2121,N_49746,N_46085);
and UO_2122 (O_2122,N_48249,N_45566);
or UO_2123 (O_2123,N_45156,N_47714);
and UO_2124 (O_2124,N_47084,N_47274);
xor UO_2125 (O_2125,N_46902,N_46432);
nand UO_2126 (O_2126,N_45687,N_49532);
or UO_2127 (O_2127,N_49376,N_48387);
xor UO_2128 (O_2128,N_48672,N_47649);
and UO_2129 (O_2129,N_49799,N_49506);
and UO_2130 (O_2130,N_47760,N_48180);
nand UO_2131 (O_2131,N_46142,N_48441);
xor UO_2132 (O_2132,N_47179,N_48810);
nand UO_2133 (O_2133,N_48702,N_48035);
nand UO_2134 (O_2134,N_49246,N_45572);
and UO_2135 (O_2135,N_45213,N_46648);
nor UO_2136 (O_2136,N_46471,N_45548);
and UO_2137 (O_2137,N_47622,N_46300);
nand UO_2138 (O_2138,N_47534,N_48884);
or UO_2139 (O_2139,N_46512,N_46242);
or UO_2140 (O_2140,N_46181,N_47427);
nor UO_2141 (O_2141,N_49091,N_48429);
nand UO_2142 (O_2142,N_47740,N_46880);
nand UO_2143 (O_2143,N_48210,N_48046);
or UO_2144 (O_2144,N_47617,N_45042);
nand UO_2145 (O_2145,N_45538,N_45837);
xor UO_2146 (O_2146,N_48164,N_49886);
xnor UO_2147 (O_2147,N_49365,N_49304);
nor UO_2148 (O_2148,N_47123,N_48654);
and UO_2149 (O_2149,N_48846,N_48638);
nand UO_2150 (O_2150,N_48009,N_45717);
or UO_2151 (O_2151,N_48155,N_45539);
xnor UO_2152 (O_2152,N_49317,N_47982);
or UO_2153 (O_2153,N_47317,N_49900);
or UO_2154 (O_2154,N_45675,N_48716);
nand UO_2155 (O_2155,N_46360,N_48676);
xor UO_2156 (O_2156,N_48578,N_45782);
nor UO_2157 (O_2157,N_46676,N_46604);
nor UO_2158 (O_2158,N_48738,N_46239);
nand UO_2159 (O_2159,N_46226,N_49513);
and UO_2160 (O_2160,N_48725,N_47311);
nand UO_2161 (O_2161,N_46005,N_46590);
nor UO_2162 (O_2162,N_49472,N_48463);
and UO_2163 (O_2163,N_46568,N_47210);
xnor UO_2164 (O_2164,N_46292,N_49324);
and UO_2165 (O_2165,N_45306,N_46912);
or UO_2166 (O_2166,N_45403,N_46699);
nand UO_2167 (O_2167,N_46113,N_48204);
xor UO_2168 (O_2168,N_47780,N_48673);
nand UO_2169 (O_2169,N_45573,N_48124);
nand UO_2170 (O_2170,N_48364,N_47547);
or UO_2171 (O_2171,N_45737,N_45948);
nor UO_2172 (O_2172,N_49162,N_46157);
or UO_2173 (O_2173,N_46842,N_46733);
nor UO_2174 (O_2174,N_48182,N_45237);
xor UO_2175 (O_2175,N_45541,N_45190);
and UO_2176 (O_2176,N_47964,N_48655);
xnor UO_2177 (O_2177,N_46329,N_47189);
nor UO_2178 (O_2178,N_49295,N_49003);
and UO_2179 (O_2179,N_49122,N_46559);
or UO_2180 (O_2180,N_49132,N_49250);
nor UO_2181 (O_2181,N_46010,N_48504);
and UO_2182 (O_2182,N_46091,N_45348);
xor UO_2183 (O_2183,N_48495,N_46139);
and UO_2184 (O_2184,N_47046,N_47597);
or UO_2185 (O_2185,N_46951,N_45786);
nor UO_2186 (O_2186,N_45695,N_49725);
and UO_2187 (O_2187,N_45145,N_48199);
nor UO_2188 (O_2188,N_48229,N_47270);
nand UO_2189 (O_2189,N_46225,N_49386);
nor UO_2190 (O_2190,N_45730,N_49098);
and UO_2191 (O_2191,N_47399,N_48596);
nand UO_2192 (O_2192,N_47540,N_48859);
nor UO_2193 (O_2193,N_49283,N_45412);
or UO_2194 (O_2194,N_46663,N_48831);
nor UO_2195 (O_2195,N_47761,N_45632);
nor UO_2196 (O_2196,N_46291,N_47472);
xor UO_2197 (O_2197,N_46020,N_46230);
xor UO_2198 (O_2198,N_49834,N_48238);
or UO_2199 (O_2199,N_45674,N_45321);
xnor UO_2200 (O_2200,N_46337,N_47519);
and UO_2201 (O_2201,N_47495,N_48131);
nor UO_2202 (O_2202,N_48173,N_48793);
xor UO_2203 (O_2203,N_45854,N_47369);
xnor UO_2204 (O_2204,N_46497,N_49165);
nor UO_2205 (O_2205,N_45133,N_48021);
or UO_2206 (O_2206,N_46519,N_49895);
xor UO_2207 (O_2207,N_45810,N_49186);
xor UO_2208 (O_2208,N_47363,N_47562);
and UO_2209 (O_2209,N_49423,N_49739);
nor UO_2210 (O_2210,N_46704,N_49526);
nand UO_2211 (O_2211,N_49897,N_49258);
nand UO_2212 (O_2212,N_46339,N_45198);
and UO_2213 (O_2213,N_45790,N_47237);
nor UO_2214 (O_2214,N_45320,N_46076);
and UO_2215 (O_2215,N_47259,N_49196);
nand UO_2216 (O_2216,N_46095,N_45290);
nand UO_2217 (O_2217,N_49738,N_47603);
nand UO_2218 (O_2218,N_47487,N_48266);
and UO_2219 (O_2219,N_46498,N_46326);
or UO_2220 (O_2220,N_46785,N_45228);
nor UO_2221 (O_2221,N_47897,N_45876);
nand UO_2222 (O_2222,N_48697,N_47549);
or UO_2223 (O_2223,N_46112,N_47712);
or UO_2224 (O_2224,N_49436,N_46460);
or UO_2225 (O_2225,N_45030,N_45338);
nor UO_2226 (O_2226,N_49148,N_49069);
and UO_2227 (O_2227,N_46656,N_47286);
and UO_2228 (O_2228,N_47146,N_48008);
xor UO_2229 (O_2229,N_46940,N_48532);
nand UO_2230 (O_2230,N_48033,N_45231);
and UO_2231 (O_2231,N_47777,N_49926);
xor UO_2232 (O_2232,N_48895,N_46909);
nand UO_2233 (O_2233,N_46247,N_47821);
nor UO_2234 (O_2234,N_46209,N_48200);
nand UO_2235 (O_2235,N_47110,N_46138);
nor UO_2236 (O_2236,N_47736,N_48661);
nand UO_2237 (O_2237,N_49629,N_48003);
and UO_2238 (O_2238,N_45609,N_46509);
xor UO_2239 (O_2239,N_47144,N_45186);
nand UO_2240 (O_2240,N_49446,N_46613);
or UO_2241 (O_2241,N_47233,N_46294);
xor UO_2242 (O_2242,N_49380,N_49240);
nand UO_2243 (O_2243,N_48255,N_49563);
or UO_2244 (O_2244,N_46024,N_46200);
nand UO_2245 (O_2245,N_49745,N_48045);
nor UO_2246 (O_2246,N_48952,N_45829);
xnor UO_2247 (O_2247,N_48953,N_46975);
or UO_2248 (O_2248,N_47963,N_45456);
or UO_2249 (O_2249,N_48457,N_48426);
nor UO_2250 (O_2250,N_45563,N_47424);
nor UO_2251 (O_2251,N_49081,N_46572);
and UO_2252 (O_2252,N_49321,N_47203);
nor UO_2253 (O_2253,N_49028,N_46586);
nand UO_2254 (O_2254,N_47475,N_48252);
nor UO_2255 (O_2255,N_46070,N_48369);
or UO_2256 (O_2256,N_46979,N_47521);
and UO_2257 (O_2257,N_45480,N_47751);
nand UO_2258 (O_2258,N_49881,N_47868);
and UO_2259 (O_2259,N_45908,N_45953);
nand UO_2260 (O_2260,N_47542,N_48154);
or UO_2261 (O_2261,N_46614,N_48471);
and UO_2262 (O_2262,N_46435,N_45144);
nor UO_2263 (O_2263,N_45142,N_47209);
nor UO_2264 (O_2264,N_47530,N_46558);
or UO_2265 (O_2265,N_45811,N_45028);
and UO_2266 (O_2266,N_48052,N_46774);
xnor UO_2267 (O_2267,N_45748,N_46609);
and UO_2268 (O_2268,N_49403,N_48373);
and UO_2269 (O_2269,N_49866,N_45929);
and UO_2270 (O_2270,N_47093,N_46039);
or UO_2271 (O_2271,N_48038,N_48466);
nand UO_2272 (O_2272,N_47808,N_46508);
xor UO_2273 (O_2273,N_47223,N_49703);
nor UO_2274 (O_2274,N_47682,N_46164);
nor UO_2275 (O_2275,N_47436,N_46749);
xnor UO_2276 (O_2276,N_45770,N_47838);
and UO_2277 (O_2277,N_48402,N_46501);
nor UO_2278 (O_2278,N_48593,N_46313);
nand UO_2279 (O_2279,N_48732,N_46937);
and UO_2280 (O_2280,N_48825,N_49552);
and UO_2281 (O_2281,N_45806,N_47710);
or UO_2282 (O_2282,N_47272,N_47739);
or UO_2283 (O_2283,N_45423,N_49690);
and UO_2284 (O_2284,N_45656,N_45905);
nor UO_2285 (O_2285,N_47411,N_49143);
xnor UO_2286 (O_2286,N_46193,N_45469);
and UO_2287 (O_2287,N_46705,N_47072);
xnor UO_2288 (O_2288,N_45188,N_49964);
nor UO_2289 (O_2289,N_45668,N_46240);
nor UO_2290 (O_2290,N_49193,N_46819);
and UO_2291 (O_2291,N_45729,N_46910);
xor UO_2292 (O_2292,N_47754,N_49232);
xnor UO_2293 (O_2293,N_49968,N_47013);
nor UO_2294 (O_2294,N_47768,N_49647);
nor UO_2295 (O_2295,N_49207,N_46310);
or UO_2296 (O_2296,N_45343,N_47068);
xor UO_2297 (O_2297,N_49932,N_46677);
nor UO_2298 (O_2298,N_47350,N_48283);
and UO_2299 (O_2299,N_49798,N_46925);
nor UO_2300 (O_2300,N_49438,N_48142);
or UO_2301 (O_2301,N_48851,N_45773);
or UO_2302 (O_2302,N_46237,N_47758);
or UO_2303 (O_2303,N_48079,N_46036);
and UO_2304 (O_2304,N_49867,N_48837);
or UO_2305 (O_2305,N_47912,N_47192);
or UO_2306 (O_2306,N_47556,N_48489);
xnor UO_2307 (O_2307,N_46317,N_48622);
nor UO_2308 (O_2308,N_46570,N_49107);
and UO_2309 (O_2309,N_45977,N_47154);
nor UO_2310 (O_2310,N_48587,N_48089);
or UO_2311 (O_2311,N_47042,N_45586);
nand UO_2312 (O_2312,N_49548,N_46093);
nand UO_2313 (O_2313,N_46554,N_46280);
or UO_2314 (O_2314,N_47301,N_45131);
or UO_2315 (O_2315,N_49272,N_49704);
xor UO_2316 (O_2316,N_47772,N_47122);
nand UO_2317 (O_2317,N_47108,N_48436);
or UO_2318 (O_2318,N_48843,N_46363);
nand UO_2319 (O_2319,N_46626,N_46661);
or UO_2320 (O_2320,N_47560,N_49300);
xor UO_2321 (O_2321,N_49734,N_48914);
nor UO_2322 (O_2322,N_46324,N_47275);
and UO_2323 (O_2323,N_49341,N_48341);
or UO_2324 (O_2324,N_45248,N_48909);
nor UO_2325 (O_2325,N_45146,N_48458);
nor UO_2326 (O_2326,N_47966,N_46615);
nor UO_2327 (O_2327,N_47492,N_47716);
xor UO_2328 (O_2328,N_47859,N_48309);
nand UO_2329 (O_2329,N_48242,N_46964);
and UO_2330 (O_2330,N_49284,N_45305);
and UO_2331 (O_2331,N_48397,N_48137);
nand UO_2332 (O_2332,N_47511,N_46518);
and UO_2333 (O_2333,N_49330,N_45636);
xor UO_2334 (O_2334,N_45149,N_46911);
or UO_2335 (O_2335,N_46603,N_45152);
or UO_2336 (O_2336,N_48219,N_46199);
or UO_2337 (O_2337,N_48642,N_47983);
xor UO_2338 (O_2338,N_47229,N_48271);
nand UO_2339 (O_2339,N_45721,N_48088);
and UO_2340 (O_2340,N_49303,N_46866);
nand UO_2341 (O_2341,N_47923,N_49684);
xor UO_2342 (O_2342,N_46415,N_47362);
or UO_2343 (O_2343,N_47027,N_45010);
nand UO_2344 (O_2344,N_45868,N_49644);
and UO_2345 (O_2345,N_46464,N_45164);
xor UO_2346 (O_2346,N_47433,N_49669);
xor UO_2347 (O_2347,N_49180,N_45389);
and UO_2348 (O_2348,N_49359,N_49998);
nand UO_2349 (O_2349,N_45615,N_48461);
or UO_2350 (O_2350,N_47412,N_46296);
nor UO_2351 (O_2351,N_45578,N_48589);
or UO_2352 (O_2352,N_48063,N_47935);
nand UO_2353 (O_2353,N_45753,N_48643);
nand UO_2354 (O_2354,N_49626,N_46578);
xor UO_2355 (O_2355,N_45518,N_48064);
nor UO_2356 (O_2356,N_48572,N_46206);
xor UO_2357 (O_2357,N_48704,N_47392);
or UO_2358 (O_2358,N_47376,N_48261);
or UO_2359 (O_2359,N_48029,N_48095);
nor UO_2360 (O_2360,N_48475,N_48296);
xor UO_2361 (O_2361,N_47402,N_47375);
and UO_2362 (O_2362,N_47918,N_45364);
and UO_2363 (O_2363,N_49785,N_46683);
or UO_2364 (O_2364,N_47010,N_46986);
or UO_2365 (O_2365,N_45601,N_45661);
nand UO_2366 (O_2366,N_49823,N_49827);
or UO_2367 (O_2367,N_49100,N_47439);
or UO_2368 (O_2368,N_46551,N_46901);
nand UO_2369 (O_2369,N_48625,N_45884);
nand UO_2370 (O_2370,N_48472,N_46918);
or UO_2371 (O_2371,N_45846,N_47895);
xor UO_2372 (O_2372,N_47097,N_49610);
nand UO_2373 (O_2373,N_47662,N_45521);
nor UO_2374 (O_2374,N_48660,N_48549);
nand UO_2375 (O_2375,N_49302,N_45243);
or UO_2376 (O_2376,N_48933,N_47340);
xor UO_2377 (O_2377,N_47221,N_48396);
and UO_2378 (O_2378,N_49407,N_46196);
nand UO_2379 (O_2379,N_48954,N_45581);
nor UO_2380 (O_2380,N_45130,N_47874);
xor UO_2381 (O_2381,N_45700,N_46021);
and UO_2382 (O_2382,N_49890,N_46149);
and UO_2383 (O_2383,N_46516,N_49443);
xor UO_2384 (O_2384,N_48821,N_46156);
or UO_2385 (O_2385,N_49367,N_49832);
and UO_2386 (O_2386,N_45344,N_48377);
or UO_2387 (O_2387,N_46702,N_48905);
nor UO_2388 (O_2388,N_47702,N_46750);
and UO_2389 (O_2389,N_49662,N_46695);
nor UO_2390 (O_2390,N_48141,N_49089);
xnor UO_2391 (O_2391,N_49682,N_45798);
nor UO_2392 (O_2392,N_46649,N_45881);
xor UO_2393 (O_2393,N_47894,N_47444);
xnor UO_2394 (O_2394,N_47053,N_49416);
nand UO_2395 (O_2395,N_47822,N_45481);
xnor UO_2396 (O_2396,N_47137,N_47723);
or UO_2397 (O_2397,N_48193,N_48547);
xor UO_2398 (O_2398,N_49596,N_46970);
or UO_2399 (O_2399,N_48653,N_48640);
or UO_2400 (O_2400,N_46672,N_48497);
xor UO_2401 (O_2401,N_45184,N_46760);
xnor UO_2402 (O_2402,N_45997,N_45844);
xor UO_2403 (O_2403,N_47490,N_47864);
nor UO_2404 (O_2404,N_49990,N_48236);
and UO_2405 (O_2405,N_47187,N_46562);
xnor UO_2406 (O_2406,N_47797,N_46838);
or UO_2407 (O_2407,N_48701,N_49287);
or UO_2408 (O_2408,N_45552,N_47564);
or UO_2409 (O_2409,N_45381,N_48376);
nand UO_2410 (O_2410,N_46330,N_49847);
xnor UO_2411 (O_2411,N_46954,N_48664);
and UO_2412 (O_2412,N_49868,N_48418);
nand UO_2413 (O_2413,N_49198,N_49138);
xnor UO_2414 (O_2414,N_48084,N_49458);
or UO_2415 (O_2415,N_46511,N_47681);
nand UO_2416 (O_2416,N_45498,N_49474);
nand UO_2417 (O_2417,N_45494,N_49921);
and UO_2418 (O_2418,N_46757,N_47566);
or UO_2419 (O_2419,N_46600,N_45201);
nor UO_2420 (O_2420,N_49820,N_45621);
or UO_2421 (O_2421,N_45002,N_47651);
or UO_2422 (O_2422,N_49899,N_48816);
xor UO_2423 (O_2423,N_46457,N_49633);
or UO_2424 (O_2424,N_45543,N_49201);
nand UO_2425 (O_2425,N_47139,N_45546);
or UO_2426 (O_2426,N_48912,N_47967);
nand UO_2427 (O_2427,N_45856,N_46743);
and UO_2428 (O_2428,N_45160,N_48433);
nor UO_2429 (O_2429,N_49400,N_48354);
xor UO_2430 (O_2430,N_49369,N_45460);
nand UO_2431 (O_2431,N_45653,N_47959);
xnor UO_2432 (O_2432,N_45604,N_49668);
nand UO_2433 (O_2433,N_48565,N_47273);
or UO_2434 (O_2434,N_45257,N_45760);
xnor UO_2435 (O_2435,N_45901,N_47222);
nand UO_2436 (O_2436,N_49835,N_49126);
nand UO_2437 (O_2437,N_48093,N_45223);
nand UO_2438 (O_2438,N_46099,N_45508);
or UO_2439 (O_2439,N_49925,N_46017);
or UO_2440 (O_2440,N_45261,N_46030);
nand UO_2441 (O_2441,N_45200,N_45075);
and UO_2442 (O_2442,N_45000,N_47509);
nor UO_2443 (O_2443,N_49461,N_49711);
or UO_2444 (O_2444,N_48695,N_49178);
or UO_2445 (O_2445,N_49216,N_46014);
and UO_2446 (O_2446,N_45039,N_48104);
and UO_2447 (O_2447,N_46483,N_49289);
xnor UO_2448 (O_2448,N_45241,N_49980);
or UO_2449 (O_2449,N_48036,N_48450);
nor UO_2450 (O_2450,N_49301,N_47654);
nand UO_2451 (O_2451,N_47453,N_47083);
or UO_2452 (O_2452,N_47044,N_46631);
nor UO_2453 (O_2453,N_45124,N_48945);
and UO_2454 (O_2454,N_48678,N_47828);
nor UO_2455 (O_2455,N_46530,N_47779);
and UO_2456 (O_2456,N_48715,N_48682);
or UO_2457 (O_2457,N_49988,N_49714);
xor UO_2458 (O_2458,N_48077,N_47269);
or UO_2459 (O_2459,N_47383,N_48662);
nor UO_2460 (O_2460,N_45875,N_45316);
and UO_2461 (O_2461,N_48477,N_46854);
and UO_2462 (O_2462,N_48379,N_47422);
nor UO_2463 (O_2463,N_47364,N_46499);
nand UO_2464 (O_2464,N_45016,N_46458);
nor UO_2465 (O_2465,N_46633,N_49950);
nand UO_2466 (O_2466,N_48322,N_47294);
nand UO_2467 (O_2467,N_47941,N_48607);
xnor UO_2468 (O_2468,N_45384,N_48190);
and UO_2469 (O_2469,N_48110,N_46177);
xor UO_2470 (O_2470,N_48553,N_45353);
nor UO_2471 (O_2471,N_45315,N_46746);
nor UO_2472 (O_2472,N_48631,N_46994);
or UO_2473 (O_2473,N_48990,N_49562);
nor UO_2474 (O_2474,N_49421,N_47943);
and UO_2475 (O_2475,N_46908,N_47853);
and UO_2476 (O_2476,N_47873,N_46058);
and UO_2477 (O_2477,N_47096,N_47958);
nand UO_2478 (O_2478,N_48942,N_48832);
or UO_2479 (O_2479,N_49323,N_46365);
xor UO_2480 (O_2480,N_45702,N_48650);
xor UO_2481 (O_2481,N_48743,N_46882);
nor UO_2482 (O_2482,N_49625,N_45108);
nand UO_2483 (O_2483,N_47113,N_46266);
nor UO_2484 (O_2484,N_45012,N_48448);
xor UO_2485 (O_2485,N_45545,N_48384);
or UO_2486 (O_2486,N_49521,N_47627);
and UO_2487 (O_2487,N_46817,N_48065);
xor UO_2488 (O_2488,N_45326,N_49234);
or UO_2489 (O_2489,N_46725,N_46490);
or UO_2490 (O_2490,N_47445,N_49962);
nor UO_2491 (O_2491,N_48926,N_45853);
nand UO_2492 (O_2492,N_48328,N_48299);
or UO_2493 (O_2493,N_46090,N_45803);
nand UO_2494 (O_2494,N_45506,N_46706);
nand UO_2495 (O_2495,N_49757,N_47420);
or UO_2496 (O_2496,N_47043,N_47057);
and UO_2497 (O_2497,N_46323,N_48424);
and UO_2498 (O_2498,N_46837,N_47769);
nor UO_2499 (O_2499,N_45172,N_47319);
nand UO_2500 (O_2500,N_47715,N_46785);
nand UO_2501 (O_2501,N_46240,N_46652);
nand UO_2502 (O_2502,N_49364,N_46204);
and UO_2503 (O_2503,N_45094,N_49632);
xnor UO_2504 (O_2504,N_49461,N_48796);
nand UO_2505 (O_2505,N_45309,N_47618);
or UO_2506 (O_2506,N_49143,N_45101);
and UO_2507 (O_2507,N_46888,N_48698);
and UO_2508 (O_2508,N_48553,N_46917);
and UO_2509 (O_2509,N_47750,N_46192);
nand UO_2510 (O_2510,N_45594,N_49111);
or UO_2511 (O_2511,N_45092,N_45242);
xor UO_2512 (O_2512,N_48962,N_47941);
xor UO_2513 (O_2513,N_46543,N_46027);
and UO_2514 (O_2514,N_49936,N_46822);
or UO_2515 (O_2515,N_46579,N_47023);
nor UO_2516 (O_2516,N_48999,N_47759);
and UO_2517 (O_2517,N_49278,N_46511);
or UO_2518 (O_2518,N_47217,N_49951);
or UO_2519 (O_2519,N_49422,N_46645);
and UO_2520 (O_2520,N_46504,N_47650);
nand UO_2521 (O_2521,N_49384,N_45664);
xor UO_2522 (O_2522,N_48489,N_46488);
or UO_2523 (O_2523,N_45746,N_46194);
xnor UO_2524 (O_2524,N_48636,N_45140);
or UO_2525 (O_2525,N_49232,N_47462);
and UO_2526 (O_2526,N_48129,N_46562);
nand UO_2527 (O_2527,N_47966,N_48026);
or UO_2528 (O_2528,N_49443,N_45488);
nor UO_2529 (O_2529,N_46235,N_48967);
nor UO_2530 (O_2530,N_47810,N_49489);
and UO_2531 (O_2531,N_46564,N_48385);
xnor UO_2532 (O_2532,N_45796,N_47938);
nand UO_2533 (O_2533,N_49042,N_48215);
nor UO_2534 (O_2534,N_48243,N_46534);
nand UO_2535 (O_2535,N_45112,N_48819);
or UO_2536 (O_2536,N_47294,N_45701);
or UO_2537 (O_2537,N_48735,N_48750);
xnor UO_2538 (O_2538,N_46765,N_47399);
and UO_2539 (O_2539,N_48556,N_45741);
nor UO_2540 (O_2540,N_45826,N_48603);
nor UO_2541 (O_2541,N_46570,N_48414);
nand UO_2542 (O_2542,N_46437,N_46530);
xnor UO_2543 (O_2543,N_47110,N_45504);
and UO_2544 (O_2544,N_48116,N_49198);
and UO_2545 (O_2545,N_49129,N_49740);
or UO_2546 (O_2546,N_45994,N_45557);
xnor UO_2547 (O_2547,N_45958,N_49191);
nand UO_2548 (O_2548,N_46072,N_45578);
or UO_2549 (O_2549,N_46988,N_47968);
nand UO_2550 (O_2550,N_47468,N_45737);
or UO_2551 (O_2551,N_48147,N_45189);
xnor UO_2552 (O_2552,N_48877,N_49987);
or UO_2553 (O_2553,N_48708,N_45007);
or UO_2554 (O_2554,N_45329,N_46064);
nor UO_2555 (O_2555,N_45674,N_47077);
nor UO_2556 (O_2556,N_48273,N_46511);
nand UO_2557 (O_2557,N_47944,N_49485);
nand UO_2558 (O_2558,N_45351,N_47697);
nor UO_2559 (O_2559,N_49593,N_46477);
nor UO_2560 (O_2560,N_48721,N_46641);
xor UO_2561 (O_2561,N_46577,N_48762);
or UO_2562 (O_2562,N_47088,N_47753);
xor UO_2563 (O_2563,N_48082,N_48758);
or UO_2564 (O_2564,N_46337,N_46421);
nor UO_2565 (O_2565,N_45380,N_46707);
and UO_2566 (O_2566,N_48876,N_48581);
nand UO_2567 (O_2567,N_46672,N_46009);
and UO_2568 (O_2568,N_48377,N_49903);
xor UO_2569 (O_2569,N_47356,N_49791);
or UO_2570 (O_2570,N_45258,N_46328);
xnor UO_2571 (O_2571,N_45709,N_46050);
and UO_2572 (O_2572,N_49344,N_49035);
nand UO_2573 (O_2573,N_46643,N_45098);
or UO_2574 (O_2574,N_47757,N_47099);
xor UO_2575 (O_2575,N_45922,N_46232);
xor UO_2576 (O_2576,N_47101,N_46045);
xor UO_2577 (O_2577,N_46197,N_47758);
nand UO_2578 (O_2578,N_46630,N_45797);
nor UO_2579 (O_2579,N_48152,N_47762);
xor UO_2580 (O_2580,N_45100,N_48793);
or UO_2581 (O_2581,N_48066,N_46788);
and UO_2582 (O_2582,N_46917,N_48213);
and UO_2583 (O_2583,N_49254,N_49067);
xnor UO_2584 (O_2584,N_45476,N_47070);
nor UO_2585 (O_2585,N_45071,N_48164);
and UO_2586 (O_2586,N_49254,N_45881);
nand UO_2587 (O_2587,N_47270,N_46216);
and UO_2588 (O_2588,N_45063,N_47262);
nor UO_2589 (O_2589,N_45769,N_48493);
nand UO_2590 (O_2590,N_48870,N_47679);
and UO_2591 (O_2591,N_46858,N_49832);
nor UO_2592 (O_2592,N_47268,N_48048);
or UO_2593 (O_2593,N_49944,N_49642);
xnor UO_2594 (O_2594,N_47312,N_48130);
nand UO_2595 (O_2595,N_45384,N_48891);
nor UO_2596 (O_2596,N_46484,N_48710);
and UO_2597 (O_2597,N_49737,N_45551);
nand UO_2598 (O_2598,N_46152,N_45187);
nand UO_2599 (O_2599,N_48891,N_47075);
and UO_2600 (O_2600,N_45619,N_49148);
nand UO_2601 (O_2601,N_45260,N_47268);
or UO_2602 (O_2602,N_48733,N_47747);
or UO_2603 (O_2603,N_47048,N_47614);
and UO_2604 (O_2604,N_45080,N_45425);
or UO_2605 (O_2605,N_45409,N_49434);
or UO_2606 (O_2606,N_49549,N_46776);
and UO_2607 (O_2607,N_46398,N_48041);
nand UO_2608 (O_2608,N_49523,N_49572);
nand UO_2609 (O_2609,N_48464,N_48614);
xnor UO_2610 (O_2610,N_48423,N_48322);
nand UO_2611 (O_2611,N_46877,N_45060);
or UO_2612 (O_2612,N_47934,N_46295);
nand UO_2613 (O_2613,N_49202,N_48305);
or UO_2614 (O_2614,N_45060,N_48864);
nor UO_2615 (O_2615,N_45752,N_48797);
nor UO_2616 (O_2616,N_49484,N_49206);
nor UO_2617 (O_2617,N_49354,N_46927);
nor UO_2618 (O_2618,N_48907,N_45787);
nand UO_2619 (O_2619,N_49639,N_49745);
nor UO_2620 (O_2620,N_46832,N_46513);
nor UO_2621 (O_2621,N_45414,N_46253);
nor UO_2622 (O_2622,N_46581,N_47739);
and UO_2623 (O_2623,N_47048,N_47224);
nand UO_2624 (O_2624,N_49542,N_47683);
xor UO_2625 (O_2625,N_45697,N_48122);
and UO_2626 (O_2626,N_48101,N_46007);
or UO_2627 (O_2627,N_46804,N_47981);
and UO_2628 (O_2628,N_48816,N_48721);
nor UO_2629 (O_2629,N_46159,N_47165);
or UO_2630 (O_2630,N_46971,N_48961);
and UO_2631 (O_2631,N_45238,N_47255);
or UO_2632 (O_2632,N_45534,N_48720);
nor UO_2633 (O_2633,N_45050,N_45846);
nor UO_2634 (O_2634,N_46582,N_45133);
nor UO_2635 (O_2635,N_46016,N_49820);
nand UO_2636 (O_2636,N_46130,N_45511);
and UO_2637 (O_2637,N_46957,N_47338);
xnor UO_2638 (O_2638,N_49992,N_49327);
nor UO_2639 (O_2639,N_48021,N_48741);
nand UO_2640 (O_2640,N_48081,N_45933);
nor UO_2641 (O_2641,N_48521,N_45521);
nand UO_2642 (O_2642,N_46240,N_48199);
or UO_2643 (O_2643,N_47667,N_46606);
and UO_2644 (O_2644,N_47100,N_45303);
xor UO_2645 (O_2645,N_49621,N_45093);
nand UO_2646 (O_2646,N_46610,N_47082);
nand UO_2647 (O_2647,N_45332,N_48560);
nand UO_2648 (O_2648,N_48236,N_49512);
and UO_2649 (O_2649,N_48423,N_48138);
nor UO_2650 (O_2650,N_45758,N_48666);
and UO_2651 (O_2651,N_49020,N_49158);
or UO_2652 (O_2652,N_47566,N_48779);
or UO_2653 (O_2653,N_48922,N_46949);
or UO_2654 (O_2654,N_47162,N_45781);
nand UO_2655 (O_2655,N_47361,N_49605);
xor UO_2656 (O_2656,N_46754,N_46642);
and UO_2657 (O_2657,N_48738,N_49913);
or UO_2658 (O_2658,N_47996,N_48469);
and UO_2659 (O_2659,N_46297,N_49508);
nand UO_2660 (O_2660,N_49630,N_47271);
and UO_2661 (O_2661,N_49304,N_47966);
or UO_2662 (O_2662,N_45893,N_48856);
xnor UO_2663 (O_2663,N_48275,N_48483);
nand UO_2664 (O_2664,N_49272,N_48416);
xor UO_2665 (O_2665,N_49024,N_47494);
and UO_2666 (O_2666,N_47829,N_46588);
xnor UO_2667 (O_2667,N_46609,N_46972);
nor UO_2668 (O_2668,N_48089,N_47637);
and UO_2669 (O_2669,N_49705,N_47498);
and UO_2670 (O_2670,N_48594,N_49046);
or UO_2671 (O_2671,N_48070,N_49187);
nand UO_2672 (O_2672,N_48413,N_48442);
and UO_2673 (O_2673,N_46116,N_45450);
xor UO_2674 (O_2674,N_46763,N_49440);
or UO_2675 (O_2675,N_49468,N_45634);
nand UO_2676 (O_2676,N_47652,N_48645);
xnor UO_2677 (O_2677,N_45520,N_49324);
xor UO_2678 (O_2678,N_46409,N_48015);
nand UO_2679 (O_2679,N_46515,N_48707);
or UO_2680 (O_2680,N_45994,N_49910);
nor UO_2681 (O_2681,N_47962,N_45614);
xor UO_2682 (O_2682,N_49295,N_46448);
or UO_2683 (O_2683,N_46151,N_46111);
nor UO_2684 (O_2684,N_46460,N_47610);
nor UO_2685 (O_2685,N_47148,N_45098);
nand UO_2686 (O_2686,N_49023,N_48558);
xnor UO_2687 (O_2687,N_45539,N_46994);
nor UO_2688 (O_2688,N_48439,N_49172);
or UO_2689 (O_2689,N_45937,N_48853);
and UO_2690 (O_2690,N_46700,N_46900);
xor UO_2691 (O_2691,N_47356,N_47157);
and UO_2692 (O_2692,N_46141,N_47391);
nor UO_2693 (O_2693,N_49619,N_46822);
xor UO_2694 (O_2694,N_46166,N_45855);
nand UO_2695 (O_2695,N_49726,N_48770);
and UO_2696 (O_2696,N_46833,N_49972);
nor UO_2697 (O_2697,N_45833,N_48423);
nand UO_2698 (O_2698,N_46566,N_47055);
xor UO_2699 (O_2699,N_49764,N_46958);
nor UO_2700 (O_2700,N_49668,N_47616);
nor UO_2701 (O_2701,N_48418,N_45052);
nor UO_2702 (O_2702,N_49520,N_47949);
or UO_2703 (O_2703,N_46706,N_45563);
nand UO_2704 (O_2704,N_48194,N_48955);
xnor UO_2705 (O_2705,N_46680,N_48343);
nor UO_2706 (O_2706,N_47501,N_47902);
and UO_2707 (O_2707,N_45634,N_49733);
xor UO_2708 (O_2708,N_47145,N_47054);
nor UO_2709 (O_2709,N_48947,N_49117);
and UO_2710 (O_2710,N_49708,N_48925);
nor UO_2711 (O_2711,N_45512,N_48760);
nand UO_2712 (O_2712,N_47033,N_46384);
nor UO_2713 (O_2713,N_46048,N_46652);
xnor UO_2714 (O_2714,N_49274,N_49682);
nand UO_2715 (O_2715,N_47952,N_48287);
nand UO_2716 (O_2716,N_46780,N_49463);
xor UO_2717 (O_2717,N_45107,N_47240);
nor UO_2718 (O_2718,N_47433,N_47713);
and UO_2719 (O_2719,N_46315,N_46639);
and UO_2720 (O_2720,N_45395,N_45294);
nand UO_2721 (O_2721,N_47258,N_47098);
or UO_2722 (O_2722,N_48076,N_45576);
xnor UO_2723 (O_2723,N_47423,N_48596);
and UO_2724 (O_2724,N_45479,N_49909);
nor UO_2725 (O_2725,N_46308,N_49261);
or UO_2726 (O_2726,N_46622,N_49006);
or UO_2727 (O_2727,N_45719,N_48483);
xor UO_2728 (O_2728,N_49364,N_46650);
and UO_2729 (O_2729,N_49573,N_48822);
nand UO_2730 (O_2730,N_46458,N_48250);
and UO_2731 (O_2731,N_46110,N_49914);
xor UO_2732 (O_2732,N_48376,N_46660);
and UO_2733 (O_2733,N_48283,N_46753);
nor UO_2734 (O_2734,N_46490,N_46807);
nor UO_2735 (O_2735,N_46413,N_45356);
xnor UO_2736 (O_2736,N_46658,N_49088);
and UO_2737 (O_2737,N_47897,N_46535);
nor UO_2738 (O_2738,N_48170,N_45761);
or UO_2739 (O_2739,N_49411,N_49939);
nor UO_2740 (O_2740,N_46404,N_49172);
and UO_2741 (O_2741,N_45989,N_46538);
or UO_2742 (O_2742,N_45065,N_46616);
nand UO_2743 (O_2743,N_46967,N_47411);
nor UO_2744 (O_2744,N_47173,N_46942);
nor UO_2745 (O_2745,N_45916,N_46882);
and UO_2746 (O_2746,N_49850,N_49983);
and UO_2747 (O_2747,N_48239,N_48764);
xnor UO_2748 (O_2748,N_49363,N_47954);
or UO_2749 (O_2749,N_45585,N_49475);
and UO_2750 (O_2750,N_46302,N_49903);
and UO_2751 (O_2751,N_46863,N_48222);
xnor UO_2752 (O_2752,N_46853,N_47053);
and UO_2753 (O_2753,N_48026,N_49300);
and UO_2754 (O_2754,N_45275,N_49407);
and UO_2755 (O_2755,N_48540,N_47660);
and UO_2756 (O_2756,N_48512,N_45705);
and UO_2757 (O_2757,N_45762,N_45619);
xnor UO_2758 (O_2758,N_46442,N_45898);
nand UO_2759 (O_2759,N_48421,N_48666);
nand UO_2760 (O_2760,N_48822,N_45328);
nand UO_2761 (O_2761,N_45322,N_49897);
and UO_2762 (O_2762,N_48936,N_46222);
xor UO_2763 (O_2763,N_46980,N_45030);
xor UO_2764 (O_2764,N_45930,N_46894);
and UO_2765 (O_2765,N_48118,N_45589);
and UO_2766 (O_2766,N_49421,N_46915);
or UO_2767 (O_2767,N_47905,N_45393);
nand UO_2768 (O_2768,N_49560,N_49772);
nor UO_2769 (O_2769,N_49134,N_48320);
nor UO_2770 (O_2770,N_45109,N_47776);
and UO_2771 (O_2771,N_49112,N_47354);
or UO_2772 (O_2772,N_48963,N_48798);
xor UO_2773 (O_2773,N_49018,N_46502);
nand UO_2774 (O_2774,N_46352,N_49707);
or UO_2775 (O_2775,N_47372,N_48265);
or UO_2776 (O_2776,N_47881,N_46875);
nand UO_2777 (O_2777,N_49465,N_49363);
nor UO_2778 (O_2778,N_45894,N_46371);
and UO_2779 (O_2779,N_46272,N_46816);
xor UO_2780 (O_2780,N_45573,N_46988);
or UO_2781 (O_2781,N_47915,N_49890);
nor UO_2782 (O_2782,N_47999,N_48246);
or UO_2783 (O_2783,N_45917,N_47060);
nand UO_2784 (O_2784,N_49804,N_49067);
and UO_2785 (O_2785,N_48312,N_46727);
xor UO_2786 (O_2786,N_47167,N_49985);
xnor UO_2787 (O_2787,N_48787,N_46031);
nor UO_2788 (O_2788,N_46206,N_48485);
and UO_2789 (O_2789,N_46179,N_45255);
nand UO_2790 (O_2790,N_46593,N_47214);
nor UO_2791 (O_2791,N_49476,N_47070);
nand UO_2792 (O_2792,N_47579,N_48252);
or UO_2793 (O_2793,N_45519,N_46211);
nor UO_2794 (O_2794,N_46806,N_48882);
nand UO_2795 (O_2795,N_45068,N_46505);
or UO_2796 (O_2796,N_46618,N_49925);
xnor UO_2797 (O_2797,N_48219,N_48070);
and UO_2798 (O_2798,N_45956,N_46172);
nor UO_2799 (O_2799,N_47146,N_45413);
or UO_2800 (O_2800,N_45052,N_48810);
nor UO_2801 (O_2801,N_46726,N_46131);
xor UO_2802 (O_2802,N_46833,N_46275);
and UO_2803 (O_2803,N_49476,N_45950);
nor UO_2804 (O_2804,N_46745,N_46256);
xor UO_2805 (O_2805,N_48215,N_45242);
or UO_2806 (O_2806,N_47505,N_48933);
xnor UO_2807 (O_2807,N_47200,N_47208);
and UO_2808 (O_2808,N_47792,N_45766);
and UO_2809 (O_2809,N_48517,N_48001);
and UO_2810 (O_2810,N_47833,N_47267);
xor UO_2811 (O_2811,N_49158,N_47396);
xor UO_2812 (O_2812,N_49681,N_48772);
and UO_2813 (O_2813,N_45738,N_45806);
xor UO_2814 (O_2814,N_45068,N_48650);
nand UO_2815 (O_2815,N_45274,N_49575);
nor UO_2816 (O_2816,N_48775,N_48722);
nand UO_2817 (O_2817,N_45211,N_47523);
or UO_2818 (O_2818,N_49961,N_49539);
nand UO_2819 (O_2819,N_49572,N_46774);
or UO_2820 (O_2820,N_49394,N_49401);
and UO_2821 (O_2821,N_47424,N_48486);
or UO_2822 (O_2822,N_48441,N_48629);
nand UO_2823 (O_2823,N_46761,N_46065);
nor UO_2824 (O_2824,N_47336,N_48892);
nand UO_2825 (O_2825,N_47806,N_46255);
nor UO_2826 (O_2826,N_45212,N_46613);
and UO_2827 (O_2827,N_48722,N_47823);
or UO_2828 (O_2828,N_47022,N_48840);
nor UO_2829 (O_2829,N_48814,N_46769);
or UO_2830 (O_2830,N_49908,N_47234);
and UO_2831 (O_2831,N_48055,N_48842);
xor UO_2832 (O_2832,N_46437,N_46518);
nor UO_2833 (O_2833,N_49128,N_46351);
and UO_2834 (O_2834,N_46546,N_45327);
xor UO_2835 (O_2835,N_48569,N_48176);
nand UO_2836 (O_2836,N_45569,N_47540);
nor UO_2837 (O_2837,N_48090,N_45684);
xnor UO_2838 (O_2838,N_49669,N_48754);
nor UO_2839 (O_2839,N_45377,N_48053);
and UO_2840 (O_2840,N_49024,N_46890);
nor UO_2841 (O_2841,N_46529,N_46875);
nor UO_2842 (O_2842,N_48215,N_47257);
and UO_2843 (O_2843,N_47462,N_45499);
nand UO_2844 (O_2844,N_46700,N_47140);
xor UO_2845 (O_2845,N_48600,N_47927);
nor UO_2846 (O_2846,N_45165,N_47462);
xor UO_2847 (O_2847,N_49078,N_46282);
xor UO_2848 (O_2848,N_48493,N_47528);
and UO_2849 (O_2849,N_47434,N_47937);
xnor UO_2850 (O_2850,N_48208,N_48152);
or UO_2851 (O_2851,N_47398,N_49958);
and UO_2852 (O_2852,N_45514,N_45666);
or UO_2853 (O_2853,N_48097,N_49237);
and UO_2854 (O_2854,N_45819,N_46989);
xnor UO_2855 (O_2855,N_46729,N_48427);
or UO_2856 (O_2856,N_48933,N_48762);
nor UO_2857 (O_2857,N_45923,N_46972);
or UO_2858 (O_2858,N_48919,N_48720);
xor UO_2859 (O_2859,N_49373,N_49066);
nor UO_2860 (O_2860,N_47653,N_45594);
xnor UO_2861 (O_2861,N_49558,N_49662);
and UO_2862 (O_2862,N_47132,N_48270);
and UO_2863 (O_2863,N_49532,N_48744);
and UO_2864 (O_2864,N_46110,N_45150);
or UO_2865 (O_2865,N_49967,N_48490);
nand UO_2866 (O_2866,N_45032,N_47612);
nor UO_2867 (O_2867,N_47470,N_49386);
or UO_2868 (O_2868,N_49552,N_46938);
nand UO_2869 (O_2869,N_46916,N_49416);
nor UO_2870 (O_2870,N_45989,N_48226);
xor UO_2871 (O_2871,N_46808,N_45888);
and UO_2872 (O_2872,N_47062,N_46938);
or UO_2873 (O_2873,N_48147,N_47014);
or UO_2874 (O_2874,N_47400,N_48707);
nand UO_2875 (O_2875,N_47007,N_45304);
and UO_2876 (O_2876,N_47087,N_48305);
and UO_2877 (O_2877,N_45209,N_49406);
nand UO_2878 (O_2878,N_48045,N_49740);
and UO_2879 (O_2879,N_46916,N_47705);
nand UO_2880 (O_2880,N_49620,N_47286);
xor UO_2881 (O_2881,N_48832,N_46576);
or UO_2882 (O_2882,N_46035,N_49026);
xor UO_2883 (O_2883,N_46767,N_45145);
xnor UO_2884 (O_2884,N_45087,N_45904);
nor UO_2885 (O_2885,N_48104,N_48425);
nor UO_2886 (O_2886,N_48696,N_45915);
xnor UO_2887 (O_2887,N_49342,N_47687);
nand UO_2888 (O_2888,N_45520,N_46256);
xnor UO_2889 (O_2889,N_47693,N_45263);
and UO_2890 (O_2890,N_45500,N_46727);
nand UO_2891 (O_2891,N_48633,N_45302);
xnor UO_2892 (O_2892,N_49653,N_47911);
or UO_2893 (O_2893,N_49206,N_45565);
nor UO_2894 (O_2894,N_48453,N_49126);
and UO_2895 (O_2895,N_49426,N_49288);
xnor UO_2896 (O_2896,N_48504,N_49395);
nand UO_2897 (O_2897,N_46531,N_47363);
nor UO_2898 (O_2898,N_45673,N_46666);
xor UO_2899 (O_2899,N_48301,N_46055);
nor UO_2900 (O_2900,N_49660,N_47326);
nand UO_2901 (O_2901,N_48165,N_46577);
nor UO_2902 (O_2902,N_48726,N_48637);
nor UO_2903 (O_2903,N_47078,N_47047);
and UO_2904 (O_2904,N_49489,N_45045);
or UO_2905 (O_2905,N_45846,N_45258);
nand UO_2906 (O_2906,N_48536,N_46286);
or UO_2907 (O_2907,N_48494,N_48767);
nor UO_2908 (O_2908,N_46530,N_45444);
xnor UO_2909 (O_2909,N_48513,N_47797);
nor UO_2910 (O_2910,N_46814,N_49223);
nor UO_2911 (O_2911,N_48091,N_49970);
and UO_2912 (O_2912,N_49787,N_49203);
nand UO_2913 (O_2913,N_45327,N_46075);
and UO_2914 (O_2914,N_47531,N_45060);
or UO_2915 (O_2915,N_49327,N_45346);
nand UO_2916 (O_2916,N_46369,N_47264);
nand UO_2917 (O_2917,N_46800,N_47850);
nor UO_2918 (O_2918,N_47789,N_46985);
and UO_2919 (O_2919,N_47838,N_47791);
and UO_2920 (O_2920,N_45972,N_49319);
or UO_2921 (O_2921,N_47855,N_45771);
xnor UO_2922 (O_2922,N_46131,N_47755);
nor UO_2923 (O_2923,N_47940,N_46875);
xnor UO_2924 (O_2924,N_46761,N_48600);
or UO_2925 (O_2925,N_46796,N_46939);
nor UO_2926 (O_2926,N_48472,N_48897);
nor UO_2927 (O_2927,N_47087,N_47468);
xor UO_2928 (O_2928,N_48018,N_46607);
nor UO_2929 (O_2929,N_49249,N_46098);
or UO_2930 (O_2930,N_45511,N_45135);
or UO_2931 (O_2931,N_45307,N_48871);
nand UO_2932 (O_2932,N_45341,N_47964);
nand UO_2933 (O_2933,N_49891,N_48979);
nor UO_2934 (O_2934,N_45523,N_48046);
nor UO_2935 (O_2935,N_46998,N_47093);
or UO_2936 (O_2936,N_47789,N_46329);
and UO_2937 (O_2937,N_48861,N_46963);
nand UO_2938 (O_2938,N_48711,N_48703);
xor UO_2939 (O_2939,N_47352,N_49544);
xnor UO_2940 (O_2940,N_46198,N_49312);
xnor UO_2941 (O_2941,N_48335,N_47485);
xor UO_2942 (O_2942,N_47397,N_48612);
and UO_2943 (O_2943,N_45808,N_48311);
or UO_2944 (O_2944,N_48149,N_45134);
and UO_2945 (O_2945,N_45898,N_47694);
and UO_2946 (O_2946,N_46154,N_46286);
xnor UO_2947 (O_2947,N_48808,N_49483);
nor UO_2948 (O_2948,N_49471,N_48237);
nor UO_2949 (O_2949,N_49053,N_45914);
or UO_2950 (O_2950,N_46239,N_47658);
nand UO_2951 (O_2951,N_49631,N_48112);
and UO_2952 (O_2952,N_48437,N_46990);
and UO_2953 (O_2953,N_49223,N_45225);
and UO_2954 (O_2954,N_48731,N_45386);
nor UO_2955 (O_2955,N_46559,N_47665);
nand UO_2956 (O_2956,N_47291,N_47343);
nand UO_2957 (O_2957,N_48456,N_46725);
nor UO_2958 (O_2958,N_49290,N_49487);
xnor UO_2959 (O_2959,N_46436,N_47003);
and UO_2960 (O_2960,N_47761,N_45895);
xnor UO_2961 (O_2961,N_46495,N_46801);
nand UO_2962 (O_2962,N_45834,N_48900);
xnor UO_2963 (O_2963,N_46103,N_48203);
or UO_2964 (O_2964,N_46699,N_46572);
or UO_2965 (O_2965,N_47178,N_45220);
and UO_2966 (O_2966,N_45250,N_49275);
xnor UO_2967 (O_2967,N_46903,N_49778);
or UO_2968 (O_2968,N_47356,N_45632);
nor UO_2969 (O_2969,N_47815,N_46893);
xnor UO_2970 (O_2970,N_48224,N_47868);
or UO_2971 (O_2971,N_47608,N_47753);
and UO_2972 (O_2972,N_48948,N_48967);
xnor UO_2973 (O_2973,N_49885,N_49431);
and UO_2974 (O_2974,N_45809,N_49953);
and UO_2975 (O_2975,N_49086,N_49769);
or UO_2976 (O_2976,N_45022,N_46292);
nand UO_2977 (O_2977,N_45795,N_47424);
nor UO_2978 (O_2978,N_45084,N_48824);
and UO_2979 (O_2979,N_49228,N_49230);
xnor UO_2980 (O_2980,N_49717,N_47516);
and UO_2981 (O_2981,N_45292,N_46884);
nor UO_2982 (O_2982,N_48533,N_49728);
nand UO_2983 (O_2983,N_49105,N_45804);
and UO_2984 (O_2984,N_49498,N_48439);
or UO_2985 (O_2985,N_49455,N_47249);
or UO_2986 (O_2986,N_45687,N_48441);
nor UO_2987 (O_2987,N_46388,N_49227);
nor UO_2988 (O_2988,N_45126,N_46419);
nor UO_2989 (O_2989,N_45113,N_47612);
nor UO_2990 (O_2990,N_46193,N_46590);
nor UO_2991 (O_2991,N_47022,N_45398);
nand UO_2992 (O_2992,N_45095,N_45992);
nor UO_2993 (O_2993,N_46017,N_45788);
nor UO_2994 (O_2994,N_46655,N_45754);
and UO_2995 (O_2995,N_46394,N_45099);
and UO_2996 (O_2996,N_49932,N_47289);
nand UO_2997 (O_2997,N_45995,N_47805);
or UO_2998 (O_2998,N_46160,N_47262);
or UO_2999 (O_2999,N_46588,N_49389);
and UO_3000 (O_3000,N_48802,N_45556);
or UO_3001 (O_3001,N_46508,N_49103);
and UO_3002 (O_3002,N_48203,N_49633);
nor UO_3003 (O_3003,N_47960,N_47576);
nor UO_3004 (O_3004,N_45443,N_45706);
and UO_3005 (O_3005,N_46349,N_49155);
or UO_3006 (O_3006,N_49248,N_47907);
xor UO_3007 (O_3007,N_47684,N_49595);
and UO_3008 (O_3008,N_46380,N_48369);
or UO_3009 (O_3009,N_47450,N_47775);
nand UO_3010 (O_3010,N_48813,N_47822);
nand UO_3011 (O_3011,N_49960,N_45369);
nand UO_3012 (O_3012,N_45181,N_46747);
xnor UO_3013 (O_3013,N_49310,N_49971);
or UO_3014 (O_3014,N_48179,N_46049);
or UO_3015 (O_3015,N_49353,N_46272);
and UO_3016 (O_3016,N_48379,N_49011);
or UO_3017 (O_3017,N_47260,N_49723);
or UO_3018 (O_3018,N_46365,N_45586);
and UO_3019 (O_3019,N_48266,N_49136);
nor UO_3020 (O_3020,N_47973,N_47196);
nor UO_3021 (O_3021,N_49744,N_45568);
nor UO_3022 (O_3022,N_45427,N_47341);
or UO_3023 (O_3023,N_45684,N_45559);
xnor UO_3024 (O_3024,N_47766,N_49114);
xor UO_3025 (O_3025,N_46945,N_48185);
nor UO_3026 (O_3026,N_48005,N_45102);
or UO_3027 (O_3027,N_48034,N_49253);
nand UO_3028 (O_3028,N_46413,N_46398);
nor UO_3029 (O_3029,N_46275,N_49185);
and UO_3030 (O_3030,N_45520,N_47391);
xor UO_3031 (O_3031,N_49266,N_45148);
and UO_3032 (O_3032,N_47315,N_46154);
or UO_3033 (O_3033,N_47871,N_49104);
and UO_3034 (O_3034,N_47231,N_49228);
nand UO_3035 (O_3035,N_48540,N_49386);
or UO_3036 (O_3036,N_48238,N_46305);
nand UO_3037 (O_3037,N_49485,N_49144);
nor UO_3038 (O_3038,N_45286,N_47778);
and UO_3039 (O_3039,N_49447,N_47105);
xnor UO_3040 (O_3040,N_45156,N_46638);
and UO_3041 (O_3041,N_47860,N_48096);
nor UO_3042 (O_3042,N_46888,N_48471);
xor UO_3043 (O_3043,N_46804,N_49972);
and UO_3044 (O_3044,N_47397,N_47054);
and UO_3045 (O_3045,N_49496,N_48155);
nand UO_3046 (O_3046,N_45588,N_47954);
nand UO_3047 (O_3047,N_47076,N_48055);
nand UO_3048 (O_3048,N_48099,N_46701);
nand UO_3049 (O_3049,N_45514,N_45751);
nor UO_3050 (O_3050,N_49102,N_49974);
xnor UO_3051 (O_3051,N_48183,N_47447);
nand UO_3052 (O_3052,N_47486,N_45247);
nand UO_3053 (O_3053,N_48175,N_47586);
and UO_3054 (O_3054,N_46339,N_48371);
or UO_3055 (O_3055,N_45689,N_47884);
nor UO_3056 (O_3056,N_49736,N_47164);
nor UO_3057 (O_3057,N_49473,N_45783);
and UO_3058 (O_3058,N_48068,N_49729);
xnor UO_3059 (O_3059,N_46749,N_49919);
nand UO_3060 (O_3060,N_47366,N_49760);
and UO_3061 (O_3061,N_45290,N_47805);
xnor UO_3062 (O_3062,N_47509,N_48601);
xor UO_3063 (O_3063,N_45737,N_46191);
and UO_3064 (O_3064,N_45303,N_47802);
xnor UO_3065 (O_3065,N_45526,N_46685);
nor UO_3066 (O_3066,N_46390,N_47138);
xnor UO_3067 (O_3067,N_48718,N_47327);
or UO_3068 (O_3068,N_49967,N_46501);
and UO_3069 (O_3069,N_47035,N_48386);
xor UO_3070 (O_3070,N_45612,N_46505);
nor UO_3071 (O_3071,N_45453,N_47061);
xnor UO_3072 (O_3072,N_45022,N_48265);
and UO_3073 (O_3073,N_46640,N_48268);
and UO_3074 (O_3074,N_45336,N_45175);
xor UO_3075 (O_3075,N_49812,N_46315);
and UO_3076 (O_3076,N_49077,N_49255);
xnor UO_3077 (O_3077,N_47674,N_45778);
and UO_3078 (O_3078,N_47808,N_45796);
and UO_3079 (O_3079,N_46683,N_47618);
xor UO_3080 (O_3080,N_46201,N_47647);
xnor UO_3081 (O_3081,N_49951,N_46736);
xor UO_3082 (O_3082,N_46672,N_45661);
xnor UO_3083 (O_3083,N_48235,N_47941);
nor UO_3084 (O_3084,N_48694,N_47931);
or UO_3085 (O_3085,N_49707,N_46569);
nor UO_3086 (O_3086,N_47601,N_49650);
nor UO_3087 (O_3087,N_49743,N_46018);
xnor UO_3088 (O_3088,N_49287,N_46176);
nor UO_3089 (O_3089,N_48030,N_49583);
xor UO_3090 (O_3090,N_45376,N_49147);
xor UO_3091 (O_3091,N_45145,N_45659);
and UO_3092 (O_3092,N_46591,N_47358);
or UO_3093 (O_3093,N_46564,N_47043);
nor UO_3094 (O_3094,N_49938,N_49673);
xnor UO_3095 (O_3095,N_46597,N_49575);
nor UO_3096 (O_3096,N_45414,N_46092);
and UO_3097 (O_3097,N_45353,N_46620);
and UO_3098 (O_3098,N_47157,N_48069);
or UO_3099 (O_3099,N_45884,N_49942);
nand UO_3100 (O_3100,N_45211,N_48725);
or UO_3101 (O_3101,N_49927,N_49498);
and UO_3102 (O_3102,N_46480,N_47066);
nor UO_3103 (O_3103,N_46608,N_48087);
nand UO_3104 (O_3104,N_47121,N_47835);
or UO_3105 (O_3105,N_48820,N_47972);
nor UO_3106 (O_3106,N_48059,N_47466);
or UO_3107 (O_3107,N_46456,N_46548);
or UO_3108 (O_3108,N_45997,N_48441);
nor UO_3109 (O_3109,N_47521,N_48610);
and UO_3110 (O_3110,N_46434,N_46358);
nor UO_3111 (O_3111,N_45722,N_49888);
nor UO_3112 (O_3112,N_48613,N_47742);
xor UO_3113 (O_3113,N_47961,N_46271);
or UO_3114 (O_3114,N_47193,N_47972);
nor UO_3115 (O_3115,N_48101,N_49315);
and UO_3116 (O_3116,N_48009,N_48668);
xnor UO_3117 (O_3117,N_48394,N_45245);
nand UO_3118 (O_3118,N_45304,N_49982);
and UO_3119 (O_3119,N_45254,N_45589);
xor UO_3120 (O_3120,N_48578,N_49990);
and UO_3121 (O_3121,N_48975,N_45949);
nand UO_3122 (O_3122,N_46185,N_48048);
and UO_3123 (O_3123,N_47568,N_47777);
nor UO_3124 (O_3124,N_47057,N_47640);
and UO_3125 (O_3125,N_49079,N_46082);
nor UO_3126 (O_3126,N_49694,N_47866);
and UO_3127 (O_3127,N_45592,N_48914);
and UO_3128 (O_3128,N_49933,N_49418);
xor UO_3129 (O_3129,N_47252,N_48073);
nand UO_3130 (O_3130,N_48143,N_48097);
or UO_3131 (O_3131,N_45215,N_46486);
or UO_3132 (O_3132,N_47906,N_49170);
nand UO_3133 (O_3133,N_49959,N_47817);
nor UO_3134 (O_3134,N_46287,N_47239);
xor UO_3135 (O_3135,N_46792,N_47218);
nand UO_3136 (O_3136,N_49012,N_46993);
nand UO_3137 (O_3137,N_47898,N_49034);
nor UO_3138 (O_3138,N_48027,N_49901);
and UO_3139 (O_3139,N_46718,N_49543);
nor UO_3140 (O_3140,N_45910,N_49467);
nand UO_3141 (O_3141,N_45397,N_46158);
and UO_3142 (O_3142,N_48829,N_45054);
nor UO_3143 (O_3143,N_45655,N_46031);
or UO_3144 (O_3144,N_45780,N_45178);
nor UO_3145 (O_3145,N_45472,N_47234);
or UO_3146 (O_3146,N_48915,N_48129);
and UO_3147 (O_3147,N_46870,N_48995);
xnor UO_3148 (O_3148,N_48092,N_49099);
nand UO_3149 (O_3149,N_48009,N_45452);
xnor UO_3150 (O_3150,N_48984,N_46917);
nor UO_3151 (O_3151,N_49319,N_47339);
nand UO_3152 (O_3152,N_47393,N_45733);
or UO_3153 (O_3153,N_49201,N_45597);
nand UO_3154 (O_3154,N_45749,N_48171);
or UO_3155 (O_3155,N_49732,N_48530);
or UO_3156 (O_3156,N_48595,N_46951);
or UO_3157 (O_3157,N_49614,N_48728);
or UO_3158 (O_3158,N_46018,N_47981);
and UO_3159 (O_3159,N_49997,N_48500);
nand UO_3160 (O_3160,N_48964,N_46826);
nand UO_3161 (O_3161,N_48759,N_46068);
and UO_3162 (O_3162,N_47828,N_45198);
xor UO_3163 (O_3163,N_46515,N_48874);
nand UO_3164 (O_3164,N_49460,N_46389);
nor UO_3165 (O_3165,N_47909,N_46035);
nor UO_3166 (O_3166,N_47619,N_48153);
nor UO_3167 (O_3167,N_48415,N_48236);
nand UO_3168 (O_3168,N_47898,N_49275);
nor UO_3169 (O_3169,N_46639,N_46344);
nor UO_3170 (O_3170,N_46957,N_49204);
nand UO_3171 (O_3171,N_48319,N_49867);
nand UO_3172 (O_3172,N_49111,N_46984);
and UO_3173 (O_3173,N_47705,N_49979);
nor UO_3174 (O_3174,N_45467,N_48606);
xor UO_3175 (O_3175,N_45752,N_47347);
or UO_3176 (O_3176,N_46581,N_46089);
or UO_3177 (O_3177,N_47376,N_47650);
nor UO_3178 (O_3178,N_49735,N_46772);
nand UO_3179 (O_3179,N_46132,N_46186);
nand UO_3180 (O_3180,N_48390,N_48194);
and UO_3181 (O_3181,N_48086,N_48796);
or UO_3182 (O_3182,N_46764,N_49533);
or UO_3183 (O_3183,N_46122,N_45610);
nand UO_3184 (O_3184,N_48258,N_48592);
xnor UO_3185 (O_3185,N_46665,N_47485);
nand UO_3186 (O_3186,N_45179,N_47895);
and UO_3187 (O_3187,N_45731,N_46562);
or UO_3188 (O_3188,N_45646,N_48014);
xnor UO_3189 (O_3189,N_49892,N_49471);
xnor UO_3190 (O_3190,N_45646,N_46739);
nand UO_3191 (O_3191,N_49573,N_47995);
or UO_3192 (O_3192,N_48964,N_49521);
and UO_3193 (O_3193,N_49436,N_49348);
nor UO_3194 (O_3194,N_47097,N_48793);
or UO_3195 (O_3195,N_45498,N_48540);
and UO_3196 (O_3196,N_45832,N_46363);
nor UO_3197 (O_3197,N_45130,N_45256);
xor UO_3198 (O_3198,N_46761,N_47513);
nand UO_3199 (O_3199,N_47011,N_48118);
and UO_3200 (O_3200,N_47583,N_46475);
nand UO_3201 (O_3201,N_45400,N_47698);
nand UO_3202 (O_3202,N_48154,N_46554);
nor UO_3203 (O_3203,N_48342,N_49312);
or UO_3204 (O_3204,N_47148,N_45606);
xnor UO_3205 (O_3205,N_48855,N_49129);
xor UO_3206 (O_3206,N_47711,N_48875);
and UO_3207 (O_3207,N_48808,N_46354);
nor UO_3208 (O_3208,N_49262,N_48901);
xnor UO_3209 (O_3209,N_47768,N_49803);
nor UO_3210 (O_3210,N_45504,N_49412);
or UO_3211 (O_3211,N_49078,N_47080);
or UO_3212 (O_3212,N_48424,N_48380);
nand UO_3213 (O_3213,N_49620,N_45167);
or UO_3214 (O_3214,N_48238,N_47123);
and UO_3215 (O_3215,N_45816,N_49473);
xnor UO_3216 (O_3216,N_46652,N_49552);
xnor UO_3217 (O_3217,N_45722,N_48257);
nand UO_3218 (O_3218,N_45160,N_45482);
or UO_3219 (O_3219,N_46353,N_46457);
and UO_3220 (O_3220,N_48206,N_45933);
nand UO_3221 (O_3221,N_47475,N_49782);
xnor UO_3222 (O_3222,N_45724,N_46445);
nand UO_3223 (O_3223,N_48496,N_46185);
nor UO_3224 (O_3224,N_45969,N_49620);
nand UO_3225 (O_3225,N_48407,N_45151);
or UO_3226 (O_3226,N_49467,N_48967);
and UO_3227 (O_3227,N_45562,N_48401);
xnor UO_3228 (O_3228,N_45585,N_47540);
xor UO_3229 (O_3229,N_46045,N_49118);
or UO_3230 (O_3230,N_45922,N_45268);
nand UO_3231 (O_3231,N_48599,N_48452);
or UO_3232 (O_3232,N_46560,N_46421);
nor UO_3233 (O_3233,N_45120,N_46766);
xor UO_3234 (O_3234,N_47102,N_48977);
nand UO_3235 (O_3235,N_46683,N_47525);
and UO_3236 (O_3236,N_47136,N_48241);
or UO_3237 (O_3237,N_46698,N_49275);
nor UO_3238 (O_3238,N_47669,N_46972);
and UO_3239 (O_3239,N_46464,N_45792);
and UO_3240 (O_3240,N_47406,N_48526);
xor UO_3241 (O_3241,N_49826,N_49080);
and UO_3242 (O_3242,N_46465,N_49002);
xor UO_3243 (O_3243,N_47509,N_47646);
xor UO_3244 (O_3244,N_47733,N_45961);
nor UO_3245 (O_3245,N_47993,N_47595);
and UO_3246 (O_3246,N_47900,N_48133);
nand UO_3247 (O_3247,N_48723,N_49867);
xnor UO_3248 (O_3248,N_47707,N_48430);
nor UO_3249 (O_3249,N_45982,N_49651);
xnor UO_3250 (O_3250,N_49696,N_46817);
nor UO_3251 (O_3251,N_47588,N_46423);
nand UO_3252 (O_3252,N_45873,N_46415);
nor UO_3253 (O_3253,N_48441,N_49391);
nand UO_3254 (O_3254,N_49988,N_48574);
or UO_3255 (O_3255,N_48843,N_47976);
xnor UO_3256 (O_3256,N_46248,N_46691);
or UO_3257 (O_3257,N_49856,N_45112);
nand UO_3258 (O_3258,N_47102,N_47301);
xnor UO_3259 (O_3259,N_45025,N_49990);
nor UO_3260 (O_3260,N_45630,N_48067);
nand UO_3261 (O_3261,N_48698,N_48837);
nand UO_3262 (O_3262,N_46839,N_46230);
nand UO_3263 (O_3263,N_47642,N_47860);
nand UO_3264 (O_3264,N_47306,N_47732);
nor UO_3265 (O_3265,N_48995,N_46261);
nand UO_3266 (O_3266,N_46029,N_49932);
nand UO_3267 (O_3267,N_45567,N_45929);
xnor UO_3268 (O_3268,N_46659,N_45085);
nor UO_3269 (O_3269,N_47455,N_45357);
xnor UO_3270 (O_3270,N_48115,N_49107);
nor UO_3271 (O_3271,N_47689,N_47022);
and UO_3272 (O_3272,N_49741,N_49678);
xnor UO_3273 (O_3273,N_45471,N_47421);
xnor UO_3274 (O_3274,N_45557,N_47035);
or UO_3275 (O_3275,N_48009,N_47881);
and UO_3276 (O_3276,N_46845,N_49530);
and UO_3277 (O_3277,N_49360,N_46841);
and UO_3278 (O_3278,N_45161,N_48233);
xor UO_3279 (O_3279,N_48547,N_45574);
nand UO_3280 (O_3280,N_45982,N_45037);
nand UO_3281 (O_3281,N_47658,N_48699);
and UO_3282 (O_3282,N_47031,N_45476);
xnor UO_3283 (O_3283,N_47584,N_48800);
nand UO_3284 (O_3284,N_49196,N_49706);
and UO_3285 (O_3285,N_47417,N_48754);
xor UO_3286 (O_3286,N_46759,N_47503);
nand UO_3287 (O_3287,N_45815,N_45871);
nor UO_3288 (O_3288,N_47625,N_48009);
nor UO_3289 (O_3289,N_47491,N_48684);
and UO_3290 (O_3290,N_47499,N_47043);
xnor UO_3291 (O_3291,N_47204,N_45672);
nand UO_3292 (O_3292,N_45562,N_48566);
nor UO_3293 (O_3293,N_47972,N_47284);
or UO_3294 (O_3294,N_47102,N_47383);
and UO_3295 (O_3295,N_49459,N_46482);
and UO_3296 (O_3296,N_45512,N_48758);
nor UO_3297 (O_3297,N_47195,N_47696);
xnor UO_3298 (O_3298,N_45700,N_49970);
and UO_3299 (O_3299,N_46637,N_46085);
or UO_3300 (O_3300,N_46063,N_47988);
and UO_3301 (O_3301,N_45170,N_45539);
xnor UO_3302 (O_3302,N_47278,N_49053);
xnor UO_3303 (O_3303,N_48541,N_45923);
or UO_3304 (O_3304,N_45083,N_49028);
and UO_3305 (O_3305,N_45335,N_48041);
or UO_3306 (O_3306,N_47642,N_46378);
and UO_3307 (O_3307,N_45692,N_48794);
or UO_3308 (O_3308,N_47167,N_49867);
nor UO_3309 (O_3309,N_49744,N_49977);
xnor UO_3310 (O_3310,N_49691,N_45368);
nand UO_3311 (O_3311,N_45295,N_46532);
nand UO_3312 (O_3312,N_47502,N_45259);
or UO_3313 (O_3313,N_48374,N_49186);
nor UO_3314 (O_3314,N_46269,N_47665);
and UO_3315 (O_3315,N_45784,N_48930);
nor UO_3316 (O_3316,N_45887,N_48061);
xnor UO_3317 (O_3317,N_47974,N_47606);
nor UO_3318 (O_3318,N_45006,N_45364);
xnor UO_3319 (O_3319,N_46070,N_45716);
or UO_3320 (O_3320,N_45656,N_49905);
xnor UO_3321 (O_3321,N_49006,N_45979);
nor UO_3322 (O_3322,N_45364,N_45368);
xor UO_3323 (O_3323,N_46585,N_45404);
and UO_3324 (O_3324,N_49599,N_47019);
nor UO_3325 (O_3325,N_49471,N_48539);
or UO_3326 (O_3326,N_47976,N_46515);
and UO_3327 (O_3327,N_49767,N_47625);
xnor UO_3328 (O_3328,N_48132,N_45821);
and UO_3329 (O_3329,N_48414,N_46593);
nand UO_3330 (O_3330,N_46468,N_46911);
nand UO_3331 (O_3331,N_45229,N_48320);
nor UO_3332 (O_3332,N_48745,N_47778);
nor UO_3333 (O_3333,N_48275,N_48010);
or UO_3334 (O_3334,N_46747,N_49385);
nand UO_3335 (O_3335,N_47456,N_49777);
xnor UO_3336 (O_3336,N_46513,N_46353);
or UO_3337 (O_3337,N_45561,N_49182);
nor UO_3338 (O_3338,N_45784,N_47804);
and UO_3339 (O_3339,N_46700,N_46893);
and UO_3340 (O_3340,N_45626,N_45775);
xnor UO_3341 (O_3341,N_48045,N_47091);
xnor UO_3342 (O_3342,N_48573,N_48154);
and UO_3343 (O_3343,N_49525,N_47298);
or UO_3344 (O_3344,N_45698,N_49840);
xor UO_3345 (O_3345,N_46436,N_45019);
nand UO_3346 (O_3346,N_45021,N_48155);
or UO_3347 (O_3347,N_48220,N_45020);
nand UO_3348 (O_3348,N_45084,N_45683);
or UO_3349 (O_3349,N_47944,N_48380);
or UO_3350 (O_3350,N_46032,N_49996);
and UO_3351 (O_3351,N_45093,N_45547);
or UO_3352 (O_3352,N_46146,N_49286);
xor UO_3353 (O_3353,N_45168,N_46802);
nand UO_3354 (O_3354,N_45828,N_49453);
and UO_3355 (O_3355,N_45615,N_45546);
nor UO_3356 (O_3356,N_47924,N_49963);
and UO_3357 (O_3357,N_48864,N_48639);
nand UO_3358 (O_3358,N_45657,N_45948);
nand UO_3359 (O_3359,N_46808,N_47445);
and UO_3360 (O_3360,N_45478,N_46090);
nand UO_3361 (O_3361,N_45395,N_47403);
nor UO_3362 (O_3362,N_47394,N_49370);
xor UO_3363 (O_3363,N_46606,N_47603);
nand UO_3364 (O_3364,N_46999,N_46443);
xnor UO_3365 (O_3365,N_49723,N_46857);
and UO_3366 (O_3366,N_49846,N_46548);
xor UO_3367 (O_3367,N_49515,N_49078);
nor UO_3368 (O_3368,N_49103,N_48940);
and UO_3369 (O_3369,N_47052,N_47545);
nor UO_3370 (O_3370,N_47574,N_48911);
and UO_3371 (O_3371,N_45095,N_45250);
nor UO_3372 (O_3372,N_49936,N_48263);
or UO_3373 (O_3373,N_48861,N_46909);
or UO_3374 (O_3374,N_46076,N_47127);
and UO_3375 (O_3375,N_46709,N_49372);
xnor UO_3376 (O_3376,N_45663,N_45779);
and UO_3377 (O_3377,N_45661,N_46713);
xnor UO_3378 (O_3378,N_46355,N_49110);
and UO_3379 (O_3379,N_47175,N_49751);
nand UO_3380 (O_3380,N_47414,N_48849);
xnor UO_3381 (O_3381,N_49743,N_48289);
xnor UO_3382 (O_3382,N_49820,N_46122);
or UO_3383 (O_3383,N_49191,N_47250);
xor UO_3384 (O_3384,N_45749,N_48434);
nor UO_3385 (O_3385,N_47916,N_45289);
nand UO_3386 (O_3386,N_47525,N_48586);
xnor UO_3387 (O_3387,N_47027,N_47877);
and UO_3388 (O_3388,N_46272,N_45229);
xor UO_3389 (O_3389,N_45923,N_49833);
and UO_3390 (O_3390,N_49126,N_48176);
or UO_3391 (O_3391,N_46662,N_45395);
and UO_3392 (O_3392,N_45228,N_47460);
and UO_3393 (O_3393,N_49422,N_48492);
and UO_3394 (O_3394,N_45758,N_47691);
or UO_3395 (O_3395,N_47781,N_46764);
xnor UO_3396 (O_3396,N_49354,N_45462);
xor UO_3397 (O_3397,N_47390,N_45437);
or UO_3398 (O_3398,N_47268,N_47101);
nor UO_3399 (O_3399,N_47716,N_45524);
and UO_3400 (O_3400,N_49202,N_49399);
nand UO_3401 (O_3401,N_48813,N_46073);
nand UO_3402 (O_3402,N_45898,N_49241);
xor UO_3403 (O_3403,N_47464,N_47935);
nor UO_3404 (O_3404,N_49623,N_47635);
nand UO_3405 (O_3405,N_45987,N_46512);
nand UO_3406 (O_3406,N_46386,N_46984);
xor UO_3407 (O_3407,N_48811,N_46044);
nor UO_3408 (O_3408,N_47000,N_48540);
xor UO_3409 (O_3409,N_45993,N_48277);
xnor UO_3410 (O_3410,N_49479,N_47857);
and UO_3411 (O_3411,N_49636,N_49871);
nand UO_3412 (O_3412,N_48497,N_46299);
and UO_3413 (O_3413,N_46918,N_47747);
xnor UO_3414 (O_3414,N_47641,N_46924);
nor UO_3415 (O_3415,N_45717,N_48490);
nand UO_3416 (O_3416,N_46792,N_45134);
or UO_3417 (O_3417,N_48805,N_47684);
and UO_3418 (O_3418,N_46143,N_47139);
nor UO_3419 (O_3419,N_46394,N_45560);
and UO_3420 (O_3420,N_45470,N_45859);
or UO_3421 (O_3421,N_49477,N_45670);
and UO_3422 (O_3422,N_46035,N_48347);
and UO_3423 (O_3423,N_45942,N_47957);
nor UO_3424 (O_3424,N_47094,N_49671);
nor UO_3425 (O_3425,N_48029,N_46160);
xor UO_3426 (O_3426,N_45249,N_46037);
xor UO_3427 (O_3427,N_48145,N_47197);
or UO_3428 (O_3428,N_47059,N_47332);
or UO_3429 (O_3429,N_48011,N_45864);
or UO_3430 (O_3430,N_46556,N_48126);
and UO_3431 (O_3431,N_49588,N_49015);
nor UO_3432 (O_3432,N_48525,N_48422);
nand UO_3433 (O_3433,N_48254,N_49682);
or UO_3434 (O_3434,N_47706,N_46746);
or UO_3435 (O_3435,N_48996,N_48151);
or UO_3436 (O_3436,N_46712,N_47997);
nand UO_3437 (O_3437,N_47501,N_45904);
nor UO_3438 (O_3438,N_45501,N_45509);
or UO_3439 (O_3439,N_47206,N_47035);
nor UO_3440 (O_3440,N_45615,N_49395);
and UO_3441 (O_3441,N_46164,N_49779);
nand UO_3442 (O_3442,N_45540,N_45828);
xor UO_3443 (O_3443,N_45361,N_48041);
nor UO_3444 (O_3444,N_47545,N_48420);
and UO_3445 (O_3445,N_49688,N_46976);
nor UO_3446 (O_3446,N_45970,N_46229);
xor UO_3447 (O_3447,N_46164,N_47514);
xnor UO_3448 (O_3448,N_48287,N_46007);
and UO_3449 (O_3449,N_48332,N_45469);
or UO_3450 (O_3450,N_48291,N_47755);
nand UO_3451 (O_3451,N_45103,N_48174);
nor UO_3452 (O_3452,N_48239,N_47646);
and UO_3453 (O_3453,N_47818,N_45614);
nand UO_3454 (O_3454,N_49833,N_46956);
and UO_3455 (O_3455,N_48648,N_46016);
nand UO_3456 (O_3456,N_46677,N_45330);
xor UO_3457 (O_3457,N_48273,N_46595);
and UO_3458 (O_3458,N_47049,N_47523);
xnor UO_3459 (O_3459,N_49993,N_47349);
nand UO_3460 (O_3460,N_47938,N_45427);
nor UO_3461 (O_3461,N_47699,N_47589);
or UO_3462 (O_3462,N_48397,N_49367);
or UO_3463 (O_3463,N_47647,N_45403);
or UO_3464 (O_3464,N_45283,N_46307);
and UO_3465 (O_3465,N_48416,N_47796);
or UO_3466 (O_3466,N_46957,N_48755);
nand UO_3467 (O_3467,N_47627,N_45996);
nand UO_3468 (O_3468,N_48096,N_49214);
nand UO_3469 (O_3469,N_49658,N_46556);
nand UO_3470 (O_3470,N_49084,N_45499);
nand UO_3471 (O_3471,N_49819,N_47423);
and UO_3472 (O_3472,N_47731,N_48802);
or UO_3473 (O_3473,N_47016,N_48946);
xnor UO_3474 (O_3474,N_49789,N_48253);
or UO_3475 (O_3475,N_45767,N_48047);
or UO_3476 (O_3476,N_45273,N_45224);
or UO_3477 (O_3477,N_47821,N_45283);
xnor UO_3478 (O_3478,N_47675,N_48521);
nand UO_3479 (O_3479,N_49658,N_45209);
or UO_3480 (O_3480,N_49120,N_47643);
nand UO_3481 (O_3481,N_48941,N_48317);
or UO_3482 (O_3482,N_46998,N_47182);
nand UO_3483 (O_3483,N_48771,N_45578);
or UO_3484 (O_3484,N_49804,N_46947);
xor UO_3485 (O_3485,N_47110,N_47866);
and UO_3486 (O_3486,N_47281,N_45831);
nor UO_3487 (O_3487,N_48689,N_47249);
nand UO_3488 (O_3488,N_46338,N_45283);
xnor UO_3489 (O_3489,N_49935,N_46234);
and UO_3490 (O_3490,N_48227,N_49522);
nand UO_3491 (O_3491,N_46115,N_45215);
nand UO_3492 (O_3492,N_45110,N_49916);
or UO_3493 (O_3493,N_48327,N_48552);
or UO_3494 (O_3494,N_46493,N_48307);
nor UO_3495 (O_3495,N_46863,N_48770);
nand UO_3496 (O_3496,N_49041,N_45325);
or UO_3497 (O_3497,N_48700,N_48490);
xnor UO_3498 (O_3498,N_49542,N_49414);
or UO_3499 (O_3499,N_46653,N_49640);
nor UO_3500 (O_3500,N_45085,N_47500);
nor UO_3501 (O_3501,N_45893,N_49708);
and UO_3502 (O_3502,N_46454,N_45110);
nor UO_3503 (O_3503,N_48005,N_47687);
or UO_3504 (O_3504,N_49892,N_48045);
nand UO_3505 (O_3505,N_47006,N_45383);
xnor UO_3506 (O_3506,N_46338,N_48439);
xnor UO_3507 (O_3507,N_45620,N_47627);
nor UO_3508 (O_3508,N_46176,N_49403);
and UO_3509 (O_3509,N_48443,N_47302);
or UO_3510 (O_3510,N_48237,N_49068);
and UO_3511 (O_3511,N_49535,N_49421);
nor UO_3512 (O_3512,N_48814,N_45154);
nor UO_3513 (O_3513,N_47251,N_49471);
nand UO_3514 (O_3514,N_49752,N_45255);
or UO_3515 (O_3515,N_48389,N_45904);
or UO_3516 (O_3516,N_48697,N_46524);
and UO_3517 (O_3517,N_48000,N_45073);
or UO_3518 (O_3518,N_49388,N_49118);
and UO_3519 (O_3519,N_45042,N_49032);
and UO_3520 (O_3520,N_46768,N_49065);
nor UO_3521 (O_3521,N_48537,N_48067);
xnor UO_3522 (O_3522,N_49134,N_47068);
nand UO_3523 (O_3523,N_46480,N_49182);
xor UO_3524 (O_3524,N_49562,N_48304);
and UO_3525 (O_3525,N_45537,N_46269);
nor UO_3526 (O_3526,N_46152,N_47317);
nor UO_3527 (O_3527,N_45706,N_47605);
and UO_3528 (O_3528,N_45936,N_49127);
nand UO_3529 (O_3529,N_48209,N_45444);
nor UO_3530 (O_3530,N_47880,N_48113);
nor UO_3531 (O_3531,N_45125,N_46923);
and UO_3532 (O_3532,N_45858,N_48194);
xnor UO_3533 (O_3533,N_46170,N_48611);
nand UO_3534 (O_3534,N_48541,N_46439);
xnor UO_3535 (O_3535,N_47958,N_47481);
nand UO_3536 (O_3536,N_49845,N_45523);
or UO_3537 (O_3537,N_47940,N_48347);
or UO_3538 (O_3538,N_47223,N_46561);
or UO_3539 (O_3539,N_47230,N_47664);
xnor UO_3540 (O_3540,N_46375,N_48055);
and UO_3541 (O_3541,N_49994,N_45524);
xnor UO_3542 (O_3542,N_46348,N_49321);
xnor UO_3543 (O_3543,N_48471,N_45181);
and UO_3544 (O_3544,N_45705,N_45406);
or UO_3545 (O_3545,N_46505,N_47069);
and UO_3546 (O_3546,N_46418,N_45927);
or UO_3547 (O_3547,N_47234,N_47152);
nand UO_3548 (O_3548,N_49584,N_48983);
xnor UO_3549 (O_3549,N_46681,N_46352);
nor UO_3550 (O_3550,N_48982,N_45143);
nand UO_3551 (O_3551,N_45257,N_46312);
nor UO_3552 (O_3552,N_45848,N_46786);
and UO_3553 (O_3553,N_46396,N_49785);
and UO_3554 (O_3554,N_46338,N_46633);
xnor UO_3555 (O_3555,N_45520,N_48741);
and UO_3556 (O_3556,N_48014,N_48401);
or UO_3557 (O_3557,N_49950,N_45259);
nor UO_3558 (O_3558,N_48575,N_49029);
and UO_3559 (O_3559,N_49548,N_49446);
xor UO_3560 (O_3560,N_48555,N_46637);
xor UO_3561 (O_3561,N_49846,N_48990);
or UO_3562 (O_3562,N_49336,N_46375);
and UO_3563 (O_3563,N_46918,N_47132);
nand UO_3564 (O_3564,N_46594,N_47978);
or UO_3565 (O_3565,N_49536,N_46454);
nor UO_3566 (O_3566,N_46392,N_45875);
nor UO_3567 (O_3567,N_48149,N_47662);
and UO_3568 (O_3568,N_49406,N_47022);
nor UO_3569 (O_3569,N_49940,N_49195);
nor UO_3570 (O_3570,N_45876,N_49981);
nor UO_3571 (O_3571,N_45391,N_45569);
and UO_3572 (O_3572,N_47533,N_49807);
nor UO_3573 (O_3573,N_47771,N_49603);
nor UO_3574 (O_3574,N_47992,N_49671);
nor UO_3575 (O_3575,N_49076,N_48123);
nand UO_3576 (O_3576,N_49173,N_45504);
nand UO_3577 (O_3577,N_46910,N_45670);
and UO_3578 (O_3578,N_46381,N_48251);
and UO_3579 (O_3579,N_48951,N_49637);
or UO_3580 (O_3580,N_46929,N_47107);
nand UO_3581 (O_3581,N_45289,N_45141);
or UO_3582 (O_3582,N_48368,N_46564);
nand UO_3583 (O_3583,N_49250,N_46127);
nand UO_3584 (O_3584,N_46848,N_45975);
nand UO_3585 (O_3585,N_48087,N_46512);
or UO_3586 (O_3586,N_49892,N_49534);
nand UO_3587 (O_3587,N_45302,N_45234);
nor UO_3588 (O_3588,N_49810,N_48269);
or UO_3589 (O_3589,N_48687,N_47977);
xnor UO_3590 (O_3590,N_49162,N_45871);
nor UO_3591 (O_3591,N_47998,N_46591);
nand UO_3592 (O_3592,N_46570,N_45486);
and UO_3593 (O_3593,N_46118,N_49419);
nor UO_3594 (O_3594,N_46352,N_45262);
and UO_3595 (O_3595,N_46839,N_46974);
xnor UO_3596 (O_3596,N_45905,N_49509);
or UO_3597 (O_3597,N_47917,N_46195);
or UO_3598 (O_3598,N_48120,N_47898);
xor UO_3599 (O_3599,N_48606,N_45270);
xor UO_3600 (O_3600,N_48336,N_47583);
nand UO_3601 (O_3601,N_46030,N_47263);
nor UO_3602 (O_3602,N_47047,N_47391);
and UO_3603 (O_3603,N_45913,N_47943);
nor UO_3604 (O_3604,N_46735,N_49493);
nor UO_3605 (O_3605,N_46262,N_47603);
nor UO_3606 (O_3606,N_49055,N_46550);
and UO_3607 (O_3607,N_48726,N_47723);
nand UO_3608 (O_3608,N_45798,N_48186);
xor UO_3609 (O_3609,N_47443,N_48212);
nand UO_3610 (O_3610,N_46864,N_47591);
xnor UO_3611 (O_3611,N_48501,N_46967);
and UO_3612 (O_3612,N_49136,N_45017);
xnor UO_3613 (O_3613,N_45597,N_45145);
nand UO_3614 (O_3614,N_46614,N_47858);
nand UO_3615 (O_3615,N_47551,N_45523);
nor UO_3616 (O_3616,N_48729,N_49017);
nor UO_3617 (O_3617,N_48658,N_45832);
or UO_3618 (O_3618,N_48661,N_46172);
or UO_3619 (O_3619,N_48997,N_46419);
xnor UO_3620 (O_3620,N_47911,N_49870);
nand UO_3621 (O_3621,N_48517,N_46592);
nor UO_3622 (O_3622,N_47969,N_46820);
xor UO_3623 (O_3623,N_48080,N_46805);
nor UO_3624 (O_3624,N_47632,N_46988);
xor UO_3625 (O_3625,N_46298,N_48557);
or UO_3626 (O_3626,N_47059,N_47318);
or UO_3627 (O_3627,N_48793,N_48345);
and UO_3628 (O_3628,N_46115,N_47998);
xor UO_3629 (O_3629,N_46861,N_48771);
xnor UO_3630 (O_3630,N_48196,N_45537);
or UO_3631 (O_3631,N_49678,N_46757);
and UO_3632 (O_3632,N_49841,N_47721);
and UO_3633 (O_3633,N_47533,N_45145);
nor UO_3634 (O_3634,N_47576,N_45226);
nor UO_3635 (O_3635,N_49283,N_47406);
nor UO_3636 (O_3636,N_45531,N_45555);
or UO_3637 (O_3637,N_48389,N_47265);
and UO_3638 (O_3638,N_49090,N_49380);
nor UO_3639 (O_3639,N_49070,N_47704);
and UO_3640 (O_3640,N_47077,N_45271);
nand UO_3641 (O_3641,N_45306,N_45576);
nand UO_3642 (O_3642,N_49639,N_45291);
or UO_3643 (O_3643,N_45936,N_48962);
nor UO_3644 (O_3644,N_46807,N_49353);
nand UO_3645 (O_3645,N_49909,N_46875);
nor UO_3646 (O_3646,N_49505,N_45278);
or UO_3647 (O_3647,N_45858,N_47206);
nor UO_3648 (O_3648,N_47492,N_49481);
and UO_3649 (O_3649,N_45305,N_48675);
or UO_3650 (O_3650,N_46720,N_46707);
nor UO_3651 (O_3651,N_46420,N_46525);
nand UO_3652 (O_3652,N_49818,N_49492);
nand UO_3653 (O_3653,N_47443,N_45865);
or UO_3654 (O_3654,N_49779,N_46776);
or UO_3655 (O_3655,N_49046,N_47441);
nand UO_3656 (O_3656,N_46277,N_45024);
and UO_3657 (O_3657,N_49402,N_45561);
nor UO_3658 (O_3658,N_46800,N_49511);
nor UO_3659 (O_3659,N_46790,N_49154);
xor UO_3660 (O_3660,N_46656,N_48419);
nand UO_3661 (O_3661,N_49539,N_47277);
nor UO_3662 (O_3662,N_49006,N_48842);
and UO_3663 (O_3663,N_45729,N_49812);
nand UO_3664 (O_3664,N_47850,N_45029);
nand UO_3665 (O_3665,N_47151,N_48586);
xnor UO_3666 (O_3666,N_47811,N_49244);
and UO_3667 (O_3667,N_45092,N_45585);
nand UO_3668 (O_3668,N_46451,N_45542);
and UO_3669 (O_3669,N_45425,N_48210);
xor UO_3670 (O_3670,N_49965,N_47094);
nand UO_3671 (O_3671,N_47709,N_45863);
or UO_3672 (O_3672,N_45904,N_47876);
or UO_3673 (O_3673,N_45833,N_45196);
or UO_3674 (O_3674,N_49759,N_49830);
and UO_3675 (O_3675,N_46184,N_46302);
or UO_3676 (O_3676,N_48940,N_49089);
nand UO_3677 (O_3677,N_47234,N_48815);
nand UO_3678 (O_3678,N_46759,N_46513);
and UO_3679 (O_3679,N_49082,N_46169);
and UO_3680 (O_3680,N_45197,N_46974);
xnor UO_3681 (O_3681,N_48455,N_45757);
or UO_3682 (O_3682,N_49978,N_45058);
nand UO_3683 (O_3683,N_49531,N_47029);
and UO_3684 (O_3684,N_46745,N_48990);
nor UO_3685 (O_3685,N_48988,N_48188);
and UO_3686 (O_3686,N_48449,N_49709);
or UO_3687 (O_3687,N_47076,N_46940);
nand UO_3688 (O_3688,N_49336,N_47849);
nand UO_3689 (O_3689,N_49440,N_47464);
and UO_3690 (O_3690,N_45265,N_46181);
nand UO_3691 (O_3691,N_45623,N_48063);
nor UO_3692 (O_3692,N_46870,N_47786);
nand UO_3693 (O_3693,N_49310,N_49799);
or UO_3694 (O_3694,N_45151,N_46628);
nor UO_3695 (O_3695,N_46312,N_46344);
or UO_3696 (O_3696,N_47738,N_49959);
and UO_3697 (O_3697,N_46168,N_49730);
nor UO_3698 (O_3698,N_46353,N_49335);
or UO_3699 (O_3699,N_49378,N_45264);
nand UO_3700 (O_3700,N_45116,N_48372);
or UO_3701 (O_3701,N_47179,N_46939);
nor UO_3702 (O_3702,N_49597,N_46296);
nand UO_3703 (O_3703,N_45237,N_45324);
and UO_3704 (O_3704,N_47063,N_49799);
nor UO_3705 (O_3705,N_47806,N_46253);
xnor UO_3706 (O_3706,N_49771,N_46919);
or UO_3707 (O_3707,N_48496,N_45402);
and UO_3708 (O_3708,N_46587,N_47974);
or UO_3709 (O_3709,N_46940,N_49277);
and UO_3710 (O_3710,N_49777,N_45696);
xor UO_3711 (O_3711,N_47697,N_45279);
or UO_3712 (O_3712,N_48025,N_45505);
and UO_3713 (O_3713,N_48553,N_45906);
and UO_3714 (O_3714,N_49467,N_47010);
or UO_3715 (O_3715,N_46433,N_49791);
or UO_3716 (O_3716,N_49023,N_45638);
nor UO_3717 (O_3717,N_49814,N_45432);
and UO_3718 (O_3718,N_49060,N_45713);
or UO_3719 (O_3719,N_49278,N_48929);
xor UO_3720 (O_3720,N_49758,N_47617);
nor UO_3721 (O_3721,N_46221,N_49546);
or UO_3722 (O_3722,N_49468,N_46277);
and UO_3723 (O_3723,N_49129,N_47956);
and UO_3724 (O_3724,N_45459,N_49155);
xor UO_3725 (O_3725,N_45050,N_47639);
xor UO_3726 (O_3726,N_49826,N_47186);
nand UO_3727 (O_3727,N_49611,N_45936);
nor UO_3728 (O_3728,N_48268,N_48647);
and UO_3729 (O_3729,N_45398,N_45468);
or UO_3730 (O_3730,N_45730,N_49075);
or UO_3731 (O_3731,N_47267,N_46572);
and UO_3732 (O_3732,N_45102,N_47215);
nor UO_3733 (O_3733,N_46255,N_45164);
and UO_3734 (O_3734,N_48331,N_48537);
or UO_3735 (O_3735,N_45101,N_47339);
xor UO_3736 (O_3736,N_48943,N_49645);
nand UO_3737 (O_3737,N_48408,N_48886);
nor UO_3738 (O_3738,N_47300,N_46390);
and UO_3739 (O_3739,N_46940,N_46698);
nor UO_3740 (O_3740,N_49470,N_47053);
or UO_3741 (O_3741,N_46527,N_47774);
or UO_3742 (O_3742,N_49431,N_48118);
nand UO_3743 (O_3743,N_48136,N_48108);
nand UO_3744 (O_3744,N_45794,N_49012);
xnor UO_3745 (O_3745,N_45118,N_49303);
or UO_3746 (O_3746,N_45598,N_49241);
nor UO_3747 (O_3747,N_48620,N_49355);
nand UO_3748 (O_3748,N_45966,N_48177);
or UO_3749 (O_3749,N_49704,N_45952);
nor UO_3750 (O_3750,N_45517,N_46528);
nor UO_3751 (O_3751,N_47766,N_49985);
nand UO_3752 (O_3752,N_46076,N_48111);
nor UO_3753 (O_3753,N_45185,N_49858);
nor UO_3754 (O_3754,N_47027,N_49434);
and UO_3755 (O_3755,N_47238,N_49981);
xor UO_3756 (O_3756,N_48241,N_48762);
or UO_3757 (O_3757,N_48673,N_47917);
nand UO_3758 (O_3758,N_45372,N_45493);
and UO_3759 (O_3759,N_48620,N_47408);
nor UO_3760 (O_3760,N_47056,N_48999);
and UO_3761 (O_3761,N_49277,N_46118);
nor UO_3762 (O_3762,N_47081,N_47858);
or UO_3763 (O_3763,N_48513,N_47375);
xnor UO_3764 (O_3764,N_46995,N_46161);
nor UO_3765 (O_3765,N_48085,N_46702);
nand UO_3766 (O_3766,N_48551,N_47100);
nor UO_3767 (O_3767,N_49494,N_47311);
nand UO_3768 (O_3768,N_49230,N_49000);
xor UO_3769 (O_3769,N_46668,N_47359);
xnor UO_3770 (O_3770,N_48201,N_46356);
and UO_3771 (O_3771,N_47546,N_46300);
and UO_3772 (O_3772,N_45262,N_45597);
or UO_3773 (O_3773,N_45180,N_47689);
xnor UO_3774 (O_3774,N_48344,N_48069);
xnor UO_3775 (O_3775,N_45850,N_45899);
and UO_3776 (O_3776,N_46564,N_46672);
or UO_3777 (O_3777,N_46379,N_45597);
and UO_3778 (O_3778,N_47474,N_45993);
nor UO_3779 (O_3779,N_48735,N_45043);
and UO_3780 (O_3780,N_45777,N_45539);
xor UO_3781 (O_3781,N_46062,N_49966);
or UO_3782 (O_3782,N_49433,N_45073);
xor UO_3783 (O_3783,N_46449,N_46317);
nor UO_3784 (O_3784,N_49141,N_46416);
xor UO_3785 (O_3785,N_47809,N_46278);
or UO_3786 (O_3786,N_47917,N_49689);
and UO_3787 (O_3787,N_48831,N_46686);
nor UO_3788 (O_3788,N_48081,N_46628);
and UO_3789 (O_3789,N_46589,N_49033);
xnor UO_3790 (O_3790,N_46386,N_46579);
nor UO_3791 (O_3791,N_48276,N_45718);
nor UO_3792 (O_3792,N_46471,N_46534);
or UO_3793 (O_3793,N_46576,N_47946);
nor UO_3794 (O_3794,N_45590,N_48427);
and UO_3795 (O_3795,N_48816,N_46608);
xnor UO_3796 (O_3796,N_46426,N_46616);
nand UO_3797 (O_3797,N_46680,N_46998);
nor UO_3798 (O_3798,N_45510,N_46983);
xor UO_3799 (O_3799,N_47635,N_45436);
xnor UO_3800 (O_3800,N_49195,N_49620);
nand UO_3801 (O_3801,N_49136,N_47753);
xnor UO_3802 (O_3802,N_48908,N_48799);
xnor UO_3803 (O_3803,N_46704,N_45189);
nor UO_3804 (O_3804,N_46898,N_47071);
nand UO_3805 (O_3805,N_48403,N_49794);
and UO_3806 (O_3806,N_47202,N_45681);
nand UO_3807 (O_3807,N_49033,N_46855);
xnor UO_3808 (O_3808,N_47851,N_45761);
nor UO_3809 (O_3809,N_45777,N_47116);
or UO_3810 (O_3810,N_47064,N_46080);
and UO_3811 (O_3811,N_47915,N_48501);
nand UO_3812 (O_3812,N_48060,N_48161);
or UO_3813 (O_3813,N_45514,N_45564);
xnor UO_3814 (O_3814,N_49268,N_46149);
or UO_3815 (O_3815,N_48976,N_48036);
nor UO_3816 (O_3816,N_47803,N_45342);
and UO_3817 (O_3817,N_49935,N_47016);
or UO_3818 (O_3818,N_46269,N_45024);
nand UO_3819 (O_3819,N_49762,N_45863);
xnor UO_3820 (O_3820,N_45956,N_47041);
xnor UO_3821 (O_3821,N_46549,N_47314);
xor UO_3822 (O_3822,N_45244,N_48010);
and UO_3823 (O_3823,N_47687,N_45062);
xnor UO_3824 (O_3824,N_47348,N_45675);
nand UO_3825 (O_3825,N_45807,N_48504);
nand UO_3826 (O_3826,N_46731,N_45519);
nand UO_3827 (O_3827,N_46401,N_45988);
xor UO_3828 (O_3828,N_47087,N_48010);
xnor UO_3829 (O_3829,N_47056,N_48910);
xnor UO_3830 (O_3830,N_46418,N_48770);
xor UO_3831 (O_3831,N_45868,N_45067);
nand UO_3832 (O_3832,N_46932,N_49966);
and UO_3833 (O_3833,N_45749,N_47903);
or UO_3834 (O_3834,N_45822,N_49993);
and UO_3835 (O_3835,N_47238,N_49776);
xnor UO_3836 (O_3836,N_47774,N_46684);
nand UO_3837 (O_3837,N_46795,N_49587);
nand UO_3838 (O_3838,N_45346,N_46839);
nand UO_3839 (O_3839,N_47142,N_47748);
xnor UO_3840 (O_3840,N_46630,N_45704);
nand UO_3841 (O_3841,N_47133,N_47587);
nand UO_3842 (O_3842,N_45871,N_49847);
and UO_3843 (O_3843,N_47345,N_49555);
nand UO_3844 (O_3844,N_47919,N_45534);
nor UO_3845 (O_3845,N_45707,N_49794);
nand UO_3846 (O_3846,N_48976,N_48285);
or UO_3847 (O_3847,N_46164,N_46613);
nor UO_3848 (O_3848,N_46215,N_47866);
nand UO_3849 (O_3849,N_49393,N_46294);
nor UO_3850 (O_3850,N_48090,N_47113);
and UO_3851 (O_3851,N_45261,N_48789);
nand UO_3852 (O_3852,N_45062,N_49273);
or UO_3853 (O_3853,N_46335,N_46872);
or UO_3854 (O_3854,N_47676,N_47336);
and UO_3855 (O_3855,N_48201,N_47550);
nand UO_3856 (O_3856,N_48775,N_48150);
or UO_3857 (O_3857,N_47782,N_49669);
or UO_3858 (O_3858,N_46413,N_48457);
nor UO_3859 (O_3859,N_45693,N_46822);
nand UO_3860 (O_3860,N_49043,N_46672);
nor UO_3861 (O_3861,N_49140,N_47353);
and UO_3862 (O_3862,N_48366,N_48194);
nor UO_3863 (O_3863,N_49175,N_46841);
and UO_3864 (O_3864,N_45108,N_49789);
xor UO_3865 (O_3865,N_45254,N_49430);
xor UO_3866 (O_3866,N_49177,N_49128);
and UO_3867 (O_3867,N_48228,N_49095);
xnor UO_3868 (O_3868,N_46846,N_48923);
or UO_3869 (O_3869,N_48263,N_46124);
and UO_3870 (O_3870,N_45980,N_45935);
nor UO_3871 (O_3871,N_46199,N_46795);
xor UO_3872 (O_3872,N_49157,N_46770);
nand UO_3873 (O_3873,N_46913,N_46648);
nand UO_3874 (O_3874,N_45584,N_47449);
or UO_3875 (O_3875,N_47249,N_45235);
nor UO_3876 (O_3876,N_46296,N_47904);
nor UO_3877 (O_3877,N_48512,N_47775);
and UO_3878 (O_3878,N_45307,N_47471);
nand UO_3879 (O_3879,N_46449,N_48102);
nand UO_3880 (O_3880,N_47195,N_45713);
nand UO_3881 (O_3881,N_47049,N_48777);
and UO_3882 (O_3882,N_48202,N_49506);
nor UO_3883 (O_3883,N_45723,N_46064);
or UO_3884 (O_3884,N_45979,N_45720);
or UO_3885 (O_3885,N_49616,N_49874);
and UO_3886 (O_3886,N_48071,N_45898);
and UO_3887 (O_3887,N_46501,N_48774);
and UO_3888 (O_3888,N_46674,N_47615);
xor UO_3889 (O_3889,N_45098,N_49186);
nand UO_3890 (O_3890,N_49897,N_49040);
or UO_3891 (O_3891,N_45928,N_46221);
nor UO_3892 (O_3892,N_46665,N_47945);
and UO_3893 (O_3893,N_49501,N_46453);
or UO_3894 (O_3894,N_46528,N_47629);
or UO_3895 (O_3895,N_47700,N_48507);
nand UO_3896 (O_3896,N_48309,N_46798);
and UO_3897 (O_3897,N_47553,N_45513);
and UO_3898 (O_3898,N_46214,N_46384);
xnor UO_3899 (O_3899,N_49215,N_49121);
nand UO_3900 (O_3900,N_47801,N_46227);
or UO_3901 (O_3901,N_49816,N_47948);
xor UO_3902 (O_3902,N_46456,N_47424);
and UO_3903 (O_3903,N_47831,N_45971);
xor UO_3904 (O_3904,N_48367,N_47127);
nor UO_3905 (O_3905,N_46317,N_47852);
nor UO_3906 (O_3906,N_49684,N_46872);
nand UO_3907 (O_3907,N_49841,N_47882);
and UO_3908 (O_3908,N_46423,N_47658);
and UO_3909 (O_3909,N_45863,N_45818);
nand UO_3910 (O_3910,N_48907,N_47168);
nand UO_3911 (O_3911,N_49406,N_48314);
nor UO_3912 (O_3912,N_46199,N_47406);
and UO_3913 (O_3913,N_47755,N_46616);
xor UO_3914 (O_3914,N_45136,N_46327);
or UO_3915 (O_3915,N_49089,N_46876);
nor UO_3916 (O_3916,N_49309,N_46309);
xnor UO_3917 (O_3917,N_47804,N_45485);
nor UO_3918 (O_3918,N_47835,N_49697);
or UO_3919 (O_3919,N_48619,N_47921);
xor UO_3920 (O_3920,N_47080,N_46454);
nor UO_3921 (O_3921,N_48303,N_49538);
xnor UO_3922 (O_3922,N_49176,N_47146);
nand UO_3923 (O_3923,N_48447,N_47565);
nor UO_3924 (O_3924,N_45934,N_48452);
nand UO_3925 (O_3925,N_49552,N_49187);
nand UO_3926 (O_3926,N_49213,N_45093);
and UO_3927 (O_3927,N_47860,N_46835);
xnor UO_3928 (O_3928,N_46098,N_48168);
xnor UO_3929 (O_3929,N_49551,N_45888);
nor UO_3930 (O_3930,N_48585,N_48064);
or UO_3931 (O_3931,N_49258,N_49433);
nor UO_3932 (O_3932,N_47798,N_49748);
xnor UO_3933 (O_3933,N_49372,N_49040);
or UO_3934 (O_3934,N_46891,N_48609);
or UO_3935 (O_3935,N_47144,N_47498);
or UO_3936 (O_3936,N_48847,N_49131);
nor UO_3937 (O_3937,N_48046,N_48923);
and UO_3938 (O_3938,N_46934,N_46606);
nand UO_3939 (O_3939,N_46247,N_46193);
or UO_3940 (O_3940,N_47829,N_46464);
nor UO_3941 (O_3941,N_46637,N_47577);
xor UO_3942 (O_3942,N_45380,N_47774);
nand UO_3943 (O_3943,N_46154,N_48948);
nor UO_3944 (O_3944,N_47850,N_49601);
or UO_3945 (O_3945,N_46538,N_46697);
xnor UO_3946 (O_3946,N_46816,N_49295);
and UO_3947 (O_3947,N_46740,N_45660);
xnor UO_3948 (O_3948,N_49396,N_45359);
or UO_3949 (O_3949,N_49044,N_46393);
nand UO_3950 (O_3950,N_47123,N_46221);
nand UO_3951 (O_3951,N_46261,N_48541);
xor UO_3952 (O_3952,N_48274,N_47881);
nand UO_3953 (O_3953,N_46920,N_47973);
nand UO_3954 (O_3954,N_46391,N_48735);
and UO_3955 (O_3955,N_48953,N_49279);
or UO_3956 (O_3956,N_49812,N_49612);
and UO_3957 (O_3957,N_47157,N_47465);
xor UO_3958 (O_3958,N_48870,N_47949);
and UO_3959 (O_3959,N_46153,N_49491);
nor UO_3960 (O_3960,N_48552,N_47431);
nor UO_3961 (O_3961,N_48375,N_47386);
nand UO_3962 (O_3962,N_45494,N_47127);
or UO_3963 (O_3963,N_48304,N_49096);
and UO_3964 (O_3964,N_48022,N_46383);
and UO_3965 (O_3965,N_49481,N_45290);
nand UO_3966 (O_3966,N_47088,N_47769);
or UO_3967 (O_3967,N_47277,N_48261);
xnor UO_3968 (O_3968,N_48041,N_46645);
xor UO_3969 (O_3969,N_45574,N_46962);
and UO_3970 (O_3970,N_45074,N_45735);
nand UO_3971 (O_3971,N_48290,N_45958);
xnor UO_3972 (O_3972,N_46729,N_46422);
or UO_3973 (O_3973,N_46129,N_48726);
nor UO_3974 (O_3974,N_49992,N_46546);
or UO_3975 (O_3975,N_48761,N_46944);
or UO_3976 (O_3976,N_47934,N_46414);
nand UO_3977 (O_3977,N_45700,N_48083);
nand UO_3978 (O_3978,N_48566,N_45163);
xor UO_3979 (O_3979,N_46109,N_49542);
nor UO_3980 (O_3980,N_45400,N_47391);
nor UO_3981 (O_3981,N_45446,N_46301);
or UO_3982 (O_3982,N_49050,N_46605);
nand UO_3983 (O_3983,N_49701,N_45246);
and UO_3984 (O_3984,N_49946,N_47510);
xor UO_3985 (O_3985,N_47552,N_48648);
and UO_3986 (O_3986,N_47709,N_49591);
and UO_3987 (O_3987,N_47934,N_48559);
nand UO_3988 (O_3988,N_47047,N_47238);
or UO_3989 (O_3989,N_49934,N_48161);
nand UO_3990 (O_3990,N_45250,N_46462);
or UO_3991 (O_3991,N_46364,N_47110);
xnor UO_3992 (O_3992,N_45190,N_49929);
or UO_3993 (O_3993,N_49863,N_49737);
and UO_3994 (O_3994,N_47812,N_47480);
or UO_3995 (O_3995,N_48497,N_49031);
or UO_3996 (O_3996,N_49620,N_47504);
nor UO_3997 (O_3997,N_46203,N_46933);
nand UO_3998 (O_3998,N_45939,N_49797);
or UO_3999 (O_3999,N_47544,N_48182);
nor UO_4000 (O_4000,N_46140,N_45226);
and UO_4001 (O_4001,N_46406,N_46884);
xor UO_4002 (O_4002,N_49997,N_48377);
xnor UO_4003 (O_4003,N_46705,N_48623);
nor UO_4004 (O_4004,N_49714,N_47838);
xor UO_4005 (O_4005,N_46353,N_47172);
nor UO_4006 (O_4006,N_48832,N_46470);
nand UO_4007 (O_4007,N_48040,N_49937);
nand UO_4008 (O_4008,N_48460,N_47518);
xnor UO_4009 (O_4009,N_47204,N_46939);
nand UO_4010 (O_4010,N_49037,N_45084);
nand UO_4011 (O_4011,N_49091,N_49577);
nor UO_4012 (O_4012,N_47838,N_49434);
xor UO_4013 (O_4013,N_48624,N_47037);
nand UO_4014 (O_4014,N_49097,N_49304);
xnor UO_4015 (O_4015,N_45555,N_46967);
or UO_4016 (O_4016,N_47912,N_46383);
nor UO_4017 (O_4017,N_48413,N_49997);
or UO_4018 (O_4018,N_47425,N_48164);
nand UO_4019 (O_4019,N_49184,N_45757);
nor UO_4020 (O_4020,N_45370,N_47159);
or UO_4021 (O_4021,N_47786,N_48819);
nand UO_4022 (O_4022,N_45004,N_45299);
nor UO_4023 (O_4023,N_47634,N_48322);
or UO_4024 (O_4024,N_46784,N_46483);
xnor UO_4025 (O_4025,N_47882,N_48598);
and UO_4026 (O_4026,N_47817,N_47993);
nand UO_4027 (O_4027,N_46639,N_45266);
nand UO_4028 (O_4028,N_49819,N_47233);
nor UO_4029 (O_4029,N_48856,N_49958);
or UO_4030 (O_4030,N_47326,N_49509);
and UO_4031 (O_4031,N_46387,N_49786);
nand UO_4032 (O_4032,N_46796,N_49453);
and UO_4033 (O_4033,N_46003,N_46771);
xnor UO_4034 (O_4034,N_49039,N_46983);
and UO_4035 (O_4035,N_48656,N_45574);
nand UO_4036 (O_4036,N_49633,N_47835);
or UO_4037 (O_4037,N_48187,N_45135);
xnor UO_4038 (O_4038,N_47321,N_48822);
and UO_4039 (O_4039,N_47884,N_49001);
or UO_4040 (O_4040,N_48919,N_49388);
nand UO_4041 (O_4041,N_49272,N_49420);
nor UO_4042 (O_4042,N_46513,N_47605);
nor UO_4043 (O_4043,N_48962,N_48180);
nor UO_4044 (O_4044,N_47418,N_46029);
nand UO_4045 (O_4045,N_48306,N_48087);
and UO_4046 (O_4046,N_47199,N_45412);
or UO_4047 (O_4047,N_46321,N_47595);
xnor UO_4048 (O_4048,N_47766,N_46599);
nand UO_4049 (O_4049,N_46691,N_45976);
nand UO_4050 (O_4050,N_45090,N_45827);
nor UO_4051 (O_4051,N_49828,N_46858);
nand UO_4052 (O_4052,N_47380,N_45484);
and UO_4053 (O_4053,N_47608,N_45744);
nor UO_4054 (O_4054,N_48014,N_47802);
nor UO_4055 (O_4055,N_46868,N_48567);
xnor UO_4056 (O_4056,N_48072,N_45250);
nand UO_4057 (O_4057,N_45225,N_48757);
xnor UO_4058 (O_4058,N_48140,N_48300);
or UO_4059 (O_4059,N_47259,N_48459);
nor UO_4060 (O_4060,N_47469,N_46067);
nor UO_4061 (O_4061,N_47307,N_48126);
and UO_4062 (O_4062,N_46512,N_47905);
nand UO_4063 (O_4063,N_45678,N_46376);
or UO_4064 (O_4064,N_45021,N_47551);
nor UO_4065 (O_4065,N_46468,N_48136);
and UO_4066 (O_4066,N_45620,N_46128);
nand UO_4067 (O_4067,N_47628,N_49982);
nand UO_4068 (O_4068,N_48797,N_45103);
xor UO_4069 (O_4069,N_45315,N_46047);
and UO_4070 (O_4070,N_47271,N_48398);
and UO_4071 (O_4071,N_48505,N_49575);
or UO_4072 (O_4072,N_49390,N_48762);
nor UO_4073 (O_4073,N_45342,N_47040);
nand UO_4074 (O_4074,N_48540,N_45848);
and UO_4075 (O_4075,N_45675,N_48940);
or UO_4076 (O_4076,N_45871,N_46208);
and UO_4077 (O_4077,N_47516,N_49613);
xor UO_4078 (O_4078,N_45986,N_47923);
nor UO_4079 (O_4079,N_49461,N_45988);
xnor UO_4080 (O_4080,N_47658,N_49107);
and UO_4081 (O_4081,N_47855,N_45170);
or UO_4082 (O_4082,N_49302,N_49445);
nor UO_4083 (O_4083,N_49887,N_49284);
and UO_4084 (O_4084,N_49860,N_48477);
nor UO_4085 (O_4085,N_48111,N_47736);
xor UO_4086 (O_4086,N_45604,N_49435);
nand UO_4087 (O_4087,N_46037,N_46454);
xnor UO_4088 (O_4088,N_45971,N_48420);
xnor UO_4089 (O_4089,N_46016,N_48080);
nand UO_4090 (O_4090,N_46515,N_48034);
and UO_4091 (O_4091,N_49259,N_48819);
or UO_4092 (O_4092,N_48361,N_49775);
xnor UO_4093 (O_4093,N_49709,N_48111);
and UO_4094 (O_4094,N_46126,N_45402);
nand UO_4095 (O_4095,N_45393,N_47661);
or UO_4096 (O_4096,N_48067,N_49670);
nand UO_4097 (O_4097,N_46134,N_47338);
nor UO_4098 (O_4098,N_46240,N_47609);
and UO_4099 (O_4099,N_46854,N_49889);
nand UO_4100 (O_4100,N_49309,N_49637);
or UO_4101 (O_4101,N_45011,N_45031);
or UO_4102 (O_4102,N_47641,N_46592);
nor UO_4103 (O_4103,N_49018,N_47330);
nand UO_4104 (O_4104,N_49123,N_47238);
xor UO_4105 (O_4105,N_48561,N_45922);
and UO_4106 (O_4106,N_47699,N_48916);
nand UO_4107 (O_4107,N_48718,N_45345);
xor UO_4108 (O_4108,N_46592,N_45525);
and UO_4109 (O_4109,N_45154,N_47451);
xor UO_4110 (O_4110,N_48072,N_49115);
or UO_4111 (O_4111,N_46170,N_46722);
xor UO_4112 (O_4112,N_46843,N_45723);
and UO_4113 (O_4113,N_45170,N_46768);
nor UO_4114 (O_4114,N_48719,N_45053);
or UO_4115 (O_4115,N_46395,N_49507);
nand UO_4116 (O_4116,N_47363,N_46648);
nand UO_4117 (O_4117,N_49625,N_48103);
nand UO_4118 (O_4118,N_46970,N_46687);
nor UO_4119 (O_4119,N_49556,N_47776);
nand UO_4120 (O_4120,N_46115,N_47764);
and UO_4121 (O_4121,N_46489,N_48869);
nor UO_4122 (O_4122,N_47065,N_47448);
nand UO_4123 (O_4123,N_48355,N_49565);
xor UO_4124 (O_4124,N_47239,N_48820);
or UO_4125 (O_4125,N_46537,N_46211);
or UO_4126 (O_4126,N_45798,N_47230);
or UO_4127 (O_4127,N_45647,N_46951);
or UO_4128 (O_4128,N_49781,N_47329);
and UO_4129 (O_4129,N_46938,N_47117);
nor UO_4130 (O_4130,N_45143,N_48838);
nor UO_4131 (O_4131,N_47528,N_47802);
or UO_4132 (O_4132,N_47078,N_47679);
or UO_4133 (O_4133,N_48770,N_45811);
xor UO_4134 (O_4134,N_45577,N_47592);
nor UO_4135 (O_4135,N_46138,N_47689);
nand UO_4136 (O_4136,N_49661,N_47552);
and UO_4137 (O_4137,N_48975,N_49530);
nand UO_4138 (O_4138,N_45347,N_45805);
nand UO_4139 (O_4139,N_47110,N_46203);
nor UO_4140 (O_4140,N_46897,N_48375);
nor UO_4141 (O_4141,N_46061,N_49194);
nor UO_4142 (O_4142,N_48185,N_46887);
nand UO_4143 (O_4143,N_47100,N_45937);
or UO_4144 (O_4144,N_46480,N_46753);
nor UO_4145 (O_4145,N_45498,N_45150);
xnor UO_4146 (O_4146,N_45356,N_48081);
and UO_4147 (O_4147,N_47129,N_49201);
xor UO_4148 (O_4148,N_49600,N_46410);
xor UO_4149 (O_4149,N_45327,N_48430);
nand UO_4150 (O_4150,N_48843,N_47904);
xnor UO_4151 (O_4151,N_46756,N_48037);
nor UO_4152 (O_4152,N_45805,N_47830);
and UO_4153 (O_4153,N_48193,N_45255);
and UO_4154 (O_4154,N_45934,N_45904);
nand UO_4155 (O_4155,N_45578,N_45631);
nor UO_4156 (O_4156,N_48027,N_49808);
or UO_4157 (O_4157,N_49773,N_47418);
nand UO_4158 (O_4158,N_47489,N_49251);
or UO_4159 (O_4159,N_45273,N_47935);
nand UO_4160 (O_4160,N_46834,N_49071);
and UO_4161 (O_4161,N_45884,N_45916);
nor UO_4162 (O_4162,N_47890,N_46514);
xnor UO_4163 (O_4163,N_49451,N_46427);
nand UO_4164 (O_4164,N_45461,N_47063);
or UO_4165 (O_4165,N_45595,N_47582);
xnor UO_4166 (O_4166,N_47709,N_45966);
nor UO_4167 (O_4167,N_45808,N_48085);
nand UO_4168 (O_4168,N_46829,N_46523);
and UO_4169 (O_4169,N_46718,N_48848);
or UO_4170 (O_4170,N_48834,N_47237);
nand UO_4171 (O_4171,N_47348,N_48819);
or UO_4172 (O_4172,N_49535,N_48208);
nor UO_4173 (O_4173,N_46020,N_47987);
nor UO_4174 (O_4174,N_49738,N_47283);
xnor UO_4175 (O_4175,N_49410,N_49091);
or UO_4176 (O_4176,N_47552,N_45002);
and UO_4177 (O_4177,N_45201,N_46504);
and UO_4178 (O_4178,N_48701,N_45510);
nand UO_4179 (O_4179,N_45424,N_46623);
and UO_4180 (O_4180,N_46828,N_49945);
xnor UO_4181 (O_4181,N_45473,N_48546);
nand UO_4182 (O_4182,N_48495,N_48677);
xnor UO_4183 (O_4183,N_49206,N_48521);
nand UO_4184 (O_4184,N_45173,N_47367);
and UO_4185 (O_4185,N_49961,N_45750);
xnor UO_4186 (O_4186,N_45928,N_49191);
and UO_4187 (O_4187,N_45943,N_49087);
or UO_4188 (O_4188,N_45327,N_47612);
or UO_4189 (O_4189,N_45879,N_47157);
xnor UO_4190 (O_4190,N_45826,N_49474);
and UO_4191 (O_4191,N_46822,N_48765);
and UO_4192 (O_4192,N_45641,N_48392);
and UO_4193 (O_4193,N_48520,N_48760);
nor UO_4194 (O_4194,N_47394,N_48999);
or UO_4195 (O_4195,N_46522,N_49012);
nand UO_4196 (O_4196,N_46667,N_49998);
nor UO_4197 (O_4197,N_48611,N_47622);
nand UO_4198 (O_4198,N_47949,N_47456);
nor UO_4199 (O_4199,N_48036,N_47836);
xor UO_4200 (O_4200,N_49892,N_46532);
and UO_4201 (O_4201,N_47469,N_47384);
or UO_4202 (O_4202,N_49103,N_46098);
or UO_4203 (O_4203,N_46979,N_45066);
or UO_4204 (O_4204,N_47630,N_49481);
and UO_4205 (O_4205,N_48058,N_46240);
nand UO_4206 (O_4206,N_49865,N_48162);
xor UO_4207 (O_4207,N_47776,N_45383);
nand UO_4208 (O_4208,N_49691,N_46720);
nand UO_4209 (O_4209,N_46054,N_48668);
nor UO_4210 (O_4210,N_46962,N_46031);
or UO_4211 (O_4211,N_49733,N_48925);
nor UO_4212 (O_4212,N_48365,N_46824);
and UO_4213 (O_4213,N_49405,N_46648);
and UO_4214 (O_4214,N_46931,N_48214);
or UO_4215 (O_4215,N_48716,N_49795);
nand UO_4216 (O_4216,N_47008,N_45863);
nor UO_4217 (O_4217,N_47483,N_46277);
xor UO_4218 (O_4218,N_46993,N_45664);
or UO_4219 (O_4219,N_45350,N_45568);
nor UO_4220 (O_4220,N_45561,N_48288);
nand UO_4221 (O_4221,N_46363,N_47723);
and UO_4222 (O_4222,N_45931,N_46369);
and UO_4223 (O_4223,N_49773,N_49541);
nand UO_4224 (O_4224,N_49234,N_46712);
or UO_4225 (O_4225,N_48371,N_47373);
xor UO_4226 (O_4226,N_46389,N_46450);
xor UO_4227 (O_4227,N_48127,N_49443);
and UO_4228 (O_4228,N_47921,N_45126);
nor UO_4229 (O_4229,N_46875,N_49786);
nor UO_4230 (O_4230,N_49297,N_49833);
nand UO_4231 (O_4231,N_46061,N_45148);
or UO_4232 (O_4232,N_45762,N_46283);
nand UO_4233 (O_4233,N_45321,N_47479);
xnor UO_4234 (O_4234,N_45143,N_46069);
nor UO_4235 (O_4235,N_48920,N_45096);
and UO_4236 (O_4236,N_45336,N_46970);
nand UO_4237 (O_4237,N_47564,N_48443);
xnor UO_4238 (O_4238,N_47484,N_46385);
nand UO_4239 (O_4239,N_47374,N_47791);
and UO_4240 (O_4240,N_46198,N_47479);
or UO_4241 (O_4241,N_48924,N_48386);
nor UO_4242 (O_4242,N_45905,N_46635);
nor UO_4243 (O_4243,N_46539,N_46301);
or UO_4244 (O_4244,N_45704,N_47488);
nor UO_4245 (O_4245,N_48496,N_47019);
nor UO_4246 (O_4246,N_48062,N_49480);
xnor UO_4247 (O_4247,N_47792,N_45535);
xor UO_4248 (O_4248,N_46753,N_48152);
nand UO_4249 (O_4249,N_48135,N_48944);
nand UO_4250 (O_4250,N_47083,N_47055);
xnor UO_4251 (O_4251,N_49712,N_49695);
nand UO_4252 (O_4252,N_47468,N_45343);
nor UO_4253 (O_4253,N_49477,N_45110);
xor UO_4254 (O_4254,N_48673,N_47140);
nor UO_4255 (O_4255,N_46480,N_49526);
nor UO_4256 (O_4256,N_45946,N_48052);
xor UO_4257 (O_4257,N_48811,N_45416);
or UO_4258 (O_4258,N_47315,N_45908);
and UO_4259 (O_4259,N_48681,N_46682);
or UO_4260 (O_4260,N_47418,N_45178);
nand UO_4261 (O_4261,N_49223,N_46847);
nor UO_4262 (O_4262,N_49169,N_46282);
and UO_4263 (O_4263,N_45924,N_48613);
and UO_4264 (O_4264,N_48357,N_47186);
nor UO_4265 (O_4265,N_47151,N_45303);
nand UO_4266 (O_4266,N_49379,N_49114);
xor UO_4267 (O_4267,N_45374,N_46236);
xor UO_4268 (O_4268,N_48663,N_46612);
and UO_4269 (O_4269,N_46001,N_45972);
nor UO_4270 (O_4270,N_49147,N_45843);
or UO_4271 (O_4271,N_47250,N_46390);
xnor UO_4272 (O_4272,N_48015,N_47296);
xor UO_4273 (O_4273,N_46165,N_46779);
nor UO_4274 (O_4274,N_49010,N_48666);
xor UO_4275 (O_4275,N_48728,N_49178);
and UO_4276 (O_4276,N_45084,N_45645);
or UO_4277 (O_4277,N_46786,N_46052);
xor UO_4278 (O_4278,N_46499,N_49288);
nand UO_4279 (O_4279,N_46059,N_49414);
nand UO_4280 (O_4280,N_47921,N_45968);
nand UO_4281 (O_4281,N_46431,N_49400);
xnor UO_4282 (O_4282,N_46717,N_49643);
xor UO_4283 (O_4283,N_49590,N_48200);
xnor UO_4284 (O_4284,N_48199,N_49418);
or UO_4285 (O_4285,N_46998,N_45448);
nor UO_4286 (O_4286,N_45216,N_46879);
nand UO_4287 (O_4287,N_46347,N_46829);
xnor UO_4288 (O_4288,N_46808,N_45922);
or UO_4289 (O_4289,N_46263,N_47811);
and UO_4290 (O_4290,N_45969,N_49754);
nand UO_4291 (O_4291,N_49698,N_49561);
xnor UO_4292 (O_4292,N_45920,N_46450);
nor UO_4293 (O_4293,N_49383,N_49563);
and UO_4294 (O_4294,N_49771,N_49734);
xor UO_4295 (O_4295,N_46779,N_49805);
or UO_4296 (O_4296,N_48251,N_48642);
nand UO_4297 (O_4297,N_48629,N_45704);
nor UO_4298 (O_4298,N_45892,N_46016);
nor UO_4299 (O_4299,N_45985,N_47098);
or UO_4300 (O_4300,N_47271,N_48539);
xor UO_4301 (O_4301,N_47962,N_49109);
nor UO_4302 (O_4302,N_47894,N_47739);
nor UO_4303 (O_4303,N_49066,N_47016);
and UO_4304 (O_4304,N_47347,N_46715);
nand UO_4305 (O_4305,N_45856,N_46550);
xor UO_4306 (O_4306,N_45697,N_45031);
or UO_4307 (O_4307,N_47959,N_49779);
nor UO_4308 (O_4308,N_45387,N_47410);
xnor UO_4309 (O_4309,N_49311,N_46758);
or UO_4310 (O_4310,N_46361,N_47176);
nand UO_4311 (O_4311,N_47892,N_47186);
and UO_4312 (O_4312,N_49314,N_47408);
nand UO_4313 (O_4313,N_47764,N_47012);
xnor UO_4314 (O_4314,N_48134,N_46442);
and UO_4315 (O_4315,N_46615,N_49059);
and UO_4316 (O_4316,N_49629,N_47294);
xnor UO_4317 (O_4317,N_45468,N_46785);
nor UO_4318 (O_4318,N_49093,N_49773);
xor UO_4319 (O_4319,N_46914,N_46043);
and UO_4320 (O_4320,N_46229,N_48496);
nor UO_4321 (O_4321,N_45670,N_49525);
or UO_4322 (O_4322,N_48721,N_48672);
xor UO_4323 (O_4323,N_47134,N_46141);
or UO_4324 (O_4324,N_47069,N_45059);
nor UO_4325 (O_4325,N_49158,N_49899);
nor UO_4326 (O_4326,N_46736,N_47987);
and UO_4327 (O_4327,N_46635,N_47019);
xor UO_4328 (O_4328,N_49130,N_49160);
or UO_4329 (O_4329,N_45305,N_47460);
nor UO_4330 (O_4330,N_49853,N_45576);
nand UO_4331 (O_4331,N_49670,N_46078);
nor UO_4332 (O_4332,N_48975,N_45866);
nor UO_4333 (O_4333,N_46429,N_45961);
and UO_4334 (O_4334,N_45849,N_47618);
nand UO_4335 (O_4335,N_49105,N_46146);
xnor UO_4336 (O_4336,N_45058,N_46561);
xnor UO_4337 (O_4337,N_47184,N_48090);
nand UO_4338 (O_4338,N_47221,N_49510);
nand UO_4339 (O_4339,N_48454,N_47826);
or UO_4340 (O_4340,N_49359,N_48775);
xnor UO_4341 (O_4341,N_46839,N_46716);
nor UO_4342 (O_4342,N_49411,N_47298);
nor UO_4343 (O_4343,N_48538,N_47056);
and UO_4344 (O_4344,N_47799,N_47627);
nand UO_4345 (O_4345,N_45754,N_45272);
nand UO_4346 (O_4346,N_48329,N_45293);
nor UO_4347 (O_4347,N_47729,N_46950);
xor UO_4348 (O_4348,N_45002,N_48049);
or UO_4349 (O_4349,N_46381,N_48589);
xor UO_4350 (O_4350,N_46702,N_45464);
nand UO_4351 (O_4351,N_49458,N_46477);
xnor UO_4352 (O_4352,N_49007,N_47524);
nand UO_4353 (O_4353,N_47584,N_47232);
and UO_4354 (O_4354,N_49200,N_48255);
nand UO_4355 (O_4355,N_48769,N_49939);
and UO_4356 (O_4356,N_48626,N_48426);
nand UO_4357 (O_4357,N_49299,N_47302);
or UO_4358 (O_4358,N_46683,N_48722);
or UO_4359 (O_4359,N_49143,N_45772);
xnor UO_4360 (O_4360,N_48917,N_49028);
nand UO_4361 (O_4361,N_46156,N_47340);
or UO_4362 (O_4362,N_49074,N_45399);
nor UO_4363 (O_4363,N_47554,N_47282);
and UO_4364 (O_4364,N_45139,N_47804);
nand UO_4365 (O_4365,N_49050,N_46488);
and UO_4366 (O_4366,N_48588,N_49072);
nand UO_4367 (O_4367,N_46148,N_46244);
or UO_4368 (O_4368,N_46498,N_46959);
nor UO_4369 (O_4369,N_49307,N_45175);
nor UO_4370 (O_4370,N_45093,N_46170);
or UO_4371 (O_4371,N_48506,N_48223);
nand UO_4372 (O_4372,N_45779,N_47034);
or UO_4373 (O_4373,N_45643,N_48214);
or UO_4374 (O_4374,N_49685,N_47432);
or UO_4375 (O_4375,N_47723,N_46301);
nor UO_4376 (O_4376,N_46803,N_47058);
nand UO_4377 (O_4377,N_45676,N_49678);
xnor UO_4378 (O_4378,N_46175,N_48630);
and UO_4379 (O_4379,N_49949,N_46731);
nor UO_4380 (O_4380,N_45356,N_47207);
xor UO_4381 (O_4381,N_49815,N_45222);
or UO_4382 (O_4382,N_48145,N_49723);
and UO_4383 (O_4383,N_46879,N_49094);
xor UO_4384 (O_4384,N_45993,N_45201);
and UO_4385 (O_4385,N_45589,N_47782);
xnor UO_4386 (O_4386,N_49178,N_49633);
and UO_4387 (O_4387,N_48257,N_49453);
xor UO_4388 (O_4388,N_48682,N_45023);
nand UO_4389 (O_4389,N_47570,N_48239);
and UO_4390 (O_4390,N_48231,N_49319);
nand UO_4391 (O_4391,N_47335,N_47552);
nor UO_4392 (O_4392,N_49463,N_49104);
and UO_4393 (O_4393,N_46401,N_48928);
xor UO_4394 (O_4394,N_48452,N_45137);
xnor UO_4395 (O_4395,N_49566,N_46672);
or UO_4396 (O_4396,N_49487,N_49028);
nor UO_4397 (O_4397,N_47260,N_45447);
and UO_4398 (O_4398,N_47752,N_49117);
or UO_4399 (O_4399,N_49440,N_45728);
nand UO_4400 (O_4400,N_45713,N_46252);
xor UO_4401 (O_4401,N_47065,N_47414);
nand UO_4402 (O_4402,N_46535,N_47345);
or UO_4403 (O_4403,N_48622,N_48561);
xnor UO_4404 (O_4404,N_45764,N_47684);
nor UO_4405 (O_4405,N_49123,N_45658);
and UO_4406 (O_4406,N_45227,N_48389);
or UO_4407 (O_4407,N_48711,N_46495);
and UO_4408 (O_4408,N_48582,N_46606);
and UO_4409 (O_4409,N_49868,N_48053);
xnor UO_4410 (O_4410,N_47740,N_48487);
or UO_4411 (O_4411,N_47663,N_46553);
nor UO_4412 (O_4412,N_46617,N_49112);
xnor UO_4413 (O_4413,N_49465,N_45804);
nand UO_4414 (O_4414,N_45291,N_47793);
and UO_4415 (O_4415,N_45833,N_49831);
and UO_4416 (O_4416,N_49240,N_46353);
and UO_4417 (O_4417,N_48806,N_47365);
xnor UO_4418 (O_4418,N_47095,N_48077);
nor UO_4419 (O_4419,N_46553,N_48086);
or UO_4420 (O_4420,N_48503,N_49222);
nor UO_4421 (O_4421,N_49303,N_45668);
xnor UO_4422 (O_4422,N_49408,N_48053);
and UO_4423 (O_4423,N_46728,N_46598);
xor UO_4424 (O_4424,N_48476,N_45638);
nor UO_4425 (O_4425,N_47639,N_48390);
nor UO_4426 (O_4426,N_49898,N_48178);
and UO_4427 (O_4427,N_49852,N_48557);
nand UO_4428 (O_4428,N_46702,N_46537);
nor UO_4429 (O_4429,N_45912,N_48872);
or UO_4430 (O_4430,N_45500,N_46102);
nand UO_4431 (O_4431,N_49179,N_46694);
or UO_4432 (O_4432,N_45313,N_47855);
or UO_4433 (O_4433,N_48406,N_47402);
or UO_4434 (O_4434,N_46819,N_47129);
xor UO_4435 (O_4435,N_48661,N_49522);
or UO_4436 (O_4436,N_49476,N_48177);
xnor UO_4437 (O_4437,N_48243,N_47827);
and UO_4438 (O_4438,N_49096,N_47686);
nand UO_4439 (O_4439,N_48266,N_46187);
and UO_4440 (O_4440,N_47692,N_48165);
nand UO_4441 (O_4441,N_45381,N_49948);
and UO_4442 (O_4442,N_47077,N_48810);
xor UO_4443 (O_4443,N_47649,N_49392);
or UO_4444 (O_4444,N_45378,N_49248);
xnor UO_4445 (O_4445,N_49463,N_45145);
nor UO_4446 (O_4446,N_47165,N_47071);
nand UO_4447 (O_4447,N_48249,N_46805);
nor UO_4448 (O_4448,N_46366,N_49423);
nor UO_4449 (O_4449,N_48111,N_45988);
nor UO_4450 (O_4450,N_45104,N_45446);
and UO_4451 (O_4451,N_47171,N_45245);
nand UO_4452 (O_4452,N_48991,N_47485);
or UO_4453 (O_4453,N_49932,N_48287);
or UO_4454 (O_4454,N_45111,N_49925);
nor UO_4455 (O_4455,N_48158,N_48215);
nor UO_4456 (O_4456,N_47266,N_45098);
nor UO_4457 (O_4457,N_48609,N_47101);
and UO_4458 (O_4458,N_48675,N_49557);
xnor UO_4459 (O_4459,N_49049,N_48401);
xor UO_4460 (O_4460,N_48898,N_45037);
and UO_4461 (O_4461,N_48973,N_45749);
xnor UO_4462 (O_4462,N_46113,N_48192);
xor UO_4463 (O_4463,N_48773,N_48149);
xnor UO_4464 (O_4464,N_49406,N_49526);
nor UO_4465 (O_4465,N_47616,N_47592);
nor UO_4466 (O_4466,N_48898,N_49730);
nor UO_4467 (O_4467,N_49659,N_45629);
nand UO_4468 (O_4468,N_45335,N_49649);
xnor UO_4469 (O_4469,N_45917,N_48921);
and UO_4470 (O_4470,N_49171,N_45150);
and UO_4471 (O_4471,N_49453,N_45353);
xnor UO_4472 (O_4472,N_49517,N_48381);
or UO_4473 (O_4473,N_46374,N_47665);
or UO_4474 (O_4474,N_48615,N_46208);
xnor UO_4475 (O_4475,N_49686,N_45316);
xor UO_4476 (O_4476,N_49209,N_48150);
xnor UO_4477 (O_4477,N_48648,N_45711);
and UO_4478 (O_4478,N_46571,N_45907);
nand UO_4479 (O_4479,N_49038,N_46585);
xnor UO_4480 (O_4480,N_47999,N_47708);
nand UO_4481 (O_4481,N_48927,N_47428);
xnor UO_4482 (O_4482,N_46496,N_47007);
or UO_4483 (O_4483,N_45571,N_46066);
xor UO_4484 (O_4484,N_45661,N_47098);
or UO_4485 (O_4485,N_47423,N_45164);
xor UO_4486 (O_4486,N_48697,N_47345);
and UO_4487 (O_4487,N_47262,N_45079);
and UO_4488 (O_4488,N_48054,N_45652);
xnor UO_4489 (O_4489,N_46150,N_47926);
or UO_4490 (O_4490,N_46683,N_45614);
nor UO_4491 (O_4491,N_47468,N_47628);
nand UO_4492 (O_4492,N_47883,N_46009);
nand UO_4493 (O_4493,N_48026,N_49626);
and UO_4494 (O_4494,N_45126,N_48580);
and UO_4495 (O_4495,N_47561,N_48462);
and UO_4496 (O_4496,N_49349,N_46490);
nor UO_4497 (O_4497,N_49176,N_49463);
nand UO_4498 (O_4498,N_45919,N_45643);
nand UO_4499 (O_4499,N_48274,N_47692);
and UO_4500 (O_4500,N_49392,N_46187);
nor UO_4501 (O_4501,N_46102,N_47830);
or UO_4502 (O_4502,N_47319,N_47581);
nand UO_4503 (O_4503,N_45946,N_46600);
and UO_4504 (O_4504,N_48803,N_48562);
xor UO_4505 (O_4505,N_49210,N_45961);
xor UO_4506 (O_4506,N_46926,N_49276);
xor UO_4507 (O_4507,N_47598,N_49497);
nor UO_4508 (O_4508,N_49689,N_48532);
or UO_4509 (O_4509,N_48672,N_46119);
xnor UO_4510 (O_4510,N_45054,N_45089);
nor UO_4511 (O_4511,N_46510,N_47678);
nand UO_4512 (O_4512,N_46451,N_46592);
and UO_4513 (O_4513,N_49417,N_48160);
or UO_4514 (O_4514,N_45026,N_49855);
nor UO_4515 (O_4515,N_46608,N_45292);
xor UO_4516 (O_4516,N_48743,N_47646);
nand UO_4517 (O_4517,N_46695,N_49317);
nor UO_4518 (O_4518,N_48432,N_49609);
and UO_4519 (O_4519,N_48911,N_47118);
or UO_4520 (O_4520,N_49798,N_48886);
xnor UO_4521 (O_4521,N_46848,N_46888);
and UO_4522 (O_4522,N_46638,N_49743);
or UO_4523 (O_4523,N_45727,N_45295);
or UO_4524 (O_4524,N_48353,N_47446);
nor UO_4525 (O_4525,N_47228,N_47248);
xor UO_4526 (O_4526,N_47357,N_48534);
xnor UO_4527 (O_4527,N_46812,N_47040);
and UO_4528 (O_4528,N_48085,N_48437);
nor UO_4529 (O_4529,N_47319,N_49149);
xor UO_4530 (O_4530,N_49794,N_45315);
xor UO_4531 (O_4531,N_45467,N_49825);
nand UO_4532 (O_4532,N_49367,N_45543);
or UO_4533 (O_4533,N_46482,N_46410);
or UO_4534 (O_4534,N_46190,N_47309);
xnor UO_4535 (O_4535,N_48162,N_45680);
nor UO_4536 (O_4536,N_49486,N_46554);
nand UO_4537 (O_4537,N_47253,N_46683);
or UO_4538 (O_4538,N_45872,N_47575);
nand UO_4539 (O_4539,N_46835,N_45769);
or UO_4540 (O_4540,N_46465,N_49317);
xnor UO_4541 (O_4541,N_47065,N_49216);
xnor UO_4542 (O_4542,N_49988,N_47774);
nor UO_4543 (O_4543,N_46864,N_48947);
and UO_4544 (O_4544,N_45472,N_46497);
nor UO_4545 (O_4545,N_45768,N_46500);
nor UO_4546 (O_4546,N_49410,N_45629);
or UO_4547 (O_4547,N_46943,N_47432);
nor UO_4548 (O_4548,N_46358,N_47767);
xor UO_4549 (O_4549,N_45071,N_45086);
xnor UO_4550 (O_4550,N_48905,N_46603);
or UO_4551 (O_4551,N_46389,N_46737);
xor UO_4552 (O_4552,N_47992,N_48943);
or UO_4553 (O_4553,N_45522,N_47854);
nor UO_4554 (O_4554,N_46582,N_45788);
and UO_4555 (O_4555,N_47972,N_48471);
nand UO_4556 (O_4556,N_46594,N_48596);
xnor UO_4557 (O_4557,N_49710,N_46710);
or UO_4558 (O_4558,N_46835,N_48019);
or UO_4559 (O_4559,N_45775,N_49674);
or UO_4560 (O_4560,N_46776,N_46786);
nand UO_4561 (O_4561,N_46124,N_48051);
and UO_4562 (O_4562,N_47606,N_45519);
and UO_4563 (O_4563,N_49061,N_47161);
nand UO_4564 (O_4564,N_45478,N_47872);
nor UO_4565 (O_4565,N_46348,N_48521);
xor UO_4566 (O_4566,N_46010,N_47855);
and UO_4567 (O_4567,N_47312,N_47962);
or UO_4568 (O_4568,N_49034,N_47810);
nand UO_4569 (O_4569,N_47751,N_48268);
nand UO_4570 (O_4570,N_46915,N_48872);
and UO_4571 (O_4571,N_48608,N_48893);
xnor UO_4572 (O_4572,N_48373,N_45172);
and UO_4573 (O_4573,N_47998,N_46708);
and UO_4574 (O_4574,N_47952,N_49929);
nand UO_4575 (O_4575,N_46753,N_49438);
nor UO_4576 (O_4576,N_49192,N_49111);
or UO_4577 (O_4577,N_48953,N_48883);
nand UO_4578 (O_4578,N_47281,N_45296);
nand UO_4579 (O_4579,N_48001,N_47238);
or UO_4580 (O_4580,N_47031,N_46492);
nand UO_4581 (O_4581,N_47844,N_47687);
nand UO_4582 (O_4582,N_45355,N_45281);
or UO_4583 (O_4583,N_45951,N_46300);
nor UO_4584 (O_4584,N_49212,N_45956);
or UO_4585 (O_4585,N_49820,N_45674);
xnor UO_4586 (O_4586,N_45040,N_45942);
and UO_4587 (O_4587,N_47817,N_46410);
xor UO_4588 (O_4588,N_47148,N_45123);
xnor UO_4589 (O_4589,N_49378,N_45612);
xor UO_4590 (O_4590,N_48825,N_46594);
xnor UO_4591 (O_4591,N_46598,N_46426);
xor UO_4592 (O_4592,N_46910,N_45123);
nor UO_4593 (O_4593,N_48617,N_48585);
and UO_4594 (O_4594,N_49687,N_48060);
nand UO_4595 (O_4595,N_49995,N_48100);
xor UO_4596 (O_4596,N_45481,N_46580);
nor UO_4597 (O_4597,N_47607,N_48274);
nor UO_4598 (O_4598,N_46394,N_45427);
nor UO_4599 (O_4599,N_45145,N_47716);
and UO_4600 (O_4600,N_49483,N_48354);
nor UO_4601 (O_4601,N_47563,N_48863);
nor UO_4602 (O_4602,N_46954,N_47357);
nor UO_4603 (O_4603,N_49522,N_46451);
nand UO_4604 (O_4604,N_45349,N_49310);
and UO_4605 (O_4605,N_46146,N_45768);
nor UO_4606 (O_4606,N_49145,N_46347);
or UO_4607 (O_4607,N_47998,N_45502);
nor UO_4608 (O_4608,N_47841,N_48810);
nand UO_4609 (O_4609,N_45685,N_45648);
and UO_4610 (O_4610,N_47165,N_46702);
nand UO_4611 (O_4611,N_46273,N_48860);
nor UO_4612 (O_4612,N_47472,N_48792);
or UO_4613 (O_4613,N_47021,N_48570);
and UO_4614 (O_4614,N_46455,N_47527);
nor UO_4615 (O_4615,N_46997,N_48122);
nand UO_4616 (O_4616,N_49962,N_47737);
or UO_4617 (O_4617,N_49202,N_49389);
and UO_4618 (O_4618,N_48990,N_49696);
xnor UO_4619 (O_4619,N_47583,N_49555);
nor UO_4620 (O_4620,N_49619,N_49009);
nand UO_4621 (O_4621,N_48801,N_46433);
nor UO_4622 (O_4622,N_45891,N_49069);
and UO_4623 (O_4623,N_49194,N_46690);
and UO_4624 (O_4624,N_48604,N_48486);
or UO_4625 (O_4625,N_47489,N_47264);
nor UO_4626 (O_4626,N_48407,N_45312);
nor UO_4627 (O_4627,N_47894,N_45943);
xnor UO_4628 (O_4628,N_47773,N_45325);
xor UO_4629 (O_4629,N_48147,N_48928);
nor UO_4630 (O_4630,N_46450,N_45202);
nand UO_4631 (O_4631,N_49562,N_47567);
xor UO_4632 (O_4632,N_47649,N_49062);
or UO_4633 (O_4633,N_46593,N_48095);
and UO_4634 (O_4634,N_46894,N_48070);
and UO_4635 (O_4635,N_46811,N_45446);
nand UO_4636 (O_4636,N_47000,N_45853);
xnor UO_4637 (O_4637,N_45312,N_45645);
and UO_4638 (O_4638,N_47136,N_47439);
nand UO_4639 (O_4639,N_49674,N_47091);
nand UO_4640 (O_4640,N_49907,N_45365);
nand UO_4641 (O_4641,N_47718,N_47464);
or UO_4642 (O_4642,N_47066,N_47555);
and UO_4643 (O_4643,N_48823,N_47779);
and UO_4644 (O_4644,N_45232,N_48295);
or UO_4645 (O_4645,N_46738,N_48934);
nand UO_4646 (O_4646,N_48758,N_48825);
or UO_4647 (O_4647,N_49341,N_47184);
nor UO_4648 (O_4648,N_46974,N_45465);
nor UO_4649 (O_4649,N_45815,N_45009);
nand UO_4650 (O_4650,N_47525,N_49904);
and UO_4651 (O_4651,N_48712,N_49435);
xor UO_4652 (O_4652,N_47897,N_49988);
xnor UO_4653 (O_4653,N_47522,N_48746);
and UO_4654 (O_4654,N_48336,N_48525);
and UO_4655 (O_4655,N_47405,N_45045);
and UO_4656 (O_4656,N_46863,N_45822);
or UO_4657 (O_4657,N_48891,N_46450);
xor UO_4658 (O_4658,N_49715,N_48138);
nand UO_4659 (O_4659,N_48618,N_48708);
and UO_4660 (O_4660,N_45388,N_45152);
xor UO_4661 (O_4661,N_45422,N_49593);
or UO_4662 (O_4662,N_45534,N_49336);
nor UO_4663 (O_4663,N_48018,N_47191);
or UO_4664 (O_4664,N_45815,N_45625);
nand UO_4665 (O_4665,N_47616,N_45783);
and UO_4666 (O_4666,N_49114,N_49835);
and UO_4667 (O_4667,N_48530,N_49799);
or UO_4668 (O_4668,N_45693,N_46686);
or UO_4669 (O_4669,N_48765,N_46608);
nor UO_4670 (O_4670,N_47532,N_49221);
xor UO_4671 (O_4671,N_47059,N_46361);
and UO_4672 (O_4672,N_48238,N_45942);
or UO_4673 (O_4673,N_49157,N_46909);
or UO_4674 (O_4674,N_48779,N_47511);
and UO_4675 (O_4675,N_49749,N_48358);
or UO_4676 (O_4676,N_48897,N_45149);
or UO_4677 (O_4677,N_48531,N_46662);
and UO_4678 (O_4678,N_46478,N_45651);
xor UO_4679 (O_4679,N_46769,N_45203);
or UO_4680 (O_4680,N_46875,N_47670);
or UO_4681 (O_4681,N_47050,N_47430);
nand UO_4682 (O_4682,N_47125,N_45092);
nor UO_4683 (O_4683,N_48355,N_46796);
and UO_4684 (O_4684,N_49553,N_46389);
nand UO_4685 (O_4685,N_46652,N_48613);
and UO_4686 (O_4686,N_46591,N_46135);
nor UO_4687 (O_4687,N_47860,N_48290);
nand UO_4688 (O_4688,N_46421,N_48164);
xor UO_4689 (O_4689,N_48057,N_48943);
xnor UO_4690 (O_4690,N_45595,N_46374);
and UO_4691 (O_4691,N_47720,N_48903);
and UO_4692 (O_4692,N_47256,N_46562);
or UO_4693 (O_4693,N_47923,N_47174);
nand UO_4694 (O_4694,N_48365,N_49241);
and UO_4695 (O_4695,N_47797,N_49000);
and UO_4696 (O_4696,N_47110,N_47740);
nor UO_4697 (O_4697,N_46235,N_48739);
nand UO_4698 (O_4698,N_49567,N_46999);
nand UO_4699 (O_4699,N_46984,N_49472);
nand UO_4700 (O_4700,N_46261,N_48173);
nand UO_4701 (O_4701,N_45227,N_45321);
xnor UO_4702 (O_4702,N_46253,N_49777);
nor UO_4703 (O_4703,N_47067,N_45232);
xor UO_4704 (O_4704,N_48571,N_45109);
nor UO_4705 (O_4705,N_45050,N_45386);
nand UO_4706 (O_4706,N_49646,N_49386);
nor UO_4707 (O_4707,N_48732,N_49328);
and UO_4708 (O_4708,N_49335,N_47167);
nand UO_4709 (O_4709,N_46404,N_45250);
nand UO_4710 (O_4710,N_46076,N_48237);
or UO_4711 (O_4711,N_47957,N_47166);
nor UO_4712 (O_4712,N_47975,N_49044);
nor UO_4713 (O_4713,N_46340,N_48867);
or UO_4714 (O_4714,N_49788,N_46408);
or UO_4715 (O_4715,N_48636,N_47294);
nand UO_4716 (O_4716,N_49785,N_45568);
nand UO_4717 (O_4717,N_48415,N_49744);
nor UO_4718 (O_4718,N_49411,N_47360);
xor UO_4719 (O_4719,N_48348,N_47609);
nor UO_4720 (O_4720,N_47231,N_46912);
and UO_4721 (O_4721,N_47324,N_46634);
xnor UO_4722 (O_4722,N_46845,N_49818);
and UO_4723 (O_4723,N_46230,N_49675);
xnor UO_4724 (O_4724,N_46732,N_49846);
nand UO_4725 (O_4725,N_45726,N_48622);
and UO_4726 (O_4726,N_46785,N_48485);
nand UO_4727 (O_4727,N_47432,N_45680);
or UO_4728 (O_4728,N_48533,N_48369);
nor UO_4729 (O_4729,N_46875,N_45578);
and UO_4730 (O_4730,N_48280,N_46565);
xor UO_4731 (O_4731,N_45579,N_45047);
nand UO_4732 (O_4732,N_46617,N_45827);
nand UO_4733 (O_4733,N_46591,N_46203);
xnor UO_4734 (O_4734,N_45913,N_45829);
or UO_4735 (O_4735,N_49079,N_46995);
nand UO_4736 (O_4736,N_46808,N_48698);
xnor UO_4737 (O_4737,N_48448,N_45305);
nand UO_4738 (O_4738,N_46935,N_46126);
or UO_4739 (O_4739,N_45002,N_46839);
nand UO_4740 (O_4740,N_46161,N_49876);
or UO_4741 (O_4741,N_45718,N_48576);
and UO_4742 (O_4742,N_45995,N_48957);
or UO_4743 (O_4743,N_47969,N_48020);
nor UO_4744 (O_4744,N_47679,N_46043);
and UO_4745 (O_4745,N_45160,N_46862);
or UO_4746 (O_4746,N_46448,N_48000);
nand UO_4747 (O_4747,N_47754,N_48521);
nand UO_4748 (O_4748,N_49096,N_47220);
or UO_4749 (O_4749,N_49599,N_45635);
or UO_4750 (O_4750,N_47221,N_46927);
nand UO_4751 (O_4751,N_47657,N_46991);
xnor UO_4752 (O_4752,N_49149,N_47169);
or UO_4753 (O_4753,N_48652,N_45827);
nor UO_4754 (O_4754,N_46779,N_45178);
nor UO_4755 (O_4755,N_49497,N_47647);
or UO_4756 (O_4756,N_45150,N_48753);
nor UO_4757 (O_4757,N_45249,N_46904);
nand UO_4758 (O_4758,N_48405,N_46501);
nand UO_4759 (O_4759,N_46836,N_47332);
xnor UO_4760 (O_4760,N_47147,N_47134);
nor UO_4761 (O_4761,N_47286,N_45980);
nor UO_4762 (O_4762,N_49509,N_47876);
or UO_4763 (O_4763,N_47306,N_48720);
nor UO_4764 (O_4764,N_45599,N_46999);
nand UO_4765 (O_4765,N_47980,N_46837);
nor UO_4766 (O_4766,N_48031,N_49036);
or UO_4767 (O_4767,N_45741,N_45821);
or UO_4768 (O_4768,N_48484,N_48311);
nor UO_4769 (O_4769,N_45821,N_47084);
xnor UO_4770 (O_4770,N_49330,N_47426);
nor UO_4771 (O_4771,N_49682,N_46964);
or UO_4772 (O_4772,N_45280,N_46959);
nand UO_4773 (O_4773,N_46239,N_47486);
xor UO_4774 (O_4774,N_49690,N_45755);
nand UO_4775 (O_4775,N_46496,N_47816);
nor UO_4776 (O_4776,N_49415,N_49000);
or UO_4777 (O_4777,N_45904,N_47567);
and UO_4778 (O_4778,N_48054,N_49974);
nand UO_4779 (O_4779,N_49573,N_48322);
xor UO_4780 (O_4780,N_48422,N_49207);
nand UO_4781 (O_4781,N_45654,N_45936);
or UO_4782 (O_4782,N_46201,N_47697);
or UO_4783 (O_4783,N_49451,N_46015);
nand UO_4784 (O_4784,N_48935,N_45531);
xor UO_4785 (O_4785,N_47153,N_47594);
nor UO_4786 (O_4786,N_47247,N_48605);
nand UO_4787 (O_4787,N_47494,N_48050);
xor UO_4788 (O_4788,N_45371,N_45599);
nand UO_4789 (O_4789,N_49147,N_49289);
nand UO_4790 (O_4790,N_47441,N_45905);
xnor UO_4791 (O_4791,N_46163,N_49263);
nand UO_4792 (O_4792,N_47208,N_47519);
xnor UO_4793 (O_4793,N_46303,N_45490);
nand UO_4794 (O_4794,N_49828,N_47019);
or UO_4795 (O_4795,N_47063,N_48741);
and UO_4796 (O_4796,N_47711,N_46044);
xnor UO_4797 (O_4797,N_49795,N_46552);
and UO_4798 (O_4798,N_46789,N_49081);
and UO_4799 (O_4799,N_47013,N_47326);
nand UO_4800 (O_4800,N_45435,N_45616);
xor UO_4801 (O_4801,N_47290,N_46177);
nor UO_4802 (O_4802,N_47367,N_46541);
nand UO_4803 (O_4803,N_46283,N_46220);
and UO_4804 (O_4804,N_45766,N_48919);
nand UO_4805 (O_4805,N_49109,N_46232);
and UO_4806 (O_4806,N_49396,N_48176);
or UO_4807 (O_4807,N_48935,N_48001);
and UO_4808 (O_4808,N_48997,N_48234);
or UO_4809 (O_4809,N_49423,N_48537);
or UO_4810 (O_4810,N_49522,N_45251);
and UO_4811 (O_4811,N_45554,N_49676);
and UO_4812 (O_4812,N_47652,N_47044);
nor UO_4813 (O_4813,N_46689,N_46213);
and UO_4814 (O_4814,N_45015,N_48104);
xnor UO_4815 (O_4815,N_49457,N_47798);
and UO_4816 (O_4816,N_47849,N_47918);
nand UO_4817 (O_4817,N_45096,N_48740);
xor UO_4818 (O_4818,N_45353,N_46691);
xor UO_4819 (O_4819,N_46167,N_45706);
or UO_4820 (O_4820,N_47830,N_48251);
and UO_4821 (O_4821,N_45178,N_46201);
or UO_4822 (O_4822,N_49404,N_47330);
and UO_4823 (O_4823,N_48237,N_45161);
nor UO_4824 (O_4824,N_45194,N_46186);
xnor UO_4825 (O_4825,N_46437,N_46595);
or UO_4826 (O_4826,N_47597,N_45765);
nor UO_4827 (O_4827,N_49854,N_47771);
xor UO_4828 (O_4828,N_47445,N_49747);
and UO_4829 (O_4829,N_49325,N_46184);
nor UO_4830 (O_4830,N_45303,N_49095);
xor UO_4831 (O_4831,N_46657,N_47332);
xnor UO_4832 (O_4832,N_46684,N_47320);
nand UO_4833 (O_4833,N_46855,N_48204);
xnor UO_4834 (O_4834,N_47475,N_45968);
and UO_4835 (O_4835,N_45264,N_48299);
or UO_4836 (O_4836,N_47011,N_48518);
and UO_4837 (O_4837,N_47901,N_48163);
or UO_4838 (O_4838,N_47233,N_45186);
or UO_4839 (O_4839,N_47138,N_47568);
nor UO_4840 (O_4840,N_47450,N_46894);
nor UO_4841 (O_4841,N_48672,N_45495);
xnor UO_4842 (O_4842,N_48433,N_48201);
and UO_4843 (O_4843,N_46916,N_45323);
xor UO_4844 (O_4844,N_45257,N_48100);
nor UO_4845 (O_4845,N_45314,N_49244);
xor UO_4846 (O_4846,N_48173,N_49579);
nand UO_4847 (O_4847,N_49128,N_49889);
xor UO_4848 (O_4848,N_49822,N_47712);
or UO_4849 (O_4849,N_48312,N_49922);
and UO_4850 (O_4850,N_48366,N_49425);
xor UO_4851 (O_4851,N_45027,N_46312);
nand UO_4852 (O_4852,N_49004,N_47349);
nor UO_4853 (O_4853,N_48782,N_45709);
nand UO_4854 (O_4854,N_46093,N_48896);
xor UO_4855 (O_4855,N_46187,N_45436);
nor UO_4856 (O_4856,N_49242,N_49574);
nand UO_4857 (O_4857,N_46591,N_46849);
nor UO_4858 (O_4858,N_49719,N_48331);
or UO_4859 (O_4859,N_46022,N_47386);
nand UO_4860 (O_4860,N_49245,N_47437);
nand UO_4861 (O_4861,N_46532,N_49619);
xnor UO_4862 (O_4862,N_45442,N_45638);
nand UO_4863 (O_4863,N_49936,N_46862);
nand UO_4864 (O_4864,N_46684,N_46506);
or UO_4865 (O_4865,N_46123,N_49650);
or UO_4866 (O_4866,N_48444,N_47669);
nor UO_4867 (O_4867,N_47400,N_46068);
xnor UO_4868 (O_4868,N_49535,N_48372);
and UO_4869 (O_4869,N_45105,N_45578);
nand UO_4870 (O_4870,N_48926,N_49805);
and UO_4871 (O_4871,N_45956,N_45418);
nand UO_4872 (O_4872,N_45572,N_49503);
or UO_4873 (O_4873,N_46169,N_48679);
xnor UO_4874 (O_4874,N_46383,N_48510);
nor UO_4875 (O_4875,N_45532,N_46007);
or UO_4876 (O_4876,N_48142,N_48320);
or UO_4877 (O_4877,N_48375,N_47097);
xnor UO_4878 (O_4878,N_47237,N_47129);
xor UO_4879 (O_4879,N_46967,N_47469);
or UO_4880 (O_4880,N_45419,N_47403);
nand UO_4881 (O_4881,N_48202,N_49902);
xnor UO_4882 (O_4882,N_49458,N_47826);
or UO_4883 (O_4883,N_45517,N_46785);
and UO_4884 (O_4884,N_48002,N_48998);
xnor UO_4885 (O_4885,N_45798,N_49582);
and UO_4886 (O_4886,N_45049,N_46134);
nor UO_4887 (O_4887,N_46059,N_49062);
xor UO_4888 (O_4888,N_45109,N_47122);
or UO_4889 (O_4889,N_47710,N_45787);
nand UO_4890 (O_4890,N_46494,N_49966);
or UO_4891 (O_4891,N_45400,N_47517);
or UO_4892 (O_4892,N_45260,N_46792);
or UO_4893 (O_4893,N_45972,N_48816);
or UO_4894 (O_4894,N_47522,N_46006);
and UO_4895 (O_4895,N_46602,N_48621);
nor UO_4896 (O_4896,N_48636,N_46104);
nand UO_4897 (O_4897,N_45799,N_45960);
xor UO_4898 (O_4898,N_48231,N_47854);
or UO_4899 (O_4899,N_49477,N_47221);
or UO_4900 (O_4900,N_48986,N_47924);
or UO_4901 (O_4901,N_48806,N_45718);
nor UO_4902 (O_4902,N_45919,N_47264);
and UO_4903 (O_4903,N_48566,N_46513);
or UO_4904 (O_4904,N_47239,N_46073);
nor UO_4905 (O_4905,N_46083,N_49540);
nand UO_4906 (O_4906,N_47891,N_46475);
and UO_4907 (O_4907,N_46540,N_48790);
and UO_4908 (O_4908,N_49756,N_49111);
or UO_4909 (O_4909,N_46493,N_49389);
nand UO_4910 (O_4910,N_47664,N_48383);
nor UO_4911 (O_4911,N_46201,N_45065);
nor UO_4912 (O_4912,N_49996,N_46344);
and UO_4913 (O_4913,N_47570,N_45710);
nand UO_4914 (O_4914,N_49459,N_49401);
or UO_4915 (O_4915,N_46883,N_45541);
nor UO_4916 (O_4916,N_45470,N_47675);
nand UO_4917 (O_4917,N_48975,N_46944);
nand UO_4918 (O_4918,N_48984,N_45492);
nand UO_4919 (O_4919,N_46880,N_49368);
xnor UO_4920 (O_4920,N_46482,N_47520);
xor UO_4921 (O_4921,N_47197,N_47842);
or UO_4922 (O_4922,N_46512,N_47316);
nand UO_4923 (O_4923,N_48575,N_47452);
nor UO_4924 (O_4924,N_46028,N_48060);
and UO_4925 (O_4925,N_45623,N_48096);
nand UO_4926 (O_4926,N_49138,N_46875);
nor UO_4927 (O_4927,N_47823,N_45534);
nor UO_4928 (O_4928,N_49763,N_47581);
or UO_4929 (O_4929,N_47632,N_49112);
nand UO_4930 (O_4930,N_45244,N_49690);
xor UO_4931 (O_4931,N_49429,N_49371);
and UO_4932 (O_4932,N_48881,N_47791);
xnor UO_4933 (O_4933,N_48399,N_47538);
or UO_4934 (O_4934,N_45719,N_47315);
nor UO_4935 (O_4935,N_49100,N_49132);
or UO_4936 (O_4936,N_46223,N_45026);
xnor UO_4937 (O_4937,N_46507,N_46356);
and UO_4938 (O_4938,N_47260,N_46527);
or UO_4939 (O_4939,N_48522,N_49694);
xnor UO_4940 (O_4940,N_45141,N_49372);
or UO_4941 (O_4941,N_49746,N_48256);
and UO_4942 (O_4942,N_47564,N_47270);
and UO_4943 (O_4943,N_47899,N_49373);
nor UO_4944 (O_4944,N_48190,N_46479);
xor UO_4945 (O_4945,N_46193,N_45877);
or UO_4946 (O_4946,N_49627,N_48107);
or UO_4947 (O_4947,N_47381,N_46258);
xor UO_4948 (O_4948,N_45182,N_49346);
nand UO_4949 (O_4949,N_48105,N_46790);
and UO_4950 (O_4950,N_48613,N_48536);
nor UO_4951 (O_4951,N_49104,N_47033);
and UO_4952 (O_4952,N_47963,N_49348);
xor UO_4953 (O_4953,N_47031,N_46858);
xor UO_4954 (O_4954,N_46575,N_47366);
or UO_4955 (O_4955,N_47981,N_47341);
or UO_4956 (O_4956,N_46586,N_48195);
and UO_4957 (O_4957,N_48320,N_45009);
nand UO_4958 (O_4958,N_47650,N_46959);
or UO_4959 (O_4959,N_47514,N_49315);
and UO_4960 (O_4960,N_46933,N_46488);
nor UO_4961 (O_4961,N_49640,N_45036);
and UO_4962 (O_4962,N_45063,N_45583);
or UO_4963 (O_4963,N_49371,N_48915);
and UO_4964 (O_4964,N_49640,N_49804);
or UO_4965 (O_4965,N_49581,N_46119);
xor UO_4966 (O_4966,N_45059,N_48380);
nand UO_4967 (O_4967,N_47021,N_46295);
nor UO_4968 (O_4968,N_47486,N_47757);
xor UO_4969 (O_4969,N_46642,N_47311);
or UO_4970 (O_4970,N_46198,N_45265);
and UO_4971 (O_4971,N_48401,N_48337);
nor UO_4972 (O_4972,N_47426,N_48512);
or UO_4973 (O_4973,N_49178,N_48630);
nand UO_4974 (O_4974,N_48123,N_48710);
or UO_4975 (O_4975,N_49827,N_47131);
nand UO_4976 (O_4976,N_49225,N_47524);
and UO_4977 (O_4977,N_49338,N_45036);
or UO_4978 (O_4978,N_49721,N_49107);
or UO_4979 (O_4979,N_47968,N_47200);
nand UO_4980 (O_4980,N_45357,N_45274);
nand UO_4981 (O_4981,N_47381,N_48459);
nand UO_4982 (O_4982,N_49595,N_46693);
and UO_4983 (O_4983,N_45043,N_49519);
and UO_4984 (O_4984,N_48517,N_48224);
nand UO_4985 (O_4985,N_47859,N_46935);
nor UO_4986 (O_4986,N_47966,N_46906);
and UO_4987 (O_4987,N_45227,N_45318);
or UO_4988 (O_4988,N_46273,N_45343);
and UO_4989 (O_4989,N_45781,N_47513);
nor UO_4990 (O_4990,N_49974,N_45452);
xor UO_4991 (O_4991,N_47454,N_49157);
and UO_4992 (O_4992,N_49613,N_46158);
or UO_4993 (O_4993,N_49078,N_45632);
xnor UO_4994 (O_4994,N_45033,N_49235);
and UO_4995 (O_4995,N_47405,N_49238);
or UO_4996 (O_4996,N_49452,N_49817);
or UO_4997 (O_4997,N_48201,N_46640);
nor UO_4998 (O_4998,N_45707,N_49949);
nand UO_4999 (O_4999,N_48986,N_48731);
endmodule