module basic_3000_30000_3500_20_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nor U0 (N_0,In_507,In_1251);
and U1 (N_1,In_2123,In_823);
xnor U2 (N_2,In_383,In_1013);
xnor U3 (N_3,In_2589,In_1472);
nand U4 (N_4,In_2328,In_1241);
nand U5 (N_5,In_2876,In_1652);
nand U6 (N_6,In_2420,In_14);
nand U7 (N_7,In_2003,In_1998);
or U8 (N_8,In_2588,In_205);
or U9 (N_9,In_1087,In_2626);
or U10 (N_10,In_1820,In_829);
and U11 (N_11,In_1059,In_1931);
and U12 (N_12,In_1044,In_2628);
nor U13 (N_13,In_2061,In_761);
xor U14 (N_14,In_2435,In_2457);
nand U15 (N_15,In_2811,In_1555);
or U16 (N_16,In_54,In_2257);
xor U17 (N_17,In_892,In_366);
nand U18 (N_18,In_296,In_1848);
or U19 (N_19,In_2385,In_2012);
nand U20 (N_20,In_1023,In_889);
and U21 (N_21,In_574,In_1563);
xnor U22 (N_22,In_938,In_1674);
nor U23 (N_23,In_1182,In_2602);
nand U24 (N_24,In_956,In_2826);
xnor U25 (N_25,In_1782,In_2750);
nor U26 (N_26,In_438,In_1447);
nand U27 (N_27,In_2646,In_1121);
xor U28 (N_28,In_2296,In_532);
xnor U29 (N_29,In_1866,In_2301);
nand U30 (N_30,In_1426,In_1637);
nor U31 (N_31,In_1539,In_2921);
and U32 (N_32,In_598,In_2065);
and U33 (N_33,In_55,In_1729);
nand U34 (N_34,In_2514,In_2007);
nor U35 (N_35,In_817,In_1794);
nand U36 (N_36,In_312,In_2358);
or U37 (N_37,In_2197,In_1409);
or U38 (N_38,In_1366,In_1961);
nor U39 (N_39,In_17,In_2576);
and U40 (N_40,In_1653,In_1672);
and U41 (N_41,In_579,In_1165);
or U42 (N_42,In_1855,In_2615);
and U43 (N_43,In_927,In_2504);
xnor U44 (N_44,In_1684,In_279);
nor U45 (N_45,In_861,In_719);
nor U46 (N_46,In_336,In_2783);
and U47 (N_47,In_1471,In_2163);
or U48 (N_48,In_2975,In_2703);
and U49 (N_49,In_2970,In_1358);
nor U50 (N_50,In_670,In_1433);
xnor U51 (N_51,In_2841,In_710);
nor U52 (N_52,In_2869,In_1244);
xnor U53 (N_53,In_2484,In_890);
or U54 (N_54,In_2530,In_1565);
nor U55 (N_55,In_2668,In_1493);
nor U56 (N_56,In_1047,In_1298);
xor U57 (N_57,In_1516,In_799);
and U58 (N_58,In_601,In_304);
and U59 (N_59,In_1970,In_1140);
nand U60 (N_60,In_391,In_2863);
xor U61 (N_61,In_2854,In_2355);
nand U62 (N_62,In_74,In_2945);
and U63 (N_63,In_2164,In_360);
xnor U64 (N_64,In_993,In_2254);
or U65 (N_65,In_2860,In_169);
nand U66 (N_66,In_1300,In_204);
nor U67 (N_67,In_197,In_129);
or U68 (N_68,In_999,In_363);
xnor U69 (N_69,In_2584,In_1091);
or U70 (N_70,In_315,In_1428);
xor U71 (N_71,In_1473,In_1261);
nand U72 (N_72,In_1751,In_2287);
or U73 (N_73,In_758,In_611);
and U74 (N_74,In_1865,In_2095);
nor U75 (N_75,In_2045,In_1499);
or U76 (N_76,In_2680,In_2511);
xor U77 (N_77,In_236,In_2746);
and U78 (N_78,In_800,In_1845);
nor U79 (N_79,In_2443,In_2232);
nor U80 (N_80,In_530,In_176);
or U81 (N_81,In_886,In_2619);
and U82 (N_82,In_2546,In_2882);
nor U83 (N_83,In_2943,In_529);
xor U84 (N_84,In_2370,In_1029);
or U85 (N_85,In_1545,In_2636);
nand U86 (N_86,In_2987,In_2684);
nand U87 (N_87,In_1993,In_930);
nand U88 (N_88,In_618,In_479);
xor U89 (N_89,In_2742,In_1785);
xor U90 (N_90,In_2275,In_994);
and U91 (N_91,In_2590,In_520);
nand U92 (N_92,In_1916,In_2521);
or U93 (N_93,In_2969,In_1895);
nor U94 (N_94,In_1700,In_584);
or U95 (N_95,In_2110,In_76);
and U96 (N_96,In_753,In_1031);
or U97 (N_97,In_456,In_634);
xnor U98 (N_98,In_688,In_119);
nand U99 (N_99,In_1245,In_1954);
xnor U100 (N_100,In_906,In_2939);
and U101 (N_101,In_2607,In_70);
and U102 (N_102,In_277,In_2167);
or U103 (N_103,In_1329,In_418);
or U104 (N_104,In_1459,In_1491);
xor U105 (N_105,In_2131,In_275);
xor U106 (N_106,In_1033,In_343);
nor U107 (N_107,In_2835,In_1211);
xnor U108 (N_108,In_2729,In_1085);
nor U109 (N_109,In_2027,In_1341);
or U110 (N_110,In_2304,In_1689);
nand U111 (N_111,In_2688,In_1922);
and U112 (N_112,In_439,In_593);
and U113 (N_113,In_2136,In_1372);
xor U114 (N_114,In_1334,In_1317);
nand U115 (N_115,In_1660,In_655);
or U116 (N_116,In_193,In_1202);
nand U117 (N_117,In_1750,In_489);
nor U118 (N_118,In_66,In_1945);
nor U119 (N_119,In_210,In_1753);
and U120 (N_120,In_2676,In_1625);
xor U121 (N_121,In_1926,In_2345);
and U122 (N_122,In_1811,In_146);
nand U123 (N_123,In_2427,In_2525);
nor U124 (N_124,In_2815,In_2694);
or U125 (N_125,In_1237,In_2940);
nor U126 (N_126,In_306,In_745);
nor U127 (N_127,In_377,In_577);
nand U128 (N_128,In_2772,In_943);
nand U129 (N_129,In_928,In_1490);
xnor U130 (N_130,In_287,In_154);
and U131 (N_131,In_258,In_522);
or U132 (N_132,In_1803,In_669);
xnor U133 (N_133,In_293,In_1614);
nand U134 (N_134,In_1139,In_2433);
nor U135 (N_135,In_2338,In_2204);
nor U136 (N_136,In_924,In_2473);
or U137 (N_137,In_1541,In_2474);
and U138 (N_138,In_2812,In_2038);
and U139 (N_139,In_61,In_2735);
and U140 (N_140,In_1159,In_945);
nand U141 (N_141,In_1407,In_2417);
or U142 (N_142,In_1369,In_867);
nor U143 (N_143,In_603,In_1512);
and U144 (N_144,In_2893,In_364);
nor U145 (N_145,In_772,In_1639);
xnor U146 (N_146,In_1870,In_1632);
nand U147 (N_147,In_971,In_255);
and U148 (N_148,In_71,In_2214);
nor U149 (N_149,In_318,In_2468);
or U150 (N_150,In_732,In_1798);
and U151 (N_151,In_1443,In_1232);
nand U152 (N_152,In_1017,In_1101);
nor U153 (N_153,In_1773,In_1109);
xor U154 (N_154,In_2864,In_2599);
xor U155 (N_155,In_1483,In_2377);
or U156 (N_156,In_623,In_724);
nand U157 (N_157,In_513,In_1209);
nand U158 (N_158,In_1401,In_2660);
nand U159 (N_159,In_1935,In_822);
nand U160 (N_160,In_1014,In_2999);
nand U161 (N_161,In_1415,In_1884);
nor U162 (N_162,In_2463,In_1791);
xor U163 (N_163,In_1707,In_1715);
nand U164 (N_164,In_173,In_2302);
and U165 (N_165,In_853,In_1011);
nand U166 (N_166,In_828,In_1021);
xor U167 (N_167,In_1966,In_1733);
and U168 (N_168,In_535,In_609);
and U169 (N_169,In_1305,In_2924);
or U170 (N_170,In_1034,In_639);
and U171 (N_171,In_1705,In_1254);
nor U172 (N_172,In_2568,In_1560);
and U173 (N_173,In_222,In_478);
and U174 (N_174,In_1188,In_733);
nor U175 (N_175,In_1214,In_441);
nand U176 (N_176,In_1243,In_2126);
nor U177 (N_177,In_2830,In_2498);
and U178 (N_178,In_1150,In_1600);
or U179 (N_179,In_1421,In_356);
xnor U180 (N_180,In_1666,In_2212);
or U181 (N_181,In_722,In_1941);
nor U182 (N_182,In_1788,In_773);
xor U183 (N_183,In_379,In_1989);
xor U184 (N_184,In_445,In_2327);
nor U185 (N_185,In_2129,In_1780);
and U186 (N_186,In_384,In_1053);
nand U187 (N_187,In_1404,In_2563);
xor U188 (N_188,In_2082,In_795);
xor U189 (N_189,In_2380,In_2566);
nor U190 (N_190,In_1892,In_2984);
and U191 (N_191,In_806,In_1082);
or U192 (N_192,In_341,In_1332);
nor U193 (N_193,In_2243,In_240);
and U194 (N_194,In_2223,In_1528);
or U195 (N_195,In_407,In_405);
or U196 (N_196,In_983,In_2579);
nand U197 (N_197,In_524,In_159);
nand U198 (N_198,In_2925,In_1740);
xor U199 (N_199,In_947,In_1362);
nor U200 (N_200,In_2393,In_201);
nand U201 (N_201,In_1032,In_40);
or U202 (N_202,In_1772,In_2536);
nand U203 (N_203,In_2887,In_1668);
nand U204 (N_204,In_43,In_1155);
nand U205 (N_205,In_2312,In_86);
or U206 (N_206,In_359,In_741);
or U207 (N_207,In_2667,In_495);
or U208 (N_208,In_189,In_1403);
xor U209 (N_209,In_1842,In_713);
nand U210 (N_210,In_2060,In_1292);
xnor U211 (N_211,In_857,In_1593);
or U212 (N_212,In_1015,In_2187);
and U213 (N_213,In_693,In_314);
and U214 (N_214,In_2567,In_1535);
and U215 (N_215,In_1641,In_1843);
or U216 (N_216,In_746,In_1546);
or U217 (N_217,In_903,In_848);
or U218 (N_218,In_1479,In_473);
xor U219 (N_219,In_1997,In_2603);
nand U220 (N_220,In_1680,In_948);
nand U221 (N_221,In_2733,In_1364);
or U222 (N_222,In_788,In_2010);
nor U223 (N_223,In_2137,In_1180);
nor U224 (N_224,In_1063,In_2872);
nand U225 (N_225,In_2934,In_250);
nand U226 (N_226,In_2832,In_1073);
nand U227 (N_227,In_152,In_2559);
or U228 (N_228,In_26,In_83);
nand U229 (N_229,In_1711,In_2333);
xnor U230 (N_230,In_1216,In_1994);
nand U231 (N_231,In_157,In_256);
nor U232 (N_232,In_301,In_2516);
xnor U233 (N_233,In_13,In_1609);
and U234 (N_234,In_2015,In_1898);
or U235 (N_235,In_2495,In_2866);
nand U236 (N_236,In_1448,In_1118);
nor U237 (N_237,In_992,In_905);
and U238 (N_238,In_2252,In_2343);
and U239 (N_239,In_1050,In_2356);
xor U240 (N_240,In_2553,In_2124);
and U241 (N_241,In_1900,In_659);
nand U242 (N_242,In_2892,In_178);
xor U243 (N_243,In_2910,In_2094);
xnor U244 (N_244,In_266,In_1571);
and U245 (N_245,In_2447,In_819);
and U246 (N_246,In_592,In_1220);
nor U247 (N_247,In_636,In_139);
or U248 (N_248,In_839,In_1460);
and U249 (N_249,In_2111,In_2165);
xnor U250 (N_250,In_712,In_1380);
or U251 (N_251,In_1702,In_1864);
nand U252 (N_252,In_481,In_2518);
or U253 (N_253,In_885,In_1919);
nor U254 (N_254,In_627,In_544);
and U255 (N_255,In_915,In_213);
and U256 (N_256,In_2141,In_998);
nor U257 (N_257,In_734,In_53);
nand U258 (N_258,In_961,In_1878);
or U259 (N_259,In_996,In_902);
and U260 (N_260,In_1899,In_1710);
and U261 (N_261,In_1889,In_1748);
xnor U262 (N_262,In_1947,In_428);
and U263 (N_263,In_2586,In_2357);
nor U264 (N_264,In_1557,In_387);
and U265 (N_265,In_2821,In_911);
and U266 (N_266,In_1985,In_1633);
or U267 (N_267,In_1877,In_2673);
or U268 (N_268,In_934,In_1186);
xnor U269 (N_269,In_2080,In_2855);
and U270 (N_270,In_1250,In_2843);
nor U271 (N_271,In_1601,In_2220);
xnor U272 (N_272,In_840,In_1390);
nor U273 (N_273,In_1869,In_324);
nor U274 (N_274,In_2743,In_1301);
nand U275 (N_275,In_1437,In_1160);
nand U276 (N_276,In_2938,In_2541);
or U277 (N_277,In_421,In_2379);
or U278 (N_278,In_671,In_470);
or U279 (N_279,In_252,In_2476);
xnor U280 (N_280,In_2701,In_2487);
xor U281 (N_281,In_2168,In_1978);
or U282 (N_282,In_973,In_2496);
or U283 (N_283,In_167,In_2090);
nand U284 (N_284,In_31,In_22);
and U285 (N_285,In_2285,In_1276);
xnor U286 (N_286,In_2051,In_1270);
or U287 (N_287,In_838,In_134);
nor U288 (N_288,In_849,In_1498);
xnor U289 (N_289,In_1282,In_163);
or U290 (N_290,In_736,In_960);
nand U291 (N_291,In_1861,In_2183);
nor U292 (N_292,In_2402,In_2410);
nor U293 (N_293,In_2177,In_2665);
and U294 (N_294,In_1697,In_1089);
nor U295 (N_295,In_1379,In_590);
and U296 (N_296,In_2436,In_1853);
or U297 (N_297,In_2316,In_540);
or U298 (N_298,In_488,In_622);
xnor U299 (N_299,In_1766,In_2499);
nand U300 (N_300,In_879,In_2886);
nor U301 (N_301,In_1543,In_717);
nand U302 (N_302,In_1141,In_2528);
nor U303 (N_303,In_11,In_2416);
and U304 (N_304,In_1620,In_881);
nor U305 (N_305,In_1808,In_1444);
xnor U306 (N_306,In_610,In_268);
nor U307 (N_307,In_1799,In_2195);
and U308 (N_308,In_2819,In_2596);
nand U309 (N_309,In_1093,In_395);
or U310 (N_310,In_1429,In_400);
xor U311 (N_311,In_2404,In_672);
or U312 (N_312,In_1475,In_376);
nand U313 (N_313,In_918,In_1984);
or U314 (N_314,In_1419,In_981);
or U315 (N_315,In_299,In_668);
nand U316 (N_316,In_1976,In_858);
xor U317 (N_317,In_2103,In_1687);
or U318 (N_318,In_1389,In_1607);
nor U319 (N_319,In_2767,In_1156);
xnor U320 (N_320,In_1096,In_1178);
and U321 (N_321,In_2942,In_1144);
nand U322 (N_322,In_1348,In_2856);
xnor U323 (N_323,In_2591,In_2612);
or U324 (N_324,In_2719,In_2524);
nand U325 (N_325,In_2083,In_1566);
nor U326 (N_326,In_2732,In_2618);
and U327 (N_327,In_2397,In_1880);
nor U328 (N_328,In_1303,In_87);
and U329 (N_329,In_2149,In_689);
xnor U330 (N_330,In_859,In_941);
or U331 (N_331,In_2229,In_2066);
xnor U332 (N_332,In_2431,In_2477);
or U333 (N_333,In_2981,In_1440);
or U334 (N_334,In_549,In_2475);
and U335 (N_335,In_2868,In_2747);
xnor U336 (N_336,In_1418,In_2079);
and U337 (N_337,In_1391,In_27);
nand U338 (N_338,In_2842,In_1965);
xor U339 (N_339,In_141,In_1646);
and U340 (N_340,In_1350,In_332);
nand U341 (N_341,In_1463,In_1293);
and U342 (N_342,In_2022,In_865);
xor U343 (N_343,In_539,In_1470);
and U344 (N_344,In_39,In_2125);
and U345 (N_345,In_2215,In_986);
nor U346 (N_346,In_1619,In_2583);
nor U347 (N_347,In_493,In_2558);
and U348 (N_348,In_2730,In_1507);
nand U349 (N_349,In_1568,In_1434);
or U350 (N_350,In_2213,In_303);
or U351 (N_351,In_2722,In_1285);
xnor U352 (N_352,In_953,In_2702);
and U353 (N_353,In_2158,In_2479);
nor U354 (N_354,In_426,In_1667);
xor U355 (N_355,In_2639,In_790);
nand U356 (N_356,In_642,In_260);
and U357 (N_357,In_1544,In_218);
xor U358 (N_358,In_1876,In_2978);
or U359 (N_359,In_122,In_643);
nor U360 (N_360,In_793,In_776);
nand U361 (N_361,In_615,In_2236);
and U362 (N_362,In_666,In_640);
and U363 (N_363,In_280,In_2874);
or U364 (N_364,In_1248,In_2894);
and U365 (N_365,In_1484,In_1222);
or U366 (N_366,In_114,In_2128);
nand U367 (N_367,In_1225,In_908);
or U368 (N_368,In_75,In_1807);
nor U369 (N_369,In_1982,In_696);
xor U370 (N_370,In_504,In_207);
and U371 (N_371,In_1360,In_1323);
xor U372 (N_372,In_1509,In_1212);
nor U373 (N_373,In_2616,In_242);
nand U374 (N_374,In_208,In_1185);
nor U375 (N_375,In_1316,In_1231);
xnor U376 (N_376,In_1163,In_675);
nor U377 (N_377,In_1929,In_2350);
nand U378 (N_378,In_2439,In_843);
and U379 (N_379,In_2162,In_1134);
nor U380 (N_380,In_436,In_1975);
xor U381 (N_381,In_136,In_2056);
and U382 (N_382,In_2481,In_2282);
xnor U383 (N_383,In_1809,In_443);
and U384 (N_384,In_912,In_585);
xnor U385 (N_385,In_272,In_2797);
nor U386 (N_386,In_465,In_1608);
or U387 (N_387,In_2268,In_2604);
or U388 (N_388,In_2310,In_1649);
and U389 (N_389,In_1712,In_2900);
nor U390 (N_390,In_449,In_980);
or U391 (N_391,In_1376,In_1797);
nand U392 (N_392,In_322,In_523);
xnor U393 (N_393,In_2523,In_1897);
or U394 (N_394,In_1005,In_2883);
or U395 (N_395,In_67,In_2754);
xor U396 (N_396,In_2960,In_116);
nor U397 (N_397,In_2537,In_1173);
or U398 (N_398,In_2573,In_491);
and U399 (N_399,In_2622,In_2363);
or U400 (N_400,In_1872,In_997);
xnor U401 (N_401,In_764,In_1765);
nor U402 (N_402,In_389,In_4);
xnor U403 (N_403,In_2251,In_1297);
or U404 (N_404,In_95,In_812);
nor U405 (N_405,In_2594,In_117);
or U406 (N_406,In_202,In_2731);
or U407 (N_407,In_2674,In_2547);
nand U408 (N_408,In_1967,In_2672);
xor U409 (N_409,In_2895,In_1955);
nand U410 (N_410,In_174,In_2793);
nor U411 (N_411,In_2844,In_1481);
nand U412 (N_412,In_647,In_417);
or U413 (N_413,In_604,In_145);
xor U414 (N_414,In_625,In_1812);
and U415 (N_415,In_687,In_47);
or U416 (N_416,In_2235,In_1344);
and U417 (N_417,In_517,In_2774);
xnor U418 (N_418,In_576,In_2552);
nor U419 (N_419,In_1943,In_2242);
nand U420 (N_420,In_2663,In_2444);
xnor U421 (N_421,In_1342,In_316);
and U422 (N_422,In_2708,In_1393);
nand U423 (N_423,In_740,In_1242);
xnor U424 (N_424,In_135,In_1757);
xnor U425 (N_425,In_1068,In_2078);
and U426 (N_426,In_2824,In_665);
or U427 (N_427,In_2419,In_1164);
nand U428 (N_428,In_2396,In_989);
nand U429 (N_429,In_1320,In_2157);
or U430 (N_430,In_106,In_2822);
xor U431 (N_431,In_1193,In_1299);
nand U432 (N_432,In_1001,In_429);
or U433 (N_433,In_1695,In_987);
nand U434 (N_434,In_2190,In_1129);
and U435 (N_435,In_177,In_2838);
nor U436 (N_436,In_2773,In_2261);
or U437 (N_437,In_1651,In_406);
xor U438 (N_438,In_2806,In_2948);
nor U439 (N_439,In_1906,In_2928);
nand U440 (N_440,In_168,In_2070);
or U441 (N_441,In_1592,In_962);
nand U442 (N_442,In_462,In_2545);
nor U443 (N_443,In_311,In_846);
and U444 (N_444,In_2432,In_1616);
nand U445 (N_445,In_1629,In_505);
or U446 (N_446,In_2845,In_2077);
nor U447 (N_447,In_2946,In_475);
nand U448 (N_448,In_1315,In_824);
and U449 (N_449,In_1815,In_920);
or U450 (N_450,In_664,In_289);
xor U451 (N_451,In_2561,In_701);
nor U452 (N_452,In_2351,In_2493);
nor U453 (N_453,In_1453,In_1526);
nand U454 (N_454,In_1048,In_2413);
nor U455 (N_455,In_319,In_2707);
or U456 (N_456,In_1774,In_2166);
xnor U457 (N_457,In_528,In_1523);
or U458 (N_458,In_1937,In_97);
nand U459 (N_459,In_1564,In_2606);
xnor U460 (N_460,In_1130,In_2671);
xnor U461 (N_461,In_412,In_2775);
xor U462 (N_462,In_706,In_2974);
nor U463 (N_463,In_2941,In_2870);
or U464 (N_464,In_2640,In_2104);
nor U465 (N_465,In_419,In_2234);
nand U466 (N_466,In_265,In_1501);
nor U467 (N_467,In_1322,In_1485);
nor U468 (N_468,In_482,In_1239);
xor U469 (N_469,In_2693,In_1020);
nor U470 (N_470,In_69,In_2318);
xor U471 (N_471,In_909,In_2852);
and U472 (N_472,In_1402,In_735);
xnor U473 (N_473,In_1558,In_2601);
nand U474 (N_474,In_219,In_2705);
and U475 (N_475,In_1430,In_108);
nand U476 (N_476,In_913,In_531);
xor U477 (N_477,In_2311,In_2112);
nand U478 (N_478,In_1515,In_678);
or U479 (N_479,In_1910,In_2076);
and U480 (N_480,In_2241,In_1204);
nor U481 (N_481,In_1191,In_1587);
and U482 (N_482,In_1795,In_1573);
or U483 (N_483,In_1787,In_802);
or U484 (N_484,In_1030,In_378);
and U485 (N_485,In_2441,In_1510);
nand U486 (N_486,In_919,In_42);
xor U487 (N_487,In_1374,In_1698);
or U488 (N_488,In_340,In_133);
xnor U489 (N_489,In_2102,In_2556);
xor U490 (N_490,In_963,In_1287);
and U491 (N_491,In_2005,In_447);
and U492 (N_492,In_1556,In_1255);
and U493 (N_493,In_1816,In_762);
or U494 (N_494,In_1284,In_1611);
nor U495 (N_495,In_803,In_1378);
nand U496 (N_496,In_286,In_1534);
nand U497 (N_497,In_1626,In_720);
and U498 (N_498,In_1420,In_241);
xnor U499 (N_499,In_1841,In_424);
nor U500 (N_500,In_621,In_2909);
and U501 (N_501,In_715,In_2609);
and U502 (N_502,In_984,In_25);
xnor U503 (N_503,In_20,In_2647);
nand U504 (N_504,In_2314,In_1950);
nor U505 (N_505,In_937,In_1406);
or U506 (N_506,In_595,In_469);
xor U507 (N_507,In_1072,In_2150);
nand U508 (N_508,In_2565,In_453);
nand U509 (N_509,In_749,In_718);
nor U510 (N_510,In_728,In_1638);
nor U511 (N_511,In_2437,In_10);
or U512 (N_512,In_533,In_160);
nor U513 (N_513,In_787,In_1745);
xor U514 (N_514,In_2074,In_1136);
xnor U515 (N_515,In_932,In_1650);
nor U516 (N_516,In_1356,In_274);
nand U517 (N_517,In_1410,In_1451);
or U518 (N_518,In_2725,In_33);
and U519 (N_519,In_1057,In_2989);
or U520 (N_520,In_2201,In_2231);
nand U521 (N_521,In_328,In_2411);
and U522 (N_522,In_2833,In_1690);
nand U523 (N_523,In_614,In_1723);
and U524 (N_524,In_2526,In_2132);
nor U525 (N_525,In_187,In_2169);
nand U526 (N_526,In_1894,In_1346);
or U527 (N_527,In_894,In_2037);
and U528 (N_528,In_1756,In_2631);
nand U529 (N_529,In_1508,In_350);
nand U530 (N_530,In_2390,In_1133);
nand U531 (N_531,In_300,In_1518);
or U532 (N_532,In_1465,In_558);
or U533 (N_533,In_2344,In_420);
or U534 (N_534,In_216,In_525);
or U535 (N_535,In_492,In_1283);
nand U536 (N_536,In_2890,In_2715);
and U537 (N_537,In_1942,In_612);
and U538 (N_538,In_617,In_775);
nand U539 (N_539,In_2689,In_755);
nor U540 (N_540,In_646,In_1613);
nand U541 (N_541,In_1114,In_267);
or U542 (N_542,In_583,In_869);
nand U543 (N_543,In_810,In_2653);
or U544 (N_544,In_15,In_2741);
nand U545 (N_545,In_1905,In_2645);
nor U546 (N_546,In_451,In_818);
nor U547 (N_547,In_34,In_2490);
or U548 (N_548,In_8,In_2638);
or U549 (N_549,In_1761,In_1233);
and U550 (N_550,In_1741,In_2483);
xor U551 (N_551,In_59,In_2283);
and U552 (N_552,In_180,In_1893);
nand U553 (N_553,In_2247,In_2494);
or U554 (N_554,In_124,In_2226);
nor U555 (N_555,In_1887,In_1883);
nor U556 (N_556,In_2240,In_402);
xnor U557 (N_557,In_1701,In_2714);
nor U558 (N_558,In_1142,In_2820);
or U559 (N_559,In_2598,In_1665);
nor U560 (N_560,In_2360,In_1223);
nor U561 (N_561,In_2717,In_284);
nor U562 (N_562,In_569,In_1128);
nor U563 (N_563,In_2392,In_2800);
xor U564 (N_564,In_1439,In_2620);
nand U565 (N_565,In_1078,In_2452);
nand U566 (N_566,In_333,In_526);
or U567 (N_567,In_866,In_2572);
nor U568 (N_568,In_1435,In_2467);
and U569 (N_569,In_1696,In_975);
xor U570 (N_570,In_2664,In_2453);
nand U571 (N_571,In_2658,In_1987);
nor U572 (N_572,In_1553,In_1201);
or U573 (N_573,In_633,In_52);
or U574 (N_574,In_2964,In_2922);
xor U575 (N_575,In_833,In_2828);
xor U576 (N_576,In_1694,In_2760);
and U577 (N_577,In_2293,In_2757);
nand U578 (N_578,In_2349,In_2176);
nand U579 (N_579,In_2801,In_1148);
nor U580 (N_580,In_2847,In_2023);
nor U581 (N_581,In_2950,In_1452);
xor U582 (N_582,In_1836,In_283);
nand U583 (N_583,In_2926,In_1271);
nand U584 (N_584,In_281,In_2237);
or U585 (N_585,In_2173,In_567);
nor U586 (N_586,In_1266,In_2686);
xnor U587 (N_587,In_1355,In_2697);
nand U588 (N_588,In_2057,In_527);
nor U589 (N_589,In_101,In_1550);
xor U590 (N_590,In_194,In_1847);
nand U591 (N_591,In_1398,In_2575);
xor U592 (N_592,In_257,In_2386);
nand U593 (N_593,In_2119,In_1281);
and U594 (N_594,In_1924,In_1599);
xnor U595 (N_595,In_200,In_2859);
xor U596 (N_596,In_226,In_2634);
and U597 (N_597,In_2353,In_2044);
nand U598 (N_598,In_2464,In_1365);
and U599 (N_599,In_1902,In_142);
nand U600 (N_600,In_786,In_2991);
and U601 (N_601,In_1436,In_2042);
nor U602 (N_602,In_2681,In_1324);
xnor U603 (N_603,In_1004,In_2560);
or U604 (N_604,In_649,In_2937);
or U605 (N_605,In_1758,In_2911);
and U606 (N_606,In_454,In_1314);
or U607 (N_607,In_373,In_2578);
xnor U608 (N_608,In_2632,In_1382);
xnor U609 (N_609,In_1062,In_1574);
xnor U610 (N_610,In_2875,In_1536);
or U611 (N_611,In_0,In_1979);
xor U612 (N_612,In_1024,In_1594);
or U613 (N_613,In_1888,In_1739);
nand U614 (N_614,In_1817,In_1487);
and U615 (N_615,In_690,In_502);
or U616 (N_616,In_2118,In_796);
xor U617 (N_617,In_1246,In_32);
and U618 (N_618,In_2017,In_2949);
or U619 (N_619,In_1946,In_503);
or U620 (N_620,In_568,In_644);
xnor U621 (N_621,In_2030,In_1036);
nand U622 (N_622,In_626,In_233);
or U623 (N_623,In_2366,In_1805);
and U624 (N_624,In_1175,In_1228);
nor U625 (N_625,In_1424,In_877);
nor U626 (N_626,In_1995,In_196);
xor U627 (N_627,In_2786,In_2548);
or U628 (N_628,In_1875,In_922);
and U629 (N_629,In_2796,In_2936);
or U630 (N_630,In_486,In_2748);
nor U631 (N_631,In_1635,In_1442);
nor U632 (N_632,In_2977,In_2053);
nor U633 (N_633,In_1736,In_895);
or U634 (N_634,In_561,In_901);
or U635 (N_635,In_1210,In_2580);
nand U636 (N_636,In_1495,In_1217);
and U637 (N_637,In_2313,In_2446);
xor U638 (N_638,In_2997,In_348);
or U639 (N_639,In_166,In_783);
and U640 (N_640,In_602,In_144);
and U641 (N_641,In_1041,In_64);
nor U642 (N_642,In_1262,In_1742);
and U643 (N_643,In_1691,In_1102);
or U644 (N_644,In_2135,In_1923);
nor U645 (N_645,In_18,In_2881);
nand U646 (N_646,In_2889,In_1097);
and U647 (N_647,In_2342,In_7);
and U648 (N_648,In_2138,In_1387);
nor U649 (N_649,In_362,In_1170);
and U650 (N_650,In_2299,In_2643);
and U651 (N_651,In_327,In_1146);
nand U652 (N_652,In_2587,In_2371);
nor U653 (N_653,In_1533,In_1007);
or U654 (N_654,In_1554,In_631);
and U655 (N_655,In_1454,In_2174);
or U656 (N_656,In_1962,In_2491);
nor U657 (N_657,In_2808,In_1933);
xnor U658 (N_658,In_1375,In_2853);
xnor U659 (N_659,In_1395,In_2535);
nand U660 (N_660,In_1703,In_1012);
and U661 (N_661,In_1309,In_104);
nor U662 (N_662,In_1213,In_2203);
xor U663 (N_663,In_550,In_630);
nor U664 (N_664,In_727,In_2046);
nor U665 (N_665,In_904,In_2758);
nand U666 (N_666,In_2320,In_1168);
or U667 (N_667,In_1113,In_2798);
or U668 (N_668,In_1502,In_2407);
xnor U669 (N_669,In_2228,In_1221);
nor U670 (N_670,In_220,In_2519);
nand U671 (N_671,In_2912,In_2685);
nand U672 (N_672,In_864,In_237);
xnor U673 (N_673,In_1480,In_1441);
nand U674 (N_674,In_1081,In_2369);
or U675 (N_675,In_685,In_698);
xnor U676 (N_676,In_269,In_624);
nor U677 (N_677,In_2244,In_1462);
or U678 (N_678,In_103,In_1458);
and U679 (N_679,In_1786,In_1354);
nand U680 (N_680,In_38,In_2315);
and U681 (N_681,In_1127,In_1657);
and U682 (N_682,In_1927,In_2706);
or U683 (N_683,In_2395,In_2337);
nor U684 (N_684,In_771,In_1006);
nor U685 (N_685,In_2877,In_575);
xnor U686 (N_686,In_1604,In_1294);
xnor U687 (N_687,In_1215,In_2266);
nand U688 (N_688,In_1455,In_591);
nor U689 (N_689,In_2971,In_2679);
nor U690 (N_690,In_2644,In_440);
or U691 (N_691,In_2768,In_580);
nor U692 (N_692,In_1981,In_1944);
nor U693 (N_693,In_2059,In_1);
nor U694 (N_694,In_1567,In_1725);
nand U695 (N_695,In_1917,In_2389);
nand U696 (N_696,In_2352,In_302);
nand U697 (N_697,In_2408,In_1265);
xnor U698 (N_698,In_1610,In_2122);
nand U699 (N_699,In_1112,In_2006);
and U700 (N_700,In_217,In_2216);
nor U701 (N_701,In_2026,In_2290);
xnor U702 (N_702,In_1514,In_2255);
nand U703 (N_703,In_781,In_1154);
nand U704 (N_704,In_1743,In_2048);
and U705 (N_705,In_2570,In_1693);
nor U706 (N_706,In_1026,In_2004);
nor U707 (N_707,In_2172,In_789);
and U708 (N_708,In_2795,In_1310);
xnor U709 (N_709,In_1110,In_2492);
or U710 (N_710,In_632,In_1060);
or U711 (N_711,In_854,In_2501);
or U712 (N_712,In_446,In_1825);
and U713 (N_713,In_2429,In_2533);
nor U714 (N_714,In_2952,In_770);
nand U715 (N_715,In_2763,In_2272);
nand U716 (N_716,In_1179,In_63);
and U717 (N_717,In_2649,In_2785);
and U718 (N_718,In_2326,In_243);
and U719 (N_719,In_1977,In_464);
and U720 (N_720,In_797,In_2873);
nand U721 (N_721,In_1971,In_1414);
or U722 (N_722,In_1717,In_2093);
nor U723 (N_723,In_968,In_2101);
nand U724 (N_724,In_403,In_331);
or U725 (N_725,In_679,In_2300);
or U726 (N_726,In_2196,In_652);
xor U727 (N_727,In_195,In_2281);
nor U728 (N_728,In_1615,In_1823);
or U729 (N_729,In_1230,In_801);
or U730 (N_730,In_2267,In_2387);
nand U731 (N_731,In_725,In_596);
or U732 (N_732,In_1912,In_1386);
nand U733 (N_733,In_738,In_35);
nor U734 (N_734,In_1520,In_1226);
or U735 (N_735,In_784,In_2221);
xnor U736 (N_736,In_691,In_1783);
xor U737 (N_737,In_1278,In_2527);
or U738 (N_738,In_1505,In_588);
xor U739 (N_739,In_1957,In_737);
nand U740 (N_740,In_455,In_2454);
xnor U741 (N_741,In_2831,In_88);
and U742 (N_742,In_1319,In_2918);
xnor U743 (N_743,In_457,In_2055);
xnor U744 (N_744,In_1003,In_2134);
nor U745 (N_745,In_2373,In_2049);
nor U746 (N_746,In_73,In_1107);
nand U747 (N_747,In_1575,In_2348);
nand U748 (N_748,In_320,In_1953);
nor U749 (N_749,In_1643,In_555);
or U750 (N_750,In_1956,In_653);
and U751 (N_751,In_566,In_1461);
nand U752 (N_752,In_1038,In_888);
nor U753 (N_753,In_2932,In_2539);
and U754 (N_754,In_2054,In_1486);
xor U755 (N_755,In_936,In_2867);
and U756 (N_756,In_791,In_1777);
xnor U757 (N_757,In_1873,In_1818);
xor U758 (N_758,In_836,In_855);
or U759 (N_759,In_2151,In_1582);
nand U760 (N_760,In_1579,In_2273);
nand U761 (N_761,In_2105,In_228);
nor U762 (N_762,In_1589,In_815);
xor U763 (N_763,In_264,In_98);
nand U764 (N_764,In_2184,In_2144);
nand U765 (N_765,In_158,In_2749);
or U766 (N_766,In_1948,In_868);
nand U767 (N_767,In_416,In_460);
or U768 (N_768,In_1769,In_1152);
xor U769 (N_769,In_2398,In_2625);
xnor U770 (N_770,In_1361,In_2133);
xnor U771 (N_771,In_2099,In_1821);
and U772 (N_772,In_425,In_444);
nor U773 (N_773,In_2372,In_2650);
or U774 (N_774,In_278,In_1174);
or U775 (N_775,In_150,In_1312);
xor U776 (N_776,In_2269,In_2289);
xor U777 (N_777,In_1411,In_164);
xor U778 (N_778,In_1308,In_2286);
xor U779 (N_779,In_2200,In_36);
nand U780 (N_780,In_743,In_1714);
xnor U781 (N_781,In_1802,In_463);
or U782 (N_782,In_510,In_143);
xor U783 (N_783,In_1903,In_1040);
xnor U784 (N_784,In_1234,In_2713);
xor U785 (N_785,In_662,In_1304);
or U786 (N_786,In_1951,In_2557);
nand U787 (N_787,In_1925,In_2325);
or U788 (N_788,In_2790,In_880);
or U789 (N_789,In_2769,In_765);
nor U790 (N_790,In_2189,In_2306);
or U791 (N_791,In_1039,In_1256);
nand U792 (N_792,In_1115,In_1099);
or U793 (N_793,In_538,In_2891);
nor U794 (N_794,In_2794,In_50);
and U795 (N_795,In_1000,In_130);
xor U796 (N_796,In_1837,In_2029);
nand U797 (N_797,In_1776,In_2359);
and U798 (N_798,In_2723,In_2555);
nand U799 (N_799,In_244,In_2648);
nand U800 (N_800,In_2140,In_769);
nand U801 (N_801,In_2551,In_1318);
xnor U802 (N_802,In_1719,In_2849);
and U803 (N_803,In_1474,In_578);
or U804 (N_804,In_2600,In_2905);
nand U805 (N_805,In_1721,In_957);
xor U806 (N_806,In_295,In_380);
nand U807 (N_807,In_1352,In_1596);
xor U808 (N_808,In_2737,In_471);
xnor U809 (N_809,In_115,In_450);
nand U810 (N_810,In_102,In_2549);
nand U811 (N_811,In_1932,In_93);
or U812 (N_812,In_21,In_1939);
and U813 (N_813,In_2430,In_1088);
nor U814 (N_814,In_1844,In_2695);
xnor U815 (N_815,In_1077,In_1670);
nor U816 (N_816,In_1500,In_2906);
xor U817 (N_817,In_374,In_1999);
nand U818 (N_818,In_2256,In_375);
and U819 (N_819,In_2406,In_1647);
or U820 (N_820,In_2335,In_1408);
nand U821 (N_821,In_79,In_2935);
nor U822 (N_822,In_437,In_2961);
nand U823 (N_823,In_1767,In_1238);
and U824 (N_824,In_434,In_1857);
xnor U825 (N_825,In_352,In_2955);
xnor U826 (N_826,In_310,In_112);
or U827 (N_827,In_110,In_2202);
nand U828 (N_828,In_1744,In_41);
or U829 (N_829,In_2529,In_203);
nand U830 (N_830,In_1413,In_2840);
nor U831 (N_831,In_484,In_1018);
or U832 (N_832,In_1686,In_1819);
xor U833 (N_833,In_1833,In_161);
nor U834 (N_834,In_2062,In_1901);
nand U835 (N_835,In_1257,In_2270);
nand U836 (N_836,In_1189,In_940);
and U837 (N_837,In_606,In_1784);
nor U838 (N_838,In_2805,In_2096);
xnor U839 (N_839,In_2507,In_1775);
nor U840 (N_840,In_1116,In_1445);
and U841 (N_841,In_682,In_368);
or U842 (N_842,In_1577,In_6);
or U843 (N_843,In_1070,In_2656);
nand U844 (N_844,In_1664,In_990);
nand U845 (N_845,In_1338,In_1291);
or U846 (N_846,In_884,In_2205);
nor U847 (N_847,In_1669,In_369);
nor U848 (N_848,In_427,In_1724);
and U849 (N_849,In_5,In_1388);
xor U850 (N_850,In_1450,In_1552);
or U851 (N_851,In_2108,In_1019);
or U852 (N_852,In_2985,In_1367);
or U853 (N_853,In_1862,In_2623);
or U854 (N_854,In_778,In_224);
nor U855 (N_855,In_2043,In_2307);
nor U856 (N_856,In_2440,In_271);
and U857 (N_857,In_2687,In_2322);
nor U858 (N_858,In_1022,In_1572);
and U859 (N_859,In_1527,In_171);
and U860 (N_860,In_96,In_1425);
nor U861 (N_861,In_92,In_261);
nand U862 (N_862,In_245,In_907);
nand U863 (N_863,In_1850,In_1618);
xnor U864 (N_864,In_1289,In_2654);
nor U865 (N_865,In_1296,In_1511);
nor U866 (N_866,In_2764,In_179);
nor U867 (N_867,In_1959,In_2690);
nand U868 (N_868,In_2246,In_1295);
or U869 (N_869,In_1302,In_2624);
and U870 (N_870,In_2011,In_342);
nor U871 (N_871,In_409,In_1054);
nor U872 (N_872,In_1083,In_926);
nand U873 (N_873,In_1673,In_1663);
or U874 (N_874,In_1153,In_827);
nand U875 (N_875,In_1337,In_2088);
nor U876 (N_876,In_2277,In_1771);
xnor U877 (N_877,In_2944,In_2544);
or U878 (N_878,In_1126,In_768);
and U879 (N_879,In_2321,In_282);
nand U880 (N_880,In_2295,In_1343);
and U881 (N_881,In_2378,In_1074);
and U882 (N_882,In_105,In_2966);
and U883 (N_883,In_499,In_2700);
and U884 (N_884,In_1904,In_2294);
and U885 (N_885,In_1796,In_490);
nand U886 (N_886,In_2424,In_571);
nand U887 (N_887,In_2739,In_345);
nand U888 (N_888,In_337,In_128);
and U889 (N_889,In_2217,In_519);
or U890 (N_890,In_1151,In_1199);
nand U891 (N_891,In_2885,In_2382);
nor U892 (N_892,In_1037,In_1247);
xor U893 (N_893,In_2250,In_1105);
or U894 (N_894,In_2040,In_1008);
and U895 (N_895,In_1648,In_2211);
nand U896 (N_896,In_2354,In_172);
or U897 (N_897,In_188,In_2914);
nor U898 (N_898,In_2383,In_1208);
nor U899 (N_899,In_656,In_2630);
and U900 (N_900,In_2253,In_731);
xnor U901 (N_901,In_118,In_834);
nor U902 (N_902,In_875,In_1871);
or U903 (N_903,In_60,In_2346);
and U904 (N_904,In_2376,In_2280);
and U905 (N_905,In_2635,In_1532);
xor U906 (N_906,In_1080,In_570);
nor U907 (N_907,In_1991,In_2091);
nand U908 (N_908,In_976,In_1960);
nand U909 (N_909,In_2608,In_1431);
xor U910 (N_910,In_1920,In_496);
and U911 (N_911,In_2271,In_1801);
or U912 (N_912,In_2765,In_1832);
and U913 (N_913,In_1958,In_2208);
and U914 (N_914,In_1279,In_2279);
or U915 (N_915,In_2569,In_1396);
and U916 (N_916,In_2823,In_448);
xor U917 (N_917,In_365,In_2146);
or U918 (N_918,In_2460,In_2682);
nand U919 (N_919,In_2520,In_1229);
nand U920 (N_920,In_2448,In_2098);
or U921 (N_921,In_148,In_2209);
nor U922 (N_922,In_767,In_1103);
and U923 (N_923,In_2907,In_2109);
nor U924 (N_924,In_2084,In_467);
and U925 (N_925,In_2884,In_887);
or U926 (N_926,In_430,In_2745);
xor U927 (N_927,In_231,In_2179);
or U928 (N_928,In_551,In_548);
nand U929 (N_929,In_1521,In_2902);
xnor U930 (N_930,In_2810,In_2879);
and U931 (N_931,In_2462,In_979);
xor U932 (N_932,In_2792,In_2919);
or U933 (N_933,In_249,In_641);
or U934 (N_934,In_1548,In_1042);
or U935 (N_935,In_1986,In_2929);
xor U936 (N_936,In_2455,In_127);
nand U937 (N_937,In_1732,In_1224);
nor U938 (N_938,In_1075,In_547);
nor U939 (N_939,In_30,In_1423);
xnor U940 (N_940,In_2956,In_863);
or U941 (N_941,In_1581,In_1353);
and U942 (N_942,In_1065,In_2092);
or U943 (N_943,In_2442,In_65);
and U944 (N_944,In_2225,In_2777);
nand U945 (N_945,In_192,In_239);
nand U946 (N_946,In_388,In_2347);
or U947 (N_947,In_2142,In_1908);
nor U948 (N_948,In_1881,In_2659);
and U949 (N_949,In_970,In_2434);
xor U950 (N_950,In_2308,In_820);
or U951 (N_951,In_2817,In_1688);
nand U952 (N_952,In_958,In_2085);
nand U953 (N_953,In_1138,In_2621);
nand U954 (N_954,In_1731,In_2362);
nand U955 (N_955,In_2605,In_842);
or U956 (N_956,In_1207,In_2677);
nand U957 (N_957,In_2503,In_1494);
nor U958 (N_958,In_2148,In_413);
xnor U959 (N_959,In_2194,In_537);
or U960 (N_960,In_651,In_432);
nand U961 (N_961,In_466,In_754);
and U962 (N_962,In_1612,In_814);
or U963 (N_963,In_874,In_1918);
nor U964 (N_964,In_1171,In_2751);
nor U965 (N_965,In_954,In_1891);
xnor U966 (N_966,In_361,In_1759);
nor U967 (N_967,In_307,In_703);
xor U968 (N_968,In_1834,In_752);
and U969 (N_969,In_335,In_935);
nand U970 (N_970,In_2193,In_1106);
and U971 (N_971,In_851,In_2506);
nor U972 (N_972,In_2219,In_589);
xnor U973 (N_973,In_2230,In_521);
nand U974 (N_974,In_254,In_1525);
and U975 (N_975,In_2188,In_560);
nor U976 (N_976,In_476,In_1789);
or U977 (N_977,In_2791,In_1131);
and U978 (N_978,In_2031,In_214);
or U979 (N_979,In_1542,In_883);
nor U980 (N_980,In_798,In_2384);
nor U981 (N_981,In_1661,In_262);
and U982 (N_982,In_1829,In_355);
nor U983 (N_983,In_48,In_2538);
or U984 (N_984,In_1313,In_2153);
or U985 (N_985,In_1531,In_2412);
nor U986 (N_986,In_608,In_1591);
or U987 (N_987,In_2486,In_1340);
or U988 (N_988,In_942,In_1738);
and U989 (N_989,In_705,In_190);
xor U990 (N_990,In_2309,In_2035);
xor U991 (N_991,In_1561,In_1349);
xor U992 (N_992,In_2238,In_1804);
nor U993 (N_993,In_2837,In_2365);
xor U994 (N_994,In_2008,In_1580);
xnor U995 (N_995,In_162,In_394);
nor U996 (N_996,In_2018,In_2336);
and U997 (N_997,In_2249,In_2629);
or U998 (N_998,In_2368,In_2032);
and U999 (N_999,In_2381,In_276);
xor U1000 (N_1000,In_2517,In_2951);
or U1001 (N_1001,In_1569,In_346);
or U1002 (N_1002,In_509,In_1492);
nor U1003 (N_1003,In_1049,In_232);
nor U1004 (N_1004,In_2262,In_2428);
xnor U1005 (N_1005,In_1384,In_1538);
xnor U1006 (N_1006,In_1111,In_1249);
nor U1007 (N_1007,In_1268,In_545);
nor U1008 (N_1008,In_2459,In_125);
xnor U1009 (N_1009,In_2013,In_9);
nand U1010 (N_1010,In_2192,In_1496);
nand U1011 (N_1011,In_2531,In_1347);
and U1012 (N_1012,In_2782,In_2522);
or U1013 (N_1013,In_1760,In_1194);
nor U1014 (N_1014,In_229,In_756);
xnor U1015 (N_1015,In_2409,In_442);
xnor U1016 (N_1016,In_28,In_967);
xnor U1017 (N_1017,In_339,In_2933);
or U1018 (N_1018,In_2662,In_2058);
nand U1019 (N_1019,In_165,In_80);
or U1020 (N_1020,In_729,In_2041);
nand U1021 (N_1021,In_1064,In_673);
nand U1022 (N_1022,In_2766,In_2534);
nor U1023 (N_1023,In_1197,In_1357);
nand U1024 (N_1024,In_138,In_1149);
and U1025 (N_1025,In_1737,In_556);
nor U1026 (N_1026,In_2641,In_452);
nor U1027 (N_1027,In_2334,In_2753);
or U1028 (N_1028,In_23,In_1145);
xnor U1029 (N_1029,In_898,In_1839);
nor U1030 (N_1030,In_2016,In_1135);
xnor U1031 (N_1031,In_57,In_2959);
xnor U1032 (N_1032,In_1052,In_2633);
nand U1033 (N_1033,In_856,In_1617);
nor U1034 (N_1034,In_988,In_1644);
or U1035 (N_1035,In_2627,In_1860);
nor U1036 (N_1036,In_1056,In_186);
nor U1037 (N_1037,In_587,In_1464);
or U1038 (N_1038,In_1227,In_317);
or U1039 (N_1039,In_2117,In_1456);
nand U1040 (N_1040,In_1100,In_140);
nor U1041 (N_1041,In_1035,In_211);
or U1042 (N_1042,In_2019,In_2807);
xor U1043 (N_1043,In_1177,In_1438);
and U1044 (N_1044,In_99,In_2367);
nor U1045 (N_1045,In_871,In_2284);
and U1046 (N_1046,In_1964,In_1814);
nand U1047 (N_1047,In_832,In_1913);
nand U1048 (N_1048,In_357,In_563);
nand U1049 (N_1049,In_1762,In_1373);
nand U1050 (N_1050,In_2923,In_230);
xnor U1051 (N_1051,In_2927,In_2052);
nor U1052 (N_1052,In_1327,In_1936);
xor U1053 (N_1053,In_1679,In_24);
nor U1054 (N_1054,In_2712,In_132);
xnor U1055 (N_1055,In_2087,In_1351);
and U1056 (N_1056,In_1466,In_2072);
nand U1057 (N_1057,In_221,In_1263);
or U1058 (N_1058,In_792,In_2976);
xnor U1059 (N_1059,In_1868,In_837);
xor U1060 (N_1060,In_1067,In_497);
nand U1061 (N_1061,In_1763,In_676);
and U1062 (N_1062,In_677,In_1624);
and U1063 (N_1063,In_564,In_206);
and U1064 (N_1064,In_1125,In_238);
nor U1065 (N_1065,In_292,In_248);
xnor U1066 (N_1066,In_1728,In_433);
nor U1067 (N_1067,In_657,In_870);
and U1068 (N_1068,In_541,In_1184);
or U1069 (N_1069,In_1119,In_2470);
nand U1070 (N_1070,In_821,In_1345);
nor U1071 (N_1071,In_2755,In_949);
nand U1072 (N_1072,In_2063,In_2480);
nand U1073 (N_1073,In_247,In_692);
nand U1074 (N_1074,In_2485,In_2564);
nor U1075 (N_1075,In_2020,In_2260);
xor U1076 (N_1076,In_1846,In_385);
nand U1077 (N_1077,In_586,In_2669);
xnor U1078 (N_1078,In_3,In_1335);
or U1079 (N_1079,In_2540,In_1909);
and U1080 (N_1080,In_1489,In_946);
and U1081 (N_1081,In_2497,In_2);
nand U1082 (N_1082,In_1009,In_2655);
nor U1083 (N_1083,In_2000,In_131);
or U1084 (N_1084,In_1468,In_386);
and U1085 (N_1085,In_2871,In_2788);
and U1086 (N_1086,In_2425,In_1940);
xor U1087 (N_1087,In_1659,In_2509);
and U1088 (N_1088,In_1826,In_2903);
or U1089 (N_1089,In_2121,In_1280);
and U1090 (N_1090,In_2947,In_435);
nor U1091 (N_1091,In_2222,In_2858);
and U1092 (N_1092,In_2968,In_2175);
nor U1093 (N_1093,In_1467,In_181);
xor U1094 (N_1094,In_2787,In_2896);
nor U1095 (N_1095,In_742,In_723);
or U1096 (N_1096,In_2857,In_779);
xnor U1097 (N_1097,In_1890,In_393);
or U1098 (N_1098,In_1907,In_2818);
and U1099 (N_1099,In_58,In_1830);
xnor U1100 (N_1100,In_916,In_1027);
and U1101 (N_1101,In_2207,In_852);
nand U1102 (N_1102,In_645,In_2466);
nand U1103 (N_1103,In_2036,In_514);
nor U1104 (N_1104,In_2069,In_694);
or U1105 (N_1105,In_1311,In_78);
or U1106 (N_1106,In_2803,In_182);
nand U1107 (N_1107,In_860,In_629);
or U1108 (N_1108,In_891,In_2908);
nor U1109 (N_1109,In_1874,In_619);
nand U1110 (N_1110,In_2698,In_600);
xnor U1111 (N_1111,In_1588,In_2185);
and U1112 (N_1112,In_500,In_347);
nand U1113 (N_1113,In_2728,In_2198);
or U1114 (N_1114,In_1258,In_2986);
nor U1115 (N_1115,In_472,In_2071);
or U1116 (N_1116,In_1713,In_1606);
nor U1117 (N_1117,In_959,In_2329);
nor U1118 (N_1118,In_2865,In_2258);
and U1119 (N_1119,In_410,In_1852);
nand U1120 (N_1120,In_2691,In_2996);
xor U1121 (N_1121,In_977,In_1662);
or U1122 (N_1122,In_2510,In_1383);
nor U1123 (N_1123,In_1974,In_2403);
and U1124 (N_1124,In_1709,In_1597);
or U1125 (N_1125,In_1930,In_964);
and U1126 (N_1126,In_900,In_2613);
and U1127 (N_1127,In_2405,In_1827);
nor U1128 (N_1128,In_2804,In_2297);
or U1129 (N_1129,In_1540,In_2039);
nor U1130 (N_1130,In_2678,In_1120);
and U1131 (N_1131,In_2917,In_305);
and U1132 (N_1132,In_897,In_209);
xnor U1133 (N_1133,In_557,In_1010);
and U1134 (N_1134,In_1192,In_191);
or U1135 (N_1135,In_969,In_94);
or U1136 (N_1136,In_1854,In_2191);
or U1137 (N_1137,In_2469,In_899);
or U1138 (N_1138,In_1273,In_2904);
nand U1139 (N_1139,In_508,In_1879);
or U1140 (N_1140,In_1562,In_921);
or U1141 (N_1141,In_876,In_1677);
nand U1142 (N_1142,In_2652,In_952);
and U1143 (N_1143,In_1095,In_2550);
xnor U1144 (N_1144,In_1286,In_1272);
nand U1145 (N_1145,In_91,In_695);
or U1146 (N_1146,In_2851,In_461);
nor U1147 (N_1147,In_893,In_1513);
nor U1148 (N_1148,In_2423,In_2116);
or U1149 (N_1149,In_235,In_2740);
and U1150 (N_1150,In_2958,In_813);
nand U1151 (N_1151,In_2562,In_2206);
nand U1152 (N_1152,In_2421,In_2227);
nor U1153 (N_1153,In_955,In_704);
nand U1154 (N_1154,In_1457,In_1549);
xnor U1155 (N_1155,In_372,In_1412);
xor U1156 (N_1156,In_44,In_674);
and U1157 (N_1157,In_804,In_2081);
or U1158 (N_1158,In_599,In_1307);
nand U1159 (N_1159,In_2152,In_1800);
xor U1160 (N_1160,In_2394,In_1397);
xnor U1161 (N_1161,In_931,In_766);
and U1162 (N_1162,In_542,In_1076);
or U1163 (N_1163,In_411,In_2776);
xnor U1164 (N_1164,In_1198,In_2814);
or U1165 (N_1165,In_707,In_2512);
nand U1166 (N_1166,In_2001,In_844);
xor U1167 (N_1167,In_978,In_873);
xor U1168 (N_1168,In_2278,In_2415);
nor U1169 (N_1169,In_1219,In_1169);
nor U1170 (N_1170,In_1584,In_512);
or U1171 (N_1171,In_2021,In_185);
and U1172 (N_1172,In_183,In_51);
and U1173 (N_1173,In_1046,In_290);
and U1174 (N_1174,In_308,In_1858);
nor U1175 (N_1175,In_835,In_2726);
and U1176 (N_1176,In_285,In_2913);
nand U1177 (N_1177,In_1576,In_534);
xnor U1178 (N_1178,In_2401,In_415);
and U1179 (N_1179,In_2100,In_2661);
and U1180 (N_1180,In_273,In_351);
or U1181 (N_1181,In_552,In_2802);
or U1182 (N_1182,In_1885,In_1749);
and U1183 (N_1183,In_1928,In_1840);
xnor U1184 (N_1184,In_1938,In_2264);
or U1185 (N_1185,In_1253,In_72);
or U1186 (N_1186,In_1746,In_637);
nand U1187 (N_1187,In_1427,In_1203);
xor U1188 (N_1188,In_1934,In_1506);
and U1189 (N_1189,In_1377,In_120);
xnor U1190 (N_1190,In_1972,In_2331);
nor U1191 (N_1191,In_1570,In_2953);
or U1192 (N_1192,In_1851,In_951);
or U1193 (N_1193,In_2899,In_2114);
or U1194 (N_1194,In_2014,In_1328);
nand U1195 (N_1195,In_156,In_2998);
or U1196 (N_1196,In_1166,In_474);
and U1197 (N_1197,In_1778,In_1598);
xor U1198 (N_1198,In_1143,In_995);
nor U1199 (N_1199,In_2593,In_2779);
or U1200 (N_1200,In_2592,In_2361);
xor U1201 (N_1201,In_2880,In_2170);
nand U1202 (N_1202,In_1524,In_1206);
nand U1203 (N_1203,In_1288,In_1326);
or U1204 (N_1204,In_2614,In_511);
nor U1205 (N_1205,In_90,In_1416);
nor U1206 (N_1206,In_581,In_982);
xor U1207 (N_1207,In_1630,In_699);
nor U1208 (N_1208,In_1519,In_2120);
nor U1209 (N_1209,In_1645,In_1187);
and U1210 (N_1210,In_726,In_2461);
or U1211 (N_1211,In_2033,In_323);
or U1212 (N_1212,In_1195,In_2505);
nor U1213 (N_1213,In_1071,In_2317);
xnor U1214 (N_1214,In_253,In_422);
and U1215 (N_1215,In_2761,In_2980);
or U1216 (N_1216,In_1368,In_2159);
nor U1217 (N_1217,In_2233,In_2709);
or U1218 (N_1218,In_1123,In_2224);
or U1219 (N_1219,In_2990,In_661);
nor U1220 (N_1220,In_1980,In_1963);
xnor U1221 (N_1221,In_2418,In_862);
xor U1222 (N_1222,In_1025,In_663);
or U1223 (N_1223,In_2154,In_2341);
or U1224 (N_1224,In_2888,In_1915);
nand U1225 (N_1225,In_1504,In_944);
and U1226 (N_1226,In_1157,In_582);
and U1227 (N_1227,In_1886,In_700);
xor U1228 (N_1228,In_2992,In_234);
and U1229 (N_1229,In_1400,In_2097);
or U1230 (N_1230,In_2738,In_760);
nand U1231 (N_1231,In_2915,In_616);
xor U1232 (N_1232,In_2799,In_2759);
nand U1233 (N_1233,In_709,In_2878);
xor U1234 (N_1234,In_270,In_1333);
nor U1235 (N_1235,In_62,In_1631);
nand U1236 (N_1236,In_2670,In_1605);
nand U1237 (N_1237,In_184,In_1988);
or U1238 (N_1238,In_635,In_401);
and U1239 (N_1239,In_2637,In_396);
and U1240 (N_1240,In_349,In_751);
nor U1241 (N_1241,In_660,In_404);
and U1242 (N_1242,In_1779,In_1079);
nand U1243 (N_1243,In_841,In_1090);
xor U1244 (N_1244,In_1092,In_2850);
xnor U1245 (N_1245,In_2445,In_1477);
and U1246 (N_1246,In_620,In_2276);
nand U1247 (N_1247,In_711,In_2716);
or U1248 (N_1248,In_29,In_1813);
nor U1249 (N_1249,In_516,In_2585);
or U1250 (N_1250,In_972,In_199);
xor U1251 (N_1251,In_2199,In_2259);
and U1252 (N_1252,In_2581,In_16);
or U1253 (N_1253,In_1867,In_1636);
and U1254 (N_1254,In_398,In_830);
xnor U1255 (N_1255,In_658,In_805);
or U1256 (N_1256,In_1086,In_914);
and U1257 (N_1257,In_1275,In_325);
or U1258 (N_1258,In_2597,In_1676);
nand U1259 (N_1259,In_2699,In_684);
or U1260 (N_1260,In_1476,In_2107);
and U1261 (N_1261,In_816,In_1683);
xnor U1262 (N_1262,In_1417,In_1708);
xnor U1263 (N_1263,In_2180,In_1642);
nor U1264 (N_1264,In_1583,In_2784);
and U1265 (N_1265,In_2305,In_1706);
and U1266 (N_1266,In_1983,In_2736);
and U1267 (N_1267,In_1449,In_2374);
nand U1268 (N_1268,In_2426,In_808);
nor U1269 (N_1269,In_494,In_605);
nand U1270 (N_1270,In_2839,In_2028);
nor U1271 (N_1271,In_1069,In_1735);
nor U1272 (N_1272,In_1104,In_1055);
or U1273 (N_1273,In_81,In_1045);
or U1274 (N_1274,In_1330,In_2542);
nor U1275 (N_1275,In_2323,In_2781);
xnor U1276 (N_1276,In_1181,In_1321);
xor U1277 (N_1277,In_1482,In_1446);
and U1278 (N_1278,In_259,In_153);
nor U1279 (N_1279,In_2489,In_917);
nor U1280 (N_1280,In_1051,In_546);
or U1281 (N_1281,In_1277,In_2931);
nor U1282 (N_1282,In_1810,In_1806);
nand U1283 (N_1283,In_344,In_2770);
xor U1284 (N_1284,In_638,In_1882);
nor U1285 (N_1285,In_399,In_974);
or U1286 (N_1286,In_2086,In_1392);
xnor U1287 (N_1287,In_483,In_2218);
nand U1288 (N_1288,In_882,In_1363);
nand U1289 (N_1289,In_151,In_2642);
xor U1290 (N_1290,In_831,In_2513);
or U1291 (N_1291,In_498,In_1381);
or U1292 (N_1292,In_850,In_309);
xor U1293 (N_1293,In_2901,In_807);
xnor U1294 (N_1294,In_1622,In_506);
or U1295 (N_1295,In_2339,In_294);
nor U1296 (N_1296,In_1952,In_910);
nand U1297 (N_1297,In_251,In_2239);
and U1298 (N_1298,In_1274,In_2089);
nor U1299 (N_1299,In_2502,In_2710);
xnor U1300 (N_1300,In_2450,In_2963);
and U1301 (N_1301,In_1692,In_2500);
nor U1302 (N_1302,In_354,In_2399);
nor U1303 (N_1303,In_2571,In_334);
nor U1304 (N_1304,In_2465,In_782);
nand U1305 (N_1305,In_811,In_326);
nor U1306 (N_1306,In_721,In_2692);
nor U1307 (N_1307,In_2995,In_1478);
nand U1308 (N_1308,In_2696,In_2554);
and U1309 (N_1309,In_1768,In_291);
xnor U1310 (N_1310,In_2827,In_2862);
xnor U1311 (N_1311,In_1603,In_1831);
nor U1312 (N_1312,In_2611,In_1537);
nor U1313 (N_1313,In_501,In_809);
nand U1314 (N_1314,In_1793,In_1517);
or U1315 (N_1315,In_1856,In_111);
and U1316 (N_1316,In_2456,In_82);
nor U1317 (N_1317,In_2657,In_1835);
or U1318 (N_1318,In_1108,In_170);
or U1319 (N_1319,In_925,In_107);
xor U1320 (N_1320,In_2651,In_84);
nor U1321 (N_1321,In_1949,In_2400);
or U1322 (N_1322,In_1969,In_2988);
nor U1323 (N_1323,In_1147,In_2666);
nor U1324 (N_1324,In_2574,In_929);
xor U1325 (N_1325,In_2813,In_45);
nand U1326 (N_1326,In_2274,In_847);
and U1327 (N_1327,In_246,In_382);
xnor U1328 (N_1328,In_1385,In_2711);
or U1329 (N_1329,In_686,In_2248);
and U1330 (N_1330,In_2288,In_371);
and U1331 (N_1331,In_215,In_2930);
nand U1332 (N_1332,In_1623,In_2422);
nor U1333 (N_1333,In_536,In_1236);
xor U1334 (N_1334,In_2816,In_367);
nand U1335 (N_1335,In_1124,In_543);
and U1336 (N_1336,In_2898,In_1896);
xor U1337 (N_1337,In_939,In_2147);
xor U1338 (N_1338,In_113,In_2752);
or U1339 (N_1339,In_263,In_2388);
xnor U1340 (N_1340,In_1043,In_175);
nor U1341 (N_1341,In_2993,In_2181);
and U1342 (N_1342,In_2789,In_1640);
and U1343 (N_1343,In_2291,In_2983);
or U1344 (N_1344,In_1530,In_2106);
nor U1345 (N_1345,In_2050,In_2265);
nor U1346 (N_1346,In_49,In_2414);
xnor U1347 (N_1347,In_1621,In_2957);
xnor U1348 (N_1348,In_2145,In_628);
and U1349 (N_1349,In_149,In_37);
xnor U1350 (N_1350,In_12,In_1183);
nor U1351 (N_1351,In_2156,In_19);
nand U1352 (N_1352,In_933,In_2292);
xnor U1353 (N_1353,In_1252,In_370);
nand U1354 (N_1354,In_2721,In_2734);
xor U1355 (N_1355,In_1828,In_1634);
nor U1356 (N_1356,In_1359,In_1595);
nand U1357 (N_1357,In_2543,In_2375);
or U1358 (N_1358,In_2836,In_1699);
xor U1359 (N_1359,In_458,In_1497);
nor U1360 (N_1360,In_1137,In_1602);
or U1361 (N_1361,In_2582,In_2068);
or U1362 (N_1362,In_123,In_845);
nor U1363 (N_1363,In_2861,In_2762);
or U1364 (N_1364,In_1264,In_1770);
or U1365 (N_1365,In_2160,In_613);
nor U1366 (N_1366,In_1973,In_109);
nor U1367 (N_1367,In_1172,In_397);
and U1368 (N_1368,In_1290,In_147);
nor U1369 (N_1369,In_1681,In_85);
and U1370 (N_1370,In_654,In_2245);
xor U1371 (N_1371,In_46,In_683);
nand U1372 (N_1372,In_1678,In_2113);
and U1373 (N_1373,In_2002,In_2025);
and U1374 (N_1374,In_1235,In_1734);
or U1375 (N_1375,In_225,In_1682);
nor U1376 (N_1376,In_1061,In_1267);
or U1377 (N_1377,In_2330,In_565);
nor U1378 (N_1378,In_2515,In_518);
or U1379 (N_1379,In_313,In_2139);
and U1380 (N_1380,In_950,In_878);
nor U1381 (N_1381,In_1260,In_1016);
xnor U1382 (N_1382,In_329,In_1240);
nand U1383 (N_1383,In_1792,In_2577);
or U1384 (N_1384,In_2508,In_2675);
or U1385 (N_1385,In_2073,In_2009);
nor U1386 (N_1386,In_2965,In_2595);
xnor U1387 (N_1387,In_826,In_2171);
nor U1388 (N_1388,In_2683,In_137);
nand U1389 (N_1389,In_100,In_77);
xnor U1390 (N_1390,In_739,In_2319);
nor U1391 (N_1391,In_2143,In_223);
nand U1392 (N_1392,In_1325,In_2778);
nor U1393 (N_1393,In_1968,In_1094);
or U1394 (N_1394,In_2916,In_2161);
nor U1395 (N_1395,In_708,In_2967);
nor U1396 (N_1396,In_212,In_1730);
nor U1397 (N_1397,In_573,In_1656);
or U1398 (N_1398,In_1996,In_56);
and U1399 (N_1399,In_353,In_1585);
xor U1400 (N_1400,In_2532,In_338);
and U1401 (N_1401,In_702,In_2186);
nand U1402 (N_1402,In_1849,In_1790);
nor U1403 (N_1403,In_1628,In_1718);
and U1404 (N_1404,In_515,In_991);
or U1405 (N_1405,In_2067,In_1914);
nor U1406 (N_1406,In_2718,In_330);
xor U1407 (N_1407,In_121,In_1722);
or U1408 (N_1408,In_1167,In_2727);
nand U1409 (N_1409,In_2771,In_777);
and U1410 (N_1410,In_321,In_198);
xor U1411 (N_1411,In_487,In_477);
and U1412 (N_1412,In_2210,In_2127);
nand U1413 (N_1413,In_89,In_2324);
nand U1414 (N_1414,In_1028,In_2178);
or U1415 (N_1415,In_714,In_2298);
nand U1416 (N_1416,In_1488,In_126);
nand U1417 (N_1417,In_1754,In_1522);
nand U1418 (N_1418,In_2064,In_697);
nor U1419 (N_1419,In_2704,In_1218);
nor U1420 (N_1420,In_1066,In_2478);
nand U1421 (N_1421,In_1727,In_2780);
nor U1422 (N_1422,In_2979,In_297);
and U1423 (N_1423,In_1370,In_1704);
or U1424 (N_1424,In_1824,In_2848);
and U1425 (N_1425,In_408,In_1161);
or U1426 (N_1426,In_2130,In_750);
xor U1427 (N_1427,In_1551,In_2438);
nand U1428 (N_1428,In_1469,In_1306);
nand U1429 (N_1429,In_1058,In_1200);
or U1430 (N_1430,In_358,In_1822);
xnor U1431 (N_1431,In_1002,In_68);
nor U1432 (N_1432,In_966,In_2391);
nand U1433 (N_1433,In_227,In_1752);
or U1434 (N_1434,In_298,In_431);
or U1435 (N_1435,In_1117,In_872);
or U1436 (N_1436,In_2263,In_1863);
or U1437 (N_1437,In_2920,In_1331);
or U1438 (N_1438,In_2024,In_2364);
nor U1439 (N_1439,In_1122,In_1990);
or U1440 (N_1440,In_1559,In_759);
nor U1441 (N_1441,In_1336,In_597);
nor U1442 (N_1442,In_680,In_480);
or U1443 (N_1443,In_2954,In_1190);
xor U1444 (N_1444,In_1781,In_896);
xnor U1445 (N_1445,In_1685,In_1405);
or U1446 (N_1446,In_1921,In_392);
or U1447 (N_1447,In_757,In_648);
or U1448 (N_1448,In_716,In_667);
nand U1449 (N_1449,In_2471,In_1716);
xnor U1450 (N_1450,In_1339,In_2825);
xor U1451 (N_1451,In_1992,In_1422);
or U1452 (N_1452,In_2834,In_2458);
xor U1453 (N_1453,In_562,In_2047);
or U1454 (N_1454,In_1259,In_485);
or U1455 (N_1455,In_1503,In_423);
nor U1456 (N_1456,In_2115,In_2182);
nor U1457 (N_1457,In_744,In_2610);
or U1458 (N_1458,In_1671,In_1162);
xor U1459 (N_1459,In_1176,In_2155);
nand U1460 (N_1460,In_1586,In_1675);
xor U1461 (N_1461,In_2994,In_1084);
xor U1462 (N_1462,In_607,In_747);
or U1463 (N_1463,In_2303,In_748);
nand U1464 (N_1464,In_2829,In_2340);
nor U1465 (N_1465,In_1590,In_2756);
nand U1466 (N_1466,In_414,In_2973);
xnor U1467 (N_1467,In_381,In_2724);
nor U1468 (N_1468,In_681,In_1196);
nor U1469 (N_1469,In_572,In_985);
and U1470 (N_1470,In_1205,In_965);
nand U1471 (N_1471,In_1755,In_1911);
nand U1472 (N_1472,In_2744,In_1132);
or U1473 (N_1473,In_553,In_2332);
or U1474 (N_1474,In_2897,In_2075);
nor U1475 (N_1475,In_1399,In_1269);
nor U1476 (N_1476,In_2617,In_1726);
or U1477 (N_1477,In_774,In_2482);
or U1478 (N_1478,In_650,In_559);
and U1479 (N_1479,In_1747,In_155);
xor U1480 (N_1480,In_794,In_1764);
xor U1481 (N_1481,In_785,In_1098);
nor U1482 (N_1482,In_730,In_2982);
and U1483 (N_1483,In_1655,In_1627);
and U1484 (N_1484,In_2972,In_390);
or U1485 (N_1485,In_1371,In_2809);
and U1486 (N_1486,In_2472,In_288);
xor U1487 (N_1487,In_825,In_1720);
or U1488 (N_1488,In_1158,In_1658);
and U1489 (N_1489,In_923,In_2034);
nor U1490 (N_1490,In_2451,In_459);
xnor U1491 (N_1491,In_2846,In_1529);
or U1492 (N_1492,In_780,In_468);
nor U1493 (N_1493,In_1859,In_1394);
or U1494 (N_1494,In_1578,In_594);
or U1495 (N_1495,In_1547,In_2449);
and U1496 (N_1496,In_2962,In_1654);
and U1497 (N_1497,In_763,In_554);
xnor U1498 (N_1498,In_1432,In_2488);
or U1499 (N_1499,In_2720,In_1838);
nor U1500 (N_1500,N_807,N_348);
xnor U1501 (N_1501,N_474,N_427);
or U1502 (N_1502,N_38,N_167);
nand U1503 (N_1503,N_1437,N_1009);
or U1504 (N_1504,N_1232,N_557);
xor U1505 (N_1505,N_859,N_1261);
xor U1506 (N_1506,N_1378,N_967);
and U1507 (N_1507,N_1499,N_892);
nand U1508 (N_1508,N_1176,N_639);
or U1509 (N_1509,N_975,N_1159);
or U1510 (N_1510,N_828,N_676);
xor U1511 (N_1511,N_624,N_784);
nor U1512 (N_1512,N_308,N_121);
xor U1513 (N_1513,N_223,N_480);
nand U1514 (N_1514,N_638,N_1097);
nor U1515 (N_1515,N_1197,N_996);
nand U1516 (N_1516,N_969,N_176);
xnor U1517 (N_1517,N_171,N_469);
and U1518 (N_1518,N_612,N_1396);
nor U1519 (N_1519,N_491,N_375);
nor U1520 (N_1520,N_725,N_622);
xor U1521 (N_1521,N_572,N_1069);
nand U1522 (N_1522,N_540,N_472);
xnor U1523 (N_1523,N_819,N_201);
nor U1524 (N_1524,N_388,N_426);
xnor U1525 (N_1525,N_1138,N_113);
or U1526 (N_1526,N_221,N_1257);
nand U1527 (N_1527,N_497,N_629);
xor U1528 (N_1528,N_988,N_157);
or U1529 (N_1529,N_724,N_900);
or U1530 (N_1530,N_92,N_991);
xnor U1531 (N_1531,N_1276,N_6);
or U1532 (N_1532,N_775,N_1120);
or U1533 (N_1533,N_1199,N_119);
xor U1534 (N_1534,N_267,N_192);
or U1535 (N_1535,N_899,N_492);
or U1536 (N_1536,N_1476,N_1479);
and U1537 (N_1537,N_760,N_650);
nand U1538 (N_1538,N_815,N_610);
nand U1539 (N_1539,N_708,N_50);
and U1540 (N_1540,N_1484,N_1077);
xor U1541 (N_1541,N_931,N_562);
nor U1542 (N_1542,N_100,N_1130);
and U1543 (N_1543,N_317,N_408);
xor U1544 (N_1544,N_1353,N_404);
and U1545 (N_1545,N_1423,N_243);
nand U1546 (N_1546,N_438,N_142);
nor U1547 (N_1547,N_1103,N_894);
xor U1548 (N_1548,N_1147,N_1288);
and U1549 (N_1549,N_699,N_1182);
and U1550 (N_1550,N_318,N_1254);
or U1551 (N_1551,N_282,N_701);
nor U1552 (N_1552,N_919,N_1487);
and U1553 (N_1553,N_358,N_65);
nor U1554 (N_1554,N_290,N_212);
or U1555 (N_1555,N_1436,N_226);
nand U1556 (N_1556,N_1498,N_1319);
or U1557 (N_1557,N_588,N_983);
or U1558 (N_1558,N_865,N_94);
nand U1559 (N_1559,N_538,N_999);
nor U1560 (N_1560,N_889,N_1128);
or U1561 (N_1561,N_286,N_233);
nor U1562 (N_1562,N_873,N_1421);
nand U1563 (N_1563,N_867,N_347);
or U1564 (N_1564,N_1329,N_1340);
nor U1565 (N_1565,N_911,N_1102);
or U1566 (N_1566,N_431,N_1286);
xor U1567 (N_1567,N_687,N_683);
nor U1568 (N_1568,N_1156,N_989);
and U1569 (N_1569,N_742,N_1282);
or U1570 (N_1570,N_1037,N_1101);
nor U1571 (N_1571,N_1453,N_102);
or U1572 (N_1572,N_583,N_363);
nor U1573 (N_1573,N_755,N_688);
nand U1574 (N_1574,N_723,N_9);
nand U1575 (N_1575,N_934,N_1265);
and U1576 (N_1576,N_1461,N_647);
and U1577 (N_1577,N_1287,N_488);
xor U1578 (N_1578,N_168,N_325);
or U1579 (N_1579,N_806,N_169);
nand U1580 (N_1580,N_501,N_1110);
nor U1581 (N_1581,N_1162,N_1115);
and U1582 (N_1582,N_643,N_385);
or U1583 (N_1583,N_662,N_916);
xnor U1584 (N_1584,N_72,N_1180);
nor U1585 (N_1585,N_679,N_703);
or U1586 (N_1586,N_37,N_231);
xor U1587 (N_1587,N_1055,N_473);
and U1588 (N_1588,N_939,N_752);
and U1589 (N_1589,N_978,N_493);
nor U1590 (N_1590,N_1035,N_834);
and U1591 (N_1591,N_147,N_332);
or U1592 (N_1592,N_1173,N_1087);
xor U1593 (N_1593,N_494,N_389);
nor U1594 (N_1594,N_864,N_710);
nor U1595 (N_1595,N_467,N_543);
xor U1596 (N_1596,N_1377,N_686);
and U1597 (N_1597,N_448,N_955);
or U1598 (N_1598,N_526,N_536);
xnor U1599 (N_1599,N_402,N_26);
and U1600 (N_1600,N_1227,N_1043);
xnor U1601 (N_1601,N_1370,N_44);
or U1602 (N_1602,N_1480,N_707);
and U1603 (N_1603,N_773,N_1497);
xor U1604 (N_1604,N_35,N_40);
and U1605 (N_1605,N_81,N_1408);
nand U1606 (N_1606,N_1252,N_531);
xor U1607 (N_1607,N_246,N_1374);
and U1608 (N_1608,N_523,N_407);
nand U1609 (N_1609,N_146,N_1468);
and U1610 (N_1610,N_258,N_613);
or U1611 (N_1611,N_125,N_596);
nand U1612 (N_1612,N_152,N_740);
and U1613 (N_1613,N_929,N_1493);
and U1614 (N_1614,N_387,N_257);
nand U1615 (N_1615,N_617,N_188);
xor U1616 (N_1616,N_750,N_165);
nand U1617 (N_1617,N_605,N_981);
nor U1618 (N_1618,N_558,N_547);
nor U1619 (N_1619,N_1414,N_933);
nor U1620 (N_1620,N_598,N_1268);
or U1621 (N_1621,N_817,N_554);
or U1622 (N_1622,N_396,N_93);
nor U1623 (N_1623,N_297,N_1417);
nand U1624 (N_1624,N_1256,N_1153);
nor U1625 (N_1625,N_261,N_1089);
and U1626 (N_1626,N_651,N_735);
nand U1627 (N_1627,N_365,N_1312);
or U1628 (N_1628,N_832,N_972);
or U1629 (N_1629,N_1072,N_449);
nand U1630 (N_1630,N_1333,N_454);
or U1631 (N_1631,N_403,N_277);
and U1632 (N_1632,N_225,N_544);
nor U1633 (N_1633,N_529,N_1415);
or U1634 (N_1634,N_938,N_684);
nand U1635 (N_1635,N_1241,N_163);
and U1636 (N_1636,N_1191,N_1220);
nor U1637 (N_1637,N_115,N_1290);
xnor U1638 (N_1638,N_640,N_542);
nand U1639 (N_1639,N_1066,N_1126);
or U1640 (N_1640,N_809,N_191);
nor U1641 (N_1641,N_421,N_127);
nor U1642 (N_1642,N_1057,N_781);
or U1643 (N_1643,N_508,N_112);
and U1644 (N_1644,N_611,N_56);
or U1645 (N_1645,N_868,N_1401);
and U1646 (N_1646,N_377,N_253);
and U1647 (N_1647,N_334,N_17);
nand U1648 (N_1648,N_757,N_133);
xor U1649 (N_1649,N_57,N_355);
xnor U1650 (N_1650,N_1008,N_1451);
nand U1651 (N_1651,N_672,N_218);
and U1652 (N_1652,N_450,N_581);
or U1653 (N_1653,N_953,N_1140);
nor U1654 (N_1654,N_1085,N_664);
and U1655 (N_1655,N_266,N_1091);
and U1656 (N_1656,N_875,N_1016);
nor U1657 (N_1657,N_685,N_534);
or U1658 (N_1658,N_1114,N_1381);
nand U1659 (N_1659,N_810,N_994);
nor U1660 (N_1660,N_578,N_974);
and U1661 (N_1661,N_76,N_1178);
nand U1662 (N_1662,N_291,N_459);
and U1663 (N_1663,N_495,N_1064);
nand U1664 (N_1664,N_522,N_1029);
and U1665 (N_1665,N_1174,N_1026);
nand U1666 (N_1666,N_310,N_719);
nand U1667 (N_1667,N_177,N_1071);
nor U1668 (N_1668,N_971,N_949);
xnor U1669 (N_1669,N_808,N_270);
nor U1670 (N_1670,N_213,N_682);
nor U1671 (N_1671,N_855,N_1465);
nor U1672 (N_1672,N_259,N_88);
or U1673 (N_1673,N_759,N_1045);
or U1674 (N_1674,N_656,N_877);
xnor U1675 (N_1675,N_843,N_97);
and U1676 (N_1676,N_1247,N_1053);
xnor U1677 (N_1677,N_1216,N_432);
or U1678 (N_1678,N_1221,N_1320);
and U1679 (N_1679,N_1013,N_715);
xor U1680 (N_1680,N_354,N_813);
or U1681 (N_1681,N_1019,N_1135);
xnor U1682 (N_1682,N_736,N_446);
nor U1683 (N_1683,N_1107,N_1278);
nand U1684 (N_1684,N_345,N_694);
or U1685 (N_1685,N_1244,N_1306);
and U1686 (N_1686,N_696,N_462);
and U1687 (N_1687,N_1277,N_1148);
and U1688 (N_1688,N_304,N_546);
nand U1689 (N_1689,N_1006,N_331);
nor U1690 (N_1690,N_1410,N_533);
nand U1691 (N_1691,N_222,N_392);
nand U1692 (N_1692,N_32,N_1127);
xnor U1693 (N_1693,N_1389,N_1462);
nor U1694 (N_1694,N_795,N_437);
nor U1695 (N_1695,N_1235,N_1266);
and U1696 (N_1696,N_1169,N_433);
and U1697 (N_1697,N_730,N_909);
nor U1698 (N_1698,N_132,N_1406);
nand U1699 (N_1699,N_316,N_573);
nand U1700 (N_1700,N_1084,N_1482);
or U1701 (N_1701,N_824,N_965);
and U1702 (N_1702,N_393,N_61);
nor U1703 (N_1703,N_1022,N_1050);
nand U1704 (N_1704,N_772,N_545);
or U1705 (N_1705,N_794,N_214);
nand U1706 (N_1706,N_768,N_1407);
nand U1707 (N_1707,N_884,N_893);
xnor U1708 (N_1708,N_504,N_681);
and U1709 (N_1709,N_702,N_591);
or U1710 (N_1710,N_926,N_879);
nor U1711 (N_1711,N_509,N_209);
or U1712 (N_1712,N_729,N_1295);
and U1713 (N_1713,N_475,N_85);
and U1714 (N_1714,N_164,N_1212);
nand U1715 (N_1715,N_1070,N_568);
nand U1716 (N_1716,N_1202,N_232);
nor U1717 (N_1717,N_771,N_942);
and U1718 (N_1718,N_138,N_663);
xor U1719 (N_1719,N_306,N_276);
and U1720 (N_1720,N_1004,N_1308);
nor U1721 (N_1721,N_766,N_745);
nor U1722 (N_1722,N_977,N_587);
or U1723 (N_1723,N_27,N_1263);
xor U1724 (N_1724,N_917,N_1301);
or U1725 (N_1725,N_626,N_296);
xor U1726 (N_1726,N_770,N_1023);
or U1727 (N_1727,N_287,N_511);
and U1728 (N_1728,N_1291,N_67);
nor U1729 (N_1729,N_985,N_1002);
and U1730 (N_1730,N_1420,N_1284);
xor U1731 (N_1731,N_930,N_273);
nand U1732 (N_1732,N_976,N_295);
and U1733 (N_1733,N_1455,N_1151);
nor U1734 (N_1734,N_507,N_42);
xnor U1735 (N_1735,N_762,N_284);
nor U1736 (N_1736,N_1303,N_799);
and U1737 (N_1737,N_269,N_886);
and U1738 (N_1738,N_1296,N_1096);
or U1739 (N_1739,N_635,N_689);
nor U1740 (N_1740,N_829,N_553);
and U1741 (N_1741,N_48,N_445);
nand U1742 (N_1742,N_122,N_1356);
nor U1743 (N_1743,N_1100,N_444);
or U1744 (N_1744,N_698,N_12);
nor U1745 (N_1745,N_1446,N_39);
xor U1746 (N_1746,N_761,N_199);
nor U1747 (N_1747,N_1259,N_118);
or U1748 (N_1748,N_1167,N_371);
and U1749 (N_1749,N_1020,N_1366);
or U1750 (N_1750,N_1113,N_461);
and U1751 (N_1751,N_1217,N_45);
nor U1752 (N_1752,N_139,N_1334);
or U1753 (N_1753,N_846,N_1478);
nand U1754 (N_1754,N_453,N_227);
and U1755 (N_1755,N_751,N_585);
nand U1756 (N_1756,N_874,N_567);
and U1757 (N_1757,N_614,N_1049);
nor U1758 (N_1758,N_344,N_435);
and U1759 (N_1759,N_872,N_47);
nand U1760 (N_1760,N_64,N_615);
nor U1761 (N_1761,N_1387,N_856);
nor U1762 (N_1762,N_506,N_1394);
and U1763 (N_1763,N_293,N_1088);
or U1764 (N_1764,N_255,N_1248);
and U1765 (N_1765,N_1208,N_619);
xnor U1766 (N_1766,N_99,N_1357);
and U1767 (N_1767,N_1315,N_1324);
or U1768 (N_1768,N_441,N_620);
or U1769 (N_1769,N_1015,N_219);
nand U1770 (N_1770,N_1444,N_1490);
nand U1771 (N_1771,N_1211,N_346);
and U1772 (N_1772,N_1441,N_527);
xor U1773 (N_1773,N_324,N_593);
nor U1774 (N_1774,N_822,N_60);
and U1775 (N_1775,N_519,N_1433);
nor U1776 (N_1776,N_1367,N_123);
or U1777 (N_1777,N_1052,N_1158);
or U1778 (N_1778,N_1432,N_1093);
nor U1779 (N_1779,N_1005,N_263);
nor U1780 (N_1780,N_1166,N_870);
nor U1781 (N_1781,N_607,N_311);
nor U1782 (N_1782,N_186,N_636);
nor U1783 (N_1783,N_55,N_3);
nand U1784 (N_1784,N_466,N_1483);
and U1785 (N_1785,N_162,N_1112);
or U1786 (N_1786,N_412,N_1350);
nand U1787 (N_1787,N_2,N_236);
nor U1788 (N_1788,N_1046,N_764);
xor U1789 (N_1789,N_950,N_1225);
xor U1790 (N_1790,N_505,N_642);
and U1791 (N_1791,N_1054,N_1214);
nor U1792 (N_1792,N_776,N_1335);
nor U1793 (N_1793,N_14,N_734);
xnor U1794 (N_1794,N_555,N_747);
nor U1795 (N_1795,N_941,N_185);
xnor U1796 (N_1796,N_997,N_78);
nor U1797 (N_1797,N_357,N_53);
nor U1798 (N_1798,N_1352,N_604);
nor U1799 (N_1799,N_535,N_802);
xnor U1800 (N_1800,N_1477,N_992);
xor U1801 (N_1801,N_43,N_584);
or U1802 (N_1802,N_849,N_1003);
xnor U1803 (N_1803,N_722,N_63);
xnor U1804 (N_1804,N_486,N_33);
and U1805 (N_1805,N_1203,N_8);
and U1806 (N_1806,N_230,N_1419);
nor U1807 (N_1807,N_630,N_1342);
nor U1808 (N_1808,N_924,N_1375);
or U1809 (N_1809,N_420,N_732);
nor U1810 (N_1810,N_204,N_1273);
and U1811 (N_1811,N_111,N_264);
or U1812 (N_1812,N_928,N_1348);
nor U1813 (N_1813,N_1080,N_1231);
xor U1814 (N_1814,N_340,N_811);
nand U1815 (N_1815,N_600,N_837);
xor U1816 (N_1816,N_397,N_1243);
or U1817 (N_1817,N_1226,N_691);
and U1818 (N_1818,N_1068,N_831);
and U1819 (N_1819,N_1144,N_1213);
nand U1820 (N_1820,N_803,N_240);
or U1821 (N_1821,N_460,N_743);
xnor U1822 (N_1822,N_1382,N_305);
or U1823 (N_1823,N_851,N_31);
nand U1824 (N_1824,N_395,N_418);
nand U1825 (N_1825,N_179,N_341);
nand U1826 (N_1826,N_825,N_183);
nand U1827 (N_1827,N_279,N_915);
xnor U1828 (N_1828,N_71,N_947);
and U1829 (N_1829,N_87,N_128);
nand U1830 (N_1830,N_484,N_1474);
or U1831 (N_1831,N_844,N_1338);
xor U1832 (N_1832,N_1081,N_883);
or U1833 (N_1833,N_4,N_1336);
xnor U1834 (N_1834,N_381,N_373);
nor U1835 (N_1835,N_549,N_510);
and U1836 (N_1836,N_439,N_1179);
and U1837 (N_1837,N_487,N_1402);
xor U1838 (N_1838,N_816,N_623);
xor U1839 (N_1839,N_13,N_443);
nand U1840 (N_1840,N_912,N_866);
and U1841 (N_1841,N_559,N_1397);
xnor U1842 (N_1842,N_602,N_1404);
or U1843 (N_1843,N_1351,N_1302);
and U1844 (N_1844,N_1447,N_590);
nand U1845 (N_1845,N_673,N_289);
and U1846 (N_1846,N_890,N_1160);
nand U1847 (N_1847,N_0,N_1428);
nor U1848 (N_1848,N_841,N_979);
nor U1849 (N_1849,N_181,N_338);
and U1850 (N_1850,N_1272,N_1466);
nand U1851 (N_1851,N_1125,N_116);
nand U1852 (N_1852,N_500,N_1289);
or U1853 (N_1853,N_1000,N_1354);
or U1854 (N_1854,N_717,N_1237);
nand U1855 (N_1855,N_1429,N_1403);
nor U1856 (N_1856,N_158,N_1281);
nor U1857 (N_1857,N_1106,N_1234);
and U1858 (N_1858,N_1327,N_54);
nand U1859 (N_1859,N_172,N_1021);
nand U1860 (N_1860,N_1017,N_927);
nor U1861 (N_1861,N_1349,N_958);
xor U1862 (N_1862,N_897,N_1196);
nand U1863 (N_1863,N_1413,N_1481);
and U1864 (N_1864,N_1332,N_173);
nor U1865 (N_1865,N_838,N_1164);
and U1866 (N_1866,N_1369,N_970);
nor U1867 (N_1867,N_28,N_1230);
and U1868 (N_1868,N_1337,N_798);
and U1869 (N_1869,N_1347,N_1393);
xnor U1870 (N_1870,N_262,N_1260);
nor U1871 (N_1871,N_203,N_582);
or U1872 (N_1872,N_1238,N_320);
and U1873 (N_1873,N_1297,N_780);
or U1874 (N_1874,N_881,N_1031);
or U1875 (N_1875,N_1470,N_69);
nor U1876 (N_1876,N_1385,N_987);
xnor U1877 (N_1877,N_1326,N_108);
or U1878 (N_1878,N_211,N_921);
xor U1879 (N_1879,N_737,N_1090);
and U1880 (N_1880,N_657,N_1034);
nand U1881 (N_1881,N_1137,N_913);
nand U1882 (N_1882,N_1450,N_1109);
nand U1883 (N_1883,N_465,N_973);
or U1884 (N_1884,N_812,N_260);
and U1885 (N_1885,N_1108,N_335);
xnor U1886 (N_1886,N_46,N_902);
xnor U1887 (N_1887,N_944,N_1434);
and U1888 (N_1888,N_1078,N_370);
xnor U1889 (N_1889,N_34,N_1359);
nor U1890 (N_1890,N_659,N_1274);
nor U1891 (N_1891,N_552,N_386);
and U1892 (N_1892,N_83,N_337);
or U1893 (N_1893,N_1345,N_485);
nor U1894 (N_1894,N_763,N_787);
nor U1895 (N_1895,N_399,N_423);
or U1896 (N_1896,N_1449,N_490);
and U1897 (N_1897,N_790,N_599);
or U1898 (N_1898,N_272,N_914);
and U1899 (N_1899,N_871,N_1012);
and U1900 (N_1900,N_1343,N_709);
xnor U1901 (N_1901,N_1188,N_948);
and U1902 (N_1902,N_1111,N_592);
xor U1903 (N_1903,N_369,N_1067);
nand U1904 (N_1904,N_654,N_109);
or U1905 (N_1905,N_966,N_525);
nor U1906 (N_1906,N_208,N_782);
nand U1907 (N_1907,N_419,N_714);
nor U1908 (N_1908,N_134,N_398);
or U1909 (N_1909,N_36,N_1205);
or U1910 (N_1910,N_577,N_792);
xor U1911 (N_1911,N_1376,N_731);
or U1912 (N_1912,N_247,N_1250);
xnor U1913 (N_1913,N_721,N_1355);
and U1914 (N_1914,N_1494,N_268);
nand U1915 (N_1915,N_11,N_51);
nor U1916 (N_1916,N_405,N_29);
nand U1917 (N_1917,N_597,N_406);
and U1918 (N_1918,N_993,N_190);
and U1919 (N_1919,N_1424,N_512);
nand U1920 (N_1920,N_1118,N_922);
xor U1921 (N_1921,N_561,N_910);
nand U1922 (N_1922,N_1195,N_514);
nor U1923 (N_1923,N_23,N_479);
xor U1924 (N_1924,N_326,N_197);
nand U1925 (N_1925,N_595,N_288);
nand U1926 (N_1926,N_52,N_248);
xor U1927 (N_1927,N_458,N_321);
nand U1928 (N_1928,N_235,N_1360);
nand U1929 (N_1929,N_130,N_678);
nor U1930 (N_1930,N_1439,N_1001);
or U1931 (N_1931,N_1042,N_1218);
xor U1932 (N_1932,N_603,N_1300);
and U1933 (N_1933,N_1007,N_1253);
xnor U1934 (N_1934,N_323,N_178);
nor U1935 (N_1935,N_476,N_66);
nand U1936 (N_1936,N_789,N_1092);
nand U1937 (N_1937,N_136,N_1467);
and U1938 (N_1938,N_1391,N_1422);
xnor U1939 (N_1939,N_895,N_563);
nand U1940 (N_1940,N_677,N_452);
xnor U1941 (N_1941,N_1177,N_954);
or U1942 (N_1942,N_104,N_1489);
nor U1943 (N_1943,N_241,N_957);
nor U1944 (N_1944,N_1242,N_470);
and U1945 (N_1945,N_379,N_150);
and U1946 (N_1946,N_1361,N_1027);
and U1947 (N_1947,N_908,N_117);
nand U1948 (N_1948,N_1154,N_842);
nor U1949 (N_1949,N_962,N_483);
xor U1950 (N_1950,N_963,N_1285);
nand U1951 (N_1951,N_1454,N_1299);
nand U1952 (N_1952,N_589,N_769);
nor U1953 (N_1953,N_618,N_114);
nand U1954 (N_1954,N_15,N_1141);
xor U1955 (N_1955,N_364,N_690);
or U1956 (N_1956,N_20,N_360);
or U1957 (N_1957,N_1309,N_413);
nand U1958 (N_1958,N_571,N_1117);
and U1959 (N_1959,N_1028,N_455);
xnor U1960 (N_1960,N_145,N_477);
or U1961 (N_1961,N_350,N_75);
or U1962 (N_1962,N_995,N_19);
and U1963 (N_1963,N_885,N_1435);
nand U1964 (N_1964,N_189,N_1175);
and U1965 (N_1965,N_372,N_706);
and U1966 (N_1966,N_503,N_1105);
nand U1967 (N_1967,N_144,N_22);
nor U1968 (N_1968,N_151,N_1317);
nand U1969 (N_1969,N_785,N_1426);
or U1970 (N_1970,N_744,N_946);
nor U1971 (N_1971,N_362,N_550);
and U1972 (N_1972,N_697,N_278);
nor U1973 (N_1973,N_1267,N_242);
xnor U1974 (N_1974,N_1443,N_1430);
nand U1975 (N_1975,N_126,N_1142);
xor U1976 (N_1976,N_1157,N_351);
xor U1977 (N_1977,N_936,N_1219);
nand U1978 (N_1978,N_481,N_129);
nor U1979 (N_1979,N_601,N_1371);
nor U1980 (N_1980,N_353,N_82);
xnor U1981 (N_1981,N_245,N_205);
or U1982 (N_1982,N_956,N_1279);
xor U1983 (N_1983,N_234,N_1486);
nor U1984 (N_1984,N_153,N_110);
or U1985 (N_1985,N_464,N_330);
xor U1986 (N_1986,N_135,N_1412);
and U1987 (N_1987,N_836,N_103);
and U1988 (N_1988,N_101,N_256);
nor U1989 (N_1989,N_160,N_1223);
or U1990 (N_1990,N_374,N_315);
nand U1991 (N_1991,N_1161,N_1200);
xor U1992 (N_1992,N_361,N_1292);
or U1993 (N_1993,N_86,N_835);
and U1994 (N_1994,N_1149,N_528);
nor U1995 (N_1995,N_539,N_1491);
nor U1996 (N_1996,N_1330,N_1331);
xor U1997 (N_1997,N_90,N_1264);
xnor U1998 (N_1998,N_502,N_671);
or U1999 (N_1999,N_1258,N_556);
nand U2000 (N_2000,N_1040,N_1036);
and U2001 (N_2001,N_565,N_1228);
nor U2002 (N_2002,N_1445,N_333);
nand U2003 (N_2003,N_1039,N_705);
or U2004 (N_2004,N_368,N_524);
or U2005 (N_2005,N_1187,N_880);
xor U2006 (N_2006,N_322,N_41);
or U2007 (N_2007,N_378,N_887);
nor U2008 (N_2008,N_239,N_658);
or U2009 (N_2009,N_516,N_1186);
and U2010 (N_2010,N_1044,N_141);
and U2011 (N_2011,N_414,N_570);
nor U2012 (N_2012,N_1011,N_401);
xnor U2013 (N_2013,N_1492,N_274);
nor U2014 (N_2014,N_314,N_309);
or U2015 (N_2015,N_210,N_896);
or U2016 (N_2016,N_1198,N_1425);
and U2017 (N_2017,N_1170,N_1146);
and U2018 (N_2018,N_728,N_746);
and U2019 (N_2019,N_935,N_7);
nand U2020 (N_2020,N_852,N_818);
or U2021 (N_2021,N_637,N_1082);
xor U2022 (N_2022,N_857,N_1368);
nor U2023 (N_2023,N_1073,N_366);
nand U2024 (N_2024,N_434,N_1409);
nor U2025 (N_2025,N_901,N_660);
nand U2026 (N_2026,N_1271,N_1121);
nor U2027 (N_2027,N_858,N_1133);
nand U2028 (N_2028,N_537,N_1472);
nand U2029 (N_2029,N_1275,N_1190);
and U2030 (N_2030,N_1452,N_847);
nand U2031 (N_2031,N_758,N_196);
nand U2032 (N_2032,N_518,N_1123);
xor U2033 (N_2033,N_1364,N_1328);
nor U2034 (N_2034,N_616,N_1440);
and U2035 (N_2035,N_1116,N_961);
nand U2036 (N_2036,N_207,N_937);
or U2037 (N_2037,N_739,N_670);
nor U2038 (N_2038,N_1083,N_1119);
and U2039 (N_2039,N_520,N_1183);
nor U2040 (N_2040,N_606,N_1384);
and U2041 (N_2041,N_1152,N_496);
and U2042 (N_2042,N_1464,N_265);
or U2043 (N_2043,N_1363,N_1163);
or U2044 (N_2044,N_436,N_1193);
and U2045 (N_2045,N_18,N_131);
and U2046 (N_2046,N_608,N_1311);
nor U2047 (N_2047,N_814,N_1262);
nand U2048 (N_2048,N_779,N_1051);
xnor U2049 (N_2049,N_194,N_695);
and U2050 (N_2050,N_586,N_237);
or U2051 (N_2051,N_1207,N_137);
xor U2052 (N_2052,N_1041,N_124);
or U2053 (N_2053,N_1204,N_652);
or U2054 (N_2054,N_1249,N_1079);
xnor U2055 (N_2055,N_1098,N_251);
nor U2056 (N_2056,N_641,N_380);
xnor U2057 (N_2057,N_1293,N_1222);
xnor U2058 (N_2058,N_727,N_1372);
xnor U2059 (N_2059,N_850,N_442);
xor U2060 (N_2060,N_84,N_1458);
and U2061 (N_2061,N_791,N_692);
or U2062 (N_2062,N_854,N_1427);
and U2063 (N_2063,N_359,N_945);
and U2064 (N_2064,N_748,N_120);
or U2065 (N_2065,N_1038,N_1024);
nor U2066 (N_2066,N_447,N_1059);
nand U2067 (N_2067,N_303,N_254);
nand U2068 (N_2068,N_1365,N_394);
xor U2069 (N_2069,N_634,N_343);
and U2070 (N_2070,N_830,N_1469);
xnor U2071 (N_2071,N_456,N_793);
xor U2072 (N_2072,N_1245,N_215);
nor U2073 (N_2073,N_280,N_430);
nor U2074 (N_2074,N_166,N_367);
nand U2075 (N_2075,N_1298,N_666);
nor U2076 (N_2076,N_409,N_1143);
xor U2077 (N_2077,N_1095,N_416);
nand U2078 (N_2078,N_95,N_1495);
or U2079 (N_2079,N_1048,N_1471);
or U2080 (N_2080,N_1339,N_1307);
xor U2081 (N_2081,N_1386,N_175);
and U2082 (N_2082,N_1316,N_1209);
or U2083 (N_2083,N_667,N_560);
nor U2084 (N_2084,N_863,N_49);
nand U2085 (N_2085,N_848,N_294);
or U2086 (N_2086,N_400,N_327);
nor U2087 (N_2087,N_1210,N_906);
or U2088 (N_2088,N_804,N_986);
and U2089 (N_2089,N_184,N_907);
nor U2090 (N_2090,N_564,N_410);
nand U2091 (N_2091,N_281,N_532);
or U2092 (N_2092,N_143,N_489);
or U2093 (N_2093,N_498,N_62);
and U2094 (N_2094,N_1310,N_1014);
or U2095 (N_2095,N_633,N_932);
and U2096 (N_2096,N_206,N_693);
nor U2097 (N_2097,N_154,N_1318);
and U2098 (N_2098,N_580,N_1229);
or U2099 (N_2099,N_882,N_457);
nand U2100 (N_2100,N_845,N_195);
xor U2101 (N_2101,N_621,N_328);
nand U2102 (N_2102,N_840,N_1270);
xnor U2103 (N_2103,N_424,N_644);
nor U2104 (N_2104,N_182,N_628);
nor U2105 (N_2105,N_105,N_876);
nor U2106 (N_2106,N_283,N_1185);
or U2107 (N_2107,N_1255,N_1442);
and U2108 (N_2108,N_1189,N_1488);
and U2109 (N_2109,N_733,N_1194);
nand U2110 (N_2110,N_440,N_713);
nor U2111 (N_2111,N_1132,N_1);
xor U2112 (N_2112,N_778,N_1362);
nor U2113 (N_2113,N_451,N_285);
xnor U2114 (N_2114,N_155,N_417);
and U2115 (N_2115,N_878,N_1416);
nand U2116 (N_2116,N_356,N_716);
and U2117 (N_2117,N_301,N_159);
nand U2118 (N_2118,N_149,N_521);
nor U2119 (N_2119,N_1463,N_1124);
nor U2120 (N_2120,N_229,N_307);
and U2121 (N_2121,N_1431,N_718);
xor U2122 (N_2122,N_579,N_777);
xor U2123 (N_2123,N_861,N_349);
xor U2124 (N_2124,N_499,N_632);
xnor U2125 (N_2125,N_275,N_1215);
and U2126 (N_2126,N_905,N_1032);
nand U2127 (N_2127,N_797,N_960);
xor U2128 (N_2128,N_376,N_1150);
xnor U2129 (N_2129,N_551,N_107);
nand U2130 (N_2130,N_250,N_79);
nor U2131 (N_2131,N_1224,N_383);
xor U2132 (N_2132,N_1395,N_823);
and U2133 (N_2133,N_224,N_1294);
or U2134 (N_2134,N_298,N_313);
or U2135 (N_2135,N_1346,N_839);
xor U2136 (N_2136,N_382,N_998);
xnor U2137 (N_2137,N_77,N_574);
xnor U2138 (N_2138,N_429,N_1056);
or U2139 (N_2139,N_156,N_720);
nand U2140 (N_2140,N_1418,N_1390);
nand U2141 (N_2141,N_1456,N_252);
and U2142 (N_2142,N_299,N_891);
nand U2143 (N_2143,N_198,N_1313);
or U2144 (N_2144,N_1206,N_704);
and U2145 (N_2145,N_390,N_788);
and U2146 (N_2146,N_1239,N_1314);
nor U2147 (N_2147,N_646,N_1392);
xor U2148 (N_2148,N_741,N_187);
or U2149 (N_2149,N_74,N_888);
and U2150 (N_2150,N_1155,N_1383);
xnor U2151 (N_2151,N_783,N_292);
xnor U2152 (N_2152,N_1321,N_959);
or U2153 (N_2153,N_96,N_1496);
nand U2154 (N_2154,N_329,N_904);
xnor U2155 (N_2155,N_517,N_594);
or U2156 (N_2156,N_220,N_648);
and U2157 (N_2157,N_569,N_566);
or U2158 (N_2158,N_726,N_513);
nor U2159 (N_2159,N_411,N_1236);
nor U2160 (N_2160,N_820,N_943);
nand U2161 (N_2161,N_1379,N_202);
and U2162 (N_2162,N_1184,N_765);
and U2163 (N_2163,N_384,N_98);
nor U2164 (N_2164,N_786,N_1018);
or U2165 (N_2165,N_1074,N_711);
or U2166 (N_2166,N_5,N_515);
or U2167 (N_2167,N_80,N_833);
and U2168 (N_2168,N_91,N_352);
nor U2169 (N_2169,N_1192,N_70);
nor U2170 (N_2170,N_336,N_767);
xor U2171 (N_2171,N_920,N_216);
or U2172 (N_2172,N_1010,N_89);
or U2173 (N_2173,N_478,N_73);
or U2174 (N_2174,N_68,N_1201);
or U2175 (N_2175,N_1134,N_1344);
nor U2176 (N_2176,N_649,N_319);
or U2177 (N_2177,N_1240,N_1325);
nand U2178 (N_2178,N_1341,N_625);
or U2179 (N_2179,N_1460,N_339);
nand U2180 (N_2180,N_1063,N_627);
xnor U2181 (N_2181,N_675,N_1136);
and U2182 (N_2182,N_1058,N_1060);
or U2183 (N_2183,N_800,N_463);
nand U2184 (N_2184,N_700,N_59);
nand U2185 (N_2185,N_25,N_1398);
nor U2186 (N_2186,N_1075,N_302);
nor U2187 (N_2187,N_980,N_148);
xor U2188 (N_2188,N_680,N_801);
xor U2189 (N_2189,N_826,N_471);
xor U2190 (N_2190,N_1251,N_1122);
nor U2191 (N_2191,N_1145,N_655);
and U2192 (N_2192,N_1411,N_753);
nand U2193 (N_2193,N_58,N_749);
nand U2194 (N_2194,N_21,N_903);
or U2195 (N_2195,N_668,N_1099);
xor U2196 (N_2196,N_170,N_821);
or U2197 (N_2197,N_1388,N_1304);
nand U2198 (N_2198,N_645,N_796);
and U2199 (N_2199,N_674,N_415);
nand U2200 (N_2200,N_541,N_952);
and U2201 (N_2201,N_984,N_300);
nand U2202 (N_2202,N_391,N_1165);
nor U2203 (N_2203,N_1094,N_1457);
xnor U2204 (N_2204,N_923,N_862);
nand U2205 (N_2205,N_1459,N_982);
xor U2206 (N_2206,N_16,N_1168);
xnor U2207 (N_2207,N_1380,N_200);
or U2208 (N_2208,N_468,N_754);
nor U2209 (N_2209,N_1322,N_1438);
nor U2210 (N_2210,N_964,N_575);
xor U2211 (N_2211,N_1131,N_1061);
nand U2212 (N_2212,N_869,N_1473);
nor U2213 (N_2213,N_712,N_1283);
nand U2214 (N_2214,N_161,N_1139);
xor U2215 (N_2215,N_951,N_1076);
nand U2216 (N_2216,N_925,N_422);
and U2217 (N_2217,N_918,N_1172);
and U2218 (N_2218,N_576,N_425);
nand U2219 (N_2219,N_193,N_342);
or U2220 (N_2220,N_1033,N_1323);
or U2221 (N_2221,N_669,N_853);
or U2222 (N_2222,N_482,N_1233);
xor U2223 (N_2223,N_548,N_249);
or U2224 (N_2224,N_805,N_653);
xnor U2225 (N_2225,N_1104,N_1485);
xor U2226 (N_2226,N_312,N_631);
or U2227 (N_2227,N_1086,N_271);
and U2228 (N_2228,N_238,N_1399);
nor U2229 (N_2229,N_860,N_180);
xor U2230 (N_2230,N_106,N_428);
or U2231 (N_2231,N_990,N_1358);
or U2232 (N_2232,N_665,N_244);
nor U2233 (N_2233,N_140,N_1171);
and U2234 (N_2234,N_738,N_1280);
and U2235 (N_2235,N_1129,N_609);
nor U2236 (N_2236,N_774,N_1062);
nor U2237 (N_2237,N_1246,N_1400);
or U2238 (N_2238,N_30,N_1405);
or U2239 (N_2239,N_24,N_968);
and U2240 (N_2240,N_228,N_898);
nor U2241 (N_2241,N_1373,N_217);
xnor U2242 (N_2242,N_756,N_1269);
nand U2243 (N_2243,N_661,N_10);
nor U2244 (N_2244,N_827,N_530);
nor U2245 (N_2245,N_940,N_1065);
and U2246 (N_2246,N_1475,N_1305);
or U2247 (N_2247,N_1181,N_1025);
nor U2248 (N_2248,N_174,N_1047);
and U2249 (N_2249,N_1448,N_1030);
or U2250 (N_2250,N_110,N_179);
nor U2251 (N_2251,N_315,N_272);
nand U2252 (N_2252,N_1279,N_599);
xnor U2253 (N_2253,N_919,N_1106);
or U2254 (N_2254,N_98,N_667);
or U2255 (N_2255,N_1244,N_854);
and U2256 (N_2256,N_1217,N_194);
or U2257 (N_2257,N_140,N_1038);
and U2258 (N_2258,N_1337,N_1152);
xor U2259 (N_2259,N_940,N_226);
and U2260 (N_2260,N_1430,N_1279);
nor U2261 (N_2261,N_1219,N_240);
nand U2262 (N_2262,N_1456,N_597);
or U2263 (N_2263,N_11,N_469);
xor U2264 (N_2264,N_830,N_684);
or U2265 (N_2265,N_945,N_1087);
nor U2266 (N_2266,N_626,N_683);
nand U2267 (N_2267,N_1026,N_755);
nor U2268 (N_2268,N_141,N_1382);
nor U2269 (N_2269,N_433,N_320);
nand U2270 (N_2270,N_1029,N_531);
xor U2271 (N_2271,N_253,N_1388);
nor U2272 (N_2272,N_1346,N_68);
xnor U2273 (N_2273,N_449,N_926);
nand U2274 (N_2274,N_461,N_848);
xor U2275 (N_2275,N_780,N_1025);
and U2276 (N_2276,N_514,N_1440);
xor U2277 (N_2277,N_1403,N_489);
or U2278 (N_2278,N_744,N_536);
or U2279 (N_2279,N_1090,N_1169);
and U2280 (N_2280,N_794,N_1433);
nand U2281 (N_2281,N_1252,N_258);
and U2282 (N_2282,N_1288,N_952);
and U2283 (N_2283,N_764,N_254);
or U2284 (N_2284,N_464,N_990);
xnor U2285 (N_2285,N_1280,N_197);
nor U2286 (N_2286,N_683,N_844);
nor U2287 (N_2287,N_655,N_1027);
or U2288 (N_2288,N_1373,N_1333);
nor U2289 (N_2289,N_560,N_130);
and U2290 (N_2290,N_790,N_757);
xnor U2291 (N_2291,N_1099,N_990);
or U2292 (N_2292,N_334,N_969);
or U2293 (N_2293,N_371,N_258);
nand U2294 (N_2294,N_1282,N_324);
and U2295 (N_2295,N_308,N_1241);
xor U2296 (N_2296,N_240,N_1018);
or U2297 (N_2297,N_641,N_1209);
or U2298 (N_2298,N_517,N_39);
and U2299 (N_2299,N_770,N_413);
and U2300 (N_2300,N_1297,N_455);
xnor U2301 (N_2301,N_857,N_712);
and U2302 (N_2302,N_1430,N_1353);
xnor U2303 (N_2303,N_1403,N_45);
xor U2304 (N_2304,N_1424,N_1224);
xnor U2305 (N_2305,N_690,N_694);
xnor U2306 (N_2306,N_1228,N_561);
xnor U2307 (N_2307,N_749,N_1260);
nor U2308 (N_2308,N_233,N_792);
xnor U2309 (N_2309,N_849,N_27);
or U2310 (N_2310,N_1250,N_192);
xnor U2311 (N_2311,N_212,N_657);
nand U2312 (N_2312,N_1245,N_735);
nand U2313 (N_2313,N_1461,N_12);
nand U2314 (N_2314,N_1229,N_1249);
nor U2315 (N_2315,N_1259,N_874);
nand U2316 (N_2316,N_723,N_1302);
and U2317 (N_2317,N_557,N_843);
nor U2318 (N_2318,N_1307,N_196);
and U2319 (N_2319,N_765,N_889);
nand U2320 (N_2320,N_1205,N_1340);
and U2321 (N_2321,N_1488,N_723);
nor U2322 (N_2322,N_644,N_1221);
xor U2323 (N_2323,N_1169,N_1074);
nand U2324 (N_2324,N_664,N_207);
xor U2325 (N_2325,N_825,N_1245);
xor U2326 (N_2326,N_1362,N_666);
nor U2327 (N_2327,N_472,N_1419);
nor U2328 (N_2328,N_518,N_876);
xnor U2329 (N_2329,N_654,N_416);
or U2330 (N_2330,N_1492,N_276);
or U2331 (N_2331,N_408,N_1091);
xnor U2332 (N_2332,N_586,N_504);
nand U2333 (N_2333,N_812,N_430);
xnor U2334 (N_2334,N_178,N_405);
nor U2335 (N_2335,N_187,N_428);
nand U2336 (N_2336,N_846,N_1228);
nor U2337 (N_2337,N_2,N_249);
nor U2338 (N_2338,N_851,N_457);
or U2339 (N_2339,N_1176,N_272);
nand U2340 (N_2340,N_701,N_684);
xor U2341 (N_2341,N_256,N_1338);
or U2342 (N_2342,N_831,N_763);
or U2343 (N_2343,N_1432,N_1212);
nand U2344 (N_2344,N_105,N_505);
nor U2345 (N_2345,N_296,N_1228);
nor U2346 (N_2346,N_1363,N_615);
xor U2347 (N_2347,N_466,N_339);
nor U2348 (N_2348,N_641,N_1378);
and U2349 (N_2349,N_273,N_672);
nand U2350 (N_2350,N_1431,N_213);
and U2351 (N_2351,N_576,N_152);
xor U2352 (N_2352,N_1496,N_330);
and U2353 (N_2353,N_243,N_145);
and U2354 (N_2354,N_1478,N_1219);
xnor U2355 (N_2355,N_817,N_1121);
and U2356 (N_2356,N_1000,N_194);
xor U2357 (N_2357,N_871,N_175);
nor U2358 (N_2358,N_1367,N_1461);
xnor U2359 (N_2359,N_63,N_902);
xnor U2360 (N_2360,N_500,N_989);
or U2361 (N_2361,N_331,N_903);
xor U2362 (N_2362,N_812,N_120);
xnor U2363 (N_2363,N_143,N_755);
or U2364 (N_2364,N_1450,N_83);
nand U2365 (N_2365,N_1266,N_171);
nor U2366 (N_2366,N_1248,N_1346);
and U2367 (N_2367,N_1093,N_589);
xor U2368 (N_2368,N_772,N_578);
or U2369 (N_2369,N_926,N_1278);
nand U2370 (N_2370,N_763,N_219);
or U2371 (N_2371,N_963,N_1459);
nand U2372 (N_2372,N_1411,N_700);
or U2373 (N_2373,N_1147,N_390);
nor U2374 (N_2374,N_555,N_650);
nor U2375 (N_2375,N_872,N_183);
or U2376 (N_2376,N_702,N_1018);
nor U2377 (N_2377,N_1438,N_810);
nor U2378 (N_2378,N_79,N_1094);
or U2379 (N_2379,N_46,N_658);
nand U2380 (N_2380,N_953,N_793);
xnor U2381 (N_2381,N_341,N_539);
nor U2382 (N_2382,N_743,N_555);
xnor U2383 (N_2383,N_1482,N_1244);
xor U2384 (N_2384,N_1111,N_1337);
or U2385 (N_2385,N_1104,N_1451);
nand U2386 (N_2386,N_812,N_1423);
xnor U2387 (N_2387,N_796,N_1083);
nand U2388 (N_2388,N_12,N_10);
or U2389 (N_2389,N_695,N_816);
xnor U2390 (N_2390,N_384,N_78);
nor U2391 (N_2391,N_465,N_105);
nor U2392 (N_2392,N_1400,N_667);
nand U2393 (N_2393,N_1457,N_1087);
nor U2394 (N_2394,N_555,N_246);
nand U2395 (N_2395,N_793,N_563);
or U2396 (N_2396,N_1471,N_1163);
xnor U2397 (N_2397,N_1245,N_1194);
and U2398 (N_2398,N_692,N_758);
or U2399 (N_2399,N_405,N_1173);
and U2400 (N_2400,N_1382,N_507);
nand U2401 (N_2401,N_751,N_941);
nor U2402 (N_2402,N_1402,N_321);
and U2403 (N_2403,N_183,N_179);
nor U2404 (N_2404,N_649,N_834);
xor U2405 (N_2405,N_436,N_228);
nand U2406 (N_2406,N_29,N_750);
and U2407 (N_2407,N_1206,N_89);
and U2408 (N_2408,N_357,N_104);
xnor U2409 (N_2409,N_1093,N_607);
and U2410 (N_2410,N_840,N_925);
nand U2411 (N_2411,N_682,N_936);
xnor U2412 (N_2412,N_407,N_1488);
nor U2413 (N_2413,N_927,N_1446);
nor U2414 (N_2414,N_610,N_176);
xor U2415 (N_2415,N_57,N_433);
xor U2416 (N_2416,N_617,N_803);
nor U2417 (N_2417,N_629,N_710);
or U2418 (N_2418,N_976,N_1273);
and U2419 (N_2419,N_1437,N_503);
nand U2420 (N_2420,N_989,N_136);
nor U2421 (N_2421,N_51,N_808);
xnor U2422 (N_2422,N_1080,N_949);
xnor U2423 (N_2423,N_1394,N_306);
and U2424 (N_2424,N_86,N_6);
and U2425 (N_2425,N_32,N_998);
xnor U2426 (N_2426,N_1211,N_70);
xnor U2427 (N_2427,N_107,N_1280);
nand U2428 (N_2428,N_205,N_1289);
nor U2429 (N_2429,N_1448,N_272);
xor U2430 (N_2430,N_1232,N_604);
and U2431 (N_2431,N_281,N_933);
and U2432 (N_2432,N_172,N_1113);
nand U2433 (N_2433,N_401,N_419);
nand U2434 (N_2434,N_1211,N_158);
nand U2435 (N_2435,N_1019,N_1064);
and U2436 (N_2436,N_352,N_261);
and U2437 (N_2437,N_756,N_23);
nand U2438 (N_2438,N_962,N_1298);
and U2439 (N_2439,N_603,N_1077);
xnor U2440 (N_2440,N_999,N_953);
nor U2441 (N_2441,N_967,N_1374);
nor U2442 (N_2442,N_1495,N_374);
or U2443 (N_2443,N_730,N_307);
xor U2444 (N_2444,N_1471,N_73);
nand U2445 (N_2445,N_1130,N_646);
or U2446 (N_2446,N_402,N_932);
xnor U2447 (N_2447,N_260,N_65);
nor U2448 (N_2448,N_1398,N_214);
xor U2449 (N_2449,N_984,N_969);
nand U2450 (N_2450,N_120,N_636);
nand U2451 (N_2451,N_1178,N_229);
or U2452 (N_2452,N_1391,N_72);
nor U2453 (N_2453,N_1472,N_726);
nor U2454 (N_2454,N_1297,N_81);
nand U2455 (N_2455,N_10,N_271);
or U2456 (N_2456,N_1484,N_1178);
nor U2457 (N_2457,N_904,N_1024);
nor U2458 (N_2458,N_624,N_215);
xor U2459 (N_2459,N_1233,N_1009);
xnor U2460 (N_2460,N_832,N_814);
or U2461 (N_2461,N_806,N_499);
xnor U2462 (N_2462,N_465,N_594);
and U2463 (N_2463,N_1028,N_678);
or U2464 (N_2464,N_392,N_444);
and U2465 (N_2465,N_716,N_1236);
xor U2466 (N_2466,N_1079,N_730);
xor U2467 (N_2467,N_1099,N_1105);
and U2468 (N_2468,N_564,N_1131);
or U2469 (N_2469,N_47,N_1240);
nand U2470 (N_2470,N_757,N_896);
and U2471 (N_2471,N_232,N_490);
xor U2472 (N_2472,N_843,N_1022);
or U2473 (N_2473,N_1170,N_1449);
nor U2474 (N_2474,N_542,N_633);
xnor U2475 (N_2475,N_277,N_177);
nand U2476 (N_2476,N_16,N_30);
xnor U2477 (N_2477,N_377,N_1341);
nand U2478 (N_2478,N_1051,N_1282);
xnor U2479 (N_2479,N_409,N_936);
nand U2480 (N_2480,N_1258,N_1456);
nor U2481 (N_2481,N_183,N_677);
and U2482 (N_2482,N_812,N_705);
and U2483 (N_2483,N_74,N_1435);
nor U2484 (N_2484,N_405,N_708);
nor U2485 (N_2485,N_12,N_497);
or U2486 (N_2486,N_1247,N_335);
and U2487 (N_2487,N_850,N_1435);
and U2488 (N_2488,N_746,N_1018);
and U2489 (N_2489,N_1262,N_616);
xor U2490 (N_2490,N_1173,N_176);
nand U2491 (N_2491,N_83,N_780);
xor U2492 (N_2492,N_26,N_952);
nor U2493 (N_2493,N_980,N_644);
nand U2494 (N_2494,N_89,N_1275);
and U2495 (N_2495,N_68,N_451);
nand U2496 (N_2496,N_965,N_134);
or U2497 (N_2497,N_74,N_10);
xor U2498 (N_2498,N_142,N_907);
and U2499 (N_2499,N_890,N_108);
or U2500 (N_2500,N_1079,N_1172);
or U2501 (N_2501,N_1267,N_277);
and U2502 (N_2502,N_772,N_1148);
and U2503 (N_2503,N_427,N_846);
nor U2504 (N_2504,N_970,N_868);
nand U2505 (N_2505,N_1214,N_1115);
nor U2506 (N_2506,N_379,N_1070);
nor U2507 (N_2507,N_411,N_172);
or U2508 (N_2508,N_1068,N_596);
nand U2509 (N_2509,N_982,N_1484);
or U2510 (N_2510,N_1011,N_289);
and U2511 (N_2511,N_1308,N_843);
nor U2512 (N_2512,N_1392,N_496);
nor U2513 (N_2513,N_266,N_1100);
xor U2514 (N_2514,N_894,N_420);
xnor U2515 (N_2515,N_282,N_1386);
nand U2516 (N_2516,N_881,N_953);
xor U2517 (N_2517,N_559,N_1320);
or U2518 (N_2518,N_394,N_841);
nor U2519 (N_2519,N_365,N_529);
and U2520 (N_2520,N_667,N_368);
nand U2521 (N_2521,N_1023,N_94);
xnor U2522 (N_2522,N_751,N_1193);
xor U2523 (N_2523,N_752,N_652);
nand U2524 (N_2524,N_930,N_1054);
nor U2525 (N_2525,N_559,N_13);
nand U2526 (N_2526,N_361,N_561);
xor U2527 (N_2527,N_555,N_1159);
and U2528 (N_2528,N_251,N_20);
or U2529 (N_2529,N_287,N_484);
xnor U2530 (N_2530,N_440,N_445);
nor U2531 (N_2531,N_214,N_908);
and U2532 (N_2532,N_937,N_251);
or U2533 (N_2533,N_274,N_1376);
nor U2534 (N_2534,N_1445,N_694);
and U2535 (N_2535,N_71,N_235);
xnor U2536 (N_2536,N_811,N_1147);
xnor U2537 (N_2537,N_1376,N_748);
and U2538 (N_2538,N_769,N_551);
xnor U2539 (N_2539,N_609,N_1331);
or U2540 (N_2540,N_814,N_596);
nand U2541 (N_2541,N_100,N_1310);
and U2542 (N_2542,N_744,N_143);
and U2543 (N_2543,N_809,N_1090);
nor U2544 (N_2544,N_999,N_1492);
xnor U2545 (N_2545,N_333,N_716);
and U2546 (N_2546,N_783,N_1175);
nor U2547 (N_2547,N_1330,N_230);
nand U2548 (N_2548,N_1202,N_43);
xor U2549 (N_2549,N_603,N_443);
or U2550 (N_2550,N_180,N_133);
xor U2551 (N_2551,N_12,N_360);
xor U2552 (N_2552,N_804,N_1216);
or U2553 (N_2553,N_116,N_71);
or U2554 (N_2554,N_213,N_1408);
nor U2555 (N_2555,N_725,N_581);
and U2556 (N_2556,N_713,N_262);
xnor U2557 (N_2557,N_1310,N_1478);
xnor U2558 (N_2558,N_559,N_1000);
nand U2559 (N_2559,N_1451,N_1070);
xor U2560 (N_2560,N_1159,N_1404);
xnor U2561 (N_2561,N_804,N_39);
nand U2562 (N_2562,N_788,N_1050);
nor U2563 (N_2563,N_1317,N_156);
or U2564 (N_2564,N_1126,N_436);
nor U2565 (N_2565,N_798,N_1469);
nand U2566 (N_2566,N_878,N_784);
nand U2567 (N_2567,N_526,N_334);
or U2568 (N_2568,N_159,N_669);
xnor U2569 (N_2569,N_1406,N_294);
nand U2570 (N_2570,N_1361,N_670);
xnor U2571 (N_2571,N_767,N_1334);
xnor U2572 (N_2572,N_1399,N_1148);
nand U2573 (N_2573,N_543,N_1452);
nor U2574 (N_2574,N_1293,N_1448);
nor U2575 (N_2575,N_313,N_769);
xor U2576 (N_2576,N_671,N_62);
xor U2577 (N_2577,N_1186,N_1428);
nand U2578 (N_2578,N_959,N_944);
or U2579 (N_2579,N_830,N_1147);
or U2580 (N_2580,N_987,N_548);
and U2581 (N_2581,N_1484,N_707);
and U2582 (N_2582,N_1006,N_505);
xor U2583 (N_2583,N_401,N_998);
nand U2584 (N_2584,N_1205,N_1308);
nor U2585 (N_2585,N_1461,N_1353);
xnor U2586 (N_2586,N_696,N_1122);
and U2587 (N_2587,N_1365,N_1279);
nand U2588 (N_2588,N_854,N_1173);
nor U2589 (N_2589,N_1488,N_437);
nand U2590 (N_2590,N_452,N_889);
xnor U2591 (N_2591,N_973,N_1200);
or U2592 (N_2592,N_86,N_294);
and U2593 (N_2593,N_212,N_588);
xor U2594 (N_2594,N_824,N_1391);
xor U2595 (N_2595,N_28,N_970);
xor U2596 (N_2596,N_1037,N_634);
nand U2597 (N_2597,N_706,N_1230);
and U2598 (N_2598,N_1012,N_1286);
nor U2599 (N_2599,N_1256,N_247);
nand U2600 (N_2600,N_472,N_1308);
nand U2601 (N_2601,N_698,N_209);
xor U2602 (N_2602,N_1313,N_88);
xor U2603 (N_2603,N_399,N_1225);
nor U2604 (N_2604,N_238,N_118);
or U2605 (N_2605,N_261,N_952);
or U2606 (N_2606,N_212,N_25);
and U2607 (N_2607,N_1361,N_920);
nor U2608 (N_2608,N_554,N_440);
or U2609 (N_2609,N_835,N_684);
nand U2610 (N_2610,N_709,N_94);
or U2611 (N_2611,N_36,N_811);
nor U2612 (N_2612,N_1370,N_695);
and U2613 (N_2613,N_1477,N_481);
or U2614 (N_2614,N_525,N_429);
or U2615 (N_2615,N_859,N_1487);
nand U2616 (N_2616,N_20,N_741);
nand U2617 (N_2617,N_1326,N_501);
nor U2618 (N_2618,N_1338,N_602);
and U2619 (N_2619,N_896,N_553);
or U2620 (N_2620,N_355,N_1058);
xnor U2621 (N_2621,N_990,N_69);
nand U2622 (N_2622,N_1275,N_1311);
nand U2623 (N_2623,N_91,N_1088);
nand U2624 (N_2624,N_256,N_677);
nand U2625 (N_2625,N_467,N_657);
nor U2626 (N_2626,N_1041,N_645);
xor U2627 (N_2627,N_1441,N_154);
nor U2628 (N_2628,N_154,N_311);
or U2629 (N_2629,N_873,N_116);
and U2630 (N_2630,N_571,N_546);
or U2631 (N_2631,N_1401,N_1346);
and U2632 (N_2632,N_1176,N_811);
xor U2633 (N_2633,N_933,N_1296);
and U2634 (N_2634,N_365,N_959);
nand U2635 (N_2635,N_192,N_1065);
and U2636 (N_2636,N_40,N_1431);
xnor U2637 (N_2637,N_955,N_617);
or U2638 (N_2638,N_154,N_762);
or U2639 (N_2639,N_77,N_443);
nand U2640 (N_2640,N_68,N_491);
xnor U2641 (N_2641,N_1222,N_1378);
nand U2642 (N_2642,N_1182,N_1040);
or U2643 (N_2643,N_954,N_1115);
nand U2644 (N_2644,N_275,N_1274);
nand U2645 (N_2645,N_399,N_479);
nor U2646 (N_2646,N_413,N_662);
nand U2647 (N_2647,N_1232,N_629);
or U2648 (N_2648,N_1394,N_355);
nand U2649 (N_2649,N_617,N_1420);
and U2650 (N_2650,N_1106,N_932);
or U2651 (N_2651,N_1073,N_452);
and U2652 (N_2652,N_1491,N_1082);
and U2653 (N_2653,N_1272,N_1322);
nand U2654 (N_2654,N_1199,N_999);
xnor U2655 (N_2655,N_1015,N_812);
nand U2656 (N_2656,N_146,N_403);
nand U2657 (N_2657,N_1425,N_898);
and U2658 (N_2658,N_532,N_536);
nand U2659 (N_2659,N_246,N_751);
nor U2660 (N_2660,N_600,N_373);
nor U2661 (N_2661,N_706,N_789);
and U2662 (N_2662,N_1313,N_273);
and U2663 (N_2663,N_1393,N_1351);
nor U2664 (N_2664,N_1375,N_499);
xor U2665 (N_2665,N_999,N_563);
or U2666 (N_2666,N_368,N_1198);
or U2667 (N_2667,N_1469,N_57);
or U2668 (N_2668,N_376,N_759);
and U2669 (N_2669,N_512,N_830);
or U2670 (N_2670,N_1441,N_1438);
xor U2671 (N_2671,N_1047,N_530);
nor U2672 (N_2672,N_528,N_418);
and U2673 (N_2673,N_184,N_947);
and U2674 (N_2674,N_50,N_834);
nand U2675 (N_2675,N_126,N_815);
nor U2676 (N_2676,N_1186,N_665);
or U2677 (N_2677,N_625,N_889);
or U2678 (N_2678,N_1091,N_1099);
or U2679 (N_2679,N_822,N_1408);
or U2680 (N_2680,N_1112,N_1213);
xnor U2681 (N_2681,N_85,N_31);
and U2682 (N_2682,N_779,N_1451);
nor U2683 (N_2683,N_829,N_115);
or U2684 (N_2684,N_718,N_262);
xor U2685 (N_2685,N_335,N_1033);
xor U2686 (N_2686,N_1191,N_689);
and U2687 (N_2687,N_1081,N_918);
and U2688 (N_2688,N_1141,N_1354);
and U2689 (N_2689,N_123,N_602);
nor U2690 (N_2690,N_654,N_403);
xnor U2691 (N_2691,N_526,N_793);
xnor U2692 (N_2692,N_245,N_982);
nand U2693 (N_2693,N_1370,N_903);
xor U2694 (N_2694,N_986,N_547);
nor U2695 (N_2695,N_104,N_753);
nand U2696 (N_2696,N_1048,N_464);
nand U2697 (N_2697,N_1047,N_935);
xor U2698 (N_2698,N_164,N_69);
nor U2699 (N_2699,N_868,N_103);
xor U2700 (N_2700,N_1052,N_306);
nor U2701 (N_2701,N_1322,N_96);
nand U2702 (N_2702,N_1421,N_437);
or U2703 (N_2703,N_237,N_1239);
nand U2704 (N_2704,N_1403,N_592);
nand U2705 (N_2705,N_819,N_294);
or U2706 (N_2706,N_86,N_1402);
xnor U2707 (N_2707,N_984,N_715);
nand U2708 (N_2708,N_1426,N_382);
xor U2709 (N_2709,N_477,N_494);
or U2710 (N_2710,N_490,N_1005);
xor U2711 (N_2711,N_587,N_1310);
xnor U2712 (N_2712,N_61,N_240);
nor U2713 (N_2713,N_1441,N_1313);
or U2714 (N_2714,N_880,N_551);
or U2715 (N_2715,N_781,N_1172);
or U2716 (N_2716,N_212,N_274);
and U2717 (N_2717,N_1038,N_1476);
nor U2718 (N_2718,N_1248,N_412);
nand U2719 (N_2719,N_1418,N_206);
and U2720 (N_2720,N_1134,N_801);
nand U2721 (N_2721,N_96,N_645);
or U2722 (N_2722,N_1254,N_993);
nor U2723 (N_2723,N_217,N_794);
and U2724 (N_2724,N_1064,N_273);
nand U2725 (N_2725,N_358,N_988);
nand U2726 (N_2726,N_1031,N_103);
and U2727 (N_2727,N_180,N_276);
or U2728 (N_2728,N_679,N_186);
xnor U2729 (N_2729,N_115,N_186);
and U2730 (N_2730,N_366,N_981);
nor U2731 (N_2731,N_1225,N_159);
nand U2732 (N_2732,N_92,N_812);
nor U2733 (N_2733,N_226,N_97);
nand U2734 (N_2734,N_769,N_217);
and U2735 (N_2735,N_1030,N_226);
or U2736 (N_2736,N_304,N_1141);
xor U2737 (N_2737,N_895,N_421);
and U2738 (N_2738,N_50,N_836);
xor U2739 (N_2739,N_477,N_359);
and U2740 (N_2740,N_1399,N_1035);
or U2741 (N_2741,N_857,N_1017);
xor U2742 (N_2742,N_961,N_1013);
or U2743 (N_2743,N_731,N_1177);
or U2744 (N_2744,N_1359,N_656);
nor U2745 (N_2745,N_178,N_511);
xor U2746 (N_2746,N_1231,N_1437);
nor U2747 (N_2747,N_1353,N_1141);
xor U2748 (N_2748,N_1362,N_234);
xor U2749 (N_2749,N_463,N_165);
nor U2750 (N_2750,N_1067,N_145);
and U2751 (N_2751,N_295,N_982);
nor U2752 (N_2752,N_201,N_821);
xor U2753 (N_2753,N_1098,N_1125);
xor U2754 (N_2754,N_409,N_539);
or U2755 (N_2755,N_420,N_1351);
nand U2756 (N_2756,N_609,N_140);
or U2757 (N_2757,N_943,N_972);
xnor U2758 (N_2758,N_1380,N_229);
or U2759 (N_2759,N_558,N_1460);
nand U2760 (N_2760,N_1214,N_250);
or U2761 (N_2761,N_276,N_147);
and U2762 (N_2762,N_688,N_1097);
or U2763 (N_2763,N_963,N_62);
xor U2764 (N_2764,N_474,N_1487);
and U2765 (N_2765,N_535,N_30);
xnor U2766 (N_2766,N_872,N_550);
nor U2767 (N_2767,N_1172,N_757);
and U2768 (N_2768,N_601,N_827);
nor U2769 (N_2769,N_123,N_262);
or U2770 (N_2770,N_1487,N_1027);
and U2771 (N_2771,N_608,N_1111);
xor U2772 (N_2772,N_532,N_106);
nand U2773 (N_2773,N_954,N_96);
or U2774 (N_2774,N_845,N_749);
nor U2775 (N_2775,N_731,N_194);
xnor U2776 (N_2776,N_727,N_944);
nor U2777 (N_2777,N_569,N_210);
xnor U2778 (N_2778,N_1065,N_1116);
or U2779 (N_2779,N_1018,N_1185);
nor U2780 (N_2780,N_541,N_1164);
nor U2781 (N_2781,N_962,N_324);
nor U2782 (N_2782,N_202,N_1154);
and U2783 (N_2783,N_1432,N_102);
and U2784 (N_2784,N_896,N_347);
or U2785 (N_2785,N_1241,N_476);
or U2786 (N_2786,N_1440,N_443);
nor U2787 (N_2787,N_1120,N_761);
nand U2788 (N_2788,N_147,N_563);
nor U2789 (N_2789,N_1490,N_371);
nor U2790 (N_2790,N_1330,N_1221);
nand U2791 (N_2791,N_1270,N_315);
xor U2792 (N_2792,N_1429,N_1234);
xnor U2793 (N_2793,N_995,N_957);
nand U2794 (N_2794,N_800,N_896);
nand U2795 (N_2795,N_482,N_731);
xor U2796 (N_2796,N_369,N_539);
nand U2797 (N_2797,N_610,N_770);
and U2798 (N_2798,N_517,N_944);
or U2799 (N_2799,N_223,N_1133);
nand U2800 (N_2800,N_830,N_880);
nand U2801 (N_2801,N_426,N_125);
and U2802 (N_2802,N_517,N_668);
nor U2803 (N_2803,N_1010,N_418);
xor U2804 (N_2804,N_22,N_1393);
nor U2805 (N_2805,N_224,N_123);
nor U2806 (N_2806,N_701,N_298);
or U2807 (N_2807,N_828,N_303);
and U2808 (N_2808,N_735,N_475);
xor U2809 (N_2809,N_145,N_15);
or U2810 (N_2810,N_235,N_1016);
xor U2811 (N_2811,N_749,N_84);
nand U2812 (N_2812,N_687,N_200);
and U2813 (N_2813,N_518,N_986);
and U2814 (N_2814,N_1241,N_1325);
or U2815 (N_2815,N_458,N_711);
nand U2816 (N_2816,N_32,N_244);
xor U2817 (N_2817,N_846,N_527);
and U2818 (N_2818,N_825,N_1225);
and U2819 (N_2819,N_2,N_782);
and U2820 (N_2820,N_549,N_398);
nand U2821 (N_2821,N_959,N_1137);
nand U2822 (N_2822,N_1174,N_593);
nand U2823 (N_2823,N_276,N_762);
and U2824 (N_2824,N_1028,N_294);
and U2825 (N_2825,N_1476,N_1336);
xnor U2826 (N_2826,N_719,N_940);
nor U2827 (N_2827,N_789,N_365);
or U2828 (N_2828,N_1152,N_501);
nor U2829 (N_2829,N_996,N_1368);
nor U2830 (N_2830,N_248,N_417);
or U2831 (N_2831,N_1053,N_1284);
nor U2832 (N_2832,N_1433,N_775);
or U2833 (N_2833,N_687,N_692);
or U2834 (N_2834,N_1035,N_1431);
nor U2835 (N_2835,N_688,N_1421);
and U2836 (N_2836,N_88,N_1470);
xnor U2837 (N_2837,N_701,N_1448);
or U2838 (N_2838,N_1093,N_1144);
xor U2839 (N_2839,N_1498,N_1140);
nor U2840 (N_2840,N_353,N_932);
nor U2841 (N_2841,N_156,N_871);
nor U2842 (N_2842,N_156,N_565);
or U2843 (N_2843,N_1300,N_718);
nor U2844 (N_2844,N_207,N_495);
nand U2845 (N_2845,N_984,N_283);
nand U2846 (N_2846,N_1325,N_1379);
or U2847 (N_2847,N_233,N_631);
or U2848 (N_2848,N_533,N_1347);
or U2849 (N_2849,N_716,N_1460);
nor U2850 (N_2850,N_49,N_650);
xnor U2851 (N_2851,N_1035,N_870);
xor U2852 (N_2852,N_1099,N_264);
and U2853 (N_2853,N_810,N_896);
nand U2854 (N_2854,N_343,N_763);
nor U2855 (N_2855,N_527,N_121);
nor U2856 (N_2856,N_667,N_251);
nand U2857 (N_2857,N_776,N_1100);
nor U2858 (N_2858,N_1164,N_464);
and U2859 (N_2859,N_1362,N_1058);
nand U2860 (N_2860,N_1077,N_361);
nand U2861 (N_2861,N_221,N_1011);
nor U2862 (N_2862,N_172,N_676);
xor U2863 (N_2863,N_1214,N_221);
nand U2864 (N_2864,N_832,N_1360);
and U2865 (N_2865,N_169,N_900);
nor U2866 (N_2866,N_875,N_1441);
nor U2867 (N_2867,N_996,N_1464);
nor U2868 (N_2868,N_343,N_508);
and U2869 (N_2869,N_998,N_1004);
xnor U2870 (N_2870,N_198,N_185);
or U2871 (N_2871,N_577,N_114);
xor U2872 (N_2872,N_1231,N_534);
or U2873 (N_2873,N_493,N_785);
and U2874 (N_2874,N_1055,N_705);
nand U2875 (N_2875,N_1396,N_1235);
or U2876 (N_2876,N_726,N_1120);
xor U2877 (N_2877,N_971,N_729);
nor U2878 (N_2878,N_228,N_186);
and U2879 (N_2879,N_94,N_819);
and U2880 (N_2880,N_286,N_361);
xnor U2881 (N_2881,N_731,N_4);
or U2882 (N_2882,N_98,N_605);
nor U2883 (N_2883,N_743,N_1235);
and U2884 (N_2884,N_1271,N_507);
nor U2885 (N_2885,N_625,N_301);
xnor U2886 (N_2886,N_132,N_397);
and U2887 (N_2887,N_936,N_1332);
xnor U2888 (N_2888,N_1276,N_1168);
and U2889 (N_2889,N_709,N_1352);
xnor U2890 (N_2890,N_1104,N_979);
and U2891 (N_2891,N_976,N_688);
nor U2892 (N_2892,N_451,N_282);
nor U2893 (N_2893,N_742,N_823);
or U2894 (N_2894,N_242,N_533);
xnor U2895 (N_2895,N_882,N_1434);
and U2896 (N_2896,N_972,N_175);
xnor U2897 (N_2897,N_258,N_1181);
or U2898 (N_2898,N_1136,N_868);
nor U2899 (N_2899,N_1401,N_923);
nor U2900 (N_2900,N_1136,N_90);
nor U2901 (N_2901,N_1064,N_1243);
nand U2902 (N_2902,N_542,N_380);
nor U2903 (N_2903,N_1050,N_659);
nand U2904 (N_2904,N_359,N_1179);
or U2905 (N_2905,N_518,N_96);
and U2906 (N_2906,N_26,N_486);
and U2907 (N_2907,N_1055,N_1498);
and U2908 (N_2908,N_606,N_904);
nor U2909 (N_2909,N_295,N_194);
or U2910 (N_2910,N_1156,N_808);
nand U2911 (N_2911,N_1141,N_71);
nand U2912 (N_2912,N_1457,N_110);
xnor U2913 (N_2913,N_1285,N_370);
nand U2914 (N_2914,N_536,N_1318);
xnor U2915 (N_2915,N_1074,N_933);
and U2916 (N_2916,N_615,N_43);
nor U2917 (N_2917,N_603,N_740);
nand U2918 (N_2918,N_194,N_636);
and U2919 (N_2919,N_1201,N_1250);
nand U2920 (N_2920,N_1251,N_823);
nor U2921 (N_2921,N_1118,N_1388);
nor U2922 (N_2922,N_534,N_108);
or U2923 (N_2923,N_89,N_1491);
or U2924 (N_2924,N_73,N_1385);
xor U2925 (N_2925,N_1395,N_879);
or U2926 (N_2926,N_310,N_970);
and U2927 (N_2927,N_551,N_1255);
or U2928 (N_2928,N_1202,N_742);
and U2929 (N_2929,N_402,N_1253);
xnor U2930 (N_2930,N_1134,N_202);
or U2931 (N_2931,N_1066,N_427);
nand U2932 (N_2932,N_640,N_140);
or U2933 (N_2933,N_1377,N_1213);
or U2934 (N_2934,N_1474,N_383);
or U2935 (N_2935,N_1011,N_135);
and U2936 (N_2936,N_754,N_1162);
and U2937 (N_2937,N_810,N_216);
or U2938 (N_2938,N_1249,N_264);
nor U2939 (N_2939,N_586,N_882);
nand U2940 (N_2940,N_1397,N_1479);
nand U2941 (N_2941,N_36,N_172);
nor U2942 (N_2942,N_1272,N_1493);
and U2943 (N_2943,N_487,N_427);
nand U2944 (N_2944,N_87,N_574);
nor U2945 (N_2945,N_348,N_332);
xor U2946 (N_2946,N_30,N_1386);
and U2947 (N_2947,N_413,N_970);
nor U2948 (N_2948,N_337,N_465);
nand U2949 (N_2949,N_1032,N_1378);
nor U2950 (N_2950,N_108,N_1321);
nor U2951 (N_2951,N_459,N_980);
nand U2952 (N_2952,N_131,N_543);
xor U2953 (N_2953,N_1342,N_233);
nand U2954 (N_2954,N_242,N_117);
xnor U2955 (N_2955,N_666,N_527);
and U2956 (N_2956,N_1045,N_833);
nor U2957 (N_2957,N_1291,N_1151);
or U2958 (N_2958,N_996,N_256);
and U2959 (N_2959,N_1413,N_676);
or U2960 (N_2960,N_774,N_1058);
and U2961 (N_2961,N_1330,N_435);
and U2962 (N_2962,N_1382,N_703);
and U2963 (N_2963,N_1119,N_911);
nand U2964 (N_2964,N_5,N_596);
or U2965 (N_2965,N_1018,N_434);
nand U2966 (N_2966,N_340,N_1170);
nand U2967 (N_2967,N_1372,N_1087);
nand U2968 (N_2968,N_838,N_1156);
nand U2969 (N_2969,N_1124,N_166);
nor U2970 (N_2970,N_652,N_1045);
xnor U2971 (N_2971,N_151,N_96);
and U2972 (N_2972,N_1011,N_396);
nor U2973 (N_2973,N_60,N_331);
xnor U2974 (N_2974,N_511,N_633);
nand U2975 (N_2975,N_399,N_536);
nor U2976 (N_2976,N_419,N_739);
and U2977 (N_2977,N_528,N_359);
nor U2978 (N_2978,N_1124,N_786);
xnor U2979 (N_2979,N_432,N_1175);
xnor U2980 (N_2980,N_998,N_653);
xor U2981 (N_2981,N_1354,N_90);
xor U2982 (N_2982,N_1197,N_1411);
or U2983 (N_2983,N_1305,N_1261);
nor U2984 (N_2984,N_1305,N_1126);
nor U2985 (N_2985,N_217,N_613);
nor U2986 (N_2986,N_1494,N_576);
or U2987 (N_2987,N_1388,N_593);
xnor U2988 (N_2988,N_158,N_1408);
xnor U2989 (N_2989,N_95,N_784);
nand U2990 (N_2990,N_1485,N_1183);
or U2991 (N_2991,N_1190,N_595);
or U2992 (N_2992,N_352,N_903);
or U2993 (N_2993,N_35,N_56);
or U2994 (N_2994,N_1070,N_79);
and U2995 (N_2995,N_282,N_36);
and U2996 (N_2996,N_1074,N_1353);
nor U2997 (N_2997,N_769,N_1342);
nand U2998 (N_2998,N_251,N_888);
nand U2999 (N_2999,N_291,N_335);
nand U3000 (N_3000,N_2076,N_2777);
or U3001 (N_3001,N_2106,N_1584);
xor U3002 (N_3002,N_2561,N_2428);
nand U3003 (N_3003,N_2673,N_1540);
or U3004 (N_3004,N_2402,N_2795);
nand U3005 (N_3005,N_1795,N_2017);
nor U3006 (N_3006,N_2277,N_2022);
nor U3007 (N_3007,N_2834,N_1714);
nor U3008 (N_3008,N_2992,N_2122);
or U3009 (N_3009,N_2606,N_2556);
nor U3010 (N_3010,N_1698,N_2393);
or U3011 (N_3011,N_1543,N_1519);
and U3012 (N_3012,N_2831,N_1921);
nand U3013 (N_3013,N_1821,N_2760);
nor U3014 (N_3014,N_1914,N_2068);
xnor U3015 (N_3015,N_1783,N_2330);
nor U3016 (N_3016,N_2750,N_2329);
nand U3017 (N_3017,N_2477,N_1516);
xor U3018 (N_3018,N_2396,N_2662);
or U3019 (N_3019,N_2256,N_1889);
or U3020 (N_3020,N_2153,N_1829);
and U3021 (N_3021,N_1624,N_1932);
xnor U3022 (N_3022,N_1637,N_2412);
nand U3023 (N_3023,N_2217,N_1562);
nor U3024 (N_3024,N_2398,N_2912);
nand U3025 (N_3025,N_1741,N_1719);
and U3026 (N_3026,N_2213,N_2843);
nand U3027 (N_3027,N_1617,N_1884);
xor U3028 (N_3028,N_2832,N_2620);
nand U3029 (N_3029,N_1920,N_2460);
nor U3030 (N_3030,N_1535,N_2778);
xor U3031 (N_3031,N_2715,N_2365);
nor U3032 (N_3032,N_1700,N_2524);
xnor U3033 (N_3033,N_2072,N_1742);
nand U3034 (N_3034,N_2056,N_2325);
xor U3035 (N_3035,N_2139,N_2573);
or U3036 (N_3036,N_1572,N_2768);
or U3037 (N_3037,N_2611,N_2497);
xor U3038 (N_3038,N_1752,N_2697);
nor U3039 (N_3039,N_2050,N_1585);
xor U3040 (N_3040,N_1588,N_2589);
nor U3041 (N_3041,N_2193,N_2819);
or U3042 (N_3042,N_2907,N_1899);
nand U3043 (N_3043,N_2609,N_2257);
xnor U3044 (N_3044,N_1806,N_2541);
xnor U3045 (N_3045,N_2227,N_2743);
and U3046 (N_3046,N_2306,N_2945);
or U3047 (N_3047,N_2592,N_1848);
or U3048 (N_3048,N_1892,N_2925);
and U3049 (N_3049,N_1552,N_1996);
or U3050 (N_3050,N_2436,N_2516);
and U3051 (N_3051,N_1680,N_1929);
xnor U3052 (N_3052,N_2356,N_2826);
and U3053 (N_3053,N_1563,N_2002);
nor U3054 (N_3054,N_1608,N_1739);
xor U3055 (N_3055,N_2132,N_1837);
nand U3056 (N_3056,N_2563,N_1715);
and U3057 (N_3057,N_2141,N_2319);
nand U3058 (N_3058,N_1604,N_2297);
nand U3059 (N_3059,N_1668,N_2560);
or U3060 (N_3060,N_2805,N_2904);
or U3061 (N_3061,N_2196,N_1747);
nor U3062 (N_3062,N_2010,N_2322);
nor U3063 (N_3063,N_1717,N_2806);
nor U3064 (N_3064,N_2271,N_2162);
nand U3065 (N_3065,N_1693,N_1626);
or U3066 (N_3066,N_2461,N_1690);
xnor U3067 (N_3067,N_2532,N_1973);
xnor U3068 (N_3068,N_2980,N_1749);
or U3069 (N_3069,N_2375,N_1520);
nor U3070 (N_3070,N_1906,N_2788);
and U3071 (N_3071,N_2966,N_2394);
or U3072 (N_3072,N_1793,N_2373);
nand U3073 (N_3073,N_2353,N_1746);
xor U3074 (N_3074,N_2995,N_1732);
nor U3075 (N_3075,N_2245,N_2440);
xor U3076 (N_3076,N_1897,N_2896);
nand U3077 (N_3077,N_1517,N_1726);
xnor U3078 (N_3078,N_1982,N_2379);
nor U3079 (N_3079,N_2618,N_2695);
nand U3080 (N_3080,N_1936,N_1578);
nand U3081 (N_3081,N_2169,N_1740);
xor U3082 (N_3082,N_1901,N_2865);
and U3083 (N_3083,N_2936,N_2200);
or U3084 (N_3084,N_2846,N_1623);
xnor U3085 (N_3085,N_1787,N_2031);
nand U3086 (N_3086,N_2565,N_1547);
and U3087 (N_3087,N_2019,N_2472);
or U3088 (N_3088,N_2442,N_1814);
xor U3089 (N_3089,N_1722,N_2228);
nand U3090 (N_3090,N_2463,N_2338);
xnor U3091 (N_3091,N_2190,N_2085);
nand U3092 (N_3092,N_2417,N_2007);
xor U3093 (N_3093,N_2352,N_1679);
and U3094 (N_3094,N_2029,N_2886);
and U3095 (N_3095,N_2130,N_2474);
nand U3096 (N_3096,N_2804,N_1734);
nor U3097 (N_3097,N_2827,N_2889);
or U3098 (N_3098,N_2575,N_1536);
and U3099 (N_3099,N_1580,N_2549);
or U3100 (N_3100,N_2158,N_1931);
xnor U3101 (N_3101,N_2685,N_2900);
or U3102 (N_3102,N_2816,N_2645);
nand U3103 (N_3103,N_2717,N_1956);
xor U3104 (N_3104,N_1810,N_2243);
xor U3105 (N_3105,N_2446,N_2374);
xor U3106 (N_3106,N_2042,N_1876);
nor U3107 (N_3107,N_2178,N_2950);
or U3108 (N_3108,N_2903,N_1620);
nor U3109 (N_3109,N_2071,N_1754);
nor U3110 (N_3110,N_2649,N_2807);
nor U3111 (N_3111,N_2439,N_2933);
xnor U3112 (N_3112,N_2792,N_2863);
and U3113 (N_3113,N_1840,N_2829);
xor U3114 (N_3114,N_2429,N_2599);
nor U3115 (N_3115,N_2756,N_1603);
nand U3116 (N_3116,N_2779,N_2718);
xnor U3117 (N_3117,N_2836,N_1774);
nor U3118 (N_3118,N_2331,N_2948);
nand U3119 (N_3119,N_1706,N_2419);
xnor U3120 (N_3120,N_1595,N_2150);
or U3121 (N_3121,N_2687,N_1720);
nand U3122 (N_3122,N_1566,N_2738);
or U3123 (N_3123,N_2958,N_2959);
xnor U3124 (N_3124,N_2894,N_2363);
and U3125 (N_3125,N_2328,N_1937);
nand U3126 (N_3126,N_2651,N_2800);
or U3127 (N_3127,N_2283,N_2005);
or U3128 (N_3128,N_2608,N_2108);
nor U3129 (N_3129,N_2437,N_2918);
xnor U3130 (N_3130,N_2411,N_1994);
xnor U3131 (N_3131,N_2164,N_2841);
nor U3132 (N_3132,N_1965,N_2521);
nand U3133 (N_3133,N_2577,N_2354);
or U3134 (N_3134,N_1805,N_2252);
nor U3135 (N_3135,N_2702,N_1970);
nand U3136 (N_3136,N_2548,N_2594);
nand U3137 (N_3137,N_1912,N_1606);
and U3138 (N_3138,N_2692,N_2910);
nand U3139 (N_3139,N_2464,N_1648);
nand U3140 (N_3140,N_2313,N_2064);
and U3141 (N_3141,N_2152,N_1511);
or U3142 (N_3142,N_2746,N_2659);
or U3143 (N_3143,N_2928,N_1775);
or U3144 (N_3144,N_2766,N_2189);
or U3145 (N_3145,N_2192,N_2110);
or U3146 (N_3146,N_1900,N_2681);
nor U3147 (N_3147,N_2047,N_2041);
or U3148 (N_3148,N_2569,N_2454);
and U3149 (N_3149,N_1716,N_2448);
nor U3150 (N_3150,N_2908,N_2091);
xor U3151 (N_3151,N_2898,N_2916);
and U3152 (N_3152,N_2345,N_2858);
xor U3153 (N_3153,N_2947,N_2961);
and U3154 (N_3154,N_2348,N_2869);
or U3155 (N_3155,N_2501,N_2057);
or U3156 (N_3156,N_2654,N_2126);
and U3157 (N_3157,N_2376,N_2597);
nand U3158 (N_3158,N_1765,N_2061);
xor U3159 (N_3159,N_1725,N_1681);
or U3160 (N_3160,N_2172,N_2989);
nand U3161 (N_3161,N_2333,N_2462);
and U3162 (N_3162,N_1735,N_2693);
nor U3163 (N_3163,N_1853,N_1873);
nand U3164 (N_3164,N_2881,N_1813);
nor U3165 (N_3165,N_2973,N_2380);
nor U3166 (N_3166,N_2775,N_1707);
or U3167 (N_3167,N_2100,N_2099);
xor U3168 (N_3168,N_1611,N_2629);
and U3169 (N_3169,N_2991,N_1660);
and U3170 (N_3170,N_1894,N_2647);
and U3171 (N_3171,N_2677,N_2390);
or U3172 (N_3172,N_2505,N_1764);
and U3173 (N_3173,N_2815,N_2929);
nor U3174 (N_3174,N_2054,N_2183);
or U3175 (N_3175,N_2246,N_1695);
xnor U3176 (N_3176,N_1812,N_2763);
and U3177 (N_3177,N_2699,N_1939);
and U3178 (N_3178,N_2730,N_2264);
nor U3179 (N_3179,N_1541,N_2711);
xnor U3180 (N_3180,N_2744,N_2906);
and U3181 (N_3181,N_1819,N_2690);
and U3182 (N_3182,N_1928,N_2784);
or U3183 (N_3183,N_1957,N_2457);
and U3184 (N_3184,N_2584,N_2737);
and U3185 (N_3185,N_2378,N_2368);
xnor U3186 (N_3186,N_2105,N_1553);
or U3187 (N_3187,N_2201,N_2239);
nor U3188 (N_3188,N_1639,N_2344);
nor U3189 (N_3189,N_1630,N_1784);
or U3190 (N_3190,N_2568,N_2403);
or U3191 (N_3191,N_2250,N_2128);
xnor U3192 (N_3192,N_1670,N_2957);
and U3193 (N_3193,N_1797,N_2926);
and U3194 (N_3194,N_1915,N_2976);
nor U3195 (N_3195,N_2159,N_2724);
and U3196 (N_3196,N_1745,N_2103);
nand U3197 (N_3197,N_2180,N_1771);
or U3198 (N_3198,N_1601,N_2721);
nand U3199 (N_3199,N_2154,N_1993);
and U3200 (N_3200,N_1594,N_1835);
nor U3201 (N_3201,N_2755,N_1654);
nand U3202 (N_3202,N_1869,N_1718);
xor U3203 (N_3203,N_2796,N_2222);
or U3204 (N_3204,N_1916,N_1788);
nand U3205 (N_3205,N_2665,N_2397);
or U3206 (N_3206,N_2013,N_2012);
or U3207 (N_3207,N_2316,N_1529);
or U3208 (N_3208,N_2281,N_2705);
and U3209 (N_3209,N_2817,N_1966);
xor U3210 (N_3210,N_2493,N_2596);
nand U3211 (N_3211,N_2850,N_1804);
and U3212 (N_3212,N_1988,N_2514);
xor U3213 (N_3213,N_2289,N_2935);
nor U3214 (N_3214,N_1583,N_1978);
nor U3215 (N_3215,N_2088,N_2294);
or U3216 (N_3216,N_2129,N_1945);
xor U3217 (N_3217,N_2234,N_2495);
or U3218 (N_3218,N_1859,N_2237);
nor U3219 (N_3219,N_2557,N_1618);
nand U3220 (N_3220,N_1977,N_1591);
nand U3221 (N_3221,N_2288,N_2102);
and U3222 (N_3222,N_2435,N_2335);
and U3223 (N_3223,N_1867,N_2707);
nor U3224 (N_3224,N_2628,N_2220);
nor U3225 (N_3225,N_1513,N_2739);
and U3226 (N_3226,N_1712,N_2955);
and U3227 (N_3227,N_2547,N_2476);
xnor U3228 (N_3228,N_2298,N_2663);
or U3229 (N_3229,N_2934,N_1832);
nand U3230 (N_3230,N_2342,N_2181);
nand U3231 (N_3231,N_1678,N_2890);
xnor U3232 (N_3232,N_2409,N_2769);
nor U3233 (N_3233,N_1697,N_2847);
or U3234 (N_3234,N_1757,N_1522);
xor U3235 (N_3235,N_2144,N_2430);
nand U3236 (N_3236,N_2602,N_1556);
xor U3237 (N_3237,N_2943,N_1801);
and U3238 (N_3238,N_1532,N_1649);
nand U3239 (N_3239,N_2350,N_2388);
nor U3240 (N_3240,N_2975,N_1587);
and U3241 (N_3241,N_2771,N_2075);
xor U3242 (N_3242,N_1908,N_2458);
and U3243 (N_3243,N_2969,N_1918);
xnor U3244 (N_3244,N_1773,N_1655);
or U3245 (N_3245,N_1568,N_2166);
nor U3246 (N_3246,N_1686,N_1694);
nor U3247 (N_3247,N_2688,N_2253);
nand U3248 (N_3248,N_2481,N_2828);
or U3249 (N_3249,N_2723,N_2299);
and U3250 (N_3250,N_1809,N_1785);
or U3251 (N_3251,N_2595,N_2094);
xor U3252 (N_3252,N_2587,N_2482);
nand U3253 (N_3253,N_2814,N_1593);
nor U3254 (N_3254,N_2679,N_1531);
xor U3255 (N_3255,N_1653,N_2445);
nand U3256 (N_3256,N_2875,N_1650);
nor U3257 (N_3257,N_1634,N_1910);
and U3258 (N_3258,N_2156,N_2490);
xor U3259 (N_3259,N_2523,N_2731);
nor U3260 (N_3260,N_1685,N_2650);
xnor U3261 (N_3261,N_2479,N_1733);
xor U3262 (N_3262,N_2372,N_2658);
nor U3263 (N_3263,N_1885,N_2116);
nand U3264 (N_3264,N_2455,N_1913);
xor U3265 (N_3265,N_2527,N_2182);
xnor U3266 (N_3266,N_2053,N_1570);
and U3267 (N_3267,N_2024,N_1909);
and U3268 (N_3268,N_2580,N_2987);
or U3269 (N_3269,N_2349,N_1811);
or U3270 (N_3270,N_2683,N_2802);
nor U3271 (N_3271,N_2623,N_1579);
or U3272 (N_3272,N_1644,N_2968);
or U3273 (N_3273,N_2552,N_2962);
or U3274 (N_3274,N_2364,N_2367);
nand U3275 (N_3275,N_2518,N_2079);
nor U3276 (N_3276,N_1687,N_2931);
xor U3277 (N_3277,N_2070,N_1709);
and U3278 (N_3278,N_2891,N_2009);
or U3279 (N_3279,N_2478,N_2515);
and U3280 (N_3280,N_1632,N_1948);
nand U3281 (N_3281,N_2612,N_1631);
nor U3282 (N_3282,N_2293,N_1628);
nor U3283 (N_3283,N_2564,N_1855);
or U3284 (N_3284,N_2536,N_1953);
or U3285 (N_3285,N_2083,N_2074);
xnor U3286 (N_3286,N_1661,N_1960);
or U3287 (N_3287,N_2276,N_1696);
xor U3288 (N_3288,N_2809,N_1665);
nand U3289 (N_3289,N_1751,N_2785);
and U3290 (N_3290,N_2972,N_2725);
nor U3291 (N_3291,N_1992,N_2058);
nand U3292 (N_3292,N_2000,N_1898);
and U3293 (N_3293,N_1565,N_2670);
or U3294 (N_3294,N_2915,N_1711);
or U3295 (N_3295,N_2418,N_1792);
xnor U3296 (N_3296,N_2242,N_2653);
xnor U3297 (N_3297,N_1807,N_2701);
nand U3298 (N_3298,N_2438,N_2320);
nor U3299 (N_3299,N_1592,N_2503);
nand U3300 (N_3300,N_1564,N_2014);
and U3301 (N_3301,N_2884,N_2055);
or U3302 (N_3302,N_2888,N_1704);
and U3303 (N_3303,N_2290,N_1575);
xnor U3304 (N_3304,N_2751,N_2346);
or U3305 (N_3305,N_2939,N_1523);
and U3306 (N_3306,N_1760,N_2032);
nand U3307 (N_3307,N_1833,N_2261);
nand U3308 (N_3308,N_2160,N_2211);
xnor U3309 (N_3309,N_2808,N_1500);
and U3310 (N_3310,N_2726,N_2332);
nor U3311 (N_3311,N_2341,N_2586);
xnor U3312 (N_3312,N_2842,N_1574);
nor U3313 (N_3313,N_2317,N_2801);
xnor U3314 (N_3314,N_1984,N_2997);
nor U3315 (N_3315,N_1769,N_2311);
and U3316 (N_3316,N_2640,N_1507);
or U3317 (N_3317,N_1895,N_2544);
xor U3318 (N_3318,N_2880,N_2840);
or U3319 (N_3319,N_1944,N_2308);
nor U3320 (N_3320,N_2913,N_2839);
nor U3321 (N_3321,N_2104,N_1951);
nand U3322 (N_3322,N_2021,N_2600);
or U3323 (N_3323,N_2639,N_1638);
or U3324 (N_3324,N_2266,N_1567);
or U3325 (N_3325,N_2698,N_2415);
or U3326 (N_3326,N_2535,N_2508);
xnor U3327 (N_3327,N_2295,N_2512);
and U3328 (N_3328,N_2231,N_2605);
nor U3329 (N_3329,N_2451,N_1605);
nand U3330 (N_3330,N_2097,N_1864);
nand U3331 (N_3331,N_1986,N_1633);
nor U3332 (N_3332,N_2305,N_2066);
nor U3333 (N_3333,N_1515,N_2893);
nor U3334 (N_3334,N_1872,N_1860);
xor U3335 (N_3335,N_2579,N_1689);
nand U3336 (N_3336,N_2835,N_1600);
nand U3337 (N_3337,N_2347,N_2984);
or U3338 (N_3338,N_2355,N_2135);
or U3339 (N_3339,N_2619,N_1822);
and U3340 (N_3340,N_2096,N_2732);
xor U3341 (N_3341,N_2638,N_1941);
nand U3342 (N_3342,N_1691,N_1673);
and U3343 (N_3343,N_2059,N_2043);
nor U3344 (N_3344,N_2525,N_1658);
and U3345 (N_3345,N_2036,N_1799);
or U3346 (N_3346,N_1907,N_1891);
xor U3347 (N_3347,N_2507,N_2080);
nand U3348 (N_3348,N_1942,N_1954);
nand U3349 (N_3349,N_2131,N_2204);
nor U3350 (N_3350,N_2336,N_2315);
and U3351 (N_3351,N_2990,N_2274);
and U3352 (N_3352,N_1607,N_2862);
xor U3353 (N_3353,N_1710,N_2044);
nor U3354 (N_3354,N_2545,N_2422);
xor U3355 (N_3355,N_1551,N_1736);
nand U3356 (N_3356,N_2845,N_2664);
or U3357 (N_3357,N_2296,N_2360);
xor U3358 (N_3358,N_2870,N_1870);
nor U3359 (N_3359,N_2185,N_2395);
or U3360 (N_3360,N_1759,N_2897);
xor U3361 (N_3361,N_2849,N_2996);
xnor U3362 (N_3362,N_2566,N_2197);
xnor U3363 (N_3363,N_2003,N_2682);
xnor U3364 (N_3364,N_1753,N_1616);
nor U3365 (N_3365,N_2033,N_1962);
xor U3366 (N_3366,N_1879,N_2956);
and U3367 (N_3367,N_1571,N_2113);
and U3368 (N_3368,N_2269,N_1713);
nor U3369 (N_3369,N_1657,N_1868);
or U3370 (N_3370,N_1850,N_1705);
and U3371 (N_3371,N_2877,N_1763);
xnor U3372 (N_3372,N_2387,N_2045);
xnor U3373 (N_3373,N_2389,N_2284);
xnor U3374 (N_3374,N_1508,N_1845);
nor U3375 (N_3375,N_2818,N_2225);
xnor U3376 (N_3376,N_2016,N_2273);
or U3377 (N_3377,N_2466,N_2520);
xnor U3378 (N_3378,N_1796,N_1619);
nand U3379 (N_3379,N_1573,N_2669);
nor U3380 (N_3380,N_2964,N_2151);
xor U3381 (N_3381,N_2291,N_2475);
and U3382 (N_3382,N_2001,N_1534);
or U3383 (N_3383,N_1998,N_2369);
xnor U3384 (N_3384,N_2526,N_1645);
and U3385 (N_3385,N_1599,N_1659);
and U3386 (N_3386,N_1526,N_2203);
or U3387 (N_3387,N_1925,N_2148);
nand U3388 (N_3388,N_2855,N_2147);
and U3389 (N_3389,N_2095,N_2517);
xor U3390 (N_3390,N_2696,N_1990);
or U3391 (N_3391,N_2138,N_2614);
and U3392 (N_3392,N_2810,N_2300);
nand U3393 (N_3393,N_1902,N_1947);
nand U3394 (N_3394,N_2255,N_2710);
nor U3395 (N_3395,N_2302,N_2876);
xnor U3396 (N_3396,N_2263,N_1502);
nor U3397 (N_3397,N_2741,N_1857);
nand U3398 (N_3398,N_1974,N_1949);
or U3399 (N_3399,N_2971,N_2830);
nor U3400 (N_3400,N_1896,N_2077);
xnor U3401 (N_3401,N_2187,N_2540);
and U3402 (N_3402,N_1961,N_1924);
nand U3403 (N_3403,N_2473,N_1952);
or U3404 (N_3404,N_1836,N_2431);
and U3405 (N_3405,N_1555,N_1817);
nand U3406 (N_3406,N_2999,N_2089);
xnor U3407 (N_3407,N_1967,N_2510);
or U3408 (N_3408,N_2981,N_1923);
nand U3409 (N_3409,N_2456,N_2616);
and U3410 (N_3410,N_2634,N_2416);
nor U3411 (N_3411,N_1770,N_2229);
nor U3412 (N_3412,N_1729,N_2408);
xor U3413 (N_3413,N_2459,N_2887);
xor U3414 (N_3414,N_2709,N_1926);
nand U3415 (N_3415,N_2661,N_2856);
nand U3416 (N_3416,N_1786,N_2381);
and U3417 (N_3417,N_2660,N_2248);
or U3418 (N_3418,N_2578,N_2254);
nor U3419 (N_3419,N_2223,N_2321);
xor U3420 (N_3420,N_1737,N_2534);
xnor U3421 (N_3421,N_1561,N_2790);
nand U3422 (N_3422,N_1981,N_2039);
or U3423 (N_3423,N_2167,N_1930);
nand U3424 (N_3424,N_2883,N_1995);
xor U3425 (N_3425,N_1688,N_1509);
xor U3426 (N_3426,N_2023,N_2757);
nor U3427 (N_3427,N_1946,N_2140);
or U3428 (N_3428,N_1767,N_2037);
nand U3429 (N_3429,N_2312,N_2528);
and U3430 (N_3430,N_2770,N_2851);
or U3431 (N_3431,N_2467,N_2864);
xor U3432 (N_3432,N_2470,N_2215);
nand U3433 (N_3433,N_1692,N_2226);
and U3434 (N_3434,N_2844,N_2538);
nand U3435 (N_3435,N_2646,N_2951);
nand U3436 (N_3436,N_2214,N_1636);
xor U3437 (N_3437,N_2424,N_2700);
and U3438 (N_3438,N_2879,N_2892);
and U3439 (N_3439,N_2601,N_2484);
nand U3440 (N_3440,N_2433,N_2452);
xnor U3441 (N_3441,N_2530,N_2798);
xnor U3442 (N_3442,N_2576,N_1979);
nor U3443 (N_3443,N_2519,N_2773);
and U3444 (N_3444,N_1544,N_1504);
or U3445 (N_3445,N_2644,N_2286);
nor U3446 (N_3446,N_1577,N_1919);
or U3447 (N_3447,N_2414,N_1789);
or U3448 (N_3448,N_1539,N_2983);
and U3449 (N_3449,N_2780,N_1514);
nor U3450 (N_3450,N_2307,N_1841);
nor U3451 (N_3451,N_2030,N_2247);
or U3452 (N_3452,N_1971,N_2413);
nand U3453 (N_3453,N_2713,N_2407);
xnor U3454 (N_3454,N_1554,N_2708);
xor U3455 (N_3455,N_2967,N_2209);
nand U3456 (N_3456,N_2531,N_1525);
xnor U3457 (N_3457,N_1596,N_2919);
or U3458 (N_3458,N_1985,N_2714);
and U3459 (N_3459,N_2781,N_1969);
and U3460 (N_3460,N_1590,N_2235);
and U3461 (N_3461,N_2018,N_1602);
or U3462 (N_3462,N_2309,N_2143);
and U3463 (N_3463,N_2668,N_2729);
xor U3464 (N_3464,N_1683,N_2598);
xnor U3465 (N_3465,N_2684,N_1675);
and U3466 (N_3466,N_1922,N_1586);
or U3467 (N_3467,N_2006,N_2868);
nand U3468 (N_3468,N_2591,N_1950);
xnor U3469 (N_3469,N_2621,N_1597);
nand U3470 (N_3470,N_2198,N_2823);
and U3471 (N_3471,N_2820,N_2613);
nor U3472 (N_3472,N_2813,N_2240);
or U3473 (N_3473,N_2405,N_2485);
nand U3474 (N_3474,N_2118,N_2207);
nand U3475 (N_3475,N_2867,N_1791);
or U3476 (N_3476,N_1802,N_2326);
xnor U3477 (N_3477,N_2086,N_1621);
xor U3478 (N_3478,N_1911,N_1987);
xnor U3479 (N_3479,N_2902,N_1524);
or U3480 (N_3480,N_1794,N_1999);
nand U3481 (N_3481,N_2028,N_2314);
xor U3482 (N_3482,N_2370,N_2655);
or U3483 (N_3483,N_1968,N_2762);
and U3484 (N_3484,N_1843,N_2443);
nor U3485 (N_3485,N_2155,N_1991);
xor U3486 (N_3486,N_2993,N_2232);
nor U3487 (N_3487,N_2206,N_2772);
and U3488 (N_3488,N_2170,N_2107);
nand U3489 (N_3489,N_2146,N_1880);
xor U3490 (N_3490,N_1779,N_1940);
nor U3491 (N_3491,N_2303,N_2791);
xor U3492 (N_3492,N_1878,N_1518);
or U3493 (N_3493,N_2069,N_2953);
nand U3494 (N_3494,N_1545,N_2421);
nand U3495 (N_3495,N_2837,N_2383);
nor U3496 (N_3496,N_2511,N_2885);
or U3497 (N_3497,N_1671,N_2944);
and U3498 (N_3498,N_2604,N_1874);
or U3499 (N_3499,N_2359,N_2504);
and U3500 (N_3500,N_1838,N_1820);
xor U3501 (N_3501,N_2607,N_2977);
or U3502 (N_3502,N_2666,N_2109);
nor U3503 (N_3503,N_1904,N_2133);
and U3504 (N_3504,N_2090,N_2543);
xor U3505 (N_3505,N_1743,N_2078);
nor U3506 (N_3506,N_1669,N_2038);
nand U3507 (N_3507,N_1849,N_1744);
xor U3508 (N_3508,N_2799,N_2753);
xor U3509 (N_3509,N_1824,N_2432);
or U3510 (N_3510,N_1877,N_2793);
nor U3511 (N_3511,N_2453,N_2994);
and U3512 (N_3512,N_2930,N_1861);
nand U3513 (N_3513,N_2674,N_1800);
nand U3514 (N_3514,N_1865,N_1980);
nand U3515 (N_3515,N_2191,N_2838);
nor U3516 (N_3516,N_1955,N_2386);
nand U3517 (N_3517,N_2093,N_1762);
xor U3518 (N_3518,N_2539,N_1782);
nor U3519 (N_3519,N_2689,N_2238);
or U3520 (N_3520,N_1672,N_2149);
nand U3521 (N_3521,N_1677,N_2425);
and U3522 (N_3522,N_2174,N_1662);
nand U3523 (N_3523,N_2179,N_2774);
or U3524 (N_3524,N_2901,N_1890);
or U3525 (N_3525,N_1846,N_2188);
xnor U3526 (N_3526,N_2233,N_2025);
nor U3527 (N_3527,N_2988,N_2171);
and U3528 (N_3528,N_1780,N_2874);
nor U3529 (N_3529,N_2195,N_1851);
nor U3530 (N_3530,N_2942,N_2854);
and U3531 (N_3531,N_1808,N_2186);
and U3532 (N_3532,N_1703,N_2940);
xor U3533 (N_3533,N_2142,N_1663);
nand U3534 (N_3534,N_2624,N_2759);
or U3535 (N_3535,N_2492,N_2447);
and U3536 (N_3536,N_2060,N_2224);
nor U3537 (N_3537,N_2671,N_2385);
and U3538 (N_3538,N_2559,N_2351);
and U3539 (N_3539,N_1724,N_2212);
or U3540 (N_3540,N_2550,N_2917);
or U3541 (N_3541,N_1528,N_1646);
nand U3542 (N_3542,N_2163,N_2570);
nor U3543 (N_3543,N_2656,N_1842);
and U3544 (N_3544,N_2026,N_2046);
nor U3545 (N_3545,N_1537,N_1903);
and U3546 (N_3546,N_1844,N_2641);
xor U3547 (N_3547,N_2377,N_2636);
xnor U3548 (N_3548,N_1614,N_1893);
or U3549 (N_3549,N_2040,N_2811);
nand U3550 (N_3550,N_2859,N_1684);
or U3551 (N_3551,N_2410,N_2765);
nor U3552 (N_3552,N_2733,N_2265);
or U3553 (N_3553,N_2905,N_2716);
nor U3554 (N_3554,N_2049,N_2735);
or U3555 (N_3555,N_2982,N_2998);
and U3556 (N_3556,N_1830,N_2287);
nand U3557 (N_3557,N_1826,N_1815);
nand U3558 (N_3558,N_1530,N_1750);
or U3559 (N_3559,N_2853,N_2282);
and U3560 (N_3560,N_1542,N_2734);
nand U3561 (N_3561,N_2084,N_2491);
xnor U3562 (N_3562,N_2496,N_1550);
or U3563 (N_3563,N_2861,N_2857);
xnor U3564 (N_3564,N_2537,N_2909);
and U3565 (N_3565,N_1748,N_2210);
nand U3566 (N_3566,N_2051,N_2567);
and U3567 (N_3567,N_1641,N_1756);
or U3568 (N_3568,N_1852,N_1613);
nor U3569 (N_3569,N_2736,N_2626);
nand U3570 (N_3570,N_2633,N_2441);
or U3571 (N_3571,N_1501,N_1576);
or U3572 (N_3572,N_2301,N_2941);
xor U3573 (N_3573,N_1510,N_1887);
nor U3574 (N_3574,N_2366,N_2092);
and U3575 (N_3575,N_2361,N_2427);
and U3576 (N_3576,N_2426,N_2337);
nor U3577 (N_3577,N_2244,N_2761);
or U3578 (N_3578,N_2275,N_2101);
nand U3579 (N_3579,N_1559,N_2062);
xor U3580 (N_3580,N_1934,N_2081);
nand U3581 (N_3581,N_2219,N_2487);
or U3582 (N_3582,N_2787,N_1560);
or U3583 (N_3583,N_2937,N_1667);
nor U3584 (N_3584,N_2748,N_2157);
nor U3585 (N_3585,N_2119,N_1625);
nand U3586 (N_3586,N_1728,N_2728);
nand U3587 (N_3587,N_1557,N_2965);
xnor U3588 (N_3588,N_1652,N_2776);
xor U3589 (N_3589,N_2480,N_1768);
nor U3590 (N_3590,N_2588,N_2067);
nand U3591 (N_3591,N_2124,N_1997);
nand U3592 (N_3592,N_2742,N_2866);
or U3593 (N_3593,N_2450,N_1856);
or U3594 (N_3594,N_2173,N_2848);
or U3595 (N_3595,N_2622,N_2382);
and U3596 (N_3596,N_2136,N_1643);
or U3597 (N_3597,N_2583,N_1642);
or U3598 (N_3598,N_2529,N_2691);
nand U3599 (N_3599,N_2015,N_2444);
nand U3600 (N_3600,N_1790,N_2749);
nor U3601 (N_3601,N_2011,N_2680);
nand U3602 (N_3602,N_2357,N_1777);
and U3603 (N_3603,N_2986,N_2558);
xor U3604 (N_3604,N_2272,N_1503);
and U3605 (N_3605,N_2176,N_2581);
and U3606 (N_3606,N_2279,N_2134);
xor U3607 (N_3607,N_2574,N_2572);
nand U3608 (N_3608,N_1871,N_1883);
xnor U3609 (N_3609,N_2642,N_2582);
xnor U3610 (N_3610,N_2938,N_1761);
xor U3611 (N_3611,N_1538,N_1702);
nand U3612 (N_3612,N_2522,N_2571);
or U3613 (N_3613,N_2978,N_1546);
xor U3614 (N_3614,N_2675,N_2509);
or U3615 (N_3615,N_1828,N_2554);
or U3616 (N_3616,N_2985,N_2920);
xor U3617 (N_3617,N_2794,N_2292);
and U3618 (N_3618,N_2324,N_2334);
nand U3619 (N_3619,N_1958,N_2082);
or U3620 (N_3620,N_1866,N_1818);
nand U3621 (N_3621,N_2686,N_2615);
nand U3622 (N_3622,N_2216,N_2752);
or U3623 (N_3623,N_1858,N_1863);
nor U3624 (N_3624,N_2924,N_2391);
and U3625 (N_3625,N_1656,N_2551);
and U3626 (N_3626,N_1598,N_1506);
and U3627 (N_3627,N_2362,N_1730);
xnor U3628 (N_3628,N_2719,N_2625);
nand U3629 (N_3629,N_2262,N_2635);
or U3630 (N_3630,N_2873,N_2471);
and U3631 (N_3631,N_1933,N_2758);
xor U3632 (N_3632,N_2643,N_1629);
or U3633 (N_3633,N_2278,N_2034);
xnor U3634 (N_3634,N_2632,N_2208);
and U3635 (N_3635,N_1558,N_2555);
or U3636 (N_3636,N_1589,N_2161);
or U3637 (N_3637,N_1615,N_1627);
or U3638 (N_3638,N_2310,N_1776);
nor U3639 (N_3639,N_2008,N_1964);
nor U3640 (N_3640,N_2465,N_2434);
nand U3641 (N_3641,N_2251,N_2676);
nand U3642 (N_3642,N_2027,N_2502);
nor U3643 (N_3643,N_2340,N_2268);
nand U3644 (N_3644,N_1976,N_2789);
nand U3645 (N_3645,N_2922,N_2199);
nor U3646 (N_3646,N_2745,N_1640);
nand U3647 (N_3647,N_2704,N_2610);
xor U3648 (N_3648,N_2168,N_1610);
or U3649 (N_3649,N_2194,N_2657);
and U3650 (N_3650,N_2921,N_1888);
or U3651 (N_3651,N_2722,N_2533);
nand U3652 (N_3652,N_1983,N_2318);
nand U3653 (N_3653,N_2327,N_1521);
xnor U3654 (N_3654,N_1647,N_2184);
nor U3655 (N_3655,N_2488,N_2630);
nand U3656 (N_3656,N_2783,N_1781);
nor U3657 (N_3657,N_1972,N_2469);
xnor U3658 (N_3658,N_1622,N_1731);
xnor U3659 (N_3659,N_1881,N_2121);
nand U3660 (N_3660,N_2678,N_2694);
nor U3661 (N_3661,N_1664,N_2952);
nand U3662 (N_3662,N_1862,N_2483);
and U3663 (N_3663,N_2617,N_1975);
or U3664 (N_3664,N_1569,N_2114);
and U3665 (N_3665,N_2120,N_2822);
and U3666 (N_3666,N_2506,N_1875);
or U3667 (N_3667,N_2065,N_2260);
or U3668 (N_3668,N_1738,N_1581);
xor U3669 (N_3669,N_1847,N_2371);
xor U3670 (N_3670,N_1989,N_2177);
nand U3671 (N_3671,N_2230,N_2970);
or U3672 (N_3672,N_2111,N_2468);
and U3673 (N_3673,N_2205,N_2399);
nor U3674 (N_3674,N_1766,N_2786);
nor U3675 (N_3675,N_2401,N_2747);
or U3676 (N_3676,N_2648,N_2882);
or U3677 (N_3677,N_2812,N_2782);
and U3678 (N_3678,N_1825,N_2954);
xnor U3679 (N_3679,N_1823,N_2499);
and U3680 (N_3680,N_2400,N_2323);
and U3681 (N_3681,N_2087,N_1721);
or U3682 (N_3682,N_2927,N_2112);
and U3683 (N_3683,N_1886,N_2703);
and U3684 (N_3684,N_2871,N_2236);
nor U3685 (N_3685,N_1803,N_1831);
or U3686 (N_3686,N_1882,N_1701);
or U3687 (N_3687,N_1666,N_1772);
or U3688 (N_3688,N_2500,N_2878);
xor U3689 (N_3689,N_2270,N_1938);
and U3690 (N_3690,N_2165,N_1827);
nand U3691 (N_3691,N_1682,N_2241);
xor U3692 (N_3692,N_2932,N_2860);
nor U3693 (N_3693,N_1854,N_2603);
or U3694 (N_3694,N_1533,N_1676);
xnor U3695 (N_3695,N_1755,N_2652);
or U3696 (N_3696,N_2593,N_2343);
and U3697 (N_3697,N_2259,N_2852);
or U3698 (N_3698,N_1512,N_1612);
or U3699 (N_3699,N_1839,N_2249);
xor U3700 (N_3700,N_1943,N_1816);
nand U3701 (N_3701,N_2895,N_2048);
nor U3702 (N_3702,N_2117,N_2052);
and U3703 (N_3703,N_2020,N_2221);
xnor U3704 (N_3704,N_1549,N_2585);
xnor U3705 (N_3705,N_2175,N_2712);
nand U3706 (N_3706,N_1798,N_1758);
nor U3707 (N_3707,N_2285,N_2667);
xor U3708 (N_3708,N_2063,N_2946);
and U3709 (N_3709,N_2404,N_2073);
or U3710 (N_3710,N_2974,N_2258);
or U3711 (N_3711,N_1778,N_2004);
xnor U3712 (N_3712,N_2137,N_2899);
nor U3713 (N_3713,N_2267,N_2631);
nand U3714 (N_3714,N_2824,N_2740);
and U3715 (N_3715,N_2486,N_2754);
nor U3716 (N_3716,N_2627,N_1527);
nand U3717 (N_3717,N_2035,N_1917);
nand U3718 (N_3718,N_2833,N_2706);
or U3719 (N_3719,N_2821,N_2115);
nor U3720 (N_3720,N_2280,N_2145);
nand U3721 (N_3721,N_2127,N_2923);
xnor U3722 (N_3722,N_1505,N_1935);
or U3723 (N_3723,N_1582,N_2125);
or U3724 (N_3724,N_2979,N_2494);
nor U3725 (N_3725,N_2553,N_2392);
or U3726 (N_3726,N_2423,N_2406);
and U3727 (N_3727,N_2304,N_2637);
and U3728 (N_3728,N_2914,N_2672);
xnor U3729 (N_3729,N_1674,N_2098);
nand U3730 (N_3730,N_1699,N_1927);
nor U3731 (N_3731,N_2546,N_1635);
and U3732 (N_3732,N_2872,N_1609);
nor U3733 (N_3733,N_2825,N_2218);
and U3734 (N_3734,N_2562,N_2420);
nand U3735 (N_3735,N_2202,N_2949);
nor U3736 (N_3736,N_2449,N_2542);
nand U3737 (N_3737,N_2513,N_1959);
nand U3738 (N_3738,N_2963,N_2590);
nand U3739 (N_3739,N_2911,N_2384);
nand U3740 (N_3740,N_2803,N_2767);
and U3741 (N_3741,N_2358,N_2498);
and U3742 (N_3742,N_1963,N_1651);
and U3743 (N_3743,N_2727,N_1548);
nand U3744 (N_3744,N_2960,N_2489);
nor U3745 (N_3745,N_1723,N_1834);
xnor U3746 (N_3746,N_2797,N_2764);
nor U3747 (N_3747,N_1708,N_1727);
nor U3748 (N_3748,N_2720,N_2339);
and U3749 (N_3749,N_2123,N_1905);
nand U3750 (N_3750,N_2050,N_1891);
or U3751 (N_3751,N_1953,N_2319);
nand U3752 (N_3752,N_2897,N_2523);
or U3753 (N_3753,N_2077,N_2240);
and U3754 (N_3754,N_2158,N_1616);
nand U3755 (N_3755,N_1714,N_2175);
or U3756 (N_3756,N_2608,N_1647);
nor U3757 (N_3757,N_1885,N_2910);
and U3758 (N_3758,N_2027,N_1677);
xor U3759 (N_3759,N_2069,N_1927);
nand U3760 (N_3760,N_1684,N_2240);
or U3761 (N_3761,N_1849,N_2887);
nand U3762 (N_3762,N_2525,N_1752);
nor U3763 (N_3763,N_2400,N_2874);
nand U3764 (N_3764,N_1985,N_1755);
or U3765 (N_3765,N_2886,N_2005);
nor U3766 (N_3766,N_2132,N_2677);
and U3767 (N_3767,N_2706,N_2598);
xor U3768 (N_3768,N_1899,N_1508);
and U3769 (N_3769,N_2538,N_1776);
xor U3770 (N_3770,N_2147,N_1650);
nor U3771 (N_3771,N_2079,N_2440);
xor U3772 (N_3772,N_1651,N_2512);
or U3773 (N_3773,N_2406,N_1681);
nand U3774 (N_3774,N_2870,N_2147);
xor U3775 (N_3775,N_1723,N_2916);
and U3776 (N_3776,N_2720,N_2248);
xnor U3777 (N_3777,N_1605,N_2160);
nand U3778 (N_3778,N_2129,N_1922);
and U3779 (N_3779,N_1884,N_1820);
nor U3780 (N_3780,N_2358,N_2882);
and U3781 (N_3781,N_2795,N_2210);
or U3782 (N_3782,N_2101,N_2359);
and U3783 (N_3783,N_2656,N_2587);
xor U3784 (N_3784,N_2344,N_2527);
nor U3785 (N_3785,N_1964,N_2018);
nand U3786 (N_3786,N_1842,N_2918);
or U3787 (N_3787,N_2678,N_1760);
nand U3788 (N_3788,N_2420,N_2063);
or U3789 (N_3789,N_1739,N_2975);
xnor U3790 (N_3790,N_2073,N_1553);
xor U3791 (N_3791,N_2421,N_1847);
and U3792 (N_3792,N_1881,N_2018);
xnor U3793 (N_3793,N_2213,N_2265);
and U3794 (N_3794,N_2135,N_2696);
or U3795 (N_3795,N_1883,N_2562);
and U3796 (N_3796,N_2538,N_2980);
and U3797 (N_3797,N_1706,N_2319);
nor U3798 (N_3798,N_1591,N_2308);
and U3799 (N_3799,N_2928,N_1740);
and U3800 (N_3800,N_2316,N_1806);
or U3801 (N_3801,N_2583,N_1843);
nor U3802 (N_3802,N_2068,N_1623);
or U3803 (N_3803,N_2114,N_2911);
xnor U3804 (N_3804,N_1765,N_2639);
and U3805 (N_3805,N_1546,N_2917);
nor U3806 (N_3806,N_2027,N_1924);
nand U3807 (N_3807,N_2549,N_2155);
nand U3808 (N_3808,N_2275,N_2161);
and U3809 (N_3809,N_1646,N_2310);
xnor U3810 (N_3810,N_2709,N_2510);
or U3811 (N_3811,N_1906,N_2513);
or U3812 (N_3812,N_1537,N_1849);
and U3813 (N_3813,N_1962,N_1506);
xnor U3814 (N_3814,N_2075,N_1912);
or U3815 (N_3815,N_2747,N_2882);
nand U3816 (N_3816,N_2345,N_1556);
nor U3817 (N_3817,N_2075,N_2881);
xor U3818 (N_3818,N_2995,N_1587);
xnor U3819 (N_3819,N_2224,N_2496);
and U3820 (N_3820,N_2224,N_1587);
nand U3821 (N_3821,N_2070,N_1882);
and U3822 (N_3822,N_2329,N_2702);
or U3823 (N_3823,N_1762,N_2036);
or U3824 (N_3824,N_1801,N_2800);
xor U3825 (N_3825,N_2960,N_2499);
or U3826 (N_3826,N_2882,N_2921);
xnor U3827 (N_3827,N_1683,N_1606);
xnor U3828 (N_3828,N_2907,N_2060);
nand U3829 (N_3829,N_1875,N_2493);
nor U3830 (N_3830,N_2954,N_2952);
nor U3831 (N_3831,N_2234,N_2375);
nor U3832 (N_3832,N_2431,N_2079);
nand U3833 (N_3833,N_2480,N_2271);
xor U3834 (N_3834,N_2594,N_1620);
nor U3835 (N_3835,N_1544,N_1550);
nor U3836 (N_3836,N_1734,N_2257);
xor U3837 (N_3837,N_2182,N_2818);
and U3838 (N_3838,N_1583,N_1845);
or U3839 (N_3839,N_2676,N_1993);
and U3840 (N_3840,N_1508,N_1882);
or U3841 (N_3841,N_2734,N_2979);
nor U3842 (N_3842,N_1786,N_2451);
nand U3843 (N_3843,N_1816,N_1641);
or U3844 (N_3844,N_2049,N_1971);
and U3845 (N_3845,N_2060,N_1824);
xor U3846 (N_3846,N_2272,N_2635);
xor U3847 (N_3847,N_2541,N_2615);
xnor U3848 (N_3848,N_2645,N_1540);
nand U3849 (N_3849,N_2440,N_2661);
or U3850 (N_3850,N_2349,N_2274);
nor U3851 (N_3851,N_2728,N_2287);
or U3852 (N_3852,N_2153,N_2210);
nand U3853 (N_3853,N_1727,N_2035);
nand U3854 (N_3854,N_2393,N_1512);
xnor U3855 (N_3855,N_2336,N_1885);
or U3856 (N_3856,N_2922,N_2411);
nor U3857 (N_3857,N_2522,N_1715);
or U3858 (N_3858,N_1974,N_2474);
nand U3859 (N_3859,N_1669,N_1805);
xor U3860 (N_3860,N_2030,N_2013);
xnor U3861 (N_3861,N_2403,N_2045);
nand U3862 (N_3862,N_2065,N_2676);
nor U3863 (N_3863,N_2542,N_1731);
xnor U3864 (N_3864,N_1642,N_1954);
or U3865 (N_3865,N_2071,N_2195);
or U3866 (N_3866,N_2482,N_2705);
and U3867 (N_3867,N_2479,N_1719);
nor U3868 (N_3868,N_2329,N_1829);
and U3869 (N_3869,N_2364,N_2347);
xor U3870 (N_3870,N_2043,N_1823);
nand U3871 (N_3871,N_2145,N_2028);
nor U3872 (N_3872,N_2036,N_1594);
or U3873 (N_3873,N_2693,N_2780);
or U3874 (N_3874,N_2668,N_1511);
and U3875 (N_3875,N_2261,N_2316);
and U3876 (N_3876,N_2416,N_2274);
and U3877 (N_3877,N_1867,N_2363);
and U3878 (N_3878,N_1774,N_1501);
and U3879 (N_3879,N_1886,N_2352);
nor U3880 (N_3880,N_2031,N_2300);
and U3881 (N_3881,N_1828,N_2885);
or U3882 (N_3882,N_2534,N_2233);
nand U3883 (N_3883,N_1835,N_1755);
and U3884 (N_3884,N_1623,N_1961);
and U3885 (N_3885,N_1666,N_1616);
xor U3886 (N_3886,N_2839,N_2480);
nand U3887 (N_3887,N_1828,N_2802);
nor U3888 (N_3888,N_2148,N_2900);
xor U3889 (N_3889,N_2586,N_1697);
nor U3890 (N_3890,N_2429,N_1689);
and U3891 (N_3891,N_2175,N_2391);
xnor U3892 (N_3892,N_2259,N_1608);
nor U3893 (N_3893,N_1876,N_2243);
nor U3894 (N_3894,N_1892,N_2973);
or U3895 (N_3895,N_2657,N_2700);
or U3896 (N_3896,N_1908,N_1833);
nand U3897 (N_3897,N_1682,N_2320);
nand U3898 (N_3898,N_1864,N_1584);
nand U3899 (N_3899,N_1537,N_1934);
and U3900 (N_3900,N_2924,N_2548);
xnor U3901 (N_3901,N_2641,N_2497);
xor U3902 (N_3902,N_2190,N_2160);
or U3903 (N_3903,N_2572,N_1802);
nand U3904 (N_3904,N_2489,N_2670);
nand U3905 (N_3905,N_1695,N_2363);
xor U3906 (N_3906,N_2288,N_1658);
or U3907 (N_3907,N_2161,N_2925);
nand U3908 (N_3908,N_1858,N_1610);
nand U3909 (N_3909,N_1928,N_2371);
and U3910 (N_3910,N_2845,N_2366);
nor U3911 (N_3911,N_2800,N_2421);
or U3912 (N_3912,N_1533,N_2877);
and U3913 (N_3913,N_2895,N_2288);
nand U3914 (N_3914,N_2604,N_2620);
nor U3915 (N_3915,N_1612,N_2795);
nor U3916 (N_3916,N_1812,N_2142);
nor U3917 (N_3917,N_2295,N_2375);
and U3918 (N_3918,N_2759,N_2884);
nand U3919 (N_3919,N_1542,N_2868);
nor U3920 (N_3920,N_1500,N_2554);
nor U3921 (N_3921,N_2279,N_2403);
nor U3922 (N_3922,N_2694,N_2571);
and U3923 (N_3923,N_2579,N_1966);
nand U3924 (N_3924,N_1937,N_2973);
xor U3925 (N_3925,N_2013,N_2238);
xor U3926 (N_3926,N_2790,N_2463);
and U3927 (N_3927,N_1933,N_1572);
nand U3928 (N_3928,N_2928,N_2945);
nor U3929 (N_3929,N_1706,N_2467);
nand U3930 (N_3930,N_2772,N_2876);
nor U3931 (N_3931,N_2106,N_1764);
xor U3932 (N_3932,N_1701,N_2986);
nor U3933 (N_3933,N_2998,N_2855);
or U3934 (N_3934,N_2340,N_2835);
and U3935 (N_3935,N_1795,N_1769);
nand U3936 (N_3936,N_2657,N_1541);
or U3937 (N_3937,N_1947,N_1601);
xor U3938 (N_3938,N_2026,N_2430);
or U3939 (N_3939,N_2292,N_1856);
or U3940 (N_3940,N_2111,N_1517);
or U3941 (N_3941,N_2128,N_1965);
and U3942 (N_3942,N_1841,N_1611);
nor U3943 (N_3943,N_2053,N_2166);
nand U3944 (N_3944,N_1779,N_2639);
or U3945 (N_3945,N_2096,N_1957);
nand U3946 (N_3946,N_2789,N_1871);
nand U3947 (N_3947,N_2477,N_2334);
nor U3948 (N_3948,N_2711,N_1940);
or U3949 (N_3949,N_1884,N_2641);
xor U3950 (N_3950,N_1630,N_1859);
nand U3951 (N_3951,N_2845,N_2697);
nand U3952 (N_3952,N_1758,N_1742);
xnor U3953 (N_3953,N_1922,N_2498);
nand U3954 (N_3954,N_1832,N_2355);
or U3955 (N_3955,N_2412,N_2039);
and U3956 (N_3956,N_1761,N_1876);
xnor U3957 (N_3957,N_1520,N_2316);
nor U3958 (N_3958,N_2982,N_2232);
or U3959 (N_3959,N_1855,N_1588);
and U3960 (N_3960,N_1900,N_1666);
xnor U3961 (N_3961,N_2978,N_1571);
xnor U3962 (N_3962,N_2123,N_2308);
nand U3963 (N_3963,N_2393,N_2768);
nand U3964 (N_3964,N_2868,N_2708);
xor U3965 (N_3965,N_1986,N_1840);
or U3966 (N_3966,N_2606,N_2406);
nor U3967 (N_3967,N_1680,N_2615);
xnor U3968 (N_3968,N_2170,N_1864);
or U3969 (N_3969,N_1564,N_2339);
or U3970 (N_3970,N_2881,N_1923);
nand U3971 (N_3971,N_1599,N_2564);
or U3972 (N_3972,N_1530,N_2858);
or U3973 (N_3973,N_2923,N_2660);
or U3974 (N_3974,N_2687,N_1748);
or U3975 (N_3975,N_2826,N_1716);
nor U3976 (N_3976,N_2116,N_2922);
nor U3977 (N_3977,N_1722,N_1795);
or U3978 (N_3978,N_2723,N_1820);
or U3979 (N_3979,N_2861,N_2212);
nand U3980 (N_3980,N_2166,N_2915);
xor U3981 (N_3981,N_2000,N_2171);
nor U3982 (N_3982,N_1583,N_1848);
or U3983 (N_3983,N_2948,N_1833);
xor U3984 (N_3984,N_1739,N_2344);
nand U3985 (N_3985,N_2664,N_2265);
and U3986 (N_3986,N_1581,N_2407);
nand U3987 (N_3987,N_2966,N_2655);
and U3988 (N_3988,N_1933,N_2956);
xnor U3989 (N_3989,N_1770,N_2781);
xnor U3990 (N_3990,N_2693,N_2960);
nand U3991 (N_3991,N_2623,N_2503);
and U3992 (N_3992,N_1745,N_2337);
and U3993 (N_3993,N_1861,N_2638);
and U3994 (N_3994,N_1956,N_2874);
xor U3995 (N_3995,N_1765,N_2562);
or U3996 (N_3996,N_2156,N_1513);
and U3997 (N_3997,N_2511,N_2654);
or U3998 (N_3998,N_2818,N_2999);
xnor U3999 (N_3999,N_2981,N_2575);
nor U4000 (N_4000,N_2250,N_1883);
nand U4001 (N_4001,N_2089,N_2328);
nand U4002 (N_4002,N_1581,N_2463);
nor U4003 (N_4003,N_2455,N_2999);
and U4004 (N_4004,N_2486,N_2784);
and U4005 (N_4005,N_2703,N_2115);
and U4006 (N_4006,N_1686,N_2306);
nand U4007 (N_4007,N_2404,N_2176);
nor U4008 (N_4008,N_2423,N_2732);
nand U4009 (N_4009,N_2737,N_2751);
xor U4010 (N_4010,N_1555,N_1678);
nor U4011 (N_4011,N_2646,N_1565);
nor U4012 (N_4012,N_1609,N_1561);
xor U4013 (N_4013,N_2799,N_2503);
and U4014 (N_4014,N_1911,N_1853);
xor U4015 (N_4015,N_2354,N_2434);
or U4016 (N_4016,N_2917,N_1646);
xnor U4017 (N_4017,N_1699,N_2493);
nor U4018 (N_4018,N_2259,N_2209);
or U4019 (N_4019,N_1654,N_2413);
and U4020 (N_4020,N_1808,N_1725);
and U4021 (N_4021,N_1888,N_2164);
and U4022 (N_4022,N_1741,N_2444);
nand U4023 (N_4023,N_2110,N_2330);
nor U4024 (N_4024,N_1561,N_2159);
or U4025 (N_4025,N_1846,N_2549);
or U4026 (N_4026,N_1596,N_1547);
nor U4027 (N_4027,N_2415,N_2833);
xor U4028 (N_4028,N_2824,N_2132);
nor U4029 (N_4029,N_2598,N_2191);
or U4030 (N_4030,N_1587,N_1838);
xor U4031 (N_4031,N_2827,N_1640);
xnor U4032 (N_4032,N_2065,N_2334);
xor U4033 (N_4033,N_2575,N_2995);
and U4034 (N_4034,N_2973,N_1501);
nor U4035 (N_4035,N_2051,N_2227);
nor U4036 (N_4036,N_2423,N_2541);
nor U4037 (N_4037,N_2734,N_1648);
nand U4038 (N_4038,N_2746,N_1676);
nor U4039 (N_4039,N_2941,N_2861);
nor U4040 (N_4040,N_1668,N_2373);
and U4041 (N_4041,N_2973,N_1683);
and U4042 (N_4042,N_1622,N_2114);
nand U4043 (N_4043,N_2466,N_2646);
and U4044 (N_4044,N_2909,N_1564);
nand U4045 (N_4045,N_2804,N_1742);
nand U4046 (N_4046,N_1660,N_2548);
and U4047 (N_4047,N_1770,N_1668);
or U4048 (N_4048,N_2156,N_1605);
nand U4049 (N_4049,N_1890,N_2606);
or U4050 (N_4050,N_2685,N_2278);
and U4051 (N_4051,N_1738,N_1503);
nor U4052 (N_4052,N_1737,N_2812);
nor U4053 (N_4053,N_2629,N_1583);
xnor U4054 (N_4054,N_1826,N_1732);
nand U4055 (N_4055,N_2742,N_1883);
xor U4056 (N_4056,N_1843,N_1998);
or U4057 (N_4057,N_2231,N_1699);
nor U4058 (N_4058,N_2250,N_2012);
and U4059 (N_4059,N_2052,N_2896);
or U4060 (N_4060,N_2979,N_2094);
and U4061 (N_4061,N_2456,N_2415);
and U4062 (N_4062,N_1959,N_1974);
xnor U4063 (N_4063,N_2266,N_2730);
nand U4064 (N_4064,N_2437,N_1692);
nand U4065 (N_4065,N_2414,N_1778);
nor U4066 (N_4066,N_2862,N_2580);
nor U4067 (N_4067,N_1816,N_1900);
or U4068 (N_4068,N_1662,N_1942);
and U4069 (N_4069,N_1805,N_2075);
or U4070 (N_4070,N_2474,N_2058);
or U4071 (N_4071,N_2277,N_1996);
xnor U4072 (N_4072,N_2495,N_2366);
and U4073 (N_4073,N_2691,N_1875);
nor U4074 (N_4074,N_2981,N_1542);
and U4075 (N_4075,N_2334,N_1858);
nand U4076 (N_4076,N_1590,N_2024);
xnor U4077 (N_4077,N_2917,N_2673);
xnor U4078 (N_4078,N_1741,N_1688);
xor U4079 (N_4079,N_2397,N_1993);
and U4080 (N_4080,N_2562,N_2341);
and U4081 (N_4081,N_2579,N_2130);
and U4082 (N_4082,N_2708,N_1871);
or U4083 (N_4083,N_2979,N_2011);
nor U4084 (N_4084,N_2959,N_2821);
nor U4085 (N_4085,N_2703,N_2561);
nand U4086 (N_4086,N_2938,N_2883);
or U4087 (N_4087,N_1676,N_2000);
xnor U4088 (N_4088,N_2365,N_2202);
and U4089 (N_4089,N_2723,N_1865);
nor U4090 (N_4090,N_2974,N_1831);
xnor U4091 (N_4091,N_2404,N_2201);
nand U4092 (N_4092,N_2500,N_2461);
nand U4093 (N_4093,N_1663,N_2071);
or U4094 (N_4094,N_2985,N_2228);
and U4095 (N_4095,N_2204,N_2693);
or U4096 (N_4096,N_2104,N_2942);
nor U4097 (N_4097,N_2610,N_2242);
or U4098 (N_4098,N_1714,N_1667);
nor U4099 (N_4099,N_2331,N_2766);
xnor U4100 (N_4100,N_1695,N_1837);
or U4101 (N_4101,N_2276,N_2436);
or U4102 (N_4102,N_2143,N_2672);
nand U4103 (N_4103,N_2917,N_2911);
xor U4104 (N_4104,N_2657,N_1592);
and U4105 (N_4105,N_1613,N_2610);
xnor U4106 (N_4106,N_1965,N_2872);
or U4107 (N_4107,N_2975,N_2479);
or U4108 (N_4108,N_2693,N_2359);
nor U4109 (N_4109,N_1530,N_2377);
xnor U4110 (N_4110,N_1971,N_2452);
or U4111 (N_4111,N_1712,N_2965);
nor U4112 (N_4112,N_1727,N_2761);
or U4113 (N_4113,N_1561,N_1727);
nor U4114 (N_4114,N_2927,N_2649);
and U4115 (N_4115,N_1771,N_2955);
nand U4116 (N_4116,N_2976,N_2655);
nand U4117 (N_4117,N_2987,N_1840);
and U4118 (N_4118,N_2558,N_2478);
and U4119 (N_4119,N_2290,N_2630);
nand U4120 (N_4120,N_1704,N_1585);
or U4121 (N_4121,N_2721,N_2572);
nor U4122 (N_4122,N_2747,N_2986);
xnor U4123 (N_4123,N_1857,N_1562);
nand U4124 (N_4124,N_2127,N_2288);
nor U4125 (N_4125,N_1966,N_2874);
nor U4126 (N_4126,N_2967,N_2636);
and U4127 (N_4127,N_2867,N_2519);
nor U4128 (N_4128,N_1705,N_1521);
nor U4129 (N_4129,N_2933,N_1557);
nand U4130 (N_4130,N_2659,N_2591);
nor U4131 (N_4131,N_1657,N_2826);
xor U4132 (N_4132,N_2211,N_2380);
and U4133 (N_4133,N_2961,N_2489);
and U4134 (N_4134,N_1600,N_2446);
or U4135 (N_4135,N_2922,N_2983);
xnor U4136 (N_4136,N_1694,N_2754);
or U4137 (N_4137,N_2689,N_1560);
nand U4138 (N_4138,N_2383,N_2202);
xnor U4139 (N_4139,N_2136,N_2174);
nand U4140 (N_4140,N_1594,N_2541);
xor U4141 (N_4141,N_1572,N_1797);
or U4142 (N_4142,N_2804,N_1867);
nor U4143 (N_4143,N_2289,N_2215);
nand U4144 (N_4144,N_2822,N_2688);
nand U4145 (N_4145,N_1964,N_1744);
xnor U4146 (N_4146,N_2633,N_2674);
nand U4147 (N_4147,N_2827,N_2477);
and U4148 (N_4148,N_2050,N_1516);
xor U4149 (N_4149,N_2727,N_2685);
nand U4150 (N_4150,N_2146,N_1713);
nand U4151 (N_4151,N_2759,N_1599);
xor U4152 (N_4152,N_1516,N_2719);
nor U4153 (N_4153,N_1890,N_2028);
and U4154 (N_4154,N_2520,N_1849);
and U4155 (N_4155,N_2838,N_2911);
and U4156 (N_4156,N_2176,N_1706);
nor U4157 (N_4157,N_2481,N_2809);
nand U4158 (N_4158,N_2080,N_1757);
nand U4159 (N_4159,N_1694,N_1847);
and U4160 (N_4160,N_2303,N_2263);
xor U4161 (N_4161,N_2511,N_1971);
and U4162 (N_4162,N_2155,N_2797);
xnor U4163 (N_4163,N_1987,N_1518);
or U4164 (N_4164,N_2199,N_1803);
and U4165 (N_4165,N_1967,N_1888);
nor U4166 (N_4166,N_2866,N_2912);
or U4167 (N_4167,N_2650,N_2726);
xnor U4168 (N_4168,N_1816,N_1840);
nor U4169 (N_4169,N_2408,N_1861);
nand U4170 (N_4170,N_2841,N_2619);
and U4171 (N_4171,N_1737,N_1838);
nor U4172 (N_4172,N_2853,N_1836);
nor U4173 (N_4173,N_2137,N_2879);
and U4174 (N_4174,N_1754,N_2843);
and U4175 (N_4175,N_1759,N_2948);
nor U4176 (N_4176,N_2119,N_1535);
or U4177 (N_4177,N_2557,N_1718);
nand U4178 (N_4178,N_2292,N_2389);
nand U4179 (N_4179,N_2208,N_2724);
nor U4180 (N_4180,N_1510,N_2983);
and U4181 (N_4181,N_2935,N_2068);
nand U4182 (N_4182,N_2368,N_2137);
xor U4183 (N_4183,N_1517,N_2665);
nand U4184 (N_4184,N_1974,N_2456);
or U4185 (N_4185,N_2253,N_2815);
or U4186 (N_4186,N_2370,N_1877);
and U4187 (N_4187,N_2091,N_2253);
or U4188 (N_4188,N_1664,N_1549);
nand U4189 (N_4189,N_1751,N_1801);
nand U4190 (N_4190,N_2530,N_2981);
nand U4191 (N_4191,N_1624,N_2528);
xnor U4192 (N_4192,N_2570,N_1959);
and U4193 (N_4193,N_2536,N_1909);
and U4194 (N_4194,N_2060,N_1764);
nor U4195 (N_4195,N_2648,N_1780);
nor U4196 (N_4196,N_2902,N_2259);
and U4197 (N_4197,N_2403,N_1615);
or U4198 (N_4198,N_2093,N_2318);
xor U4199 (N_4199,N_2439,N_2259);
or U4200 (N_4200,N_1796,N_1950);
nand U4201 (N_4201,N_2930,N_1586);
nand U4202 (N_4202,N_1802,N_2053);
xnor U4203 (N_4203,N_1739,N_2849);
xnor U4204 (N_4204,N_2541,N_2159);
and U4205 (N_4205,N_2707,N_2025);
and U4206 (N_4206,N_2821,N_2126);
or U4207 (N_4207,N_2491,N_1600);
nand U4208 (N_4208,N_2139,N_2750);
nand U4209 (N_4209,N_1920,N_2227);
nor U4210 (N_4210,N_2974,N_1539);
nand U4211 (N_4211,N_1950,N_2229);
and U4212 (N_4212,N_2942,N_1962);
xnor U4213 (N_4213,N_2781,N_2406);
xnor U4214 (N_4214,N_1826,N_2486);
xnor U4215 (N_4215,N_1612,N_1562);
and U4216 (N_4216,N_2953,N_2318);
nand U4217 (N_4217,N_2415,N_1978);
xnor U4218 (N_4218,N_2879,N_2123);
nand U4219 (N_4219,N_1996,N_2760);
and U4220 (N_4220,N_1646,N_2288);
nor U4221 (N_4221,N_2062,N_1817);
nor U4222 (N_4222,N_2259,N_1941);
xnor U4223 (N_4223,N_2844,N_2936);
nand U4224 (N_4224,N_1563,N_2541);
xnor U4225 (N_4225,N_2602,N_1950);
xor U4226 (N_4226,N_2746,N_2057);
or U4227 (N_4227,N_2863,N_2801);
nand U4228 (N_4228,N_2697,N_2807);
xor U4229 (N_4229,N_2305,N_2461);
xor U4230 (N_4230,N_2307,N_1814);
xnor U4231 (N_4231,N_2243,N_2198);
or U4232 (N_4232,N_2127,N_2599);
and U4233 (N_4233,N_2067,N_2402);
nand U4234 (N_4234,N_2720,N_1960);
nor U4235 (N_4235,N_2052,N_1965);
xor U4236 (N_4236,N_2891,N_1782);
nand U4237 (N_4237,N_2117,N_2808);
and U4238 (N_4238,N_2627,N_2276);
and U4239 (N_4239,N_2349,N_2857);
xnor U4240 (N_4240,N_2558,N_2779);
xnor U4241 (N_4241,N_2231,N_2857);
nand U4242 (N_4242,N_2747,N_2287);
nand U4243 (N_4243,N_2929,N_1840);
or U4244 (N_4244,N_1810,N_2664);
xnor U4245 (N_4245,N_2402,N_2954);
and U4246 (N_4246,N_2081,N_2808);
and U4247 (N_4247,N_2918,N_2375);
xor U4248 (N_4248,N_2839,N_2169);
nor U4249 (N_4249,N_2407,N_2423);
xor U4250 (N_4250,N_2085,N_2948);
xnor U4251 (N_4251,N_1707,N_2458);
and U4252 (N_4252,N_2262,N_2435);
nor U4253 (N_4253,N_2550,N_1659);
and U4254 (N_4254,N_1889,N_1841);
or U4255 (N_4255,N_1875,N_1886);
and U4256 (N_4256,N_2107,N_2275);
nor U4257 (N_4257,N_2572,N_1656);
xor U4258 (N_4258,N_2829,N_1622);
nor U4259 (N_4259,N_2104,N_2863);
xnor U4260 (N_4260,N_2937,N_2853);
or U4261 (N_4261,N_2922,N_2274);
nor U4262 (N_4262,N_1541,N_1733);
xnor U4263 (N_4263,N_2374,N_1503);
xor U4264 (N_4264,N_2856,N_1817);
xnor U4265 (N_4265,N_1703,N_1794);
nor U4266 (N_4266,N_1562,N_1840);
and U4267 (N_4267,N_2465,N_2260);
or U4268 (N_4268,N_1678,N_2262);
nand U4269 (N_4269,N_2141,N_1929);
nand U4270 (N_4270,N_2308,N_2936);
xor U4271 (N_4271,N_2876,N_1887);
and U4272 (N_4272,N_1566,N_2794);
xor U4273 (N_4273,N_2897,N_1703);
nor U4274 (N_4274,N_1631,N_1586);
nor U4275 (N_4275,N_1969,N_1665);
nand U4276 (N_4276,N_2992,N_2806);
or U4277 (N_4277,N_2191,N_2091);
nand U4278 (N_4278,N_1684,N_2512);
nand U4279 (N_4279,N_2239,N_1771);
nor U4280 (N_4280,N_2128,N_2679);
xor U4281 (N_4281,N_2582,N_1607);
or U4282 (N_4282,N_2694,N_1915);
xnor U4283 (N_4283,N_2888,N_2123);
xnor U4284 (N_4284,N_2327,N_2685);
xnor U4285 (N_4285,N_2651,N_2294);
xor U4286 (N_4286,N_1640,N_2757);
nand U4287 (N_4287,N_2641,N_2709);
nor U4288 (N_4288,N_2198,N_2641);
or U4289 (N_4289,N_2556,N_2853);
and U4290 (N_4290,N_1720,N_1695);
nor U4291 (N_4291,N_2386,N_1981);
and U4292 (N_4292,N_1957,N_2353);
nand U4293 (N_4293,N_2072,N_1829);
nor U4294 (N_4294,N_2310,N_2628);
and U4295 (N_4295,N_1671,N_2237);
nor U4296 (N_4296,N_2795,N_1725);
or U4297 (N_4297,N_1896,N_2304);
and U4298 (N_4298,N_2337,N_2454);
and U4299 (N_4299,N_1727,N_2888);
or U4300 (N_4300,N_2697,N_2338);
or U4301 (N_4301,N_2812,N_2776);
xor U4302 (N_4302,N_2912,N_2086);
nand U4303 (N_4303,N_2853,N_2691);
and U4304 (N_4304,N_1682,N_2589);
nand U4305 (N_4305,N_2241,N_2757);
or U4306 (N_4306,N_2382,N_1617);
and U4307 (N_4307,N_2119,N_2284);
nand U4308 (N_4308,N_2949,N_2069);
and U4309 (N_4309,N_2506,N_1528);
nand U4310 (N_4310,N_1815,N_2549);
and U4311 (N_4311,N_1908,N_2628);
and U4312 (N_4312,N_2190,N_2779);
xor U4313 (N_4313,N_2295,N_2223);
and U4314 (N_4314,N_2533,N_2848);
xor U4315 (N_4315,N_2622,N_2474);
or U4316 (N_4316,N_2986,N_2524);
nor U4317 (N_4317,N_1944,N_1789);
or U4318 (N_4318,N_2265,N_1507);
nand U4319 (N_4319,N_1740,N_1510);
and U4320 (N_4320,N_2524,N_2318);
xor U4321 (N_4321,N_2199,N_2655);
nand U4322 (N_4322,N_2764,N_2660);
nand U4323 (N_4323,N_1896,N_2767);
nand U4324 (N_4324,N_2975,N_1585);
and U4325 (N_4325,N_2932,N_2031);
nand U4326 (N_4326,N_1847,N_1839);
and U4327 (N_4327,N_2359,N_2512);
nor U4328 (N_4328,N_2126,N_2063);
nor U4329 (N_4329,N_2463,N_1763);
nor U4330 (N_4330,N_2348,N_2521);
nor U4331 (N_4331,N_1821,N_2845);
or U4332 (N_4332,N_1659,N_2868);
xnor U4333 (N_4333,N_2502,N_1623);
nor U4334 (N_4334,N_2817,N_2536);
nor U4335 (N_4335,N_2982,N_2473);
xnor U4336 (N_4336,N_1916,N_1844);
and U4337 (N_4337,N_2646,N_2257);
or U4338 (N_4338,N_2787,N_2426);
xnor U4339 (N_4339,N_1528,N_2985);
or U4340 (N_4340,N_1587,N_1772);
or U4341 (N_4341,N_1694,N_2954);
nor U4342 (N_4342,N_2062,N_2462);
nand U4343 (N_4343,N_2964,N_2097);
and U4344 (N_4344,N_2653,N_2747);
and U4345 (N_4345,N_2724,N_1544);
xnor U4346 (N_4346,N_2930,N_1576);
xor U4347 (N_4347,N_2988,N_2102);
or U4348 (N_4348,N_1636,N_1833);
nand U4349 (N_4349,N_2891,N_1607);
xor U4350 (N_4350,N_2320,N_2538);
xnor U4351 (N_4351,N_2714,N_2133);
and U4352 (N_4352,N_1728,N_2932);
nand U4353 (N_4353,N_2716,N_2766);
xnor U4354 (N_4354,N_2015,N_1825);
xnor U4355 (N_4355,N_2701,N_1876);
xnor U4356 (N_4356,N_2991,N_2177);
xnor U4357 (N_4357,N_2993,N_2815);
and U4358 (N_4358,N_2511,N_1704);
or U4359 (N_4359,N_1905,N_2827);
nor U4360 (N_4360,N_2219,N_1900);
xnor U4361 (N_4361,N_1818,N_2446);
and U4362 (N_4362,N_1641,N_2196);
xnor U4363 (N_4363,N_2373,N_2796);
xnor U4364 (N_4364,N_2266,N_2639);
or U4365 (N_4365,N_2243,N_1626);
nor U4366 (N_4366,N_2847,N_1896);
and U4367 (N_4367,N_2545,N_1657);
or U4368 (N_4368,N_2360,N_1873);
nor U4369 (N_4369,N_1695,N_2054);
xor U4370 (N_4370,N_2600,N_2147);
xor U4371 (N_4371,N_2494,N_1636);
xor U4372 (N_4372,N_2312,N_2534);
nand U4373 (N_4373,N_1665,N_1902);
and U4374 (N_4374,N_2328,N_2193);
xnor U4375 (N_4375,N_1779,N_2295);
xnor U4376 (N_4376,N_2877,N_2295);
or U4377 (N_4377,N_2649,N_1632);
xnor U4378 (N_4378,N_2219,N_2080);
nor U4379 (N_4379,N_2966,N_2088);
and U4380 (N_4380,N_2796,N_1858);
nor U4381 (N_4381,N_1795,N_2200);
nor U4382 (N_4382,N_1514,N_2717);
nand U4383 (N_4383,N_2524,N_2482);
nand U4384 (N_4384,N_2383,N_1707);
and U4385 (N_4385,N_2894,N_2193);
nor U4386 (N_4386,N_1916,N_1627);
and U4387 (N_4387,N_2497,N_1908);
nand U4388 (N_4388,N_2522,N_2507);
or U4389 (N_4389,N_2175,N_2884);
nor U4390 (N_4390,N_1590,N_2387);
and U4391 (N_4391,N_2642,N_2557);
xor U4392 (N_4392,N_2655,N_2376);
nand U4393 (N_4393,N_2465,N_2026);
nor U4394 (N_4394,N_2133,N_1892);
nand U4395 (N_4395,N_1693,N_2126);
nor U4396 (N_4396,N_2771,N_2952);
and U4397 (N_4397,N_2014,N_2602);
nor U4398 (N_4398,N_2139,N_2294);
nor U4399 (N_4399,N_2371,N_1999);
nor U4400 (N_4400,N_2237,N_2672);
or U4401 (N_4401,N_1624,N_1667);
and U4402 (N_4402,N_2663,N_2311);
and U4403 (N_4403,N_1506,N_2716);
nor U4404 (N_4404,N_2118,N_2945);
or U4405 (N_4405,N_1607,N_2817);
nor U4406 (N_4406,N_1709,N_2054);
xor U4407 (N_4407,N_2526,N_2291);
nand U4408 (N_4408,N_2083,N_2117);
or U4409 (N_4409,N_2480,N_1803);
nor U4410 (N_4410,N_2191,N_1756);
nand U4411 (N_4411,N_2645,N_2203);
or U4412 (N_4412,N_1836,N_2584);
xnor U4413 (N_4413,N_2075,N_2903);
nand U4414 (N_4414,N_1846,N_1974);
nand U4415 (N_4415,N_2885,N_2185);
and U4416 (N_4416,N_2823,N_2676);
and U4417 (N_4417,N_2178,N_1869);
nand U4418 (N_4418,N_2382,N_2774);
and U4419 (N_4419,N_1874,N_2642);
and U4420 (N_4420,N_1701,N_2859);
or U4421 (N_4421,N_1714,N_1888);
and U4422 (N_4422,N_2064,N_2976);
nand U4423 (N_4423,N_1698,N_2987);
xnor U4424 (N_4424,N_2942,N_2241);
xnor U4425 (N_4425,N_1809,N_2318);
xnor U4426 (N_4426,N_2957,N_2524);
nand U4427 (N_4427,N_2157,N_2069);
nor U4428 (N_4428,N_2674,N_2225);
nor U4429 (N_4429,N_2826,N_2709);
nand U4430 (N_4430,N_2104,N_2235);
nor U4431 (N_4431,N_2335,N_1613);
or U4432 (N_4432,N_2788,N_2337);
nand U4433 (N_4433,N_2190,N_2636);
or U4434 (N_4434,N_2808,N_2138);
nand U4435 (N_4435,N_2389,N_1659);
xnor U4436 (N_4436,N_2249,N_2586);
and U4437 (N_4437,N_2849,N_2439);
and U4438 (N_4438,N_1963,N_2598);
nor U4439 (N_4439,N_1957,N_1717);
and U4440 (N_4440,N_1669,N_2645);
xnor U4441 (N_4441,N_2017,N_2500);
or U4442 (N_4442,N_2983,N_2065);
nand U4443 (N_4443,N_2972,N_2015);
and U4444 (N_4444,N_2409,N_2547);
nor U4445 (N_4445,N_2237,N_1636);
nand U4446 (N_4446,N_2424,N_2324);
xnor U4447 (N_4447,N_1538,N_1565);
and U4448 (N_4448,N_1791,N_1870);
nand U4449 (N_4449,N_2630,N_1531);
nor U4450 (N_4450,N_2975,N_2452);
and U4451 (N_4451,N_1762,N_2482);
or U4452 (N_4452,N_1871,N_2549);
and U4453 (N_4453,N_2687,N_1572);
nand U4454 (N_4454,N_1520,N_2735);
or U4455 (N_4455,N_2678,N_1959);
or U4456 (N_4456,N_2211,N_2041);
xnor U4457 (N_4457,N_2967,N_2497);
or U4458 (N_4458,N_1630,N_1540);
and U4459 (N_4459,N_2902,N_2782);
xnor U4460 (N_4460,N_2776,N_1959);
xor U4461 (N_4461,N_2162,N_2026);
nor U4462 (N_4462,N_2986,N_2245);
and U4463 (N_4463,N_1814,N_2640);
or U4464 (N_4464,N_2031,N_2507);
xor U4465 (N_4465,N_2251,N_2888);
or U4466 (N_4466,N_2607,N_2506);
xor U4467 (N_4467,N_1608,N_2530);
xor U4468 (N_4468,N_2219,N_2614);
and U4469 (N_4469,N_1723,N_2595);
nand U4470 (N_4470,N_1632,N_2604);
and U4471 (N_4471,N_2109,N_2729);
and U4472 (N_4472,N_2305,N_1526);
and U4473 (N_4473,N_2689,N_1848);
nor U4474 (N_4474,N_2804,N_2772);
nand U4475 (N_4475,N_1599,N_2827);
or U4476 (N_4476,N_1888,N_2167);
xnor U4477 (N_4477,N_1591,N_2633);
xor U4478 (N_4478,N_2664,N_1914);
xnor U4479 (N_4479,N_2185,N_2617);
or U4480 (N_4480,N_1837,N_1571);
nor U4481 (N_4481,N_2317,N_2336);
nor U4482 (N_4482,N_2208,N_2164);
and U4483 (N_4483,N_2564,N_1680);
nand U4484 (N_4484,N_1799,N_2244);
or U4485 (N_4485,N_1866,N_2619);
xor U4486 (N_4486,N_2994,N_2047);
nor U4487 (N_4487,N_1542,N_2296);
nand U4488 (N_4488,N_1798,N_1879);
and U4489 (N_4489,N_2431,N_2679);
nor U4490 (N_4490,N_2267,N_2088);
nand U4491 (N_4491,N_2890,N_1501);
xnor U4492 (N_4492,N_2022,N_2750);
nand U4493 (N_4493,N_1887,N_2128);
xor U4494 (N_4494,N_1694,N_2122);
nor U4495 (N_4495,N_2919,N_2945);
nor U4496 (N_4496,N_1785,N_2108);
nor U4497 (N_4497,N_2780,N_2034);
xnor U4498 (N_4498,N_1642,N_2311);
nand U4499 (N_4499,N_2580,N_1785);
or U4500 (N_4500,N_3718,N_3847);
or U4501 (N_4501,N_4464,N_3835);
xor U4502 (N_4502,N_3923,N_3999);
nand U4503 (N_4503,N_3065,N_3230);
and U4504 (N_4504,N_4162,N_4133);
or U4505 (N_4505,N_3788,N_4434);
or U4506 (N_4506,N_4174,N_3586);
or U4507 (N_4507,N_3077,N_4123);
or U4508 (N_4508,N_3031,N_4167);
nand U4509 (N_4509,N_4176,N_3855);
nor U4510 (N_4510,N_3531,N_4299);
nand U4511 (N_4511,N_3188,N_3389);
and U4512 (N_4512,N_3904,N_3454);
nand U4513 (N_4513,N_3189,N_4352);
and U4514 (N_4514,N_4189,N_4110);
xor U4515 (N_4515,N_3623,N_3499);
nand U4516 (N_4516,N_4365,N_3351);
and U4517 (N_4517,N_3288,N_3284);
and U4518 (N_4518,N_3975,N_3983);
xor U4519 (N_4519,N_3332,N_3916);
nor U4520 (N_4520,N_4276,N_3674);
and U4521 (N_4521,N_4079,N_3010);
or U4522 (N_4522,N_4171,N_3604);
or U4523 (N_4523,N_3627,N_3142);
or U4524 (N_4524,N_3930,N_3283);
or U4525 (N_4525,N_3812,N_4437);
nand U4526 (N_4526,N_3785,N_3101);
nor U4527 (N_4527,N_4408,N_4168);
nand U4528 (N_4528,N_3607,N_4487);
nor U4529 (N_4529,N_3967,N_3509);
and U4530 (N_4530,N_3908,N_4127);
xnor U4531 (N_4531,N_3068,N_3996);
and U4532 (N_4532,N_3701,N_3635);
and U4533 (N_4533,N_3472,N_4083);
and U4534 (N_4534,N_3676,N_3338);
nor U4535 (N_4535,N_4204,N_3191);
xnor U4536 (N_4536,N_4294,N_3337);
nand U4537 (N_4537,N_3845,N_4052);
nor U4538 (N_4538,N_3544,N_3846);
xor U4539 (N_4539,N_3715,N_3605);
and U4540 (N_4540,N_3662,N_3998);
and U4541 (N_4541,N_4423,N_3979);
xor U4542 (N_4542,N_3315,N_3504);
or U4543 (N_4543,N_4376,N_3938);
and U4544 (N_4544,N_3181,N_4497);
nand U4545 (N_4545,N_3083,N_4484);
nor U4546 (N_4546,N_3682,N_4111);
and U4547 (N_4547,N_3611,N_4337);
or U4548 (N_4548,N_3932,N_3954);
or U4549 (N_4549,N_3046,N_3969);
xnor U4550 (N_4550,N_4067,N_3203);
xnor U4551 (N_4551,N_3539,N_4201);
and U4552 (N_4552,N_3208,N_3141);
and U4553 (N_4553,N_4438,N_3327);
and U4554 (N_4554,N_3574,N_3167);
xnor U4555 (N_4555,N_3244,N_3296);
nor U4556 (N_4556,N_3583,N_3480);
nand U4557 (N_4557,N_3392,N_4192);
xor U4558 (N_4558,N_3970,N_3778);
and U4559 (N_4559,N_3793,N_3640);
or U4560 (N_4560,N_3311,N_3196);
nor U4561 (N_4561,N_3724,N_3849);
nor U4562 (N_4562,N_3395,N_3433);
nand U4563 (N_4563,N_4030,N_3872);
nor U4564 (N_4564,N_3731,N_4141);
or U4565 (N_4565,N_3949,N_4129);
or U4566 (N_4566,N_3575,N_3224);
nor U4567 (N_4567,N_3385,N_4452);
and U4568 (N_4568,N_3685,N_3494);
xor U4569 (N_4569,N_4314,N_4406);
or U4570 (N_4570,N_4125,N_4471);
or U4571 (N_4571,N_4383,N_3099);
nand U4572 (N_4572,N_4463,N_3442);
or U4573 (N_4573,N_4293,N_3707);
xnor U4574 (N_4574,N_4004,N_3261);
nand U4575 (N_4575,N_3383,N_3056);
nor U4576 (N_4576,N_4009,N_3787);
nor U4577 (N_4577,N_4350,N_4336);
and U4578 (N_4578,N_3100,N_3647);
xor U4579 (N_4579,N_3137,N_4298);
nand U4580 (N_4580,N_4234,N_3738);
or U4581 (N_4581,N_3824,N_4287);
xor U4582 (N_4582,N_4218,N_3760);
and U4583 (N_4583,N_3255,N_4451);
xor U4584 (N_4584,N_3764,N_3781);
xnor U4585 (N_4585,N_3741,N_3800);
nand U4586 (N_4586,N_4026,N_4065);
and U4587 (N_4587,N_3393,N_3609);
or U4588 (N_4588,N_4394,N_3613);
nand U4589 (N_4589,N_3811,N_3792);
nand U4590 (N_4590,N_3834,N_3709);
nand U4591 (N_4591,N_4388,N_3844);
xnor U4592 (N_4592,N_4245,N_4428);
and U4593 (N_4593,N_3508,N_3298);
xnor U4594 (N_4594,N_3696,N_3522);
nand U4595 (N_4595,N_4296,N_3915);
nor U4596 (N_4596,N_3773,N_4309);
and U4597 (N_4597,N_3020,N_3153);
xor U4598 (N_4598,N_4242,N_3643);
or U4599 (N_4599,N_4040,N_3677);
xor U4600 (N_4600,N_3132,N_3269);
nand U4601 (N_4601,N_3201,N_3403);
xor U4602 (N_4602,N_4163,N_3743);
nor U4603 (N_4603,N_3394,N_3352);
and U4604 (N_4604,N_3889,N_3532);
and U4605 (N_4605,N_3551,N_3193);
or U4606 (N_4606,N_3219,N_3946);
nand U4607 (N_4607,N_3270,N_3651);
nand U4608 (N_4608,N_4013,N_4165);
xor U4609 (N_4609,N_4116,N_3815);
nor U4610 (N_4610,N_4332,N_3036);
or U4611 (N_4611,N_3645,N_3873);
nor U4612 (N_4612,N_3693,N_3429);
nand U4613 (N_4613,N_3919,N_4285);
nand U4614 (N_4614,N_3276,N_3626);
nand U4615 (N_4615,N_3728,N_3683);
or U4616 (N_4616,N_3450,N_3059);
and U4617 (N_4617,N_3250,N_3665);
xor U4618 (N_4618,N_4033,N_4448);
and U4619 (N_4619,N_3906,N_3826);
and U4620 (N_4620,N_3152,N_3241);
and U4621 (N_4621,N_3816,N_4445);
nand U4622 (N_4622,N_3408,N_4290);
xor U4623 (N_4623,N_4048,N_4098);
or U4624 (N_4624,N_3285,N_4476);
nand U4625 (N_4625,N_3636,N_3940);
nand U4626 (N_4626,N_4202,N_3516);
or U4627 (N_4627,N_3777,N_3094);
nor U4628 (N_4628,N_4372,N_3652);
nor U4629 (N_4629,N_4334,N_3076);
or U4630 (N_4630,N_3837,N_3624);
and U4631 (N_4631,N_3328,N_3529);
nor U4632 (N_4632,N_3121,N_3038);
nor U4633 (N_4633,N_3519,N_3015);
nor U4634 (N_4634,N_3356,N_4459);
nand U4635 (N_4635,N_3014,N_3466);
or U4636 (N_4636,N_4398,N_3373);
or U4637 (N_4637,N_3972,N_4301);
or U4638 (N_4638,N_3510,N_4144);
or U4639 (N_4639,N_3411,N_4082);
nand U4640 (N_4640,N_3251,N_3390);
or U4641 (N_4641,N_3857,N_3007);
or U4642 (N_4642,N_3440,N_3012);
xor U4643 (N_4643,N_4235,N_3671);
or U4644 (N_4644,N_3354,N_3111);
and U4645 (N_4645,N_3037,N_3123);
xor U4646 (N_4646,N_3618,N_3143);
xnor U4647 (N_4647,N_3415,N_3317);
nand U4648 (N_4648,N_3122,N_3286);
xnor U4649 (N_4649,N_4231,N_4000);
nor U4650 (N_4650,N_3089,N_4243);
nor U4651 (N_4651,N_3981,N_3673);
nor U4652 (N_4652,N_4327,N_3183);
or U4653 (N_4653,N_4213,N_3880);
or U4654 (N_4654,N_3971,N_3937);
nand U4655 (N_4655,N_3515,N_3309);
nand U4656 (N_4656,N_4489,N_3874);
or U4657 (N_4657,N_4279,N_3488);
xor U4658 (N_4658,N_3161,N_4090);
or U4659 (N_4659,N_3573,N_4330);
nand U4660 (N_4660,N_3560,N_3348);
xnor U4661 (N_4661,N_4099,N_3506);
and U4662 (N_4662,N_3882,N_4077);
nand U4663 (N_4663,N_3173,N_4232);
nand U4664 (N_4664,N_4429,N_4343);
or U4665 (N_4665,N_3610,N_4321);
nand U4666 (N_4666,N_3911,N_3799);
nor U4667 (N_4667,N_3747,N_3144);
and U4668 (N_4668,N_4379,N_3710);
or U4669 (N_4669,N_3482,N_4399);
and U4670 (N_4670,N_4105,N_3150);
nand U4671 (N_4671,N_3939,N_3303);
or U4672 (N_4672,N_3236,N_4087);
or U4673 (N_4673,N_3655,N_3853);
and U4674 (N_4674,N_3871,N_3809);
or U4675 (N_4675,N_3806,N_3469);
xnor U4676 (N_4676,N_4302,N_3865);
nand U4677 (N_4677,N_3424,N_3737);
nand U4678 (N_4678,N_3216,N_3293);
or U4679 (N_4679,N_3115,N_3905);
or U4680 (N_4680,N_4166,N_3430);
or U4681 (N_4681,N_3473,N_3331);
or U4682 (N_4682,N_3520,N_3186);
and U4683 (N_4683,N_3571,N_3320);
and U4684 (N_4684,N_3124,N_4233);
nand U4685 (N_4685,N_3767,N_3190);
xnor U4686 (N_4686,N_4173,N_3098);
nor U4687 (N_4687,N_4430,N_4016);
nand U4688 (N_4688,N_3514,N_3563);
xnor U4689 (N_4689,N_4253,N_4361);
nor U4690 (N_4690,N_3802,N_3814);
nor U4691 (N_4691,N_3714,N_3085);
nand U4692 (N_4692,N_4441,N_3592);
and U4693 (N_4693,N_4465,N_4136);
xor U4694 (N_4694,N_3585,N_4325);
nand U4695 (N_4695,N_4342,N_4022);
nand U4696 (N_4696,N_3438,N_4442);
nor U4697 (N_4697,N_4057,N_3187);
nand U4698 (N_4698,N_3796,N_4023);
or U4699 (N_4699,N_3368,N_3172);
or U4700 (N_4700,N_3692,N_3663);
nor U4701 (N_4701,N_3176,N_3698);
or U4702 (N_4702,N_4300,N_3476);
xor U4703 (N_4703,N_3289,N_4102);
or U4704 (N_4704,N_3040,N_3061);
xor U4705 (N_4705,N_3165,N_3256);
or U4706 (N_4706,N_3989,N_3479);
nor U4707 (N_4707,N_4366,N_4260);
nor U4708 (N_4708,N_4240,N_3088);
xor U4709 (N_4709,N_3263,N_3615);
nand U4710 (N_4710,N_3689,N_3774);
and U4711 (N_4711,N_4095,N_4074);
and U4712 (N_4712,N_4130,N_4313);
xor U4713 (N_4713,N_3436,N_3029);
xor U4714 (N_4714,N_4209,N_4108);
or U4715 (N_4715,N_3481,N_3599);
nor U4716 (N_4716,N_4432,N_4122);
nand U4717 (N_4717,N_3060,N_4289);
and U4718 (N_4718,N_3159,N_3326);
nand U4719 (N_4719,N_3246,N_3541);
nor U4720 (N_4720,N_3247,N_4024);
nor U4721 (N_4721,N_3723,N_3362);
and U4722 (N_4722,N_4206,N_3420);
and U4723 (N_4723,N_3112,N_3725);
and U4724 (N_4724,N_3034,N_3726);
nor U4725 (N_4725,N_3895,N_4257);
or U4726 (N_4726,N_3017,N_3071);
and U4727 (N_4727,N_3470,N_4303);
or U4728 (N_4728,N_4272,N_3517);
xor U4729 (N_4729,N_4094,N_3217);
nand U4730 (N_4730,N_4247,N_3266);
and U4731 (N_4731,N_3681,N_4075);
nor U4732 (N_4732,N_3067,N_3678);
xor U4733 (N_4733,N_3232,N_3295);
xor U4734 (N_4734,N_3924,N_4207);
or U4735 (N_4735,N_4416,N_3242);
nor U4736 (N_4736,N_3075,N_4138);
or U4737 (N_4737,N_3058,N_3307);
or U4738 (N_4738,N_3210,N_3513);
xnor U4739 (N_4739,N_4373,N_3090);
nor U4740 (N_4740,N_3739,N_3818);
and U4741 (N_4741,N_3943,N_3850);
nor U4742 (N_4742,N_3866,N_4374);
and U4743 (N_4743,N_4146,N_3062);
nor U4744 (N_4744,N_3301,N_3754);
nand U4745 (N_4745,N_3490,N_4409);
nor U4746 (N_4746,N_4252,N_3021);
nand U4747 (N_4747,N_3340,N_3898);
xor U4748 (N_4748,N_4046,N_3547);
xor U4749 (N_4749,N_3486,N_3556);
and U4750 (N_4750,N_3237,N_3982);
nand U4751 (N_4751,N_4080,N_3661);
and U4752 (N_4752,N_3598,N_3041);
and U4753 (N_4753,N_3658,N_3893);
nand U4754 (N_4754,N_3576,N_4284);
nand U4755 (N_4755,N_3033,N_4045);
or U4756 (N_4756,N_3002,N_3366);
or U4757 (N_4757,N_3157,N_4205);
nor U4758 (N_4758,N_3282,N_3192);
xor U4759 (N_4759,N_3903,N_3310);
nand U4760 (N_4760,N_4324,N_3458);
or U4761 (N_4761,N_3240,N_3521);
nand U4762 (N_4762,N_4368,N_4469);
nand U4763 (N_4763,N_3776,N_3711);
and U4764 (N_4764,N_3164,N_4227);
nor U4765 (N_4765,N_3084,N_4224);
nor U4766 (N_4766,N_3997,N_3942);
nor U4767 (N_4767,N_4344,N_3974);
nor U4768 (N_4768,N_4482,N_4404);
nand U4769 (N_4769,N_4104,N_3406);
nand U4770 (N_4770,N_3955,N_3823);
nand U4771 (N_4771,N_4073,N_3732);
or U4772 (N_4772,N_3195,N_3933);
nor U4773 (N_4773,N_3103,N_3439);
nor U4774 (N_4774,N_3091,N_3434);
xnor U4775 (N_4775,N_3006,N_3491);
or U4776 (N_4776,N_3578,N_4028);
xor U4777 (N_4777,N_3018,N_4160);
and U4778 (N_4778,N_3452,N_3670);
or U4779 (N_4779,N_3158,N_4086);
xor U4780 (N_4780,N_3238,N_3957);
nor U4781 (N_4781,N_3446,N_4049);
nand U4782 (N_4782,N_3225,N_3281);
nor U4783 (N_4783,N_3786,N_3253);
nor U4784 (N_4784,N_3134,N_3708);
nand U4785 (N_4785,N_4228,N_3211);
or U4786 (N_4786,N_3881,N_3736);
or U4787 (N_4787,N_4262,N_4119);
nor U4788 (N_4788,N_3876,N_3330);
xor U4789 (N_4789,N_3047,N_3043);
nand U4790 (N_4790,N_3966,N_3465);
nor U4791 (N_4791,N_3218,N_3220);
nand U4792 (N_4792,N_4450,N_4066);
nor U4793 (N_4793,N_3909,N_3222);
nor U4794 (N_4794,N_3028,N_3024);
and U4795 (N_4795,N_3080,N_4084);
nor U4796 (N_4796,N_4397,N_3428);
and U4797 (N_4797,N_3110,N_3536);
and U4798 (N_4798,N_3254,N_4270);
nand U4799 (N_4799,N_4217,N_4357);
nor U4800 (N_4800,N_3593,N_4191);
or U4801 (N_4801,N_3603,N_3935);
and U4802 (N_4802,N_3313,N_4003);
or U4803 (N_4803,N_3496,N_3695);
nand U4804 (N_4804,N_4107,N_3422);
nor U4805 (N_4805,N_3988,N_3595);
or U4806 (N_4806,N_4269,N_4051);
and U4807 (N_4807,N_3455,N_4059);
nor U4808 (N_4808,N_3730,N_4153);
and U4809 (N_4809,N_3828,N_3412);
xnor U4810 (N_4810,N_3052,N_4490);
or U4811 (N_4811,N_3780,N_3746);
xor U4812 (N_4812,N_3782,N_4312);
or U4813 (N_4813,N_4387,N_3808);
or U4814 (N_4814,N_3562,N_4170);
xnor U4815 (N_4815,N_4216,N_3474);
nand U4816 (N_4816,N_3401,N_3435);
and U4817 (N_4817,N_3807,N_4367);
or U4818 (N_4818,N_3334,N_3171);
nor U4819 (N_4819,N_3827,N_3464);
and U4820 (N_4820,N_3205,N_3622);
and U4821 (N_4821,N_3092,N_3821);
or U4822 (N_4822,N_3441,N_4055);
nor U4823 (N_4823,N_3264,N_4076);
nor U4824 (N_4824,N_3257,N_3267);
xor U4825 (N_4825,N_3820,N_4044);
nor U4826 (N_4826,N_3891,N_4011);
and U4827 (N_4827,N_3180,N_4317);
nand U4828 (N_4828,N_4188,N_4422);
xor U4829 (N_4829,N_3910,N_3104);
xnor U4830 (N_4830,N_3934,N_3045);
xor U4831 (N_4831,N_3892,N_3883);
xor U4832 (N_4832,N_4197,N_3249);
xor U4833 (N_4833,N_3596,N_3680);
nor U4834 (N_4834,N_4225,N_4185);
xnor U4835 (N_4835,N_3527,N_3492);
or U4836 (N_4836,N_4280,N_3762);
nor U4837 (N_4837,N_3960,N_4395);
xnor U4838 (N_4838,N_3497,N_3750);
or U4839 (N_4839,N_4151,N_3928);
or U4840 (N_4840,N_3659,N_3748);
nor U4841 (N_4841,N_3437,N_3641);
nand U4842 (N_4842,N_4058,N_3638);
or U4843 (N_4843,N_4433,N_4392);
nand U4844 (N_4844,N_4311,N_4060);
xor U4845 (N_4845,N_3962,N_4156);
and U4846 (N_4846,N_3292,N_3105);
nand U4847 (N_4847,N_4021,N_3489);
xor U4848 (N_4848,N_3869,N_4346);
nand U4849 (N_4849,N_3794,N_3477);
nand U4850 (N_4850,N_3961,N_3859);
nand U4851 (N_4851,N_4050,N_3319);
and U4852 (N_4852,N_4483,N_3400);
nand U4853 (N_4853,N_3557,N_3601);
nor U4854 (N_4854,N_4412,N_3644);
xnor U4855 (N_4855,N_3361,N_3372);
nor U4856 (N_4856,N_3064,N_3637);
and U4857 (N_4857,N_4472,N_3279);
nand U4858 (N_4858,N_3130,N_3565);
nand U4859 (N_4859,N_3765,N_3300);
or U4860 (N_4860,N_4158,N_3215);
or U4861 (N_4861,N_3117,N_4458);
and U4862 (N_4862,N_3810,N_4488);
xnor U4863 (N_4863,N_3822,N_3550);
nand U4864 (N_4864,N_4027,N_3375);
nand U4865 (N_4865,N_4477,N_3380);
xnor U4866 (N_4866,N_3177,N_4249);
xor U4867 (N_4867,N_3213,N_3913);
and U4868 (N_4868,N_4275,N_3761);
or U4869 (N_4869,N_3417,N_3475);
nand U4870 (N_4870,N_3081,N_3646);
or U4871 (N_4871,N_3174,N_4149);
nand U4872 (N_4872,N_3146,N_3170);
nand U4873 (N_4873,N_3798,N_4386);
nor U4874 (N_4874,N_4440,N_4467);
xor U4875 (N_4875,N_3931,N_4281);
nor U4876 (N_4876,N_3397,N_3066);
or U4877 (N_4877,N_3323,N_3095);
nand U4878 (N_4878,N_3617,N_3032);
and U4879 (N_4879,N_3302,N_4268);
nand U4880 (N_4880,N_4172,N_3022);
nand U4881 (N_4881,N_4186,N_3591);
and U4882 (N_4882,N_4499,N_4389);
xor U4883 (N_4883,N_3369,N_3048);
nand U4884 (N_4884,N_3291,N_3227);
xor U4885 (N_4885,N_3921,N_3569);
or U4886 (N_4886,N_3752,N_3495);
or U4887 (N_4887,N_3287,N_4359);
nand U4888 (N_4888,N_4179,N_4425);
nor U4889 (N_4889,N_3070,N_4431);
xnor U4890 (N_4890,N_4401,N_3306);
nor U4891 (N_4891,N_4152,N_3443);
and U4892 (N_4892,N_3003,N_4328);
nand U4893 (N_4893,N_3462,N_3936);
and U4894 (N_4894,N_3280,N_3779);
and U4895 (N_4895,N_3318,N_4148);
nand U4896 (N_4896,N_4297,N_3484);
nand U4897 (N_4897,N_3890,N_4345);
nor U4898 (N_4898,N_4274,N_4005);
xor U4899 (N_4899,N_4203,N_4193);
and U4900 (N_4900,N_3852,N_4335);
nor U4901 (N_4901,N_3233,N_4208);
nor U4902 (N_4902,N_4042,N_3648);
or U4903 (N_4903,N_3344,N_3457);
xnor U4904 (N_4904,N_3290,N_4447);
nand U4905 (N_4905,N_3713,N_3907);
nand U4906 (N_4906,N_4029,N_3019);
nor U4907 (N_4907,N_3538,N_3135);
nand U4908 (N_4908,N_3483,N_4147);
nor U4909 (N_4909,N_3087,N_3376);
and U4910 (N_4910,N_3096,N_4363);
or U4911 (N_4911,N_3769,N_3775);
nor U4912 (N_4912,N_4126,N_3580);
or U4913 (N_4913,N_3699,N_4143);
xnor U4914 (N_4914,N_4391,N_3456);
xor U4915 (N_4915,N_3353,N_4237);
or U4916 (N_4916,N_3262,N_3705);
nor U4917 (N_4917,N_3228,N_3831);
nor U4918 (N_4918,N_3004,N_4093);
nand U4919 (N_4919,N_4256,N_3404);
or U4920 (N_4920,N_3642,N_3448);
xnor U4921 (N_4921,N_3026,N_3825);
nor U4922 (N_4922,N_3629,N_3941);
or U4923 (N_4923,N_4053,N_4474);
xnor U4924 (N_4924,N_3063,N_3168);
or U4925 (N_4925,N_4455,N_3757);
nand U4926 (N_4926,N_3606,N_4113);
or U4927 (N_4927,N_4360,N_4351);
xnor U4928 (N_4928,N_3977,N_3675);
or U4929 (N_4929,N_4085,N_3667);
or U4930 (N_4930,N_3343,N_3133);
and U4931 (N_4931,N_3719,N_3740);
xor U4932 (N_4932,N_3964,N_3860);
and U4933 (N_4933,N_3386,N_3023);
or U4934 (N_4934,N_3097,N_3733);
and U4935 (N_4935,N_4427,N_4498);
or U4936 (N_4936,N_3868,N_3929);
and U4937 (N_4937,N_3425,N_3803);
nor U4938 (N_4938,N_3734,N_3973);
nand U4939 (N_4939,N_3453,N_4064);
and U4940 (N_4940,N_3727,N_3314);
and U4941 (N_4941,N_4068,N_3407);
nor U4942 (N_4942,N_3324,N_3347);
or U4943 (N_4943,N_4316,N_3468);
and U4944 (N_4944,N_3114,N_3577);
or U4945 (N_4945,N_4362,N_3273);
xnor U4946 (N_4946,N_3008,N_3387);
and U4947 (N_4947,N_3268,N_3836);
and U4948 (N_4948,N_4037,N_4400);
and U4949 (N_4949,N_3630,N_3182);
and U4950 (N_4950,N_4385,N_4196);
nand U4951 (N_4951,N_3588,N_3856);
nor U4952 (N_4952,N_3487,N_4140);
or U4953 (N_4953,N_3772,N_3235);
nor U4954 (N_4954,N_3325,N_3952);
and U4955 (N_4955,N_4056,N_3633);
nor U4956 (N_4956,N_3953,N_3399);
or U4957 (N_4957,N_4453,N_3763);
xor U4958 (N_4958,N_3357,N_3621);
nand U4959 (N_4959,N_3505,N_3951);
nor U4960 (N_4960,N_3149,N_3669);
and U4961 (N_4961,N_3756,N_3418);
or U4962 (N_4962,N_3523,N_4380);
nor U4963 (N_4963,N_3140,N_3231);
nand U4964 (N_4964,N_3833,N_4306);
nand U4965 (N_4965,N_3947,N_3365);
and U4966 (N_4966,N_4286,N_4230);
and U4967 (N_4967,N_3234,N_3278);
nor U4968 (N_4968,N_4415,N_3546);
and U4969 (N_4969,N_3958,N_4112);
nor U4970 (N_4970,N_3414,N_4492);
and U4971 (N_4971,N_4012,N_3316);
nor U4972 (N_4972,N_4019,N_3275);
and U4973 (N_4973,N_3572,N_4248);
or U4974 (N_4974,N_4263,N_3795);
or U4975 (N_4975,N_3447,N_4277);
nand U4976 (N_4976,N_3650,N_4106);
nor U4977 (N_4977,N_3185,N_3363);
and U4978 (N_4978,N_3867,N_4264);
nor U4979 (N_4979,N_3841,N_3305);
nand U4980 (N_4980,N_3700,N_4323);
nor U4981 (N_4981,N_3398,N_3129);
and U4982 (N_4982,N_3691,N_4419);
xnor U4983 (N_4983,N_4114,N_3877);
nand U4984 (N_4984,N_3154,N_3771);
xor U4985 (N_4985,N_3248,N_4475);
nor U4986 (N_4986,N_4241,N_3925);
xnor U4987 (N_4987,N_3570,N_3207);
nor U4988 (N_4988,N_4396,N_3136);
nand U4989 (N_4989,N_3843,N_3742);
and U4990 (N_4990,N_4246,N_4480);
nor U4991 (N_4991,N_4061,N_3634);
and U4992 (N_4992,N_4155,N_4182);
xnor U4993 (N_4993,N_4364,N_3703);
or U4994 (N_4994,N_3206,N_3993);
or U4995 (N_4995,N_3223,N_3978);
or U4996 (N_4996,N_3959,N_3870);
xor U4997 (N_4997,N_3759,N_3374);
nor U4998 (N_4998,N_3148,N_3920);
nand U4999 (N_4999,N_3566,N_3553);
nor U5000 (N_5000,N_3801,N_3963);
and U5001 (N_5001,N_3864,N_3156);
and U5002 (N_5002,N_3359,N_4039);
xnor U5003 (N_5003,N_4142,N_3459);
xnor U5004 (N_5004,N_4215,N_3590);
nor U5005 (N_5005,N_4353,N_4486);
xor U5006 (N_5006,N_3042,N_3832);
nand U5007 (N_5007,N_4025,N_3886);
xnor U5008 (N_5008,N_3976,N_3013);
and U5009 (N_5009,N_3649,N_4134);
or U5010 (N_5010,N_4417,N_3545);
nand U5011 (N_5011,N_3057,N_3405);
xor U5012 (N_5012,N_3770,N_4238);
xor U5013 (N_5013,N_3030,N_4071);
nand U5014 (N_5014,N_3579,N_3884);
xor U5015 (N_5015,N_3914,N_3639);
xnor U5016 (N_5016,N_4444,N_3887);
or U5017 (N_5017,N_3118,N_3897);
nor U5018 (N_5018,N_3355,N_4007);
xor U5019 (N_5019,N_3199,N_3339);
nand U5020 (N_5020,N_3745,N_3126);
or U5021 (N_5021,N_3533,N_3688);
nand U5022 (N_5022,N_3768,N_3568);
nand U5023 (N_5023,N_4347,N_3530);
xor U5024 (N_5024,N_3367,N_4457);
xor U5025 (N_5025,N_3653,N_3819);
or U5026 (N_5026,N_3668,N_3848);
xor U5027 (N_5027,N_3402,N_3053);
nor U5028 (N_5028,N_3956,N_4340);
nor U5029 (N_5029,N_3986,N_3106);
nand U5030 (N_5030,N_3830,N_4115);
xor U5031 (N_5031,N_4069,N_3702);
xnor U5032 (N_5032,N_3888,N_3214);
nand U5033 (N_5033,N_3790,N_3184);
or U5034 (N_5034,N_3069,N_3512);
xnor U5035 (N_5035,N_3861,N_4255);
xor U5036 (N_5036,N_4020,N_3086);
and U5037 (N_5037,N_4435,N_4456);
and U5038 (N_5038,N_3755,N_3277);
nand U5039 (N_5039,N_3044,N_4091);
nand U5040 (N_5040,N_3965,N_3984);
or U5041 (N_5041,N_4015,N_3243);
nand U5042 (N_5042,N_3471,N_3994);
xnor U5043 (N_5043,N_3107,N_3239);
or U5044 (N_5044,N_3697,N_3011);
xor U5045 (N_5045,N_3660,N_4118);
xnor U5046 (N_5046,N_3274,N_4222);
nand U5047 (N_5047,N_3335,N_3346);
xor U5048 (N_5048,N_4305,N_3602);
nand U5049 (N_5049,N_3444,N_3524);
or U5050 (N_5050,N_4032,N_4239);
or U5051 (N_5051,N_4390,N_3178);
and U5052 (N_5052,N_3294,N_4333);
xor U5053 (N_5053,N_3322,N_4410);
and U5054 (N_5054,N_3054,N_3501);
or U5055 (N_5055,N_4031,N_3147);
and U5056 (N_5056,N_3783,N_3500);
and U5057 (N_5057,N_3345,N_3619);
xor U5058 (N_5058,N_4063,N_4291);
nand U5059 (N_5059,N_3535,N_3628);
and U5060 (N_5060,N_3463,N_4411);
and U5061 (N_5061,N_3050,N_3991);
xor U5062 (N_5062,N_3005,N_4322);
or U5063 (N_5063,N_3537,N_4449);
and U5064 (N_5064,N_3534,N_3297);
and U5065 (N_5065,N_4101,N_3507);
nand U5066 (N_5066,N_4132,N_4088);
or U5067 (N_5067,N_4288,N_4041);
xnor U5068 (N_5068,N_4375,N_4405);
xor U5069 (N_5069,N_3840,N_4078);
nor U5070 (N_5070,N_3016,N_4219);
nand U5071 (N_5071,N_4103,N_3001);
xor U5072 (N_5072,N_3364,N_3612);
and U5073 (N_5073,N_3431,N_3687);
xor U5074 (N_5074,N_4154,N_3093);
nand U5075 (N_5075,N_3116,N_4493);
nand U5076 (N_5076,N_3885,N_3555);
nand U5077 (N_5077,N_4421,N_4251);
and U5078 (N_5078,N_3427,N_4164);
and U5079 (N_5079,N_3039,N_3049);
and U5080 (N_5080,N_3329,N_3654);
xnor U5081 (N_5081,N_3051,N_3567);
xnor U5082 (N_5082,N_3944,N_3554);
xor U5083 (N_5083,N_3616,N_3035);
or U5084 (N_5084,N_4035,N_3922);
xor U5085 (N_5085,N_3614,N_4377);
xnor U5086 (N_5086,N_4008,N_3055);
xor U5087 (N_5087,N_3419,N_4338);
or U5088 (N_5088,N_3179,N_3252);
and U5089 (N_5089,N_3525,N_3901);
nor U5090 (N_5090,N_3721,N_4295);
or U5091 (N_5091,N_4308,N_4393);
nor U5092 (N_5092,N_3594,N_4047);
and U5093 (N_5093,N_3766,N_4348);
nor U5094 (N_5094,N_4354,N_3502);
nand U5095 (N_5095,N_4161,N_3461);
nor U5096 (N_5096,N_4292,N_4036);
and U5097 (N_5097,N_3912,N_3125);
and U5098 (N_5098,N_4439,N_3917);
nand U5099 (N_5099,N_3899,N_3712);
and U5100 (N_5100,N_4491,N_4339);
and U5101 (N_5101,N_3694,N_4200);
xnor U5102 (N_5102,N_4378,N_3145);
xnor U5103 (N_5103,N_3259,N_4420);
and U5104 (N_5104,N_3162,N_3980);
or U5105 (N_5105,N_4461,N_3072);
nor U5106 (N_5106,N_3258,N_3729);
nand U5107 (N_5107,N_3265,N_4426);
nand U5108 (N_5108,N_3839,N_3109);
and U5109 (N_5109,N_4265,N_4014);
xor U5110 (N_5110,N_4259,N_4180);
nand U5111 (N_5111,N_3272,N_4214);
and U5112 (N_5112,N_3212,N_3817);
nand U5113 (N_5113,N_3160,N_3838);
xnor U5114 (N_5114,N_4054,N_3460);
xnor U5115 (N_5115,N_4250,N_3226);
and U5116 (N_5116,N_3632,N_3842);
nor U5117 (N_5117,N_3879,N_4244);
xor U5118 (N_5118,N_3758,N_3449);
nor U5119 (N_5119,N_4424,N_4271);
and U5120 (N_5120,N_3379,N_4006);
and U5121 (N_5121,N_3992,N_4436);
nand U5122 (N_5122,N_4034,N_3498);
nor U5123 (N_5123,N_3478,N_3197);
nand U5124 (N_5124,N_4261,N_3175);
nand U5125 (N_5125,N_4307,N_4454);
nand U5126 (N_5126,N_3625,N_4121);
nor U5127 (N_5127,N_3308,N_3558);
or U5128 (N_5128,N_4210,N_3945);
nor U5129 (N_5129,N_3735,N_3608);
or U5130 (N_5130,N_4195,N_4258);
nor U5131 (N_5131,N_4157,N_4462);
nand U5132 (N_5132,N_4169,N_3416);
nand U5133 (N_5133,N_3720,N_3990);
and U5134 (N_5134,N_4199,N_3127);
and U5135 (N_5135,N_4283,N_3410);
nor U5136 (N_5136,N_3716,N_3421);
and U5137 (N_5137,N_3666,N_3209);
nor U5138 (N_5138,N_3078,N_3657);
nor U5139 (N_5139,N_3511,N_4175);
nand U5140 (N_5140,N_3493,N_3025);
nor U5141 (N_5141,N_3467,N_4190);
xnor U5142 (N_5142,N_3894,N_4355);
xnor U5143 (N_5143,N_3995,N_3138);
nand U5144 (N_5144,N_3854,N_4473);
xor U5145 (N_5145,N_4267,N_3350);
nor U5146 (N_5146,N_3009,N_4495);
xnor U5147 (N_5147,N_3968,N_3271);
nand U5148 (N_5148,N_3918,N_3163);
or U5149 (N_5149,N_3552,N_3299);
or U5150 (N_5150,N_3342,N_3672);
nand U5151 (N_5151,N_3749,N_3396);
or U5152 (N_5152,N_3631,N_4131);
nor U5153 (N_5153,N_4273,N_4468);
and U5154 (N_5154,N_3336,N_4331);
and U5155 (N_5155,N_3950,N_3503);
nor U5156 (N_5156,N_3128,N_3027);
xor U5157 (N_5157,N_4254,N_4494);
or U5158 (N_5158,N_3717,N_3900);
nand U5159 (N_5159,N_3528,N_3829);
xor U5160 (N_5160,N_3896,N_3656);
nor U5161 (N_5161,N_4043,N_3858);
and U5162 (N_5162,N_3744,N_3797);
nand U5163 (N_5163,N_3202,N_3597);
and U5164 (N_5164,N_4370,N_4478);
and U5165 (N_5165,N_3391,N_4184);
nor U5166 (N_5166,N_3378,N_4018);
nand U5167 (N_5167,N_3073,N_4181);
nand U5168 (N_5168,N_3321,N_3582);
xnor U5169 (N_5169,N_4326,N_4315);
nor U5170 (N_5170,N_4318,N_4349);
or U5171 (N_5171,N_4120,N_4282);
xnor U5172 (N_5172,N_3079,N_4407);
nor U5173 (N_5173,N_4072,N_3664);
and U5174 (N_5174,N_3863,N_3423);
or U5175 (N_5175,N_3540,N_3198);
and U5176 (N_5176,N_4017,N_3985);
or U5177 (N_5177,N_4414,N_4092);
xor U5178 (N_5178,N_4481,N_3686);
xnor U5179 (N_5179,N_3381,N_3371);
or U5180 (N_5180,N_3722,N_3113);
xor U5181 (N_5181,N_4381,N_4369);
and U5182 (N_5182,N_4226,N_4236);
and U5183 (N_5183,N_4221,N_3102);
xnor U5184 (N_5184,N_4371,N_4183);
nand U5185 (N_5185,N_3987,N_3948);
and U5186 (N_5186,N_4124,N_3119);
nand U5187 (N_5187,N_3409,N_3542);
or U5188 (N_5188,N_3384,N_3451);
and U5189 (N_5189,N_4413,N_3584);
and U5190 (N_5190,N_3108,N_3426);
nand U5191 (N_5191,N_3581,N_3804);
or U5192 (N_5192,N_4402,N_4097);
nor U5193 (N_5193,N_3260,N_3358);
or U5194 (N_5194,N_3564,N_3902);
xnor U5195 (N_5195,N_3155,N_3341);
and U5196 (N_5196,N_4229,N_3166);
xnor U5197 (N_5197,N_3349,N_4496);
or U5198 (N_5198,N_3194,N_3245);
and U5199 (N_5199,N_3518,N_3333);
nand U5200 (N_5200,N_4329,N_3312);
nand U5201 (N_5201,N_3862,N_4211);
and U5202 (N_5202,N_4384,N_4089);
nand U5203 (N_5203,N_4117,N_3485);
nor U5204 (N_5204,N_3791,N_4150);
nor U5205 (N_5205,N_3413,N_3878);
xor U5206 (N_5206,N_3229,N_3388);
and U5207 (N_5207,N_3751,N_4460);
nor U5208 (N_5208,N_4320,N_3600);
and U5209 (N_5209,N_3706,N_3548);
nand U5210 (N_5210,N_3587,N_3526);
nand U5211 (N_5211,N_3927,N_4220);
nand U5212 (N_5212,N_3139,N_4137);
nor U5213 (N_5213,N_3789,N_4341);
nand U5214 (N_5214,N_3559,N_3169);
nor U5215 (N_5215,N_3684,N_3000);
and U5216 (N_5216,N_4178,N_3561);
and U5217 (N_5217,N_4187,N_4479);
or U5218 (N_5218,N_3690,N_3543);
nand U5219 (N_5219,N_3377,N_3151);
and U5220 (N_5220,N_4198,N_3204);
nand U5221 (N_5221,N_3753,N_4109);
or U5222 (N_5222,N_3370,N_4135);
and U5223 (N_5223,N_3221,N_4038);
or U5224 (N_5224,N_3432,N_4356);
nand U5225 (N_5225,N_3926,N_3620);
nand U5226 (N_5226,N_3589,N_3200);
or U5227 (N_5227,N_3784,N_4466);
or U5228 (N_5228,N_4403,N_4177);
and U5229 (N_5229,N_3805,N_4304);
or U5230 (N_5230,N_3704,N_4223);
xnor U5231 (N_5231,N_3120,N_4100);
xor U5232 (N_5232,N_4212,N_3074);
nand U5233 (N_5233,N_4145,N_4358);
and U5234 (N_5234,N_3679,N_3549);
nand U5235 (N_5235,N_4002,N_4266);
nor U5236 (N_5236,N_3813,N_4139);
nor U5237 (N_5237,N_4485,N_3082);
or U5238 (N_5238,N_4070,N_3304);
or U5239 (N_5239,N_4128,N_4062);
and U5240 (N_5240,N_4382,N_3445);
and U5241 (N_5241,N_4319,N_4446);
nor U5242 (N_5242,N_4443,N_3131);
xnor U5243 (N_5243,N_4096,N_4001);
and U5244 (N_5244,N_3851,N_3382);
and U5245 (N_5245,N_3360,N_4470);
nand U5246 (N_5246,N_4010,N_4194);
xor U5247 (N_5247,N_4159,N_4278);
and U5248 (N_5248,N_4081,N_3875);
or U5249 (N_5249,N_4310,N_4418);
nand U5250 (N_5250,N_4069,N_3350);
xor U5251 (N_5251,N_3749,N_4499);
and U5252 (N_5252,N_3134,N_3260);
nand U5253 (N_5253,N_4442,N_3562);
or U5254 (N_5254,N_3257,N_4164);
nand U5255 (N_5255,N_4390,N_3899);
or U5256 (N_5256,N_3606,N_3691);
or U5257 (N_5257,N_3887,N_3087);
nand U5258 (N_5258,N_3127,N_3263);
nor U5259 (N_5259,N_4434,N_3558);
or U5260 (N_5260,N_3004,N_3470);
or U5261 (N_5261,N_3713,N_3993);
and U5262 (N_5262,N_3347,N_3740);
or U5263 (N_5263,N_4067,N_3538);
and U5264 (N_5264,N_4286,N_3048);
xnor U5265 (N_5265,N_4431,N_3254);
or U5266 (N_5266,N_3313,N_4269);
xnor U5267 (N_5267,N_3368,N_4327);
xor U5268 (N_5268,N_3958,N_3130);
xor U5269 (N_5269,N_3790,N_4491);
xnor U5270 (N_5270,N_3130,N_3594);
xnor U5271 (N_5271,N_3785,N_3857);
nor U5272 (N_5272,N_3851,N_3396);
nor U5273 (N_5273,N_3111,N_3705);
xor U5274 (N_5274,N_4367,N_3620);
nand U5275 (N_5275,N_4466,N_4234);
nor U5276 (N_5276,N_4337,N_3503);
and U5277 (N_5277,N_4263,N_3833);
xor U5278 (N_5278,N_4297,N_3758);
and U5279 (N_5279,N_3279,N_3459);
xor U5280 (N_5280,N_3682,N_4113);
xnor U5281 (N_5281,N_3113,N_4318);
and U5282 (N_5282,N_4374,N_4191);
xor U5283 (N_5283,N_3689,N_3039);
xnor U5284 (N_5284,N_4461,N_3064);
xor U5285 (N_5285,N_3879,N_3468);
nand U5286 (N_5286,N_3713,N_4461);
nor U5287 (N_5287,N_3842,N_3476);
or U5288 (N_5288,N_4193,N_3155);
or U5289 (N_5289,N_3622,N_3441);
nor U5290 (N_5290,N_3043,N_4193);
xnor U5291 (N_5291,N_3255,N_3767);
or U5292 (N_5292,N_4206,N_3978);
nand U5293 (N_5293,N_3971,N_3218);
nand U5294 (N_5294,N_4491,N_4154);
or U5295 (N_5295,N_4025,N_3382);
nor U5296 (N_5296,N_4349,N_4143);
and U5297 (N_5297,N_3830,N_3250);
and U5298 (N_5298,N_3010,N_3434);
and U5299 (N_5299,N_4200,N_3984);
xor U5300 (N_5300,N_3290,N_4083);
xor U5301 (N_5301,N_3586,N_3133);
xor U5302 (N_5302,N_3212,N_3652);
or U5303 (N_5303,N_3357,N_3551);
nand U5304 (N_5304,N_4379,N_4276);
and U5305 (N_5305,N_3301,N_4163);
nor U5306 (N_5306,N_3955,N_3805);
or U5307 (N_5307,N_3516,N_4229);
and U5308 (N_5308,N_4028,N_3159);
xnor U5309 (N_5309,N_3204,N_4233);
nor U5310 (N_5310,N_3888,N_4058);
and U5311 (N_5311,N_3226,N_4065);
nor U5312 (N_5312,N_3142,N_4107);
xor U5313 (N_5313,N_3672,N_4066);
and U5314 (N_5314,N_3264,N_3683);
or U5315 (N_5315,N_3298,N_4102);
xnor U5316 (N_5316,N_3685,N_4352);
or U5317 (N_5317,N_3597,N_4351);
nand U5318 (N_5318,N_4037,N_4193);
xor U5319 (N_5319,N_3869,N_3800);
or U5320 (N_5320,N_3024,N_3073);
or U5321 (N_5321,N_3092,N_3190);
nand U5322 (N_5322,N_3167,N_3469);
or U5323 (N_5323,N_3588,N_3938);
nand U5324 (N_5324,N_4089,N_3828);
and U5325 (N_5325,N_3761,N_3178);
nor U5326 (N_5326,N_3357,N_3067);
nor U5327 (N_5327,N_4263,N_3876);
nor U5328 (N_5328,N_4391,N_3504);
and U5329 (N_5329,N_4246,N_3418);
or U5330 (N_5330,N_3925,N_3540);
or U5331 (N_5331,N_3318,N_4018);
or U5332 (N_5332,N_3494,N_3442);
or U5333 (N_5333,N_4049,N_3756);
xnor U5334 (N_5334,N_3855,N_3986);
nor U5335 (N_5335,N_4313,N_3214);
and U5336 (N_5336,N_3118,N_3177);
and U5337 (N_5337,N_3363,N_4123);
nor U5338 (N_5338,N_3878,N_3751);
xnor U5339 (N_5339,N_3264,N_3273);
or U5340 (N_5340,N_3790,N_4278);
and U5341 (N_5341,N_3396,N_4133);
nor U5342 (N_5342,N_4057,N_4196);
or U5343 (N_5343,N_3807,N_3645);
or U5344 (N_5344,N_4487,N_3977);
and U5345 (N_5345,N_3688,N_3087);
or U5346 (N_5346,N_3720,N_3962);
nor U5347 (N_5347,N_3339,N_3447);
and U5348 (N_5348,N_4029,N_3353);
nor U5349 (N_5349,N_3678,N_3894);
xor U5350 (N_5350,N_4404,N_3507);
xor U5351 (N_5351,N_3351,N_3608);
nor U5352 (N_5352,N_3250,N_4318);
xor U5353 (N_5353,N_3156,N_3078);
nor U5354 (N_5354,N_4285,N_3708);
or U5355 (N_5355,N_4414,N_3299);
nor U5356 (N_5356,N_3137,N_3743);
nor U5357 (N_5357,N_4041,N_3361);
nand U5358 (N_5358,N_4363,N_3538);
xnor U5359 (N_5359,N_3172,N_3853);
nor U5360 (N_5360,N_3743,N_3837);
or U5361 (N_5361,N_3596,N_4413);
nor U5362 (N_5362,N_3867,N_4498);
or U5363 (N_5363,N_3238,N_4175);
or U5364 (N_5364,N_3483,N_4225);
and U5365 (N_5365,N_3686,N_3555);
nor U5366 (N_5366,N_3660,N_3695);
and U5367 (N_5367,N_4197,N_3409);
nor U5368 (N_5368,N_3977,N_3196);
xnor U5369 (N_5369,N_4139,N_4165);
nand U5370 (N_5370,N_3489,N_3960);
xor U5371 (N_5371,N_4375,N_4075);
nor U5372 (N_5372,N_4278,N_4452);
nor U5373 (N_5373,N_3106,N_3171);
and U5374 (N_5374,N_4357,N_3315);
nor U5375 (N_5375,N_3371,N_3611);
or U5376 (N_5376,N_4027,N_3818);
or U5377 (N_5377,N_3770,N_3755);
xor U5378 (N_5378,N_3900,N_3177);
xor U5379 (N_5379,N_3674,N_3824);
and U5380 (N_5380,N_4319,N_3445);
nand U5381 (N_5381,N_4489,N_4196);
or U5382 (N_5382,N_3207,N_4075);
xor U5383 (N_5383,N_3124,N_3187);
xor U5384 (N_5384,N_3839,N_3197);
nor U5385 (N_5385,N_3356,N_4208);
and U5386 (N_5386,N_3907,N_3272);
nor U5387 (N_5387,N_3723,N_3856);
or U5388 (N_5388,N_3400,N_3148);
xnor U5389 (N_5389,N_4244,N_3240);
nand U5390 (N_5390,N_3307,N_3249);
nand U5391 (N_5391,N_4383,N_3602);
nand U5392 (N_5392,N_3775,N_3086);
or U5393 (N_5393,N_3240,N_3456);
nor U5394 (N_5394,N_3093,N_3584);
nand U5395 (N_5395,N_3508,N_3195);
and U5396 (N_5396,N_3427,N_3324);
xor U5397 (N_5397,N_3846,N_3018);
nor U5398 (N_5398,N_4435,N_3227);
xnor U5399 (N_5399,N_3414,N_3452);
nand U5400 (N_5400,N_3530,N_4209);
xnor U5401 (N_5401,N_3235,N_3471);
nand U5402 (N_5402,N_4010,N_3447);
and U5403 (N_5403,N_3066,N_4105);
nor U5404 (N_5404,N_3013,N_3398);
nand U5405 (N_5405,N_3474,N_3094);
nand U5406 (N_5406,N_3257,N_4431);
xor U5407 (N_5407,N_4177,N_3967);
nand U5408 (N_5408,N_3940,N_3218);
nand U5409 (N_5409,N_3324,N_3946);
xnor U5410 (N_5410,N_3356,N_4299);
xor U5411 (N_5411,N_3573,N_4126);
or U5412 (N_5412,N_4042,N_3934);
or U5413 (N_5413,N_4070,N_4135);
and U5414 (N_5414,N_3660,N_3858);
nor U5415 (N_5415,N_4337,N_3528);
nand U5416 (N_5416,N_3091,N_4178);
nand U5417 (N_5417,N_3223,N_3502);
nand U5418 (N_5418,N_3468,N_4171);
and U5419 (N_5419,N_3900,N_3297);
nor U5420 (N_5420,N_3941,N_3993);
nor U5421 (N_5421,N_3736,N_4357);
nand U5422 (N_5422,N_4209,N_3198);
or U5423 (N_5423,N_3936,N_4316);
xor U5424 (N_5424,N_3090,N_3935);
nor U5425 (N_5425,N_3159,N_3504);
nand U5426 (N_5426,N_3735,N_3081);
and U5427 (N_5427,N_4230,N_3290);
or U5428 (N_5428,N_3266,N_4045);
xnor U5429 (N_5429,N_3293,N_4270);
xor U5430 (N_5430,N_4298,N_3537);
xnor U5431 (N_5431,N_3765,N_4428);
nand U5432 (N_5432,N_3748,N_4441);
and U5433 (N_5433,N_3195,N_3504);
nor U5434 (N_5434,N_4321,N_4371);
or U5435 (N_5435,N_3246,N_3765);
nand U5436 (N_5436,N_3274,N_3617);
xnor U5437 (N_5437,N_3071,N_3945);
nor U5438 (N_5438,N_3903,N_3353);
and U5439 (N_5439,N_3306,N_4484);
xnor U5440 (N_5440,N_4086,N_3832);
and U5441 (N_5441,N_4485,N_4119);
xor U5442 (N_5442,N_4330,N_3007);
or U5443 (N_5443,N_3654,N_3948);
nand U5444 (N_5444,N_3761,N_3770);
nor U5445 (N_5445,N_3578,N_4142);
xnor U5446 (N_5446,N_3678,N_3497);
or U5447 (N_5447,N_4211,N_4350);
or U5448 (N_5448,N_3381,N_3916);
and U5449 (N_5449,N_4108,N_4306);
xnor U5450 (N_5450,N_3834,N_4023);
nor U5451 (N_5451,N_3818,N_4425);
or U5452 (N_5452,N_4358,N_3533);
nand U5453 (N_5453,N_3707,N_4042);
nand U5454 (N_5454,N_3759,N_3271);
nor U5455 (N_5455,N_3415,N_3913);
or U5456 (N_5456,N_3486,N_3883);
and U5457 (N_5457,N_3561,N_3829);
or U5458 (N_5458,N_4464,N_4431);
and U5459 (N_5459,N_3517,N_4461);
and U5460 (N_5460,N_4498,N_4227);
xor U5461 (N_5461,N_4043,N_4256);
and U5462 (N_5462,N_4179,N_3404);
nor U5463 (N_5463,N_3113,N_3742);
and U5464 (N_5464,N_3532,N_3751);
or U5465 (N_5465,N_3140,N_3938);
or U5466 (N_5466,N_4281,N_3912);
nand U5467 (N_5467,N_4221,N_3162);
nand U5468 (N_5468,N_3919,N_3152);
xor U5469 (N_5469,N_3253,N_3060);
or U5470 (N_5470,N_4116,N_3085);
xnor U5471 (N_5471,N_4030,N_3988);
xnor U5472 (N_5472,N_4471,N_4183);
nor U5473 (N_5473,N_4306,N_3852);
xor U5474 (N_5474,N_3996,N_3468);
nor U5475 (N_5475,N_3211,N_3182);
nor U5476 (N_5476,N_4492,N_4048);
xnor U5477 (N_5477,N_3399,N_3662);
or U5478 (N_5478,N_4044,N_4096);
nor U5479 (N_5479,N_3894,N_3167);
and U5480 (N_5480,N_4041,N_3116);
nand U5481 (N_5481,N_3650,N_4323);
or U5482 (N_5482,N_3934,N_4494);
xor U5483 (N_5483,N_3549,N_4151);
and U5484 (N_5484,N_4416,N_3183);
nand U5485 (N_5485,N_3109,N_3578);
and U5486 (N_5486,N_3643,N_4390);
nor U5487 (N_5487,N_4052,N_3866);
nor U5488 (N_5488,N_3687,N_3283);
or U5489 (N_5489,N_3659,N_4434);
nand U5490 (N_5490,N_3223,N_3886);
xor U5491 (N_5491,N_4332,N_3632);
nand U5492 (N_5492,N_4070,N_3450);
nor U5493 (N_5493,N_4426,N_4001);
nand U5494 (N_5494,N_4229,N_4401);
xnor U5495 (N_5495,N_4251,N_3227);
nand U5496 (N_5496,N_3070,N_3540);
or U5497 (N_5497,N_3356,N_3093);
or U5498 (N_5498,N_3360,N_3454);
nor U5499 (N_5499,N_3604,N_3090);
nand U5500 (N_5500,N_3226,N_4292);
and U5501 (N_5501,N_4068,N_3275);
nor U5502 (N_5502,N_3034,N_4182);
and U5503 (N_5503,N_3161,N_3728);
nand U5504 (N_5504,N_3601,N_3742);
xnor U5505 (N_5505,N_3881,N_3021);
and U5506 (N_5506,N_3446,N_3774);
xor U5507 (N_5507,N_3639,N_3995);
and U5508 (N_5508,N_3489,N_3469);
or U5509 (N_5509,N_3548,N_3384);
nor U5510 (N_5510,N_3884,N_3957);
and U5511 (N_5511,N_4358,N_3951);
and U5512 (N_5512,N_3314,N_4156);
or U5513 (N_5513,N_3627,N_3421);
nor U5514 (N_5514,N_3069,N_3647);
nand U5515 (N_5515,N_4259,N_4291);
and U5516 (N_5516,N_3391,N_3767);
xor U5517 (N_5517,N_3313,N_3811);
or U5518 (N_5518,N_3647,N_3467);
nand U5519 (N_5519,N_3608,N_3385);
xnor U5520 (N_5520,N_3901,N_3143);
xnor U5521 (N_5521,N_3422,N_4444);
nand U5522 (N_5522,N_3723,N_4130);
nor U5523 (N_5523,N_3365,N_3109);
or U5524 (N_5524,N_3561,N_3715);
xnor U5525 (N_5525,N_4373,N_3347);
nor U5526 (N_5526,N_3153,N_3899);
and U5527 (N_5527,N_3301,N_3483);
and U5528 (N_5528,N_4081,N_3904);
or U5529 (N_5529,N_3739,N_3882);
xor U5530 (N_5530,N_4254,N_3089);
xor U5531 (N_5531,N_4005,N_4155);
or U5532 (N_5532,N_4341,N_4051);
nor U5533 (N_5533,N_4265,N_3086);
nor U5534 (N_5534,N_3903,N_4275);
nand U5535 (N_5535,N_3968,N_3239);
nor U5536 (N_5536,N_3837,N_3060);
nor U5537 (N_5537,N_3639,N_3086);
nand U5538 (N_5538,N_4028,N_3520);
or U5539 (N_5539,N_3569,N_3230);
xor U5540 (N_5540,N_3471,N_3673);
nor U5541 (N_5541,N_4377,N_3622);
or U5542 (N_5542,N_4458,N_4178);
or U5543 (N_5543,N_3639,N_3141);
nand U5544 (N_5544,N_3247,N_4082);
nand U5545 (N_5545,N_3716,N_4499);
and U5546 (N_5546,N_4127,N_4305);
xor U5547 (N_5547,N_3034,N_3426);
or U5548 (N_5548,N_3474,N_3375);
nand U5549 (N_5549,N_3972,N_3929);
and U5550 (N_5550,N_3227,N_3344);
and U5551 (N_5551,N_3697,N_3103);
nand U5552 (N_5552,N_3799,N_4014);
xnor U5553 (N_5553,N_3138,N_3106);
and U5554 (N_5554,N_3011,N_4254);
nor U5555 (N_5555,N_4139,N_4408);
or U5556 (N_5556,N_3697,N_3112);
and U5557 (N_5557,N_3232,N_4318);
nor U5558 (N_5558,N_4341,N_3181);
nor U5559 (N_5559,N_3639,N_4230);
or U5560 (N_5560,N_4021,N_3086);
and U5561 (N_5561,N_4267,N_3655);
or U5562 (N_5562,N_3603,N_3536);
nor U5563 (N_5563,N_3262,N_3648);
nand U5564 (N_5564,N_3806,N_3880);
nand U5565 (N_5565,N_3982,N_3815);
xnor U5566 (N_5566,N_3915,N_4126);
and U5567 (N_5567,N_3665,N_3163);
and U5568 (N_5568,N_3314,N_3160);
nor U5569 (N_5569,N_4324,N_3854);
xor U5570 (N_5570,N_3110,N_4389);
nand U5571 (N_5571,N_4055,N_4226);
xor U5572 (N_5572,N_3055,N_3592);
and U5573 (N_5573,N_3078,N_3606);
nor U5574 (N_5574,N_3997,N_3683);
nor U5575 (N_5575,N_3555,N_4342);
nand U5576 (N_5576,N_3644,N_4335);
nor U5577 (N_5577,N_3357,N_3514);
nand U5578 (N_5578,N_3689,N_4432);
nand U5579 (N_5579,N_4419,N_3291);
xor U5580 (N_5580,N_4191,N_3753);
nand U5581 (N_5581,N_4297,N_3116);
nor U5582 (N_5582,N_3100,N_3704);
and U5583 (N_5583,N_3606,N_3127);
nor U5584 (N_5584,N_4466,N_3244);
and U5585 (N_5585,N_3337,N_4389);
and U5586 (N_5586,N_3296,N_3580);
xor U5587 (N_5587,N_3202,N_4373);
and U5588 (N_5588,N_3880,N_3535);
nor U5589 (N_5589,N_3447,N_4040);
or U5590 (N_5590,N_3035,N_3984);
nor U5591 (N_5591,N_3051,N_4174);
nand U5592 (N_5592,N_3947,N_3952);
nand U5593 (N_5593,N_3911,N_3005);
nor U5594 (N_5594,N_3971,N_3690);
or U5595 (N_5595,N_3312,N_4261);
or U5596 (N_5596,N_4210,N_3292);
nor U5597 (N_5597,N_4378,N_3277);
nand U5598 (N_5598,N_3665,N_3383);
nand U5599 (N_5599,N_3710,N_4453);
nand U5600 (N_5600,N_3384,N_4460);
and U5601 (N_5601,N_3960,N_3138);
nand U5602 (N_5602,N_3318,N_3398);
and U5603 (N_5603,N_4193,N_4372);
nand U5604 (N_5604,N_4107,N_4234);
or U5605 (N_5605,N_4195,N_3578);
xnor U5606 (N_5606,N_3431,N_4178);
nand U5607 (N_5607,N_3335,N_4315);
and U5608 (N_5608,N_3751,N_3012);
nand U5609 (N_5609,N_3223,N_3536);
xor U5610 (N_5610,N_3845,N_3101);
and U5611 (N_5611,N_3664,N_3630);
nand U5612 (N_5612,N_3495,N_4481);
xor U5613 (N_5613,N_4286,N_3793);
and U5614 (N_5614,N_3552,N_3034);
nand U5615 (N_5615,N_4283,N_3906);
and U5616 (N_5616,N_3743,N_3005);
or U5617 (N_5617,N_3734,N_3809);
nor U5618 (N_5618,N_3793,N_3637);
and U5619 (N_5619,N_3761,N_3465);
xor U5620 (N_5620,N_3239,N_4194);
or U5621 (N_5621,N_3011,N_3476);
nand U5622 (N_5622,N_4401,N_4430);
xor U5623 (N_5623,N_3910,N_4430);
nor U5624 (N_5624,N_3307,N_3391);
nand U5625 (N_5625,N_4285,N_3196);
or U5626 (N_5626,N_4007,N_4112);
nor U5627 (N_5627,N_4439,N_3233);
or U5628 (N_5628,N_4419,N_3233);
or U5629 (N_5629,N_3100,N_4420);
nand U5630 (N_5630,N_3423,N_3708);
and U5631 (N_5631,N_4446,N_4226);
xnor U5632 (N_5632,N_4231,N_3933);
or U5633 (N_5633,N_3981,N_4144);
and U5634 (N_5634,N_3159,N_3378);
and U5635 (N_5635,N_3386,N_4138);
xor U5636 (N_5636,N_4117,N_3648);
and U5637 (N_5637,N_4475,N_3926);
xor U5638 (N_5638,N_4313,N_3574);
or U5639 (N_5639,N_3674,N_3717);
nand U5640 (N_5640,N_3654,N_4420);
nand U5641 (N_5641,N_4027,N_3657);
nor U5642 (N_5642,N_4007,N_4286);
nand U5643 (N_5643,N_3345,N_3659);
nand U5644 (N_5644,N_3008,N_4319);
or U5645 (N_5645,N_3163,N_3980);
nor U5646 (N_5646,N_3167,N_4378);
nand U5647 (N_5647,N_3894,N_3107);
nand U5648 (N_5648,N_3703,N_3251);
nor U5649 (N_5649,N_3364,N_3904);
or U5650 (N_5650,N_3982,N_4123);
xnor U5651 (N_5651,N_3883,N_3405);
or U5652 (N_5652,N_4018,N_3577);
nand U5653 (N_5653,N_3634,N_3760);
and U5654 (N_5654,N_4242,N_4234);
and U5655 (N_5655,N_4432,N_3927);
nand U5656 (N_5656,N_3130,N_3719);
or U5657 (N_5657,N_4177,N_4356);
xnor U5658 (N_5658,N_3113,N_3760);
or U5659 (N_5659,N_3334,N_3064);
or U5660 (N_5660,N_4154,N_4264);
and U5661 (N_5661,N_3386,N_3040);
or U5662 (N_5662,N_3372,N_3191);
and U5663 (N_5663,N_3692,N_4370);
or U5664 (N_5664,N_3951,N_3463);
nor U5665 (N_5665,N_3913,N_3079);
or U5666 (N_5666,N_3711,N_4235);
xor U5667 (N_5667,N_3629,N_4152);
xor U5668 (N_5668,N_3795,N_3640);
nor U5669 (N_5669,N_4100,N_3829);
and U5670 (N_5670,N_3915,N_3826);
nand U5671 (N_5671,N_3830,N_4410);
xor U5672 (N_5672,N_3582,N_3041);
and U5673 (N_5673,N_4252,N_4195);
xnor U5674 (N_5674,N_3905,N_3577);
nand U5675 (N_5675,N_3643,N_4206);
or U5676 (N_5676,N_4085,N_3139);
xor U5677 (N_5677,N_3354,N_3199);
nor U5678 (N_5678,N_3337,N_4218);
nand U5679 (N_5679,N_4078,N_4204);
or U5680 (N_5680,N_3493,N_3001);
nor U5681 (N_5681,N_3877,N_3526);
nor U5682 (N_5682,N_3489,N_3910);
xnor U5683 (N_5683,N_3879,N_4377);
and U5684 (N_5684,N_3965,N_3710);
or U5685 (N_5685,N_4295,N_3817);
nor U5686 (N_5686,N_4453,N_3505);
nand U5687 (N_5687,N_4202,N_3682);
nor U5688 (N_5688,N_4417,N_4010);
xor U5689 (N_5689,N_4102,N_4369);
and U5690 (N_5690,N_4477,N_3396);
xnor U5691 (N_5691,N_3589,N_3503);
and U5692 (N_5692,N_4206,N_3604);
xor U5693 (N_5693,N_4430,N_3921);
nor U5694 (N_5694,N_4487,N_4362);
xor U5695 (N_5695,N_3997,N_4086);
and U5696 (N_5696,N_3235,N_3079);
nand U5697 (N_5697,N_3372,N_3938);
xor U5698 (N_5698,N_3647,N_3788);
nor U5699 (N_5699,N_3843,N_3988);
or U5700 (N_5700,N_3782,N_3245);
nand U5701 (N_5701,N_4156,N_3674);
nand U5702 (N_5702,N_3691,N_4245);
nand U5703 (N_5703,N_3672,N_4253);
xnor U5704 (N_5704,N_3138,N_3891);
or U5705 (N_5705,N_3621,N_3840);
and U5706 (N_5706,N_3501,N_4040);
and U5707 (N_5707,N_4056,N_3672);
and U5708 (N_5708,N_3654,N_4040);
nor U5709 (N_5709,N_3570,N_4387);
nor U5710 (N_5710,N_3435,N_3388);
nand U5711 (N_5711,N_3529,N_3729);
nor U5712 (N_5712,N_4135,N_3205);
xnor U5713 (N_5713,N_4133,N_3319);
or U5714 (N_5714,N_3041,N_4382);
and U5715 (N_5715,N_4118,N_3328);
or U5716 (N_5716,N_4025,N_3708);
nor U5717 (N_5717,N_4396,N_3233);
nand U5718 (N_5718,N_3052,N_3403);
nor U5719 (N_5719,N_4309,N_3982);
xor U5720 (N_5720,N_3598,N_3668);
xnor U5721 (N_5721,N_3178,N_4042);
and U5722 (N_5722,N_3815,N_4246);
and U5723 (N_5723,N_4204,N_3473);
xnor U5724 (N_5724,N_3575,N_3838);
nor U5725 (N_5725,N_3213,N_3771);
nand U5726 (N_5726,N_4202,N_4026);
xor U5727 (N_5727,N_3638,N_3299);
and U5728 (N_5728,N_3472,N_3218);
xnor U5729 (N_5729,N_3900,N_4050);
nand U5730 (N_5730,N_4369,N_3963);
or U5731 (N_5731,N_3029,N_3974);
and U5732 (N_5732,N_3901,N_4057);
xor U5733 (N_5733,N_3062,N_3322);
or U5734 (N_5734,N_3085,N_4401);
and U5735 (N_5735,N_3013,N_3321);
or U5736 (N_5736,N_4210,N_4328);
nor U5737 (N_5737,N_3234,N_3384);
or U5738 (N_5738,N_3685,N_4250);
xor U5739 (N_5739,N_4483,N_4333);
or U5740 (N_5740,N_3028,N_3427);
nor U5741 (N_5741,N_3380,N_3475);
nand U5742 (N_5742,N_3552,N_4116);
nand U5743 (N_5743,N_3367,N_3664);
xor U5744 (N_5744,N_3495,N_3208);
nand U5745 (N_5745,N_4158,N_3446);
and U5746 (N_5746,N_3847,N_3169);
or U5747 (N_5747,N_3291,N_3113);
and U5748 (N_5748,N_3923,N_4477);
nand U5749 (N_5749,N_3546,N_3462);
nand U5750 (N_5750,N_4488,N_3095);
or U5751 (N_5751,N_3497,N_3336);
nand U5752 (N_5752,N_3611,N_3031);
nor U5753 (N_5753,N_3676,N_3688);
xnor U5754 (N_5754,N_4265,N_3764);
nand U5755 (N_5755,N_3607,N_4200);
and U5756 (N_5756,N_3716,N_3140);
xnor U5757 (N_5757,N_4367,N_3124);
nand U5758 (N_5758,N_3335,N_3019);
nand U5759 (N_5759,N_4124,N_3539);
and U5760 (N_5760,N_3118,N_3037);
xnor U5761 (N_5761,N_4266,N_3239);
nand U5762 (N_5762,N_3895,N_4205);
xnor U5763 (N_5763,N_4490,N_4497);
or U5764 (N_5764,N_4293,N_3927);
nand U5765 (N_5765,N_4054,N_3513);
or U5766 (N_5766,N_3253,N_3347);
nor U5767 (N_5767,N_4250,N_3390);
and U5768 (N_5768,N_3666,N_4418);
nand U5769 (N_5769,N_3069,N_3251);
or U5770 (N_5770,N_3887,N_3041);
and U5771 (N_5771,N_4466,N_3973);
and U5772 (N_5772,N_3401,N_4327);
and U5773 (N_5773,N_3832,N_4234);
nor U5774 (N_5774,N_4270,N_4395);
nor U5775 (N_5775,N_4033,N_3333);
and U5776 (N_5776,N_3556,N_3521);
nand U5777 (N_5777,N_3155,N_4326);
nor U5778 (N_5778,N_4123,N_3352);
and U5779 (N_5779,N_3954,N_4205);
or U5780 (N_5780,N_4211,N_3116);
nor U5781 (N_5781,N_3745,N_3026);
xor U5782 (N_5782,N_4246,N_3858);
xor U5783 (N_5783,N_4206,N_3221);
nand U5784 (N_5784,N_4350,N_3185);
nor U5785 (N_5785,N_3118,N_3509);
or U5786 (N_5786,N_3239,N_3976);
or U5787 (N_5787,N_3564,N_4194);
or U5788 (N_5788,N_3853,N_3201);
or U5789 (N_5789,N_3082,N_3353);
and U5790 (N_5790,N_4096,N_3585);
xnor U5791 (N_5791,N_3083,N_3306);
and U5792 (N_5792,N_4033,N_3165);
nor U5793 (N_5793,N_4309,N_3679);
or U5794 (N_5794,N_3313,N_4223);
nor U5795 (N_5795,N_3006,N_3132);
and U5796 (N_5796,N_3479,N_4211);
xor U5797 (N_5797,N_3326,N_3025);
and U5798 (N_5798,N_3653,N_4253);
or U5799 (N_5799,N_3556,N_3923);
nand U5800 (N_5800,N_3861,N_3294);
or U5801 (N_5801,N_3249,N_4136);
and U5802 (N_5802,N_4333,N_3865);
or U5803 (N_5803,N_3376,N_3834);
xnor U5804 (N_5804,N_4153,N_3886);
or U5805 (N_5805,N_4484,N_3130);
xnor U5806 (N_5806,N_3442,N_4440);
and U5807 (N_5807,N_4210,N_3513);
nor U5808 (N_5808,N_4101,N_3068);
nand U5809 (N_5809,N_4404,N_3191);
nand U5810 (N_5810,N_3902,N_3422);
and U5811 (N_5811,N_3085,N_3487);
xor U5812 (N_5812,N_3994,N_3101);
nand U5813 (N_5813,N_3272,N_3958);
or U5814 (N_5814,N_4313,N_3824);
xnor U5815 (N_5815,N_3192,N_3104);
nor U5816 (N_5816,N_3580,N_4135);
nand U5817 (N_5817,N_4393,N_3331);
xor U5818 (N_5818,N_3389,N_3108);
xnor U5819 (N_5819,N_3137,N_4160);
nor U5820 (N_5820,N_3406,N_4247);
xnor U5821 (N_5821,N_4259,N_4475);
and U5822 (N_5822,N_3662,N_4344);
xnor U5823 (N_5823,N_3652,N_4015);
nand U5824 (N_5824,N_3784,N_4343);
and U5825 (N_5825,N_4280,N_3674);
xor U5826 (N_5826,N_4108,N_3220);
xor U5827 (N_5827,N_4456,N_4144);
xor U5828 (N_5828,N_4318,N_3368);
and U5829 (N_5829,N_4400,N_3872);
nor U5830 (N_5830,N_4268,N_4458);
xor U5831 (N_5831,N_3504,N_3680);
and U5832 (N_5832,N_3273,N_4271);
and U5833 (N_5833,N_4035,N_4376);
xor U5834 (N_5834,N_4310,N_3917);
and U5835 (N_5835,N_3257,N_3983);
or U5836 (N_5836,N_4006,N_4211);
and U5837 (N_5837,N_3857,N_4330);
and U5838 (N_5838,N_4359,N_3568);
xor U5839 (N_5839,N_4172,N_3086);
nand U5840 (N_5840,N_3054,N_4293);
xnor U5841 (N_5841,N_4136,N_4064);
nand U5842 (N_5842,N_4053,N_3079);
nand U5843 (N_5843,N_3209,N_3609);
nor U5844 (N_5844,N_3529,N_4028);
and U5845 (N_5845,N_4404,N_3725);
xor U5846 (N_5846,N_4253,N_3469);
nor U5847 (N_5847,N_3440,N_3278);
or U5848 (N_5848,N_4089,N_3354);
or U5849 (N_5849,N_4301,N_4482);
and U5850 (N_5850,N_4181,N_3019);
nand U5851 (N_5851,N_3456,N_4165);
nor U5852 (N_5852,N_3831,N_3102);
nand U5853 (N_5853,N_3517,N_4331);
nand U5854 (N_5854,N_3518,N_4185);
or U5855 (N_5855,N_3328,N_3233);
nand U5856 (N_5856,N_3542,N_3797);
nand U5857 (N_5857,N_3215,N_4316);
and U5858 (N_5858,N_3063,N_4079);
and U5859 (N_5859,N_4340,N_3949);
nand U5860 (N_5860,N_4414,N_3912);
and U5861 (N_5861,N_4181,N_3569);
nor U5862 (N_5862,N_3119,N_3215);
and U5863 (N_5863,N_4227,N_4372);
or U5864 (N_5864,N_3427,N_3570);
xnor U5865 (N_5865,N_3811,N_3719);
or U5866 (N_5866,N_4195,N_3637);
and U5867 (N_5867,N_3365,N_3935);
xor U5868 (N_5868,N_4048,N_3125);
nor U5869 (N_5869,N_3245,N_3870);
or U5870 (N_5870,N_4103,N_4343);
nand U5871 (N_5871,N_3515,N_4499);
nor U5872 (N_5872,N_4391,N_3956);
nand U5873 (N_5873,N_3196,N_4314);
or U5874 (N_5874,N_3382,N_3034);
or U5875 (N_5875,N_3528,N_3520);
nor U5876 (N_5876,N_4038,N_3111);
nand U5877 (N_5877,N_3091,N_3235);
xnor U5878 (N_5878,N_3969,N_4064);
nand U5879 (N_5879,N_3018,N_3912);
and U5880 (N_5880,N_3278,N_4362);
nand U5881 (N_5881,N_3575,N_3830);
and U5882 (N_5882,N_4169,N_4350);
and U5883 (N_5883,N_3318,N_3431);
and U5884 (N_5884,N_3842,N_3110);
and U5885 (N_5885,N_3306,N_3716);
xnor U5886 (N_5886,N_3093,N_3205);
nor U5887 (N_5887,N_3702,N_4103);
and U5888 (N_5888,N_4496,N_3262);
nand U5889 (N_5889,N_4043,N_4090);
nor U5890 (N_5890,N_4300,N_3842);
or U5891 (N_5891,N_3719,N_3235);
and U5892 (N_5892,N_4494,N_4158);
or U5893 (N_5893,N_3800,N_3998);
and U5894 (N_5894,N_4337,N_3999);
nor U5895 (N_5895,N_4463,N_3217);
nand U5896 (N_5896,N_3419,N_4122);
or U5897 (N_5897,N_3895,N_3595);
and U5898 (N_5898,N_3901,N_4329);
and U5899 (N_5899,N_4336,N_3462);
nor U5900 (N_5900,N_3258,N_3344);
nand U5901 (N_5901,N_3064,N_4071);
and U5902 (N_5902,N_4473,N_4246);
or U5903 (N_5903,N_4383,N_3633);
or U5904 (N_5904,N_3449,N_3154);
nor U5905 (N_5905,N_4303,N_3928);
xnor U5906 (N_5906,N_3567,N_3578);
nand U5907 (N_5907,N_3252,N_3329);
and U5908 (N_5908,N_4001,N_3359);
nor U5909 (N_5909,N_3760,N_3120);
xor U5910 (N_5910,N_4162,N_3691);
xor U5911 (N_5911,N_3808,N_3021);
and U5912 (N_5912,N_4307,N_3334);
nor U5913 (N_5913,N_4107,N_3241);
nand U5914 (N_5914,N_3545,N_3851);
nor U5915 (N_5915,N_4138,N_3323);
xor U5916 (N_5916,N_3982,N_4439);
xor U5917 (N_5917,N_3369,N_3312);
nor U5918 (N_5918,N_4323,N_3801);
nor U5919 (N_5919,N_3284,N_4150);
xor U5920 (N_5920,N_3641,N_3967);
nand U5921 (N_5921,N_3764,N_3782);
or U5922 (N_5922,N_4302,N_4454);
nor U5923 (N_5923,N_3091,N_3063);
nor U5924 (N_5924,N_3997,N_4421);
or U5925 (N_5925,N_3833,N_3813);
or U5926 (N_5926,N_3371,N_4268);
nand U5927 (N_5927,N_3452,N_3030);
nor U5928 (N_5928,N_3086,N_3814);
nor U5929 (N_5929,N_4468,N_4381);
and U5930 (N_5930,N_3743,N_3930);
nor U5931 (N_5931,N_3779,N_3424);
nand U5932 (N_5932,N_3586,N_4111);
xor U5933 (N_5933,N_3980,N_3446);
or U5934 (N_5934,N_4032,N_4130);
or U5935 (N_5935,N_3442,N_3987);
nor U5936 (N_5936,N_3567,N_4124);
nor U5937 (N_5937,N_4401,N_4423);
or U5938 (N_5938,N_3195,N_4209);
nor U5939 (N_5939,N_4359,N_4267);
and U5940 (N_5940,N_4068,N_3485);
nand U5941 (N_5941,N_3676,N_3694);
nand U5942 (N_5942,N_4304,N_4045);
and U5943 (N_5943,N_3921,N_4017);
xnor U5944 (N_5944,N_3891,N_4087);
and U5945 (N_5945,N_3154,N_3020);
xnor U5946 (N_5946,N_4351,N_4106);
nand U5947 (N_5947,N_3596,N_3911);
xor U5948 (N_5948,N_3423,N_3242);
or U5949 (N_5949,N_4457,N_4466);
xor U5950 (N_5950,N_3630,N_3338);
nand U5951 (N_5951,N_4188,N_4179);
nand U5952 (N_5952,N_4089,N_3390);
or U5953 (N_5953,N_3874,N_3267);
nand U5954 (N_5954,N_3804,N_3326);
nor U5955 (N_5955,N_3979,N_4346);
xnor U5956 (N_5956,N_3288,N_4306);
nand U5957 (N_5957,N_3432,N_4395);
or U5958 (N_5958,N_4182,N_3243);
xnor U5959 (N_5959,N_3652,N_4342);
or U5960 (N_5960,N_3973,N_4028);
and U5961 (N_5961,N_3953,N_4046);
or U5962 (N_5962,N_3147,N_3452);
nand U5963 (N_5963,N_3498,N_4151);
xnor U5964 (N_5964,N_3758,N_3558);
and U5965 (N_5965,N_3212,N_3147);
nand U5966 (N_5966,N_3179,N_3023);
nor U5967 (N_5967,N_3642,N_4343);
and U5968 (N_5968,N_4113,N_3774);
nand U5969 (N_5969,N_3713,N_3386);
nand U5970 (N_5970,N_3773,N_3974);
xnor U5971 (N_5971,N_3351,N_3556);
nor U5972 (N_5972,N_4214,N_4473);
and U5973 (N_5973,N_3923,N_4100);
and U5974 (N_5974,N_3268,N_4294);
xor U5975 (N_5975,N_4006,N_3360);
xor U5976 (N_5976,N_4048,N_3782);
nand U5977 (N_5977,N_3482,N_4295);
or U5978 (N_5978,N_3962,N_3195);
nor U5979 (N_5979,N_3679,N_4226);
and U5980 (N_5980,N_3583,N_4022);
or U5981 (N_5981,N_3453,N_3454);
xnor U5982 (N_5982,N_3420,N_3782);
nor U5983 (N_5983,N_3512,N_3760);
or U5984 (N_5984,N_3530,N_4497);
and U5985 (N_5985,N_4476,N_4050);
or U5986 (N_5986,N_3494,N_3809);
nor U5987 (N_5987,N_3041,N_4097);
or U5988 (N_5988,N_4315,N_3903);
nor U5989 (N_5989,N_3489,N_3801);
nand U5990 (N_5990,N_4462,N_3539);
or U5991 (N_5991,N_4303,N_3680);
nand U5992 (N_5992,N_3354,N_3580);
and U5993 (N_5993,N_3183,N_3674);
nand U5994 (N_5994,N_3400,N_3364);
xnor U5995 (N_5995,N_3852,N_3897);
and U5996 (N_5996,N_3138,N_3695);
nand U5997 (N_5997,N_3985,N_3816);
nor U5998 (N_5998,N_4142,N_3127);
nor U5999 (N_5999,N_4413,N_3116);
xnor U6000 (N_6000,N_4927,N_5343);
nor U6001 (N_6001,N_4683,N_4892);
or U6002 (N_6002,N_4619,N_4844);
xor U6003 (N_6003,N_5455,N_5276);
or U6004 (N_6004,N_4591,N_4880);
nor U6005 (N_6005,N_5175,N_5417);
nand U6006 (N_6006,N_5333,N_5541);
xor U6007 (N_6007,N_4560,N_5006);
nand U6008 (N_6008,N_4748,N_5353);
nor U6009 (N_6009,N_4868,N_5387);
nor U6010 (N_6010,N_5802,N_5344);
and U6011 (N_6011,N_5866,N_4674);
nand U6012 (N_6012,N_5976,N_4825);
nand U6013 (N_6013,N_5349,N_4548);
xor U6014 (N_6014,N_4506,N_5862);
nor U6015 (N_6015,N_4830,N_4753);
nor U6016 (N_6016,N_5314,N_4948);
xor U6017 (N_6017,N_4607,N_5169);
nor U6018 (N_6018,N_5577,N_5003);
or U6019 (N_6019,N_4514,N_5555);
nor U6020 (N_6020,N_5717,N_5610);
nor U6021 (N_6021,N_4966,N_5737);
or U6022 (N_6022,N_4983,N_5328);
xnor U6023 (N_6023,N_5616,N_5882);
nor U6024 (N_6024,N_5659,N_4552);
nor U6025 (N_6025,N_4920,N_5670);
nand U6026 (N_6026,N_4905,N_5162);
nand U6027 (N_6027,N_4944,N_4550);
or U6028 (N_6028,N_4863,N_5423);
or U6029 (N_6029,N_5507,N_5485);
nand U6030 (N_6030,N_5028,N_5161);
nor U6031 (N_6031,N_5655,N_5518);
and U6032 (N_6032,N_4798,N_5641);
nor U6033 (N_6033,N_4803,N_4818);
or U6034 (N_6034,N_5547,N_4677);
and U6035 (N_6035,N_5823,N_5563);
nand U6036 (N_6036,N_5639,N_4510);
nor U6037 (N_6037,N_5439,N_5415);
xor U6038 (N_6038,N_4543,N_4605);
and U6039 (N_6039,N_5073,N_5200);
or U6040 (N_6040,N_4931,N_4744);
nand U6041 (N_6041,N_5826,N_5571);
nand U6042 (N_6042,N_4870,N_5032);
and U6043 (N_6043,N_4565,N_5024);
nand U6044 (N_6044,N_5489,N_5953);
xnor U6045 (N_6045,N_5725,N_4616);
xnor U6046 (N_6046,N_5047,N_5868);
xnor U6047 (N_6047,N_5752,N_5171);
nor U6048 (N_6048,N_5474,N_4918);
xor U6049 (N_6049,N_5891,N_5093);
xor U6050 (N_6050,N_4529,N_5568);
xnor U6051 (N_6051,N_4789,N_5560);
and U6052 (N_6052,N_5100,N_5755);
xor U6053 (N_6053,N_5926,N_5111);
nor U6054 (N_6054,N_4501,N_5935);
and U6055 (N_6055,N_5844,N_5742);
nor U6056 (N_6056,N_4910,N_5875);
nand U6057 (N_6057,N_5115,N_5722);
and U6058 (N_6058,N_5812,N_4846);
and U6059 (N_6059,N_4553,N_4866);
and U6060 (N_6060,N_5818,N_5089);
or U6061 (N_6061,N_5222,N_5011);
or U6062 (N_6062,N_5512,N_4559);
and U6063 (N_6063,N_5787,N_4557);
nor U6064 (N_6064,N_5174,N_5786);
or U6065 (N_6065,N_5870,N_5217);
xor U6066 (N_6066,N_5720,N_5471);
and U6067 (N_6067,N_5556,N_5388);
and U6068 (N_6068,N_5550,N_5012);
and U6069 (N_6069,N_5470,N_5905);
and U6070 (N_6070,N_5257,N_4572);
nor U6071 (N_6071,N_4740,N_4782);
xor U6072 (N_6072,N_4581,N_5376);
and U6073 (N_6073,N_5767,N_4979);
or U6074 (N_6074,N_5298,N_5989);
nand U6075 (N_6075,N_5973,N_5212);
and U6076 (N_6076,N_4522,N_5052);
nor U6077 (N_6077,N_5040,N_5498);
and U6078 (N_6078,N_5484,N_5183);
xor U6079 (N_6079,N_5061,N_5098);
xor U6080 (N_6080,N_4662,N_4624);
nor U6081 (N_6081,N_4837,N_4615);
or U6082 (N_6082,N_5405,N_5180);
xor U6083 (N_6083,N_4527,N_5954);
nand U6084 (N_6084,N_4511,N_4673);
and U6085 (N_6085,N_4609,N_5460);
nand U6086 (N_6086,N_5766,N_5119);
nor U6087 (N_6087,N_5749,N_5172);
nand U6088 (N_6088,N_4909,N_5969);
and U6089 (N_6089,N_4823,N_5790);
nor U6090 (N_6090,N_4856,N_4541);
nand U6091 (N_6091,N_4586,N_4785);
or U6092 (N_6092,N_4596,N_5132);
nand U6093 (N_6093,N_5635,N_5943);
nand U6094 (N_6094,N_5126,N_5562);
xor U6095 (N_6095,N_5038,N_5553);
nor U6096 (N_6096,N_5207,N_4932);
nand U6097 (N_6097,N_4643,N_5760);
xnor U6098 (N_6098,N_4638,N_5253);
xnor U6099 (N_6099,N_4639,N_4562);
nand U6100 (N_6100,N_5661,N_5385);
and U6101 (N_6101,N_5480,N_5150);
nor U6102 (N_6102,N_4998,N_5004);
xnor U6103 (N_6103,N_5532,N_5227);
nor U6104 (N_6104,N_5962,N_5805);
or U6105 (N_6105,N_5998,N_4915);
and U6106 (N_6106,N_5667,N_4808);
xnor U6107 (N_6107,N_5194,N_5690);
or U6108 (N_6108,N_5522,N_4841);
and U6109 (N_6109,N_4623,N_5016);
or U6110 (N_6110,N_5595,N_5108);
or U6111 (N_6111,N_5205,N_5339);
nor U6112 (N_6112,N_5289,N_5116);
or U6113 (N_6113,N_4922,N_5516);
xnor U6114 (N_6114,N_4791,N_5352);
or U6115 (N_6115,N_4690,N_5380);
or U6116 (N_6116,N_5929,N_5015);
or U6117 (N_6117,N_5808,N_5819);
or U6118 (N_6118,N_5127,N_4908);
nand U6119 (N_6119,N_5963,N_5366);
nor U6120 (N_6120,N_5420,N_5859);
or U6121 (N_6121,N_4987,N_5481);
or U6122 (N_6122,N_5318,N_5846);
nand U6123 (N_6123,N_4821,N_4843);
or U6124 (N_6124,N_5465,N_4804);
or U6125 (N_6125,N_4579,N_5793);
and U6126 (N_6126,N_5817,N_4847);
nor U6127 (N_6127,N_5564,N_5338);
nor U6128 (N_6128,N_5806,N_5216);
xor U6129 (N_6129,N_5649,N_5694);
nor U6130 (N_6130,N_4574,N_5546);
or U6131 (N_6131,N_5299,N_4730);
and U6132 (N_6132,N_5753,N_4786);
and U6133 (N_6133,N_4681,N_4877);
xor U6134 (N_6134,N_4864,N_5219);
nand U6135 (N_6135,N_5626,N_5296);
nand U6136 (N_6136,N_5874,N_5794);
nand U6137 (N_6137,N_5734,N_5033);
nand U6138 (N_6138,N_4968,N_4770);
xnor U6139 (N_6139,N_4771,N_5044);
and U6140 (N_6140,N_4584,N_5199);
nor U6141 (N_6141,N_4715,N_5744);
xor U6142 (N_6142,N_4967,N_5966);
nand U6143 (N_6143,N_5260,N_5091);
or U6144 (N_6144,N_4589,N_5952);
or U6145 (N_6145,N_4959,N_5261);
nand U6146 (N_6146,N_4721,N_5377);
nor U6147 (N_6147,N_4942,N_5596);
and U6148 (N_6148,N_5020,N_5582);
nor U6149 (N_6149,N_4689,N_5195);
nor U6150 (N_6150,N_5579,N_5074);
or U6151 (N_6151,N_5906,N_5209);
or U6152 (N_6152,N_5167,N_5580);
nor U6153 (N_6153,N_5182,N_5660);
nor U6154 (N_6154,N_5988,N_5406);
or U6155 (N_6155,N_5431,N_5039);
nand U6156 (N_6156,N_5208,N_5304);
or U6157 (N_6157,N_5928,N_5751);
and U6158 (N_6158,N_5046,N_5715);
or U6159 (N_6159,N_5910,N_5113);
nor U6160 (N_6160,N_5697,N_5773);
nor U6161 (N_6161,N_4859,N_5849);
or U6162 (N_6162,N_5210,N_5588);
or U6163 (N_6163,N_5775,N_4928);
nand U6164 (N_6164,N_5457,N_5202);
and U6165 (N_6165,N_5931,N_4564);
and U6166 (N_6166,N_4884,N_5852);
nor U6167 (N_6167,N_5325,N_4984);
nor U6168 (N_6168,N_5869,N_4815);
and U6169 (N_6169,N_5757,N_5159);
xor U6170 (N_6170,N_5683,N_4593);
nor U6171 (N_6171,N_5668,N_5548);
xnor U6172 (N_6172,N_5398,N_5565);
xor U6173 (N_6173,N_5663,N_4570);
xor U6174 (N_6174,N_4537,N_4814);
xor U6175 (N_6175,N_5394,N_5414);
nor U6176 (N_6176,N_4929,N_5477);
xnor U6177 (N_6177,N_4536,N_5648);
xnor U6178 (N_6178,N_5357,N_5136);
nor U6179 (N_6179,N_5590,N_4861);
or U6180 (N_6180,N_5919,N_5673);
or U6181 (N_6181,N_5251,N_4760);
xor U6182 (N_6182,N_4865,N_4601);
nand U6183 (N_6183,N_4737,N_5425);
and U6184 (N_6184,N_5315,N_5619);
or U6185 (N_6185,N_5176,N_5206);
or U6186 (N_6186,N_5832,N_5959);
xnor U6187 (N_6187,N_5416,N_5982);
nand U6188 (N_6188,N_4777,N_4535);
nor U6189 (N_6189,N_5043,N_4679);
nor U6190 (N_6190,N_5572,N_4653);
nand U6191 (N_6191,N_5955,N_5835);
and U6192 (N_6192,N_5429,N_5599);
and U6193 (N_6193,N_5501,N_5008);
or U6194 (N_6194,N_5486,N_5441);
xor U6195 (N_6195,N_5552,N_5201);
xor U6196 (N_6196,N_5784,N_4568);
nor U6197 (N_6197,N_5068,N_5809);
nor U6198 (N_6198,N_4997,N_4993);
and U6199 (N_6199,N_4576,N_5937);
xor U6200 (N_6200,N_5083,N_5123);
or U6201 (N_6201,N_4508,N_5324);
xor U6202 (N_6202,N_5137,N_5204);
and U6203 (N_6203,N_4954,N_5031);
and U6204 (N_6204,N_5699,N_5617);
nand U6205 (N_6205,N_5591,N_5252);
nand U6206 (N_6206,N_4819,N_4802);
nand U6207 (N_6207,N_5458,N_5393);
or U6208 (N_6208,N_4577,N_5373);
xnor U6209 (N_6209,N_5271,N_4888);
and U6210 (N_6210,N_4829,N_5903);
and U6211 (N_6211,N_4627,N_5232);
nand U6212 (N_6212,N_5993,N_5569);
xor U6213 (N_6213,N_5270,N_5493);
xor U6214 (N_6214,N_5965,N_5614);
or U6215 (N_6215,N_5469,N_5007);
nand U6216 (N_6216,N_4783,N_5983);
xor U6217 (N_6217,N_5129,N_4569);
xnor U6218 (N_6218,N_5765,N_4608);
or U6219 (N_6219,N_4648,N_4772);
nor U6220 (N_6220,N_5292,N_4806);
nor U6221 (N_6221,N_5782,N_4886);
or U6222 (N_6222,N_5428,N_4551);
nor U6223 (N_6223,N_5278,N_5778);
or U6224 (N_6224,N_5535,N_4943);
or U6225 (N_6225,N_5144,N_5403);
nand U6226 (N_6226,N_5155,N_5951);
and U6227 (N_6227,N_5769,N_5070);
nand U6228 (N_6228,N_4645,N_4755);
nand U6229 (N_6229,N_4519,N_5118);
and U6230 (N_6230,N_5491,N_4745);
and U6231 (N_6231,N_5130,N_4917);
nor U6232 (N_6232,N_4528,N_4710);
nand U6233 (N_6233,N_5371,N_4796);
or U6234 (N_6234,N_4545,N_5308);
xnor U6235 (N_6235,N_4556,N_4775);
xnor U6236 (N_6236,N_5504,N_5029);
and U6237 (N_6237,N_5597,N_5886);
nand U6238 (N_6238,N_5446,N_4986);
nand U6239 (N_6239,N_5559,N_5598);
and U6240 (N_6240,N_5770,N_4764);
and U6241 (N_6241,N_4539,N_5710);
and U6242 (N_6242,N_5402,N_4630);
or U6243 (N_6243,N_5510,N_5379);
and U6244 (N_6244,N_5382,N_4538);
xnor U6245 (N_6245,N_4692,N_5305);
or U6246 (N_6246,N_5804,N_5059);
and U6247 (N_6247,N_5917,N_5848);
and U6248 (N_6248,N_5783,N_5702);
xor U6249 (N_6249,N_5438,N_4733);
nand U6250 (N_6250,N_5482,N_5017);
or U6251 (N_6251,N_4575,N_4716);
and U6252 (N_6252,N_5689,N_5600);
or U6253 (N_6253,N_5506,N_4502);
nand U6254 (N_6254,N_5593,N_5358);
or U6255 (N_6255,N_4773,N_4622);
nor U6256 (N_6256,N_4598,N_5570);
and U6257 (N_6257,N_5221,N_4707);
and U6258 (N_6258,N_5440,N_5378);
nor U6259 (N_6259,N_5688,N_4895);
and U6260 (N_6260,N_5631,N_4784);
nand U6261 (N_6261,N_5754,N_5154);
xor U6262 (N_6262,N_4774,N_4874);
nor U6263 (N_6263,N_5107,N_5013);
or U6264 (N_6264,N_5211,N_4792);
and U6265 (N_6265,N_5407,N_5229);
and U6266 (N_6266,N_5777,N_5367);
or U6267 (N_6267,N_5899,N_4995);
nand U6268 (N_6268,N_5307,N_5185);
nor U6269 (N_6269,N_5146,N_4835);
and U6270 (N_6270,N_5258,N_5791);
xnor U6271 (N_6271,N_4580,N_4851);
nand U6272 (N_6272,N_4686,N_5992);
xor U6273 (N_6273,N_5291,N_5530);
nor U6274 (N_6274,N_5274,N_5459);
xor U6275 (N_6275,N_5948,N_4824);
nor U6276 (N_6276,N_4964,N_4972);
xnor U6277 (N_6277,N_5540,N_5728);
nand U6278 (N_6278,N_5557,N_4566);
or U6279 (N_6279,N_5938,N_5190);
and U6280 (N_6280,N_5657,N_4695);
and U6281 (N_6281,N_5424,N_5601);
nor U6282 (N_6282,N_5500,N_5288);
or U6283 (N_6283,N_4743,N_4655);
and U6284 (N_6284,N_5283,N_5196);
and U6285 (N_6285,N_4694,N_5084);
and U6286 (N_6286,N_4853,N_5476);
and U6287 (N_6287,N_5748,N_5233);
nand U6288 (N_6288,N_5456,N_5691);
nand U6289 (N_6289,N_5957,N_5079);
xnor U6290 (N_6290,N_5566,N_5860);
nand U6291 (N_6291,N_4963,N_4980);
nor U6292 (N_6292,N_5188,N_5418);
nor U6293 (N_6293,N_5633,N_5226);
and U6294 (N_6294,N_4661,N_5589);
nor U6295 (N_6295,N_4751,N_4769);
and U6296 (N_6296,N_5234,N_4684);
nand U6297 (N_6297,N_5490,N_5995);
nand U6298 (N_6298,N_4911,N_5511);
nand U6299 (N_6299,N_5912,N_5764);
nor U6300 (N_6300,N_5716,N_5762);
and U6301 (N_6301,N_4820,N_5192);
nand U6302 (N_6302,N_5365,N_5825);
xor U6303 (N_6303,N_5273,N_4691);
or U6304 (N_6304,N_5574,N_5300);
nor U6305 (N_6305,N_5679,N_5133);
nand U6306 (N_6306,N_5065,N_4667);
nor U6307 (N_6307,N_5904,N_5356);
nand U6308 (N_6308,N_5450,N_4595);
and U6309 (N_6309,N_4664,N_5181);
or U6310 (N_6310,N_5166,N_4842);
nand U6311 (N_6311,N_5723,N_4649);
and U6312 (N_6312,N_5220,N_5096);
or U6313 (N_6313,N_5974,N_5242);
nand U6314 (N_6314,N_5950,N_4646);
and U6315 (N_6315,N_5301,N_5121);
or U6316 (N_6316,N_5836,N_4946);
or U6317 (N_6317,N_5051,N_5768);
nor U6318 (N_6318,N_4947,N_5411);
and U6319 (N_6319,N_5733,N_5279);
nor U6320 (N_6320,N_5309,N_4500);
xor U6321 (N_6321,N_5368,N_4885);
nand U6322 (N_6322,N_5243,N_5104);
xor U6323 (N_6323,N_5985,N_4604);
nor U6324 (N_6324,N_5256,N_5987);
and U6325 (N_6325,N_5055,N_5090);
nor U6326 (N_6326,N_4869,N_5864);
and U6327 (N_6327,N_4520,N_5853);
nor U6328 (N_6328,N_5796,N_5224);
xnor U6329 (N_6329,N_5592,N_5922);
or U6330 (N_6330,N_4765,N_4708);
nand U6331 (N_6331,N_5395,N_4778);
xor U6332 (N_6332,N_5152,N_4613);
or U6333 (N_6333,N_4614,N_5514);
nand U6334 (N_6334,N_4898,N_5933);
nand U6335 (N_6335,N_4780,N_5410);
xor U6336 (N_6336,N_5294,N_5035);
or U6337 (N_6337,N_4982,N_5030);
and U6338 (N_6338,N_4533,N_5637);
nor U6339 (N_6339,N_4962,N_5980);
or U6340 (N_6340,N_5524,N_5719);
or U6341 (N_6341,N_4938,N_5293);
nor U6342 (N_6342,N_5627,N_5581);
nand U6343 (N_6343,N_5671,N_5505);
and U6344 (N_6344,N_4878,N_5942);
or U6345 (N_6345,N_5878,N_5156);
xnor U6346 (N_6346,N_5134,N_5932);
nand U6347 (N_6347,N_4587,N_5363);
nand U6348 (N_6348,N_5454,N_5827);
nand U6349 (N_6349,N_4992,N_5462);
and U6350 (N_6350,N_5269,N_5014);
and U6351 (N_6351,N_5117,N_4845);
nor U6352 (N_6352,N_4704,N_5731);
nand U6353 (N_6353,N_5771,N_5189);
xnor U6354 (N_6354,N_4642,N_5975);
nor U6355 (N_6355,N_5551,N_4554);
and U6356 (N_6356,N_5163,N_5643);
nor U6357 (N_6357,N_5392,N_4700);
and U6358 (N_6358,N_5676,N_4629);
nand U6359 (N_6359,N_4530,N_5002);
nand U6360 (N_6360,N_4882,N_5005);
nor U6361 (N_6361,N_4717,N_5529);
nor U6362 (N_6362,N_5718,N_4939);
and U6363 (N_6363,N_5941,N_5828);
or U6364 (N_6364,N_4526,N_4610);
xnor U6365 (N_6365,N_5884,N_5434);
nand U6366 (N_6366,N_5544,N_4881);
nand U6367 (N_6367,N_4836,N_5348);
nand U6368 (N_6368,N_4752,N_5698);
and U6369 (N_6369,N_5058,N_4805);
xor U6370 (N_6370,N_5545,N_5543);
nand U6371 (N_6371,N_5889,N_4670);
and U6372 (N_6372,N_4600,N_5803);
xnor U6373 (N_6373,N_5607,N_4631);
xnor U6374 (N_6374,N_5897,N_4549);
xor U6375 (N_6375,N_5409,N_4725);
or U6376 (N_6376,N_4750,N_5082);
xor U6377 (N_6377,N_5756,N_5654);
or U6378 (N_6378,N_5094,N_5374);
and U6379 (N_6379,N_5923,N_5936);
or U6380 (N_6380,N_4936,N_5843);
nor U6381 (N_6381,N_5714,N_5665);
and U6382 (N_6382,N_4656,N_5186);
nand U6383 (N_6383,N_4872,N_5426);
xor U6384 (N_6384,N_4517,N_4933);
nor U6385 (N_6385,N_5779,N_5968);
or U6386 (N_6386,N_4887,N_4926);
nand U6387 (N_6387,N_5263,N_5726);
xor U6388 (N_6388,N_5537,N_5620);
xnor U6389 (N_6389,N_5704,N_4563);
xnor U6390 (N_6390,N_4761,N_5534);
and U6391 (N_6391,N_5022,N_4894);
nor U6392 (N_6392,N_5785,N_4719);
nand U6393 (N_6393,N_5647,N_5443);
or U6394 (N_6394,N_5266,N_4665);
nor U6395 (N_6395,N_5277,N_4970);
and U6396 (N_6396,N_5245,N_5527);
or U6397 (N_6397,N_5850,N_5845);
nor U6398 (N_6398,N_5622,N_4883);
nor U6399 (N_6399,N_5023,N_4916);
and U6400 (N_6400,N_4741,N_4612);
and U6401 (N_6401,N_4834,N_5509);
nand U6402 (N_6402,N_4594,N_5452);
or U6403 (N_6403,N_4810,N_5990);
and U6404 (N_6404,N_5911,N_5453);
and U6405 (N_6405,N_5422,N_5795);
nor U6406 (N_6406,N_5179,N_5867);
nand U6407 (N_6407,N_5930,N_5890);
nor U6408 (N_6408,N_4636,N_5542);
or U6409 (N_6409,N_5686,N_5427);
xor U6410 (N_6410,N_4583,N_4523);
or U6411 (N_6411,N_5473,N_5855);
nand U6412 (N_6412,N_4961,N_4697);
and U6413 (N_6413,N_5198,N_4831);
nand U6414 (N_6414,N_4923,N_5822);
and U6415 (N_6415,N_4973,N_5321);
or U6416 (N_6416,N_4663,N_4809);
or U6417 (N_6417,N_4779,N_5970);
or U6418 (N_6418,N_5057,N_4971);
and U6419 (N_6419,N_5645,N_4641);
and U6420 (N_6420,N_5228,N_4937);
or U6421 (N_6421,N_5447,N_5684);
nand U6422 (N_6422,N_5240,N_5513);
xnor U6423 (N_6423,N_5075,N_5743);
nand U6424 (N_6424,N_5451,N_5799);
xnor U6425 (N_6425,N_5624,N_4941);
or U6426 (N_6426,N_5048,N_4921);
or U6427 (N_6427,N_5608,N_5721);
and U6428 (N_6428,N_4713,N_5267);
nand U6429 (N_6429,N_5238,N_5881);
or U6430 (N_6430,N_5036,N_5246);
nand U6431 (N_6431,N_5488,N_4904);
xor U6432 (N_6432,N_5064,N_5323);
nor U6433 (N_6433,N_5042,N_5322);
nand U6434 (N_6434,N_5861,N_5508);
or U6435 (N_6435,N_4757,N_5067);
nand U6436 (N_6436,N_5781,N_4678);
xnor U6437 (N_6437,N_4860,N_5112);
nand U6438 (N_6438,N_4729,N_5184);
nor U6439 (N_6439,N_5887,N_5705);
nand U6440 (N_6440,N_4685,N_4759);
nor U6441 (N_6441,N_5110,N_4647);
and U6442 (N_6442,N_5739,N_5468);
and U6443 (N_6443,N_5062,N_5960);
or U6444 (N_6444,N_5173,N_4666);
nor U6445 (N_6445,N_5400,N_5583);
xor U6446 (N_6446,N_5713,N_5401);
nand U6447 (N_6447,N_4901,N_5494);
nor U6448 (N_6448,N_5609,N_5311);
nor U6449 (N_6449,N_5312,N_5341);
nand U6450 (N_6450,N_4722,N_4531);
nand U6451 (N_6451,N_5895,N_5214);
xor U6452 (N_6452,N_5105,N_5863);
xnor U6453 (N_6453,N_4633,N_4567);
and U6454 (N_6454,N_5114,N_5297);
nor U6455 (N_6455,N_4746,N_5525);
xnor U6456 (N_6456,N_4893,N_4816);
nor U6457 (N_6457,N_4990,N_4788);
nand U6458 (N_6458,N_4723,N_5384);
and U6459 (N_6459,N_5254,N_5262);
nor U6460 (N_6460,N_5165,N_5241);
or U6461 (N_6461,N_4701,N_4524);
nor U6462 (N_6462,N_4668,N_5711);
xor U6463 (N_6463,N_5539,N_4891);
and U6464 (N_6464,N_5807,N_5010);
or U6465 (N_6465,N_4658,N_5902);
nor U6466 (N_6466,N_4875,N_5037);
or U6467 (N_6467,N_5124,N_5317);
nand U6468 (N_6468,N_5644,N_5709);
nor U6469 (N_6469,N_4505,N_5792);
nand U6470 (N_6470,N_5788,N_5847);
or U6471 (N_6471,N_5034,N_4738);
nand U6472 (N_6472,N_4513,N_4699);
and U6473 (N_6473,N_4900,N_5140);
nand U6474 (N_6474,N_5138,N_4976);
nand U6475 (N_6475,N_4768,N_4611);
and U6476 (N_6476,N_5613,N_5724);
xor U6477 (N_6477,N_5203,N_5914);
xnor U6478 (N_6478,N_5880,N_5106);
xor U6479 (N_6479,N_5466,N_5833);
nor U6480 (N_6480,N_5148,N_5681);
xor U6481 (N_6481,N_5223,N_5888);
or U6482 (N_6482,N_5528,N_5369);
or U6483 (N_6483,N_5628,N_5638);
or U6484 (N_6484,N_5730,N_5419);
xnor U6485 (N_6485,N_4763,N_4637);
nand U6486 (N_6486,N_4827,N_4634);
and U6487 (N_6487,N_4698,N_5893);
nor U6488 (N_6488,N_5894,N_4999);
and U6489 (N_6489,N_5615,N_4521);
xor U6490 (N_6490,N_5153,N_5909);
and U6491 (N_6491,N_5829,N_5934);
and U6492 (N_6492,N_5268,N_5230);
nor U6493 (N_6493,N_4956,N_5801);
nor U6494 (N_6494,N_5800,N_4687);
nor U6495 (N_6495,N_5896,N_4935);
xor U6496 (N_6496,N_4732,N_5576);
xnor U6497 (N_6497,N_4654,N_5877);
xor U6498 (N_6498,N_4912,N_4512);
nor U6499 (N_6499,N_5280,N_5247);
nand U6500 (N_6500,N_5746,N_5000);
nand U6501 (N_6501,N_4807,N_5287);
and U6502 (N_6502,N_5109,N_4588);
and U6503 (N_6503,N_5538,N_5674);
or U6504 (N_6504,N_5856,N_5873);
xor U6505 (N_6505,N_4822,N_4602);
nor U6506 (N_6506,N_5102,N_5834);
nor U6507 (N_6507,N_5021,N_5701);
or U6508 (N_6508,N_5696,N_5449);
nand U6509 (N_6509,N_4925,N_5669);
nor U6510 (N_6510,N_4534,N_5467);
nand U6511 (N_6511,N_5141,N_4945);
nor U6512 (N_6512,N_4731,N_5533);
xnor U6513 (N_6513,N_5977,N_5646);
and U6514 (N_6514,N_5774,N_5445);
xor U6515 (N_6515,N_5071,N_5871);
or U6516 (N_6516,N_5054,N_5630);
xor U6517 (N_6517,N_5264,N_5072);
xor U6518 (N_6518,N_4702,N_5675);
and U6519 (N_6519,N_5160,N_4902);
and U6520 (N_6520,N_5840,N_5789);
and U6521 (N_6521,N_4659,N_5945);
or U6522 (N_6522,N_5077,N_4800);
nor U6523 (N_6523,N_5421,N_5355);
nor U6524 (N_6524,N_4766,N_5404);
nor U6525 (N_6525,N_4532,N_5430);
and U6526 (N_6526,N_5603,N_5947);
xor U6527 (N_6527,N_5883,N_4828);
nor U6528 (N_6528,N_5685,N_5095);
or U6529 (N_6529,N_5284,N_4924);
xnor U6530 (N_6530,N_5125,N_5636);
and U6531 (N_6531,N_4906,N_5907);
nand U6532 (N_6532,N_4981,N_5282);
and U6533 (N_6533,N_5259,N_4991);
nand U6534 (N_6534,N_4838,N_5526);
nand U6535 (N_6535,N_4867,N_5060);
nand U6536 (N_6536,N_5360,N_4706);
nand U6537 (N_6537,N_5732,N_5944);
nand U6538 (N_6538,N_5080,N_4736);
or U6539 (N_6539,N_4975,N_4776);
nor U6540 (N_6540,N_5585,N_5841);
and U6541 (N_6541,N_5142,N_4606);
xnor U6542 (N_6542,N_5170,N_5026);
nor U6543 (N_6543,N_5340,N_5265);
and U6544 (N_6544,N_4590,N_5049);
and U6545 (N_6545,N_5536,N_5521);
or U6546 (N_6546,N_5285,N_5984);
or U6547 (N_6547,N_4504,N_5120);
xor U6548 (N_6548,N_5250,N_5900);
nor U6549 (N_6549,N_5244,N_5345);
nand U6550 (N_6550,N_5503,N_5390);
and U6551 (N_6551,N_5295,N_5197);
nor U6552 (N_6552,N_5978,N_5361);
nand U6553 (N_6553,N_4714,N_4896);
or U6554 (N_6554,N_4985,N_5213);
xnor U6555 (N_6555,N_4903,N_5330);
nor U6556 (N_6556,N_5397,N_5139);
xnor U6557 (N_6557,N_5949,N_5687);
nor U6558 (N_6558,N_5097,N_5391);
and U6559 (N_6559,N_4546,N_5492);
or U6560 (N_6560,N_5329,N_5830);
and U6561 (N_6561,N_4794,N_4994);
xnor U6562 (N_6562,N_4754,N_4813);
or U6563 (N_6563,N_5103,N_5326);
and U6564 (N_6564,N_5351,N_4592);
xor U6565 (N_6565,N_5961,N_5502);
nor U6566 (N_6566,N_5815,N_5193);
xnor U6567 (N_6567,N_5359,N_5692);
xor U6568 (N_6568,N_4762,N_5303);
or U6569 (N_6569,N_5736,N_4675);
nor U6570 (N_6570,N_5621,N_4507);
or U6571 (N_6571,N_5085,N_4735);
and U6572 (N_6572,N_4817,N_5763);
or U6573 (N_6573,N_4709,N_4907);
nor U6574 (N_6574,N_4618,N_5249);
nor U6575 (N_6575,N_4724,N_5248);
and U6576 (N_6576,N_4951,N_5901);
nor U6577 (N_6577,N_5479,N_5442);
and U6578 (N_6578,N_5735,N_5706);
nand U6579 (N_6579,N_5086,N_4988);
nand U6580 (N_6580,N_5231,N_4540);
nor U6581 (N_6581,N_5342,N_5650);
xnor U6582 (N_6582,N_5337,N_5399);
xor U6583 (N_6583,N_5745,N_5939);
xor U6584 (N_6584,N_4728,N_4897);
nand U6585 (N_6585,N_4669,N_4657);
or U6586 (N_6586,N_5996,N_5302);
xor U6587 (N_6587,N_4930,N_5001);
nor U6588 (N_6588,N_4515,N_4758);
and U6589 (N_6589,N_4958,N_4749);
and U6590 (N_6590,N_5370,N_5478);
nand U6591 (N_6591,N_5549,N_4635);
and U6592 (N_6592,N_4632,N_4525);
or U6593 (N_6593,N_5350,N_5019);
nand U6594 (N_6594,N_5281,N_5759);
nand U6595 (N_6595,N_4652,N_5306);
and U6596 (N_6596,N_4793,N_5517);
nor U6597 (N_6597,N_4582,N_5916);
nor U6598 (N_6598,N_4857,N_4739);
xnor U6599 (N_6599,N_5956,N_5772);
nand U6600 (N_6600,N_5851,N_4855);
nand U6601 (N_6601,N_4651,N_5483);
nor U6602 (N_6602,N_5389,N_5320);
nand U6603 (N_6603,N_5149,N_5837);
nor U6604 (N_6604,N_5412,N_5168);
nor U6605 (N_6605,N_4934,N_5623);
nor U6606 (N_6606,N_5346,N_5994);
or U6607 (N_6607,N_4871,N_4850);
nand U6608 (N_6608,N_4795,N_5131);
xor U6609 (N_6609,N_5432,N_5332);
xor U6610 (N_6610,N_4585,N_4949);
or U6611 (N_6611,N_5741,N_5255);
or U6612 (N_6612,N_4811,N_5237);
nor U6613 (N_6613,N_4571,N_5472);
nand U6614 (N_6614,N_5239,N_4889);
nand U6615 (N_6615,N_4876,N_5997);
nand U6616 (N_6616,N_5215,N_4626);
and U6617 (N_6617,N_5813,N_5319);
or U6618 (N_6618,N_5761,N_5816);
nor U6619 (N_6619,N_5386,N_5629);
nor U6620 (N_6620,N_5865,N_4561);
nor U6621 (N_6621,N_5811,N_5558);
or U6622 (N_6622,N_5913,N_5972);
and U6623 (N_6623,N_5433,N_5499);
or U6624 (N_6624,N_4693,N_5700);
or U6625 (N_6625,N_5918,N_5758);
nand U6626 (N_6626,N_5464,N_5707);
and U6627 (N_6627,N_4781,N_5740);
and U6628 (N_6628,N_4977,N_5087);
or U6629 (N_6629,N_5680,N_5876);
or U6630 (N_6630,N_4712,N_5858);
nor U6631 (N_6631,N_4978,N_4848);
and U6632 (N_6632,N_5151,N_5437);
xor U6633 (N_6633,N_4660,N_5682);
and U6634 (N_6634,N_5053,N_4950);
nand U6635 (N_6635,N_4696,N_5747);
xnor U6636 (N_6636,N_5653,N_4797);
or U6637 (N_6637,N_5041,N_5729);
nor U6638 (N_6638,N_4858,N_4965);
and U6639 (N_6639,N_5413,N_5776);
and U6640 (N_6640,N_5157,N_5727);
and U6641 (N_6641,N_5435,N_5408);
or U6642 (N_6642,N_5523,N_5396);
xor U6643 (N_6643,N_5018,N_4862);
or U6644 (N_6644,N_5712,N_5940);
xor U6645 (N_6645,N_5463,N_5336);
xor U6646 (N_6646,N_4542,N_5567);
and U6647 (N_6647,N_5313,N_4555);
xnor U6648 (N_6648,N_5971,N_4671);
or U6649 (N_6649,N_5986,N_4955);
or U6650 (N_6650,N_5892,N_5225);
nor U6651 (N_6651,N_5991,N_4989);
nor U6652 (N_6652,N_5236,N_5708);
nor U6653 (N_6653,N_4705,N_4573);
nor U6654 (N_6654,N_5066,N_5286);
and U6655 (N_6655,N_5857,N_4974);
nand U6656 (N_6656,N_5981,N_5316);
and U6657 (N_6657,N_5898,N_5143);
or U6658 (N_6658,N_4832,N_4680);
or U6659 (N_6659,N_5612,N_5921);
and U6660 (N_6660,N_5738,N_5842);
xor U6661 (N_6661,N_5088,N_4952);
nand U6662 (N_6662,N_5814,N_5327);
nor U6663 (N_6663,N_5496,N_5958);
xor U6664 (N_6664,N_4840,N_4682);
nor U6665 (N_6665,N_4960,N_4726);
xor U6666 (N_6666,N_4756,N_5586);
nor U6667 (N_6667,N_4599,N_5750);
nand U6668 (N_6668,N_4672,N_4711);
and U6669 (N_6669,N_4913,N_5964);
nand U6670 (N_6670,N_5235,N_4747);
and U6671 (N_6671,N_5448,N_5611);
nand U6672 (N_6672,N_5693,N_5798);
xor U6673 (N_6673,N_4799,N_5651);
xnor U6674 (N_6674,N_5436,N_5666);
nor U6675 (N_6675,N_5854,N_4621);
and U6676 (N_6676,N_5497,N_5575);
nand U6677 (N_6677,N_4578,N_4969);
nand U6678 (N_6678,N_4603,N_4718);
nor U6679 (N_6679,N_5810,N_5561);
and U6680 (N_6680,N_5063,N_5640);
and U6681 (N_6681,N_5584,N_5475);
xor U6682 (N_6682,N_5652,N_4852);
nor U6683 (N_6683,N_4644,N_5078);
and U6684 (N_6684,N_5618,N_5587);
xor U6685 (N_6685,N_5594,N_5128);
and U6686 (N_6686,N_5461,N_4727);
or U6687 (N_6687,N_4597,N_5520);
and U6688 (N_6688,N_4812,N_4787);
nand U6689 (N_6689,N_4790,N_4628);
or U6690 (N_6690,N_5920,N_5147);
xnor U6691 (N_6691,N_5310,N_5158);
and U6692 (N_6692,N_5554,N_4509);
nor U6693 (N_6693,N_5531,N_4734);
and U6694 (N_6694,N_5218,N_4996);
nor U6695 (N_6695,N_5824,N_5444);
or U6696 (N_6696,N_5967,N_5573);
nand U6697 (N_6697,N_5495,N_5335);
xor U6698 (N_6698,N_5578,N_4742);
xor U6699 (N_6699,N_5664,N_5872);
xnor U6700 (N_6700,N_5656,N_4957);
xnor U6701 (N_6701,N_5362,N_4879);
and U6702 (N_6702,N_5381,N_4833);
or U6703 (N_6703,N_4688,N_5178);
and U6704 (N_6704,N_5677,N_5908);
and U6705 (N_6705,N_5519,N_5672);
nor U6706 (N_6706,N_5347,N_4617);
and U6707 (N_6707,N_5027,N_5354);
xnor U6708 (N_6708,N_4899,N_5099);
and U6709 (N_6709,N_4516,N_4914);
and U6710 (N_6710,N_4839,N_5838);
nor U6711 (N_6711,N_5604,N_5331);
and U6712 (N_6712,N_5695,N_5839);
xor U6713 (N_6713,N_5364,N_5797);
xnor U6714 (N_6714,N_4854,N_4640);
nand U6715 (N_6715,N_5334,N_5372);
nor U6716 (N_6716,N_5383,N_5821);
nand U6717 (N_6717,N_5925,N_4547);
and U6718 (N_6718,N_4890,N_5045);
or U6719 (N_6719,N_5606,N_5290);
and U6720 (N_6720,N_5658,N_4650);
xnor U6721 (N_6721,N_5642,N_5092);
nand U6722 (N_6722,N_5101,N_5056);
and U6723 (N_6723,N_5515,N_4625);
or U6724 (N_6724,N_4703,N_5164);
nor U6725 (N_6725,N_5924,N_5625);
or U6726 (N_6726,N_4518,N_5025);
xnor U6727 (N_6727,N_5191,N_5081);
or U6728 (N_6728,N_5634,N_4801);
nand U6729 (N_6729,N_5780,N_4544);
or U6730 (N_6730,N_4940,N_5831);
nand U6731 (N_6731,N_5662,N_5069);
nand U6732 (N_6732,N_5050,N_4503);
xor U6733 (N_6733,N_5999,N_5879);
nand U6734 (N_6734,N_4873,N_5375);
nor U6735 (N_6735,N_5946,N_5076);
or U6736 (N_6736,N_5605,N_5187);
nor U6737 (N_6737,N_5145,N_5122);
nand U6738 (N_6738,N_5632,N_4620);
and U6739 (N_6739,N_5272,N_5009);
nor U6740 (N_6740,N_5703,N_5885);
xnor U6741 (N_6741,N_5275,N_5820);
and U6742 (N_6742,N_4676,N_4849);
and U6743 (N_6743,N_5602,N_4767);
or U6744 (N_6744,N_5135,N_5915);
or U6745 (N_6745,N_4953,N_4919);
or U6746 (N_6746,N_5177,N_4826);
nor U6747 (N_6747,N_4558,N_5487);
nor U6748 (N_6748,N_5979,N_5678);
and U6749 (N_6749,N_5927,N_4720);
and U6750 (N_6750,N_5844,N_4704);
xnor U6751 (N_6751,N_5255,N_4526);
nor U6752 (N_6752,N_5059,N_4517);
xor U6753 (N_6753,N_5942,N_5006);
or U6754 (N_6754,N_4788,N_5324);
nor U6755 (N_6755,N_4913,N_5441);
nor U6756 (N_6756,N_5278,N_4952);
xor U6757 (N_6757,N_5449,N_5992);
and U6758 (N_6758,N_4635,N_5195);
nand U6759 (N_6759,N_5294,N_5589);
xnor U6760 (N_6760,N_5711,N_4720);
nor U6761 (N_6761,N_5946,N_5580);
xor U6762 (N_6762,N_5914,N_5553);
nand U6763 (N_6763,N_5052,N_5175);
or U6764 (N_6764,N_4863,N_5548);
or U6765 (N_6765,N_5410,N_5629);
nor U6766 (N_6766,N_4960,N_5816);
xnor U6767 (N_6767,N_4539,N_5022);
and U6768 (N_6768,N_4556,N_4790);
nor U6769 (N_6769,N_5642,N_5227);
and U6770 (N_6770,N_5676,N_5540);
nand U6771 (N_6771,N_5104,N_5136);
and U6772 (N_6772,N_5864,N_5973);
and U6773 (N_6773,N_4650,N_5338);
and U6774 (N_6774,N_5103,N_5521);
nand U6775 (N_6775,N_5489,N_4541);
nand U6776 (N_6776,N_4956,N_5097);
nor U6777 (N_6777,N_5984,N_4525);
nand U6778 (N_6778,N_4929,N_4738);
and U6779 (N_6779,N_4725,N_5432);
nand U6780 (N_6780,N_4834,N_5650);
xnor U6781 (N_6781,N_4703,N_5812);
nor U6782 (N_6782,N_5039,N_5023);
xor U6783 (N_6783,N_4734,N_5459);
xnor U6784 (N_6784,N_5191,N_4794);
or U6785 (N_6785,N_5122,N_4640);
and U6786 (N_6786,N_5386,N_5930);
nand U6787 (N_6787,N_4736,N_4536);
nor U6788 (N_6788,N_5131,N_5225);
nor U6789 (N_6789,N_4791,N_5234);
nor U6790 (N_6790,N_5003,N_5085);
nor U6791 (N_6791,N_5331,N_5625);
or U6792 (N_6792,N_5989,N_5115);
or U6793 (N_6793,N_4643,N_5552);
xnor U6794 (N_6794,N_5423,N_5995);
and U6795 (N_6795,N_4927,N_4731);
nor U6796 (N_6796,N_5249,N_5368);
nor U6797 (N_6797,N_5660,N_5150);
nor U6798 (N_6798,N_4797,N_4709);
or U6799 (N_6799,N_4564,N_5558);
or U6800 (N_6800,N_5446,N_5411);
and U6801 (N_6801,N_5751,N_5806);
xor U6802 (N_6802,N_5530,N_4733);
nand U6803 (N_6803,N_4735,N_5709);
nand U6804 (N_6804,N_5500,N_5263);
nand U6805 (N_6805,N_5595,N_4847);
and U6806 (N_6806,N_5157,N_4910);
or U6807 (N_6807,N_5054,N_4531);
xnor U6808 (N_6808,N_4979,N_4746);
and U6809 (N_6809,N_5273,N_5185);
or U6810 (N_6810,N_5973,N_5913);
nor U6811 (N_6811,N_5227,N_4813);
and U6812 (N_6812,N_5008,N_5213);
and U6813 (N_6813,N_4619,N_5731);
nand U6814 (N_6814,N_4983,N_5565);
or U6815 (N_6815,N_4713,N_5706);
or U6816 (N_6816,N_5454,N_5258);
xor U6817 (N_6817,N_5134,N_5276);
and U6818 (N_6818,N_5921,N_4773);
or U6819 (N_6819,N_5134,N_5046);
and U6820 (N_6820,N_5594,N_5273);
or U6821 (N_6821,N_5714,N_4880);
xor U6822 (N_6822,N_4957,N_4730);
and U6823 (N_6823,N_5401,N_5179);
and U6824 (N_6824,N_5568,N_4853);
or U6825 (N_6825,N_4779,N_5163);
or U6826 (N_6826,N_5208,N_5062);
xnor U6827 (N_6827,N_5285,N_4556);
nor U6828 (N_6828,N_5262,N_5581);
xnor U6829 (N_6829,N_5122,N_4772);
and U6830 (N_6830,N_5539,N_5723);
or U6831 (N_6831,N_5087,N_4613);
nor U6832 (N_6832,N_5269,N_5108);
or U6833 (N_6833,N_5806,N_5074);
xor U6834 (N_6834,N_5972,N_4790);
xnor U6835 (N_6835,N_5983,N_5240);
or U6836 (N_6836,N_5030,N_4881);
and U6837 (N_6837,N_5672,N_5983);
or U6838 (N_6838,N_5408,N_5175);
or U6839 (N_6839,N_5906,N_5664);
and U6840 (N_6840,N_5529,N_5540);
nand U6841 (N_6841,N_5406,N_5973);
and U6842 (N_6842,N_5660,N_5407);
xnor U6843 (N_6843,N_4886,N_5760);
xnor U6844 (N_6844,N_5625,N_4507);
nor U6845 (N_6845,N_4683,N_5771);
and U6846 (N_6846,N_4711,N_5796);
or U6847 (N_6847,N_5541,N_4560);
nand U6848 (N_6848,N_4983,N_4670);
or U6849 (N_6849,N_5864,N_5995);
nor U6850 (N_6850,N_5946,N_5813);
nor U6851 (N_6851,N_4810,N_4866);
nand U6852 (N_6852,N_5377,N_4855);
or U6853 (N_6853,N_4540,N_5100);
and U6854 (N_6854,N_5612,N_4732);
or U6855 (N_6855,N_4842,N_5876);
xnor U6856 (N_6856,N_5846,N_5818);
and U6857 (N_6857,N_5846,N_5249);
xor U6858 (N_6858,N_4831,N_4646);
or U6859 (N_6859,N_5855,N_5505);
or U6860 (N_6860,N_5679,N_4812);
xor U6861 (N_6861,N_5517,N_5980);
nor U6862 (N_6862,N_5155,N_5841);
xnor U6863 (N_6863,N_4894,N_4791);
xnor U6864 (N_6864,N_4931,N_5295);
or U6865 (N_6865,N_5351,N_4937);
nor U6866 (N_6866,N_4502,N_4611);
or U6867 (N_6867,N_5089,N_5433);
nand U6868 (N_6868,N_4770,N_4769);
and U6869 (N_6869,N_5768,N_4705);
or U6870 (N_6870,N_4681,N_5733);
nand U6871 (N_6871,N_5612,N_4723);
and U6872 (N_6872,N_5550,N_5140);
nor U6873 (N_6873,N_4996,N_5144);
or U6874 (N_6874,N_5388,N_4724);
nand U6875 (N_6875,N_4910,N_4599);
nand U6876 (N_6876,N_5290,N_4862);
nor U6877 (N_6877,N_4761,N_5569);
xor U6878 (N_6878,N_4894,N_4656);
nand U6879 (N_6879,N_5803,N_5456);
xor U6880 (N_6880,N_5728,N_4805);
nor U6881 (N_6881,N_4598,N_4967);
nand U6882 (N_6882,N_5450,N_4943);
nand U6883 (N_6883,N_5859,N_5483);
nor U6884 (N_6884,N_5198,N_5926);
nor U6885 (N_6885,N_5755,N_5174);
and U6886 (N_6886,N_5564,N_5028);
and U6887 (N_6887,N_5352,N_5751);
or U6888 (N_6888,N_5069,N_5421);
or U6889 (N_6889,N_5981,N_5845);
and U6890 (N_6890,N_5598,N_5153);
nand U6891 (N_6891,N_5431,N_5178);
and U6892 (N_6892,N_4597,N_4770);
nand U6893 (N_6893,N_5152,N_5260);
xnor U6894 (N_6894,N_4790,N_5307);
nor U6895 (N_6895,N_5078,N_4796);
nor U6896 (N_6896,N_5676,N_5365);
nor U6897 (N_6897,N_4840,N_5965);
and U6898 (N_6898,N_4879,N_4841);
and U6899 (N_6899,N_5453,N_4654);
xnor U6900 (N_6900,N_4983,N_5624);
nand U6901 (N_6901,N_5726,N_5272);
nor U6902 (N_6902,N_4937,N_5475);
and U6903 (N_6903,N_5807,N_4552);
nand U6904 (N_6904,N_5077,N_5092);
or U6905 (N_6905,N_5759,N_5262);
nand U6906 (N_6906,N_5009,N_4674);
or U6907 (N_6907,N_4827,N_5499);
or U6908 (N_6908,N_4846,N_5795);
or U6909 (N_6909,N_5638,N_5803);
or U6910 (N_6910,N_5688,N_4510);
or U6911 (N_6911,N_5371,N_5993);
nor U6912 (N_6912,N_5530,N_4549);
nand U6913 (N_6913,N_4856,N_5840);
nand U6914 (N_6914,N_5878,N_4688);
xnor U6915 (N_6915,N_4777,N_5408);
nor U6916 (N_6916,N_4586,N_4796);
or U6917 (N_6917,N_4822,N_5552);
xor U6918 (N_6918,N_5343,N_4664);
nand U6919 (N_6919,N_5920,N_5498);
or U6920 (N_6920,N_5202,N_5223);
or U6921 (N_6921,N_5974,N_4694);
xor U6922 (N_6922,N_5043,N_5083);
xor U6923 (N_6923,N_5905,N_4518);
or U6924 (N_6924,N_4624,N_5936);
nor U6925 (N_6925,N_5132,N_4757);
nand U6926 (N_6926,N_5842,N_5245);
and U6927 (N_6927,N_5524,N_4982);
nand U6928 (N_6928,N_5518,N_5873);
nor U6929 (N_6929,N_5247,N_5849);
xnor U6930 (N_6930,N_5478,N_5458);
xor U6931 (N_6931,N_4608,N_5354);
nor U6932 (N_6932,N_5886,N_5255);
and U6933 (N_6933,N_4843,N_4782);
xnor U6934 (N_6934,N_4947,N_5695);
and U6935 (N_6935,N_4653,N_5180);
xor U6936 (N_6936,N_5302,N_5283);
nor U6937 (N_6937,N_5501,N_4944);
nor U6938 (N_6938,N_5048,N_5379);
and U6939 (N_6939,N_5265,N_5866);
nand U6940 (N_6940,N_4717,N_5384);
and U6941 (N_6941,N_5903,N_4601);
and U6942 (N_6942,N_5677,N_5982);
and U6943 (N_6943,N_5412,N_4712);
nand U6944 (N_6944,N_4666,N_5539);
and U6945 (N_6945,N_4973,N_4955);
xnor U6946 (N_6946,N_5262,N_5526);
or U6947 (N_6947,N_5990,N_5035);
xnor U6948 (N_6948,N_5771,N_5669);
and U6949 (N_6949,N_5575,N_5686);
nor U6950 (N_6950,N_5795,N_5705);
xnor U6951 (N_6951,N_5440,N_5892);
and U6952 (N_6952,N_5068,N_5427);
and U6953 (N_6953,N_5030,N_4669);
or U6954 (N_6954,N_5804,N_4824);
and U6955 (N_6955,N_5582,N_4557);
and U6956 (N_6956,N_5783,N_5114);
xor U6957 (N_6957,N_5133,N_4918);
xor U6958 (N_6958,N_5364,N_5528);
nor U6959 (N_6959,N_5620,N_5521);
xnor U6960 (N_6960,N_4730,N_5712);
nand U6961 (N_6961,N_5590,N_4756);
nor U6962 (N_6962,N_4883,N_5429);
and U6963 (N_6963,N_5751,N_5693);
xor U6964 (N_6964,N_5679,N_4993);
nor U6965 (N_6965,N_4926,N_5398);
nor U6966 (N_6966,N_5395,N_5137);
and U6967 (N_6967,N_5378,N_5373);
nand U6968 (N_6968,N_5138,N_5855);
nand U6969 (N_6969,N_5169,N_5706);
nor U6970 (N_6970,N_5638,N_5766);
and U6971 (N_6971,N_4655,N_5524);
and U6972 (N_6972,N_5333,N_5912);
and U6973 (N_6973,N_5157,N_5505);
nor U6974 (N_6974,N_5792,N_5061);
xnor U6975 (N_6975,N_5970,N_4986);
xor U6976 (N_6976,N_5391,N_5703);
or U6977 (N_6977,N_5615,N_5222);
nand U6978 (N_6978,N_4603,N_4561);
nand U6979 (N_6979,N_5299,N_5256);
nand U6980 (N_6980,N_4610,N_5582);
and U6981 (N_6981,N_5722,N_5301);
nand U6982 (N_6982,N_5105,N_5601);
and U6983 (N_6983,N_5484,N_5664);
nand U6984 (N_6984,N_5396,N_5123);
nand U6985 (N_6985,N_5000,N_5493);
nor U6986 (N_6986,N_4766,N_4657);
nor U6987 (N_6987,N_4770,N_4621);
xnor U6988 (N_6988,N_5546,N_4578);
nand U6989 (N_6989,N_5413,N_5742);
xnor U6990 (N_6990,N_4710,N_5936);
nor U6991 (N_6991,N_5292,N_4805);
and U6992 (N_6992,N_5708,N_5387);
xor U6993 (N_6993,N_5641,N_5250);
or U6994 (N_6994,N_5662,N_5638);
and U6995 (N_6995,N_5490,N_5222);
nor U6996 (N_6996,N_5717,N_5003);
nor U6997 (N_6997,N_5212,N_5687);
xor U6998 (N_6998,N_4852,N_5756);
xnor U6999 (N_6999,N_4671,N_5538);
nand U7000 (N_7000,N_4671,N_5486);
nand U7001 (N_7001,N_4707,N_5171);
nand U7002 (N_7002,N_4736,N_5845);
nand U7003 (N_7003,N_5848,N_4730);
nor U7004 (N_7004,N_5496,N_4567);
or U7005 (N_7005,N_4950,N_5133);
and U7006 (N_7006,N_4502,N_5084);
and U7007 (N_7007,N_4744,N_4882);
and U7008 (N_7008,N_5844,N_5886);
nand U7009 (N_7009,N_4755,N_5606);
nor U7010 (N_7010,N_5938,N_4964);
and U7011 (N_7011,N_5529,N_5259);
or U7012 (N_7012,N_5686,N_5023);
or U7013 (N_7013,N_4635,N_5232);
nand U7014 (N_7014,N_4729,N_5024);
and U7015 (N_7015,N_5105,N_4951);
and U7016 (N_7016,N_5510,N_5355);
nor U7017 (N_7017,N_4778,N_5780);
nor U7018 (N_7018,N_4794,N_4808);
nor U7019 (N_7019,N_5317,N_5327);
xor U7020 (N_7020,N_4842,N_4506);
xnor U7021 (N_7021,N_4671,N_5956);
nor U7022 (N_7022,N_5576,N_5883);
or U7023 (N_7023,N_5696,N_5477);
or U7024 (N_7024,N_5739,N_5384);
and U7025 (N_7025,N_5881,N_4938);
nand U7026 (N_7026,N_5920,N_4843);
xor U7027 (N_7027,N_5093,N_5606);
nand U7028 (N_7028,N_5769,N_4890);
nor U7029 (N_7029,N_5402,N_5817);
xnor U7030 (N_7030,N_5531,N_4739);
nand U7031 (N_7031,N_5917,N_4966);
xnor U7032 (N_7032,N_4589,N_5896);
and U7033 (N_7033,N_5535,N_4627);
or U7034 (N_7034,N_5289,N_5423);
nand U7035 (N_7035,N_4865,N_4561);
nand U7036 (N_7036,N_5681,N_5308);
xor U7037 (N_7037,N_4579,N_5922);
or U7038 (N_7038,N_5843,N_5584);
nand U7039 (N_7039,N_5211,N_4572);
nand U7040 (N_7040,N_4942,N_5864);
or U7041 (N_7041,N_4857,N_5364);
or U7042 (N_7042,N_5518,N_5724);
and U7043 (N_7043,N_5839,N_4686);
and U7044 (N_7044,N_4862,N_5359);
and U7045 (N_7045,N_5945,N_4944);
nor U7046 (N_7046,N_5690,N_4681);
nor U7047 (N_7047,N_5296,N_5824);
xnor U7048 (N_7048,N_5224,N_5847);
and U7049 (N_7049,N_5498,N_5999);
or U7050 (N_7050,N_5437,N_4732);
nor U7051 (N_7051,N_5717,N_4869);
or U7052 (N_7052,N_5099,N_5640);
xnor U7053 (N_7053,N_5908,N_5400);
nor U7054 (N_7054,N_4523,N_5247);
xor U7055 (N_7055,N_5447,N_5965);
nand U7056 (N_7056,N_5000,N_5357);
or U7057 (N_7057,N_5390,N_5688);
or U7058 (N_7058,N_4937,N_5374);
or U7059 (N_7059,N_4558,N_5281);
or U7060 (N_7060,N_5907,N_5352);
xor U7061 (N_7061,N_5705,N_4956);
nand U7062 (N_7062,N_5583,N_5899);
and U7063 (N_7063,N_4919,N_5789);
nor U7064 (N_7064,N_5214,N_5743);
nand U7065 (N_7065,N_4620,N_5210);
and U7066 (N_7066,N_4653,N_5833);
and U7067 (N_7067,N_5178,N_4939);
nor U7068 (N_7068,N_5874,N_5617);
nand U7069 (N_7069,N_4634,N_5351);
xnor U7070 (N_7070,N_5171,N_5874);
and U7071 (N_7071,N_4842,N_4826);
xnor U7072 (N_7072,N_4759,N_5105);
and U7073 (N_7073,N_5958,N_4933);
or U7074 (N_7074,N_5155,N_4743);
nand U7075 (N_7075,N_5988,N_5054);
xor U7076 (N_7076,N_4571,N_4618);
nand U7077 (N_7077,N_5393,N_5954);
xnor U7078 (N_7078,N_5763,N_5631);
nor U7079 (N_7079,N_5484,N_4836);
or U7080 (N_7080,N_5441,N_4670);
nand U7081 (N_7081,N_5530,N_5946);
xor U7082 (N_7082,N_5761,N_4571);
nor U7083 (N_7083,N_5700,N_5482);
nor U7084 (N_7084,N_5477,N_5995);
nor U7085 (N_7085,N_5122,N_5630);
nand U7086 (N_7086,N_4878,N_5248);
nand U7087 (N_7087,N_4663,N_5362);
nor U7088 (N_7088,N_5314,N_5519);
or U7089 (N_7089,N_4990,N_5902);
or U7090 (N_7090,N_5143,N_5328);
and U7091 (N_7091,N_5263,N_4837);
xnor U7092 (N_7092,N_5376,N_5137);
or U7093 (N_7093,N_4566,N_5323);
and U7094 (N_7094,N_5028,N_4545);
or U7095 (N_7095,N_4692,N_5784);
nor U7096 (N_7096,N_5799,N_5092);
or U7097 (N_7097,N_4595,N_5426);
xor U7098 (N_7098,N_5128,N_5373);
or U7099 (N_7099,N_5090,N_5404);
nor U7100 (N_7100,N_5567,N_5937);
nor U7101 (N_7101,N_5974,N_5984);
nand U7102 (N_7102,N_4656,N_5808);
or U7103 (N_7103,N_5857,N_4726);
xnor U7104 (N_7104,N_4748,N_5514);
nand U7105 (N_7105,N_5946,N_5607);
nor U7106 (N_7106,N_5929,N_4947);
and U7107 (N_7107,N_5014,N_4696);
or U7108 (N_7108,N_5052,N_4650);
nor U7109 (N_7109,N_5604,N_5698);
nor U7110 (N_7110,N_4624,N_5171);
nand U7111 (N_7111,N_5269,N_4603);
xnor U7112 (N_7112,N_5872,N_5938);
or U7113 (N_7113,N_5535,N_4611);
nor U7114 (N_7114,N_4589,N_5536);
or U7115 (N_7115,N_5149,N_5758);
or U7116 (N_7116,N_5321,N_4801);
and U7117 (N_7117,N_5796,N_5639);
nor U7118 (N_7118,N_5747,N_5703);
xnor U7119 (N_7119,N_5960,N_5355);
or U7120 (N_7120,N_5151,N_4758);
or U7121 (N_7121,N_5525,N_5514);
xor U7122 (N_7122,N_4810,N_4697);
xnor U7123 (N_7123,N_5677,N_5324);
and U7124 (N_7124,N_5814,N_5513);
and U7125 (N_7125,N_4603,N_5669);
or U7126 (N_7126,N_5918,N_5704);
xor U7127 (N_7127,N_4747,N_5089);
nor U7128 (N_7128,N_5382,N_4725);
nor U7129 (N_7129,N_4905,N_5657);
nand U7130 (N_7130,N_5044,N_5482);
xor U7131 (N_7131,N_5060,N_5559);
nand U7132 (N_7132,N_5033,N_5242);
nor U7133 (N_7133,N_5639,N_4604);
and U7134 (N_7134,N_4561,N_5339);
xor U7135 (N_7135,N_4743,N_5877);
and U7136 (N_7136,N_5069,N_4895);
and U7137 (N_7137,N_5805,N_4541);
xnor U7138 (N_7138,N_4932,N_5995);
nor U7139 (N_7139,N_4636,N_5347);
nand U7140 (N_7140,N_5412,N_5748);
nand U7141 (N_7141,N_4658,N_5497);
and U7142 (N_7142,N_5295,N_4530);
or U7143 (N_7143,N_5298,N_5568);
nor U7144 (N_7144,N_5297,N_5905);
xor U7145 (N_7145,N_5831,N_5000);
nand U7146 (N_7146,N_4695,N_5743);
and U7147 (N_7147,N_5882,N_4839);
nand U7148 (N_7148,N_4979,N_5174);
and U7149 (N_7149,N_5382,N_4632);
or U7150 (N_7150,N_4509,N_4653);
xor U7151 (N_7151,N_4551,N_5929);
or U7152 (N_7152,N_5201,N_5130);
or U7153 (N_7153,N_4835,N_5380);
nor U7154 (N_7154,N_5870,N_4958);
xor U7155 (N_7155,N_5796,N_5631);
and U7156 (N_7156,N_5711,N_5217);
xnor U7157 (N_7157,N_5980,N_5233);
nand U7158 (N_7158,N_4757,N_5296);
nand U7159 (N_7159,N_4820,N_5564);
or U7160 (N_7160,N_5788,N_4557);
or U7161 (N_7161,N_5869,N_5311);
nor U7162 (N_7162,N_4988,N_4655);
nor U7163 (N_7163,N_5523,N_5383);
or U7164 (N_7164,N_5827,N_5931);
nand U7165 (N_7165,N_5942,N_5753);
nor U7166 (N_7166,N_5860,N_4990);
nand U7167 (N_7167,N_5227,N_5947);
nor U7168 (N_7168,N_5777,N_4526);
xor U7169 (N_7169,N_4536,N_4912);
and U7170 (N_7170,N_5428,N_5746);
and U7171 (N_7171,N_5494,N_5763);
nor U7172 (N_7172,N_5464,N_5951);
nor U7173 (N_7173,N_4850,N_5386);
or U7174 (N_7174,N_5533,N_4586);
xor U7175 (N_7175,N_5601,N_4501);
or U7176 (N_7176,N_5540,N_4656);
or U7177 (N_7177,N_5082,N_4548);
xnor U7178 (N_7178,N_4711,N_5560);
nand U7179 (N_7179,N_5735,N_4768);
or U7180 (N_7180,N_5539,N_5022);
or U7181 (N_7181,N_4778,N_4590);
or U7182 (N_7182,N_5137,N_5825);
xnor U7183 (N_7183,N_5559,N_5087);
xnor U7184 (N_7184,N_5096,N_5117);
xor U7185 (N_7185,N_5375,N_5171);
nand U7186 (N_7186,N_4965,N_4799);
xor U7187 (N_7187,N_5654,N_5018);
and U7188 (N_7188,N_5879,N_5769);
or U7189 (N_7189,N_5545,N_5458);
or U7190 (N_7190,N_5532,N_5854);
nor U7191 (N_7191,N_5859,N_4515);
nand U7192 (N_7192,N_4759,N_5159);
nor U7193 (N_7193,N_5532,N_5398);
xor U7194 (N_7194,N_5938,N_5758);
and U7195 (N_7195,N_5388,N_4587);
nor U7196 (N_7196,N_4575,N_5811);
xor U7197 (N_7197,N_5478,N_5571);
nand U7198 (N_7198,N_5018,N_5267);
xnor U7199 (N_7199,N_5951,N_5150);
nand U7200 (N_7200,N_4872,N_5592);
nor U7201 (N_7201,N_5029,N_4660);
xnor U7202 (N_7202,N_5249,N_5606);
nor U7203 (N_7203,N_4854,N_4990);
nor U7204 (N_7204,N_5756,N_4708);
nor U7205 (N_7205,N_4714,N_5353);
or U7206 (N_7206,N_4829,N_5030);
xnor U7207 (N_7207,N_4731,N_5809);
nand U7208 (N_7208,N_4821,N_4894);
xnor U7209 (N_7209,N_5569,N_5527);
xnor U7210 (N_7210,N_5467,N_4621);
nand U7211 (N_7211,N_5681,N_5668);
or U7212 (N_7212,N_5154,N_4763);
nor U7213 (N_7213,N_5287,N_5355);
xor U7214 (N_7214,N_5923,N_5738);
nor U7215 (N_7215,N_4849,N_4781);
and U7216 (N_7216,N_5259,N_5716);
nor U7217 (N_7217,N_5810,N_5495);
nand U7218 (N_7218,N_5696,N_5912);
nor U7219 (N_7219,N_5619,N_5013);
nand U7220 (N_7220,N_5316,N_5060);
nand U7221 (N_7221,N_4982,N_5335);
nand U7222 (N_7222,N_5865,N_5725);
or U7223 (N_7223,N_5313,N_5044);
nand U7224 (N_7224,N_5747,N_5850);
nor U7225 (N_7225,N_5854,N_5539);
nand U7226 (N_7226,N_5521,N_5955);
or U7227 (N_7227,N_5359,N_4790);
nand U7228 (N_7228,N_4713,N_5274);
and U7229 (N_7229,N_5011,N_4809);
nor U7230 (N_7230,N_5327,N_5444);
or U7231 (N_7231,N_4508,N_5411);
and U7232 (N_7232,N_4992,N_4902);
nand U7233 (N_7233,N_5829,N_5029);
nand U7234 (N_7234,N_5089,N_5451);
and U7235 (N_7235,N_5388,N_5507);
nor U7236 (N_7236,N_5824,N_4840);
nor U7237 (N_7237,N_4920,N_4885);
nand U7238 (N_7238,N_5803,N_4927);
nor U7239 (N_7239,N_5052,N_5717);
nand U7240 (N_7240,N_5010,N_5026);
or U7241 (N_7241,N_5521,N_5823);
nand U7242 (N_7242,N_4903,N_5510);
and U7243 (N_7243,N_4844,N_5594);
or U7244 (N_7244,N_4758,N_5722);
nand U7245 (N_7245,N_4519,N_5182);
nand U7246 (N_7246,N_5795,N_4748);
xor U7247 (N_7247,N_5020,N_5922);
or U7248 (N_7248,N_5632,N_5769);
or U7249 (N_7249,N_4675,N_4571);
nand U7250 (N_7250,N_4884,N_4990);
xnor U7251 (N_7251,N_4901,N_5521);
nand U7252 (N_7252,N_5590,N_5793);
nor U7253 (N_7253,N_4593,N_5519);
and U7254 (N_7254,N_5579,N_5950);
or U7255 (N_7255,N_5417,N_5924);
xnor U7256 (N_7256,N_5828,N_5452);
and U7257 (N_7257,N_4679,N_4857);
nand U7258 (N_7258,N_5786,N_5092);
and U7259 (N_7259,N_4804,N_4575);
nor U7260 (N_7260,N_5257,N_5379);
and U7261 (N_7261,N_5441,N_5903);
and U7262 (N_7262,N_4751,N_4538);
xor U7263 (N_7263,N_5995,N_5349);
and U7264 (N_7264,N_5692,N_4674);
and U7265 (N_7265,N_5993,N_5975);
and U7266 (N_7266,N_4683,N_4647);
nand U7267 (N_7267,N_4686,N_5522);
nor U7268 (N_7268,N_4820,N_5362);
or U7269 (N_7269,N_4776,N_5591);
nand U7270 (N_7270,N_5662,N_4585);
nand U7271 (N_7271,N_5921,N_4754);
nand U7272 (N_7272,N_5467,N_5046);
nand U7273 (N_7273,N_5568,N_5865);
nor U7274 (N_7274,N_5629,N_5270);
xnor U7275 (N_7275,N_5959,N_5141);
nor U7276 (N_7276,N_4696,N_4687);
nand U7277 (N_7277,N_5991,N_5355);
xor U7278 (N_7278,N_5064,N_5628);
xnor U7279 (N_7279,N_5329,N_4520);
nand U7280 (N_7280,N_5900,N_4677);
nor U7281 (N_7281,N_5205,N_5858);
or U7282 (N_7282,N_4738,N_4803);
or U7283 (N_7283,N_4607,N_5452);
and U7284 (N_7284,N_5993,N_5311);
nor U7285 (N_7285,N_4905,N_4642);
nand U7286 (N_7286,N_4918,N_5366);
xnor U7287 (N_7287,N_5321,N_5439);
nand U7288 (N_7288,N_4879,N_5311);
nand U7289 (N_7289,N_5601,N_5789);
nand U7290 (N_7290,N_4674,N_5543);
xnor U7291 (N_7291,N_4944,N_5648);
and U7292 (N_7292,N_5021,N_4655);
and U7293 (N_7293,N_5112,N_4756);
xnor U7294 (N_7294,N_5543,N_4673);
xor U7295 (N_7295,N_5702,N_5219);
xnor U7296 (N_7296,N_4768,N_5385);
nand U7297 (N_7297,N_4648,N_4502);
and U7298 (N_7298,N_5562,N_5121);
and U7299 (N_7299,N_5658,N_4888);
xnor U7300 (N_7300,N_4759,N_5240);
or U7301 (N_7301,N_5229,N_4651);
nand U7302 (N_7302,N_5896,N_4697);
xnor U7303 (N_7303,N_5330,N_5078);
or U7304 (N_7304,N_5593,N_5220);
nand U7305 (N_7305,N_5366,N_5740);
xor U7306 (N_7306,N_4789,N_5320);
xor U7307 (N_7307,N_5545,N_4664);
xor U7308 (N_7308,N_5909,N_5346);
and U7309 (N_7309,N_5975,N_5560);
nor U7310 (N_7310,N_5335,N_5840);
nand U7311 (N_7311,N_5265,N_4603);
or U7312 (N_7312,N_4547,N_5308);
and U7313 (N_7313,N_5960,N_4949);
and U7314 (N_7314,N_5790,N_5659);
and U7315 (N_7315,N_4999,N_4696);
nand U7316 (N_7316,N_5640,N_5317);
xor U7317 (N_7317,N_5054,N_5093);
and U7318 (N_7318,N_4701,N_5655);
nor U7319 (N_7319,N_4911,N_5302);
nor U7320 (N_7320,N_4677,N_4770);
nand U7321 (N_7321,N_4588,N_5044);
nor U7322 (N_7322,N_5659,N_5143);
and U7323 (N_7323,N_5329,N_4659);
xnor U7324 (N_7324,N_4851,N_5405);
xor U7325 (N_7325,N_5405,N_5233);
nand U7326 (N_7326,N_5026,N_4863);
xor U7327 (N_7327,N_4583,N_5372);
and U7328 (N_7328,N_4926,N_4945);
or U7329 (N_7329,N_4575,N_5549);
and U7330 (N_7330,N_5338,N_4503);
xor U7331 (N_7331,N_5574,N_4963);
and U7332 (N_7332,N_5725,N_4701);
or U7333 (N_7333,N_5714,N_5140);
nor U7334 (N_7334,N_4595,N_5644);
xor U7335 (N_7335,N_4515,N_5484);
or U7336 (N_7336,N_5295,N_5061);
or U7337 (N_7337,N_4759,N_5785);
nand U7338 (N_7338,N_5795,N_5715);
and U7339 (N_7339,N_5337,N_4630);
and U7340 (N_7340,N_4553,N_5073);
nor U7341 (N_7341,N_5720,N_5537);
nor U7342 (N_7342,N_5237,N_4976);
nor U7343 (N_7343,N_5857,N_5756);
nand U7344 (N_7344,N_4578,N_5768);
or U7345 (N_7345,N_5424,N_5687);
nand U7346 (N_7346,N_4818,N_5897);
and U7347 (N_7347,N_4689,N_5557);
xnor U7348 (N_7348,N_4511,N_4677);
or U7349 (N_7349,N_4518,N_5176);
or U7350 (N_7350,N_5537,N_4749);
and U7351 (N_7351,N_4585,N_5398);
xor U7352 (N_7352,N_5447,N_4845);
xnor U7353 (N_7353,N_4551,N_5951);
nor U7354 (N_7354,N_5023,N_4917);
and U7355 (N_7355,N_5103,N_4780);
nand U7356 (N_7356,N_5731,N_4569);
nor U7357 (N_7357,N_5525,N_5876);
nand U7358 (N_7358,N_5667,N_5530);
or U7359 (N_7359,N_5160,N_4634);
nor U7360 (N_7360,N_5410,N_5031);
xnor U7361 (N_7361,N_4513,N_4603);
xnor U7362 (N_7362,N_5504,N_5285);
nand U7363 (N_7363,N_4510,N_5862);
or U7364 (N_7364,N_5984,N_5606);
nand U7365 (N_7365,N_5351,N_5125);
nor U7366 (N_7366,N_4982,N_5313);
nor U7367 (N_7367,N_5053,N_5232);
or U7368 (N_7368,N_4608,N_5193);
nand U7369 (N_7369,N_5234,N_5505);
nor U7370 (N_7370,N_4903,N_5867);
or U7371 (N_7371,N_5014,N_5705);
nand U7372 (N_7372,N_4610,N_5568);
and U7373 (N_7373,N_4643,N_4746);
xnor U7374 (N_7374,N_4501,N_4666);
xor U7375 (N_7375,N_4933,N_4659);
and U7376 (N_7376,N_4952,N_5811);
nor U7377 (N_7377,N_4526,N_5024);
and U7378 (N_7378,N_5385,N_5927);
or U7379 (N_7379,N_5393,N_5056);
xor U7380 (N_7380,N_5962,N_4507);
or U7381 (N_7381,N_4613,N_4891);
xnor U7382 (N_7382,N_4876,N_4924);
xnor U7383 (N_7383,N_4727,N_4592);
and U7384 (N_7384,N_4659,N_4671);
or U7385 (N_7385,N_4897,N_5428);
nor U7386 (N_7386,N_5560,N_5860);
and U7387 (N_7387,N_5451,N_4593);
nor U7388 (N_7388,N_5519,N_5975);
and U7389 (N_7389,N_5342,N_5044);
xor U7390 (N_7390,N_5031,N_5866);
nand U7391 (N_7391,N_5217,N_4745);
or U7392 (N_7392,N_5698,N_5002);
or U7393 (N_7393,N_5284,N_5043);
nor U7394 (N_7394,N_5089,N_4822);
nand U7395 (N_7395,N_4552,N_4618);
or U7396 (N_7396,N_5123,N_5018);
nand U7397 (N_7397,N_5718,N_5659);
nor U7398 (N_7398,N_5054,N_5935);
nor U7399 (N_7399,N_4910,N_5769);
and U7400 (N_7400,N_5160,N_5485);
xor U7401 (N_7401,N_5413,N_5778);
xor U7402 (N_7402,N_4678,N_4658);
and U7403 (N_7403,N_5481,N_5546);
or U7404 (N_7404,N_5701,N_5927);
xor U7405 (N_7405,N_5706,N_5576);
xnor U7406 (N_7406,N_5930,N_5903);
or U7407 (N_7407,N_4769,N_5154);
or U7408 (N_7408,N_5412,N_5314);
and U7409 (N_7409,N_4660,N_5508);
nor U7410 (N_7410,N_4995,N_5845);
or U7411 (N_7411,N_5803,N_4564);
or U7412 (N_7412,N_5372,N_5212);
xnor U7413 (N_7413,N_4580,N_5445);
nor U7414 (N_7414,N_5563,N_4621);
and U7415 (N_7415,N_5213,N_5470);
nand U7416 (N_7416,N_5812,N_5092);
xnor U7417 (N_7417,N_4704,N_5772);
nor U7418 (N_7418,N_4574,N_5560);
nor U7419 (N_7419,N_4596,N_5471);
xnor U7420 (N_7420,N_4990,N_5032);
nor U7421 (N_7421,N_5701,N_5751);
nand U7422 (N_7422,N_5959,N_4746);
nand U7423 (N_7423,N_4961,N_5812);
nand U7424 (N_7424,N_5429,N_4661);
nor U7425 (N_7425,N_5022,N_4890);
xnor U7426 (N_7426,N_5217,N_5257);
xor U7427 (N_7427,N_5160,N_5578);
xor U7428 (N_7428,N_5133,N_5967);
xnor U7429 (N_7429,N_5227,N_5186);
nor U7430 (N_7430,N_5722,N_4914);
nand U7431 (N_7431,N_5300,N_5001);
nand U7432 (N_7432,N_5973,N_4775);
and U7433 (N_7433,N_4561,N_5478);
and U7434 (N_7434,N_4809,N_5050);
xor U7435 (N_7435,N_5133,N_4795);
and U7436 (N_7436,N_5864,N_4940);
nand U7437 (N_7437,N_5102,N_5196);
and U7438 (N_7438,N_4930,N_4853);
xnor U7439 (N_7439,N_5955,N_5319);
xor U7440 (N_7440,N_5014,N_5155);
xor U7441 (N_7441,N_4916,N_4703);
xnor U7442 (N_7442,N_5688,N_5649);
and U7443 (N_7443,N_4784,N_5852);
xnor U7444 (N_7444,N_4510,N_5326);
nand U7445 (N_7445,N_5014,N_5596);
and U7446 (N_7446,N_4964,N_5229);
nand U7447 (N_7447,N_4715,N_5971);
nand U7448 (N_7448,N_5277,N_4666);
nand U7449 (N_7449,N_4896,N_4954);
nor U7450 (N_7450,N_5729,N_5031);
xnor U7451 (N_7451,N_5415,N_4538);
xor U7452 (N_7452,N_4541,N_5056);
xor U7453 (N_7453,N_4533,N_4538);
xnor U7454 (N_7454,N_4651,N_5568);
or U7455 (N_7455,N_5794,N_4852);
and U7456 (N_7456,N_5370,N_5574);
xor U7457 (N_7457,N_4918,N_5754);
xor U7458 (N_7458,N_5712,N_4545);
xnor U7459 (N_7459,N_5208,N_5326);
nor U7460 (N_7460,N_4705,N_4505);
nor U7461 (N_7461,N_5295,N_5682);
and U7462 (N_7462,N_5800,N_4536);
nand U7463 (N_7463,N_5796,N_4843);
xor U7464 (N_7464,N_5706,N_4911);
nand U7465 (N_7465,N_5625,N_5627);
nor U7466 (N_7466,N_4946,N_4575);
or U7467 (N_7467,N_5729,N_5709);
and U7468 (N_7468,N_5987,N_4889);
and U7469 (N_7469,N_4552,N_4851);
or U7470 (N_7470,N_5529,N_5823);
xnor U7471 (N_7471,N_4968,N_4962);
and U7472 (N_7472,N_4983,N_5297);
xnor U7473 (N_7473,N_5750,N_5137);
and U7474 (N_7474,N_5848,N_5177);
and U7475 (N_7475,N_5839,N_4510);
or U7476 (N_7476,N_4576,N_4926);
xnor U7477 (N_7477,N_4776,N_5424);
nand U7478 (N_7478,N_5827,N_4763);
nand U7479 (N_7479,N_5596,N_5964);
or U7480 (N_7480,N_4760,N_5665);
or U7481 (N_7481,N_5753,N_5409);
and U7482 (N_7482,N_5201,N_5187);
and U7483 (N_7483,N_5307,N_5455);
or U7484 (N_7484,N_5755,N_5140);
xnor U7485 (N_7485,N_4743,N_4779);
and U7486 (N_7486,N_4855,N_4565);
xnor U7487 (N_7487,N_4898,N_5305);
nor U7488 (N_7488,N_5654,N_4537);
xnor U7489 (N_7489,N_4596,N_5291);
xor U7490 (N_7490,N_5002,N_4652);
nand U7491 (N_7491,N_5505,N_4766);
nand U7492 (N_7492,N_5137,N_5136);
and U7493 (N_7493,N_5497,N_5711);
and U7494 (N_7494,N_5504,N_4733);
and U7495 (N_7495,N_5342,N_5407);
nand U7496 (N_7496,N_5705,N_5101);
nor U7497 (N_7497,N_5299,N_5880);
or U7498 (N_7498,N_5300,N_4738);
xnor U7499 (N_7499,N_4795,N_5593);
xor U7500 (N_7500,N_7336,N_7217);
xor U7501 (N_7501,N_7433,N_6510);
or U7502 (N_7502,N_7112,N_6593);
xor U7503 (N_7503,N_6693,N_6490);
nand U7504 (N_7504,N_6332,N_6461);
and U7505 (N_7505,N_6955,N_7042);
and U7506 (N_7506,N_6360,N_6058);
xnor U7507 (N_7507,N_7454,N_6975);
xnor U7508 (N_7508,N_7090,N_6178);
or U7509 (N_7509,N_7301,N_7121);
xor U7510 (N_7510,N_6962,N_6493);
or U7511 (N_7511,N_7131,N_7388);
and U7512 (N_7512,N_6006,N_7200);
or U7513 (N_7513,N_6701,N_6543);
xor U7514 (N_7514,N_7476,N_6044);
and U7515 (N_7515,N_6748,N_6207);
or U7516 (N_7516,N_7171,N_6891);
or U7517 (N_7517,N_7108,N_6610);
nor U7518 (N_7518,N_7417,N_6934);
and U7519 (N_7519,N_6276,N_7403);
xor U7520 (N_7520,N_7367,N_7236);
nor U7521 (N_7521,N_6579,N_6434);
nand U7522 (N_7522,N_7369,N_6477);
xor U7523 (N_7523,N_7187,N_7292);
nand U7524 (N_7524,N_7496,N_6895);
xnor U7525 (N_7525,N_7157,N_6268);
xnor U7526 (N_7526,N_6395,N_7457);
nand U7527 (N_7527,N_7359,N_6738);
and U7528 (N_7528,N_7068,N_7310);
and U7529 (N_7529,N_7287,N_6181);
nor U7530 (N_7530,N_7041,N_6481);
nand U7531 (N_7531,N_6985,N_6994);
or U7532 (N_7532,N_7159,N_6845);
nand U7533 (N_7533,N_6781,N_7240);
nor U7534 (N_7534,N_6068,N_6015);
xor U7535 (N_7535,N_6079,N_6894);
and U7536 (N_7536,N_7396,N_7362);
nand U7537 (N_7537,N_7306,N_6864);
nand U7538 (N_7538,N_6464,N_6407);
nor U7539 (N_7539,N_6812,N_6870);
or U7540 (N_7540,N_6088,N_6148);
nand U7541 (N_7541,N_6502,N_6007);
nor U7542 (N_7542,N_6711,N_6762);
or U7543 (N_7543,N_6304,N_6730);
xor U7544 (N_7544,N_6650,N_7429);
xnor U7545 (N_7545,N_7133,N_6496);
nor U7546 (N_7546,N_6688,N_7030);
xor U7547 (N_7547,N_7009,N_6888);
xnor U7548 (N_7548,N_7286,N_7486);
or U7549 (N_7549,N_6430,N_6445);
nand U7550 (N_7550,N_7186,N_6678);
or U7551 (N_7551,N_6999,N_7373);
or U7552 (N_7552,N_6746,N_6056);
nand U7553 (N_7553,N_7463,N_6797);
and U7554 (N_7554,N_6644,N_7272);
xor U7555 (N_7555,N_7044,N_7389);
nor U7556 (N_7556,N_7479,N_6011);
xnor U7557 (N_7557,N_6474,N_7246);
nor U7558 (N_7558,N_6990,N_6214);
nand U7559 (N_7559,N_6336,N_6694);
xor U7560 (N_7560,N_6151,N_6583);
xnor U7561 (N_7561,N_6083,N_6270);
nand U7562 (N_7562,N_6731,N_6414);
xnor U7563 (N_7563,N_7071,N_6715);
and U7564 (N_7564,N_6780,N_7181);
nor U7565 (N_7565,N_7218,N_6288);
xor U7566 (N_7566,N_6317,N_6908);
or U7567 (N_7567,N_6102,N_6292);
nand U7568 (N_7568,N_6863,N_6790);
and U7569 (N_7569,N_7166,N_6334);
xor U7570 (N_7570,N_7151,N_6252);
nor U7571 (N_7571,N_6032,N_6147);
nor U7572 (N_7572,N_6002,N_6501);
and U7573 (N_7573,N_6622,N_6974);
and U7574 (N_7574,N_7224,N_7448);
xor U7575 (N_7575,N_7216,N_6358);
xor U7576 (N_7576,N_6145,N_6760);
xor U7577 (N_7577,N_7449,N_6967);
or U7578 (N_7578,N_6375,N_6896);
or U7579 (N_7579,N_7494,N_6699);
and U7580 (N_7580,N_7352,N_7118);
and U7581 (N_7581,N_6514,N_6843);
nand U7582 (N_7582,N_6728,N_6824);
or U7583 (N_7583,N_6233,N_7414);
or U7584 (N_7584,N_7179,N_6695);
nor U7585 (N_7585,N_6751,N_6783);
or U7586 (N_7586,N_7266,N_6259);
xnor U7587 (N_7587,N_6261,N_6476);
xor U7588 (N_7588,N_7168,N_6480);
nand U7589 (N_7589,N_6884,N_7124);
or U7590 (N_7590,N_7105,N_6067);
xor U7591 (N_7591,N_6373,N_7278);
nand U7592 (N_7592,N_7125,N_6383);
xnor U7593 (N_7593,N_6112,N_6979);
nor U7594 (N_7594,N_7464,N_7205);
or U7595 (N_7595,N_6499,N_7334);
nand U7596 (N_7596,N_7309,N_7196);
xor U7597 (N_7597,N_6813,N_6826);
nand U7598 (N_7598,N_6833,N_6902);
nand U7599 (N_7599,N_6568,N_6177);
nand U7600 (N_7600,N_6330,N_6584);
nand U7601 (N_7601,N_6471,N_7273);
and U7602 (N_7602,N_6662,N_6633);
nor U7603 (N_7603,N_7355,N_7184);
or U7604 (N_7604,N_7004,N_6462);
nand U7605 (N_7605,N_6498,N_7360);
xor U7606 (N_7606,N_6084,N_6885);
nor U7607 (N_7607,N_7234,N_6192);
nand U7608 (N_7608,N_6241,N_7130);
xnor U7609 (N_7609,N_6388,N_6577);
xor U7610 (N_7610,N_6237,N_6786);
and U7611 (N_7611,N_7317,N_6054);
nand U7612 (N_7612,N_6160,N_6025);
xor U7613 (N_7613,N_6131,N_7017);
or U7614 (N_7614,N_6681,N_6115);
nor U7615 (N_7615,N_6318,N_6630);
and U7616 (N_7616,N_6071,N_6931);
and U7617 (N_7617,N_6779,N_6647);
xnor U7618 (N_7618,N_6676,N_6114);
xnor U7619 (N_7619,N_6784,N_6046);
nand U7620 (N_7620,N_6950,N_6823);
nor U7621 (N_7621,N_7138,N_6907);
and U7622 (N_7622,N_7113,N_7320);
or U7623 (N_7623,N_6628,N_6980);
nor U7624 (N_7624,N_6665,N_7357);
or U7625 (N_7625,N_6544,N_7192);
nor U7626 (N_7626,N_6886,N_6713);
nor U7627 (N_7627,N_6216,N_6314);
xor U7628 (N_7628,N_6369,N_6286);
or U7629 (N_7629,N_6134,N_6101);
or U7630 (N_7630,N_6904,N_6599);
and U7631 (N_7631,N_7338,N_6653);
nor U7632 (N_7632,N_7328,N_6224);
nand U7633 (N_7633,N_6053,N_6277);
nor U7634 (N_7634,N_6322,N_6364);
and U7635 (N_7635,N_7458,N_6109);
and U7636 (N_7636,N_6850,N_6897);
or U7637 (N_7637,N_6768,N_6554);
and U7638 (N_7638,N_7390,N_6413);
xor U7639 (N_7639,N_7230,N_6637);
xnor U7640 (N_7640,N_6608,N_7145);
xnor U7641 (N_7641,N_6656,N_7208);
and U7642 (N_7642,N_6486,N_6909);
nand U7643 (N_7643,N_7488,N_7165);
and U7644 (N_7644,N_6242,N_7180);
and U7645 (N_7645,N_6700,N_6307);
nor U7646 (N_7646,N_6732,N_7487);
and U7647 (N_7647,N_7032,N_6840);
nand U7648 (N_7648,N_6774,N_6235);
or U7649 (N_7649,N_7249,N_6572);
and U7650 (N_7650,N_7239,N_7421);
nand U7651 (N_7651,N_6319,N_6411);
and U7652 (N_7652,N_6150,N_7087);
or U7653 (N_7653,N_7387,N_7086);
nor U7654 (N_7654,N_6977,N_7285);
nor U7655 (N_7655,N_6116,N_7128);
xnor U7656 (N_7656,N_7482,N_6403);
nor U7657 (N_7657,N_6100,N_6542);
and U7658 (N_7658,N_7252,N_6794);
xnor U7659 (N_7659,N_7470,N_6218);
xor U7660 (N_7660,N_7380,N_7141);
xor U7661 (N_7661,N_7412,N_6925);
and U7662 (N_7662,N_7258,N_6459);
or U7663 (N_7663,N_6141,N_7061);
nor U7664 (N_7664,N_6515,N_7024);
xor U7665 (N_7665,N_6368,N_6918);
nand U7666 (N_7666,N_7035,N_6377);
nand U7667 (N_7667,N_7423,N_7007);
nor U7668 (N_7668,N_7314,N_7099);
xnor U7669 (N_7669,N_6191,N_6533);
nand U7670 (N_7670,N_6356,N_6851);
or U7671 (N_7671,N_6454,N_6726);
and U7672 (N_7672,N_6537,N_6488);
xnor U7673 (N_7673,N_7049,N_6170);
and U7674 (N_7674,N_7177,N_6799);
and U7675 (N_7675,N_6272,N_6744);
nand U7676 (N_7676,N_6303,N_6697);
or U7677 (N_7677,N_7191,N_6816);
nor U7678 (N_7678,N_6031,N_6301);
nor U7679 (N_7679,N_6457,N_7075);
nor U7680 (N_7680,N_6226,N_7443);
nor U7681 (N_7681,N_7144,N_6956);
and U7682 (N_7682,N_6539,N_7394);
nor U7683 (N_7683,N_6070,N_6211);
and U7684 (N_7684,N_6952,N_6857);
xor U7685 (N_7685,N_7284,N_6519);
and U7686 (N_7686,N_7148,N_6418);
nor U7687 (N_7687,N_6405,N_6624);
nor U7688 (N_7688,N_6529,N_6924);
and U7689 (N_7689,N_6926,N_6353);
nand U7690 (N_7690,N_6775,N_7327);
nor U7691 (N_7691,N_6337,N_6815);
or U7692 (N_7692,N_6040,N_7424);
or U7693 (N_7693,N_6466,N_7103);
nor U7694 (N_7694,N_6335,N_7185);
and U7695 (N_7695,N_7139,N_6366);
nand U7696 (N_7696,N_6094,N_7193);
or U7697 (N_7697,N_6901,N_6659);
nor U7698 (N_7698,N_7023,N_7472);
nor U7699 (N_7699,N_6538,N_7100);
and U7700 (N_7700,N_6463,N_7440);
nand U7701 (N_7701,N_7221,N_6964);
nor U7702 (N_7702,N_7422,N_7435);
and U7703 (N_7703,N_6789,N_6119);
and U7704 (N_7704,N_6846,N_6961);
and U7705 (N_7705,N_6168,N_7307);
or U7706 (N_7706,N_7361,N_7462);
or U7707 (N_7707,N_6588,N_6839);
xor U7708 (N_7708,N_6201,N_7093);
nand U7709 (N_7709,N_7415,N_6323);
xnor U7710 (N_7710,N_6692,N_6600);
or U7711 (N_7711,N_7228,N_6995);
or U7712 (N_7712,N_6944,N_7325);
or U7713 (N_7713,N_6295,N_6485);
and U7714 (N_7714,N_7436,N_6844);
and U7715 (N_7715,N_6282,N_6887);
and U7716 (N_7716,N_7297,N_6427);
or U7717 (N_7717,N_6431,N_6449);
nor U7718 (N_7718,N_7289,N_7295);
xnor U7719 (N_7719,N_6299,N_7247);
nand U7720 (N_7720,N_6657,N_6777);
nor U7721 (N_7721,N_6540,N_7109);
or U7722 (N_7722,N_7120,N_6014);
nor U7723 (N_7723,N_7003,N_7382);
nor U7724 (N_7724,N_7135,N_6889);
xnor U7725 (N_7725,N_6171,N_6667);
xnor U7726 (N_7726,N_7060,N_6852);
nand U7727 (N_7727,N_6144,N_6039);
or U7728 (N_7728,N_6574,N_6422);
nor U7729 (N_7729,N_6140,N_6293);
nand U7730 (N_7730,N_6984,N_6387);
and U7731 (N_7731,N_6338,N_7465);
xor U7732 (N_7732,N_6219,N_6012);
nand U7733 (N_7733,N_6120,N_7152);
nor U7734 (N_7734,N_6047,N_6123);
nand U7735 (N_7735,N_6569,N_6442);
or U7736 (N_7736,N_6664,N_6257);
nand U7737 (N_7737,N_6029,N_7259);
nor U7738 (N_7738,N_7451,N_6167);
xor U7739 (N_7739,N_7401,N_6722);
xor U7740 (N_7740,N_7340,N_7447);
nor U7741 (N_7741,N_6500,N_6076);
or U7742 (N_7742,N_7210,N_6865);
and U7743 (N_7743,N_6346,N_6856);
nor U7744 (N_7744,N_7413,N_6055);
xor U7745 (N_7745,N_6398,N_6595);
nor U7746 (N_7746,N_6180,N_6787);
and U7747 (N_7747,N_6671,N_6443);
nand U7748 (N_7748,N_6832,N_6260);
nor U7749 (N_7749,N_7364,N_6796);
xor U7750 (N_7750,N_6525,N_6196);
nor U7751 (N_7751,N_6565,N_7257);
nand U7752 (N_7752,N_6792,N_6808);
nand U7753 (N_7753,N_6279,N_6429);
or U7754 (N_7754,N_6670,N_6757);
and U7755 (N_7755,N_7046,N_7083);
nor U7756 (N_7756,N_6194,N_7268);
nand U7757 (N_7757,N_6139,N_6996);
nand U7758 (N_7758,N_6673,N_7256);
or U7759 (N_7759,N_7303,N_6973);
nor U7760 (N_7760,N_7375,N_6831);
and U7761 (N_7761,N_6928,N_6878);
nor U7762 (N_7762,N_6234,N_7220);
xor U7763 (N_7763,N_6423,N_6987);
nand U7764 (N_7764,N_6549,N_6993);
or U7765 (N_7765,N_6080,N_6210);
or U7766 (N_7766,N_6215,N_6328);
xnor U7767 (N_7767,N_7232,N_6696);
or U7768 (N_7768,N_6448,N_7022);
and U7769 (N_7769,N_6426,N_7163);
nor U7770 (N_7770,N_6158,N_7214);
or U7771 (N_7771,N_7402,N_6698);
nand U7772 (N_7772,N_7053,N_6021);
nand U7773 (N_7773,N_6793,N_7491);
and U7774 (N_7774,N_6061,N_7263);
nor U7775 (N_7775,N_7203,N_6157);
nor U7776 (N_7776,N_7484,N_6484);
nor U7777 (N_7777,N_6626,N_7034);
or U7778 (N_7778,N_7377,N_6290);
nand U7779 (N_7779,N_6034,N_6174);
or U7780 (N_7780,N_6154,N_6737);
and U7781 (N_7781,N_6264,N_7197);
and U7782 (N_7782,N_6706,N_6853);
nand U7783 (N_7783,N_6024,N_6954);
and U7784 (N_7784,N_7194,N_6175);
nor U7785 (N_7785,N_7223,N_7097);
and U7786 (N_7786,N_6221,N_6617);
and U7787 (N_7787,N_6892,N_6655);
xor U7788 (N_7788,N_7119,N_7250);
or U7789 (N_7789,N_6509,N_6818);
or U7790 (N_7790,N_6893,N_6169);
nor U7791 (N_7791,N_7335,N_6858);
and U7792 (N_7792,N_7069,N_6129);
or U7793 (N_7793,N_6351,N_6385);
or U7794 (N_7794,N_7190,N_6077);
xnor U7795 (N_7795,N_6921,N_6208);
and U7796 (N_7796,N_6854,N_6912);
or U7797 (N_7797,N_7372,N_7043);
nand U7798 (N_7798,N_7226,N_6827);
or U7799 (N_7799,N_7419,N_7158);
xnor U7800 (N_7800,N_6776,N_7432);
nor U7801 (N_7801,N_6804,N_7005);
nand U7802 (N_7802,N_7073,N_7404);
nand U7803 (N_7803,N_7241,N_6478);
nand U7804 (N_7804,N_6597,N_7091);
xor U7805 (N_7805,N_6381,N_7170);
xnor U7806 (N_7806,N_7495,N_6450);
nand U7807 (N_7807,N_7400,N_6153);
nand U7808 (N_7808,N_7195,N_6313);
nand U7809 (N_7809,N_7027,N_6193);
nor U7810 (N_7810,N_6672,N_6527);
nand U7811 (N_7811,N_6524,N_7254);
nand U7812 (N_7812,N_6275,N_6458);
or U7813 (N_7813,N_6042,N_6045);
xor U7814 (N_7814,N_7173,N_7441);
nand U7815 (N_7815,N_6048,N_6842);
nor U7816 (N_7816,N_6410,N_6957);
xnor U7817 (N_7817,N_7153,N_7013);
nor U7818 (N_7818,N_6773,N_6531);
nor U7819 (N_7819,N_7425,N_6666);
nand U7820 (N_7820,N_6714,N_6370);
or U7821 (N_7821,N_6640,N_6755);
nor U7822 (N_7822,N_7288,N_6651);
and U7823 (N_7823,N_7174,N_6278);
nand U7824 (N_7824,N_7311,N_6986);
nor U7825 (N_7825,N_6258,N_6229);
nand U7826 (N_7826,N_7204,N_6942);
or U7827 (N_7827,N_6805,N_6801);
nand U7828 (N_7828,N_6915,N_6765);
or U7829 (N_7829,N_6689,N_6482);
or U7830 (N_7830,N_6828,N_6451);
nand U7831 (N_7831,N_6447,N_6406);
nor U7832 (N_7832,N_6562,N_7067);
nand U7833 (N_7833,N_6217,N_6709);
or U7834 (N_7834,N_6740,N_6619);
nand U7835 (N_7835,N_6236,N_7350);
nor U7836 (N_7836,N_6325,N_6872);
or U7837 (N_7837,N_7444,N_7383);
nand U7838 (N_7838,N_7167,N_7384);
xnor U7839 (N_7839,N_6036,N_6312);
nand U7840 (N_7840,N_6612,N_6057);
and U7841 (N_7841,N_7021,N_6273);
nor U7842 (N_7842,N_6587,N_6747);
or U7843 (N_7843,N_7363,N_6770);
nor U7844 (N_7844,N_6380,N_6598);
xor U7845 (N_7845,N_6038,N_7248);
xnor U7846 (N_7846,N_6248,N_7242);
nand U7847 (N_7847,N_6933,N_7480);
nand U7848 (N_7848,N_6750,N_7172);
nand U7849 (N_7849,N_6707,N_7074);
and U7850 (N_7850,N_6329,N_6274);
nand U7851 (N_7851,N_6350,N_7446);
xor U7852 (N_7852,N_6017,N_6625);
nand U7853 (N_7853,N_7341,N_7082);
and U7854 (N_7854,N_6511,N_6641);
nand U7855 (N_7855,N_6124,N_6195);
nand U7856 (N_7856,N_7331,N_6105);
xnor U7857 (N_7857,N_7420,N_7142);
or U7858 (N_7858,N_6530,N_6734);
nand U7859 (N_7859,N_6880,N_6165);
xnor U7860 (N_7860,N_7453,N_7057);
xnor U7861 (N_7861,N_6315,N_6310);
xor U7862 (N_7862,N_6004,N_6761);
nand U7863 (N_7863,N_7452,N_6735);
nor U7864 (N_7864,N_7198,N_6555);
and U7865 (N_7865,N_6382,N_6717);
and U7866 (N_7866,N_7321,N_6627);
or U7867 (N_7867,N_6016,N_6075);
xnor U7868 (N_7868,N_6010,N_6404);
and U7869 (N_7869,N_7215,N_7008);
and U7870 (N_7870,N_6691,N_7346);
xor U7871 (N_7871,N_6103,N_6108);
or U7872 (N_7872,N_7081,N_6809);
nor U7873 (N_7873,N_6877,N_6679);
nand U7874 (N_7874,N_6283,N_6631);
or U7875 (N_7875,N_7262,N_7026);
xor U7876 (N_7876,N_7048,N_6089);
xor U7877 (N_7877,N_7147,N_7156);
nor U7878 (N_7878,N_6415,N_6674);
or U7879 (N_7879,N_7342,N_6372);
xnor U7880 (N_7880,N_6397,N_7302);
and U7881 (N_7881,N_6172,N_6620);
nor U7882 (N_7882,N_6365,N_6795);
and U7883 (N_7883,N_6913,N_6914);
and U7884 (N_7884,N_6232,N_6348);
or U7885 (N_7885,N_6409,N_6118);
or U7886 (N_7886,N_6998,N_6836);
xnor U7887 (N_7887,N_6677,N_6206);
nor U7888 (N_7888,N_6309,N_7182);
or U7889 (N_7889,N_7326,N_6263);
nor U7890 (N_7890,N_6362,N_6199);
nand U7891 (N_7891,N_7466,N_7343);
nand U7892 (N_7892,N_6564,N_6374);
nand U7893 (N_7893,N_7291,N_6590);
xor U7894 (N_7894,N_6342,N_6817);
and U7895 (N_7895,N_6417,N_6663);
xor U7896 (N_7896,N_6632,N_7481);
and U7897 (N_7897,N_6528,N_6687);
xnor U7898 (N_7898,N_6135,N_6352);
nand U7899 (N_7899,N_6300,N_6585);
nand U7900 (N_7900,N_6030,N_6830);
xnor U7901 (N_7901,N_6764,N_7498);
xor U7902 (N_7902,N_6495,N_6615);
and U7903 (N_7903,N_6298,N_6550);
nand U7904 (N_7904,N_6333,N_6473);
xnor U7905 (N_7905,N_7054,N_6561);
nor U7906 (N_7906,N_7127,N_6008);
or U7907 (N_7907,N_6384,N_6560);
or U7908 (N_7908,N_7227,N_6269);
and U7909 (N_7909,N_6092,N_6861);
and U7910 (N_7910,N_6341,N_7146);
xor U7911 (N_7911,N_6517,N_7475);
nor U7912 (N_7912,N_7011,N_6161);
nor U7913 (N_7913,N_7033,N_6183);
nor U7914 (N_7914,N_7202,N_7237);
nor U7915 (N_7915,N_7366,N_7304);
and U7916 (N_7916,N_6113,N_6376);
or U7917 (N_7917,N_6802,N_6062);
nand U7918 (N_7918,N_7040,N_6197);
and U7919 (N_7919,N_7442,N_6825);
xnor U7920 (N_7920,N_6978,N_6073);
nand U7921 (N_7921,N_7395,N_7489);
and U7922 (N_7922,N_6654,N_7025);
and U7923 (N_7923,N_6200,N_6354);
nor U7924 (N_7924,N_7418,N_6204);
nand U7925 (N_7925,N_7055,N_6306);
nor U7926 (N_7926,N_7374,N_6874);
or U7927 (N_7927,N_7000,N_6690);
and U7928 (N_7928,N_6188,N_6899);
and U7929 (N_7929,N_6660,N_7492);
and U7930 (N_7930,N_6771,N_7010);
and U7931 (N_7931,N_7238,N_7376);
xor U7932 (N_7932,N_6271,N_6629);
and U7933 (N_7933,N_6037,N_7316);
or U7934 (N_7934,N_7102,N_7207);
nand U7935 (N_7935,N_7323,N_7381);
nor U7936 (N_7936,N_6041,N_6882);
and U7937 (N_7937,N_6091,N_7426);
xnor U7938 (N_7938,N_7260,N_6769);
or U7939 (N_7939,N_7299,N_6189);
and U7940 (N_7940,N_7150,N_6126);
nor U7941 (N_7941,N_6834,N_6652);
and U7942 (N_7942,N_6661,N_6308);
and U7943 (N_7943,N_6685,N_6910);
or U7944 (N_7944,N_6623,N_6548);
and U7945 (N_7945,N_6604,N_6951);
nand U7946 (N_7946,N_6251,N_6492);
or U7947 (N_7947,N_7267,N_6876);
nor U7948 (N_7948,N_6541,N_6439);
or U7949 (N_7949,N_6117,N_7308);
or U7950 (N_7950,N_6649,N_7070);
nor U7951 (N_7951,N_6327,N_6645);
and U7952 (N_7952,N_6149,N_6922);
and U7953 (N_7953,N_7365,N_7134);
nor U7954 (N_7954,N_6324,N_7019);
and U7955 (N_7955,N_7149,N_6020);
and U7956 (N_7956,N_7438,N_6110);
nand U7957 (N_7957,N_7430,N_6552);
xor U7958 (N_7958,N_6121,N_7276);
or U7959 (N_7959,N_6494,N_7499);
nand U7960 (N_7960,N_6820,N_7235);
and U7961 (N_7961,N_7371,N_6708);
and U7962 (N_7962,N_7461,N_6349);
nor U7963 (N_7963,N_6347,N_6256);
nand U7964 (N_7964,N_7175,N_6621);
nand U7965 (N_7965,N_6396,N_6096);
or U7966 (N_7966,N_7368,N_6111);
or U7967 (N_7967,N_7012,N_7379);
or U7968 (N_7968,N_7445,N_7183);
nand U7969 (N_7969,N_6069,N_6758);
xor U7970 (N_7970,N_7076,N_6142);
and U7971 (N_7971,N_6386,N_6001);
or U7972 (N_7972,N_7264,N_6586);
and U7973 (N_7973,N_6847,N_6465);
xnor U7974 (N_7974,N_6606,N_7161);
xor U7975 (N_7975,N_6719,N_7279);
nand U7976 (N_7976,N_7271,N_7261);
or U7977 (N_7977,N_6163,N_6436);
or U7978 (N_7978,N_7098,N_6971);
and U7979 (N_7979,N_7493,N_6785);
or U7980 (N_7980,N_6320,N_6821);
xnor U7981 (N_7981,N_7409,N_6782);
and U7982 (N_7982,N_6575,N_7092);
and U7983 (N_7983,N_6835,N_7162);
or U7984 (N_7984,N_7459,N_6592);
or U7985 (N_7985,N_6855,N_6359);
and U7986 (N_7986,N_6456,N_6203);
nand U7987 (N_7987,N_6723,N_6455);
xnor U7988 (N_7988,N_6052,N_6222);
and U7989 (N_7989,N_6085,N_7085);
or U7990 (N_7990,N_6166,N_6159);
nand U7991 (N_7991,N_6508,N_6246);
or U7992 (N_7992,N_6727,N_6223);
xor U7993 (N_7993,N_6532,N_6937);
or U7994 (N_7994,N_7225,N_6280);
and U7995 (N_7995,N_7282,N_6098);
and U7996 (N_7996,N_6402,N_6064);
xnor U7997 (N_7997,N_7002,N_7468);
xor U7998 (N_7998,N_6883,N_6146);
nand U7999 (N_7999,N_7045,N_6960);
or U8000 (N_8000,N_6939,N_6090);
nor U8001 (N_8001,N_6250,N_6611);
or U8002 (N_8002,N_7330,N_7416);
and U8003 (N_8003,N_6534,N_6739);
nor U8004 (N_8004,N_6551,N_6989);
or U8005 (N_8005,N_6302,N_6868);
or U8006 (N_8006,N_6616,N_6243);
nor U8007 (N_8007,N_6097,N_6582);
nor U8008 (N_8008,N_6022,N_7251);
or U8009 (N_8009,N_6803,N_6253);
and U8010 (N_8010,N_6202,N_7222);
nand U8011 (N_8011,N_7104,N_6906);
nand U8012 (N_8012,N_6609,N_7107);
nand U8013 (N_8013,N_7111,N_6390);
nor U8014 (N_8014,N_6106,N_6389);
and U8015 (N_8015,N_6571,N_6866);
nand U8016 (N_8016,N_7080,N_6841);
or U8017 (N_8017,N_6753,N_6547);
or U8018 (N_8018,N_6618,N_6573);
or U8019 (N_8019,N_7332,N_6355);
nor U8020 (N_8020,N_7243,N_6441);
xnor U8021 (N_8021,N_6213,N_6911);
or U8022 (N_8022,N_6743,N_7305);
or U8023 (N_8023,N_6953,N_7140);
nand U8024 (N_8024,N_6505,N_7293);
or U8025 (N_8025,N_7066,N_7231);
nand U8026 (N_8026,N_6176,N_7037);
and U8027 (N_8027,N_6535,N_6479);
and U8028 (N_8028,N_6972,N_6557);
or U8029 (N_8029,N_6668,N_7122);
nor U8030 (N_8030,N_7201,N_6491);
nor U8031 (N_8031,N_6287,N_7137);
xor U8032 (N_8032,N_6043,N_7116);
nor U8033 (N_8033,N_6078,N_7385);
or U8034 (N_8034,N_7213,N_7407);
xor U8035 (N_8035,N_6965,N_6507);
nand U8036 (N_8036,N_7001,N_7020);
and U8037 (N_8037,N_6187,N_6143);
and U8038 (N_8038,N_6412,N_6000);
or U8039 (N_8039,N_6297,N_7391);
xor U8040 (N_8040,N_6703,N_7312);
nor U8041 (N_8041,N_6523,N_6220);
nor U8042 (N_8042,N_6992,N_7349);
and U8043 (N_8043,N_7039,N_6066);
nor U8044 (N_8044,N_7006,N_6742);
nor U8045 (N_8045,N_7255,N_7209);
xor U8046 (N_8046,N_6982,N_7199);
nor U8047 (N_8047,N_6898,N_7126);
nor U8048 (N_8048,N_6033,N_6005);
nand U8049 (N_8049,N_6281,N_7245);
xnor U8050 (N_8050,N_6567,N_6578);
or U8051 (N_8051,N_6838,N_6050);
xnor U8052 (N_8052,N_6262,N_7353);
and U8053 (N_8053,N_6859,N_7450);
xor U8054 (N_8054,N_6756,N_7176);
or U8055 (N_8055,N_6553,N_6453);
nor U8056 (N_8056,N_7094,N_6772);
xnor U8057 (N_8057,N_6945,N_7160);
or U8058 (N_8058,N_7397,N_6682);
xor U8059 (N_8059,N_6049,N_7280);
nand U8060 (N_8060,N_6475,N_6563);
or U8061 (N_8061,N_6483,N_6470);
nand U8062 (N_8062,N_7129,N_7283);
or U8063 (N_8063,N_7253,N_6026);
nand U8064 (N_8064,N_6968,N_6745);
nor U8065 (N_8065,N_7078,N_6357);
or U8066 (N_8066,N_7333,N_6254);
xnor U8067 (N_8067,N_6059,N_6240);
nor U8068 (N_8068,N_6581,N_6638);
xnor U8069 (N_8069,N_6721,N_6467);
xor U8070 (N_8070,N_7485,N_7322);
and U8071 (N_8071,N_6741,N_6340);
nand U8072 (N_8072,N_6130,N_7274);
nand U8073 (N_8073,N_6936,N_6291);
nor U8074 (N_8074,N_7298,N_6512);
or U8075 (N_8075,N_6035,N_6074);
and U8076 (N_8076,N_7339,N_6930);
nand U8077 (N_8077,N_6634,N_6546);
nor U8078 (N_8078,N_7212,N_6605);
and U8079 (N_8079,N_7018,N_6704);
and U8080 (N_8080,N_7398,N_6122);
xor U8081 (N_8081,N_6943,N_6027);
nand U8082 (N_8082,N_7188,N_6733);
or U8083 (N_8083,N_6503,N_6518);
nand U8084 (N_8084,N_6736,N_6400);
nor U8085 (N_8085,N_6917,N_6446);
and U8086 (N_8086,N_6244,N_6255);
or U8087 (N_8087,N_6513,N_7490);
or U8088 (N_8088,N_7428,N_7028);
or U8089 (N_8089,N_6752,N_6227);
nand U8090 (N_8090,N_7483,N_7132);
or U8091 (N_8091,N_6890,N_7431);
and U8092 (N_8092,N_6594,N_7467);
xnor U8093 (N_8093,N_6522,N_7056);
nor U8094 (N_8094,N_7393,N_6879);
nor U8095 (N_8095,N_6468,N_6249);
nand U8096 (N_8096,N_6104,N_6545);
nand U8097 (N_8097,N_6162,N_7300);
nand U8098 (N_8098,N_6469,N_6435);
or U8099 (N_8099,N_6558,N_6576);
xor U8100 (N_8100,N_7277,N_6391);
or U8101 (N_8101,N_6935,N_7324);
xnor U8102 (N_8102,N_7088,N_7106);
nand U8103 (N_8103,N_6099,N_6788);
or U8104 (N_8104,N_6186,N_7456);
and U8105 (N_8105,N_7029,N_6156);
or U8106 (N_8106,N_6959,N_6399);
nor U8107 (N_8107,N_6339,N_6862);
xnor U8108 (N_8108,N_7244,N_6829);
nor U8109 (N_8109,N_6095,N_6003);
nand U8110 (N_8110,N_6729,N_6013);
nor U8111 (N_8111,N_7290,N_6343);
nand U8112 (N_8112,N_7358,N_6873);
nand U8113 (N_8113,N_6127,N_6401);
nor U8114 (N_8114,N_6392,N_6432);
and U8115 (N_8115,N_6536,N_6822);
and U8116 (N_8116,N_6311,N_7015);
and U8117 (N_8117,N_6023,N_6230);
or U8118 (N_8118,N_6393,N_6602);
nand U8119 (N_8119,N_7123,N_6763);
and U8120 (N_8120,N_7281,N_6559);
or U8121 (N_8121,N_6132,N_6966);
nor U8122 (N_8122,N_7370,N_7047);
nand U8123 (N_8123,N_7406,N_6869);
nor U8124 (N_8124,N_7233,N_7319);
or U8125 (N_8125,N_6881,N_7354);
xnor U8126 (N_8126,N_6452,N_6718);
xor U8127 (N_8127,N_7497,N_6648);
xor U8128 (N_8128,N_7434,N_7471);
nor U8129 (N_8129,N_7294,N_7265);
nor U8130 (N_8130,N_6806,N_6981);
nand U8131 (N_8131,N_6239,N_6988);
nor U8132 (N_8132,N_6344,N_6556);
and U8133 (N_8133,N_7439,N_6316);
xor U8134 (N_8134,N_7206,N_7399);
or U8135 (N_8135,N_6296,N_6636);
nand U8136 (N_8136,N_6428,N_6072);
xnor U8137 (N_8137,N_6419,N_7392);
or U8138 (N_8138,N_6504,N_6521);
and U8139 (N_8139,N_7058,N_6173);
or U8140 (N_8140,N_6983,N_6009);
nand U8141 (N_8141,N_6716,N_6408);
or U8142 (N_8142,N_7050,N_6378);
xor U8143 (N_8143,N_6367,N_7345);
xor U8144 (N_8144,N_7211,N_6416);
nand U8145 (N_8145,N_6238,N_6970);
xnor U8146 (N_8146,N_6028,N_6289);
nand U8147 (N_8147,N_6603,N_6155);
xor U8148 (N_8148,N_7115,N_6916);
or U8149 (N_8149,N_6639,N_6093);
nor U8150 (N_8150,N_7064,N_7169);
nand U8151 (N_8151,N_7337,N_6754);
nor U8152 (N_8152,N_7178,N_7079);
nand U8153 (N_8153,N_6019,N_7089);
and U8154 (N_8154,N_6848,N_6596);
or U8155 (N_8155,N_6345,N_7410);
or U8156 (N_8156,N_7052,N_7062);
or U8157 (N_8157,N_6190,N_6712);
xor U8158 (N_8158,N_6958,N_6497);
nand U8159 (N_8159,N_7117,N_7408);
and U8160 (N_8160,N_6580,N_6976);
and U8161 (N_8161,N_7348,N_6489);
nand U8162 (N_8162,N_6438,N_6212);
and U8163 (N_8163,N_7427,N_7275);
or U8164 (N_8164,N_6063,N_7315);
nand U8165 (N_8165,N_7269,N_6819);
or U8166 (N_8166,N_6963,N_6705);
or U8167 (N_8167,N_7110,N_7155);
nor U8168 (N_8168,N_6138,N_6516);
xor U8169 (N_8169,N_6520,N_6205);
nand U8170 (N_8170,N_7143,N_7478);
nor U8171 (N_8171,N_6228,N_6394);
xor U8172 (N_8172,N_6683,N_6710);
and U8173 (N_8173,N_7136,N_6903);
nand U8174 (N_8174,N_6997,N_6371);
xnor U8175 (N_8175,N_7329,N_7437);
nor U8176 (N_8176,N_6940,N_7016);
and U8177 (N_8177,N_7077,N_6460);
nand U8178 (N_8178,N_6184,N_6472);
and U8179 (N_8179,N_6720,N_7229);
nor U8180 (N_8180,N_6128,N_6927);
or U8181 (N_8181,N_6231,N_6946);
and U8182 (N_8182,N_6433,N_6294);
nand U8183 (N_8183,N_6152,N_6607);
nor U8184 (N_8184,N_6321,N_7405);
nand U8185 (N_8185,N_7101,N_6900);
xnor U8186 (N_8186,N_6949,N_7460);
nor U8187 (N_8187,N_6642,N_6810);
nand U8188 (N_8188,N_7296,N_6800);
nor U8189 (N_8189,N_6591,N_7344);
nor U8190 (N_8190,N_6182,N_7065);
or U8191 (N_8191,N_6440,N_6749);
or U8192 (N_8192,N_6421,N_6929);
xnor U8193 (N_8193,N_6566,N_6209);
nand U8194 (N_8194,N_6991,N_6526);
xnor U8195 (N_8195,N_7114,N_6225);
and U8196 (N_8196,N_7063,N_6245);
and U8197 (N_8197,N_6807,N_7378);
xnor U8198 (N_8198,N_6305,N_6860);
xnor U8199 (N_8199,N_6051,N_6082);
and U8200 (N_8200,N_7059,N_6871);
and U8201 (N_8201,N_6185,N_7219);
and U8202 (N_8202,N_7038,N_6635);
or U8203 (N_8203,N_6589,N_6923);
and U8204 (N_8204,N_6136,N_6646);
or U8205 (N_8205,N_7154,N_6198);
xor U8206 (N_8206,N_7051,N_6613);
and U8207 (N_8207,N_6331,N_6849);
nand U8208 (N_8208,N_6948,N_7014);
xor U8209 (N_8209,N_6614,N_6658);
or U8210 (N_8210,N_6060,N_6107);
or U8211 (N_8211,N_6675,N_6164);
or U8212 (N_8212,N_7270,N_7072);
nand U8213 (N_8213,N_7411,N_6506);
xnor U8214 (N_8214,N_7473,N_7386);
or U8215 (N_8215,N_6444,N_6125);
nor U8216 (N_8216,N_7031,N_6766);
or U8217 (N_8217,N_6437,N_6379);
and U8218 (N_8218,N_6087,N_6081);
or U8219 (N_8219,N_6798,N_7164);
xor U8220 (N_8220,N_6363,N_6947);
nor U8221 (N_8221,N_6684,N_7351);
or U8222 (N_8222,N_7313,N_6247);
xor U8223 (N_8223,N_6875,N_6767);
and U8224 (N_8224,N_6267,N_7096);
nand U8225 (N_8225,N_6814,N_6086);
or U8226 (N_8226,N_6487,N_6137);
and U8227 (N_8227,N_7036,N_6420);
xnor U8228 (N_8228,N_6778,N_6265);
or U8229 (N_8229,N_6702,N_6759);
nand U8230 (N_8230,N_7084,N_6643);
and U8231 (N_8231,N_6425,N_6920);
and U8232 (N_8232,N_7474,N_6941);
and U8233 (N_8233,N_7477,N_6867);
nor U8234 (N_8234,N_6724,N_6285);
nand U8235 (N_8235,N_7189,N_7347);
and U8236 (N_8236,N_6179,N_6284);
nor U8237 (N_8237,N_7469,N_6680);
xor U8238 (N_8238,N_6969,N_6791);
or U8239 (N_8239,N_7356,N_6601);
or U8240 (N_8240,N_6919,N_6570);
nand U8241 (N_8241,N_6938,N_7095);
nor U8242 (N_8242,N_7318,N_6905);
or U8243 (N_8243,N_6686,N_6932);
and U8244 (N_8244,N_6811,N_6326);
nand U8245 (N_8245,N_6133,N_6065);
nand U8246 (N_8246,N_6837,N_6669);
or U8247 (N_8247,N_7455,N_6361);
nand U8248 (N_8248,N_6266,N_6725);
and U8249 (N_8249,N_6018,N_6424);
or U8250 (N_8250,N_6420,N_7476);
nor U8251 (N_8251,N_6281,N_7329);
or U8252 (N_8252,N_7022,N_6330);
and U8253 (N_8253,N_6503,N_7075);
xnor U8254 (N_8254,N_7121,N_6345);
xor U8255 (N_8255,N_6824,N_6251);
xor U8256 (N_8256,N_6520,N_7299);
nor U8257 (N_8257,N_6914,N_7189);
and U8258 (N_8258,N_6699,N_7490);
nand U8259 (N_8259,N_7369,N_7404);
and U8260 (N_8260,N_6708,N_7065);
and U8261 (N_8261,N_6482,N_6425);
nor U8262 (N_8262,N_6457,N_6962);
nor U8263 (N_8263,N_7084,N_6019);
xnor U8264 (N_8264,N_6329,N_6999);
or U8265 (N_8265,N_6959,N_6765);
or U8266 (N_8266,N_6960,N_6752);
and U8267 (N_8267,N_6278,N_6369);
nor U8268 (N_8268,N_7391,N_6425);
or U8269 (N_8269,N_7199,N_6294);
or U8270 (N_8270,N_7029,N_6590);
nand U8271 (N_8271,N_6577,N_7132);
xor U8272 (N_8272,N_7493,N_7348);
nand U8273 (N_8273,N_6952,N_7083);
and U8274 (N_8274,N_6409,N_6368);
nand U8275 (N_8275,N_6208,N_6828);
xnor U8276 (N_8276,N_6214,N_6032);
or U8277 (N_8277,N_6835,N_6203);
nand U8278 (N_8278,N_7429,N_6876);
or U8279 (N_8279,N_7482,N_6373);
or U8280 (N_8280,N_6670,N_7400);
or U8281 (N_8281,N_6091,N_7333);
and U8282 (N_8282,N_7263,N_6845);
nor U8283 (N_8283,N_7075,N_6851);
and U8284 (N_8284,N_6248,N_6630);
nor U8285 (N_8285,N_6516,N_7421);
nor U8286 (N_8286,N_6538,N_6361);
or U8287 (N_8287,N_6848,N_7196);
nand U8288 (N_8288,N_6261,N_6055);
nand U8289 (N_8289,N_6262,N_7273);
xor U8290 (N_8290,N_6661,N_6361);
nor U8291 (N_8291,N_7492,N_7178);
and U8292 (N_8292,N_6276,N_7489);
xnor U8293 (N_8293,N_7082,N_7171);
nand U8294 (N_8294,N_6928,N_7324);
and U8295 (N_8295,N_7458,N_6660);
nand U8296 (N_8296,N_7283,N_6846);
nand U8297 (N_8297,N_6883,N_6362);
xor U8298 (N_8298,N_6017,N_7365);
nor U8299 (N_8299,N_7356,N_7328);
xnor U8300 (N_8300,N_6736,N_7304);
or U8301 (N_8301,N_7362,N_7275);
xnor U8302 (N_8302,N_6636,N_6087);
or U8303 (N_8303,N_6002,N_6140);
or U8304 (N_8304,N_6995,N_7044);
nor U8305 (N_8305,N_6176,N_6375);
xnor U8306 (N_8306,N_7347,N_6520);
or U8307 (N_8307,N_6513,N_6967);
or U8308 (N_8308,N_6556,N_6248);
nor U8309 (N_8309,N_6751,N_6403);
xnor U8310 (N_8310,N_7082,N_6608);
and U8311 (N_8311,N_6304,N_6334);
nor U8312 (N_8312,N_7041,N_7168);
nand U8313 (N_8313,N_6610,N_6669);
or U8314 (N_8314,N_6408,N_6660);
nor U8315 (N_8315,N_6939,N_6608);
nand U8316 (N_8316,N_6852,N_7036);
nor U8317 (N_8317,N_6290,N_6162);
nor U8318 (N_8318,N_7295,N_7414);
nor U8319 (N_8319,N_7028,N_6046);
nor U8320 (N_8320,N_6183,N_7207);
or U8321 (N_8321,N_6228,N_6882);
and U8322 (N_8322,N_6025,N_7158);
nor U8323 (N_8323,N_6333,N_7399);
and U8324 (N_8324,N_6651,N_6735);
and U8325 (N_8325,N_7485,N_6706);
xnor U8326 (N_8326,N_6500,N_7495);
and U8327 (N_8327,N_6478,N_7182);
nor U8328 (N_8328,N_6314,N_7351);
and U8329 (N_8329,N_6370,N_7181);
or U8330 (N_8330,N_7138,N_7373);
and U8331 (N_8331,N_6604,N_7297);
xnor U8332 (N_8332,N_7108,N_6993);
or U8333 (N_8333,N_6442,N_7467);
and U8334 (N_8334,N_6572,N_6303);
xnor U8335 (N_8335,N_6022,N_7263);
nand U8336 (N_8336,N_7464,N_6825);
nand U8337 (N_8337,N_6929,N_6681);
xor U8338 (N_8338,N_7166,N_6199);
xor U8339 (N_8339,N_6613,N_6386);
nand U8340 (N_8340,N_7495,N_6103);
nand U8341 (N_8341,N_7369,N_7175);
nor U8342 (N_8342,N_6179,N_6938);
nor U8343 (N_8343,N_6250,N_6538);
nor U8344 (N_8344,N_6101,N_6179);
xnor U8345 (N_8345,N_7031,N_6719);
xor U8346 (N_8346,N_7181,N_6169);
nand U8347 (N_8347,N_6913,N_6864);
and U8348 (N_8348,N_6468,N_6832);
and U8349 (N_8349,N_6594,N_6211);
nor U8350 (N_8350,N_6892,N_6869);
and U8351 (N_8351,N_6988,N_6386);
or U8352 (N_8352,N_6675,N_6021);
or U8353 (N_8353,N_6779,N_6743);
or U8354 (N_8354,N_6296,N_7116);
xnor U8355 (N_8355,N_7185,N_6092);
nor U8356 (N_8356,N_6402,N_7409);
or U8357 (N_8357,N_6398,N_6153);
and U8358 (N_8358,N_7073,N_6236);
and U8359 (N_8359,N_7120,N_7306);
or U8360 (N_8360,N_6396,N_6139);
and U8361 (N_8361,N_6507,N_6559);
and U8362 (N_8362,N_6427,N_7229);
and U8363 (N_8363,N_6765,N_6106);
or U8364 (N_8364,N_6933,N_6381);
xor U8365 (N_8365,N_6397,N_6665);
xnor U8366 (N_8366,N_6201,N_6430);
nor U8367 (N_8367,N_7076,N_6249);
nor U8368 (N_8368,N_6661,N_6070);
nor U8369 (N_8369,N_7066,N_7222);
or U8370 (N_8370,N_7261,N_7375);
nor U8371 (N_8371,N_6245,N_7019);
nor U8372 (N_8372,N_6417,N_7153);
and U8373 (N_8373,N_7128,N_6722);
nor U8374 (N_8374,N_6664,N_6893);
xnor U8375 (N_8375,N_7457,N_6443);
xor U8376 (N_8376,N_6716,N_6131);
nor U8377 (N_8377,N_6799,N_6228);
nand U8378 (N_8378,N_7407,N_7421);
and U8379 (N_8379,N_6115,N_7143);
or U8380 (N_8380,N_7003,N_6525);
xor U8381 (N_8381,N_6943,N_6192);
or U8382 (N_8382,N_7372,N_7397);
xor U8383 (N_8383,N_6708,N_7376);
nand U8384 (N_8384,N_6140,N_6690);
xnor U8385 (N_8385,N_6673,N_6687);
nand U8386 (N_8386,N_7042,N_6485);
or U8387 (N_8387,N_6843,N_6715);
or U8388 (N_8388,N_6903,N_6010);
or U8389 (N_8389,N_6841,N_6247);
nand U8390 (N_8390,N_6262,N_7274);
nand U8391 (N_8391,N_6776,N_7205);
nor U8392 (N_8392,N_6274,N_7105);
nor U8393 (N_8393,N_7149,N_6071);
nor U8394 (N_8394,N_7444,N_6788);
nor U8395 (N_8395,N_7251,N_6926);
or U8396 (N_8396,N_7364,N_6268);
or U8397 (N_8397,N_7255,N_6312);
and U8398 (N_8398,N_7429,N_6448);
nor U8399 (N_8399,N_6477,N_6729);
or U8400 (N_8400,N_6789,N_6892);
or U8401 (N_8401,N_6420,N_6381);
xor U8402 (N_8402,N_6479,N_6492);
nor U8403 (N_8403,N_6573,N_7253);
or U8404 (N_8404,N_6177,N_6283);
nand U8405 (N_8405,N_6477,N_6961);
nor U8406 (N_8406,N_6153,N_6298);
xor U8407 (N_8407,N_7193,N_6275);
nor U8408 (N_8408,N_6274,N_6575);
or U8409 (N_8409,N_6662,N_7101);
or U8410 (N_8410,N_6093,N_6999);
xor U8411 (N_8411,N_6114,N_7069);
and U8412 (N_8412,N_7299,N_7051);
and U8413 (N_8413,N_6563,N_7311);
or U8414 (N_8414,N_7324,N_6965);
nor U8415 (N_8415,N_7074,N_6116);
or U8416 (N_8416,N_6294,N_6953);
nand U8417 (N_8417,N_6597,N_7375);
and U8418 (N_8418,N_6579,N_6609);
nor U8419 (N_8419,N_6719,N_6604);
and U8420 (N_8420,N_6834,N_7125);
or U8421 (N_8421,N_6028,N_7304);
or U8422 (N_8422,N_6860,N_7129);
nand U8423 (N_8423,N_6728,N_6156);
nor U8424 (N_8424,N_6504,N_6758);
nand U8425 (N_8425,N_6451,N_7193);
nor U8426 (N_8426,N_6631,N_6491);
xor U8427 (N_8427,N_6988,N_6161);
nor U8428 (N_8428,N_6103,N_7377);
nor U8429 (N_8429,N_6430,N_6252);
and U8430 (N_8430,N_7131,N_6191);
or U8431 (N_8431,N_7317,N_7023);
and U8432 (N_8432,N_7015,N_7303);
xor U8433 (N_8433,N_7033,N_7054);
nand U8434 (N_8434,N_7099,N_6635);
nand U8435 (N_8435,N_7143,N_6439);
nand U8436 (N_8436,N_7175,N_6761);
xor U8437 (N_8437,N_6517,N_6616);
nor U8438 (N_8438,N_6733,N_6244);
or U8439 (N_8439,N_6207,N_6795);
nand U8440 (N_8440,N_6669,N_7378);
xnor U8441 (N_8441,N_7077,N_6227);
or U8442 (N_8442,N_6829,N_6712);
or U8443 (N_8443,N_6989,N_6143);
and U8444 (N_8444,N_6173,N_6667);
nand U8445 (N_8445,N_6365,N_7076);
nor U8446 (N_8446,N_6515,N_6611);
xor U8447 (N_8447,N_7470,N_6415);
nand U8448 (N_8448,N_6902,N_6512);
and U8449 (N_8449,N_6091,N_6994);
nand U8450 (N_8450,N_6772,N_6003);
or U8451 (N_8451,N_6651,N_7474);
or U8452 (N_8452,N_7434,N_7061);
and U8453 (N_8453,N_6533,N_7337);
or U8454 (N_8454,N_6799,N_6931);
nand U8455 (N_8455,N_6619,N_6959);
and U8456 (N_8456,N_7158,N_6591);
nand U8457 (N_8457,N_6062,N_6597);
nand U8458 (N_8458,N_6908,N_6247);
or U8459 (N_8459,N_7220,N_6661);
or U8460 (N_8460,N_6106,N_7062);
xnor U8461 (N_8461,N_7270,N_6776);
xor U8462 (N_8462,N_6789,N_7157);
nand U8463 (N_8463,N_7047,N_7452);
nor U8464 (N_8464,N_6601,N_7227);
and U8465 (N_8465,N_7021,N_7396);
or U8466 (N_8466,N_6148,N_7394);
nor U8467 (N_8467,N_6143,N_6319);
and U8468 (N_8468,N_6695,N_6048);
and U8469 (N_8469,N_6511,N_6000);
xnor U8470 (N_8470,N_6880,N_7225);
and U8471 (N_8471,N_7416,N_6788);
or U8472 (N_8472,N_7203,N_6530);
nand U8473 (N_8473,N_6113,N_7215);
and U8474 (N_8474,N_6094,N_6319);
nor U8475 (N_8475,N_7292,N_7179);
or U8476 (N_8476,N_7250,N_6804);
nand U8477 (N_8477,N_7129,N_6861);
nor U8478 (N_8478,N_6268,N_7217);
xor U8479 (N_8479,N_6102,N_7097);
nand U8480 (N_8480,N_6187,N_6624);
nor U8481 (N_8481,N_7430,N_7301);
xor U8482 (N_8482,N_7382,N_6272);
and U8483 (N_8483,N_6141,N_6556);
nand U8484 (N_8484,N_6162,N_6338);
xor U8485 (N_8485,N_6085,N_7126);
xnor U8486 (N_8486,N_6629,N_6942);
or U8487 (N_8487,N_7119,N_6068);
xor U8488 (N_8488,N_6909,N_6297);
nand U8489 (N_8489,N_6632,N_6542);
nand U8490 (N_8490,N_6077,N_7036);
nor U8491 (N_8491,N_6394,N_6012);
or U8492 (N_8492,N_6861,N_6113);
xnor U8493 (N_8493,N_7494,N_6094);
and U8494 (N_8494,N_6152,N_6907);
xnor U8495 (N_8495,N_6562,N_6200);
nand U8496 (N_8496,N_6320,N_6400);
and U8497 (N_8497,N_6915,N_7354);
xor U8498 (N_8498,N_6632,N_6199);
nor U8499 (N_8499,N_6075,N_7064);
and U8500 (N_8500,N_6821,N_7154);
nor U8501 (N_8501,N_6171,N_7363);
or U8502 (N_8502,N_6340,N_7141);
and U8503 (N_8503,N_6244,N_6621);
and U8504 (N_8504,N_7461,N_6872);
nand U8505 (N_8505,N_7076,N_7307);
nor U8506 (N_8506,N_6056,N_6772);
and U8507 (N_8507,N_7384,N_6372);
and U8508 (N_8508,N_6264,N_6583);
or U8509 (N_8509,N_6690,N_6373);
nand U8510 (N_8510,N_6385,N_6239);
or U8511 (N_8511,N_6044,N_7011);
and U8512 (N_8512,N_6533,N_6153);
nor U8513 (N_8513,N_6834,N_7235);
nor U8514 (N_8514,N_6843,N_6014);
xnor U8515 (N_8515,N_6616,N_6238);
nor U8516 (N_8516,N_7199,N_6039);
nand U8517 (N_8517,N_6389,N_6091);
or U8518 (N_8518,N_6452,N_6184);
or U8519 (N_8519,N_6122,N_7493);
nand U8520 (N_8520,N_7376,N_7284);
xnor U8521 (N_8521,N_6706,N_7242);
xnor U8522 (N_8522,N_6169,N_7452);
or U8523 (N_8523,N_7350,N_6604);
nand U8524 (N_8524,N_6298,N_6417);
nor U8525 (N_8525,N_6768,N_7491);
nor U8526 (N_8526,N_6626,N_7390);
and U8527 (N_8527,N_7069,N_7207);
and U8528 (N_8528,N_7212,N_6071);
xnor U8529 (N_8529,N_6905,N_6171);
nor U8530 (N_8530,N_7490,N_6711);
or U8531 (N_8531,N_7176,N_6670);
nand U8532 (N_8532,N_6187,N_7338);
xor U8533 (N_8533,N_6370,N_6015);
or U8534 (N_8534,N_6373,N_7087);
nand U8535 (N_8535,N_6967,N_7492);
xor U8536 (N_8536,N_6095,N_6754);
or U8537 (N_8537,N_7369,N_6523);
or U8538 (N_8538,N_6617,N_7099);
and U8539 (N_8539,N_6828,N_6540);
and U8540 (N_8540,N_7375,N_6876);
xnor U8541 (N_8541,N_6934,N_6799);
nand U8542 (N_8542,N_6701,N_7126);
nand U8543 (N_8543,N_7020,N_6447);
nand U8544 (N_8544,N_6381,N_6510);
nor U8545 (N_8545,N_7241,N_7456);
or U8546 (N_8546,N_6479,N_6304);
nand U8547 (N_8547,N_6252,N_6103);
or U8548 (N_8548,N_7240,N_6814);
nor U8549 (N_8549,N_6623,N_6018);
xor U8550 (N_8550,N_6074,N_6966);
nand U8551 (N_8551,N_7367,N_6589);
nand U8552 (N_8552,N_7471,N_7146);
or U8553 (N_8553,N_6908,N_7026);
nand U8554 (N_8554,N_7071,N_6496);
and U8555 (N_8555,N_6793,N_7035);
nand U8556 (N_8556,N_6117,N_7341);
nor U8557 (N_8557,N_7267,N_6196);
and U8558 (N_8558,N_6284,N_6128);
nand U8559 (N_8559,N_6052,N_6539);
xnor U8560 (N_8560,N_6796,N_7234);
or U8561 (N_8561,N_6869,N_7454);
nand U8562 (N_8562,N_7229,N_7460);
xnor U8563 (N_8563,N_6666,N_7474);
xor U8564 (N_8564,N_7466,N_6574);
nand U8565 (N_8565,N_6743,N_7018);
nand U8566 (N_8566,N_6521,N_7100);
nor U8567 (N_8567,N_6138,N_7380);
and U8568 (N_8568,N_6946,N_6170);
xor U8569 (N_8569,N_6075,N_6436);
xor U8570 (N_8570,N_7427,N_6893);
and U8571 (N_8571,N_6589,N_7198);
nand U8572 (N_8572,N_7003,N_7412);
nor U8573 (N_8573,N_6579,N_7450);
nand U8574 (N_8574,N_6071,N_7242);
and U8575 (N_8575,N_7445,N_7150);
or U8576 (N_8576,N_7242,N_7213);
and U8577 (N_8577,N_6759,N_6108);
xnor U8578 (N_8578,N_6161,N_7256);
xor U8579 (N_8579,N_7062,N_6296);
nor U8580 (N_8580,N_7182,N_6212);
nor U8581 (N_8581,N_6062,N_7244);
or U8582 (N_8582,N_6092,N_6536);
nor U8583 (N_8583,N_6164,N_7095);
and U8584 (N_8584,N_6661,N_7321);
or U8585 (N_8585,N_7328,N_6662);
nand U8586 (N_8586,N_6423,N_7230);
nand U8587 (N_8587,N_7222,N_7168);
and U8588 (N_8588,N_6845,N_7248);
xor U8589 (N_8589,N_6635,N_7466);
xor U8590 (N_8590,N_6147,N_7424);
and U8591 (N_8591,N_6666,N_6236);
xor U8592 (N_8592,N_7263,N_6828);
xnor U8593 (N_8593,N_7193,N_6153);
nor U8594 (N_8594,N_6874,N_6319);
nand U8595 (N_8595,N_6619,N_6585);
nand U8596 (N_8596,N_6018,N_6461);
xnor U8597 (N_8597,N_6842,N_6699);
nor U8598 (N_8598,N_7354,N_7305);
xnor U8599 (N_8599,N_6740,N_6478);
nand U8600 (N_8600,N_6609,N_6092);
or U8601 (N_8601,N_6425,N_6637);
xnor U8602 (N_8602,N_7101,N_7090);
or U8603 (N_8603,N_7000,N_6662);
nand U8604 (N_8604,N_6690,N_6743);
xor U8605 (N_8605,N_6122,N_7148);
xor U8606 (N_8606,N_7008,N_6798);
and U8607 (N_8607,N_7322,N_7424);
and U8608 (N_8608,N_7137,N_7362);
xor U8609 (N_8609,N_6705,N_6102);
nor U8610 (N_8610,N_7101,N_7135);
nand U8611 (N_8611,N_6951,N_6838);
or U8612 (N_8612,N_7111,N_6503);
nand U8613 (N_8613,N_6918,N_7448);
nor U8614 (N_8614,N_6405,N_7258);
and U8615 (N_8615,N_7019,N_6755);
and U8616 (N_8616,N_6449,N_7000);
or U8617 (N_8617,N_7298,N_6769);
or U8618 (N_8618,N_7153,N_7129);
nand U8619 (N_8619,N_7377,N_7108);
nand U8620 (N_8620,N_6543,N_7054);
xnor U8621 (N_8621,N_6370,N_6388);
xnor U8622 (N_8622,N_7161,N_6618);
nor U8623 (N_8623,N_6617,N_6969);
or U8624 (N_8624,N_7165,N_7124);
nor U8625 (N_8625,N_7248,N_6835);
nor U8626 (N_8626,N_6370,N_6789);
or U8627 (N_8627,N_6104,N_7052);
xor U8628 (N_8628,N_6348,N_7443);
xor U8629 (N_8629,N_6619,N_7362);
nor U8630 (N_8630,N_6418,N_6933);
or U8631 (N_8631,N_6128,N_7157);
or U8632 (N_8632,N_7388,N_6173);
nor U8633 (N_8633,N_6998,N_7454);
nand U8634 (N_8634,N_6046,N_6702);
xor U8635 (N_8635,N_6088,N_6268);
or U8636 (N_8636,N_6520,N_6098);
xnor U8637 (N_8637,N_6938,N_7180);
nor U8638 (N_8638,N_6501,N_7322);
or U8639 (N_8639,N_6194,N_6477);
nor U8640 (N_8640,N_7226,N_6857);
nor U8641 (N_8641,N_6721,N_6498);
and U8642 (N_8642,N_6738,N_7282);
and U8643 (N_8643,N_6467,N_6659);
or U8644 (N_8644,N_6895,N_6540);
nand U8645 (N_8645,N_7275,N_6303);
xor U8646 (N_8646,N_7032,N_6265);
nand U8647 (N_8647,N_6518,N_6822);
or U8648 (N_8648,N_7489,N_6614);
and U8649 (N_8649,N_7271,N_6641);
and U8650 (N_8650,N_6636,N_6627);
and U8651 (N_8651,N_7347,N_6122);
xor U8652 (N_8652,N_7410,N_6936);
or U8653 (N_8653,N_6336,N_7323);
nand U8654 (N_8654,N_7276,N_6718);
xor U8655 (N_8655,N_7355,N_7391);
and U8656 (N_8656,N_7481,N_6211);
xor U8657 (N_8657,N_6266,N_7275);
and U8658 (N_8658,N_6402,N_6393);
or U8659 (N_8659,N_6279,N_6344);
and U8660 (N_8660,N_6752,N_6338);
or U8661 (N_8661,N_6990,N_6100);
nand U8662 (N_8662,N_6274,N_6736);
or U8663 (N_8663,N_6599,N_6489);
and U8664 (N_8664,N_6883,N_6050);
and U8665 (N_8665,N_6001,N_6851);
or U8666 (N_8666,N_6621,N_6333);
xor U8667 (N_8667,N_7442,N_6157);
xnor U8668 (N_8668,N_6526,N_7295);
nor U8669 (N_8669,N_6631,N_6679);
or U8670 (N_8670,N_6022,N_6444);
xnor U8671 (N_8671,N_7159,N_6353);
nor U8672 (N_8672,N_7339,N_7133);
nor U8673 (N_8673,N_6383,N_7217);
xnor U8674 (N_8674,N_7153,N_6778);
nor U8675 (N_8675,N_6447,N_6265);
or U8676 (N_8676,N_7055,N_6749);
and U8677 (N_8677,N_7477,N_7094);
and U8678 (N_8678,N_6197,N_6256);
nor U8679 (N_8679,N_7216,N_6447);
nand U8680 (N_8680,N_6467,N_6510);
nand U8681 (N_8681,N_7138,N_6732);
and U8682 (N_8682,N_7000,N_7465);
and U8683 (N_8683,N_6464,N_6024);
and U8684 (N_8684,N_7114,N_7342);
nand U8685 (N_8685,N_7136,N_7134);
nor U8686 (N_8686,N_7292,N_6152);
and U8687 (N_8687,N_7367,N_6314);
and U8688 (N_8688,N_7194,N_7141);
nor U8689 (N_8689,N_6202,N_7117);
nor U8690 (N_8690,N_6604,N_6340);
nor U8691 (N_8691,N_6449,N_7352);
xnor U8692 (N_8692,N_6828,N_7172);
nand U8693 (N_8693,N_6308,N_7111);
nor U8694 (N_8694,N_7211,N_6503);
and U8695 (N_8695,N_6608,N_6934);
and U8696 (N_8696,N_6938,N_6886);
nand U8697 (N_8697,N_7424,N_6008);
nand U8698 (N_8698,N_7119,N_6440);
xor U8699 (N_8699,N_7302,N_7180);
nand U8700 (N_8700,N_7303,N_7157);
xor U8701 (N_8701,N_6881,N_6528);
nand U8702 (N_8702,N_6263,N_6222);
nand U8703 (N_8703,N_7150,N_7251);
and U8704 (N_8704,N_6612,N_7342);
xor U8705 (N_8705,N_7031,N_6812);
or U8706 (N_8706,N_6975,N_7010);
nor U8707 (N_8707,N_7392,N_7165);
nand U8708 (N_8708,N_6449,N_7134);
nand U8709 (N_8709,N_6079,N_6169);
nor U8710 (N_8710,N_6563,N_7282);
or U8711 (N_8711,N_7161,N_7473);
xnor U8712 (N_8712,N_7058,N_7440);
or U8713 (N_8713,N_6718,N_6555);
nor U8714 (N_8714,N_6874,N_7409);
xor U8715 (N_8715,N_6960,N_6468);
or U8716 (N_8716,N_7172,N_6339);
xor U8717 (N_8717,N_6652,N_7125);
nand U8718 (N_8718,N_6893,N_6192);
nor U8719 (N_8719,N_6605,N_6156);
nand U8720 (N_8720,N_6146,N_7444);
or U8721 (N_8721,N_6066,N_6565);
nand U8722 (N_8722,N_6148,N_6158);
xor U8723 (N_8723,N_6845,N_7476);
or U8724 (N_8724,N_6946,N_6389);
xor U8725 (N_8725,N_7167,N_7378);
or U8726 (N_8726,N_6728,N_7287);
nand U8727 (N_8727,N_7364,N_6020);
xor U8728 (N_8728,N_6270,N_6364);
xor U8729 (N_8729,N_7282,N_7462);
nor U8730 (N_8730,N_6769,N_6490);
nand U8731 (N_8731,N_7029,N_6719);
nor U8732 (N_8732,N_6012,N_6744);
xnor U8733 (N_8733,N_6382,N_6119);
or U8734 (N_8734,N_6659,N_6680);
nor U8735 (N_8735,N_7459,N_6318);
or U8736 (N_8736,N_6674,N_6579);
and U8737 (N_8737,N_6515,N_6333);
xnor U8738 (N_8738,N_7270,N_6104);
xor U8739 (N_8739,N_6473,N_6061);
nand U8740 (N_8740,N_7095,N_6788);
and U8741 (N_8741,N_6572,N_6124);
nor U8742 (N_8742,N_6813,N_6096);
xnor U8743 (N_8743,N_6572,N_6693);
and U8744 (N_8744,N_6661,N_6328);
xor U8745 (N_8745,N_6367,N_6546);
nor U8746 (N_8746,N_6480,N_6309);
nor U8747 (N_8747,N_6637,N_6847);
or U8748 (N_8748,N_7221,N_6680);
and U8749 (N_8749,N_6975,N_7391);
xnor U8750 (N_8750,N_6170,N_6238);
and U8751 (N_8751,N_7135,N_6377);
nor U8752 (N_8752,N_6296,N_7102);
nand U8753 (N_8753,N_6140,N_6740);
xor U8754 (N_8754,N_6274,N_7018);
or U8755 (N_8755,N_6470,N_7263);
or U8756 (N_8756,N_6567,N_6260);
xor U8757 (N_8757,N_6821,N_6759);
nand U8758 (N_8758,N_6287,N_7043);
xor U8759 (N_8759,N_7015,N_7189);
nor U8760 (N_8760,N_7035,N_6819);
xnor U8761 (N_8761,N_6878,N_6081);
nand U8762 (N_8762,N_6418,N_6654);
nor U8763 (N_8763,N_6841,N_6276);
or U8764 (N_8764,N_6314,N_6684);
and U8765 (N_8765,N_7374,N_6835);
nand U8766 (N_8766,N_6122,N_7260);
nor U8767 (N_8767,N_7011,N_6318);
or U8768 (N_8768,N_6385,N_6145);
or U8769 (N_8769,N_6000,N_7283);
or U8770 (N_8770,N_6477,N_6396);
and U8771 (N_8771,N_6298,N_7084);
nand U8772 (N_8772,N_7425,N_6176);
and U8773 (N_8773,N_6833,N_7032);
nor U8774 (N_8774,N_6687,N_6086);
xor U8775 (N_8775,N_7131,N_6085);
or U8776 (N_8776,N_7095,N_6641);
xor U8777 (N_8777,N_6573,N_7477);
or U8778 (N_8778,N_6748,N_6255);
nand U8779 (N_8779,N_6695,N_7490);
nand U8780 (N_8780,N_7289,N_6345);
and U8781 (N_8781,N_7254,N_6664);
xnor U8782 (N_8782,N_6595,N_6467);
xnor U8783 (N_8783,N_7253,N_7391);
and U8784 (N_8784,N_6060,N_6353);
nor U8785 (N_8785,N_6207,N_7139);
nor U8786 (N_8786,N_6490,N_6598);
xnor U8787 (N_8787,N_7491,N_7421);
or U8788 (N_8788,N_7415,N_6316);
nand U8789 (N_8789,N_6532,N_7187);
nand U8790 (N_8790,N_7100,N_6579);
or U8791 (N_8791,N_6811,N_7433);
xnor U8792 (N_8792,N_6562,N_6649);
and U8793 (N_8793,N_7030,N_6990);
nor U8794 (N_8794,N_7496,N_6286);
or U8795 (N_8795,N_7053,N_6879);
nor U8796 (N_8796,N_7145,N_6888);
nor U8797 (N_8797,N_6054,N_6804);
nand U8798 (N_8798,N_6764,N_6682);
and U8799 (N_8799,N_6098,N_6530);
nor U8800 (N_8800,N_7032,N_6101);
and U8801 (N_8801,N_7011,N_7133);
and U8802 (N_8802,N_6347,N_7389);
and U8803 (N_8803,N_6273,N_6472);
and U8804 (N_8804,N_6899,N_6771);
nor U8805 (N_8805,N_7363,N_6893);
xor U8806 (N_8806,N_7137,N_7310);
and U8807 (N_8807,N_6522,N_6885);
nand U8808 (N_8808,N_7310,N_6734);
or U8809 (N_8809,N_6391,N_6713);
nor U8810 (N_8810,N_6543,N_6965);
nand U8811 (N_8811,N_6893,N_7491);
and U8812 (N_8812,N_7319,N_7420);
and U8813 (N_8813,N_6612,N_6275);
nand U8814 (N_8814,N_6203,N_6522);
nor U8815 (N_8815,N_6730,N_7062);
xnor U8816 (N_8816,N_6351,N_7039);
and U8817 (N_8817,N_6297,N_6978);
or U8818 (N_8818,N_6818,N_7377);
and U8819 (N_8819,N_6814,N_6737);
or U8820 (N_8820,N_7471,N_6169);
and U8821 (N_8821,N_7487,N_7309);
nand U8822 (N_8822,N_6519,N_6796);
or U8823 (N_8823,N_6595,N_7364);
nand U8824 (N_8824,N_7207,N_6349);
or U8825 (N_8825,N_6909,N_6204);
xnor U8826 (N_8826,N_6484,N_6769);
and U8827 (N_8827,N_6228,N_6012);
xnor U8828 (N_8828,N_6725,N_6540);
nand U8829 (N_8829,N_6902,N_7050);
or U8830 (N_8830,N_7119,N_6584);
or U8831 (N_8831,N_7404,N_6920);
xnor U8832 (N_8832,N_6943,N_7364);
and U8833 (N_8833,N_6547,N_6119);
nand U8834 (N_8834,N_6211,N_6265);
or U8835 (N_8835,N_7262,N_6275);
nor U8836 (N_8836,N_7334,N_6678);
or U8837 (N_8837,N_7016,N_6586);
nor U8838 (N_8838,N_6608,N_7076);
or U8839 (N_8839,N_6095,N_6199);
xnor U8840 (N_8840,N_6512,N_6014);
or U8841 (N_8841,N_6157,N_7346);
xnor U8842 (N_8842,N_7170,N_7407);
xnor U8843 (N_8843,N_7474,N_6087);
nand U8844 (N_8844,N_6487,N_7014);
or U8845 (N_8845,N_6769,N_6873);
nand U8846 (N_8846,N_6373,N_6727);
nand U8847 (N_8847,N_6936,N_6500);
and U8848 (N_8848,N_6776,N_6530);
and U8849 (N_8849,N_6525,N_6613);
nand U8850 (N_8850,N_6726,N_7485);
nor U8851 (N_8851,N_6003,N_7393);
nand U8852 (N_8852,N_6573,N_6919);
xnor U8853 (N_8853,N_7447,N_6326);
nand U8854 (N_8854,N_7456,N_7134);
xnor U8855 (N_8855,N_7238,N_6776);
and U8856 (N_8856,N_7389,N_6825);
and U8857 (N_8857,N_6530,N_6819);
nor U8858 (N_8858,N_7402,N_7440);
or U8859 (N_8859,N_7344,N_7192);
nor U8860 (N_8860,N_6052,N_6718);
xnor U8861 (N_8861,N_7253,N_7460);
or U8862 (N_8862,N_6374,N_7101);
or U8863 (N_8863,N_7173,N_6546);
xor U8864 (N_8864,N_7094,N_6088);
nor U8865 (N_8865,N_6371,N_6538);
nand U8866 (N_8866,N_6301,N_6843);
and U8867 (N_8867,N_7478,N_6471);
xnor U8868 (N_8868,N_7321,N_7051);
or U8869 (N_8869,N_7021,N_7037);
and U8870 (N_8870,N_6585,N_6035);
nand U8871 (N_8871,N_7428,N_6224);
xnor U8872 (N_8872,N_7369,N_7340);
or U8873 (N_8873,N_6239,N_7256);
and U8874 (N_8874,N_6786,N_6433);
or U8875 (N_8875,N_6064,N_7093);
and U8876 (N_8876,N_6408,N_7303);
nand U8877 (N_8877,N_7054,N_6656);
and U8878 (N_8878,N_6302,N_6157);
nor U8879 (N_8879,N_7059,N_6956);
and U8880 (N_8880,N_6189,N_6289);
and U8881 (N_8881,N_7149,N_7387);
nor U8882 (N_8882,N_6883,N_6973);
and U8883 (N_8883,N_6615,N_6792);
and U8884 (N_8884,N_7396,N_6094);
or U8885 (N_8885,N_7006,N_6904);
nand U8886 (N_8886,N_6802,N_6467);
nand U8887 (N_8887,N_6802,N_6615);
xor U8888 (N_8888,N_6140,N_6963);
and U8889 (N_8889,N_6631,N_6866);
nor U8890 (N_8890,N_7154,N_6997);
nand U8891 (N_8891,N_6783,N_6247);
nor U8892 (N_8892,N_7254,N_7413);
nor U8893 (N_8893,N_6364,N_7429);
xnor U8894 (N_8894,N_7196,N_6871);
or U8895 (N_8895,N_7409,N_6039);
or U8896 (N_8896,N_6871,N_6063);
or U8897 (N_8897,N_7320,N_6847);
nand U8898 (N_8898,N_6029,N_6467);
nor U8899 (N_8899,N_6019,N_6141);
xnor U8900 (N_8900,N_7059,N_6271);
xor U8901 (N_8901,N_7398,N_6415);
nor U8902 (N_8902,N_6774,N_6681);
nand U8903 (N_8903,N_7292,N_7433);
xnor U8904 (N_8904,N_7114,N_7270);
nor U8905 (N_8905,N_6204,N_6690);
nor U8906 (N_8906,N_7070,N_6610);
or U8907 (N_8907,N_6331,N_7144);
and U8908 (N_8908,N_7231,N_6789);
nand U8909 (N_8909,N_7028,N_7372);
or U8910 (N_8910,N_6150,N_7334);
xor U8911 (N_8911,N_6264,N_6796);
and U8912 (N_8912,N_7466,N_6968);
nor U8913 (N_8913,N_7444,N_6125);
nand U8914 (N_8914,N_7025,N_6930);
or U8915 (N_8915,N_6924,N_6506);
or U8916 (N_8916,N_6795,N_7084);
nor U8917 (N_8917,N_6075,N_6396);
or U8918 (N_8918,N_6889,N_6308);
nor U8919 (N_8919,N_7433,N_6727);
and U8920 (N_8920,N_6336,N_6206);
nor U8921 (N_8921,N_6152,N_7034);
xnor U8922 (N_8922,N_7326,N_7144);
xor U8923 (N_8923,N_6293,N_6451);
or U8924 (N_8924,N_6824,N_7122);
xnor U8925 (N_8925,N_6064,N_7405);
or U8926 (N_8926,N_6926,N_6475);
xor U8927 (N_8927,N_6248,N_6168);
nand U8928 (N_8928,N_6697,N_6288);
nand U8929 (N_8929,N_6375,N_7479);
and U8930 (N_8930,N_6794,N_6228);
xor U8931 (N_8931,N_6513,N_6028);
xor U8932 (N_8932,N_7374,N_6362);
nor U8933 (N_8933,N_6903,N_7017);
nor U8934 (N_8934,N_7419,N_7347);
xnor U8935 (N_8935,N_6214,N_6989);
nor U8936 (N_8936,N_6279,N_7047);
xor U8937 (N_8937,N_7436,N_6723);
xnor U8938 (N_8938,N_7446,N_6164);
nor U8939 (N_8939,N_7190,N_6844);
or U8940 (N_8940,N_6908,N_6370);
and U8941 (N_8941,N_6170,N_7374);
nor U8942 (N_8942,N_6545,N_6897);
and U8943 (N_8943,N_7157,N_6680);
nand U8944 (N_8944,N_6447,N_6949);
or U8945 (N_8945,N_7366,N_6542);
and U8946 (N_8946,N_6363,N_6748);
xor U8947 (N_8947,N_6755,N_6088);
or U8948 (N_8948,N_6952,N_7317);
xor U8949 (N_8949,N_7339,N_7235);
nor U8950 (N_8950,N_6754,N_6005);
or U8951 (N_8951,N_6533,N_7301);
xnor U8952 (N_8952,N_6864,N_7414);
or U8953 (N_8953,N_7463,N_6546);
nand U8954 (N_8954,N_6349,N_6905);
nor U8955 (N_8955,N_6766,N_6218);
or U8956 (N_8956,N_7051,N_6352);
and U8957 (N_8957,N_6312,N_6762);
nor U8958 (N_8958,N_6912,N_7081);
nand U8959 (N_8959,N_6824,N_6199);
nor U8960 (N_8960,N_7295,N_7273);
or U8961 (N_8961,N_7417,N_6534);
xor U8962 (N_8962,N_6069,N_6379);
and U8963 (N_8963,N_6536,N_7007);
and U8964 (N_8964,N_6016,N_7242);
nor U8965 (N_8965,N_7226,N_6608);
xnor U8966 (N_8966,N_7467,N_6193);
nor U8967 (N_8967,N_6236,N_7254);
nor U8968 (N_8968,N_6921,N_6393);
and U8969 (N_8969,N_7125,N_6836);
xor U8970 (N_8970,N_6969,N_6330);
xor U8971 (N_8971,N_6640,N_7439);
or U8972 (N_8972,N_6049,N_6367);
nand U8973 (N_8973,N_6941,N_6592);
nor U8974 (N_8974,N_6755,N_7130);
nand U8975 (N_8975,N_6795,N_7400);
nor U8976 (N_8976,N_6739,N_6773);
nand U8977 (N_8977,N_7305,N_6884);
nand U8978 (N_8978,N_7318,N_6299);
nand U8979 (N_8979,N_7133,N_6863);
nand U8980 (N_8980,N_6157,N_7421);
nand U8981 (N_8981,N_7004,N_6661);
nor U8982 (N_8982,N_7352,N_7326);
or U8983 (N_8983,N_7181,N_6056);
and U8984 (N_8984,N_6314,N_7021);
nor U8985 (N_8985,N_6759,N_6664);
xor U8986 (N_8986,N_7127,N_7073);
nand U8987 (N_8987,N_6576,N_6071);
and U8988 (N_8988,N_6269,N_6613);
nor U8989 (N_8989,N_6617,N_7162);
xor U8990 (N_8990,N_6458,N_6340);
nand U8991 (N_8991,N_7111,N_6472);
or U8992 (N_8992,N_6535,N_7010);
xnor U8993 (N_8993,N_7001,N_7295);
and U8994 (N_8994,N_7176,N_7425);
nand U8995 (N_8995,N_6973,N_6653);
and U8996 (N_8996,N_6698,N_6348);
or U8997 (N_8997,N_6518,N_6782);
or U8998 (N_8998,N_7282,N_6379);
xnor U8999 (N_8999,N_6498,N_6655);
xnor U9000 (N_9000,N_8694,N_7860);
nand U9001 (N_9001,N_8228,N_8376);
or U9002 (N_9002,N_8186,N_8935);
or U9003 (N_9003,N_7530,N_7780);
nor U9004 (N_9004,N_7713,N_8462);
or U9005 (N_9005,N_8374,N_7735);
or U9006 (N_9006,N_8303,N_8050);
nand U9007 (N_9007,N_8887,N_7580);
and U9008 (N_9008,N_8721,N_8889);
and U9009 (N_9009,N_7682,N_7851);
and U9010 (N_9010,N_7595,N_8018);
nand U9011 (N_9011,N_8079,N_8795);
nand U9012 (N_9012,N_8827,N_8443);
nand U9013 (N_9013,N_8032,N_8099);
nor U9014 (N_9014,N_8354,N_7912);
nor U9015 (N_9015,N_8253,N_7862);
xnor U9016 (N_9016,N_7703,N_7610);
and U9017 (N_9017,N_7736,N_8541);
and U9018 (N_9018,N_8966,N_7650);
or U9019 (N_9019,N_8671,N_8956);
xnor U9020 (N_9020,N_7819,N_8092);
xor U9021 (N_9021,N_8572,N_8449);
nand U9022 (N_9022,N_7627,N_8038);
nand U9023 (N_9023,N_7845,N_8825);
nand U9024 (N_9024,N_7803,N_8182);
and U9025 (N_9025,N_7984,N_8703);
or U9026 (N_9026,N_8548,N_7507);
nor U9027 (N_9027,N_8619,N_8237);
and U9028 (N_9028,N_7747,N_8390);
xor U9029 (N_9029,N_8418,N_8134);
or U9030 (N_9030,N_7714,N_7718);
nand U9031 (N_9031,N_8755,N_7857);
or U9032 (N_9032,N_8178,N_7756);
and U9033 (N_9033,N_7670,N_8869);
xor U9034 (N_9034,N_7847,N_8275);
or U9035 (N_9035,N_8080,N_7503);
nand U9036 (N_9036,N_8739,N_7581);
nor U9037 (N_9037,N_7568,N_8738);
nor U9038 (N_9038,N_8817,N_8709);
nor U9039 (N_9039,N_7908,N_7547);
nor U9040 (N_9040,N_7890,N_8369);
and U9041 (N_9041,N_8782,N_7935);
nor U9042 (N_9042,N_8534,N_7828);
and U9043 (N_9043,N_8302,N_7525);
xor U9044 (N_9044,N_8898,N_8830);
nand U9045 (N_9045,N_7611,N_8505);
and U9046 (N_9046,N_7913,N_7877);
and U9047 (N_9047,N_7961,N_8125);
nand U9048 (N_9048,N_7830,N_7769);
and U9049 (N_9049,N_8024,N_8300);
or U9050 (N_9050,N_8364,N_8413);
or U9051 (N_9051,N_8072,N_8326);
or U9052 (N_9052,N_8392,N_7812);
xor U9053 (N_9053,N_7757,N_8803);
nand U9054 (N_9054,N_8381,N_7986);
and U9055 (N_9055,N_7881,N_8842);
nor U9056 (N_9056,N_7844,N_8144);
and U9057 (N_9057,N_8289,N_8028);
and U9058 (N_9058,N_8566,N_8511);
nand U9059 (N_9059,N_8547,N_8821);
and U9060 (N_9060,N_7774,N_8805);
or U9061 (N_9061,N_8532,N_7596);
nor U9062 (N_9062,N_8812,N_7576);
or U9063 (N_9063,N_8840,N_8508);
or U9064 (N_9064,N_7981,N_8081);
and U9065 (N_9065,N_7560,N_7741);
xnor U9066 (N_9066,N_8603,N_7527);
and U9067 (N_9067,N_8873,N_7737);
nand U9068 (N_9068,N_8398,N_8098);
and U9069 (N_9069,N_8667,N_8843);
nor U9070 (N_9070,N_8618,N_8758);
xor U9071 (N_9071,N_8331,N_7658);
and U9072 (N_9072,N_7573,N_8415);
nand U9073 (N_9073,N_8642,N_8191);
nand U9074 (N_9074,N_8991,N_8939);
and U9075 (N_9075,N_7708,N_7827);
nand U9076 (N_9076,N_7927,N_8052);
nand U9077 (N_9077,N_8702,N_8067);
nor U9078 (N_9078,N_8714,N_8586);
nor U9079 (N_9079,N_8617,N_7592);
xor U9080 (N_9080,N_7975,N_7821);
nor U9081 (N_9081,N_8061,N_8672);
xor U9082 (N_9082,N_7716,N_8922);
xnor U9083 (N_9083,N_8864,N_7623);
and U9084 (N_9084,N_8652,N_7807);
or U9085 (N_9085,N_8324,N_7502);
nand U9086 (N_9086,N_8666,N_8199);
xnor U9087 (N_9087,N_8635,N_7938);
or U9088 (N_9088,N_7782,N_7802);
or U9089 (N_9089,N_8330,N_8184);
nand U9090 (N_9090,N_8095,N_8035);
nand U9091 (N_9091,N_8172,N_7850);
or U9092 (N_9092,N_8693,N_7750);
nor U9093 (N_9093,N_8342,N_8501);
or U9094 (N_9094,N_8692,N_7659);
nand U9095 (N_9095,N_8409,N_8202);
xnor U9096 (N_9096,N_8114,N_7691);
xnor U9097 (N_9097,N_8733,N_7728);
nor U9098 (N_9098,N_8744,N_8433);
xnor U9099 (N_9099,N_8411,N_8814);
nor U9100 (N_9100,N_8216,N_7668);
xor U9101 (N_9101,N_7848,N_8489);
xor U9102 (N_9102,N_8159,N_8696);
or U9103 (N_9103,N_8767,N_8707);
or U9104 (N_9104,N_8871,N_7726);
xnor U9105 (N_9105,N_8565,N_7826);
and U9106 (N_9106,N_8288,N_8798);
or U9107 (N_9107,N_8404,N_8245);
nand U9108 (N_9108,N_8620,N_8244);
or U9109 (N_9109,N_8160,N_7515);
or U9110 (N_9110,N_8256,N_8003);
or U9111 (N_9111,N_8664,N_8914);
nand U9112 (N_9112,N_8025,N_7787);
xnor U9113 (N_9113,N_7964,N_7727);
nand U9114 (N_9114,N_8568,N_8529);
nand U9115 (N_9115,N_8950,N_8234);
nor U9116 (N_9116,N_8713,N_8639);
xnor U9117 (N_9117,N_8530,N_7715);
nand U9118 (N_9118,N_8471,N_8021);
xnor U9119 (N_9119,N_7648,N_8044);
xnor U9120 (N_9120,N_8093,N_8488);
xor U9121 (N_9121,N_8339,N_8352);
and U9122 (N_9122,N_7840,N_7865);
and U9123 (N_9123,N_8372,N_8687);
nand U9124 (N_9124,N_8203,N_8185);
and U9125 (N_9125,N_8752,N_8661);
nor U9126 (N_9126,N_8929,N_8011);
xnor U9127 (N_9127,N_7858,N_7838);
nand U9128 (N_9128,N_8453,N_7645);
nor U9129 (N_9129,N_7730,N_7585);
nand U9130 (N_9130,N_8792,N_8150);
xor U9131 (N_9131,N_7810,N_8341);
nor U9132 (N_9132,N_8612,N_7678);
nand U9133 (N_9133,N_7980,N_7696);
xor U9134 (N_9134,N_8347,N_8378);
xor U9135 (N_9135,N_7570,N_7962);
or U9136 (N_9136,N_8883,N_8085);
xnor U9137 (N_9137,N_8148,N_8796);
nor U9138 (N_9138,N_7823,N_8282);
xnor U9139 (N_9139,N_8581,N_8512);
or U9140 (N_9140,N_8304,N_7504);
or U9141 (N_9141,N_8832,N_8408);
xnor U9142 (N_9142,N_7704,N_7720);
xor U9143 (N_9143,N_7545,N_8732);
xnor U9144 (N_9144,N_7534,N_8387);
and U9145 (N_9145,N_7959,N_8167);
nor U9146 (N_9146,N_8906,N_7766);
nor U9147 (N_9147,N_8899,N_8344);
nand U9148 (N_9148,N_7613,N_8560);
nor U9149 (N_9149,N_8957,N_7591);
and U9150 (N_9150,N_8273,N_8868);
xor U9151 (N_9151,N_8502,N_8528);
or U9152 (N_9152,N_7712,N_7542);
xor U9153 (N_9153,N_8087,N_7604);
or U9154 (N_9154,N_8490,N_7921);
nor U9155 (N_9155,N_8031,N_8269);
or U9156 (N_9156,N_8596,N_8059);
or U9157 (N_9157,N_7677,N_8880);
or U9158 (N_9158,N_8001,N_7898);
nand U9159 (N_9159,N_7942,N_8251);
nand U9160 (N_9160,N_8239,N_8622);
xor U9161 (N_9161,N_8046,N_8006);
and U9162 (N_9162,N_8121,N_8007);
or U9163 (N_9163,N_7781,N_8804);
and U9164 (N_9164,N_8473,N_8507);
nand U9165 (N_9165,N_8838,N_8564);
xnor U9166 (N_9166,N_7778,N_8506);
or U9167 (N_9167,N_7761,N_8002);
and U9168 (N_9168,N_8570,N_8708);
and U9169 (N_9169,N_7630,N_7520);
and U9170 (N_9170,N_8466,N_8297);
xor U9171 (N_9171,N_7588,N_7866);
or U9172 (N_9172,N_8075,N_8987);
nand U9173 (N_9173,N_7639,N_8014);
and U9174 (N_9174,N_8437,N_8416);
xor U9175 (N_9175,N_8115,N_7794);
or U9176 (N_9176,N_8766,N_7663);
or U9177 (N_9177,N_8590,N_8686);
nand U9178 (N_9178,N_8695,N_8784);
xnor U9179 (N_9179,N_8246,N_8822);
or U9180 (N_9180,N_8674,N_7894);
nand U9181 (N_9181,N_8478,N_7939);
xor U9182 (N_9182,N_7559,N_8145);
nand U9183 (N_9183,N_8320,N_7614);
or U9184 (N_9184,N_8919,N_7829);
nand U9185 (N_9185,N_8120,N_7552);
nand U9186 (N_9186,N_8673,N_8384);
and U9187 (N_9187,N_7606,N_8557);
nor U9188 (N_9188,N_7979,N_8054);
xor U9189 (N_9189,N_8467,N_8229);
xor U9190 (N_9190,N_8977,N_8625);
or U9191 (N_9191,N_8335,N_7949);
nand U9192 (N_9192,N_8070,N_7690);
nor U9193 (N_9193,N_7952,N_7544);
or U9194 (N_9194,N_7679,N_8894);
nor U9195 (N_9195,N_8811,N_7751);
nor U9196 (N_9196,N_7886,N_8220);
nor U9197 (N_9197,N_8214,N_7738);
or U9198 (N_9198,N_7833,N_7540);
nor U9199 (N_9199,N_8606,N_7876);
or U9200 (N_9200,N_7872,N_7548);
or U9201 (N_9201,N_8600,N_8809);
xor U9202 (N_9202,N_8383,N_8412);
and U9203 (N_9203,N_7667,N_8004);
and U9204 (N_9204,N_8876,N_7764);
nand U9205 (N_9205,N_8238,N_8458);
and U9206 (N_9206,N_8110,N_8662);
xor U9207 (N_9207,N_8360,N_8975);
and U9208 (N_9208,N_7684,N_7638);
or U9209 (N_9209,N_8893,N_7861);
nand U9210 (N_9210,N_8201,N_7644);
and U9211 (N_9211,N_7578,N_7879);
xor U9212 (N_9212,N_8047,N_8469);
or U9213 (N_9213,N_7689,N_7923);
nand U9214 (N_9214,N_8867,N_7887);
and U9215 (N_9215,N_8903,N_8187);
nand U9216 (N_9216,N_8649,N_8902);
xor U9217 (N_9217,N_8648,N_8951);
nand U9218 (N_9218,N_7688,N_7683);
or U9219 (N_9219,N_8980,N_8224);
xnor U9220 (N_9220,N_8104,N_8520);
and U9221 (N_9221,N_7546,N_8040);
nand U9222 (N_9222,N_8858,N_8322);
xor U9223 (N_9223,N_8278,N_7768);
and U9224 (N_9224,N_8371,N_7892);
nor U9225 (N_9225,N_7569,N_8292);
or U9226 (N_9226,N_7918,N_8343);
nor U9227 (N_9227,N_7524,N_8180);
nor U9228 (N_9228,N_7672,N_8853);
nor U9229 (N_9229,N_8386,N_8263);
and U9230 (N_9230,N_7811,N_8475);
or U9231 (N_9231,N_7722,N_8362);
xor U9232 (N_9232,N_8169,N_8571);
nor U9233 (N_9233,N_8112,N_8395);
and U9234 (N_9234,N_8774,N_8117);
nand U9235 (N_9235,N_8680,N_8573);
and U9236 (N_9236,N_8992,N_8118);
xor U9237 (N_9237,N_7759,N_8389);
nor U9238 (N_9238,N_8034,N_8794);
nor U9239 (N_9239,N_8139,N_8773);
nand U9240 (N_9240,N_8497,N_7995);
or U9241 (N_9241,N_8158,N_7501);
and U9242 (N_9242,N_8365,N_8474);
nor U9243 (N_9243,N_8317,N_8585);
xnor U9244 (N_9244,N_8852,N_8623);
nor U9245 (N_9245,N_8682,N_8742);
and U9246 (N_9246,N_8333,N_8720);
nor U9247 (N_9247,N_7919,N_7740);
and U9248 (N_9248,N_8439,N_8097);
and U9249 (N_9249,N_7796,N_8550);
and U9250 (N_9250,N_7705,N_8074);
and U9251 (N_9251,N_7561,N_8311);
or U9252 (N_9252,N_7567,N_7583);
and U9253 (N_9253,N_8525,N_8051);
or U9254 (N_9254,N_8227,N_7752);
xor U9255 (N_9255,N_8928,N_8510);
nand U9256 (N_9256,N_8785,N_7600);
nor U9257 (N_9257,N_8434,N_8319);
or U9258 (N_9258,N_8559,N_7805);
xor U9259 (N_9259,N_7529,N_8751);
and U9260 (N_9260,N_8424,N_7909);
and U9261 (N_9261,N_8663,N_8283);
or U9262 (N_9262,N_8700,N_7863);
nand U9263 (N_9263,N_7601,N_8427);
and U9264 (N_9264,N_8677,N_7748);
nor U9265 (N_9265,N_8770,N_8069);
and U9266 (N_9266,N_7513,N_7603);
or U9267 (N_9267,N_8296,N_8233);
nor U9268 (N_9268,N_8105,N_8829);
and U9269 (N_9269,N_7977,N_7773);
and U9270 (N_9270,N_8900,N_7510);
nand U9271 (N_9271,N_8996,N_7589);
and U9272 (N_9272,N_8351,N_8291);
nand U9273 (N_9273,N_8461,N_7706);
nand U9274 (N_9274,N_8176,N_8135);
nand U9275 (N_9275,N_7744,N_7885);
or U9276 (N_9276,N_7549,N_8388);
xnor U9277 (N_9277,N_8293,N_8281);
nand U9278 (N_9278,N_8665,N_8756);
or U9279 (N_9279,N_8915,N_8310);
or U9280 (N_9280,N_8946,N_8043);
nor U9281 (N_9281,N_7686,N_7695);
xnor U9282 (N_9282,N_8198,N_7932);
nand U9283 (N_9283,N_8940,N_8685);
nor U9284 (N_9284,N_8429,N_8405);
and U9285 (N_9285,N_8918,N_8923);
nor U9286 (N_9286,N_7767,N_8628);
nor U9287 (N_9287,N_7571,N_7822);
or U9288 (N_9288,N_8601,N_7920);
or U9289 (N_9289,N_8621,N_7665);
nand U9290 (N_9290,N_8020,N_7575);
xor U9291 (N_9291,N_7514,N_8219);
nor U9292 (N_9292,N_8740,N_8428);
xnor U9293 (N_9293,N_8598,N_7526);
nor U9294 (N_9294,N_8494,N_8971);
or U9295 (N_9295,N_8523,N_8763);
nor U9296 (N_9296,N_8760,N_8106);
nor U9297 (N_9297,N_8810,N_7924);
and U9298 (N_9298,N_8932,N_8688);
xor U9299 (N_9299,N_7777,N_8057);
and U9300 (N_9300,N_8724,N_8926);
and U9301 (N_9301,N_8726,N_8042);
nand U9302 (N_9302,N_7967,N_8334);
and U9303 (N_9303,N_7558,N_7701);
and U9304 (N_9304,N_8147,N_8772);
or U9305 (N_9305,N_8775,N_8213);
nand U9306 (N_9306,N_7651,N_7929);
or U9307 (N_9307,N_8848,N_7599);
and U9308 (N_9308,N_8062,N_8563);
or U9309 (N_9309,N_8235,N_8470);
or U9310 (N_9310,N_8000,N_8457);
or U9311 (N_9311,N_7901,N_8514);
xor U9312 (N_9312,N_7676,N_8657);
nand U9313 (N_9313,N_8472,N_7572);
or U9314 (N_9314,N_8323,N_8402);
or U9315 (N_9315,N_8353,N_8259);
nand U9316 (N_9316,N_7841,N_8553);
xnor U9317 (N_9317,N_8927,N_7931);
xnor U9318 (N_9318,N_8636,N_8232);
or U9319 (N_9319,N_8985,N_7616);
and U9320 (N_9320,N_8328,N_8196);
or U9321 (N_9321,N_8192,N_7762);
nand U9322 (N_9322,N_8668,N_8123);
nand U9323 (N_9323,N_7903,N_8616);
nor U9324 (N_9324,N_7699,N_8527);
and U9325 (N_9325,N_8254,N_8400);
xnor U9326 (N_9326,N_8790,N_8938);
nor U9327 (N_9327,N_8165,N_7732);
nand U9328 (N_9328,N_7801,N_8998);
nor U9329 (N_9329,N_8500,N_7911);
and U9330 (N_9330,N_8698,N_8277);
or U9331 (N_9331,N_8771,N_8890);
and U9332 (N_9332,N_8498,N_7897);
and U9333 (N_9333,N_8456,N_8911);
nor U9334 (N_9334,N_7790,N_7617);
nand U9335 (N_9335,N_7905,N_8904);
xor U9336 (N_9336,N_7631,N_8460);
and U9337 (N_9337,N_7789,N_7869);
nor U9338 (N_9338,N_7618,N_8325);
xor U9339 (N_9339,N_8264,N_7835);
and U9340 (N_9340,N_8704,N_8200);
and U9341 (N_9341,N_7926,N_7698);
or U9342 (N_9342,N_8096,N_8967);
xnor U9343 (N_9343,N_8068,N_8023);
or U9344 (N_9344,N_8305,N_7673);
or U9345 (N_9345,N_8819,N_8874);
nor U9346 (N_9346,N_8653,N_8654);
nand U9347 (N_9347,N_8857,N_8683);
and U9348 (N_9348,N_8670,N_7936);
nand U9349 (N_9349,N_8438,N_8567);
xor U9350 (N_9350,N_8689,N_7795);
or U9351 (N_9351,N_8716,N_8631);
nand U9352 (N_9352,N_8624,N_8363);
xnor U9353 (N_9353,N_7966,N_7820);
nor U9354 (N_9354,N_7671,N_8077);
and U9355 (N_9355,N_8016,N_7622);
nand U9356 (N_9356,N_7893,N_8820);
or U9357 (N_9357,N_7516,N_8658);
or U9358 (N_9358,N_7993,N_8109);
nor U9359 (N_9359,N_8806,N_8361);
and U9360 (N_9360,N_8982,N_8509);
and U9361 (N_9361,N_8337,N_8850);
and U9362 (N_9362,N_8442,N_8197);
or U9363 (N_9363,N_8808,N_8211);
xnor U9364 (N_9364,N_8964,N_7632);
nor U9365 (N_9365,N_8551,N_8299);
or U9366 (N_9366,N_8161,N_7896);
or U9367 (N_9367,N_8540,N_7710);
or U9368 (N_9368,N_8205,N_8223);
xnor U9369 (N_9369,N_8558,N_8086);
and U9370 (N_9370,N_7958,N_8945);
nor U9371 (N_9371,N_7753,N_8285);
xor U9372 (N_9372,N_8284,N_8513);
nor U9373 (N_9373,N_8249,N_8860);
or U9374 (N_9374,N_7878,N_8406);
xnor U9375 (N_9375,N_7535,N_8204);
or U9376 (N_9376,N_7652,N_8504);
nor U9377 (N_9377,N_8485,N_7649);
nor U9378 (N_9378,N_8878,N_8518);
nand U9379 (N_9379,N_7765,N_8990);
xnor U9380 (N_9380,N_8066,N_8608);
and U9381 (N_9381,N_8613,N_7853);
xor U9382 (N_9382,N_8599,N_8272);
nor U9383 (N_9383,N_8206,N_8454);
nor U9384 (N_9384,N_8749,N_8152);
xor U9385 (N_9385,N_7904,N_8678);
nand U9386 (N_9386,N_7656,N_7808);
nand U9387 (N_9387,N_8717,N_7772);
nor U9388 (N_9388,N_8729,N_8701);
nand U9389 (N_9389,N_8882,N_8725);
or U9390 (N_9390,N_8270,N_7721);
and U9391 (N_9391,N_8242,N_8986);
nand U9392 (N_9392,N_8009,N_8357);
nor U9393 (N_9393,N_7729,N_7839);
nand U9394 (N_9394,N_7587,N_7831);
or U9395 (N_9395,N_8562,N_7989);
xnor U9396 (N_9396,N_8747,N_8884);
xor U9397 (N_9397,N_8955,N_7666);
and U9398 (N_9398,N_7934,N_8157);
xor U9399 (N_9399,N_8949,N_8958);
nand U9400 (N_9400,N_7957,N_8151);
nand U9401 (N_9401,N_7607,N_8816);
or U9402 (N_9402,N_7697,N_8451);
and U9403 (N_9403,N_8156,N_7594);
xor U9404 (N_9404,N_8988,N_8972);
and U9405 (N_9405,N_8602,N_7760);
or U9406 (N_9406,N_8516,N_7797);
and U9407 (N_9407,N_8968,N_8373);
or U9408 (N_9408,N_8421,N_8866);
nand U9409 (N_9409,N_8634,N_8426);
nor U9410 (N_9410,N_8012,N_8491);
nand U9411 (N_9411,N_7621,N_7968);
and U9412 (N_9412,N_8380,N_7798);
and U9413 (N_9413,N_8944,N_8644);
xor U9414 (N_9414,N_8886,N_8247);
or U9415 (N_9415,N_7956,N_7978);
or U9416 (N_9416,N_8979,N_8515);
xor U9417 (N_9417,N_7868,N_7948);
xnor U9418 (N_9418,N_7597,N_8941);
nand U9419 (N_9419,N_8633,N_8286);
and U9420 (N_9420,N_8538,N_8129);
nand U9421 (N_9421,N_8800,N_8005);
or U9422 (N_9422,N_7551,N_8218);
nand U9423 (N_9423,N_7849,N_8268);
nor U9424 (N_9424,N_8423,N_7517);
nor U9425 (N_9425,N_8768,N_8582);
and U9426 (N_9426,N_8676,N_8632);
or U9427 (N_9427,N_8358,N_7537);
nor U9428 (N_9428,N_8791,N_8897);
and U9429 (N_9429,N_8446,N_7916);
or U9430 (N_9430,N_8645,N_8905);
and U9431 (N_9431,N_7799,N_8403);
xnor U9432 (N_9432,N_8124,N_8954);
nand U9433 (N_9433,N_7702,N_7971);
and U9434 (N_9434,N_8119,N_8823);
nand U9435 (N_9435,N_7554,N_8769);
xnor U9436 (N_9436,N_8989,N_8435);
or U9437 (N_9437,N_8807,N_7816);
or U9438 (N_9438,N_8745,N_8391);
or U9439 (N_9439,N_8659,N_8916);
and U9440 (N_9440,N_7654,N_8138);
nor U9441 (N_9441,N_7969,N_8230);
xnor U9442 (N_9442,N_7634,N_8126);
nand U9443 (N_9443,N_8332,N_8855);
and U9444 (N_9444,N_8313,N_8522);
or U9445 (N_9445,N_7859,N_8813);
and U9446 (N_9446,N_8584,N_8545);
nand U9447 (N_9447,N_8789,N_7694);
or U9448 (N_9448,N_7906,N_8496);
nor U9449 (N_9449,N_8824,N_8569);
or U9450 (N_9450,N_7994,N_8452);
or U9451 (N_9451,N_7800,N_8818);
or U9452 (N_9452,N_8177,N_8141);
or U9453 (N_9453,N_8183,N_7937);
nand U9454 (N_9454,N_8041,N_8641);
or U9455 (N_9455,N_7771,N_8710);
nor U9456 (N_9456,N_7974,N_8131);
or U9457 (N_9457,N_8209,N_7963);
nand U9458 (N_9458,N_8195,N_8295);
nor U9459 (N_9459,N_8976,N_7758);
and U9460 (N_9460,N_8103,N_8394);
nor U9461 (N_9461,N_7813,N_8166);
nand U9462 (N_9462,N_7500,N_8013);
xor U9463 (N_9463,N_8217,N_8477);
xor U9464 (N_9464,N_7687,N_8675);
or U9465 (N_9465,N_8519,N_8962);
xor U9466 (N_9466,N_8764,N_7674);
or U9467 (N_9467,N_8948,N_8879);
xnor U9468 (N_9468,N_7528,N_8797);
or U9469 (N_9469,N_8741,N_8039);
nor U9470 (N_9470,N_8901,N_8937);
nand U9471 (N_9471,N_8399,N_8594);
nand U9472 (N_9472,N_7598,N_8350);
or U9473 (N_9473,N_8930,N_8753);
and U9474 (N_9474,N_8626,N_8638);
nand U9475 (N_9475,N_8276,N_8257);
nor U9476 (N_9476,N_8260,N_7999);
or U9477 (N_9477,N_7565,N_8063);
and U9478 (N_9478,N_8073,N_8656);
nand U9479 (N_9479,N_7692,N_8917);
xnor U9480 (N_9480,N_8377,N_7856);
nand U9481 (N_9481,N_8045,N_8348);
nand U9482 (N_9482,N_8318,N_8801);
nor U9483 (N_9483,N_7685,N_7941);
and U9484 (N_9484,N_8761,N_8647);
or U9485 (N_9485,N_8856,N_8107);
nor U9486 (N_9486,N_8910,N_8609);
and U9487 (N_9487,N_8316,N_8091);
or U9488 (N_9488,N_8521,N_8419);
xor U9489 (N_9489,N_7846,N_7635);
nor U9490 (N_9490,N_8370,N_7804);
or U9491 (N_9491,N_7538,N_8846);
nor U9492 (N_9492,N_7985,N_8327);
nor U9493 (N_9493,N_7586,N_8604);
xnor U9494 (N_9494,N_8605,N_8920);
and U9495 (N_9495,N_7745,N_8215);
xor U9496 (N_9496,N_8615,N_7947);
xor U9497 (N_9497,N_8019,N_7824);
or U9498 (N_9498,N_8111,N_8250);
or U9499 (N_9499,N_8430,N_8321);
nor U9500 (N_9500,N_8271,N_7940);
nand U9501 (N_9501,N_8146,N_8963);
xnor U9502 (N_9502,N_8142,N_7628);
nor U9503 (N_9503,N_7990,N_7873);
xnor U9504 (N_9504,N_8484,N_8793);
xnor U9505 (N_9505,N_8925,N_8503);
or U9506 (N_9506,N_8681,N_8844);
or U9507 (N_9507,N_8346,N_7593);
and U9508 (N_9508,N_7700,N_7619);
nor U9509 (N_9509,N_8248,N_8587);
and U9510 (N_9510,N_7953,N_8969);
or U9511 (N_9511,N_8465,N_8546);
nand U9512 (N_9512,N_8274,N_7625);
or U9513 (N_9513,N_8375,N_8891);
and U9514 (N_9514,N_8909,N_7646);
and U9515 (N_9515,N_7577,N_8385);
and U9516 (N_9516,N_7541,N_8459);
and U9517 (N_9517,N_8448,N_8651);
xor U9518 (N_9518,N_7723,N_8715);
nand U9519 (N_9519,N_8450,N_8113);
nand U9520 (N_9520,N_8089,N_7992);
or U9521 (N_9521,N_8854,N_8580);
nand U9522 (N_9522,N_7874,N_8290);
or U9523 (N_9523,N_8684,N_8379);
and U9524 (N_9524,N_8155,N_7950);
nor U9525 (N_9525,N_7556,N_8207);
nor U9526 (N_9526,N_8049,N_8154);
and U9527 (N_9527,N_8583,N_8441);
or U9528 (N_9528,N_7998,N_8912);
nand U9529 (N_9529,N_8646,N_8338);
or U9530 (N_9530,N_8447,N_8163);
and U9531 (N_9531,N_8788,N_8947);
xor U9532 (N_9532,N_8368,N_8776);
nor U9533 (N_9533,N_8464,N_8637);
or U9534 (N_9534,N_8723,N_8179);
or U9535 (N_9535,N_7945,N_7788);
nand U9536 (N_9536,N_8728,N_8895);
nor U9537 (N_9537,N_8863,N_7724);
or U9538 (N_9538,N_8543,N_8595);
and U9539 (N_9539,N_7608,N_8934);
and U9540 (N_9540,N_7605,N_7900);
and U9541 (N_9541,N_8936,N_8100);
and U9542 (N_9542,N_7602,N_8088);
and U9543 (N_9543,N_8978,N_7910);
nor U9544 (N_9544,N_7522,N_7543);
or U9545 (N_9545,N_7566,N_7711);
nor U9546 (N_9546,N_7655,N_8959);
nand U9547 (N_9547,N_8577,N_8588);
nand U9548 (N_9548,N_8487,N_8828);
nand U9549 (N_9549,N_8140,N_8836);
nand U9550 (N_9550,N_8862,N_8189);
nand U9551 (N_9551,N_8190,N_8549);
or U9552 (N_9552,N_8593,N_8679);
nand U9553 (N_9553,N_7505,N_8865);
xnor U9554 (N_9554,N_7664,N_8875);
nor U9555 (N_9555,N_8287,N_7925);
nor U9556 (N_9556,N_7653,N_8690);
xnor U9557 (N_9557,N_7642,N_8839);
xnor U9558 (N_9558,N_7612,N_7834);
or U9559 (N_9559,N_8630,N_8243);
xor U9560 (N_9560,N_7629,N_8425);
xnor U9561 (N_9561,N_8960,N_8255);
nand U9562 (N_9562,N_7982,N_7557);
and U9563 (N_9563,N_7864,N_8555);
or U9564 (N_9564,N_8306,N_7662);
or U9565 (N_9565,N_8885,N_7818);
xor U9566 (N_9566,N_8414,N_8589);
xor U9567 (N_9567,N_7518,N_8143);
xor U9568 (N_9568,N_7996,N_8483);
and U9569 (N_9569,N_8307,N_8759);
nand U9570 (N_9570,N_8065,N_7976);
and U9571 (N_9571,N_7709,N_8783);
and U9572 (N_9572,N_7815,N_7902);
nand U9573 (N_9573,N_7770,N_7883);
or U9574 (N_9574,N_8535,N_7531);
nor U9575 (N_9575,N_8084,N_7755);
nand U9576 (N_9576,N_7533,N_8309);
nor U9577 (N_9577,N_8222,N_7574);
nand U9578 (N_9578,N_8952,N_8090);
nor U9579 (N_9579,N_8640,N_7553);
or U9580 (N_9580,N_7609,N_7707);
nor U9581 (N_9581,N_8815,N_8102);
xor U9582 (N_9582,N_8008,N_8531);
and U9583 (N_9583,N_8942,N_8931);
and U9584 (N_9584,N_8845,N_7637);
nor U9585 (N_9585,N_8961,N_8017);
and U9586 (N_9586,N_8746,N_8877);
and U9587 (N_9587,N_8162,N_8033);
or U9588 (N_9588,N_8750,N_8837);
and U9589 (N_9589,N_7922,N_7640);
xor U9590 (N_9590,N_7965,N_8480);
or U9591 (N_9591,N_8266,N_7523);
and U9592 (N_9592,N_7763,N_8356);
xnor U9593 (N_9593,N_8479,N_7972);
or U9594 (N_9594,N_8101,N_8053);
and U9595 (N_9595,N_7987,N_8533);
nor U9596 (N_9596,N_7582,N_7681);
or U9597 (N_9597,N_8994,N_8280);
or U9598 (N_9598,N_8554,N_8781);
or U9599 (N_9599,N_8279,N_8913);
nand U9600 (N_9600,N_8349,N_8737);
nor U9601 (N_9601,N_7973,N_8336);
and U9602 (N_9602,N_7564,N_8078);
nor U9603 (N_9603,N_8831,N_8226);
nand U9604 (N_9604,N_8777,N_7854);
nor U9605 (N_9605,N_7590,N_7643);
and U9606 (N_9606,N_8431,N_8312);
xnor U9607 (N_9607,N_7754,N_8727);
and U9608 (N_9608,N_8212,N_8921);
or U9609 (N_9609,N_8892,N_8933);
or U9610 (N_9610,N_7930,N_7786);
or U9611 (N_9611,N_8730,N_7842);
and U9612 (N_9612,N_8655,N_8258);
or U9613 (N_9613,N_8896,N_8762);
nor U9614 (N_9614,N_7888,N_8669);
nor U9615 (N_9615,N_8410,N_8340);
nand U9616 (N_9616,N_8517,N_8030);
and U9617 (N_9617,N_8168,N_8181);
xor U9618 (N_9618,N_8736,N_7825);
or U9619 (N_9619,N_8267,N_8924);
xnor U9620 (N_9620,N_8544,N_7809);
nor U9621 (N_9621,N_8444,N_8482);
nor U9622 (N_9622,N_8083,N_8591);
xor U9623 (N_9623,N_8128,N_7717);
nor U9624 (N_9624,N_8122,N_8026);
or U9625 (N_9625,N_8579,N_8943);
or U9626 (N_9626,N_8231,N_7954);
nor U9627 (N_9627,N_8786,N_7743);
nand U9628 (N_9628,N_7512,N_8643);
nor U9629 (N_9629,N_8614,N_8164);
nor U9630 (N_9630,N_8722,N_8973);
or U9631 (N_9631,N_7814,N_8997);
nor U9632 (N_9632,N_8241,N_8436);
and U9633 (N_9633,N_8440,N_7895);
or U9634 (N_9634,N_7508,N_8393);
nor U9635 (N_9635,N_8974,N_8076);
nand U9636 (N_9636,N_7955,N_7855);
nand U9637 (N_9637,N_8711,N_8486);
or U9638 (N_9638,N_7991,N_8748);
nor U9639 (N_9639,N_8455,N_8493);
and U9640 (N_9640,N_8799,N_8308);
or U9641 (N_9641,N_8965,N_7970);
nand U9642 (N_9642,N_8432,N_8366);
xor U9643 (N_9643,N_8757,N_8401);
and U9644 (N_9644,N_8037,N_7867);
xnor U9645 (N_9645,N_7776,N_7615);
or U9646 (N_9646,N_8888,N_7775);
nand U9647 (N_9647,N_8778,N_8022);
and U9648 (N_9648,N_7647,N_8705);
nor U9649 (N_9649,N_8629,N_8208);
xor U9650 (N_9650,N_7960,N_7899);
and U9651 (N_9651,N_8048,N_7836);
and U9652 (N_9652,N_8094,N_8137);
nor U9653 (N_9653,N_8870,N_7792);
or U9654 (N_9654,N_7536,N_7739);
nor U9655 (N_9655,N_8132,N_8420);
xor U9656 (N_9656,N_7946,N_8780);
xnor U9657 (N_9657,N_8610,N_8575);
or U9658 (N_9658,N_7914,N_7783);
and U9659 (N_9659,N_8970,N_8802);
xnor U9660 (N_9660,N_7731,N_8225);
or U9661 (N_9661,N_8849,N_8697);
nand U9662 (N_9662,N_8556,N_7563);
nor U9663 (N_9663,N_7871,N_8881);
or U9664 (N_9664,N_7988,N_7719);
xor U9665 (N_9665,N_7579,N_8301);
xnor U9666 (N_9666,N_8174,N_8542);
nand U9667 (N_9667,N_7785,N_8847);
or U9668 (N_9668,N_7943,N_7793);
or U9669 (N_9669,N_8314,N_8607);
and U9670 (N_9670,N_7519,N_8574);
and U9671 (N_9671,N_8660,N_8153);
xnor U9672 (N_9672,N_8524,N_7669);
xor U9673 (N_9673,N_7742,N_8552);
xnor U9674 (N_9674,N_8834,N_7693);
and U9675 (N_9675,N_8236,N_8526);
nor U9676 (N_9676,N_8699,N_8995);
nand U9677 (N_9677,N_8578,N_8261);
and U9678 (N_9678,N_7870,N_7661);
and U9679 (N_9679,N_8468,N_8481);
nand U9680 (N_9680,N_7915,N_8981);
and U9681 (N_9681,N_7889,N_8127);
xnor U9682 (N_9682,N_8993,N_8765);
and U9683 (N_9683,N_8367,N_8499);
xnor U9684 (N_9684,N_8650,N_8859);
or U9685 (N_9685,N_7791,N_8718);
nand U9686 (N_9686,N_8265,N_7680);
nor U9687 (N_9687,N_7997,N_8627);
nor U9688 (N_9688,N_7928,N_8953);
nor U9689 (N_9689,N_7636,N_8712);
nor U9690 (N_9690,N_8826,N_8445);
nand U9691 (N_9691,N_7675,N_7817);
xor U9692 (N_9692,N_7852,N_8495);
nor U9693 (N_9693,N_7550,N_7733);
xnor U9694 (N_9694,N_7641,N_8058);
or U9695 (N_9695,N_8706,N_7506);
or U9696 (N_9696,N_8060,N_8476);
or U9697 (N_9697,N_8835,N_8315);
or U9698 (N_9698,N_7511,N_8262);
nand U9699 (N_9699,N_8536,N_8329);
or U9700 (N_9700,N_8210,N_7837);
nor U9701 (N_9701,N_8015,N_8984);
or U9702 (N_9702,N_7521,N_7907);
or U9703 (N_9703,N_7832,N_8735);
nor U9704 (N_9704,N_7562,N_8240);
or U9705 (N_9705,N_8734,N_8173);
nand U9706 (N_9706,N_8787,N_7657);
xor U9707 (N_9707,N_8355,N_8833);
or U9708 (N_9708,N_8221,N_8194);
or U9709 (N_9709,N_8908,N_8193);
nand U9710 (N_9710,N_8492,N_7891);
nor U9711 (N_9711,N_8907,N_7509);
nand U9712 (N_9712,N_8064,N_8010);
and U9713 (N_9713,N_8027,N_8754);
and U9714 (N_9714,N_7532,N_7734);
and U9715 (N_9715,N_8397,N_7884);
xnor U9716 (N_9716,N_8691,N_8056);
xor U9717 (N_9717,N_7882,N_7539);
nor U9718 (N_9718,N_8082,N_7555);
and U9719 (N_9719,N_7951,N_7779);
or U9720 (N_9720,N_7917,N_8407);
or U9721 (N_9721,N_7620,N_8731);
and U9722 (N_9722,N_7660,N_8175);
nand U9723 (N_9723,N_7843,N_8861);
xor U9724 (N_9724,N_8872,N_7880);
xor U9725 (N_9725,N_8539,N_8359);
nand U9726 (N_9726,N_8611,N_7624);
and U9727 (N_9727,N_8116,N_8133);
xnor U9728 (N_9728,N_8841,N_7584);
or U9729 (N_9729,N_8136,N_8417);
nor U9730 (N_9730,N_8382,N_7749);
and U9731 (N_9731,N_7633,N_8999);
xor U9732 (N_9732,N_8171,N_8463);
nor U9733 (N_9733,N_8561,N_7806);
and U9734 (N_9734,N_8779,N_8345);
nand U9735 (N_9735,N_8743,N_7725);
nand U9736 (N_9736,N_7784,N_8188);
and U9737 (N_9737,N_8130,N_8422);
or U9738 (N_9738,N_8983,N_8294);
nor U9739 (N_9739,N_8298,N_8071);
nand U9740 (N_9740,N_8396,N_8108);
xor U9741 (N_9741,N_7933,N_8592);
xnor U9742 (N_9742,N_7626,N_7944);
and U9743 (N_9743,N_8576,N_8055);
or U9744 (N_9744,N_8029,N_7746);
nor U9745 (N_9745,N_7875,N_8036);
xor U9746 (N_9746,N_8537,N_8597);
nor U9747 (N_9747,N_7983,N_8170);
and U9748 (N_9748,N_8851,N_8719);
nor U9749 (N_9749,N_8149,N_8252);
and U9750 (N_9750,N_8434,N_7526);
or U9751 (N_9751,N_7874,N_8629);
nor U9752 (N_9752,N_8920,N_8298);
and U9753 (N_9753,N_7645,N_7683);
or U9754 (N_9754,N_8642,N_7800);
and U9755 (N_9755,N_8322,N_8221);
nand U9756 (N_9756,N_8805,N_7933);
or U9757 (N_9757,N_7580,N_7649);
nand U9758 (N_9758,N_8766,N_8093);
or U9759 (N_9759,N_8864,N_8998);
and U9760 (N_9760,N_8089,N_8019);
or U9761 (N_9761,N_8499,N_7589);
nand U9762 (N_9762,N_8845,N_8336);
nand U9763 (N_9763,N_8705,N_7914);
and U9764 (N_9764,N_8844,N_7687);
xnor U9765 (N_9765,N_8433,N_7574);
and U9766 (N_9766,N_8244,N_8350);
or U9767 (N_9767,N_7953,N_8562);
and U9768 (N_9768,N_8815,N_7719);
or U9769 (N_9769,N_8431,N_7964);
nor U9770 (N_9770,N_8820,N_8585);
nand U9771 (N_9771,N_8657,N_8359);
nand U9772 (N_9772,N_8240,N_8439);
and U9773 (N_9773,N_7664,N_7820);
nor U9774 (N_9774,N_8881,N_8491);
nand U9775 (N_9775,N_8283,N_8377);
nor U9776 (N_9776,N_8562,N_8234);
xor U9777 (N_9777,N_8448,N_7663);
xnor U9778 (N_9778,N_7847,N_7742);
xor U9779 (N_9779,N_8227,N_8860);
xor U9780 (N_9780,N_8107,N_8544);
and U9781 (N_9781,N_8280,N_8540);
and U9782 (N_9782,N_8294,N_7682);
nor U9783 (N_9783,N_8995,N_7527);
nand U9784 (N_9784,N_8322,N_7716);
and U9785 (N_9785,N_8475,N_8563);
or U9786 (N_9786,N_8038,N_8767);
and U9787 (N_9787,N_8101,N_8692);
nor U9788 (N_9788,N_8378,N_7871);
xor U9789 (N_9789,N_8303,N_8861);
or U9790 (N_9790,N_8635,N_8231);
nand U9791 (N_9791,N_8898,N_8573);
or U9792 (N_9792,N_7884,N_7647);
and U9793 (N_9793,N_7830,N_8069);
nor U9794 (N_9794,N_7737,N_8738);
nor U9795 (N_9795,N_7559,N_7965);
nor U9796 (N_9796,N_7779,N_8368);
nor U9797 (N_9797,N_8084,N_8510);
or U9798 (N_9798,N_8032,N_8036);
nand U9799 (N_9799,N_8956,N_8879);
xor U9800 (N_9800,N_8582,N_7915);
nor U9801 (N_9801,N_8522,N_7579);
and U9802 (N_9802,N_8906,N_7897);
nor U9803 (N_9803,N_7767,N_8708);
nor U9804 (N_9804,N_8061,N_8945);
and U9805 (N_9805,N_8667,N_7597);
xnor U9806 (N_9806,N_8180,N_7760);
and U9807 (N_9807,N_7791,N_7857);
nand U9808 (N_9808,N_8929,N_7814);
or U9809 (N_9809,N_7629,N_8545);
and U9810 (N_9810,N_8192,N_7542);
or U9811 (N_9811,N_8124,N_8256);
and U9812 (N_9812,N_8607,N_7770);
and U9813 (N_9813,N_8325,N_8709);
or U9814 (N_9814,N_8838,N_7767);
or U9815 (N_9815,N_7781,N_8654);
nand U9816 (N_9816,N_8606,N_8214);
nor U9817 (N_9817,N_8731,N_7526);
nand U9818 (N_9818,N_8809,N_8992);
nand U9819 (N_9819,N_8984,N_7732);
xnor U9820 (N_9820,N_8410,N_7725);
nand U9821 (N_9821,N_8653,N_8638);
or U9822 (N_9822,N_8908,N_8467);
nor U9823 (N_9823,N_8531,N_8092);
and U9824 (N_9824,N_8545,N_7549);
or U9825 (N_9825,N_8477,N_8382);
xnor U9826 (N_9826,N_7629,N_7668);
xor U9827 (N_9827,N_8988,N_8956);
nor U9828 (N_9828,N_7599,N_7520);
nand U9829 (N_9829,N_8157,N_8136);
or U9830 (N_9830,N_8653,N_8136);
and U9831 (N_9831,N_7551,N_7734);
or U9832 (N_9832,N_7995,N_8352);
xnor U9833 (N_9833,N_8279,N_8101);
or U9834 (N_9834,N_8500,N_8389);
and U9835 (N_9835,N_7538,N_7862);
nor U9836 (N_9836,N_8785,N_7678);
or U9837 (N_9837,N_7623,N_7765);
nand U9838 (N_9838,N_8519,N_8438);
nand U9839 (N_9839,N_8787,N_7955);
and U9840 (N_9840,N_8457,N_8148);
nor U9841 (N_9841,N_7870,N_7859);
nor U9842 (N_9842,N_7612,N_8834);
xor U9843 (N_9843,N_8978,N_8048);
or U9844 (N_9844,N_8648,N_7766);
xnor U9845 (N_9845,N_8400,N_8734);
and U9846 (N_9846,N_7635,N_8188);
nand U9847 (N_9847,N_7872,N_7982);
nor U9848 (N_9848,N_8646,N_7675);
nor U9849 (N_9849,N_8774,N_8051);
nand U9850 (N_9850,N_8326,N_8399);
nand U9851 (N_9851,N_7898,N_8639);
or U9852 (N_9852,N_8889,N_7910);
xnor U9853 (N_9853,N_8587,N_7688);
nand U9854 (N_9854,N_8093,N_7552);
and U9855 (N_9855,N_8381,N_8322);
and U9856 (N_9856,N_8031,N_8956);
nand U9857 (N_9857,N_8570,N_8292);
xnor U9858 (N_9858,N_8510,N_7501);
nor U9859 (N_9859,N_7627,N_8348);
or U9860 (N_9860,N_8009,N_7968);
nand U9861 (N_9861,N_8446,N_8487);
nor U9862 (N_9862,N_8338,N_8618);
xor U9863 (N_9863,N_7767,N_7864);
nand U9864 (N_9864,N_8934,N_8719);
xor U9865 (N_9865,N_8501,N_7890);
nand U9866 (N_9866,N_8566,N_8512);
or U9867 (N_9867,N_8179,N_8191);
and U9868 (N_9868,N_8860,N_8976);
and U9869 (N_9869,N_8542,N_7990);
nor U9870 (N_9870,N_8828,N_8189);
xnor U9871 (N_9871,N_8840,N_7658);
and U9872 (N_9872,N_7894,N_8815);
nor U9873 (N_9873,N_8574,N_7783);
nand U9874 (N_9874,N_8529,N_8700);
and U9875 (N_9875,N_8728,N_8950);
xnor U9876 (N_9876,N_8681,N_8717);
nand U9877 (N_9877,N_8437,N_7704);
nand U9878 (N_9878,N_8500,N_8643);
and U9879 (N_9879,N_8938,N_8415);
nor U9880 (N_9880,N_8548,N_7684);
xor U9881 (N_9881,N_8892,N_8371);
nand U9882 (N_9882,N_8317,N_8678);
nand U9883 (N_9883,N_8525,N_7594);
nand U9884 (N_9884,N_7560,N_7525);
xnor U9885 (N_9885,N_7537,N_8369);
nor U9886 (N_9886,N_8342,N_8274);
xnor U9887 (N_9887,N_8966,N_8322);
nor U9888 (N_9888,N_8070,N_8945);
xor U9889 (N_9889,N_8092,N_8320);
or U9890 (N_9890,N_8629,N_8873);
and U9891 (N_9891,N_8799,N_7649);
xnor U9892 (N_9892,N_8981,N_7858);
and U9893 (N_9893,N_7818,N_7937);
and U9894 (N_9894,N_7639,N_7931);
and U9895 (N_9895,N_7902,N_7808);
xor U9896 (N_9896,N_7685,N_8806);
or U9897 (N_9897,N_8857,N_7691);
or U9898 (N_9898,N_7580,N_7627);
nand U9899 (N_9899,N_8736,N_8279);
xnor U9900 (N_9900,N_8676,N_8421);
nor U9901 (N_9901,N_7894,N_7512);
and U9902 (N_9902,N_8570,N_7897);
and U9903 (N_9903,N_8684,N_7550);
and U9904 (N_9904,N_8655,N_8264);
nand U9905 (N_9905,N_7982,N_8138);
xnor U9906 (N_9906,N_8513,N_8552);
and U9907 (N_9907,N_8915,N_8182);
and U9908 (N_9908,N_8440,N_8881);
nor U9909 (N_9909,N_8719,N_8233);
or U9910 (N_9910,N_8361,N_8009);
nand U9911 (N_9911,N_8807,N_8179);
nor U9912 (N_9912,N_7563,N_8810);
nand U9913 (N_9913,N_8232,N_8771);
nor U9914 (N_9914,N_8087,N_7971);
xor U9915 (N_9915,N_8767,N_8285);
xor U9916 (N_9916,N_7772,N_7712);
and U9917 (N_9917,N_7509,N_8171);
or U9918 (N_9918,N_8303,N_8524);
nor U9919 (N_9919,N_8911,N_8421);
xor U9920 (N_9920,N_8842,N_7526);
nand U9921 (N_9921,N_7946,N_8824);
nor U9922 (N_9922,N_8468,N_7995);
or U9923 (N_9923,N_8687,N_8978);
xor U9924 (N_9924,N_8998,N_8663);
nor U9925 (N_9925,N_8433,N_7904);
and U9926 (N_9926,N_8445,N_7703);
and U9927 (N_9927,N_8442,N_8071);
nand U9928 (N_9928,N_8254,N_8675);
xor U9929 (N_9929,N_8383,N_8937);
or U9930 (N_9930,N_7644,N_8671);
nand U9931 (N_9931,N_8845,N_8475);
and U9932 (N_9932,N_8637,N_8215);
nand U9933 (N_9933,N_8323,N_8699);
or U9934 (N_9934,N_8968,N_8489);
or U9935 (N_9935,N_8814,N_8216);
xnor U9936 (N_9936,N_7844,N_8857);
and U9937 (N_9937,N_8489,N_7618);
nand U9938 (N_9938,N_8131,N_7716);
xor U9939 (N_9939,N_7937,N_7677);
nor U9940 (N_9940,N_7770,N_8896);
or U9941 (N_9941,N_8008,N_8514);
nand U9942 (N_9942,N_7686,N_8954);
and U9943 (N_9943,N_7734,N_8348);
or U9944 (N_9944,N_8344,N_8097);
nand U9945 (N_9945,N_8149,N_7906);
and U9946 (N_9946,N_8686,N_7601);
xor U9947 (N_9947,N_7661,N_8899);
nor U9948 (N_9948,N_7821,N_8024);
nor U9949 (N_9949,N_8021,N_7689);
and U9950 (N_9950,N_7961,N_8856);
or U9951 (N_9951,N_8942,N_7990);
nor U9952 (N_9952,N_8124,N_8005);
or U9953 (N_9953,N_8329,N_8222);
nor U9954 (N_9954,N_8205,N_8695);
and U9955 (N_9955,N_7643,N_8572);
nand U9956 (N_9956,N_7992,N_7842);
or U9957 (N_9957,N_7719,N_7688);
nand U9958 (N_9958,N_7650,N_8931);
and U9959 (N_9959,N_8847,N_8333);
and U9960 (N_9960,N_8380,N_8428);
xnor U9961 (N_9961,N_7651,N_8474);
nand U9962 (N_9962,N_8714,N_7683);
or U9963 (N_9963,N_8382,N_8272);
nand U9964 (N_9964,N_8598,N_8646);
and U9965 (N_9965,N_7659,N_8024);
nand U9966 (N_9966,N_7749,N_7588);
or U9967 (N_9967,N_7949,N_8714);
and U9968 (N_9968,N_8631,N_7926);
or U9969 (N_9969,N_8194,N_8865);
nand U9970 (N_9970,N_8441,N_7930);
or U9971 (N_9971,N_8425,N_8297);
nand U9972 (N_9972,N_8390,N_8287);
nand U9973 (N_9973,N_8900,N_8478);
xnor U9974 (N_9974,N_8414,N_8829);
xnor U9975 (N_9975,N_7759,N_8336);
or U9976 (N_9976,N_8164,N_7902);
nor U9977 (N_9977,N_8316,N_8454);
and U9978 (N_9978,N_8823,N_8406);
and U9979 (N_9979,N_8060,N_8203);
nor U9980 (N_9980,N_8805,N_8729);
xor U9981 (N_9981,N_8072,N_7614);
nand U9982 (N_9982,N_7888,N_8029);
xor U9983 (N_9983,N_8120,N_7714);
and U9984 (N_9984,N_7982,N_8094);
xor U9985 (N_9985,N_8278,N_8296);
or U9986 (N_9986,N_8834,N_8065);
xor U9987 (N_9987,N_8472,N_7857);
nand U9988 (N_9988,N_8232,N_8775);
nor U9989 (N_9989,N_8583,N_8210);
nand U9990 (N_9990,N_8593,N_8001);
xor U9991 (N_9991,N_7950,N_8585);
and U9992 (N_9992,N_8753,N_8102);
xor U9993 (N_9993,N_8716,N_8670);
xnor U9994 (N_9994,N_8085,N_8701);
and U9995 (N_9995,N_8687,N_7582);
and U9996 (N_9996,N_8399,N_8200);
nand U9997 (N_9997,N_8705,N_8149);
nor U9998 (N_9998,N_8903,N_8121);
and U9999 (N_9999,N_8259,N_8717);
nand U10000 (N_10000,N_8763,N_8148);
or U10001 (N_10001,N_7595,N_8491);
xor U10002 (N_10002,N_8804,N_8520);
xor U10003 (N_10003,N_8686,N_8837);
or U10004 (N_10004,N_7568,N_8149);
nor U10005 (N_10005,N_7891,N_7841);
nand U10006 (N_10006,N_7683,N_7644);
nand U10007 (N_10007,N_8926,N_7917);
or U10008 (N_10008,N_8899,N_8842);
and U10009 (N_10009,N_7819,N_7992);
and U10010 (N_10010,N_8514,N_8552);
and U10011 (N_10011,N_7839,N_8384);
xnor U10012 (N_10012,N_8147,N_8740);
nor U10013 (N_10013,N_8625,N_7894);
and U10014 (N_10014,N_7689,N_7963);
nand U10015 (N_10015,N_8112,N_7748);
nand U10016 (N_10016,N_8885,N_7686);
xnor U10017 (N_10017,N_7554,N_8269);
or U10018 (N_10018,N_7653,N_8214);
xor U10019 (N_10019,N_8790,N_7882);
or U10020 (N_10020,N_8492,N_7869);
and U10021 (N_10021,N_8150,N_8989);
xnor U10022 (N_10022,N_7746,N_7761);
and U10023 (N_10023,N_8104,N_8467);
and U10024 (N_10024,N_7868,N_8469);
xor U10025 (N_10025,N_8646,N_8870);
nor U10026 (N_10026,N_8008,N_7739);
nor U10027 (N_10027,N_7741,N_8238);
or U10028 (N_10028,N_8538,N_8104);
xnor U10029 (N_10029,N_8955,N_7765);
xnor U10030 (N_10030,N_8312,N_8358);
nor U10031 (N_10031,N_8338,N_8532);
xnor U10032 (N_10032,N_8755,N_8957);
nor U10033 (N_10033,N_8563,N_8874);
nand U10034 (N_10034,N_8225,N_8479);
xnor U10035 (N_10035,N_8527,N_7831);
xor U10036 (N_10036,N_7713,N_8485);
nor U10037 (N_10037,N_7937,N_8932);
nor U10038 (N_10038,N_7595,N_7757);
xnor U10039 (N_10039,N_7592,N_8529);
and U10040 (N_10040,N_7757,N_8610);
and U10041 (N_10041,N_8511,N_8845);
nor U10042 (N_10042,N_7769,N_7653);
and U10043 (N_10043,N_7883,N_7996);
nor U10044 (N_10044,N_7867,N_8348);
nor U10045 (N_10045,N_8482,N_8712);
xnor U10046 (N_10046,N_7931,N_8540);
or U10047 (N_10047,N_8748,N_7735);
xor U10048 (N_10048,N_8324,N_7525);
and U10049 (N_10049,N_8222,N_7766);
nor U10050 (N_10050,N_8020,N_8769);
or U10051 (N_10051,N_8384,N_7540);
xnor U10052 (N_10052,N_7679,N_8566);
nor U10053 (N_10053,N_8938,N_8808);
nor U10054 (N_10054,N_8685,N_8362);
nor U10055 (N_10055,N_8715,N_8533);
nor U10056 (N_10056,N_8804,N_7811);
nor U10057 (N_10057,N_8710,N_8293);
or U10058 (N_10058,N_7671,N_8376);
xnor U10059 (N_10059,N_8231,N_8090);
or U10060 (N_10060,N_8077,N_7608);
xnor U10061 (N_10061,N_7698,N_8611);
or U10062 (N_10062,N_8038,N_7553);
and U10063 (N_10063,N_7968,N_8846);
and U10064 (N_10064,N_7721,N_8988);
and U10065 (N_10065,N_7874,N_8797);
nor U10066 (N_10066,N_7798,N_8687);
nand U10067 (N_10067,N_8812,N_8706);
or U10068 (N_10068,N_8488,N_7864);
nor U10069 (N_10069,N_7752,N_8657);
nand U10070 (N_10070,N_8586,N_7673);
or U10071 (N_10071,N_8523,N_7599);
and U10072 (N_10072,N_7544,N_8779);
nor U10073 (N_10073,N_8407,N_7857);
nand U10074 (N_10074,N_7914,N_7969);
or U10075 (N_10075,N_8978,N_8240);
and U10076 (N_10076,N_7506,N_7523);
xnor U10077 (N_10077,N_8666,N_7903);
nand U10078 (N_10078,N_8034,N_8277);
xnor U10079 (N_10079,N_8687,N_8635);
or U10080 (N_10080,N_7735,N_8891);
xnor U10081 (N_10081,N_8231,N_8734);
and U10082 (N_10082,N_8989,N_7549);
nand U10083 (N_10083,N_8586,N_8867);
nand U10084 (N_10084,N_8932,N_8698);
and U10085 (N_10085,N_8209,N_8517);
xor U10086 (N_10086,N_8052,N_7550);
xor U10087 (N_10087,N_7876,N_8160);
nand U10088 (N_10088,N_8512,N_7995);
or U10089 (N_10089,N_8238,N_8680);
and U10090 (N_10090,N_7957,N_8291);
xor U10091 (N_10091,N_7863,N_8820);
and U10092 (N_10092,N_7588,N_8754);
nand U10093 (N_10093,N_8137,N_7887);
or U10094 (N_10094,N_8439,N_7706);
or U10095 (N_10095,N_8256,N_8481);
and U10096 (N_10096,N_7766,N_7795);
xor U10097 (N_10097,N_8811,N_8910);
nor U10098 (N_10098,N_7847,N_8883);
or U10099 (N_10099,N_7696,N_7805);
or U10100 (N_10100,N_8703,N_7557);
nand U10101 (N_10101,N_7966,N_7669);
nand U10102 (N_10102,N_7552,N_7500);
xnor U10103 (N_10103,N_8127,N_7931);
and U10104 (N_10104,N_7952,N_8003);
and U10105 (N_10105,N_8959,N_8123);
or U10106 (N_10106,N_8964,N_8306);
xnor U10107 (N_10107,N_8989,N_8568);
nand U10108 (N_10108,N_8110,N_7818);
or U10109 (N_10109,N_8080,N_7617);
nor U10110 (N_10110,N_8789,N_7827);
or U10111 (N_10111,N_8809,N_8124);
xnor U10112 (N_10112,N_8225,N_7612);
and U10113 (N_10113,N_8272,N_8229);
xnor U10114 (N_10114,N_7649,N_7537);
nor U10115 (N_10115,N_8454,N_8347);
or U10116 (N_10116,N_8366,N_8409);
or U10117 (N_10117,N_8105,N_8898);
or U10118 (N_10118,N_7862,N_7848);
nor U10119 (N_10119,N_7929,N_8200);
nand U10120 (N_10120,N_8562,N_8890);
and U10121 (N_10121,N_8081,N_7885);
xor U10122 (N_10122,N_8251,N_7892);
nand U10123 (N_10123,N_7714,N_8504);
nand U10124 (N_10124,N_8770,N_8717);
and U10125 (N_10125,N_8103,N_8285);
nor U10126 (N_10126,N_8146,N_8450);
and U10127 (N_10127,N_8447,N_7804);
or U10128 (N_10128,N_7726,N_7603);
and U10129 (N_10129,N_8727,N_7985);
nor U10130 (N_10130,N_7739,N_8499);
nand U10131 (N_10131,N_8141,N_8617);
nand U10132 (N_10132,N_7934,N_7513);
nand U10133 (N_10133,N_8150,N_8165);
or U10134 (N_10134,N_8822,N_7969);
nor U10135 (N_10135,N_7633,N_8830);
xnor U10136 (N_10136,N_7743,N_8307);
xnor U10137 (N_10137,N_8660,N_8712);
nand U10138 (N_10138,N_7855,N_8317);
nand U10139 (N_10139,N_8108,N_8443);
xnor U10140 (N_10140,N_7578,N_8638);
and U10141 (N_10141,N_8345,N_8271);
nand U10142 (N_10142,N_8623,N_7725);
nor U10143 (N_10143,N_8641,N_7710);
xnor U10144 (N_10144,N_8595,N_8711);
xor U10145 (N_10145,N_8096,N_8959);
or U10146 (N_10146,N_7833,N_8826);
nand U10147 (N_10147,N_8648,N_8958);
nand U10148 (N_10148,N_7577,N_8619);
nor U10149 (N_10149,N_7981,N_7696);
nor U10150 (N_10150,N_8224,N_8639);
xnor U10151 (N_10151,N_8789,N_8417);
or U10152 (N_10152,N_8548,N_8123);
nand U10153 (N_10153,N_8398,N_8621);
or U10154 (N_10154,N_8559,N_8874);
nor U10155 (N_10155,N_8934,N_8034);
and U10156 (N_10156,N_8658,N_8085);
xnor U10157 (N_10157,N_8592,N_8690);
or U10158 (N_10158,N_8984,N_8543);
and U10159 (N_10159,N_8869,N_8362);
or U10160 (N_10160,N_8669,N_8679);
xnor U10161 (N_10161,N_8149,N_8355);
or U10162 (N_10162,N_7635,N_8300);
nand U10163 (N_10163,N_8811,N_8820);
nand U10164 (N_10164,N_7857,N_8894);
or U10165 (N_10165,N_8476,N_8488);
xnor U10166 (N_10166,N_8234,N_8014);
or U10167 (N_10167,N_7762,N_8624);
nand U10168 (N_10168,N_7984,N_7610);
xnor U10169 (N_10169,N_8035,N_8118);
nand U10170 (N_10170,N_8879,N_7983);
or U10171 (N_10171,N_7630,N_7828);
nor U10172 (N_10172,N_8721,N_8019);
or U10173 (N_10173,N_7801,N_8981);
nand U10174 (N_10174,N_7981,N_7942);
nand U10175 (N_10175,N_7852,N_8322);
and U10176 (N_10176,N_7852,N_8024);
xor U10177 (N_10177,N_7792,N_8663);
or U10178 (N_10178,N_8566,N_8889);
and U10179 (N_10179,N_8767,N_7532);
xor U10180 (N_10180,N_8946,N_8379);
or U10181 (N_10181,N_7615,N_7810);
nand U10182 (N_10182,N_7858,N_7744);
or U10183 (N_10183,N_8886,N_8698);
nor U10184 (N_10184,N_7686,N_7671);
or U10185 (N_10185,N_8831,N_8903);
nand U10186 (N_10186,N_8844,N_8332);
xnor U10187 (N_10187,N_8604,N_8377);
nor U10188 (N_10188,N_7737,N_7592);
xor U10189 (N_10189,N_8646,N_8833);
nor U10190 (N_10190,N_7885,N_8286);
or U10191 (N_10191,N_8385,N_8166);
and U10192 (N_10192,N_8951,N_8275);
or U10193 (N_10193,N_8257,N_8647);
and U10194 (N_10194,N_8915,N_8071);
or U10195 (N_10195,N_7616,N_7975);
nand U10196 (N_10196,N_8226,N_7765);
nand U10197 (N_10197,N_8197,N_8413);
and U10198 (N_10198,N_8029,N_8379);
nor U10199 (N_10199,N_7912,N_7867);
nor U10200 (N_10200,N_7912,N_8029);
and U10201 (N_10201,N_7546,N_8954);
xnor U10202 (N_10202,N_7565,N_8935);
and U10203 (N_10203,N_8840,N_7562);
and U10204 (N_10204,N_8249,N_8323);
and U10205 (N_10205,N_8592,N_7792);
and U10206 (N_10206,N_8488,N_7750);
xor U10207 (N_10207,N_8043,N_8024);
xor U10208 (N_10208,N_8210,N_8467);
nor U10209 (N_10209,N_8312,N_8721);
nor U10210 (N_10210,N_8403,N_8434);
or U10211 (N_10211,N_8377,N_8590);
and U10212 (N_10212,N_7937,N_7679);
xor U10213 (N_10213,N_8158,N_7607);
xnor U10214 (N_10214,N_8725,N_8745);
nor U10215 (N_10215,N_7653,N_7596);
xnor U10216 (N_10216,N_8191,N_8182);
and U10217 (N_10217,N_8724,N_8175);
and U10218 (N_10218,N_8942,N_8021);
xnor U10219 (N_10219,N_7557,N_7546);
and U10220 (N_10220,N_8870,N_8733);
nand U10221 (N_10221,N_7784,N_7788);
and U10222 (N_10222,N_8121,N_7856);
nor U10223 (N_10223,N_7764,N_8947);
and U10224 (N_10224,N_7876,N_8962);
nor U10225 (N_10225,N_8157,N_7799);
nor U10226 (N_10226,N_7857,N_8956);
or U10227 (N_10227,N_7715,N_8955);
and U10228 (N_10228,N_8204,N_7554);
and U10229 (N_10229,N_8474,N_8424);
nor U10230 (N_10230,N_7926,N_7639);
xor U10231 (N_10231,N_7986,N_8886);
xnor U10232 (N_10232,N_7894,N_8887);
nand U10233 (N_10233,N_8862,N_8606);
and U10234 (N_10234,N_8840,N_7851);
xor U10235 (N_10235,N_8852,N_7924);
xor U10236 (N_10236,N_8505,N_8605);
or U10237 (N_10237,N_7862,N_8331);
or U10238 (N_10238,N_7882,N_8985);
nor U10239 (N_10239,N_8741,N_7532);
nor U10240 (N_10240,N_7725,N_8614);
nor U10241 (N_10241,N_7917,N_8074);
or U10242 (N_10242,N_7598,N_7970);
nand U10243 (N_10243,N_7790,N_7689);
and U10244 (N_10244,N_8077,N_8936);
nor U10245 (N_10245,N_8303,N_8152);
nor U10246 (N_10246,N_7794,N_7927);
xnor U10247 (N_10247,N_7727,N_7568);
nand U10248 (N_10248,N_8271,N_8257);
xnor U10249 (N_10249,N_8330,N_7996);
xor U10250 (N_10250,N_8628,N_8517);
or U10251 (N_10251,N_8246,N_8965);
and U10252 (N_10252,N_8947,N_7642);
and U10253 (N_10253,N_7865,N_8724);
nor U10254 (N_10254,N_8671,N_7823);
nor U10255 (N_10255,N_8415,N_8263);
nand U10256 (N_10256,N_8410,N_8028);
nor U10257 (N_10257,N_8977,N_8206);
or U10258 (N_10258,N_8629,N_8135);
and U10259 (N_10259,N_7537,N_7945);
and U10260 (N_10260,N_7775,N_8008);
nor U10261 (N_10261,N_8561,N_7657);
or U10262 (N_10262,N_7828,N_8451);
or U10263 (N_10263,N_7964,N_8138);
and U10264 (N_10264,N_8778,N_8281);
and U10265 (N_10265,N_8567,N_8118);
or U10266 (N_10266,N_8675,N_8371);
nand U10267 (N_10267,N_8633,N_8203);
or U10268 (N_10268,N_7961,N_8139);
and U10269 (N_10269,N_8155,N_8184);
xnor U10270 (N_10270,N_8771,N_8550);
or U10271 (N_10271,N_8744,N_8326);
xnor U10272 (N_10272,N_8998,N_8772);
and U10273 (N_10273,N_8168,N_7766);
xnor U10274 (N_10274,N_7601,N_8637);
and U10275 (N_10275,N_8677,N_8243);
nor U10276 (N_10276,N_8776,N_8430);
nor U10277 (N_10277,N_8114,N_7650);
nor U10278 (N_10278,N_8173,N_7785);
and U10279 (N_10279,N_8059,N_8574);
and U10280 (N_10280,N_8167,N_8284);
and U10281 (N_10281,N_8471,N_8350);
and U10282 (N_10282,N_7521,N_7930);
xnor U10283 (N_10283,N_8595,N_8429);
nand U10284 (N_10284,N_8538,N_8400);
and U10285 (N_10285,N_8144,N_8412);
and U10286 (N_10286,N_7730,N_8419);
xor U10287 (N_10287,N_8202,N_7881);
xor U10288 (N_10288,N_8392,N_8889);
or U10289 (N_10289,N_8962,N_8525);
xor U10290 (N_10290,N_8531,N_8691);
or U10291 (N_10291,N_7534,N_8616);
xor U10292 (N_10292,N_8833,N_8482);
nor U10293 (N_10293,N_8178,N_8473);
nor U10294 (N_10294,N_7953,N_8620);
nor U10295 (N_10295,N_8599,N_8582);
and U10296 (N_10296,N_8235,N_8685);
and U10297 (N_10297,N_8361,N_7672);
and U10298 (N_10298,N_7807,N_7522);
and U10299 (N_10299,N_7771,N_7890);
and U10300 (N_10300,N_8455,N_8001);
nand U10301 (N_10301,N_8028,N_8076);
or U10302 (N_10302,N_8454,N_8562);
xor U10303 (N_10303,N_8989,N_8580);
xnor U10304 (N_10304,N_8000,N_7650);
or U10305 (N_10305,N_8110,N_8071);
and U10306 (N_10306,N_8738,N_7523);
xor U10307 (N_10307,N_8737,N_8426);
or U10308 (N_10308,N_7778,N_8251);
xnor U10309 (N_10309,N_8249,N_7673);
xnor U10310 (N_10310,N_8283,N_7632);
or U10311 (N_10311,N_7887,N_7613);
xor U10312 (N_10312,N_7502,N_8838);
or U10313 (N_10313,N_8318,N_8931);
nand U10314 (N_10314,N_8696,N_7790);
nor U10315 (N_10315,N_7876,N_8061);
nand U10316 (N_10316,N_8168,N_8258);
nor U10317 (N_10317,N_7785,N_7886);
nor U10318 (N_10318,N_8432,N_7510);
or U10319 (N_10319,N_7928,N_8036);
nor U10320 (N_10320,N_7685,N_8051);
nor U10321 (N_10321,N_8997,N_8963);
xor U10322 (N_10322,N_7834,N_8637);
and U10323 (N_10323,N_8508,N_8428);
and U10324 (N_10324,N_8670,N_8198);
or U10325 (N_10325,N_7798,N_8411);
or U10326 (N_10326,N_8709,N_8792);
nand U10327 (N_10327,N_7759,N_7702);
nor U10328 (N_10328,N_8517,N_7751);
xnor U10329 (N_10329,N_8165,N_8866);
xor U10330 (N_10330,N_8428,N_7879);
and U10331 (N_10331,N_8872,N_7879);
nand U10332 (N_10332,N_7844,N_8451);
nor U10333 (N_10333,N_7538,N_7615);
nor U10334 (N_10334,N_7950,N_7652);
or U10335 (N_10335,N_7585,N_8691);
nor U10336 (N_10336,N_7785,N_8225);
nand U10337 (N_10337,N_7702,N_7659);
or U10338 (N_10338,N_8841,N_8615);
or U10339 (N_10339,N_7758,N_7970);
nor U10340 (N_10340,N_7805,N_8112);
or U10341 (N_10341,N_8032,N_8069);
nor U10342 (N_10342,N_7871,N_7895);
nor U10343 (N_10343,N_7637,N_7770);
nor U10344 (N_10344,N_7721,N_8692);
xor U10345 (N_10345,N_8779,N_8675);
nand U10346 (N_10346,N_8453,N_8488);
nand U10347 (N_10347,N_8802,N_8075);
or U10348 (N_10348,N_8748,N_8499);
or U10349 (N_10349,N_7889,N_8398);
xnor U10350 (N_10350,N_8914,N_8996);
or U10351 (N_10351,N_7727,N_7856);
xor U10352 (N_10352,N_8967,N_7623);
and U10353 (N_10353,N_7934,N_7539);
nor U10354 (N_10354,N_7575,N_7562);
nand U10355 (N_10355,N_7904,N_8140);
nor U10356 (N_10356,N_8139,N_8045);
nand U10357 (N_10357,N_8190,N_7765);
or U10358 (N_10358,N_8112,N_8177);
and U10359 (N_10359,N_8816,N_8614);
and U10360 (N_10360,N_8040,N_8076);
nand U10361 (N_10361,N_7994,N_7938);
xor U10362 (N_10362,N_8483,N_8734);
xnor U10363 (N_10363,N_8075,N_8309);
nor U10364 (N_10364,N_7859,N_8943);
nand U10365 (N_10365,N_7718,N_7936);
xor U10366 (N_10366,N_8423,N_8773);
xor U10367 (N_10367,N_8332,N_8585);
nand U10368 (N_10368,N_8431,N_8090);
nor U10369 (N_10369,N_8014,N_8000);
and U10370 (N_10370,N_8742,N_7525);
xnor U10371 (N_10371,N_8237,N_7684);
and U10372 (N_10372,N_8784,N_8354);
nand U10373 (N_10373,N_7582,N_7835);
nor U10374 (N_10374,N_8941,N_8329);
nor U10375 (N_10375,N_7785,N_8894);
nand U10376 (N_10376,N_8317,N_8142);
xor U10377 (N_10377,N_8848,N_8240);
or U10378 (N_10378,N_8092,N_8755);
and U10379 (N_10379,N_7666,N_8945);
nand U10380 (N_10380,N_8837,N_7646);
and U10381 (N_10381,N_8243,N_8045);
or U10382 (N_10382,N_8371,N_8767);
and U10383 (N_10383,N_7563,N_7960);
and U10384 (N_10384,N_7957,N_8994);
nand U10385 (N_10385,N_8559,N_8870);
nor U10386 (N_10386,N_7854,N_8402);
or U10387 (N_10387,N_7925,N_8460);
nor U10388 (N_10388,N_7921,N_7522);
or U10389 (N_10389,N_8059,N_7617);
or U10390 (N_10390,N_7622,N_8463);
xor U10391 (N_10391,N_8398,N_7906);
and U10392 (N_10392,N_7670,N_8016);
nand U10393 (N_10393,N_8012,N_7867);
and U10394 (N_10394,N_7805,N_8134);
xor U10395 (N_10395,N_7854,N_8794);
and U10396 (N_10396,N_8558,N_8378);
nor U10397 (N_10397,N_7585,N_8911);
nor U10398 (N_10398,N_8134,N_8422);
nand U10399 (N_10399,N_8197,N_7610);
or U10400 (N_10400,N_8955,N_7962);
nor U10401 (N_10401,N_8037,N_8636);
or U10402 (N_10402,N_8993,N_7727);
or U10403 (N_10403,N_8183,N_8240);
nor U10404 (N_10404,N_8319,N_8189);
xnor U10405 (N_10405,N_8224,N_7533);
nor U10406 (N_10406,N_8383,N_7615);
xor U10407 (N_10407,N_7735,N_8468);
and U10408 (N_10408,N_8994,N_7644);
and U10409 (N_10409,N_8752,N_8442);
or U10410 (N_10410,N_7725,N_7807);
nor U10411 (N_10411,N_8264,N_7537);
xor U10412 (N_10412,N_8334,N_8871);
and U10413 (N_10413,N_7947,N_8152);
nor U10414 (N_10414,N_8213,N_8407);
nand U10415 (N_10415,N_8408,N_8697);
nor U10416 (N_10416,N_8270,N_8726);
nor U10417 (N_10417,N_8538,N_8825);
nor U10418 (N_10418,N_8097,N_8985);
nor U10419 (N_10419,N_8536,N_8025);
or U10420 (N_10420,N_8162,N_8942);
nor U10421 (N_10421,N_8496,N_8843);
and U10422 (N_10422,N_7998,N_7966);
and U10423 (N_10423,N_8966,N_8831);
xnor U10424 (N_10424,N_8450,N_7620);
and U10425 (N_10425,N_7626,N_8137);
nor U10426 (N_10426,N_8819,N_8210);
or U10427 (N_10427,N_8017,N_8129);
nor U10428 (N_10428,N_8714,N_8269);
and U10429 (N_10429,N_8115,N_7512);
and U10430 (N_10430,N_8959,N_7915);
nand U10431 (N_10431,N_8418,N_8692);
and U10432 (N_10432,N_8516,N_8170);
and U10433 (N_10433,N_8763,N_8907);
and U10434 (N_10434,N_8005,N_7760);
xor U10435 (N_10435,N_8303,N_7802);
xor U10436 (N_10436,N_7918,N_8003);
or U10437 (N_10437,N_8105,N_8646);
or U10438 (N_10438,N_8298,N_8240);
xor U10439 (N_10439,N_8538,N_7605);
xnor U10440 (N_10440,N_7701,N_8348);
and U10441 (N_10441,N_7963,N_7970);
and U10442 (N_10442,N_8361,N_7795);
nor U10443 (N_10443,N_8368,N_8446);
xor U10444 (N_10444,N_8964,N_7659);
nand U10445 (N_10445,N_7892,N_7786);
nand U10446 (N_10446,N_8657,N_8201);
or U10447 (N_10447,N_8284,N_8006);
nor U10448 (N_10448,N_8194,N_8073);
and U10449 (N_10449,N_7809,N_7525);
nor U10450 (N_10450,N_8833,N_8147);
nand U10451 (N_10451,N_8336,N_8833);
nor U10452 (N_10452,N_8619,N_7935);
and U10453 (N_10453,N_8521,N_8554);
or U10454 (N_10454,N_7958,N_8221);
nand U10455 (N_10455,N_8915,N_7915);
or U10456 (N_10456,N_8812,N_8209);
and U10457 (N_10457,N_7608,N_8782);
or U10458 (N_10458,N_8880,N_8054);
or U10459 (N_10459,N_8000,N_7516);
and U10460 (N_10460,N_8249,N_7741);
or U10461 (N_10461,N_8247,N_8135);
nand U10462 (N_10462,N_8686,N_8365);
and U10463 (N_10463,N_8256,N_7722);
nand U10464 (N_10464,N_8629,N_8572);
xor U10465 (N_10465,N_8871,N_8886);
xnor U10466 (N_10466,N_8500,N_8789);
and U10467 (N_10467,N_8121,N_7605);
and U10468 (N_10468,N_8015,N_8275);
and U10469 (N_10469,N_8408,N_8869);
or U10470 (N_10470,N_8656,N_8765);
xor U10471 (N_10471,N_7627,N_7768);
and U10472 (N_10472,N_8278,N_7671);
nor U10473 (N_10473,N_8272,N_8489);
nor U10474 (N_10474,N_8617,N_8466);
nor U10475 (N_10475,N_7667,N_7740);
nand U10476 (N_10476,N_8942,N_8478);
nand U10477 (N_10477,N_8227,N_8356);
xnor U10478 (N_10478,N_8428,N_8990);
xor U10479 (N_10479,N_8913,N_8169);
and U10480 (N_10480,N_7766,N_7978);
xnor U10481 (N_10481,N_7672,N_8918);
nor U10482 (N_10482,N_7643,N_7948);
xor U10483 (N_10483,N_8218,N_8701);
nor U10484 (N_10484,N_8040,N_7951);
and U10485 (N_10485,N_8108,N_8479);
nor U10486 (N_10486,N_8294,N_7812);
or U10487 (N_10487,N_7866,N_8077);
or U10488 (N_10488,N_8236,N_8188);
or U10489 (N_10489,N_8832,N_8421);
xor U10490 (N_10490,N_8478,N_8473);
or U10491 (N_10491,N_8645,N_8594);
nor U10492 (N_10492,N_8126,N_8117);
nor U10493 (N_10493,N_8161,N_8932);
nor U10494 (N_10494,N_8118,N_8675);
or U10495 (N_10495,N_8296,N_7637);
xor U10496 (N_10496,N_8448,N_7511);
or U10497 (N_10497,N_8135,N_8220);
nand U10498 (N_10498,N_7781,N_8487);
xnor U10499 (N_10499,N_8956,N_8146);
or U10500 (N_10500,N_9051,N_9575);
xnor U10501 (N_10501,N_10248,N_9700);
nor U10502 (N_10502,N_9909,N_9769);
nor U10503 (N_10503,N_9445,N_9174);
nor U10504 (N_10504,N_10387,N_9164);
and U10505 (N_10505,N_9163,N_10272);
or U10506 (N_10506,N_9841,N_9449);
and U10507 (N_10507,N_9736,N_10128);
nor U10508 (N_10508,N_10361,N_9530);
nand U10509 (N_10509,N_9443,N_9652);
or U10510 (N_10510,N_9246,N_9797);
or U10511 (N_10511,N_9107,N_9810);
nor U10512 (N_10512,N_9552,N_9074);
and U10513 (N_10513,N_10348,N_9819);
or U10514 (N_10514,N_9504,N_9434);
nand U10515 (N_10515,N_9308,N_10098);
nor U10516 (N_10516,N_10150,N_9430);
xnor U10517 (N_10517,N_9390,N_10154);
xor U10518 (N_10518,N_9265,N_9648);
and U10519 (N_10519,N_9191,N_9153);
nor U10520 (N_10520,N_10041,N_9774);
nand U10521 (N_10521,N_9050,N_9245);
or U10522 (N_10522,N_9803,N_9507);
or U10523 (N_10523,N_9101,N_10261);
and U10524 (N_10524,N_9440,N_9744);
xnor U10525 (N_10525,N_10290,N_9302);
nand U10526 (N_10526,N_9478,N_9137);
and U10527 (N_10527,N_9852,N_9953);
or U10528 (N_10528,N_9776,N_10453);
or U10529 (N_10529,N_9113,N_9637);
nand U10530 (N_10530,N_9655,N_10179);
or U10531 (N_10531,N_9379,N_10198);
nand U10532 (N_10532,N_10223,N_10412);
xor U10533 (N_10533,N_9503,N_9068);
xnor U10534 (N_10534,N_9377,N_9004);
xnor U10535 (N_10535,N_9871,N_10149);
or U10536 (N_10536,N_9709,N_10447);
xor U10537 (N_10537,N_9666,N_10492);
and U10538 (N_10538,N_9340,N_10095);
xnor U10539 (N_10539,N_10202,N_9018);
nor U10540 (N_10540,N_9956,N_10277);
or U10541 (N_10541,N_9509,N_10424);
nor U10542 (N_10542,N_9404,N_9121);
xnor U10543 (N_10543,N_9321,N_9179);
nor U10544 (N_10544,N_9830,N_9347);
xor U10545 (N_10545,N_9498,N_10350);
or U10546 (N_10546,N_10006,N_10423);
and U10547 (N_10547,N_9543,N_9537);
and U10548 (N_10548,N_9866,N_9924);
or U10549 (N_10549,N_9026,N_9234);
nor U10550 (N_10550,N_10431,N_9927);
nor U10551 (N_10551,N_9562,N_9737);
xor U10552 (N_10552,N_9664,N_9313);
or U10553 (N_10553,N_10273,N_9385);
xnor U10554 (N_10554,N_9998,N_9111);
or U10555 (N_10555,N_9186,N_9640);
xnor U10556 (N_10556,N_9786,N_9919);
or U10557 (N_10557,N_10384,N_9046);
and U10558 (N_10558,N_10059,N_9554);
xnor U10559 (N_10559,N_10125,N_9447);
xnor U10560 (N_10560,N_9991,N_9337);
nand U10561 (N_10561,N_9999,N_9886);
nand U10562 (N_10562,N_10123,N_10168);
and U10563 (N_10563,N_9820,N_10218);
or U10564 (N_10564,N_9785,N_9044);
and U10565 (N_10565,N_10260,N_9255);
or U10566 (N_10566,N_9954,N_9353);
nand U10567 (N_10567,N_9861,N_10340);
or U10568 (N_10568,N_9192,N_10274);
or U10569 (N_10569,N_9077,N_10490);
xnor U10570 (N_10570,N_9043,N_10382);
nor U10571 (N_10571,N_10334,N_9407);
and U10572 (N_10572,N_10430,N_9903);
nand U10573 (N_10573,N_9361,N_10081);
xor U10574 (N_10574,N_9633,N_9715);
nor U10575 (N_10575,N_9789,N_9423);
xnor U10576 (N_10576,N_9060,N_9942);
nand U10577 (N_10577,N_9100,N_9446);
and U10578 (N_10578,N_10079,N_10498);
or U10579 (N_10579,N_9396,N_9695);
nor U10580 (N_10580,N_10239,N_9398);
or U10581 (N_10581,N_9968,N_10421);
nand U10582 (N_10582,N_9030,N_9740);
xnor U10583 (N_10583,N_9222,N_10313);
and U10584 (N_10584,N_10271,N_10156);
nor U10585 (N_10585,N_10300,N_9099);
and U10586 (N_10586,N_9105,N_9873);
nand U10587 (N_10587,N_9611,N_9657);
and U10588 (N_10588,N_10344,N_9704);
and U10589 (N_10589,N_9817,N_9489);
xnor U10590 (N_10590,N_9822,N_9807);
xor U10591 (N_10591,N_9758,N_10297);
xnor U10592 (N_10592,N_10325,N_10388);
or U10593 (N_10593,N_10103,N_10312);
xor U10594 (N_10594,N_9135,N_9836);
xnor U10595 (N_10595,N_9808,N_9545);
and U10596 (N_10596,N_9225,N_9485);
or U10597 (N_10597,N_10220,N_10178);
nor U10598 (N_10598,N_9252,N_10242);
nand U10599 (N_10599,N_10365,N_9124);
nor U10600 (N_10600,N_9865,N_9452);
or U10601 (N_10601,N_9471,N_9600);
and U10602 (N_10602,N_9804,N_9754);
nor U10603 (N_10603,N_9818,N_9196);
nor U10604 (N_10604,N_9607,N_9437);
nor U10605 (N_10605,N_10358,N_9875);
xnor U10606 (N_10606,N_10296,N_10426);
xor U10607 (N_10607,N_10152,N_9676);
nor U10608 (N_10608,N_10204,N_9921);
nand U10609 (N_10609,N_10285,N_9370);
nand U10610 (N_10610,N_10039,N_9933);
or U10611 (N_10611,N_10134,N_10457);
xor U10612 (N_10612,N_10011,N_9006);
xnor U10613 (N_10613,N_9948,N_9592);
nor U10614 (N_10614,N_9049,N_9949);
nor U10615 (N_10615,N_9232,N_10449);
and U10616 (N_10616,N_10222,N_9891);
or U10617 (N_10617,N_9708,N_9734);
or U10618 (N_10618,N_10473,N_9605);
nor U10619 (N_10619,N_9168,N_10064);
and U10620 (N_10620,N_10063,N_9173);
or U10621 (N_10621,N_9380,N_9767);
nand U10622 (N_10622,N_9667,N_9867);
nand U10623 (N_10623,N_9297,N_9966);
or U10624 (N_10624,N_9585,N_9596);
nor U10625 (N_10625,N_10488,N_9765);
xnor U10626 (N_10626,N_9188,N_10166);
nand U10627 (N_10627,N_10108,N_10427);
nand U10628 (N_10628,N_10065,N_10475);
or U10629 (N_10629,N_10336,N_9905);
xor U10630 (N_10630,N_10302,N_9123);
or U10631 (N_10631,N_9923,N_10416);
or U10632 (N_10632,N_9036,N_10293);
xnor U10633 (N_10633,N_9488,N_9180);
xor U10634 (N_10634,N_9809,N_10180);
and U10635 (N_10635,N_9925,N_9939);
and U10636 (N_10636,N_9969,N_9209);
nor U10637 (N_10637,N_9112,N_10053);
or U10638 (N_10638,N_10048,N_9974);
nand U10639 (N_10639,N_9609,N_9242);
or U10640 (N_10640,N_10376,N_9499);
xor U10641 (N_10641,N_10107,N_9851);
nor U10642 (N_10642,N_9895,N_10253);
or U10643 (N_10643,N_10197,N_9182);
xor U10644 (N_10644,N_9813,N_10176);
and U10645 (N_10645,N_10240,N_10200);
nor U10646 (N_10646,N_9079,N_9687);
or U10647 (N_10647,N_9915,N_9210);
xor U10648 (N_10648,N_9730,N_10385);
and U10649 (N_10649,N_9799,N_10170);
and U10650 (N_10650,N_9673,N_9720);
nor U10651 (N_10651,N_9951,N_9500);
or U10652 (N_10652,N_10441,N_10339);
and U10653 (N_10653,N_9862,N_10395);
xnor U10654 (N_10654,N_9868,N_9037);
nor U10655 (N_10655,N_10030,N_9229);
or U10656 (N_10656,N_10052,N_9955);
nor U10657 (N_10657,N_9344,N_9181);
nor U10658 (N_10658,N_9978,N_9747);
nand U10659 (N_10659,N_9087,N_10330);
and U10660 (N_10660,N_9620,N_9271);
xnor U10661 (N_10661,N_9343,N_9680);
or U10662 (N_10662,N_9965,N_10034);
nor U10663 (N_10663,N_9461,N_9055);
or U10664 (N_10664,N_9384,N_9349);
xnor U10665 (N_10665,N_9269,N_9047);
nand U10666 (N_10666,N_9669,N_9928);
nor U10667 (N_10667,N_9106,N_9635);
xor U10668 (N_10668,N_9878,N_10035);
or U10669 (N_10669,N_9062,N_10148);
and U10670 (N_10670,N_10480,N_10213);
xnor U10671 (N_10671,N_9206,N_10363);
xnor U10672 (N_10672,N_10458,N_9763);
and U10673 (N_10673,N_9967,N_9301);
nor U10674 (N_10674,N_9063,N_9548);
xnor U10675 (N_10675,N_9364,N_10143);
nor U10676 (N_10676,N_9475,N_9490);
nor U10677 (N_10677,N_9457,N_9663);
xnor U10678 (N_10678,N_9355,N_10189);
xnor U10679 (N_10679,N_10489,N_9023);
or U10680 (N_10680,N_9299,N_10016);
and U10681 (N_10681,N_9712,N_9568);
nand U10682 (N_10682,N_10028,N_9165);
nand U10683 (N_10683,N_10493,N_10215);
or U10684 (N_10684,N_9595,N_9574);
and U10685 (N_10685,N_9354,N_9638);
nand U10686 (N_10686,N_10433,N_9703);
or U10687 (N_10687,N_9358,N_9617);
nor U10688 (N_10688,N_10280,N_10468);
or U10689 (N_10689,N_9336,N_9288);
nor U10690 (N_10690,N_9899,N_9801);
and U10691 (N_10691,N_10378,N_9439);
nand U10692 (N_10692,N_10194,N_10258);
nor U10693 (N_10693,N_10338,N_10046);
nand U10694 (N_10694,N_9567,N_9015);
xor U10695 (N_10695,N_9646,N_9685);
nor U10696 (N_10696,N_9913,N_9551);
xor U10697 (N_10697,N_9535,N_9368);
or U10698 (N_10698,N_10229,N_10354);
or U10699 (N_10699,N_9144,N_9997);
nor U10700 (N_10700,N_9127,N_9166);
and U10701 (N_10701,N_10131,N_9076);
xor U10702 (N_10702,N_9802,N_9952);
xnor U10703 (N_10703,N_9413,N_9155);
nand U10704 (N_10704,N_10368,N_10130);
and U10705 (N_10705,N_9083,N_9096);
nor U10706 (N_10706,N_9834,N_9395);
and U10707 (N_10707,N_9946,N_9244);
xnor U10708 (N_10708,N_9837,N_9701);
nor U10709 (N_10709,N_9001,N_9022);
and U10710 (N_10710,N_10422,N_10076);
and U10711 (N_10711,N_9787,N_9415);
or U10712 (N_10712,N_9938,N_10235);
xnor U10713 (N_10713,N_10404,N_9492);
nand U10714 (N_10714,N_9738,N_10055);
nand U10715 (N_10715,N_10083,N_10446);
nor U10716 (N_10716,N_10209,N_10124);
and U10717 (N_10717,N_9081,N_9156);
xor U10718 (N_10718,N_10397,N_10392);
nand U10719 (N_10719,N_9352,N_10097);
or U10720 (N_10720,N_9133,N_9702);
nand U10721 (N_10721,N_10310,N_10283);
or U10722 (N_10722,N_9872,N_10331);
xnor U10723 (N_10723,N_9178,N_9326);
nand U10724 (N_10724,N_9989,N_9311);
xnor U10725 (N_10725,N_9777,N_9278);
nand U10726 (N_10726,N_10038,N_10352);
xnor U10727 (N_10727,N_10225,N_9713);
or U10728 (N_10728,N_9661,N_10276);
or U10729 (N_10729,N_10318,N_9464);
and U10730 (N_10730,N_9070,N_9456);
and U10731 (N_10731,N_9973,N_9421);
and U10732 (N_10732,N_10356,N_9745);
and U10733 (N_10733,N_9935,N_10205);
and U10734 (N_10734,N_9943,N_10085);
nand U10735 (N_10735,N_10221,N_10173);
xor U10736 (N_10736,N_9118,N_9177);
nand U10737 (N_10737,N_9645,N_9389);
or U10738 (N_10738,N_9084,N_9618);
xor U10739 (N_10739,N_9858,N_9816);
xor U10740 (N_10740,N_9002,N_10461);
xor U10741 (N_10741,N_9435,N_9020);
xnor U10742 (N_10742,N_10266,N_10469);
nand U10743 (N_10743,N_9850,N_10369);
nor U10744 (N_10744,N_9573,N_9760);
or U10745 (N_10745,N_9205,N_9912);
or U10746 (N_10746,N_9406,N_9069);
nor U10747 (N_10747,N_9835,N_10137);
xor U10748 (N_10748,N_9040,N_9262);
xnor U10749 (N_10749,N_9114,N_9298);
xnor U10750 (N_10750,N_9920,N_9305);
nor U10751 (N_10751,N_9134,N_9937);
xor U10752 (N_10752,N_9863,N_10144);
and U10753 (N_10753,N_9204,N_10443);
nand U10754 (N_10754,N_10036,N_10005);
nand U10755 (N_10755,N_9587,N_9828);
or U10756 (N_10756,N_9468,N_9932);
and U10757 (N_10757,N_9211,N_9272);
xor U10758 (N_10758,N_10249,N_10316);
nor U10759 (N_10759,N_10074,N_9699);
nor U10760 (N_10760,N_10259,N_9710);
or U10761 (N_10761,N_9294,N_9593);
and U10762 (N_10762,N_9463,N_9625);
nand U10763 (N_10763,N_9682,N_10307);
and U10764 (N_10764,N_10136,N_9735);
nor U10765 (N_10765,N_9724,N_9557);
nand U10766 (N_10766,N_9523,N_9258);
nand U10767 (N_10767,N_9743,N_9926);
nand U10768 (N_10768,N_9986,N_10432);
and U10769 (N_10769,N_9675,N_9860);
xor U10770 (N_10770,N_10379,N_9003);
and U10771 (N_10771,N_9541,N_9529);
or U10772 (N_10772,N_10419,N_9911);
and U10773 (N_10773,N_9300,N_9581);
xor U10774 (N_10774,N_10265,N_9483);
nor U10775 (N_10775,N_10210,N_10304);
and U10776 (N_10776,N_10286,N_10017);
nor U10777 (N_10777,N_9442,N_10349);
nor U10778 (N_10778,N_10459,N_10429);
or U10779 (N_10779,N_9629,N_9260);
or U10780 (N_10780,N_9125,N_9280);
and U10781 (N_10781,N_9533,N_10037);
nor U10782 (N_10782,N_9591,N_10138);
nand U10783 (N_10783,N_9908,N_9285);
or U10784 (N_10784,N_9132,N_9613);
or U10785 (N_10785,N_9947,N_9658);
nand U10786 (N_10786,N_9782,N_10027);
nand U10787 (N_10787,N_9256,N_10428);
nor U10788 (N_10788,N_9750,N_9520);
xor U10789 (N_10789,N_9580,N_9189);
nor U10790 (N_10790,N_9433,N_9399);
xnor U10791 (N_10791,N_9846,N_9513);
nand U10792 (N_10792,N_10303,N_9459);
nor U10793 (N_10793,N_9462,N_9171);
nor U10794 (N_10794,N_9091,N_9547);
or U10795 (N_10795,N_10263,N_9831);
or U10796 (N_10796,N_9167,N_10184);
and U10797 (N_10797,N_9486,N_10279);
or U10798 (N_10798,N_9103,N_9427);
and U10799 (N_10799,N_10346,N_9012);
and U10800 (N_10800,N_9825,N_9469);
nand U10801 (N_10801,N_9185,N_9603);
or U10802 (N_10802,N_10077,N_10452);
nor U10803 (N_10803,N_9008,N_9628);
xor U10804 (N_10804,N_9792,N_9630);
nand U10805 (N_10805,N_9668,N_9233);
nor U10806 (N_10806,N_9052,N_9221);
nor U10807 (N_10807,N_10024,N_9264);
nand U10808 (N_10808,N_9849,N_9705);
nor U10809 (N_10809,N_10116,N_9881);
or U10810 (N_10810,N_10256,N_9304);
or U10811 (N_10811,N_9555,N_9054);
nand U10812 (N_10812,N_9844,N_10466);
and U10813 (N_10813,N_9634,N_9239);
nor U10814 (N_10814,N_9508,N_10401);
nor U10815 (N_10815,N_10439,N_10435);
nand U10816 (N_10816,N_9323,N_10377);
nor U10817 (N_10817,N_9829,N_9553);
nand U10818 (N_10818,N_10090,N_10127);
or U10819 (N_10819,N_10414,N_10174);
or U10820 (N_10820,N_10371,N_9403);
and U10821 (N_10821,N_10407,N_9606);
and U10822 (N_10822,N_9146,N_10022);
or U10823 (N_10823,N_9296,N_9429);
nand U10824 (N_10824,N_9654,N_9770);
nor U10825 (N_10825,N_10391,N_9170);
nand U10826 (N_10826,N_9152,N_9778);
nand U10827 (N_10827,N_9139,N_9546);
xor U10828 (N_10828,N_10450,N_9572);
nand U10829 (N_10829,N_9130,N_9856);
and U10830 (N_10830,N_10456,N_10402);
and U10831 (N_10831,N_9350,N_9746);
or U10832 (N_10832,N_9309,N_10483);
and U10833 (N_10833,N_9267,N_9408);
and U10834 (N_10834,N_9882,N_9798);
and U10835 (N_10835,N_9821,N_10362);
nor U10836 (N_10836,N_9249,N_9987);
nor U10837 (N_10837,N_10374,N_9162);
xor U10838 (N_10838,N_9277,N_9193);
nand U10839 (N_10839,N_9073,N_10115);
xnor U10840 (N_10840,N_9436,N_9711);
nor U10841 (N_10841,N_9197,N_9080);
or U10842 (N_10842,N_9394,N_9386);
or U10843 (N_10843,N_10417,N_9108);
and U10844 (N_10844,N_10002,N_9346);
nor U10845 (N_10845,N_10494,N_9303);
nand U10846 (N_10846,N_10084,N_9088);
nor U10847 (N_10847,N_9674,N_9450);
or U10848 (N_10848,N_10111,N_10070);
nor U10849 (N_10849,N_10162,N_9348);
or U10850 (N_10850,N_10282,N_10003);
nand U10851 (N_10851,N_10066,N_9160);
and U10852 (N_10852,N_9345,N_9010);
xor U10853 (N_10853,N_9092,N_9307);
or U10854 (N_10854,N_10275,N_10324);
xor U10855 (N_10855,N_10224,N_9980);
or U10856 (N_10856,N_10298,N_9129);
or U10857 (N_10857,N_10231,N_9733);
xnor U10858 (N_10858,N_9894,N_9382);
xnor U10859 (N_10859,N_9597,N_10051);
nor U10860 (N_10860,N_9254,N_9961);
xnor U10861 (N_10861,N_10216,N_9757);
and U10862 (N_10862,N_10117,N_9200);
nand U10863 (N_10863,N_9870,N_9219);
or U10864 (N_10864,N_10009,N_10093);
nand U10865 (N_10865,N_9612,N_9731);
and U10866 (N_10866,N_9332,N_9138);
and U10867 (N_10867,N_10230,N_9161);
nor U10868 (N_10868,N_9588,N_10021);
or U10869 (N_10869,N_9996,N_9522);
nor U10870 (N_10870,N_9158,N_9110);
or U10871 (N_10871,N_9212,N_10314);
nor U10872 (N_10872,N_10114,N_10445);
xor U10873 (N_10873,N_9071,N_9501);
xor U10874 (N_10874,N_9482,N_9692);
and U10875 (N_10875,N_10477,N_10212);
or U10876 (N_10876,N_10106,N_10467);
nand U10877 (N_10877,N_9287,N_10135);
xnor U10878 (N_10878,N_9218,N_9647);
or U10879 (N_10879,N_9534,N_10185);
xnor U10880 (N_10880,N_9729,N_9075);
nand U10881 (N_10881,N_9257,N_10031);
and U10882 (N_10882,N_10153,N_9217);
or U10883 (N_10883,N_9698,N_10370);
nand U10884 (N_10884,N_10351,N_10418);
nor U10885 (N_10885,N_9914,N_9838);
or U10886 (N_10886,N_9684,N_10262);
nor U10887 (N_10887,N_9237,N_9791);
nand U10888 (N_10888,N_9815,N_9024);
nor U10889 (N_10889,N_9678,N_9615);
nor U10890 (N_10890,N_10019,N_9454);
nand U10891 (N_10891,N_9985,N_10381);
or U10892 (N_10892,N_9560,N_9335);
nand U10893 (N_10893,N_9072,N_10470);
nor U10894 (N_10894,N_9276,N_9610);
xor U10895 (N_10895,N_9544,N_9418);
and U10896 (N_10896,N_9683,N_10169);
xor U10897 (N_10897,N_9689,N_9558);
nor U10898 (N_10898,N_9827,N_9086);
or U10899 (N_10899,N_9511,N_9274);
or U10900 (N_10900,N_10147,N_10284);
and U10901 (N_10901,N_10410,N_9800);
or U10902 (N_10902,N_9842,N_9643);
xnor U10903 (N_10903,N_9251,N_9425);
xnor U10904 (N_10904,N_9169,N_10245);
nand U10905 (N_10905,N_9016,N_9283);
nor U10906 (N_10906,N_9314,N_9889);
nor U10907 (N_10907,N_9465,N_9960);
and U10908 (N_10908,N_10207,N_9962);
xor U10909 (N_10909,N_9972,N_9320);
and U10910 (N_10910,N_9780,N_9616);
and U10911 (N_10911,N_10434,N_10020);
or U10912 (N_10912,N_9794,N_9929);
nor U10913 (N_10913,N_10061,N_10342);
xnor U10914 (N_10914,N_10438,N_10139);
xnor U10915 (N_10915,N_9467,N_9248);
xor U10916 (N_10916,N_9119,N_10243);
nor U10917 (N_10917,N_9795,N_9325);
nand U10918 (N_10918,N_9496,N_10484);
nor U10919 (N_10919,N_9273,N_10025);
and U10920 (N_10920,N_9141,N_10321);
or U10921 (N_10921,N_9401,N_9126);
nor U10922 (N_10922,N_9775,N_9608);
and U10923 (N_10923,N_9491,N_10383);
nand U10924 (N_10924,N_9330,N_10012);
xnor U10925 (N_10925,N_9565,N_9172);
nor U10926 (N_10926,N_10192,N_9227);
and U10927 (N_10927,N_9027,N_10393);
xor U10928 (N_10928,N_10499,N_10015);
or U10929 (N_10929,N_9397,N_10269);
and U10930 (N_10930,N_9832,N_10102);
nor U10931 (N_10931,N_10415,N_9417);
and U10932 (N_10932,N_10305,N_9066);
nand U10933 (N_10933,N_10403,N_9128);
or U10934 (N_10934,N_9621,N_10478);
nand U10935 (N_10935,N_9662,N_9039);
nand U10936 (N_10936,N_9788,N_9145);
nor U10937 (N_10937,N_10058,N_9224);
xor U10938 (N_10938,N_9723,N_9341);
nor U10939 (N_10939,N_9975,N_9057);
and U10940 (N_10940,N_9214,N_10080);
xor U10941 (N_10941,N_9749,N_9958);
and U10942 (N_10942,N_10238,N_9466);
nor U10943 (N_10943,N_9388,N_10161);
nand U10944 (N_10944,N_10399,N_9028);
nor U10945 (N_10945,N_10167,N_9725);
xor U10946 (N_10946,N_9516,N_9266);
xor U10947 (N_10947,N_9916,N_9065);
xor U10948 (N_10948,N_9755,N_9041);
nor U10949 (N_10949,N_9532,N_9202);
or U10950 (N_10950,N_9582,N_9104);
or U10951 (N_10951,N_9451,N_9426);
or U10952 (N_10952,N_9893,N_9011);
xnor U10953 (N_10953,N_9990,N_9253);
and U10954 (N_10954,N_9624,N_9563);
or U10955 (N_10955,N_9586,N_9814);
or U10956 (N_10956,N_9374,N_9781);
or U10957 (N_10957,N_10236,N_9383);
and U10958 (N_10958,N_10267,N_9556);
and U10959 (N_10959,N_10250,N_10068);
or U10960 (N_10960,N_10232,N_9142);
nor U10961 (N_10961,N_10317,N_9679);
and U10962 (N_10962,N_9005,N_9897);
and U10963 (N_10963,N_10437,N_10219);
nor U10964 (N_10964,N_9448,N_10217);
xor U10965 (N_10965,N_10355,N_9009);
and U10966 (N_10966,N_10050,N_9869);
or U10967 (N_10967,N_9766,N_10196);
xor U10968 (N_10968,N_9157,N_9007);
and U10969 (N_10969,N_10233,N_9306);
or U10970 (N_10970,N_9823,N_9531);
nand U10971 (N_10971,N_10040,N_9539);
nor U10972 (N_10972,N_9375,N_9422);
xor U10973 (N_10973,N_9497,N_9651);
xnor U10974 (N_10974,N_10182,N_10246);
nand U10975 (N_10975,N_10485,N_9067);
xnor U10976 (N_10976,N_9095,N_10113);
and U10977 (N_10977,N_10201,N_10159);
and U10978 (N_10978,N_10056,N_9477);
or U10979 (N_10979,N_9268,N_9742);
nand U10980 (N_10980,N_10241,N_9732);
or U10981 (N_10981,N_9690,N_9512);
nor U10982 (N_10982,N_10251,N_9601);
or U10983 (N_10983,N_10448,N_9247);
xnor U10984 (N_10984,N_9085,N_9453);
and U10985 (N_10985,N_9056,N_9292);
nand U10986 (N_10986,N_9331,N_10425);
or U10987 (N_10987,N_10023,N_9082);
nor U10988 (N_10988,N_10082,N_9098);
nand U10989 (N_10989,N_9589,N_9324);
xor U10990 (N_10990,N_9506,N_10146);
and U10991 (N_10991,N_9090,N_10013);
and U10992 (N_10992,N_9363,N_10100);
and U10993 (N_10993,N_9691,N_9263);
xor U10994 (N_10994,N_10078,N_9578);
and U10995 (N_10995,N_9874,N_10069);
nor U10996 (N_10996,N_9898,N_9412);
nand U10997 (N_10997,N_9151,N_9149);
and U10998 (N_10998,N_9312,N_10455);
xnor U10999 (N_10999,N_9751,N_9688);
xnor U11000 (N_11000,N_9930,N_9627);
nor U11001 (N_11001,N_9502,N_10440);
xnor U11002 (N_11002,N_10033,N_9526);
nand U11003 (N_11003,N_9286,N_9566);
xor U11004 (N_11004,N_9727,N_9964);
and U11005 (N_11005,N_9226,N_10105);
and U11006 (N_11006,N_10306,N_9892);
xnor U11007 (N_11007,N_9722,N_9971);
xnor U11008 (N_11008,N_9569,N_9726);
or U11009 (N_11009,N_9681,N_9333);
nor U11010 (N_11010,N_10026,N_9359);
or U11011 (N_11011,N_10175,N_10386);
nor U11012 (N_11012,N_9660,N_9035);
or U11013 (N_11013,N_9896,N_9025);
and U11014 (N_11014,N_9672,N_9362);
nand U11015 (N_11015,N_10380,N_9031);
nor U11016 (N_11016,N_9201,N_9904);
nor U11017 (N_11017,N_10032,N_10479);
xnor U11018 (N_11018,N_9641,N_9431);
nor U11019 (N_11019,N_9061,N_9579);
nor U11020 (N_11020,N_9476,N_10089);
or U11021 (N_11021,N_9243,N_10367);
or U11022 (N_11022,N_10311,N_9639);
or U11023 (N_11023,N_10129,N_10472);
nand U11024 (N_11024,N_9282,N_10244);
nor U11025 (N_11025,N_9979,N_9000);
and U11026 (N_11026,N_10375,N_9014);
or U11027 (N_11027,N_9848,N_9538);
or U11028 (N_11028,N_9982,N_10188);
nor U11029 (N_11029,N_10181,N_9183);
nor U11030 (N_11030,N_10491,N_10287);
xor U11031 (N_11031,N_9017,N_10206);
and U11032 (N_11032,N_10291,N_9604);
xor U11033 (N_11033,N_9032,N_10214);
and U11034 (N_11034,N_10164,N_9470);
xnor U11035 (N_11035,N_10288,N_9038);
or U11036 (N_11036,N_10411,N_9756);
nand U11037 (N_11037,N_9405,N_10463);
and U11038 (N_11038,N_9988,N_9619);
xor U11039 (N_11039,N_9369,N_9753);
nand U11040 (N_11040,N_10014,N_10270);
nand U11041 (N_11041,N_10301,N_10254);
and U11042 (N_11042,N_9131,N_9599);
and U11043 (N_11043,N_9381,N_10299);
and U11044 (N_11044,N_10208,N_9887);
nand U11045 (N_11045,N_9474,N_10289);
and U11046 (N_11046,N_10308,N_10398);
xnor U11047 (N_11047,N_10073,N_9393);
xor U11048 (N_11048,N_10327,N_10442);
and U11049 (N_11049,N_9880,N_10018);
nand U11050 (N_11050,N_10122,N_10186);
nand U11051 (N_11051,N_10360,N_9295);
nand U11052 (N_11052,N_10373,N_10482);
nor U11053 (N_11053,N_9826,N_9120);
nor U11054 (N_11054,N_10062,N_9045);
nand U11055 (N_11055,N_9934,N_9857);
or U11056 (N_11056,N_9356,N_10474);
and U11057 (N_11057,N_9190,N_9706);
nand U11058 (N_11058,N_9339,N_9697);
nor U11059 (N_11059,N_9334,N_9402);
xnor U11060 (N_11060,N_10497,N_10054);
nor U11061 (N_11061,N_9550,N_9042);
nor U11062 (N_11062,N_9910,N_9293);
or U11063 (N_11063,N_10158,N_10165);
and U11064 (N_11064,N_10195,N_9472);
or U11065 (N_11065,N_9441,N_9940);
xnor U11066 (N_11066,N_9316,N_9428);
or U11067 (N_11067,N_10155,N_10451);
nand U11068 (N_11068,N_9784,N_9931);
nand U11069 (N_11069,N_9718,N_10000);
nor U11070 (N_11070,N_9484,N_9481);
nor U11071 (N_11071,N_9117,N_9717);
nor U11072 (N_11072,N_9576,N_9093);
nand U11073 (N_11073,N_9208,N_9235);
nand U11074 (N_11074,N_9365,N_9290);
xor U11075 (N_11075,N_9549,N_9884);
xor U11076 (N_11076,N_9216,N_9854);
nand U11077 (N_11077,N_9322,N_10049);
xor U11078 (N_11078,N_9116,N_9716);
nand U11079 (N_11079,N_10183,N_9455);
nand U11080 (N_11080,N_9571,N_9671);
and U11081 (N_11081,N_9371,N_9864);
and U11082 (N_11082,N_9400,N_9626);
nor U11083 (N_11083,N_9976,N_9059);
and U11084 (N_11084,N_9411,N_9420);
or U11085 (N_11085,N_9632,N_9458);
nor U11086 (N_11086,N_10087,N_10043);
nor U11087 (N_11087,N_9064,N_9994);
nor U11088 (N_11088,N_9525,N_10126);
xnor U11089 (N_11089,N_9840,N_9888);
xor U11090 (N_11090,N_9877,N_9310);
or U11091 (N_11091,N_10140,N_10007);
nor U11092 (N_11092,N_9416,N_10044);
or U11093 (N_11093,N_10400,N_9847);
nand U11094 (N_11094,N_10145,N_9950);
nor U11095 (N_11095,N_9741,N_10343);
and U11096 (N_11096,N_9622,N_9665);
xnor U11097 (N_11097,N_9696,N_9876);
nor U11098 (N_11098,N_10057,N_9029);
nor U11099 (N_11099,N_9521,N_10389);
and U11100 (N_11100,N_10092,N_9570);
and U11101 (N_11101,N_9559,N_9315);
and U11102 (N_11102,N_9194,N_9241);
nor U11103 (N_11103,N_9279,N_9944);
nor U11104 (N_11104,N_10151,N_9759);
and U11105 (N_11105,N_9518,N_10086);
or U11106 (N_11106,N_10464,N_9236);
nand U11107 (N_11107,N_9670,N_9366);
or U11108 (N_11108,N_9094,N_10228);
nor U11109 (N_11109,N_9824,N_10390);
and U11110 (N_11110,N_9270,N_9318);
or U11111 (N_11111,N_10071,N_10315);
nor U11112 (N_11112,N_9577,N_9631);
nor U11113 (N_11113,N_9959,N_9367);
or U11114 (N_11114,N_10211,N_10460);
and U11115 (N_11115,N_9811,N_9650);
or U11116 (N_11116,N_9762,N_10326);
xnor U11117 (N_11117,N_9136,N_10104);
nand U11118 (N_11118,N_9392,N_10295);
and U11119 (N_11119,N_10091,N_10142);
or U11120 (N_11120,N_10394,N_9783);
nor U11121 (N_11121,N_10255,N_9686);
nor U11122 (N_11122,N_9514,N_9203);
and U11123 (N_11123,N_9147,N_9941);
xor U11124 (N_11124,N_9957,N_9021);
and U11125 (N_11125,N_10454,N_9414);
nor U11126 (N_11126,N_9424,N_10323);
and U11127 (N_11127,N_10405,N_9289);
nand U11128 (N_11128,N_9779,N_9376);
nand U11129 (N_11129,N_9109,N_10436);
or U11130 (N_11130,N_9019,N_10281);
nand U11131 (N_11131,N_10364,N_9176);
nand U11132 (N_11132,N_9089,N_10096);
nand U11133 (N_11133,N_9378,N_9372);
nor U11134 (N_11134,N_9228,N_10112);
nand U11135 (N_11135,N_10237,N_9790);
nand U11136 (N_11136,N_9906,N_9519);
or U11137 (N_11137,N_9859,N_9728);
nand U11138 (N_11138,N_9444,N_10226);
nand U11139 (N_11139,N_9739,N_9199);
nor U11140 (N_11140,N_9291,N_9721);
nand U11141 (N_11141,N_9772,N_10413);
nand U11142 (N_11142,N_10193,N_10075);
nand U11143 (N_11143,N_10444,N_10004);
or U11144 (N_11144,N_9473,N_10029);
and U11145 (N_11145,N_9907,N_9855);
nor U11146 (N_11146,N_9839,N_9993);
nor U11147 (N_11147,N_10171,N_9207);
xor U11148 (N_11148,N_9707,N_10088);
and U11149 (N_11149,N_9719,N_9410);
and U11150 (N_11150,N_9261,N_9812);
nor U11151 (N_11151,N_9479,N_10190);
nor U11152 (N_11152,N_10163,N_9584);
or U11153 (N_11153,N_9885,N_9154);
and U11154 (N_11154,N_10101,N_10118);
xnor U11155 (N_11155,N_10347,N_10257);
xnor U11156 (N_11156,N_9231,N_10047);
and U11157 (N_11157,N_10353,N_9238);
and U11158 (N_11158,N_9527,N_9714);
and U11159 (N_11159,N_9936,N_9773);
and U11160 (N_11160,N_9983,N_10172);
or U11161 (N_11161,N_9223,N_9122);
nand U11162 (N_11162,N_9034,N_9373);
or U11163 (N_11163,N_9495,N_9598);
or U11164 (N_11164,N_9220,N_10060);
xnor U11165 (N_11165,N_9159,N_10408);
xnor U11166 (N_11166,N_9143,N_10319);
or U11167 (N_11167,N_10010,N_10268);
nand U11168 (N_11168,N_9677,N_10372);
nor U11169 (N_11169,N_10072,N_9977);
xnor U11170 (N_11170,N_9187,N_9917);
xor U11171 (N_11171,N_10481,N_9636);
nand U11172 (N_11172,N_9748,N_9259);
nor U11173 (N_11173,N_9694,N_9493);
or U11174 (N_11174,N_9902,N_9432);
nor U11175 (N_11175,N_9771,N_9752);
and U11176 (N_11176,N_9329,N_9487);
and U11177 (N_11177,N_10462,N_9984);
or U11178 (N_11178,N_10121,N_9564);
nand U11179 (N_11179,N_10252,N_10120);
nor U11180 (N_11180,N_10001,N_9213);
and U11181 (N_11181,N_10341,N_9583);
nand U11182 (N_11182,N_10141,N_10203);
and U11183 (N_11183,N_9494,N_10322);
or U11184 (N_11184,N_10487,N_9653);
nand U11185 (N_11185,N_9460,N_9013);
and U11186 (N_11186,N_10366,N_10359);
nor U11187 (N_11187,N_9843,N_9945);
xnor U11188 (N_11188,N_9536,N_10406);
xnor U11189 (N_11189,N_10357,N_9901);
and U11190 (N_11190,N_10471,N_9515);
or U11191 (N_11191,N_9900,N_10495);
and U11192 (N_11192,N_9806,N_9796);
nor U11193 (N_11193,N_9642,N_10333);
nand U11194 (N_11194,N_9328,N_10110);
xnor U11195 (N_11195,N_9480,N_9097);
nor U11196 (N_11196,N_9995,N_10099);
xor U11197 (N_11197,N_9761,N_10008);
nor U11198 (N_11198,N_10094,N_9198);
nand U11199 (N_11199,N_10496,N_9793);
or U11200 (N_11200,N_9240,N_9419);
or U11201 (N_11201,N_9561,N_9879);
and U11202 (N_11202,N_9883,N_9391);
xnor U11203 (N_11203,N_9140,N_9524);
and U11204 (N_11204,N_10345,N_10177);
and U11205 (N_11205,N_9281,N_10332);
nor U11206 (N_11206,N_9970,N_9357);
and U11207 (N_11207,N_9215,N_9053);
xnor U11208 (N_11208,N_9387,N_9805);
nand U11209 (N_11209,N_10294,N_10187);
nor U11210 (N_11210,N_9890,N_9409);
nor U11211 (N_11211,N_9992,N_10320);
xnor U11212 (N_11212,N_9048,N_9623);
nand U11213 (N_11213,N_10109,N_10264);
and U11214 (N_11214,N_9590,N_9150);
and U11215 (N_11215,N_9505,N_10227);
nand U11216 (N_11216,N_9319,N_9058);
nand U11217 (N_11217,N_10199,N_9922);
nand U11218 (N_11218,N_9649,N_9342);
or U11219 (N_11219,N_10157,N_9327);
xnor U11220 (N_11220,N_9768,N_9764);
nor U11221 (N_11221,N_9918,N_9644);
or U11222 (N_11222,N_10476,N_9360);
or U11223 (N_11223,N_10329,N_10465);
and U11224 (N_11224,N_9148,N_9175);
or U11225 (N_11225,N_9845,N_10328);
nor U11226 (N_11226,N_10042,N_9540);
and U11227 (N_11227,N_10119,N_9517);
nor U11228 (N_11228,N_10045,N_10234);
xnor U11229 (N_11229,N_9195,N_9284);
and U11230 (N_11230,N_10337,N_9656);
or U11231 (N_11231,N_9033,N_9078);
nor U11232 (N_11232,N_9102,N_10132);
or U11233 (N_11233,N_9510,N_9981);
or U11234 (N_11234,N_9338,N_9250);
nand U11235 (N_11235,N_10396,N_9230);
or U11236 (N_11236,N_9853,N_10409);
nor U11237 (N_11237,N_9594,N_9693);
xor U11238 (N_11238,N_9833,N_9602);
or U11239 (N_11239,N_10292,N_9115);
nand U11240 (N_11240,N_9963,N_10191);
and U11241 (N_11241,N_10278,N_9275);
or U11242 (N_11242,N_10067,N_10309);
nand U11243 (N_11243,N_9317,N_9351);
xnor U11244 (N_11244,N_10247,N_10420);
xnor U11245 (N_11245,N_9438,N_10486);
nor U11246 (N_11246,N_9542,N_9614);
nand U11247 (N_11247,N_10133,N_10160);
and U11248 (N_11248,N_9659,N_9528);
or U11249 (N_11249,N_10335,N_9184);
nor U11250 (N_11250,N_9190,N_9262);
nor U11251 (N_11251,N_9097,N_10472);
xnor U11252 (N_11252,N_10060,N_9057);
nor U11253 (N_11253,N_9518,N_9751);
nand U11254 (N_11254,N_9107,N_9513);
nor U11255 (N_11255,N_10428,N_9191);
xor U11256 (N_11256,N_9598,N_9914);
or U11257 (N_11257,N_9581,N_9058);
nor U11258 (N_11258,N_9833,N_9036);
or U11259 (N_11259,N_10242,N_9606);
xnor U11260 (N_11260,N_9857,N_10213);
xnor U11261 (N_11261,N_9385,N_9333);
xor U11262 (N_11262,N_9730,N_9067);
nor U11263 (N_11263,N_9220,N_9074);
nand U11264 (N_11264,N_10158,N_10428);
nand U11265 (N_11265,N_9541,N_9619);
nor U11266 (N_11266,N_10330,N_9227);
xor U11267 (N_11267,N_9214,N_10227);
and U11268 (N_11268,N_9505,N_10077);
and U11269 (N_11269,N_9392,N_10085);
nand U11270 (N_11270,N_9703,N_9370);
and U11271 (N_11271,N_9455,N_9910);
nand U11272 (N_11272,N_10169,N_9942);
nand U11273 (N_11273,N_9369,N_9672);
nand U11274 (N_11274,N_9774,N_9500);
or U11275 (N_11275,N_10225,N_10055);
nand U11276 (N_11276,N_9478,N_10172);
nand U11277 (N_11277,N_10094,N_9877);
or U11278 (N_11278,N_9000,N_9999);
or U11279 (N_11279,N_9719,N_10178);
nand U11280 (N_11280,N_9285,N_9775);
nor U11281 (N_11281,N_9483,N_9504);
nand U11282 (N_11282,N_9793,N_9035);
xor U11283 (N_11283,N_10006,N_9212);
xor U11284 (N_11284,N_9792,N_10391);
nor U11285 (N_11285,N_9637,N_9077);
nand U11286 (N_11286,N_9691,N_10114);
nor U11287 (N_11287,N_10343,N_9399);
or U11288 (N_11288,N_9541,N_10270);
nand U11289 (N_11289,N_9209,N_9370);
xnor U11290 (N_11290,N_9431,N_9930);
nor U11291 (N_11291,N_9389,N_10126);
xor U11292 (N_11292,N_10474,N_10098);
and U11293 (N_11293,N_10069,N_9830);
nand U11294 (N_11294,N_9397,N_9265);
or U11295 (N_11295,N_9573,N_9374);
nor U11296 (N_11296,N_9026,N_9672);
nor U11297 (N_11297,N_9405,N_9716);
nand U11298 (N_11298,N_9643,N_9852);
nand U11299 (N_11299,N_9541,N_9397);
xnor U11300 (N_11300,N_9672,N_9050);
or U11301 (N_11301,N_10169,N_9066);
xor U11302 (N_11302,N_9264,N_9929);
xor U11303 (N_11303,N_9642,N_9362);
nand U11304 (N_11304,N_10318,N_9641);
xnor U11305 (N_11305,N_10417,N_9572);
nor U11306 (N_11306,N_9906,N_9811);
nor U11307 (N_11307,N_10282,N_9061);
nor U11308 (N_11308,N_9988,N_9075);
and U11309 (N_11309,N_9951,N_9035);
xnor U11310 (N_11310,N_10372,N_9287);
nor U11311 (N_11311,N_10367,N_10187);
nand U11312 (N_11312,N_9242,N_9362);
nor U11313 (N_11313,N_10116,N_10368);
and U11314 (N_11314,N_10478,N_10049);
nand U11315 (N_11315,N_10374,N_9084);
xor U11316 (N_11316,N_9574,N_9476);
and U11317 (N_11317,N_10104,N_9509);
nor U11318 (N_11318,N_9244,N_9203);
nand U11319 (N_11319,N_10093,N_9663);
nand U11320 (N_11320,N_9967,N_9493);
nand U11321 (N_11321,N_9976,N_9002);
and U11322 (N_11322,N_10177,N_9931);
or U11323 (N_11323,N_10239,N_10065);
nor U11324 (N_11324,N_10353,N_10147);
xor U11325 (N_11325,N_9301,N_10465);
xor U11326 (N_11326,N_9873,N_10317);
or U11327 (N_11327,N_10342,N_9377);
and U11328 (N_11328,N_10310,N_9875);
nand U11329 (N_11329,N_9702,N_9547);
and U11330 (N_11330,N_9484,N_10015);
xnor U11331 (N_11331,N_10289,N_9908);
nand U11332 (N_11332,N_9281,N_10368);
nor U11333 (N_11333,N_9544,N_9840);
nor U11334 (N_11334,N_10012,N_9301);
nor U11335 (N_11335,N_9251,N_9431);
nor U11336 (N_11336,N_10065,N_9268);
nand U11337 (N_11337,N_9699,N_9441);
xnor U11338 (N_11338,N_10472,N_9553);
nor U11339 (N_11339,N_9415,N_9432);
or U11340 (N_11340,N_9883,N_9357);
nand U11341 (N_11341,N_9943,N_9890);
and U11342 (N_11342,N_9165,N_9727);
nand U11343 (N_11343,N_9735,N_9775);
or U11344 (N_11344,N_10136,N_10326);
xor U11345 (N_11345,N_9505,N_9124);
and U11346 (N_11346,N_9933,N_10303);
nand U11347 (N_11347,N_10145,N_9688);
nand U11348 (N_11348,N_10441,N_9225);
nor U11349 (N_11349,N_9439,N_9602);
nand U11350 (N_11350,N_9455,N_10238);
nand U11351 (N_11351,N_9732,N_10487);
and U11352 (N_11352,N_9529,N_10344);
or U11353 (N_11353,N_10287,N_9878);
and U11354 (N_11354,N_9501,N_10100);
and U11355 (N_11355,N_9427,N_10191);
nor U11356 (N_11356,N_9672,N_10086);
and U11357 (N_11357,N_9667,N_9646);
nor U11358 (N_11358,N_9897,N_10436);
xnor U11359 (N_11359,N_10085,N_10001);
nor U11360 (N_11360,N_10270,N_9752);
nor U11361 (N_11361,N_9917,N_9708);
or U11362 (N_11362,N_9639,N_9713);
xnor U11363 (N_11363,N_10296,N_9364);
nor U11364 (N_11364,N_9061,N_9768);
xor U11365 (N_11365,N_9262,N_10153);
nor U11366 (N_11366,N_10380,N_9349);
and U11367 (N_11367,N_9460,N_9412);
nand U11368 (N_11368,N_9544,N_9309);
xnor U11369 (N_11369,N_9568,N_10078);
nor U11370 (N_11370,N_9287,N_9720);
or U11371 (N_11371,N_9776,N_9151);
and U11372 (N_11372,N_9640,N_9038);
or U11373 (N_11373,N_9388,N_9770);
and U11374 (N_11374,N_9276,N_10129);
nand U11375 (N_11375,N_9604,N_9780);
nand U11376 (N_11376,N_9256,N_9966);
nand U11377 (N_11377,N_9017,N_9551);
and U11378 (N_11378,N_9987,N_9033);
xnor U11379 (N_11379,N_9087,N_9142);
nor U11380 (N_11380,N_9702,N_10143);
or U11381 (N_11381,N_10357,N_9436);
or U11382 (N_11382,N_9007,N_9804);
nor U11383 (N_11383,N_10098,N_10019);
and U11384 (N_11384,N_9067,N_10328);
and U11385 (N_11385,N_9038,N_9053);
xnor U11386 (N_11386,N_9130,N_9391);
nand U11387 (N_11387,N_10434,N_10388);
or U11388 (N_11388,N_9324,N_9247);
xor U11389 (N_11389,N_9478,N_9346);
nand U11390 (N_11390,N_9125,N_10299);
nand U11391 (N_11391,N_10141,N_10419);
and U11392 (N_11392,N_10276,N_10028);
xnor U11393 (N_11393,N_9111,N_9866);
nor U11394 (N_11394,N_10496,N_9506);
or U11395 (N_11395,N_10112,N_10187);
nor U11396 (N_11396,N_10073,N_9577);
xnor U11397 (N_11397,N_9375,N_10057);
nand U11398 (N_11398,N_9336,N_10030);
nand U11399 (N_11399,N_10158,N_9263);
nand U11400 (N_11400,N_9654,N_9782);
or U11401 (N_11401,N_10009,N_9286);
and U11402 (N_11402,N_10189,N_9458);
or U11403 (N_11403,N_9878,N_9756);
nand U11404 (N_11404,N_9043,N_9379);
nand U11405 (N_11405,N_10134,N_9911);
or U11406 (N_11406,N_10457,N_10245);
nand U11407 (N_11407,N_9872,N_10283);
and U11408 (N_11408,N_10099,N_9021);
nand U11409 (N_11409,N_9166,N_9874);
and U11410 (N_11410,N_10387,N_10014);
xor U11411 (N_11411,N_9291,N_9371);
and U11412 (N_11412,N_9541,N_10403);
and U11413 (N_11413,N_9151,N_10039);
xnor U11414 (N_11414,N_9181,N_10232);
xnor U11415 (N_11415,N_9373,N_9809);
or U11416 (N_11416,N_9541,N_9431);
or U11417 (N_11417,N_9282,N_10477);
or U11418 (N_11418,N_9048,N_9822);
and U11419 (N_11419,N_9236,N_9349);
nand U11420 (N_11420,N_9546,N_9892);
xor U11421 (N_11421,N_9370,N_9291);
nand U11422 (N_11422,N_9798,N_9455);
nor U11423 (N_11423,N_9827,N_9141);
nand U11424 (N_11424,N_9483,N_9660);
or U11425 (N_11425,N_9121,N_9150);
xor U11426 (N_11426,N_9034,N_10423);
or U11427 (N_11427,N_9474,N_9947);
and U11428 (N_11428,N_9382,N_10401);
or U11429 (N_11429,N_10090,N_9094);
and U11430 (N_11430,N_9658,N_9458);
nand U11431 (N_11431,N_9265,N_9492);
nor U11432 (N_11432,N_9135,N_9463);
xnor U11433 (N_11433,N_10207,N_10021);
nand U11434 (N_11434,N_10017,N_10409);
nand U11435 (N_11435,N_9281,N_9082);
nor U11436 (N_11436,N_10198,N_10298);
nand U11437 (N_11437,N_9500,N_9136);
nand U11438 (N_11438,N_10392,N_10430);
xnor U11439 (N_11439,N_10156,N_10297);
nand U11440 (N_11440,N_9617,N_9652);
and U11441 (N_11441,N_9914,N_10209);
and U11442 (N_11442,N_9211,N_9354);
nand U11443 (N_11443,N_9023,N_10419);
xor U11444 (N_11444,N_10460,N_9432);
and U11445 (N_11445,N_9258,N_9255);
or U11446 (N_11446,N_10204,N_9206);
nand U11447 (N_11447,N_9748,N_9004);
nand U11448 (N_11448,N_9547,N_9518);
nor U11449 (N_11449,N_9704,N_10328);
or U11450 (N_11450,N_9205,N_10194);
and U11451 (N_11451,N_9657,N_10223);
or U11452 (N_11452,N_10082,N_9892);
nor U11453 (N_11453,N_9479,N_10208);
xor U11454 (N_11454,N_9576,N_9877);
nor U11455 (N_11455,N_9729,N_9676);
nand U11456 (N_11456,N_9321,N_9238);
or U11457 (N_11457,N_9088,N_9197);
nand U11458 (N_11458,N_10346,N_10285);
nor U11459 (N_11459,N_9060,N_9541);
or U11460 (N_11460,N_10329,N_9661);
or U11461 (N_11461,N_9720,N_10270);
and U11462 (N_11462,N_9538,N_9827);
nor U11463 (N_11463,N_10347,N_10173);
xnor U11464 (N_11464,N_9316,N_9596);
nand U11465 (N_11465,N_9867,N_10335);
nand U11466 (N_11466,N_9142,N_9243);
xor U11467 (N_11467,N_10170,N_10484);
or U11468 (N_11468,N_9489,N_9529);
nand U11469 (N_11469,N_9333,N_10224);
or U11470 (N_11470,N_9792,N_9049);
nand U11471 (N_11471,N_10270,N_9909);
xor U11472 (N_11472,N_10060,N_9050);
xnor U11473 (N_11473,N_9982,N_10204);
and U11474 (N_11474,N_9446,N_10234);
xnor U11475 (N_11475,N_9076,N_9985);
nor U11476 (N_11476,N_9858,N_9822);
and U11477 (N_11477,N_9618,N_9927);
nand U11478 (N_11478,N_9397,N_9401);
and U11479 (N_11479,N_9225,N_9462);
xnor U11480 (N_11480,N_10271,N_9940);
and U11481 (N_11481,N_10078,N_10393);
or U11482 (N_11482,N_9513,N_9974);
and U11483 (N_11483,N_9145,N_9823);
nand U11484 (N_11484,N_10285,N_9393);
xor U11485 (N_11485,N_10431,N_9088);
nor U11486 (N_11486,N_10480,N_9109);
or U11487 (N_11487,N_9247,N_9424);
xor U11488 (N_11488,N_9450,N_9780);
or U11489 (N_11489,N_9420,N_9442);
nor U11490 (N_11490,N_9741,N_10083);
nand U11491 (N_11491,N_9223,N_9692);
or U11492 (N_11492,N_9211,N_9425);
or U11493 (N_11493,N_9022,N_9116);
nand U11494 (N_11494,N_9872,N_10420);
nand U11495 (N_11495,N_9188,N_9928);
nand U11496 (N_11496,N_9983,N_9994);
and U11497 (N_11497,N_9942,N_9972);
or U11498 (N_11498,N_10146,N_9500);
nand U11499 (N_11499,N_9521,N_9256);
nor U11500 (N_11500,N_9558,N_9366);
xnor U11501 (N_11501,N_9997,N_9639);
and U11502 (N_11502,N_9897,N_9949);
nor U11503 (N_11503,N_10332,N_9495);
or U11504 (N_11504,N_9141,N_10312);
and U11505 (N_11505,N_9275,N_9313);
xor U11506 (N_11506,N_10441,N_9356);
xor U11507 (N_11507,N_9876,N_9481);
nand U11508 (N_11508,N_10116,N_10406);
or U11509 (N_11509,N_10034,N_10086);
nor U11510 (N_11510,N_9828,N_9476);
xnor U11511 (N_11511,N_10396,N_10000);
and U11512 (N_11512,N_9404,N_9662);
or U11513 (N_11513,N_9252,N_10101);
nand U11514 (N_11514,N_9444,N_9963);
and U11515 (N_11515,N_9715,N_9996);
nand U11516 (N_11516,N_10356,N_9235);
nand U11517 (N_11517,N_9563,N_9956);
xor U11518 (N_11518,N_9321,N_9192);
nor U11519 (N_11519,N_9702,N_9904);
or U11520 (N_11520,N_9688,N_9121);
xor U11521 (N_11521,N_9788,N_10046);
or U11522 (N_11522,N_9617,N_9846);
nor U11523 (N_11523,N_9637,N_10033);
nor U11524 (N_11524,N_9135,N_9037);
nor U11525 (N_11525,N_9118,N_9381);
xor U11526 (N_11526,N_9009,N_9513);
xnor U11527 (N_11527,N_10077,N_9811);
and U11528 (N_11528,N_9387,N_9202);
nand U11529 (N_11529,N_9622,N_9454);
or U11530 (N_11530,N_10097,N_9390);
nand U11531 (N_11531,N_9642,N_9123);
and U11532 (N_11532,N_9230,N_9332);
nor U11533 (N_11533,N_9337,N_9023);
and U11534 (N_11534,N_9716,N_10041);
xor U11535 (N_11535,N_9639,N_9906);
nor U11536 (N_11536,N_9882,N_9893);
and U11537 (N_11537,N_9426,N_9714);
and U11538 (N_11538,N_9874,N_9853);
and U11539 (N_11539,N_10084,N_9557);
nand U11540 (N_11540,N_9184,N_10047);
xnor U11541 (N_11541,N_10319,N_10143);
or U11542 (N_11542,N_10195,N_9758);
nor U11543 (N_11543,N_10345,N_9492);
or U11544 (N_11544,N_9454,N_10184);
or U11545 (N_11545,N_10346,N_9651);
or U11546 (N_11546,N_10107,N_10418);
nor U11547 (N_11547,N_9638,N_10316);
nor U11548 (N_11548,N_10197,N_9506);
nand U11549 (N_11549,N_10254,N_9082);
xor U11550 (N_11550,N_9002,N_10482);
or U11551 (N_11551,N_9928,N_10484);
nand U11552 (N_11552,N_10091,N_9711);
and U11553 (N_11553,N_10019,N_9793);
nor U11554 (N_11554,N_9434,N_9127);
xor U11555 (N_11555,N_9288,N_9999);
nand U11556 (N_11556,N_10095,N_9636);
or U11557 (N_11557,N_10390,N_9915);
xor U11558 (N_11558,N_10293,N_9678);
nand U11559 (N_11559,N_10067,N_9792);
and U11560 (N_11560,N_10021,N_10061);
or U11561 (N_11561,N_10163,N_9970);
and U11562 (N_11562,N_9878,N_10189);
nand U11563 (N_11563,N_9108,N_10291);
and U11564 (N_11564,N_10411,N_9400);
xor U11565 (N_11565,N_10342,N_10487);
or U11566 (N_11566,N_10232,N_10226);
nand U11567 (N_11567,N_9169,N_10361);
and U11568 (N_11568,N_9605,N_9925);
nor U11569 (N_11569,N_9670,N_9919);
nor U11570 (N_11570,N_9483,N_9009);
nand U11571 (N_11571,N_9166,N_9715);
or U11572 (N_11572,N_9098,N_10000);
and U11573 (N_11573,N_9440,N_10239);
xor U11574 (N_11574,N_9321,N_10347);
nand U11575 (N_11575,N_10362,N_9214);
nand U11576 (N_11576,N_9350,N_10474);
nor U11577 (N_11577,N_9147,N_9472);
nor U11578 (N_11578,N_10097,N_9658);
nor U11579 (N_11579,N_9339,N_9587);
nor U11580 (N_11580,N_10083,N_9785);
or U11581 (N_11581,N_9077,N_9557);
nor U11582 (N_11582,N_10015,N_9036);
or U11583 (N_11583,N_10160,N_9281);
nand U11584 (N_11584,N_9612,N_9352);
and U11585 (N_11585,N_9292,N_9865);
and U11586 (N_11586,N_9903,N_9898);
xor U11587 (N_11587,N_9312,N_9495);
or U11588 (N_11588,N_10390,N_10275);
nor U11589 (N_11589,N_9554,N_9957);
nor U11590 (N_11590,N_9735,N_9327);
and U11591 (N_11591,N_9719,N_9049);
nor U11592 (N_11592,N_10289,N_9345);
xnor U11593 (N_11593,N_10328,N_9923);
nand U11594 (N_11594,N_9096,N_9444);
xor U11595 (N_11595,N_10401,N_10493);
nor U11596 (N_11596,N_10451,N_10039);
nor U11597 (N_11597,N_9409,N_9903);
nor U11598 (N_11598,N_9195,N_9000);
or U11599 (N_11599,N_9409,N_9730);
nor U11600 (N_11600,N_9361,N_9937);
xnor U11601 (N_11601,N_9737,N_9591);
xor U11602 (N_11602,N_10274,N_9049);
or U11603 (N_11603,N_9119,N_9882);
or U11604 (N_11604,N_9412,N_9588);
nor U11605 (N_11605,N_9055,N_10204);
nand U11606 (N_11606,N_10432,N_10064);
and U11607 (N_11607,N_9310,N_9646);
nor U11608 (N_11608,N_10169,N_9186);
or U11609 (N_11609,N_9322,N_10339);
nand U11610 (N_11610,N_9259,N_9792);
xnor U11611 (N_11611,N_9767,N_9605);
xor U11612 (N_11612,N_9184,N_10466);
xnor U11613 (N_11613,N_9109,N_9935);
xnor U11614 (N_11614,N_9586,N_9633);
nor U11615 (N_11615,N_10074,N_9051);
or U11616 (N_11616,N_9357,N_9028);
or U11617 (N_11617,N_9407,N_10339);
or U11618 (N_11618,N_9817,N_9110);
nand U11619 (N_11619,N_9315,N_9482);
or U11620 (N_11620,N_10273,N_9013);
nor U11621 (N_11621,N_9451,N_10325);
and U11622 (N_11622,N_9211,N_9477);
and U11623 (N_11623,N_9121,N_10097);
or U11624 (N_11624,N_9129,N_10431);
nand U11625 (N_11625,N_10075,N_9532);
or U11626 (N_11626,N_9573,N_9289);
nand U11627 (N_11627,N_9500,N_9517);
or U11628 (N_11628,N_9028,N_9003);
or U11629 (N_11629,N_9758,N_9392);
xnor U11630 (N_11630,N_9556,N_9850);
and U11631 (N_11631,N_9424,N_10110);
xor U11632 (N_11632,N_9976,N_10466);
and U11633 (N_11633,N_10443,N_9643);
xor U11634 (N_11634,N_10131,N_9671);
and U11635 (N_11635,N_9159,N_9806);
nor U11636 (N_11636,N_10036,N_9816);
nand U11637 (N_11637,N_9284,N_9741);
or U11638 (N_11638,N_10333,N_10109);
and U11639 (N_11639,N_9294,N_9045);
xor U11640 (N_11640,N_9785,N_10233);
or U11641 (N_11641,N_9915,N_9492);
nor U11642 (N_11642,N_9217,N_9816);
xor U11643 (N_11643,N_9061,N_9045);
or U11644 (N_11644,N_9911,N_9203);
xnor U11645 (N_11645,N_9290,N_9703);
and U11646 (N_11646,N_9168,N_10476);
nor U11647 (N_11647,N_9691,N_10049);
or U11648 (N_11648,N_9728,N_9928);
or U11649 (N_11649,N_9724,N_9841);
nor U11650 (N_11650,N_9315,N_10450);
nor U11651 (N_11651,N_9558,N_9359);
or U11652 (N_11652,N_9291,N_10450);
and U11653 (N_11653,N_10037,N_9434);
nand U11654 (N_11654,N_9400,N_10174);
nor U11655 (N_11655,N_9445,N_9225);
xor U11656 (N_11656,N_9929,N_10077);
or U11657 (N_11657,N_9879,N_10026);
and U11658 (N_11658,N_9564,N_10495);
or U11659 (N_11659,N_10017,N_10330);
xnor U11660 (N_11660,N_10356,N_9103);
nor U11661 (N_11661,N_9804,N_9489);
nor U11662 (N_11662,N_9131,N_9523);
or U11663 (N_11663,N_10339,N_9780);
xor U11664 (N_11664,N_9027,N_9494);
and U11665 (N_11665,N_9706,N_10240);
or U11666 (N_11666,N_9865,N_9449);
and U11667 (N_11667,N_9050,N_9087);
xnor U11668 (N_11668,N_9545,N_9681);
nand U11669 (N_11669,N_9197,N_9121);
or U11670 (N_11670,N_9991,N_9742);
or U11671 (N_11671,N_10373,N_9362);
xor U11672 (N_11672,N_10354,N_10446);
xnor U11673 (N_11673,N_10121,N_9452);
xor U11674 (N_11674,N_10368,N_9623);
nand U11675 (N_11675,N_10150,N_9570);
or U11676 (N_11676,N_9784,N_9418);
or U11677 (N_11677,N_9723,N_10012);
and U11678 (N_11678,N_9126,N_9835);
or U11679 (N_11679,N_10398,N_10181);
nor U11680 (N_11680,N_9309,N_10481);
nor U11681 (N_11681,N_9797,N_10029);
and U11682 (N_11682,N_10012,N_10390);
xnor U11683 (N_11683,N_10160,N_9991);
nand U11684 (N_11684,N_9623,N_9339);
nor U11685 (N_11685,N_9470,N_9665);
nand U11686 (N_11686,N_9947,N_9682);
and U11687 (N_11687,N_10471,N_9791);
and U11688 (N_11688,N_9871,N_9620);
nor U11689 (N_11689,N_9939,N_9142);
xor U11690 (N_11690,N_9702,N_9347);
nand U11691 (N_11691,N_10146,N_10235);
xnor U11692 (N_11692,N_9983,N_9996);
or U11693 (N_11693,N_10311,N_9565);
and U11694 (N_11694,N_9491,N_10291);
or U11695 (N_11695,N_9863,N_10213);
or U11696 (N_11696,N_9455,N_9537);
nand U11697 (N_11697,N_10099,N_10349);
nor U11698 (N_11698,N_10457,N_10485);
nor U11699 (N_11699,N_9052,N_10342);
or U11700 (N_11700,N_10294,N_9478);
and U11701 (N_11701,N_9898,N_9986);
xor U11702 (N_11702,N_10109,N_9945);
nor U11703 (N_11703,N_9728,N_10231);
nand U11704 (N_11704,N_9319,N_9611);
nor U11705 (N_11705,N_9039,N_9399);
nor U11706 (N_11706,N_10210,N_9201);
xor U11707 (N_11707,N_9208,N_9469);
and U11708 (N_11708,N_9631,N_9564);
xnor U11709 (N_11709,N_9329,N_9518);
and U11710 (N_11710,N_9800,N_10015);
nand U11711 (N_11711,N_9241,N_9834);
or U11712 (N_11712,N_9398,N_9627);
or U11713 (N_11713,N_9737,N_9300);
nand U11714 (N_11714,N_9181,N_9517);
nor U11715 (N_11715,N_9534,N_9348);
or U11716 (N_11716,N_9420,N_10105);
nand U11717 (N_11717,N_9508,N_9685);
nand U11718 (N_11718,N_10075,N_10422);
or U11719 (N_11719,N_9008,N_10172);
nand U11720 (N_11720,N_10219,N_9799);
and U11721 (N_11721,N_9149,N_9738);
nor U11722 (N_11722,N_9990,N_9371);
nand U11723 (N_11723,N_9409,N_9873);
xnor U11724 (N_11724,N_9312,N_9580);
or U11725 (N_11725,N_9723,N_9143);
nor U11726 (N_11726,N_10366,N_10091);
nand U11727 (N_11727,N_9621,N_9654);
or U11728 (N_11728,N_9581,N_10260);
and U11729 (N_11729,N_9244,N_10150);
nor U11730 (N_11730,N_10112,N_10079);
nor U11731 (N_11731,N_9463,N_9756);
xor U11732 (N_11732,N_9903,N_9672);
xnor U11733 (N_11733,N_10498,N_9236);
nand U11734 (N_11734,N_9987,N_9986);
nor U11735 (N_11735,N_9456,N_10060);
and U11736 (N_11736,N_9399,N_10040);
xnor U11737 (N_11737,N_10445,N_9709);
or U11738 (N_11738,N_10261,N_10421);
or U11739 (N_11739,N_10010,N_9480);
xor U11740 (N_11740,N_9751,N_9623);
and U11741 (N_11741,N_9889,N_10161);
nor U11742 (N_11742,N_10183,N_9341);
and U11743 (N_11743,N_9150,N_10270);
nand U11744 (N_11744,N_10011,N_9853);
nand U11745 (N_11745,N_9562,N_10152);
xnor U11746 (N_11746,N_10280,N_9550);
and U11747 (N_11747,N_10209,N_10059);
nand U11748 (N_11748,N_9658,N_9572);
nand U11749 (N_11749,N_10024,N_10017);
xnor U11750 (N_11750,N_9030,N_9398);
nand U11751 (N_11751,N_9762,N_9307);
nand U11752 (N_11752,N_10458,N_10051);
and U11753 (N_11753,N_9967,N_9182);
and U11754 (N_11754,N_9523,N_9661);
and U11755 (N_11755,N_9136,N_9889);
and U11756 (N_11756,N_10306,N_9866);
xnor U11757 (N_11757,N_9324,N_10369);
or U11758 (N_11758,N_9801,N_10207);
or U11759 (N_11759,N_9619,N_9826);
or U11760 (N_11760,N_10251,N_10173);
nand U11761 (N_11761,N_10124,N_10055);
xnor U11762 (N_11762,N_9797,N_9693);
nor U11763 (N_11763,N_10457,N_9658);
xnor U11764 (N_11764,N_9287,N_9882);
and U11765 (N_11765,N_10334,N_9461);
and U11766 (N_11766,N_10460,N_9112);
nand U11767 (N_11767,N_9951,N_10104);
xor U11768 (N_11768,N_9849,N_9046);
or U11769 (N_11769,N_9660,N_10114);
and U11770 (N_11770,N_9503,N_9405);
or U11771 (N_11771,N_9849,N_9168);
or U11772 (N_11772,N_10150,N_9887);
and U11773 (N_11773,N_10019,N_9288);
or U11774 (N_11774,N_9014,N_9092);
nor U11775 (N_11775,N_9202,N_9858);
or U11776 (N_11776,N_10477,N_10114);
nand U11777 (N_11777,N_9907,N_9736);
nand U11778 (N_11778,N_9143,N_9067);
xnor U11779 (N_11779,N_10313,N_9903);
and U11780 (N_11780,N_9427,N_9093);
nor U11781 (N_11781,N_10477,N_9310);
nand U11782 (N_11782,N_10143,N_10306);
nor U11783 (N_11783,N_9368,N_10267);
xor U11784 (N_11784,N_9692,N_9218);
nand U11785 (N_11785,N_9836,N_10363);
xor U11786 (N_11786,N_9928,N_9478);
or U11787 (N_11787,N_9709,N_10129);
and U11788 (N_11788,N_9134,N_10160);
and U11789 (N_11789,N_9301,N_10074);
or U11790 (N_11790,N_9538,N_10226);
nor U11791 (N_11791,N_9704,N_9821);
and U11792 (N_11792,N_10120,N_10186);
or U11793 (N_11793,N_9760,N_10296);
and U11794 (N_11794,N_9882,N_9325);
and U11795 (N_11795,N_10275,N_9514);
nor U11796 (N_11796,N_9288,N_10355);
nor U11797 (N_11797,N_9850,N_10188);
nor U11798 (N_11798,N_9448,N_9338);
xnor U11799 (N_11799,N_9569,N_9125);
nand U11800 (N_11800,N_10202,N_9700);
or U11801 (N_11801,N_9971,N_9198);
nor U11802 (N_11802,N_10253,N_10351);
xor U11803 (N_11803,N_10249,N_10095);
nand U11804 (N_11804,N_10497,N_9446);
xnor U11805 (N_11805,N_9039,N_10081);
nor U11806 (N_11806,N_9764,N_9936);
nor U11807 (N_11807,N_10293,N_10295);
or U11808 (N_11808,N_9211,N_9498);
xnor U11809 (N_11809,N_10238,N_10345);
nand U11810 (N_11810,N_10154,N_10350);
nor U11811 (N_11811,N_10025,N_9842);
nand U11812 (N_11812,N_9321,N_10487);
xnor U11813 (N_11813,N_9722,N_9584);
nand U11814 (N_11814,N_9133,N_10414);
or U11815 (N_11815,N_10220,N_9203);
xnor U11816 (N_11816,N_10431,N_9807);
nor U11817 (N_11817,N_9976,N_9997);
or U11818 (N_11818,N_10489,N_9640);
or U11819 (N_11819,N_9448,N_10136);
or U11820 (N_11820,N_9645,N_9372);
and U11821 (N_11821,N_10006,N_10498);
or U11822 (N_11822,N_9070,N_10469);
or U11823 (N_11823,N_9389,N_10195);
or U11824 (N_11824,N_9842,N_9349);
nand U11825 (N_11825,N_9515,N_9581);
xnor U11826 (N_11826,N_9347,N_9811);
nor U11827 (N_11827,N_9601,N_9630);
nand U11828 (N_11828,N_10213,N_10151);
xor U11829 (N_11829,N_10017,N_10190);
or U11830 (N_11830,N_9492,N_10343);
or U11831 (N_11831,N_9030,N_9713);
nand U11832 (N_11832,N_9295,N_9750);
and U11833 (N_11833,N_9785,N_9374);
or U11834 (N_11834,N_10220,N_9266);
xor U11835 (N_11835,N_9570,N_9197);
nand U11836 (N_11836,N_9676,N_10437);
nand U11837 (N_11837,N_10342,N_9288);
nand U11838 (N_11838,N_9287,N_10115);
nand U11839 (N_11839,N_9488,N_10163);
xnor U11840 (N_11840,N_9972,N_10085);
xor U11841 (N_11841,N_9952,N_9063);
xnor U11842 (N_11842,N_10423,N_9797);
nor U11843 (N_11843,N_10427,N_9594);
or U11844 (N_11844,N_9322,N_10043);
or U11845 (N_11845,N_10310,N_9909);
or U11846 (N_11846,N_9849,N_9590);
xnor U11847 (N_11847,N_10319,N_9679);
nand U11848 (N_11848,N_9059,N_9301);
nand U11849 (N_11849,N_9957,N_9203);
or U11850 (N_11850,N_10443,N_9144);
nor U11851 (N_11851,N_9175,N_9395);
xnor U11852 (N_11852,N_9965,N_9041);
nor U11853 (N_11853,N_9577,N_9933);
or U11854 (N_11854,N_9035,N_9023);
and U11855 (N_11855,N_9216,N_9594);
nor U11856 (N_11856,N_10164,N_10000);
and U11857 (N_11857,N_9455,N_9215);
nor U11858 (N_11858,N_9619,N_9383);
and U11859 (N_11859,N_9040,N_10185);
xnor U11860 (N_11860,N_10362,N_10023);
nand U11861 (N_11861,N_10427,N_9875);
and U11862 (N_11862,N_9184,N_9140);
xnor U11863 (N_11863,N_10140,N_9337);
nand U11864 (N_11864,N_9350,N_9817);
nor U11865 (N_11865,N_9009,N_9536);
or U11866 (N_11866,N_10264,N_10076);
xor U11867 (N_11867,N_10182,N_9070);
xnor U11868 (N_11868,N_9486,N_9290);
and U11869 (N_11869,N_9608,N_9946);
xnor U11870 (N_11870,N_9743,N_9918);
or U11871 (N_11871,N_10043,N_9662);
nor U11872 (N_11872,N_9646,N_9693);
xnor U11873 (N_11873,N_9465,N_9562);
and U11874 (N_11874,N_9406,N_9738);
nor U11875 (N_11875,N_9263,N_9951);
nand U11876 (N_11876,N_9831,N_10317);
or U11877 (N_11877,N_9133,N_9203);
nand U11878 (N_11878,N_10423,N_9997);
or U11879 (N_11879,N_9492,N_10292);
xor U11880 (N_11880,N_9658,N_10307);
and U11881 (N_11881,N_9493,N_9139);
xor U11882 (N_11882,N_10386,N_10346);
nor U11883 (N_11883,N_9757,N_10324);
xor U11884 (N_11884,N_10004,N_9140);
nand U11885 (N_11885,N_10332,N_9313);
nand U11886 (N_11886,N_9086,N_9732);
nor U11887 (N_11887,N_10293,N_10074);
nor U11888 (N_11888,N_9133,N_9560);
or U11889 (N_11889,N_9151,N_10035);
nand U11890 (N_11890,N_10226,N_10010);
or U11891 (N_11891,N_9246,N_9800);
and U11892 (N_11892,N_9444,N_10415);
xnor U11893 (N_11893,N_9728,N_9457);
nor U11894 (N_11894,N_10050,N_10182);
nand U11895 (N_11895,N_10266,N_9573);
xnor U11896 (N_11896,N_9005,N_10423);
and U11897 (N_11897,N_9825,N_10172);
nor U11898 (N_11898,N_9658,N_10180);
nand U11899 (N_11899,N_10321,N_10047);
nor U11900 (N_11900,N_9277,N_9026);
and U11901 (N_11901,N_9753,N_10170);
nand U11902 (N_11902,N_9995,N_9484);
nand U11903 (N_11903,N_9868,N_9724);
nor U11904 (N_11904,N_10201,N_9218);
nand U11905 (N_11905,N_9956,N_10343);
xnor U11906 (N_11906,N_10419,N_9722);
xnor U11907 (N_11907,N_10019,N_10108);
and U11908 (N_11908,N_9833,N_9285);
nand U11909 (N_11909,N_9491,N_9537);
xor U11910 (N_11910,N_9806,N_9162);
or U11911 (N_11911,N_9087,N_9600);
nor U11912 (N_11912,N_9266,N_9268);
and U11913 (N_11913,N_9627,N_9635);
or U11914 (N_11914,N_10054,N_9721);
nand U11915 (N_11915,N_9922,N_9468);
nor U11916 (N_11916,N_10452,N_10260);
nor U11917 (N_11917,N_10284,N_9844);
nor U11918 (N_11918,N_9581,N_9129);
nor U11919 (N_11919,N_9832,N_9638);
nand U11920 (N_11920,N_10441,N_9459);
nor U11921 (N_11921,N_9051,N_9936);
nor U11922 (N_11922,N_9788,N_9370);
or U11923 (N_11923,N_9947,N_9453);
and U11924 (N_11924,N_9516,N_10338);
xor U11925 (N_11925,N_9757,N_10224);
nor U11926 (N_11926,N_10353,N_9193);
nand U11927 (N_11927,N_9308,N_10266);
nand U11928 (N_11928,N_9885,N_10278);
or U11929 (N_11929,N_9768,N_10052);
or U11930 (N_11930,N_9364,N_9889);
and U11931 (N_11931,N_9581,N_10346);
and U11932 (N_11932,N_9768,N_9945);
nor U11933 (N_11933,N_10165,N_10317);
xor U11934 (N_11934,N_9489,N_9316);
xnor U11935 (N_11935,N_9861,N_10158);
or U11936 (N_11936,N_10437,N_9836);
and U11937 (N_11937,N_10362,N_10061);
nor U11938 (N_11938,N_10018,N_10475);
xor U11939 (N_11939,N_10421,N_10117);
xnor U11940 (N_11940,N_10231,N_10499);
and U11941 (N_11941,N_10347,N_9544);
and U11942 (N_11942,N_9384,N_9615);
nor U11943 (N_11943,N_9042,N_10139);
or U11944 (N_11944,N_9768,N_10375);
or U11945 (N_11945,N_9258,N_10147);
or U11946 (N_11946,N_9588,N_9021);
nand U11947 (N_11947,N_9637,N_9977);
nor U11948 (N_11948,N_10302,N_9146);
xnor U11949 (N_11949,N_9647,N_10081);
nor U11950 (N_11950,N_10070,N_9171);
and U11951 (N_11951,N_9437,N_9309);
nor U11952 (N_11952,N_9218,N_9492);
and U11953 (N_11953,N_10394,N_9299);
or U11954 (N_11954,N_10148,N_9595);
and U11955 (N_11955,N_10157,N_10114);
and U11956 (N_11956,N_9015,N_9098);
nand U11957 (N_11957,N_9334,N_9085);
xnor U11958 (N_11958,N_9444,N_10496);
nand U11959 (N_11959,N_10069,N_9602);
nand U11960 (N_11960,N_9106,N_10165);
or U11961 (N_11961,N_10293,N_10061);
or U11962 (N_11962,N_9955,N_10174);
nor U11963 (N_11963,N_9238,N_9012);
xnor U11964 (N_11964,N_9373,N_10044);
nand U11965 (N_11965,N_9367,N_9385);
or U11966 (N_11966,N_9730,N_10373);
nor U11967 (N_11967,N_9288,N_9455);
or U11968 (N_11968,N_9015,N_9836);
xor U11969 (N_11969,N_9435,N_10220);
or U11970 (N_11970,N_10185,N_10383);
and U11971 (N_11971,N_10006,N_9353);
or U11972 (N_11972,N_10306,N_9343);
nor U11973 (N_11973,N_10183,N_9231);
xor U11974 (N_11974,N_10013,N_9182);
or U11975 (N_11975,N_9592,N_9812);
xnor U11976 (N_11976,N_9787,N_9365);
xor U11977 (N_11977,N_9239,N_9782);
or U11978 (N_11978,N_9054,N_9535);
or U11979 (N_11979,N_10254,N_10171);
nor U11980 (N_11980,N_9994,N_10346);
nor U11981 (N_11981,N_9784,N_10425);
nand U11982 (N_11982,N_9676,N_9452);
and U11983 (N_11983,N_10486,N_9551);
or U11984 (N_11984,N_10147,N_9861);
or U11985 (N_11985,N_9222,N_10389);
and U11986 (N_11986,N_10210,N_9932);
nand U11987 (N_11987,N_9521,N_9031);
nand U11988 (N_11988,N_9862,N_10287);
xor U11989 (N_11989,N_10159,N_9267);
or U11990 (N_11990,N_9697,N_10214);
nand U11991 (N_11991,N_9194,N_9933);
or U11992 (N_11992,N_9088,N_9280);
nor U11993 (N_11993,N_9451,N_9508);
and U11994 (N_11994,N_10279,N_9951);
or U11995 (N_11995,N_9941,N_9105);
and U11996 (N_11996,N_9321,N_9978);
nand U11997 (N_11997,N_9134,N_10196);
or U11998 (N_11998,N_9845,N_10216);
or U11999 (N_11999,N_9905,N_9652);
and U12000 (N_12000,N_10785,N_11378);
xor U12001 (N_12001,N_10654,N_11614);
nand U12002 (N_12002,N_10902,N_10598);
or U12003 (N_12003,N_11600,N_10587);
or U12004 (N_12004,N_10814,N_11247);
or U12005 (N_12005,N_10683,N_11363);
nor U12006 (N_12006,N_10991,N_10925);
nor U12007 (N_12007,N_10512,N_11842);
or U12008 (N_12008,N_11664,N_10866);
and U12009 (N_12009,N_11811,N_10642);
nand U12010 (N_12010,N_11311,N_10890);
xor U12011 (N_12011,N_10873,N_11776);
xor U12012 (N_12012,N_11018,N_11075);
and U12013 (N_12013,N_10623,N_11472);
nand U12014 (N_12014,N_11610,N_11398);
nand U12015 (N_12015,N_11772,N_11318);
xor U12016 (N_12016,N_10947,N_10561);
nor U12017 (N_12017,N_10787,N_11441);
xor U12018 (N_12018,N_10772,N_11178);
xor U12019 (N_12019,N_10593,N_10580);
and U12020 (N_12020,N_11386,N_10556);
and U12021 (N_12021,N_11846,N_11701);
and U12022 (N_12022,N_10907,N_11929);
nand U12023 (N_12023,N_11790,N_10673);
or U12024 (N_12024,N_11146,N_11115);
nand U12025 (N_12025,N_10732,N_10637);
and U12026 (N_12026,N_11061,N_11280);
xnor U12027 (N_12027,N_11332,N_11888);
xor U12028 (N_12028,N_11496,N_11465);
and U12029 (N_12029,N_11934,N_11053);
and U12030 (N_12030,N_11968,N_10663);
or U12031 (N_12031,N_11380,N_11905);
xnor U12032 (N_12032,N_11414,N_11913);
xor U12033 (N_12033,N_11249,N_11365);
and U12034 (N_12034,N_11826,N_11911);
and U12035 (N_12035,N_11523,N_11252);
xor U12036 (N_12036,N_11016,N_11397);
xnor U12037 (N_12037,N_11302,N_11801);
nor U12038 (N_12038,N_11983,N_10900);
xnor U12039 (N_12039,N_10685,N_10942);
nand U12040 (N_12040,N_10562,N_10566);
nor U12041 (N_12041,N_11855,N_11727);
or U12042 (N_12042,N_10851,N_10993);
and U12043 (N_12043,N_11008,N_11305);
and U12044 (N_12044,N_11840,N_11338);
xnor U12045 (N_12045,N_11341,N_10628);
nor U12046 (N_12046,N_10624,N_11513);
nand U12047 (N_12047,N_11782,N_11735);
or U12048 (N_12048,N_11781,N_11731);
nand U12049 (N_12049,N_11323,N_11538);
or U12050 (N_12050,N_10727,N_10794);
or U12051 (N_12051,N_11005,N_11350);
and U12052 (N_12052,N_10974,N_10763);
or U12053 (N_12053,N_10889,N_11742);
and U12054 (N_12054,N_11308,N_11946);
or U12055 (N_12055,N_10746,N_11549);
nand U12056 (N_12056,N_11462,N_11299);
or U12057 (N_12057,N_11029,N_11509);
nand U12058 (N_12058,N_11474,N_11721);
nor U12059 (N_12059,N_11133,N_11389);
xor U12060 (N_12060,N_11738,N_11999);
and U12061 (N_12061,N_11981,N_11090);
or U12062 (N_12062,N_11932,N_10741);
nor U12063 (N_12063,N_11966,N_11511);
and U12064 (N_12064,N_11073,N_10842);
nand U12065 (N_12065,N_11851,N_11637);
nor U12066 (N_12066,N_11896,N_10548);
xnor U12067 (N_12067,N_11704,N_11835);
nor U12068 (N_12068,N_11942,N_10543);
or U12069 (N_12069,N_10844,N_11223);
nor U12070 (N_12070,N_10857,N_11215);
and U12071 (N_12071,N_10575,N_11428);
or U12072 (N_12072,N_11202,N_10809);
nor U12073 (N_12073,N_11762,N_11454);
xor U12074 (N_12074,N_11181,N_11271);
xnor U12075 (N_12075,N_11489,N_11371);
and U12076 (N_12076,N_10606,N_10953);
or U12077 (N_12077,N_11931,N_11793);
xor U12078 (N_12078,N_10714,N_10766);
nand U12079 (N_12079,N_10748,N_10643);
nand U12080 (N_12080,N_10616,N_11900);
nor U12081 (N_12081,N_11477,N_11922);
and U12082 (N_12082,N_11370,N_10992);
or U12083 (N_12083,N_11971,N_10863);
xor U12084 (N_12084,N_11187,N_11996);
nor U12085 (N_12085,N_11829,N_10754);
xnor U12086 (N_12086,N_10538,N_11147);
xor U12087 (N_12087,N_11125,N_10705);
nor U12088 (N_12088,N_11697,N_11961);
and U12089 (N_12089,N_11765,N_11965);
and U12090 (N_12090,N_11006,N_10681);
nand U12091 (N_12091,N_11953,N_11225);
xor U12092 (N_12092,N_11036,N_11186);
xnor U12093 (N_12093,N_11325,N_11702);
nand U12094 (N_12094,N_11194,N_11530);
nor U12095 (N_12095,N_11915,N_11410);
xnor U12096 (N_12096,N_10796,N_10817);
nand U12097 (N_12097,N_10740,N_11486);
and U12098 (N_12098,N_10718,N_10771);
nand U12099 (N_12099,N_10911,N_11060);
xor U12100 (N_12100,N_10668,N_10504);
and U12101 (N_12101,N_10567,N_11122);
xnor U12102 (N_12102,N_10941,N_11129);
nor U12103 (N_12103,N_10508,N_11969);
and U12104 (N_12104,N_10525,N_11789);
nor U12105 (N_12105,N_11967,N_11403);
or U12106 (N_12106,N_11169,N_10865);
and U12107 (N_12107,N_10872,N_10854);
nand U12108 (N_12108,N_11524,N_10610);
or U12109 (N_12109,N_11645,N_11933);
xnor U12110 (N_12110,N_11027,N_10896);
nand U12111 (N_12111,N_10965,N_11049);
and U12112 (N_12112,N_10584,N_10664);
and U12113 (N_12113,N_11559,N_11611);
nor U12114 (N_12114,N_10943,N_11110);
and U12115 (N_12115,N_10996,N_11992);
nor U12116 (N_12116,N_10641,N_11551);
nand U12117 (N_12117,N_11213,N_11691);
nor U12118 (N_12118,N_11886,N_11553);
and U12119 (N_12119,N_11291,N_11510);
or U12120 (N_12120,N_10666,N_10577);
or U12121 (N_12121,N_10530,N_11642);
or U12122 (N_12122,N_10722,N_11847);
or U12123 (N_12123,N_11392,N_10743);
xor U12124 (N_12124,N_11381,N_10975);
nor U12125 (N_12125,N_10927,N_11505);
or U12126 (N_12126,N_11051,N_11670);
nor U12127 (N_12127,N_10630,N_11345);
and U12128 (N_12128,N_11884,N_10679);
or U12129 (N_12129,N_11984,N_11035);
nand U12130 (N_12130,N_10523,N_11165);
nor U12131 (N_12131,N_10858,N_11173);
nor U12132 (N_12132,N_10632,N_11991);
nor U12133 (N_12133,N_10946,N_11809);
xnor U12134 (N_12134,N_11460,N_11166);
nand U12135 (N_12135,N_10536,N_11248);
nand U12136 (N_12136,N_11543,N_11787);
xor U12137 (N_12137,N_11607,N_11872);
xnor U12138 (N_12138,N_11909,N_11042);
nand U12139 (N_12139,N_11820,N_11621);
or U12140 (N_12140,N_10825,N_10886);
and U12141 (N_12141,N_10834,N_11232);
xor U12142 (N_12142,N_11055,N_11279);
xnor U12143 (N_12143,N_10997,N_10861);
and U12144 (N_12144,N_11815,N_11679);
or U12145 (N_12145,N_11072,N_10841);
nand U12146 (N_12146,N_11724,N_11528);
and U12147 (N_12147,N_11723,N_11502);
xnor U12148 (N_12148,N_11092,N_11405);
nand U12149 (N_12149,N_10960,N_11425);
or U12150 (N_12150,N_11023,N_11944);
nand U12151 (N_12151,N_11373,N_10573);
nand U12152 (N_12152,N_11164,N_10651);
nor U12153 (N_12153,N_10591,N_11424);
xnor U12154 (N_12154,N_10962,N_11429);
xnor U12155 (N_12155,N_10609,N_10867);
or U12156 (N_12156,N_11268,N_10912);
nand U12157 (N_12157,N_10777,N_11960);
or U12158 (N_12158,N_11764,N_11245);
and U12159 (N_12159,N_10586,N_11868);
nand U12160 (N_12160,N_11666,N_10626);
and U12161 (N_12161,N_11289,N_10999);
xor U12162 (N_12162,N_11858,N_11678);
nand U12163 (N_12163,N_11955,N_10830);
xnor U12164 (N_12164,N_10773,N_10676);
nor U12165 (N_12165,N_11040,N_11880);
nand U12166 (N_12166,N_11567,N_11116);
and U12167 (N_12167,N_11628,N_11198);
xnor U12168 (N_12168,N_11824,N_11834);
and U12169 (N_12169,N_11574,N_11962);
and U12170 (N_12170,N_11217,N_11879);
nand U12171 (N_12171,N_11587,N_11032);
nand U12172 (N_12172,N_10747,N_11033);
nor U12173 (N_12173,N_10551,N_10607);
or U12174 (N_12174,N_11799,N_10824);
xnor U12175 (N_12175,N_11438,N_10533);
xnor U12176 (N_12176,N_11748,N_10839);
xor U12177 (N_12177,N_10933,N_10919);
xor U12178 (N_12178,N_11914,N_10932);
and U12179 (N_12179,N_11171,N_10513);
and U12180 (N_12180,N_11746,N_11798);
xnor U12181 (N_12181,N_10786,N_11185);
nor U12182 (N_12182,N_11100,N_11810);
or U12183 (N_12183,N_11716,N_10726);
xor U12184 (N_12184,N_10876,N_11596);
or U12185 (N_12185,N_10819,N_10614);
nand U12186 (N_12186,N_10686,N_11416);
nor U12187 (N_12187,N_10646,N_10874);
xor U12188 (N_12188,N_11466,N_10967);
nor U12189 (N_12189,N_11493,N_11795);
nand U12190 (N_12190,N_11277,N_10915);
nor U12191 (N_12191,N_11584,N_11594);
nand U12192 (N_12192,N_11191,N_11867);
or U12193 (N_12193,N_11558,N_10524);
nor U12194 (N_12194,N_10675,N_11206);
or U12195 (N_12195,N_11265,N_10955);
xor U12196 (N_12196,N_10592,N_10784);
or U12197 (N_12197,N_11836,N_11025);
xnor U12198 (N_12198,N_11803,N_11703);
nand U12199 (N_12199,N_11572,N_11830);
nor U12200 (N_12200,N_10680,N_11445);
nor U12201 (N_12201,N_11891,N_11095);
or U12202 (N_12202,N_11887,N_10826);
nor U12203 (N_12203,N_11504,N_11862);
xor U12204 (N_12204,N_11327,N_11714);
nand U12205 (N_12205,N_11705,N_11157);
and U12206 (N_12206,N_10723,N_11358);
or U12207 (N_12207,N_11333,N_11168);
and U12208 (N_12208,N_11593,N_11402);
nand U12209 (N_12209,N_11203,N_11156);
and U12210 (N_12210,N_11937,N_11952);
nand U12211 (N_12211,N_11713,N_10547);
nand U12212 (N_12212,N_11537,N_10944);
and U12213 (N_12213,N_11155,N_11526);
or U12214 (N_12214,N_11238,N_11508);
xor U12215 (N_12215,N_11595,N_11521);
or U12216 (N_12216,N_10696,N_11000);
nand U12217 (N_12217,N_11082,N_11417);
or U12218 (N_12218,N_10712,N_11087);
or U12219 (N_12219,N_11658,N_10698);
or U12220 (N_12220,N_11687,N_11009);
xor U12221 (N_12221,N_11451,N_10621);
nand U12222 (N_12222,N_11631,N_11089);
or U12223 (N_12223,N_11737,N_10897);
or U12224 (N_12224,N_10936,N_11176);
or U12225 (N_12225,N_10620,N_10979);
nand U12226 (N_12226,N_11512,N_10868);
nor U12227 (N_12227,N_11336,N_11885);
xnor U12228 (N_12228,N_10719,N_11833);
and U12229 (N_12229,N_10811,N_11604);
xor U12230 (N_12230,N_11818,N_10550);
or U12231 (N_12231,N_10542,N_11151);
xor U12232 (N_12232,N_11069,N_11956);
or U12233 (N_12233,N_11276,N_11076);
xor U12234 (N_12234,N_10973,N_10658);
xor U12235 (N_12235,N_10831,N_10820);
xor U12236 (N_12236,N_11749,N_10769);
nand U12237 (N_12237,N_11272,N_11629);
and U12238 (N_12238,N_10849,N_11605);
nand U12239 (N_12239,N_10644,N_10846);
xnor U12240 (N_12240,N_10682,N_11845);
nand U12241 (N_12241,N_10708,N_11640);
nor U12242 (N_12242,N_10667,N_10564);
and U12243 (N_12243,N_11406,N_11004);
nor U12244 (N_12244,N_10730,N_10576);
xnor U12245 (N_12245,N_11831,N_11419);
nand U12246 (N_12246,N_11665,N_10959);
and U12247 (N_12247,N_10869,N_11501);
xnor U12248 (N_12248,N_11487,N_10724);
or U12249 (N_12249,N_11792,N_11753);
or U12250 (N_12250,N_11093,N_11431);
and U12251 (N_12251,N_11024,N_11145);
nand U12252 (N_12252,N_10793,N_11759);
xnor U12253 (N_12253,N_11368,N_11432);
xor U12254 (N_12254,N_11662,N_11037);
and U12255 (N_12255,N_11893,N_11261);
and U12256 (N_12256,N_10828,N_11693);
nor U12257 (N_12257,N_10559,N_11455);
nor U12258 (N_12258,N_11927,N_11152);
nor U12259 (N_12259,N_11812,N_10950);
nand U12260 (N_12260,N_11492,N_11676);
xnor U12261 (N_12261,N_10703,N_11266);
xor U12262 (N_12262,N_10790,N_11415);
nand U12263 (N_12263,N_11582,N_10758);
or U12264 (N_12264,N_10905,N_11695);
or U12265 (N_12265,N_10986,N_11189);
or U12266 (N_12266,N_11190,N_10653);
or U12267 (N_12267,N_11433,N_11334);
nor U12268 (N_12268,N_10717,N_11517);
nand U12269 (N_12269,N_11550,N_10937);
and U12270 (N_12270,N_10760,N_11104);
and U12271 (N_12271,N_10870,N_11344);
nand U12272 (N_12272,N_11136,N_11747);
xor U12273 (N_12273,N_11010,N_10994);
xor U12274 (N_12274,N_11571,N_10835);
nor U12275 (N_12275,N_11850,N_11852);
or U12276 (N_12276,N_10563,N_11453);
or U12277 (N_12277,N_10805,N_11434);
xor U12278 (N_12278,N_10534,N_10840);
and U12279 (N_12279,N_11297,N_10880);
and U12280 (N_12280,N_11774,N_10509);
nand U12281 (N_12281,N_11064,N_10829);
xnor U12282 (N_12282,N_11907,N_10898);
xor U12283 (N_12283,N_11457,N_11897);
or U12284 (N_12284,N_11177,N_11507);
nand U12285 (N_12285,N_11728,N_11158);
and U12286 (N_12286,N_10529,N_11692);
xor U12287 (N_12287,N_11007,N_11356);
nor U12288 (N_12288,N_10594,N_11951);
or U12289 (N_12289,N_11566,N_11207);
xor U12290 (N_12290,N_11963,N_11870);
nor U12291 (N_12291,N_11167,N_11118);
nor U12292 (N_12292,N_11026,N_10710);
xor U12293 (N_12293,N_10948,N_11562);
or U12294 (N_12294,N_11889,N_10600);
xnor U12295 (N_12295,N_10971,N_11674);
or U12296 (N_12296,N_10906,N_11542);
xor U12297 (N_12297,N_11160,N_11581);
xor U12298 (N_12298,N_10501,N_11615);
nor U12299 (N_12299,N_11123,N_10978);
and U12300 (N_12300,N_10583,N_10983);
and U12301 (N_12301,N_11257,N_11794);
and U12302 (N_12302,N_10541,N_11226);
nor U12303 (N_12303,N_11828,N_11844);
and U12304 (N_12304,N_11015,N_11339);
nand U12305 (N_12305,N_11390,N_11763);
or U12306 (N_12306,N_11618,N_11337);
xnor U12307 (N_12307,N_11654,N_11319);
and U12308 (N_12308,N_11838,N_11921);
nand U12309 (N_12309,N_10735,N_11802);
nand U12310 (N_12310,N_10510,N_11568);
and U12311 (N_12311,N_11387,N_11564);
and U12312 (N_12312,N_11488,N_11456);
or U12313 (N_12313,N_11459,N_11686);
nor U12314 (N_12314,N_11011,N_11139);
or U12315 (N_12315,N_11943,N_11324);
and U12316 (N_12316,N_11575,N_11876);
xor U12317 (N_12317,N_10980,N_11912);
nor U12318 (N_12318,N_10531,N_11430);
xor U12319 (N_12319,N_10875,N_11668);
or U12320 (N_12320,N_11395,N_11320);
nor U12321 (N_12321,N_11780,N_10818);
xor U12322 (N_12322,N_11864,N_11503);
nand U12323 (N_12323,N_10633,N_11988);
xnor U12324 (N_12324,N_11925,N_11755);
or U12325 (N_12325,N_11813,N_10882);
xor U12326 (N_12326,N_11903,N_11673);
nand U12327 (N_12327,N_11047,N_11105);
nand U12328 (N_12328,N_11583,N_11340);
nand U12329 (N_12329,N_11698,N_11126);
xnor U12330 (N_12330,N_10806,N_10952);
or U12331 (N_12331,N_10837,N_10969);
and U12332 (N_12332,N_11899,N_10612);
nand U12333 (N_12333,N_10742,N_10888);
or U12334 (N_12334,N_11119,N_10926);
xnor U12335 (N_12335,N_10568,N_11985);
or U12336 (N_12336,N_11262,N_11527);
and U12337 (N_12337,N_11290,N_11957);
xor U12338 (N_12338,N_11439,N_11014);
and U12339 (N_12339,N_11726,N_11643);
nor U12340 (N_12340,N_10764,N_10711);
nor U12341 (N_12341,N_11468,N_10690);
nor U12342 (N_12342,N_10756,N_10549);
and U12343 (N_12343,N_11536,N_11366);
xor U12344 (N_12344,N_11841,N_11304);
nor U12345 (N_12345,N_11141,N_11849);
xor U12346 (N_12346,N_10701,N_10776);
xnor U12347 (N_12347,N_11860,N_10921);
nand U12348 (N_12348,N_11744,N_10914);
nand U12349 (N_12349,N_10982,N_11709);
or U12350 (N_12350,N_10923,N_11739);
xnor U12351 (N_12351,N_11200,N_11906);
nor U12352 (N_12352,N_10877,N_11067);
nand U12353 (N_12353,N_11352,N_11919);
nor U12354 (N_12354,N_11039,N_11883);
xnor U12355 (N_12355,N_11633,N_11625);
xor U12356 (N_12356,N_11938,N_11783);
nand U12357 (N_12357,N_10761,N_10908);
xnor U12358 (N_12358,N_11875,N_11470);
or U12359 (N_12359,N_11140,N_11646);
and U12360 (N_12360,N_11132,N_11396);
and U12361 (N_12361,N_11636,N_11585);
and U12362 (N_12362,N_10954,N_10636);
and U12363 (N_12363,N_11210,N_11547);
and U12364 (N_12364,N_11056,N_11978);
xnor U12365 (N_12365,N_10739,N_11315);
nand U12366 (N_12366,N_11597,N_11295);
or U12367 (N_12367,N_11800,N_10845);
or U12368 (N_12368,N_11443,N_11760);
and U12369 (N_12369,N_11233,N_11231);
nand U12370 (N_12370,N_11535,N_11446);
and U12371 (N_12371,N_11590,N_11557);
or U12372 (N_12372,N_10572,N_11260);
and U12373 (N_12373,N_10611,N_11275);
or U12374 (N_12374,N_11606,N_11522);
or U12375 (N_12375,N_11577,N_11554);
and U12376 (N_12376,N_11580,N_11103);
and U12377 (N_12377,N_10693,N_11630);
or U12378 (N_12378,N_11684,N_11661);
and U12379 (N_12379,N_11993,N_11690);
and U12380 (N_12380,N_11719,N_11881);
or U12381 (N_12381,N_10765,N_11284);
xor U12382 (N_12382,N_11068,N_10970);
nand U12383 (N_12383,N_11329,N_10627);
or U12384 (N_12384,N_10687,N_11250);
nand U12385 (N_12385,N_10972,N_11349);
nor U12386 (N_12386,N_11939,N_11134);
nand U12387 (N_12387,N_11017,N_11873);
nand U12388 (N_12388,N_11591,N_10887);
or U12389 (N_12389,N_10571,N_11494);
nor U12390 (N_12390,N_10847,N_10601);
or U12391 (N_12391,N_11030,N_11948);
xnor U12392 (N_12392,N_10848,N_10884);
xnor U12393 (N_12393,N_11979,N_11808);
or U12394 (N_12394,N_11987,N_10535);
nor U12395 (N_12395,N_11372,N_11256);
xnor U12396 (N_12396,N_10622,N_11699);
nor U12397 (N_12397,N_10506,N_11239);
nand U12398 (N_12398,N_11696,N_11548);
xnor U12399 (N_12399,N_11361,N_11720);
nor U12400 (N_12400,N_10913,N_10958);
and U12401 (N_12401,N_11570,N_11436);
nor U12402 (N_12402,N_10555,N_11561);
and U12403 (N_12403,N_11639,N_11193);
or U12404 (N_12404,N_10949,N_11563);
nor U12405 (N_12405,N_10904,N_11375);
nand U12406 (N_12406,N_11806,N_11940);
or U12407 (N_12407,N_11052,N_11998);
or U12408 (N_12408,N_11479,N_10545);
nor U12409 (N_12409,N_11651,N_11400);
xnor U12410 (N_12410,N_11990,N_10581);
nor U12411 (N_12411,N_10895,N_11667);
and U12412 (N_12412,N_10985,N_10843);
nand U12413 (N_12413,N_11255,N_11612);
and U12414 (N_12414,N_11745,N_11081);
and U12415 (N_12415,N_10578,N_10729);
or U12416 (N_12416,N_11314,N_10516);
xor U12417 (N_12417,N_10780,N_11317);
and U12418 (N_12418,N_11222,N_11074);
or U12419 (N_12419,N_11211,N_11552);
nand U12420 (N_12420,N_11094,N_10546);
nor U12421 (N_12421,N_11143,N_11994);
nand U12422 (N_12422,N_10517,N_11234);
xnor U12423 (N_12423,N_11229,N_11878);
or U12424 (N_12424,N_11857,N_10521);
and U12425 (N_12425,N_11058,N_11458);
nand U12426 (N_12426,N_11775,N_10862);
nand U12427 (N_12427,N_10599,N_11534);
nor U12428 (N_12428,N_10779,N_11022);
xnor U12429 (N_12429,N_11253,N_11989);
and U12430 (N_12430,N_10565,N_10990);
nor U12431 (N_12431,N_11469,N_11863);
and U12432 (N_12432,N_11916,N_10553);
nor U12433 (N_12433,N_11149,N_11672);
nor U12434 (N_12434,N_11895,N_11449);
xor U12435 (N_12435,N_10963,N_10588);
or U12436 (N_12436,N_10755,N_11218);
nand U12437 (N_12437,N_11278,N_11224);
nand U12438 (N_12438,N_10639,N_11038);
and U12439 (N_12439,N_11054,N_11769);
xnor U12440 (N_12440,N_11099,N_11463);
nand U12441 (N_12441,N_11997,N_11917);
nand U12442 (N_12442,N_11740,N_11354);
nand U12443 (N_12443,N_10838,N_11285);
and U12444 (N_12444,N_10881,N_11388);
or U12445 (N_12445,N_10816,N_11346);
nand U12446 (N_12446,N_11142,N_10655);
nor U12447 (N_12447,N_10570,N_10995);
xor U12448 (N_12448,N_10532,N_11565);
or U12449 (N_12449,N_10976,N_11683);
nor U12450 (N_12450,N_10928,N_11601);
and U12451 (N_12451,N_11694,N_11411);
or U12452 (N_12452,N_11865,N_10715);
nor U12453 (N_12453,N_11677,N_11221);
or U12454 (N_12454,N_10605,N_11288);
nand U12455 (N_12455,N_11652,N_10706);
and U12456 (N_12456,N_11079,N_11188);
nor U12457 (N_12457,N_10656,N_11404);
nor U12458 (N_12458,N_11130,N_10956);
xnor U12459 (N_12459,N_10585,N_10770);
xor U12460 (N_12460,N_11588,N_10892);
and U12461 (N_12461,N_10752,N_11205);
or U12462 (N_12462,N_10514,N_11569);
nand U12463 (N_12463,N_11786,N_11822);
and U12464 (N_12464,N_10799,N_11954);
or U12465 (N_12465,N_10757,N_10702);
nor U12466 (N_12466,N_10659,N_11263);
nor U12467 (N_12467,N_10540,N_11958);
xnor U12468 (N_12468,N_11347,N_11062);
and U12469 (N_12469,N_11482,N_11586);
or U12470 (N_12470,N_11418,N_10855);
xor U12471 (N_12471,N_11741,N_10853);
nor U12472 (N_12472,N_10528,N_11296);
nand U12473 (N_12473,N_11484,N_11201);
xnor U12474 (N_12474,N_11498,N_11773);
nor U12475 (N_12475,N_11663,N_11532);
and U12476 (N_12476,N_11420,N_11766);
nor U12477 (N_12477,N_11080,N_10823);
nand U12478 (N_12478,N_11096,N_11480);
or U12479 (N_12479,N_10694,N_11473);
and U12480 (N_12480,N_10836,N_11982);
nand U12481 (N_12481,N_11241,N_11950);
and U12482 (N_12482,N_11768,N_11127);
nor U12483 (N_12483,N_11385,N_10697);
nor U12484 (N_12484,N_11084,N_11920);
nand U12485 (N_12485,N_11031,N_11028);
nand U12486 (N_12486,N_11973,N_10939);
or U12487 (N_12487,N_11335,N_10684);
nand U12488 (N_12488,N_10792,N_10984);
nor U12489 (N_12489,N_11689,N_11926);
and U12490 (N_12490,N_11578,N_11274);
nand U12491 (N_12491,N_10822,N_10803);
nor U12492 (N_12492,N_11376,N_11722);
nand U12493 (N_12493,N_10856,N_11182);
nor U12494 (N_12494,N_10768,N_10751);
or U12495 (N_12495,N_11227,N_11246);
nor U12496 (N_12496,N_10629,N_11779);
xnor U12497 (N_12497,N_11121,N_10966);
or U12498 (N_12498,N_11001,N_10734);
and U12499 (N_12499,N_11540,N_11150);
nor U12500 (N_12500,N_11321,N_11882);
xor U12501 (N_12501,N_11598,N_11506);
xor U12502 (N_12502,N_11180,N_11359);
nand U12503 (N_12503,N_10917,N_10569);
nand U12504 (N_12504,N_11048,N_11854);
or U12505 (N_12505,N_10736,N_10775);
nand U12506 (N_12506,N_11467,N_10511);
xor U12507 (N_12507,N_10850,N_11447);
nor U12508 (N_12508,N_11219,N_11367);
xnor U12509 (N_12509,N_11959,N_11647);
xnor U12510 (N_12510,N_10910,N_10597);
or U12511 (N_12511,N_11947,N_11623);
or U12512 (N_12512,N_10977,N_11240);
and U12513 (N_12513,N_11326,N_10859);
nand U12514 (N_12514,N_10692,N_10579);
xnor U12515 (N_12515,N_11251,N_10810);
or U12516 (N_12516,N_11409,N_11065);
xnor U12517 (N_12517,N_11382,N_11653);
and U12518 (N_12518,N_10934,N_11708);
nor U12519 (N_12519,N_11819,N_11413);
nand U12520 (N_12520,N_10798,N_11301);
nand U12521 (N_12521,N_11374,N_10893);
xor U12522 (N_12522,N_11977,N_10801);
and U12523 (N_12523,N_11148,N_11097);
or U12524 (N_12524,N_10631,N_10725);
nand U12525 (N_12525,N_11330,N_10713);
nand U12526 (N_12526,N_11821,N_11945);
nand U12527 (N_12527,N_11717,N_10901);
nand U12528 (N_12528,N_10922,N_10608);
or U12529 (N_12529,N_11519,N_10669);
xor U12530 (N_12530,N_11784,N_11242);
or U12531 (N_12531,N_10670,N_11649);
nand U12532 (N_12532,N_11012,N_11609);
xnor U12533 (N_12533,N_10527,N_11294);
xnor U12534 (N_12534,N_11412,N_11660);
or U12535 (N_12535,N_11273,N_11270);
xnor U12536 (N_12536,N_11791,N_11603);
nand U12537 (N_12537,N_11675,N_11310);
xor U12538 (N_12538,N_10645,N_10981);
nor U12539 (N_12539,N_11102,N_11733);
or U12540 (N_12540,N_10744,N_11706);
xnor U12541 (N_12541,N_10700,N_11805);
nor U12542 (N_12542,N_10699,N_11877);
nor U12543 (N_12543,N_10558,N_10903);
xor U12544 (N_12544,N_10852,N_11485);
or U12545 (N_12545,N_11286,N_11797);
xor U12546 (N_12546,N_10957,N_10619);
or U12547 (N_12547,N_11101,N_10728);
nand U12548 (N_12548,N_11539,N_11109);
xor U12549 (N_12549,N_11871,N_10613);
nand U12550 (N_12550,N_10964,N_10731);
xor U12551 (N_12551,N_11576,N_10891);
nor U12552 (N_12552,N_10930,N_10661);
xnor U12553 (N_12553,N_10665,N_11949);
xor U12554 (N_12554,N_11254,N_10635);
and U12555 (N_12555,N_11827,N_10657);
and U12556 (N_12556,N_11183,N_11313);
nand U12557 (N_12557,N_11837,N_10652);
or U12558 (N_12558,N_11624,N_11063);
nand U12559 (N_12559,N_11154,N_10762);
and U12560 (N_12560,N_11902,N_11778);
or U12561 (N_12561,N_10745,N_11711);
nand U12562 (N_12562,N_10704,N_11970);
and U12563 (N_12563,N_10808,N_11796);
and U12564 (N_12564,N_10721,N_11159);
or U12565 (N_12565,N_11408,N_11085);
or U12566 (N_12566,N_11153,N_11244);
nor U12567 (N_12567,N_10500,N_11613);
nand U12568 (N_12568,N_11995,N_11353);
xnor U12569 (N_12569,N_11235,N_10968);
xnor U12570 (N_12570,N_11756,N_11490);
nor U12571 (N_12571,N_11657,N_11120);
nand U12572 (N_12572,N_10759,N_11179);
or U12573 (N_12573,N_11743,N_11444);
nor U12574 (N_12574,N_10707,N_10918);
nand U12575 (N_12575,N_11322,N_11137);
and U12576 (N_12576,N_11935,N_11823);
or U12577 (N_12577,N_11573,N_11736);
nor U12578 (N_12578,N_11659,N_11758);
xor U12579 (N_12579,N_11700,N_10502);
and U12580 (N_12580,N_11499,N_11369);
nor U12581 (N_12581,N_10883,N_11476);
xor U12582 (N_12582,N_11908,N_11898);
or U12583 (N_12583,N_10671,N_11230);
and U12584 (N_12584,N_11825,N_10590);
nand U12585 (N_12585,N_11685,N_11208);
nand U12586 (N_12586,N_11632,N_11113);
xnor U12587 (N_12587,N_11751,N_11560);
or U12588 (N_12588,N_11114,N_11450);
nand U12589 (N_12589,N_10827,N_11269);
nor U12590 (N_12590,N_10603,N_11682);
and U12591 (N_12591,N_11832,N_10916);
xor U12592 (N_12592,N_10720,N_11264);
nand U12593 (N_12593,N_11975,N_10589);
xor U12594 (N_12594,N_10615,N_10649);
and U12595 (N_12595,N_10899,N_11083);
xnor U12596 (N_12596,N_10662,N_10650);
xnor U12597 (N_12597,N_10507,N_11710);
xnor U12598 (N_12598,N_11656,N_10674);
or U12599 (N_12599,N_11712,N_11918);
nor U12600 (N_12600,N_10864,N_11771);
and U12601 (N_12601,N_11237,N_11599);
nand U12602 (N_12602,N_10909,N_11078);
nor U12603 (N_12603,N_11041,N_11303);
nor U12604 (N_12604,N_11448,N_11757);
nand U12605 (N_12605,N_11399,N_10522);
xnor U12606 (N_12606,N_11214,N_10660);
nand U12607 (N_12607,N_10782,N_11106);
xnor U12608 (N_12608,N_10783,N_11715);
or U12609 (N_12609,N_11091,N_10800);
nor U12610 (N_12610,N_11752,N_11111);
xor U12611 (N_12611,N_11175,N_11807);
xor U12612 (N_12612,N_10813,N_11525);
or U12613 (N_12613,N_11481,N_11750);
and U12614 (N_12614,N_11483,N_11440);
or U12615 (N_12615,N_11620,N_10774);
xnor U12616 (N_12616,N_11309,N_11383);
and U12617 (N_12617,N_11754,N_10879);
nand U12618 (N_12618,N_11627,N_10945);
xnor U12619 (N_12619,N_11066,N_10929);
xor U12620 (N_12620,N_11848,N_10709);
nor U12621 (N_12621,N_11013,N_11282);
nor U12622 (N_12622,N_11520,N_11904);
xor U12623 (N_12623,N_11401,N_10526);
nand U12624 (N_12624,N_11437,N_11228);
nor U12625 (N_12625,N_11859,N_10544);
nand U12626 (N_12626,N_10749,N_11174);
and U12627 (N_12627,N_11500,N_11421);
nand U12628 (N_12628,N_10931,N_11258);
or U12629 (N_12629,N_10678,N_11843);
or U12630 (N_12630,N_11292,N_11088);
nor U12631 (N_12631,N_11343,N_11377);
and U12632 (N_12632,N_11098,N_11394);
nand U12633 (N_12633,N_10537,N_11046);
and U12634 (N_12634,N_11059,N_10560);
and U12635 (N_12635,N_11804,N_11788);
nand U12636 (N_12636,N_11974,N_11635);
nor U12637 (N_12637,N_10596,N_11003);
xor U12638 (N_12638,N_11427,N_11901);
nor U12639 (N_12639,N_10951,N_11874);
or U12640 (N_12640,N_11161,N_11216);
nand U12641 (N_12641,N_11220,N_11497);
xor U12642 (N_12642,N_11923,N_11461);
nor U12643 (N_12643,N_11077,N_10695);
xor U12644 (N_12644,N_10832,N_11423);
nand U12645 (N_12645,N_11767,N_11034);
or U12646 (N_12646,N_11044,N_10924);
xnor U12647 (N_12647,N_11287,N_11928);
or U12648 (N_12648,N_11648,N_11283);
or U12649 (N_12649,N_10640,N_10920);
nand U12650 (N_12650,N_11243,N_11300);
or U12651 (N_12651,N_11360,N_11546);
xor U12652 (N_12652,N_10648,N_11172);
nand U12653 (N_12653,N_11533,N_11734);
or U12654 (N_12654,N_11357,N_11785);
xor U12655 (N_12655,N_11545,N_11212);
or U12656 (N_12656,N_11729,N_10604);
and U12657 (N_12657,N_10894,N_10505);
xor U12658 (N_12658,N_10987,N_11681);
nor U12659 (N_12659,N_11112,N_11236);
or U12660 (N_12660,N_11196,N_11644);
or U12661 (N_12661,N_11422,N_10574);
nand U12662 (N_12662,N_10688,N_10733);
xor U12663 (N_12663,N_11608,N_10753);
or U12664 (N_12664,N_11199,N_11331);
nand U12665 (N_12665,N_11589,N_10737);
xor U12666 (N_12666,N_10767,N_10795);
nand U12667 (N_12667,N_10738,N_10691);
nand U12668 (N_12668,N_11869,N_11163);
or U12669 (N_12669,N_11680,N_11622);
xor U12670 (N_12670,N_11348,N_11839);
nor U12671 (N_12671,N_11355,N_11986);
xor U12672 (N_12672,N_11592,N_11316);
and U12673 (N_12673,N_10797,N_10638);
nor U12674 (N_12674,N_11298,N_11555);
xor U12675 (N_12675,N_11021,N_11531);
nand U12676 (N_12676,N_11435,N_10788);
xor U12677 (N_12677,N_11162,N_11976);
xor U12678 (N_12678,N_11980,N_11391);
xor U12679 (N_12679,N_10582,N_11579);
and U12680 (N_12680,N_10520,N_11086);
or U12681 (N_12681,N_11495,N_11892);
nor U12682 (N_12682,N_11638,N_11379);
xnor U12683 (N_12683,N_11941,N_11362);
and U12684 (N_12684,N_10940,N_11124);
nand U12685 (N_12685,N_10672,N_10804);
xnor U12686 (N_12686,N_10689,N_10750);
and U12687 (N_12687,N_11814,N_10961);
and U12688 (N_12688,N_11655,N_10781);
xnor U12689 (N_12689,N_11135,N_10989);
and U12690 (N_12690,N_11602,N_10802);
nor U12691 (N_12691,N_11117,N_11688);
nor U12692 (N_12692,N_11138,N_11267);
nand U12693 (N_12693,N_10860,N_11407);
and U12694 (N_12694,N_11328,N_11544);
or U12695 (N_12695,N_11816,N_10677);
or U12696 (N_12696,N_11936,N_11634);
nor U12697 (N_12697,N_11144,N_11641);
nand U12698 (N_12698,N_10618,N_11364);
nand U12699 (N_12699,N_11890,N_11761);
or U12700 (N_12700,N_11516,N_11930);
nand U12701 (N_12701,N_10998,N_11045);
nor U12702 (N_12702,N_11626,N_11964);
nand U12703 (N_12703,N_11128,N_10815);
xor U12704 (N_12704,N_11617,N_11108);
or U12705 (N_12705,N_10871,N_11491);
and U12706 (N_12706,N_10515,N_11184);
or U12707 (N_12707,N_11924,N_10617);
nand U12708 (N_12708,N_10634,N_10539);
and U12709 (N_12709,N_10519,N_11043);
and U12710 (N_12710,N_11770,N_10647);
and U12711 (N_12711,N_11866,N_11452);
and U12712 (N_12712,N_10812,N_11019);
or U12713 (N_12713,N_11732,N_10988);
xor U12714 (N_12714,N_11020,N_11475);
nand U12715 (N_12715,N_11195,N_11131);
or U12716 (N_12716,N_10789,N_11204);
and U12717 (N_12717,N_11894,N_11529);
nor U12718 (N_12718,N_11671,N_10791);
or U12719 (N_12719,N_11515,N_10807);
xnor U12720 (N_12720,N_11718,N_11471);
nor U12721 (N_12721,N_11478,N_11725);
or U12722 (N_12722,N_10518,N_11518);
and U12723 (N_12723,N_10503,N_11197);
nand U12724 (N_12724,N_10595,N_11650);
and U12725 (N_12725,N_11070,N_11861);
nor U12726 (N_12726,N_11293,N_11050);
and U12727 (N_12727,N_11464,N_10938);
nor U12728 (N_12728,N_11071,N_11853);
and U12729 (N_12729,N_11514,N_11393);
and U12730 (N_12730,N_11306,N_11817);
nor U12731 (N_12731,N_11669,N_11259);
and U12732 (N_12732,N_11342,N_10554);
xnor U12733 (N_12733,N_11192,N_11616);
nor U12734 (N_12734,N_11856,N_11281);
and U12735 (N_12735,N_11619,N_10885);
and U12736 (N_12736,N_11730,N_11556);
nor U12737 (N_12737,N_10557,N_11972);
nor U12738 (N_12738,N_11170,N_11777);
nor U12739 (N_12739,N_11426,N_11312);
and U12740 (N_12740,N_11541,N_11107);
xnor U12741 (N_12741,N_11442,N_10821);
nor U12742 (N_12742,N_10778,N_11384);
nor U12743 (N_12743,N_10716,N_11910);
or U12744 (N_12744,N_10878,N_10552);
nor U12745 (N_12745,N_11209,N_10935);
xnor U12746 (N_12746,N_11307,N_10625);
and U12747 (N_12747,N_11707,N_11351);
or U12748 (N_12748,N_11002,N_11057);
or U12749 (N_12749,N_10602,N_10833);
nand U12750 (N_12750,N_11748,N_10653);
and U12751 (N_12751,N_11636,N_10836);
and U12752 (N_12752,N_11936,N_10744);
xnor U12753 (N_12753,N_11231,N_10738);
xor U12754 (N_12754,N_11256,N_10521);
nor U12755 (N_12755,N_10552,N_10806);
nor U12756 (N_12756,N_11141,N_10560);
xnor U12757 (N_12757,N_10968,N_11959);
nor U12758 (N_12758,N_11267,N_11964);
nand U12759 (N_12759,N_11896,N_11108);
xnor U12760 (N_12760,N_10895,N_11269);
nand U12761 (N_12761,N_10864,N_10603);
xor U12762 (N_12762,N_10929,N_10648);
xnor U12763 (N_12763,N_10591,N_11850);
xnor U12764 (N_12764,N_10859,N_10897);
and U12765 (N_12765,N_10504,N_11655);
or U12766 (N_12766,N_11431,N_11660);
xor U12767 (N_12767,N_11315,N_11655);
nor U12768 (N_12768,N_11048,N_11746);
nor U12769 (N_12769,N_11094,N_11960);
and U12770 (N_12770,N_10692,N_10783);
or U12771 (N_12771,N_10501,N_11343);
xor U12772 (N_12772,N_10676,N_11293);
or U12773 (N_12773,N_11051,N_11945);
and U12774 (N_12774,N_11796,N_10789);
or U12775 (N_12775,N_11295,N_10669);
nand U12776 (N_12776,N_10555,N_11281);
or U12777 (N_12777,N_11293,N_11540);
nor U12778 (N_12778,N_10560,N_11784);
or U12779 (N_12779,N_11028,N_11410);
xor U12780 (N_12780,N_10862,N_10642);
or U12781 (N_12781,N_11815,N_11312);
and U12782 (N_12782,N_10659,N_11681);
and U12783 (N_12783,N_11977,N_11863);
or U12784 (N_12784,N_11234,N_11011);
nor U12785 (N_12785,N_11778,N_11201);
and U12786 (N_12786,N_11012,N_11087);
and U12787 (N_12787,N_11470,N_11929);
xor U12788 (N_12788,N_10878,N_11245);
and U12789 (N_12789,N_11160,N_11548);
nand U12790 (N_12790,N_10690,N_11804);
or U12791 (N_12791,N_11177,N_11437);
nor U12792 (N_12792,N_11916,N_11341);
and U12793 (N_12793,N_11792,N_10876);
nand U12794 (N_12794,N_10720,N_11119);
and U12795 (N_12795,N_10530,N_11144);
nand U12796 (N_12796,N_11436,N_11975);
and U12797 (N_12797,N_11269,N_11131);
or U12798 (N_12798,N_11713,N_10738);
or U12799 (N_12799,N_11998,N_11832);
nor U12800 (N_12800,N_11882,N_11331);
nor U12801 (N_12801,N_11887,N_11909);
nand U12802 (N_12802,N_11826,N_11928);
or U12803 (N_12803,N_10776,N_10911);
or U12804 (N_12804,N_11443,N_10721);
or U12805 (N_12805,N_11249,N_11267);
nand U12806 (N_12806,N_11183,N_10782);
nor U12807 (N_12807,N_11722,N_11209);
and U12808 (N_12808,N_10599,N_10827);
and U12809 (N_12809,N_11625,N_11530);
xor U12810 (N_12810,N_10500,N_11195);
and U12811 (N_12811,N_11318,N_11803);
nand U12812 (N_12812,N_11566,N_11256);
nand U12813 (N_12813,N_11281,N_11626);
and U12814 (N_12814,N_11250,N_11386);
or U12815 (N_12815,N_11418,N_10930);
or U12816 (N_12816,N_10524,N_11041);
nand U12817 (N_12817,N_10804,N_10616);
xnor U12818 (N_12818,N_11237,N_11642);
or U12819 (N_12819,N_11589,N_11247);
xor U12820 (N_12820,N_10872,N_11313);
nand U12821 (N_12821,N_10520,N_11132);
or U12822 (N_12822,N_11322,N_10703);
xor U12823 (N_12823,N_11771,N_11042);
xnor U12824 (N_12824,N_11101,N_11289);
and U12825 (N_12825,N_10649,N_11088);
and U12826 (N_12826,N_11286,N_10630);
and U12827 (N_12827,N_11607,N_11669);
or U12828 (N_12828,N_11012,N_11187);
or U12829 (N_12829,N_10887,N_10988);
xor U12830 (N_12830,N_11739,N_11400);
xor U12831 (N_12831,N_10779,N_11679);
nand U12832 (N_12832,N_10597,N_10774);
or U12833 (N_12833,N_11164,N_11608);
nand U12834 (N_12834,N_11683,N_11492);
nand U12835 (N_12835,N_11801,N_11944);
or U12836 (N_12836,N_11378,N_11753);
and U12837 (N_12837,N_11623,N_10592);
nor U12838 (N_12838,N_10541,N_11352);
nand U12839 (N_12839,N_10939,N_10534);
nor U12840 (N_12840,N_10840,N_11153);
and U12841 (N_12841,N_10902,N_11464);
and U12842 (N_12842,N_11067,N_11185);
nand U12843 (N_12843,N_11758,N_11035);
xor U12844 (N_12844,N_11394,N_11800);
or U12845 (N_12845,N_10609,N_10840);
xor U12846 (N_12846,N_11708,N_10682);
or U12847 (N_12847,N_11114,N_11145);
or U12848 (N_12848,N_11805,N_11858);
and U12849 (N_12849,N_10745,N_11478);
nor U12850 (N_12850,N_11166,N_11826);
nand U12851 (N_12851,N_10660,N_10982);
or U12852 (N_12852,N_11943,N_11740);
nor U12853 (N_12853,N_11156,N_11597);
and U12854 (N_12854,N_10625,N_10858);
and U12855 (N_12855,N_11194,N_10906);
xnor U12856 (N_12856,N_11567,N_10932);
and U12857 (N_12857,N_10508,N_10839);
or U12858 (N_12858,N_10673,N_10960);
and U12859 (N_12859,N_11735,N_11475);
xor U12860 (N_12860,N_11852,N_11688);
or U12861 (N_12861,N_11179,N_11517);
or U12862 (N_12862,N_10665,N_11672);
nor U12863 (N_12863,N_10660,N_11445);
or U12864 (N_12864,N_11344,N_11400);
xor U12865 (N_12865,N_10587,N_11191);
xor U12866 (N_12866,N_11110,N_11387);
nor U12867 (N_12867,N_10567,N_11311);
nor U12868 (N_12868,N_10982,N_11973);
nor U12869 (N_12869,N_11382,N_11392);
and U12870 (N_12870,N_11133,N_10838);
and U12871 (N_12871,N_11739,N_10694);
nor U12872 (N_12872,N_10505,N_11125);
nand U12873 (N_12873,N_10904,N_11908);
and U12874 (N_12874,N_10803,N_11010);
nand U12875 (N_12875,N_11800,N_10793);
and U12876 (N_12876,N_11465,N_11626);
nand U12877 (N_12877,N_10783,N_10900);
xnor U12878 (N_12878,N_11698,N_11850);
or U12879 (N_12879,N_11983,N_11043);
nand U12880 (N_12880,N_10890,N_11766);
xor U12881 (N_12881,N_11478,N_11240);
nand U12882 (N_12882,N_11252,N_11829);
nand U12883 (N_12883,N_11242,N_11971);
xnor U12884 (N_12884,N_11200,N_11488);
and U12885 (N_12885,N_10588,N_10543);
or U12886 (N_12886,N_11452,N_11119);
and U12887 (N_12887,N_11907,N_11923);
or U12888 (N_12888,N_11280,N_11681);
and U12889 (N_12889,N_11284,N_11418);
or U12890 (N_12890,N_11569,N_10858);
and U12891 (N_12891,N_11515,N_11400);
xor U12892 (N_12892,N_11321,N_10689);
and U12893 (N_12893,N_10657,N_11162);
nand U12894 (N_12894,N_11815,N_11428);
xnor U12895 (N_12895,N_11233,N_11463);
nor U12896 (N_12896,N_11968,N_10641);
or U12897 (N_12897,N_10717,N_11896);
nor U12898 (N_12898,N_11590,N_10667);
or U12899 (N_12899,N_10678,N_11460);
nor U12900 (N_12900,N_11576,N_10584);
and U12901 (N_12901,N_10906,N_11229);
xnor U12902 (N_12902,N_11373,N_11827);
or U12903 (N_12903,N_11934,N_11294);
or U12904 (N_12904,N_10675,N_10632);
or U12905 (N_12905,N_11567,N_11347);
xor U12906 (N_12906,N_11393,N_11438);
xnor U12907 (N_12907,N_11710,N_11782);
nor U12908 (N_12908,N_10590,N_10908);
xor U12909 (N_12909,N_11460,N_11076);
and U12910 (N_12910,N_10757,N_10932);
xor U12911 (N_12911,N_10865,N_11636);
nand U12912 (N_12912,N_10661,N_11571);
xor U12913 (N_12913,N_11568,N_10784);
xor U12914 (N_12914,N_11930,N_11712);
or U12915 (N_12915,N_10514,N_11108);
xor U12916 (N_12916,N_10528,N_11078);
xnor U12917 (N_12917,N_11201,N_11326);
nand U12918 (N_12918,N_11550,N_11095);
or U12919 (N_12919,N_11248,N_11867);
nor U12920 (N_12920,N_10954,N_11509);
and U12921 (N_12921,N_11619,N_11518);
or U12922 (N_12922,N_11648,N_11785);
xnor U12923 (N_12923,N_11193,N_10545);
nor U12924 (N_12924,N_10503,N_11054);
xnor U12925 (N_12925,N_11271,N_11297);
xnor U12926 (N_12926,N_11826,N_10760);
nor U12927 (N_12927,N_11479,N_10984);
nor U12928 (N_12928,N_10977,N_11078);
nor U12929 (N_12929,N_11449,N_11870);
or U12930 (N_12930,N_10511,N_11890);
or U12931 (N_12931,N_11218,N_11355);
nand U12932 (N_12932,N_11861,N_10996);
nand U12933 (N_12933,N_11367,N_11712);
nor U12934 (N_12934,N_11288,N_10792);
nor U12935 (N_12935,N_10672,N_11593);
nor U12936 (N_12936,N_10639,N_11128);
and U12937 (N_12937,N_11225,N_11134);
nand U12938 (N_12938,N_11596,N_11108);
nor U12939 (N_12939,N_11412,N_11265);
nor U12940 (N_12940,N_11994,N_10763);
or U12941 (N_12941,N_11625,N_10621);
and U12942 (N_12942,N_10853,N_10913);
xor U12943 (N_12943,N_11728,N_10954);
and U12944 (N_12944,N_11743,N_11425);
and U12945 (N_12945,N_11977,N_11910);
nor U12946 (N_12946,N_11780,N_11167);
nor U12947 (N_12947,N_10820,N_11433);
xnor U12948 (N_12948,N_11934,N_11059);
nor U12949 (N_12949,N_10662,N_11290);
nor U12950 (N_12950,N_10638,N_11315);
nand U12951 (N_12951,N_11536,N_11266);
xnor U12952 (N_12952,N_11318,N_11272);
nand U12953 (N_12953,N_10618,N_10836);
nand U12954 (N_12954,N_11409,N_10852);
or U12955 (N_12955,N_11976,N_10918);
nand U12956 (N_12956,N_11189,N_11607);
and U12957 (N_12957,N_10599,N_10760);
or U12958 (N_12958,N_10740,N_11340);
xnor U12959 (N_12959,N_11692,N_10849);
or U12960 (N_12960,N_10546,N_11648);
or U12961 (N_12961,N_11141,N_10527);
and U12962 (N_12962,N_11208,N_11131);
xor U12963 (N_12963,N_10576,N_11122);
nor U12964 (N_12964,N_11347,N_10843);
nand U12965 (N_12965,N_11345,N_11737);
nor U12966 (N_12966,N_11966,N_11076);
and U12967 (N_12967,N_11903,N_11893);
xor U12968 (N_12968,N_11541,N_11307);
xnor U12969 (N_12969,N_11907,N_11580);
nand U12970 (N_12970,N_11806,N_11845);
xnor U12971 (N_12971,N_10807,N_11985);
xnor U12972 (N_12972,N_11451,N_11069);
or U12973 (N_12973,N_10757,N_11157);
nand U12974 (N_12974,N_11777,N_11461);
and U12975 (N_12975,N_11308,N_10707);
and U12976 (N_12976,N_11654,N_11614);
nor U12977 (N_12977,N_11348,N_11167);
and U12978 (N_12978,N_11929,N_11339);
nor U12979 (N_12979,N_11300,N_11131);
or U12980 (N_12980,N_10524,N_10672);
and U12981 (N_12981,N_10657,N_11552);
and U12982 (N_12982,N_11959,N_10782);
xnor U12983 (N_12983,N_10851,N_11202);
or U12984 (N_12984,N_10945,N_11455);
nand U12985 (N_12985,N_11899,N_10680);
and U12986 (N_12986,N_11915,N_11124);
and U12987 (N_12987,N_11727,N_11631);
nand U12988 (N_12988,N_11672,N_11379);
or U12989 (N_12989,N_11760,N_11506);
and U12990 (N_12990,N_10815,N_11899);
nand U12991 (N_12991,N_11731,N_11108);
and U12992 (N_12992,N_11847,N_11385);
or U12993 (N_12993,N_10976,N_11733);
xnor U12994 (N_12994,N_11122,N_11868);
xor U12995 (N_12995,N_10578,N_11091);
nand U12996 (N_12996,N_11552,N_11628);
and U12997 (N_12997,N_11647,N_11424);
nand U12998 (N_12998,N_10747,N_11915);
nand U12999 (N_12999,N_10563,N_11218);
or U13000 (N_13000,N_10519,N_10664);
and U13001 (N_13001,N_11072,N_11788);
nand U13002 (N_13002,N_11223,N_11417);
or U13003 (N_13003,N_11820,N_11255);
and U13004 (N_13004,N_11563,N_11718);
nor U13005 (N_13005,N_10884,N_11408);
nand U13006 (N_13006,N_11476,N_11131);
or U13007 (N_13007,N_11091,N_11172);
nand U13008 (N_13008,N_11217,N_10892);
nor U13009 (N_13009,N_11963,N_11710);
nor U13010 (N_13010,N_11783,N_10565);
nor U13011 (N_13011,N_10501,N_11200);
and U13012 (N_13012,N_11566,N_10690);
or U13013 (N_13013,N_11778,N_11730);
or U13014 (N_13014,N_10992,N_11799);
or U13015 (N_13015,N_10513,N_11465);
nor U13016 (N_13016,N_11032,N_11939);
nand U13017 (N_13017,N_11331,N_10964);
and U13018 (N_13018,N_11236,N_11627);
and U13019 (N_13019,N_10526,N_11673);
or U13020 (N_13020,N_10886,N_11288);
or U13021 (N_13021,N_11018,N_11933);
xor U13022 (N_13022,N_11705,N_10504);
nor U13023 (N_13023,N_11331,N_10858);
xor U13024 (N_13024,N_11111,N_11887);
and U13025 (N_13025,N_10528,N_10709);
nor U13026 (N_13026,N_11398,N_11256);
or U13027 (N_13027,N_11219,N_10652);
or U13028 (N_13028,N_11239,N_11638);
nor U13029 (N_13029,N_11379,N_11328);
or U13030 (N_13030,N_10835,N_11834);
nor U13031 (N_13031,N_10521,N_11996);
or U13032 (N_13032,N_11256,N_11678);
or U13033 (N_13033,N_10870,N_10658);
nand U13034 (N_13034,N_11625,N_10819);
xnor U13035 (N_13035,N_11838,N_10528);
or U13036 (N_13036,N_11935,N_11704);
or U13037 (N_13037,N_10904,N_10727);
xor U13038 (N_13038,N_11714,N_10673);
nor U13039 (N_13039,N_10709,N_11785);
or U13040 (N_13040,N_11560,N_11658);
and U13041 (N_13041,N_11406,N_10852);
nand U13042 (N_13042,N_11152,N_11307);
nand U13043 (N_13043,N_11330,N_11211);
or U13044 (N_13044,N_10996,N_11566);
nor U13045 (N_13045,N_11570,N_11724);
or U13046 (N_13046,N_10880,N_11705);
nand U13047 (N_13047,N_11526,N_11681);
nor U13048 (N_13048,N_10689,N_11249);
xnor U13049 (N_13049,N_11773,N_10685);
nand U13050 (N_13050,N_10990,N_10837);
or U13051 (N_13051,N_11989,N_11841);
and U13052 (N_13052,N_11101,N_10630);
and U13053 (N_13053,N_11253,N_11686);
nor U13054 (N_13054,N_10751,N_11069);
xnor U13055 (N_13055,N_11563,N_11881);
and U13056 (N_13056,N_11481,N_11189);
nand U13057 (N_13057,N_10824,N_11631);
xor U13058 (N_13058,N_10858,N_11966);
and U13059 (N_13059,N_10779,N_10988);
xor U13060 (N_13060,N_11357,N_11193);
xnor U13061 (N_13061,N_11847,N_11570);
or U13062 (N_13062,N_11141,N_10772);
xor U13063 (N_13063,N_11867,N_10861);
or U13064 (N_13064,N_11381,N_11886);
nand U13065 (N_13065,N_11092,N_10753);
or U13066 (N_13066,N_10982,N_11135);
and U13067 (N_13067,N_11298,N_10796);
nor U13068 (N_13068,N_11462,N_11177);
or U13069 (N_13069,N_11547,N_11984);
xnor U13070 (N_13070,N_11253,N_10576);
or U13071 (N_13071,N_11280,N_11387);
nor U13072 (N_13072,N_10567,N_11307);
nand U13073 (N_13073,N_10847,N_11260);
nor U13074 (N_13074,N_10674,N_11569);
and U13075 (N_13075,N_10663,N_11674);
or U13076 (N_13076,N_10753,N_10659);
or U13077 (N_13077,N_11339,N_10968);
xnor U13078 (N_13078,N_11679,N_11610);
nor U13079 (N_13079,N_11815,N_11436);
nor U13080 (N_13080,N_11216,N_11709);
or U13081 (N_13081,N_11823,N_11811);
or U13082 (N_13082,N_10614,N_10923);
nand U13083 (N_13083,N_11041,N_10959);
nor U13084 (N_13084,N_11821,N_11478);
and U13085 (N_13085,N_11205,N_11601);
nand U13086 (N_13086,N_10718,N_11358);
xor U13087 (N_13087,N_11483,N_11825);
or U13088 (N_13088,N_10751,N_11196);
xnor U13089 (N_13089,N_10506,N_10916);
nor U13090 (N_13090,N_11693,N_11796);
or U13091 (N_13091,N_11627,N_11872);
xor U13092 (N_13092,N_10603,N_11161);
xor U13093 (N_13093,N_11954,N_11084);
nand U13094 (N_13094,N_11439,N_11121);
and U13095 (N_13095,N_10606,N_11229);
xnor U13096 (N_13096,N_10907,N_11192);
nor U13097 (N_13097,N_11303,N_11546);
and U13098 (N_13098,N_11707,N_11621);
or U13099 (N_13099,N_11103,N_11006);
xnor U13100 (N_13100,N_11583,N_11523);
and U13101 (N_13101,N_11766,N_11892);
and U13102 (N_13102,N_10618,N_11150);
and U13103 (N_13103,N_11937,N_11277);
nand U13104 (N_13104,N_11147,N_11322);
and U13105 (N_13105,N_10542,N_11809);
xnor U13106 (N_13106,N_11236,N_11354);
or U13107 (N_13107,N_10644,N_11358);
xor U13108 (N_13108,N_10754,N_11437);
nor U13109 (N_13109,N_11943,N_10897);
xnor U13110 (N_13110,N_11006,N_10689);
nand U13111 (N_13111,N_10926,N_10836);
xnor U13112 (N_13112,N_10925,N_11541);
or U13113 (N_13113,N_11399,N_10963);
and U13114 (N_13114,N_10966,N_11517);
nor U13115 (N_13115,N_11498,N_10804);
and U13116 (N_13116,N_10986,N_10899);
or U13117 (N_13117,N_10535,N_10948);
xnor U13118 (N_13118,N_11095,N_11483);
nand U13119 (N_13119,N_11423,N_10645);
xor U13120 (N_13120,N_11464,N_10884);
or U13121 (N_13121,N_10870,N_11508);
or U13122 (N_13122,N_11814,N_10978);
and U13123 (N_13123,N_11820,N_10533);
xnor U13124 (N_13124,N_11051,N_11585);
nor U13125 (N_13125,N_10527,N_10551);
or U13126 (N_13126,N_11321,N_11135);
nand U13127 (N_13127,N_11205,N_10910);
and U13128 (N_13128,N_10988,N_11600);
or U13129 (N_13129,N_11610,N_10803);
xnor U13130 (N_13130,N_11234,N_10849);
or U13131 (N_13131,N_10753,N_10729);
or U13132 (N_13132,N_11641,N_11472);
and U13133 (N_13133,N_11392,N_10986);
and U13134 (N_13134,N_11314,N_11598);
or U13135 (N_13135,N_11852,N_11174);
or U13136 (N_13136,N_11554,N_11329);
nand U13137 (N_13137,N_11967,N_11637);
and U13138 (N_13138,N_10721,N_11525);
and U13139 (N_13139,N_10915,N_10549);
nor U13140 (N_13140,N_10930,N_10600);
nand U13141 (N_13141,N_11557,N_10864);
xnor U13142 (N_13142,N_11258,N_10927);
and U13143 (N_13143,N_10990,N_10925);
nand U13144 (N_13144,N_11313,N_11729);
and U13145 (N_13145,N_11567,N_11510);
nand U13146 (N_13146,N_11301,N_11809);
nand U13147 (N_13147,N_10915,N_11435);
or U13148 (N_13148,N_11682,N_11800);
xnor U13149 (N_13149,N_11729,N_10920);
and U13150 (N_13150,N_10811,N_11598);
nand U13151 (N_13151,N_10992,N_11904);
nand U13152 (N_13152,N_10609,N_11130);
nand U13153 (N_13153,N_11211,N_11452);
or U13154 (N_13154,N_10549,N_11430);
or U13155 (N_13155,N_11646,N_11990);
nor U13156 (N_13156,N_10907,N_10651);
nand U13157 (N_13157,N_11677,N_10844);
nor U13158 (N_13158,N_10892,N_10792);
nor U13159 (N_13159,N_10710,N_11471);
or U13160 (N_13160,N_11918,N_11555);
nand U13161 (N_13161,N_10861,N_11492);
nor U13162 (N_13162,N_11805,N_11303);
or U13163 (N_13163,N_11324,N_11883);
xnor U13164 (N_13164,N_11148,N_11864);
nand U13165 (N_13165,N_11523,N_11287);
or U13166 (N_13166,N_11590,N_11065);
nor U13167 (N_13167,N_11148,N_10816);
xor U13168 (N_13168,N_11394,N_11273);
and U13169 (N_13169,N_10840,N_11326);
or U13170 (N_13170,N_10645,N_11157);
nor U13171 (N_13171,N_10821,N_10648);
nand U13172 (N_13172,N_10778,N_11105);
and U13173 (N_13173,N_11528,N_11754);
and U13174 (N_13174,N_10572,N_10620);
nand U13175 (N_13175,N_10668,N_11781);
xor U13176 (N_13176,N_11485,N_10545);
nand U13177 (N_13177,N_10706,N_11266);
or U13178 (N_13178,N_11134,N_11342);
nor U13179 (N_13179,N_11561,N_10949);
and U13180 (N_13180,N_11177,N_11207);
or U13181 (N_13181,N_11563,N_11944);
nand U13182 (N_13182,N_10673,N_11893);
or U13183 (N_13183,N_10567,N_10579);
xnor U13184 (N_13184,N_11138,N_11261);
nand U13185 (N_13185,N_10600,N_11468);
nor U13186 (N_13186,N_11892,N_11765);
nand U13187 (N_13187,N_11614,N_11400);
nand U13188 (N_13188,N_11575,N_11681);
nand U13189 (N_13189,N_11931,N_10504);
and U13190 (N_13190,N_11423,N_11650);
nand U13191 (N_13191,N_10530,N_11778);
nor U13192 (N_13192,N_10703,N_10588);
xor U13193 (N_13193,N_11420,N_11483);
and U13194 (N_13194,N_11759,N_11432);
xor U13195 (N_13195,N_10635,N_10892);
xor U13196 (N_13196,N_11532,N_11451);
or U13197 (N_13197,N_11551,N_11595);
xor U13198 (N_13198,N_10506,N_11931);
and U13199 (N_13199,N_11358,N_11631);
or U13200 (N_13200,N_11299,N_11171);
xnor U13201 (N_13201,N_11400,N_10721);
nand U13202 (N_13202,N_10566,N_11156);
nor U13203 (N_13203,N_10615,N_11508);
and U13204 (N_13204,N_10533,N_11735);
nor U13205 (N_13205,N_11815,N_10557);
or U13206 (N_13206,N_11005,N_11932);
and U13207 (N_13207,N_11073,N_11523);
and U13208 (N_13208,N_11471,N_10517);
or U13209 (N_13209,N_10826,N_10832);
nor U13210 (N_13210,N_11501,N_11903);
nand U13211 (N_13211,N_11328,N_11926);
nand U13212 (N_13212,N_11578,N_11049);
nand U13213 (N_13213,N_11314,N_10802);
xor U13214 (N_13214,N_10773,N_11560);
nand U13215 (N_13215,N_11551,N_11041);
or U13216 (N_13216,N_11233,N_10952);
and U13217 (N_13217,N_11771,N_10542);
nor U13218 (N_13218,N_10732,N_11203);
or U13219 (N_13219,N_11855,N_11866);
nor U13220 (N_13220,N_11327,N_11652);
and U13221 (N_13221,N_11345,N_11328);
and U13222 (N_13222,N_11746,N_10865);
nor U13223 (N_13223,N_11815,N_10649);
nand U13224 (N_13224,N_11596,N_11379);
xnor U13225 (N_13225,N_10703,N_11989);
nand U13226 (N_13226,N_11775,N_10670);
and U13227 (N_13227,N_11697,N_10956);
xnor U13228 (N_13228,N_10794,N_10571);
and U13229 (N_13229,N_11894,N_10632);
nand U13230 (N_13230,N_10573,N_11981);
nor U13231 (N_13231,N_11369,N_11297);
and U13232 (N_13232,N_11513,N_11230);
nand U13233 (N_13233,N_10658,N_11121);
nor U13234 (N_13234,N_10916,N_10606);
and U13235 (N_13235,N_10662,N_10827);
nand U13236 (N_13236,N_10734,N_10778);
xor U13237 (N_13237,N_10548,N_10990);
nand U13238 (N_13238,N_11238,N_11503);
xnor U13239 (N_13239,N_11864,N_11189);
and U13240 (N_13240,N_10989,N_10850);
nand U13241 (N_13241,N_11628,N_11063);
or U13242 (N_13242,N_10580,N_11981);
nand U13243 (N_13243,N_11131,N_11008);
nand U13244 (N_13244,N_11977,N_10585);
and U13245 (N_13245,N_11220,N_11206);
nor U13246 (N_13246,N_10782,N_10553);
nand U13247 (N_13247,N_10514,N_11178);
and U13248 (N_13248,N_11547,N_11691);
and U13249 (N_13249,N_11022,N_11305);
nor U13250 (N_13250,N_10740,N_10854);
and U13251 (N_13251,N_11395,N_10740);
nor U13252 (N_13252,N_10517,N_10761);
xnor U13253 (N_13253,N_11967,N_10717);
nor U13254 (N_13254,N_11587,N_11110);
nand U13255 (N_13255,N_11281,N_10798);
nand U13256 (N_13256,N_10831,N_10871);
nand U13257 (N_13257,N_11973,N_10541);
xor U13258 (N_13258,N_10732,N_11554);
and U13259 (N_13259,N_11451,N_11692);
nor U13260 (N_13260,N_11093,N_11602);
nor U13261 (N_13261,N_11813,N_10959);
and U13262 (N_13262,N_11326,N_11539);
or U13263 (N_13263,N_11232,N_11723);
or U13264 (N_13264,N_11174,N_11309);
nor U13265 (N_13265,N_11152,N_11286);
nor U13266 (N_13266,N_11789,N_11942);
nor U13267 (N_13267,N_10646,N_11950);
and U13268 (N_13268,N_10551,N_11198);
xor U13269 (N_13269,N_11251,N_11012);
xnor U13270 (N_13270,N_11571,N_11671);
xor U13271 (N_13271,N_10587,N_10584);
or U13272 (N_13272,N_11373,N_10700);
nand U13273 (N_13273,N_10899,N_11626);
or U13274 (N_13274,N_11713,N_10526);
nand U13275 (N_13275,N_11544,N_11248);
or U13276 (N_13276,N_11828,N_11754);
nor U13277 (N_13277,N_10829,N_11272);
nor U13278 (N_13278,N_10696,N_10603);
nor U13279 (N_13279,N_11599,N_11318);
xnor U13280 (N_13280,N_10667,N_10791);
or U13281 (N_13281,N_11707,N_11625);
nand U13282 (N_13282,N_11438,N_11972);
nor U13283 (N_13283,N_11118,N_11713);
xnor U13284 (N_13284,N_11831,N_11758);
xor U13285 (N_13285,N_11993,N_10887);
nor U13286 (N_13286,N_10604,N_11657);
nor U13287 (N_13287,N_11726,N_10858);
or U13288 (N_13288,N_11384,N_11304);
and U13289 (N_13289,N_11746,N_10593);
nand U13290 (N_13290,N_11231,N_11144);
nand U13291 (N_13291,N_11315,N_10977);
and U13292 (N_13292,N_11357,N_10601);
or U13293 (N_13293,N_10860,N_11843);
nand U13294 (N_13294,N_11833,N_11141);
and U13295 (N_13295,N_11905,N_10803);
and U13296 (N_13296,N_11227,N_10606);
or U13297 (N_13297,N_11632,N_11684);
or U13298 (N_13298,N_10920,N_10608);
xnor U13299 (N_13299,N_10581,N_10510);
nand U13300 (N_13300,N_10976,N_11471);
and U13301 (N_13301,N_11650,N_11442);
nand U13302 (N_13302,N_10549,N_11161);
nor U13303 (N_13303,N_10905,N_11501);
xor U13304 (N_13304,N_11581,N_10747);
or U13305 (N_13305,N_11816,N_11006);
nand U13306 (N_13306,N_11187,N_11010);
xor U13307 (N_13307,N_11030,N_11817);
and U13308 (N_13308,N_11625,N_11601);
xnor U13309 (N_13309,N_11461,N_11678);
nor U13310 (N_13310,N_11316,N_11885);
or U13311 (N_13311,N_10546,N_11276);
nand U13312 (N_13312,N_11898,N_10813);
nor U13313 (N_13313,N_11583,N_10733);
nand U13314 (N_13314,N_11563,N_11608);
xor U13315 (N_13315,N_11341,N_11464);
or U13316 (N_13316,N_11528,N_11272);
nor U13317 (N_13317,N_11786,N_11827);
or U13318 (N_13318,N_11602,N_11556);
and U13319 (N_13319,N_11321,N_11301);
nor U13320 (N_13320,N_10962,N_10996);
nor U13321 (N_13321,N_11904,N_11718);
or U13322 (N_13322,N_11920,N_11209);
nor U13323 (N_13323,N_11464,N_11174);
nand U13324 (N_13324,N_10909,N_11659);
xnor U13325 (N_13325,N_10872,N_11130);
and U13326 (N_13326,N_11399,N_11515);
or U13327 (N_13327,N_11119,N_11321);
nor U13328 (N_13328,N_10522,N_10838);
nand U13329 (N_13329,N_11840,N_11712);
or U13330 (N_13330,N_10985,N_11945);
nand U13331 (N_13331,N_10699,N_11979);
or U13332 (N_13332,N_11566,N_11389);
xnor U13333 (N_13333,N_11089,N_11990);
nand U13334 (N_13334,N_11927,N_11461);
nand U13335 (N_13335,N_11440,N_10601);
and U13336 (N_13336,N_11869,N_11587);
nand U13337 (N_13337,N_10764,N_11439);
or U13338 (N_13338,N_11083,N_10691);
nand U13339 (N_13339,N_11783,N_10527);
or U13340 (N_13340,N_11267,N_10817);
nand U13341 (N_13341,N_11159,N_10518);
nor U13342 (N_13342,N_11757,N_11702);
and U13343 (N_13343,N_10764,N_10845);
nor U13344 (N_13344,N_11345,N_11337);
or U13345 (N_13345,N_10705,N_10721);
nand U13346 (N_13346,N_10951,N_11843);
xnor U13347 (N_13347,N_10534,N_10922);
or U13348 (N_13348,N_11632,N_10780);
or U13349 (N_13349,N_11208,N_10825);
and U13350 (N_13350,N_11512,N_11579);
nor U13351 (N_13351,N_10965,N_10824);
nand U13352 (N_13352,N_11213,N_10966);
or U13353 (N_13353,N_11805,N_10677);
nor U13354 (N_13354,N_10567,N_10800);
nor U13355 (N_13355,N_10855,N_11616);
xor U13356 (N_13356,N_10843,N_10943);
xor U13357 (N_13357,N_10584,N_11358);
nor U13358 (N_13358,N_11684,N_11020);
or U13359 (N_13359,N_11491,N_10788);
nor U13360 (N_13360,N_10625,N_11246);
and U13361 (N_13361,N_11328,N_11321);
or U13362 (N_13362,N_11089,N_11682);
nand U13363 (N_13363,N_10738,N_11348);
xnor U13364 (N_13364,N_10909,N_11849);
nor U13365 (N_13365,N_11635,N_11933);
or U13366 (N_13366,N_11148,N_10620);
or U13367 (N_13367,N_11894,N_11206);
nor U13368 (N_13368,N_10954,N_10686);
nor U13369 (N_13369,N_10954,N_11964);
xor U13370 (N_13370,N_11396,N_10917);
and U13371 (N_13371,N_11390,N_11201);
nor U13372 (N_13372,N_11065,N_11216);
nor U13373 (N_13373,N_11045,N_10996);
and U13374 (N_13374,N_10562,N_10766);
and U13375 (N_13375,N_11330,N_10983);
xor U13376 (N_13376,N_10890,N_11117);
nand U13377 (N_13377,N_11737,N_10601);
nand U13378 (N_13378,N_11102,N_10696);
xor U13379 (N_13379,N_10966,N_10644);
and U13380 (N_13380,N_11645,N_11142);
nor U13381 (N_13381,N_11187,N_10647);
nand U13382 (N_13382,N_11470,N_10950);
xnor U13383 (N_13383,N_10978,N_11660);
nand U13384 (N_13384,N_11545,N_10693);
nor U13385 (N_13385,N_11811,N_11817);
and U13386 (N_13386,N_10599,N_10784);
and U13387 (N_13387,N_11585,N_11901);
nand U13388 (N_13388,N_11060,N_11748);
nand U13389 (N_13389,N_11570,N_11109);
nand U13390 (N_13390,N_11567,N_11285);
or U13391 (N_13391,N_11556,N_10535);
nor U13392 (N_13392,N_11988,N_11598);
nor U13393 (N_13393,N_11147,N_11745);
xor U13394 (N_13394,N_11670,N_11690);
nand U13395 (N_13395,N_10540,N_10650);
and U13396 (N_13396,N_11357,N_11611);
xor U13397 (N_13397,N_11328,N_10565);
nand U13398 (N_13398,N_11271,N_10825);
nor U13399 (N_13399,N_11127,N_11536);
xnor U13400 (N_13400,N_11324,N_11403);
xnor U13401 (N_13401,N_11609,N_11180);
or U13402 (N_13402,N_11108,N_11654);
nand U13403 (N_13403,N_11025,N_11277);
nand U13404 (N_13404,N_11951,N_10728);
nor U13405 (N_13405,N_11788,N_11298);
nand U13406 (N_13406,N_11559,N_11447);
nor U13407 (N_13407,N_11641,N_11568);
or U13408 (N_13408,N_10635,N_11596);
nand U13409 (N_13409,N_11412,N_11541);
nor U13410 (N_13410,N_11946,N_11321);
or U13411 (N_13411,N_11406,N_11396);
and U13412 (N_13412,N_10957,N_11735);
and U13413 (N_13413,N_11723,N_10948);
or U13414 (N_13414,N_11260,N_11947);
nand U13415 (N_13415,N_11338,N_11466);
nand U13416 (N_13416,N_11785,N_10519);
nor U13417 (N_13417,N_10573,N_11216);
nand U13418 (N_13418,N_10730,N_11564);
and U13419 (N_13419,N_11710,N_10633);
and U13420 (N_13420,N_11877,N_11090);
or U13421 (N_13421,N_11408,N_10968);
and U13422 (N_13422,N_11028,N_10872);
nand U13423 (N_13423,N_10869,N_11168);
nand U13424 (N_13424,N_11393,N_11384);
nor U13425 (N_13425,N_11977,N_11611);
and U13426 (N_13426,N_11114,N_11516);
or U13427 (N_13427,N_11401,N_11074);
and U13428 (N_13428,N_11641,N_11111);
nand U13429 (N_13429,N_11601,N_11690);
or U13430 (N_13430,N_11423,N_10996);
or U13431 (N_13431,N_10833,N_10767);
or U13432 (N_13432,N_10693,N_11831);
or U13433 (N_13433,N_11917,N_10516);
and U13434 (N_13434,N_11991,N_10947);
nor U13435 (N_13435,N_10825,N_11986);
and U13436 (N_13436,N_10844,N_11333);
nand U13437 (N_13437,N_11304,N_11720);
nand U13438 (N_13438,N_11220,N_10594);
nor U13439 (N_13439,N_11130,N_10858);
nor U13440 (N_13440,N_11449,N_10830);
xnor U13441 (N_13441,N_10865,N_11409);
nand U13442 (N_13442,N_10642,N_11975);
nor U13443 (N_13443,N_11152,N_11478);
nand U13444 (N_13444,N_11968,N_11326);
or U13445 (N_13445,N_11824,N_10965);
xnor U13446 (N_13446,N_11107,N_11905);
or U13447 (N_13447,N_10790,N_11533);
nand U13448 (N_13448,N_11960,N_10662);
nor U13449 (N_13449,N_11018,N_11622);
nor U13450 (N_13450,N_11026,N_11682);
xor U13451 (N_13451,N_11963,N_11905);
and U13452 (N_13452,N_10510,N_11424);
and U13453 (N_13453,N_11719,N_11150);
nor U13454 (N_13454,N_11532,N_10564);
nand U13455 (N_13455,N_10571,N_10593);
nand U13456 (N_13456,N_11400,N_10740);
nor U13457 (N_13457,N_11378,N_11002);
and U13458 (N_13458,N_11608,N_10997);
nor U13459 (N_13459,N_10583,N_11643);
xor U13460 (N_13460,N_11166,N_10583);
and U13461 (N_13461,N_11361,N_11904);
and U13462 (N_13462,N_11272,N_11574);
and U13463 (N_13463,N_10981,N_10620);
nand U13464 (N_13464,N_10766,N_11743);
or U13465 (N_13465,N_11185,N_11299);
xnor U13466 (N_13466,N_11129,N_11748);
nand U13467 (N_13467,N_10885,N_11887);
nand U13468 (N_13468,N_11858,N_10516);
xnor U13469 (N_13469,N_11501,N_11803);
and U13470 (N_13470,N_11220,N_11812);
nor U13471 (N_13471,N_10730,N_10621);
nor U13472 (N_13472,N_11332,N_11515);
or U13473 (N_13473,N_10607,N_11825);
xnor U13474 (N_13474,N_11535,N_11635);
xor U13475 (N_13475,N_10555,N_11891);
xor U13476 (N_13476,N_11523,N_10566);
nor U13477 (N_13477,N_10786,N_11275);
nor U13478 (N_13478,N_11212,N_10775);
or U13479 (N_13479,N_11061,N_11480);
xor U13480 (N_13480,N_11811,N_11211);
nand U13481 (N_13481,N_11307,N_11599);
xnor U13482 (N_13482,N_10993,N_11019);
nand U13483 (N_13483,N_11733,N_10935);
nor U13484 (N_13484,N_10828,N_11143);
and U13485 (N_13485,N_11418,N_11895);
or U13486 (N_13486,N_11239,N_10756);
or U13487 (N_13487,N_10745,N_11021);
nand U13488 (N_13488,N_11285,N_11167);
nor U13489 (N_13489,N_11518,N_11786);
nand U13490 (N_13490,N_11849,N_11172);
and U13491 (N_13491,N_11492,N_11890);
or U13492 (N_13492,N_11839,N_11158);
nor U13493 (N_13493,N_11194,N_10716);
xor U13494 (N_13494,N_11604,N_10582);
nor U13495 (N_13495,N_11485,N_11745);
xnor U13496 (N_13496,N_10868,N_11841);
xnor U13497 (N_13497,N_11488,N_11829);
xor U13498 (N_13498,N_11438,N_11992);
nor U13499 (N_13499,N_10606,N_10871);
nand U13500 (N_13500,N_13046,N_12126);
and U13501 (N_13501,N_13312,N_13211);
nor U13502 (N_13502,N_13339,N_13220);
xnor U13503 (N_13503,N_12374,N_13152);
and U13504 (N_13504,N_12460,N_12343);
and U13505 (N_13505,N_12244,N_12507);
or U13506 (N_13506,N_12956,N_13428);
xor U13507 (N_13507,N_12446,N_13116);
and U13508 (N_13508,N_12425,N_12058);
and U13509 (N_13509,N_12540,N_12825);
and U13510 (N_13510,N_12055,N_13385);
xnor U13511 (N_13511,N_12490,N_13283);
or U13512 (N_13512,N_13307,N_12672);
xnor U13513 (N_13513,N_12225,N_12255);
nor U13514 (N_13514,N_13272,N_12711);
or U13515 (N_13515,N_12959,N_12164);
nor U13516 (N_13516,N_12045,N_12091);
xor U13517 (N_13517,N_13285,N_12533);
nor U13518 (N_13518,N_12954,N_13384);
or U13519 (N_13519,N_13224,N_12110);
xnor U13520 (N_13520,N_12757,N_13070);
nand U13521 (N_13521,N_12938,N_12386);
nand U13522 (N_13522,N_12319,N_12382);
or U13523 (N_13523,N_12048,N_12564);
nand U13524 (N_13524,N_12526,N_13026);
or U13525 (N_13525,N_12367,N_12114);
or U13526 (N_13526,N_12310,N_12655);
nand U13527 (N_13527,N_12732,N_13136);
or U13528 (N_13528,N_12301,N_13126);
nor U13529 (N_13529,N_12714,N_12153);
nor U13530 (N_13530,N_12095,N_12669);
or U13531 (N_13531,N_12147,N_13147);
nand U13532 (N_13532,N_12200,N_13228);
and U13533 (N_13533,N_13076,N_13368);
nor U13534 (N_13534,N_13037,N_13370);
nor U13535 (N_13535,N_12359,N_12270);
nand U13536 (N_13536,N_13437,N_13178);
and U13537 (N_13537,N_12432,N_13436);
and U13538 (N_13538,N_12330,N_12828);
nor U13539 (N_13539,N_12589,N_12239);
nor U13540 (N_13540,N_12154,N_12890);
xnor U13541 (N_13541,N_12884,N_13474);
nand U13542 (N_13542,N_13476,N_12149);
nor U13543 (N_13543,N_12298,N_13114);
and U13544 (N_13544,N_12749,N_12824);
and U13545 (N_13545,N_12391,N_12903);
and U13546 (N_13546,N_13260,N_13498);
nor U13547 (N_13547,N_13462,N_13081);
and U13548 (N_13548,N_12447,N_12028);
nor U13549 (N_13549,N_12519,N_13180);
or U13550 (N_13550,N_12313,N_13214);
or U13551 (N_13551,N_12668,N_12934);
nor U13552 (N_13552,N_12217,N_13488);
nor U13553 (N_13553,N_13215,N_12292);
and U13554 (N_13554,N_13458,N_12839);
nor U13555 (N_13555,N_12013,N_12053);
xor U13556 (N_13556,N_12069,N_12582);
xor U13557 (N_13557,N_12872,N_12812);
and U13558 (N_13558,N_12505,N_12222);
nand U13559 (N_13559,N_12761,N_12322);
and U13560 (N_13560,N_12776,N_13455);
or U13561 (N_13561,N_12614,N_13128);
nor U13562 (N_13562,N_13298,N_13068);
nor U13563 (N_13563,N_12573,N_12285);
xnor U13564 (N_13564,N_12510,N_13030);
and U13565 (N_13565,N_12556,N_12034);
nand U13566 (N_13566,N_12652,N_13181);
nand U13567 (N_13567,N_12532,N_13022);
nand U13568 (N_13568,N_12373,N_12978);
and U13569 (N_13569,N_13487,N_12724);
nand U13570 (N_13570,N_13445,N_12883);
nor U13571 (N_13571,N_12616,N_13150);
or U13572 (N_13572,N_13057,N_12945);
xor U13573 (N_13573,N_12770,N_13222);
or U13574 (N_13574,N_12245,N_12809);
nand U13575 (N_13575,N_12312,N_13266);
or U13576 (N_13576,N_12849,N_12554);
xor U13577 (N_13577,N_12356,N_12602);
nand U13578 (N_13578,N_12986,N_12415);
nand U13579 (N_13579,N_13088,N_12414);
and U13580 (N_13580,N_12501,N_12413);
nand U13581 (N_13581,N_12950,N_13041);
or U13582 (N_13582,N_13139,N_12326);
or U13583 (N_13583,N_12102,N_13375);
and U13584 (N_13584,N_13452,N_13051);
and U13585 (N_13585,N_12187,N_12471);
xor U13586 (N_13586,N_13361,N_12644);
nand U13587 (N_13587,N_12705,N_12898);
xnor U13588 (N_13588,N_12317,N_12957);
nand U13589 (N_13589,N_12429,N_12656);
xnor U13590 (N_13590,N_12767,N_12731);
nand U13591 (N_13591,N_12947,N_12097);
nor U13592 (N_13592,N_13376,N_13015);
and U13593 (N_13593,N_12104,N_12900);
nand U13594 (N_13594,N_12891,N_12393);
and U13595 (N_13595,N_12269,N_13159);
and U13596 (N_13596,N_13156,N_12547);
or U13597 (N_13597,N_12930,N_12228);
and U13598 (N_13598,N_12988,N_13130);
nand U13599 (N_13599,N_13393,N_13111);
nor U13600 (N_13600,N_12129,N_12494);
or U13601 (N_13601,N_12975,N_12256);
nor U13602 (N_13602,N_12468,N_13472);
xor U13603 (N_13603,N_13499,N_12160);
or U13604 (N_13604,N_13407,N_13047);
or U13605 (N_13605,N_12161,N_13110);
xor U13606 (N_13606,N_12340,N_13148);
and U13607 (N_13607,N_13466,N_12998);
or U13608 (N_13608,N_12262,N_12846);
xor U13609 (N_13609,N_12569,N_12834);
nor U13610 (N_13610,N_12976,N_13104);
xor U13611 (N_13611,N_12766,N_12831);
and U13612 (N_13612,N_12911,N_12679);
nor U13613 (N_13613,N_12662,N_13197);
nand U13614 (N_13614,N_13480,N_13035);
and U13615 (N_13615,N_12401,N_12605);
xnor U13616 (N_13616,N_12191,N_13300);
nor U13617 (N_13617,N_12787,N_12138);
nand U13618 (N_13618,N_12733,N_13245);
or U13619 (N_13619,N_12005,N_13271);
and U13620 (N_13620,N_12037,N_13240);
nand U13621 (N_13621,N_12880,N_13225);
and U13622 (N_13622,N_13018,N_12933);
xor U13623 (N_13623,N_13170,N_12372);
xnor U13624 (N_13624,N_12212,N_13131);
nand U13625 (N_13625,N_12789,N_12021);
nand U13626 (N_13626,N_13431,N_13288);
or U13627 (N_13627,N_12280,N_12194);
and U13628 (N_13628,N_13188,N_12328);
nor U13629 (N_13629,N_12558,N_12250);
nand U13630 (N_13630,N_12017,N_12964);
nand U13631 (N_13631,N_12075,N_12735);
nor U13632 (N_13632,N_12049,N_13430);
nand U13633 (N_13633,N_13415,N_12719);
nand U13634 (N_13634,N_13161,N_12248);
and U13635 (N_13635,N_13036,N_12738);
and U13636 (N_13636,N_13183,N_12213);
xnor U13637 (N_13637,N_12162,N_13241);
xor U13638 (N_13638,N_12018,N_12113);
xnor U13639 (N_13639,N_12769,N_13014);
or U13640 (N_13640,N_12083,N_12546);
nand U13641 (N_13641,N_13395,N_13117);
nor U13642 (N_13642,N_12543,N_12035);
nor U13643 (N_13643,N_12072,N_12675);
xnor U13644 (N_13644,N_12867,N_13213);
nor U13645 (N_13645,N_12908,N_13157);
nand U13646 (N_13646,N_12932,N_13091);
nand U13647 (N_13647,N_12286,N_13149);
nor U13648 (N_13648,N_12455,N_12741);
or U13649 (N_13649,N_12167,N_12671);
nor U13650 (N_13650,N_12463,N_12708);
or U13651 (N_13651,N_12350,N_12620);
and U13652 (N_13652,N_12297,N_13492);
and U13653 (N_13653,N_13365,N_13059);
or U13654 (N_13654,N_13281,N_12051);
and U13655 (N_13655,N_13009,N_13421);
nor U13656 (N_13656,N_12044,N_13084);
xor U13657 (N_13657,N_12858,N_13282);
nor U13658 (N_13658,N_12640,N_13200);
nor U13659 (N_13659,N_13348,N_12529);
nand U13660 (N_13660,N_13229,N_12765);
nand U13661 (N_13661,N_12196,N_13102);
nor U13662 (N_13662,N_12387,N_13005);
or U13663 (N_13663,N_12970,N_12520);
nor U13664 (N_13664,N_13324,N_13297);
nand U13665 (N_13665,N_12365,N_13082);
and U13666 (N_13666,N_13001,N_12331);
nor U13667 (N_13667,N_13302,N_13287);
and U13668 (N_13668,N_12647,N_13244);
or U13669 (N_13669,N_12060,N_12531);
xnor U13670 (N_13670,N_12188,N_12008);
and U13671 (N_13671,N_12628,N_12728);
nand U13672 (N_13672,N_12779,N_12666);
or U13673 (N_13673,N_12445,N_13294);
xor U13674 (N_13674,N_12944,N_13173);
xor U13675 (N_13675,N_12031,N_12878);
xnor U13676 (N_13676,N_12337,N_12555);
xor U13677 (N_13677,N_12023,N_12026);
or U13678 (N_13678,N_12958,N_12922);
nand U13679 (N_13679,N_13179,N_13249);
xor U13680 (N_13680,N_13337,N_12462);
or U13681 (N_13681,N_13329,N_12452);
and U13682 (N_13682,N_12388,N_12363);
nor U13683 (N_13683,N_12946,N_12132);
and U13684 (N_13684,N_12660,N_12253);
and U13685 (N_13685,N_12702,N_12124);
nand U13686 (N_13686,N_13098,N_12430);
xor U13687 (N_13687,N_12107,N_12249);
nand U13688 (N_13688,N_12865,N_13099);
xnor U13689 (N_13689,N_12506,N_12901);
xnor U13690 (N_13690,N_13343,N_12346);
nand U13691 (N_13691,N_12973,N_12426);
and U13692 (N_13692,N_12683,N_12392);
xnor U13693 (N_13693,N_13406,N_12477);
xnor U13694 (N_13694,N_12804,N_13203);
or U13695 (N_13695,N_12498,N_12033);
and U13696 (N_13696,N_12536,N_12693);
and U13697 (N_13697,N_12276,N_12838);
nand U13698 (N_13698,N_13394,N_12324);
xnor U13699 (N_13699,N_13304,N_12175);
nor U13700 (N_13700,N_12806,N_12145);
nand U13701 (N_13701,N_12994,N_12420);
and U13702 (N_13702,N_12739,N_12659);
nor U13703 (N_13703,N_12720,N_12349);
or U13704 (N_13704,N_12295,N_12389);
and U13705 (N_13705,N_13118,N_12856);
nand U13706 (N_13706,N_12151,N_12985);
nor U13707 (N_13707,N_12619,N_13290);
xnor U13708 (N_13708,N_13109,N_13032);
xor U13709 (N_13709,N_13345,N_12822);
or U13710 (N_13710,N_12261,N_12300);
and U13711 (N_13711,N_12299,N_13079);
xnor U13712 (N_13712,N_13083,N_13247);
or U13713 (N_13713,N_13105,N_13494);
xor U13714 (N_13714,N_12692,N_12265);
nor U13715 (N_13715,N_12586,N_13112);
nand U13716 (N_13716,N_12074,N_12886);
or U13717 (N_13717,N_12635,N_13469);
and U13718 (N_13718,N_12530,N_12150);
and U13719 (N_13719,N_13325,N_13023);
nand U13720 (N_13720,N_13177,N_12137);
xnor U13721 (N_13721,N_12159,N_12036);
or U13722 (N_13722,N_13253,N_12544);
nand U13723 (N_13723,N_13311,N_12704);
xor U13724 (N_13724,N_12820,N_13291);
or U13725 (N_13725,N_12718,N_12246);
nand U13726 (N_13726,N_13264,N_12928);
or U13727 (N_13727,N_12351,N_13400);
and U13728 (N_13728,N_13425,N_12918);
and U13729 (N_13729,N_12314,N_12525);
nor U13730 (N_13730,N_12603,N_13061);
or U13731 (N_13731,N_12198,N_13024);
nor U13732 (N_13732,N_12370,N_12700);
or U13733 (N_13733,N_13449,N_12009);
or U13734 (N_13734,N_12362,N_12682);
or U13735 (N_13735,N_12513,N_12271);
xor U13736 (N_13736,N_13333,N_12862);
and U13737 (N_13737,N_12534,N_13419);
xnor U13738 (N_13738,N_12813,N_13349);
and U13739 (N_13739,N_12949,N_12797);
or U13740 (N_13740,N_13243,N_12987);
and U13741 (N_13741,N_12354,N_13490);
and U13742 (N_13742,N_12966,N_12518);
or U13743 (N_13743,N_13378,N_13184);
nand U13744 (N_13744,N_12054,N_12829);
nand U13745 (N_13745,N_12006,N_12484);
or U13746 (N_13746,N_12277,N_12570);
xor U13747 (N_13747,N_12565,N_13199);
or U13748 (N_13748,N_12642,N_12951);
xor U13749 (N_13749,N_12606,N_12979);
or U13750 (N_13750,N_12968,N_12868);
nand U13751 (N_13751,N_12219,N_12119);
or U13752 (N_13752,N_13473,N_12991);
nor U13753 (N_13753,N_12487,N_12716);
or U13754 (N_13754,N_12041,N_13404);
xor U13755 (N_13755,N_12764,N_12254);
nor U13756 (N_13756,N_12011,N_12892);
and U13757 (N_13757,N_13450,N_13048);
xnor U13758 (N_13758,N_12407,N_12844);
or U13759 (N_13759,N_13386,N_12783);
and U13760 (N_13760,N_12238,N_12293);
and U13761 (N_13761,N_13192,N_13232);
and U13762 (N_13762,N_13497,N_12090);
nor U13763 (N_13763,N_13465,N_12101);
nand U13764 (N_13764,N_13468,N_13003);
or U13765 (N_13765,N_13467,N_12791);
nand U13766 (N_13766,N_12752,N_12740);
or U13767 (N_13767,N_12768,N_12989);
nand U13768 (N_13768,N_13399,N_13137);
nand U13769 (N_13769,N_12889,N_13134);
nor U13770 (N_13770,N_12476,N_12121);
nor U13771 (N_13771,N_12087,N_13133);
nand U13772 (N_13772,N_12550,N_13382);
or U13773 (N_13773,N_12073,N_13350);
and U13774 (N_13774,N_12877,N_13427);
or U13775 (N_13775,N_13416,N_12627);
or U13776 (N_13776,N_12172,N_13422);
or U13777 (N_13777,N_13187,N_12168);
xor U13778 (N_13778,N_12542,N_13176);
xnor U13779 (N_13779,N_13326,N_12698);
nor U13780 (N_13780,N_13080,N_12940);
xnor U13781 (N_13781,N_12843,N_12885);
and U13782 (N_13782,N_13231,N_12327);
and U13783 (N_13783,N_13040,N_12371);
and U13784 (N_13784,N_13043,N_12524);
nand U13785 (N_13785,N_12144,N_12869);
nand U13786 (N_13786,N_12472,N_12674);
xnor U13787 (N_13787,N_12962,N_12438);
and U13788 (N_13788,N_13234,N_12805);
or U13789 (N_13789,N_13265,N_13408);
and U13790 (N_13790,N_12252,N_12268);
nand U13791 (N_13791,N_12795,N_12631);
nand U13792 (N_13792,N_12706,N_12123);
nand U13793 (N_13793,N_12552,N_13489);
or U13794 (N_13794,N_12624,N_12093);
xnor U13795 (N_13795,N_12961,N_12112);
or U13796 (N_13796,N_12197,N_12587);
xnor U13797 (N_13797,N_12177,N_12406);
xnor U13798 (N_13798,N_13191,N_12808);
xnor U13799 (N_13799,N_13056,N_12667);
nor U13800 (N_13800,N_12777,N_13064);
xnor U13801 (N_13801,N_12007,N_12052);
nand U13802 (N_13802,N_12439,N_13078);
nor U13803 (N_13803,N_12306,N_13323);
xnor U13804 (N_13804,N_12729,N_12459);
nand U13805 (N_13805,N_13162,N_12133);
xnor U13806 (N_13806,N_12592,N_12341);
nor U13807 (N_13807,N_12431,N_13089);
nor U13808 (N_13808,N_12399,N_12135);
xnor U13809 (N_13809,N_13223,N_12279);
and U13810 (N_13810,N_12338,N_12836);
nand U13811 (N_13811,N_13280,N_13146);
or U13812 (N_13812,N_12909,N_13309);
or U13813 (N_13813,N_13461,N_12830);
nor U13814 (N_13814,N_12636,N_12062);
nand U13815 (N_13815,N_12456,N_12851);
nor U13816 (N_13816,N_13097,N_12881);
and U13817 (N_13817,N_12888,N_12166);
or U13818 (N_13818,N_12444,N_12260);
or U13819 (N_13819,N_13052,N_12325);
nor U13820 (N_13820,N_12527,N_12709);
and U13821 (N_13821,N_13357,N_12854);
nand U13822 (N_13822,N_12068,N_13012);
and U13823 (N_13823,N_13107,N_13336);
or U13824 (N_13824,N_12515,N_12567);
and U13825 (N_13825,N_13226,N_12971);
or U13826 (N_13826,N_12015,N_13113);
xor U13827 (N_13827,N_12014,N_13276);
and U13828 (N_13828,N_13346,N_12377);
nand U13829 (N_13829,N_12503,N_12850);
nand U13830 (N_13830,N_12697,N_13250);
nor U13831 (N_13831,N_13209,N_13259);
or U13832 (N_13832,N_12321,N_12493);
nand U13833 (N_13833,N_12591,N_12082);
or U13834 (N_13834,N_13058,N_13295);
xor U13835 (N_13835,N_13219,N_12189);
and U13836 (N_13836,N_12304,N_12722);
nor U13837 (N_13837,N_13478,N_12193);
nor U13838 (N_13838,N_12220,N_12939);
nand U13839 (N_13839,N_13206,N_12274);
or U13840 (N_13840,N_12423,N_13355);
and U13841 (N_13841,N_12027,N_12109);
nor U13842 (N_13842,N_12980,N_12247);
nand U13843 (N_13843,N_13366,N_12233);
nand U13844 (N_13844,N_13444,N_12593);
nor U13845 (N_13845,N_12024,N_12383);
and U13846 (N_13846,N_12848,N_12875);
xor U13847 (N_13847,N_13447,N_12173);
nand U13848 (N_13848,N_12678,N_12290);
xor U13849 (N_13849,N_12726,N_13432);
xnor U13850 (N_13850,N_12223,N_13257);
xor U13851 (N_13851,N_12861,N_13420);
and U13852 (N_13852,N_12019,N_12915);
nor U13853 (N_13853,N_12897,N_13060);
nor U13854 (N_13854,N_12925,N_12288);
nor U13855 (N_13855,N_13426,N_12169);
or U13856 (N_13856,N_12491,N_12977);
xnor U13857 (N_13857,N_12466,N_12760);
xnor U13858 (N_13858,N_12369,N_13320);
nor U13859 (N_13859,N_12342,N_12514);
and U13860 (N_13860,N_13208,N_12334);
and U13861 (N_13861,N_12066,N_12641);
or U13862 (N_13862,N_13354,N_12264);
xnor U13863 (N_13863,N_12863,N_13486);
xor U13864 (N_13864,N_12874,N_12793);
or U13865 (N_13865,N_13074,N_13409);
xnor U13866 (N_13866,N_12899,N_12816);
xor U13867 (N_13867,N_13453,N_13062);
xnor U13868 (N_13868,N_12786,N_12106);
nand U13869 (N_13869,N_12818,N_13402);
and U13870 (N_13870,N_13085,N_12237);
and U13871 (N_13871,N_12557,N_12411);
xnor U13872 (N_13872,N_12100,N_12105);
nand U13873 (N_13873,N_12384,N_12996);
and U13874 (N_13874,N_13207,N_12782);
xor U13875 (N_13875,N_12479,N_13353);
nand U13876 (N_13876,N_13202,N_12645);
nor U13877 (N_13877,N_12483,N_12545);
nand U13878 (N_13878,N_12012,N_12381);
nor U13879 (N_13879,N_13362,N_12042);
and U13880 (N_13880,N_12664,N_12376);
or U13881 (N_13881,N_13189,N_13115);
or U13882 (N_13882,N_12549,N_12136);
nor U13883 (N_13883,N_12296,N_12676);
and U13884 (N_13884,N_12873,N_12584);
nor U13885 (N_13885,N_13417,N_13172);
nor U13886 (N_13886,N_13356,N_12730);
xor U13887 (N_13887,N_12418,N_13360);
or U13888 (N_13888,N_12663,N_13190);
and U13889 (N_13889,N_12919,N_12202);
xor U13890 (N_13890,N_12409,N_12753);
xor U13891 (N_13891,N_12344,N_13477);
nand U13892 (N_13892,N_12229,N_12917);
and U13893 (N_13893,N_12002,N_13021);
nor U13894 (N_13894,N_13459,N_12611);
or U13895 (N_13895,N_12574,N_13069);
nand U13896 (N_13896,N_12819,N_12071);
or U13897 (N_13897,N_13484,N_12500);
nor U13898 (N_13898,N_12499,N_13479);
or U13899 (N_13899,N_12067,N_13075);
nand U13900 (N_13900,N_12302,N_12802);
and U13901 (N_13901,N_12092,N_13155);
or U13902 (N_13902,N_12241,N_12522);
or U13903 (N_13903,N_12379,N_12785);
nand U13904 (N_13904,N_12427,N_13013);
nor U13905 (N_13905,N_13334,N_12568);
xnor U13906 (N_13906,N_12983,N_12470);
and U13907 (N_13907,N_12896,N_13359);
nor U13908 (N_13908,N_12163,N_12879);
and U13909 (N_13909,N_12712,N_12030);
and U13910 (N_13910,N_13296,N_13090);
xnor U13911 (N_13911,N_12778,N_12598);
nor U13912 (N_13912,N_12999,N_13204);
nand U13913 (N_13913,N_12453,N_12440);
and U13914 (N_13914,N_12864,N_12099);
nor U13915 (N_13915,N_13316,N_13168);
or U13916 (N_13916,N_12355,N_13380);
or U13917 (N_13917,N_12981,N_12581);
xnor U13918 (N_13918,N_12303,N_12451);
or U13919 (N_13919,N_12590,N_13347);
nor U13920 (N_13920,N_13166,N_12118);
xor U13921 (N_13921,N_12358,N_12774);
nor U13922 (N_13922,N_12128,N_13195);
nor U13923 (N_13923,N_12853,N_13293);
and U13924 (N_13924,N_12771,N_12583);
or U13925 (N_13925,N_12174,N_13185);
nor U13926 (N_13926,N_12639,N_12405);
nand U13927 (N_13927,N_12743,N_12242);
nor U13928 (N_13928,N_13094,N_13143);
and U13929 (N_13929,N_13418,N_12308);
nand U13930 (N_13930,N_12230,N_13121);
xnor U13931 (N_13931,N_12204,N_13433);
and U13932 (N_13932,N_12195,N_12906);
nand U13933 (N_13933,N_12857,N_13194);
or U13934 (N_13934,N_12870,N_13086);
nand U13935 (N_13935,N_13008,N_12117);
or U13936 (N_13936,N_13025,N_12615);
nor U13937 (N_13937,N_12366,N_12142);
nand U13938 (N_13938,N_13303,N_12199);
and U13939 (N_13939,N_12993,N_12116);
xor U13940 (N_13940,N_12004,N_13328);
and U13941 (N_13941,N_13065,N_12375);
xor U13942 (N_13942,N_12604,N_12412);
and U13943 (N_13943,N_12953,N_12650);
xnor U13944 (N_13944,N_13038,N_12390);
or U13945 (N_13945,N_12224,N_13205);
and U13946 (N_13946,N_13413,N_13438);
or U13947 (N_13947,N_12461,N_12206);
and U13948 (N_13948,N_12969,N_13135);
nand U13949 (N_13949,N_12275,N_12032);
or U13950 (N_13950,N_12156,N_12311);
nor U13951 (N_13951,N_12929,N_12579);
xor U13952 (N_13952,N_12715,N_12673);
xnor U13953 (N_13953,N_12096,N_12378);
xor U13954 (N_13954,N_12385,N_13031);
nand U13955 (N_13955,N_12665,N_12357);
nand U13956 (N_13956,N_12772,N_12841);
nor U13957 (N_13957,N_13122,N_13258);
xnor U13958 (N_13958,N_12205,N_12921);
nor U13959 (N_13959,N_12832,N_13154);
nor U13960 (N_13960,N_12677,N_13125);
and U13961 (N_13961,N_13267,N_12907);
nor U13962 (N_13962,N_13481,N_12600);
and U13963 (N_13963,N_12089,N_13138);
or U13964 (N_13964,N_12185,N_13218);
xor U13965 (N_13965,N_13401,N_12685);
nor U13966 (N_13966,N_12203,N_12638);
and U13967 (N_13967,N_13451,N_13363);
or U13968 (N_13968,N_12625,N_12654);
nand U13969 (N_13969,N_12022,N_13096);
or U13970 (N_13970,N_13002,N_12535);
nor U13971 (N_13971,N_12762,N_12422);
nand U13972 (N_13972,N_12686,N_12360);
and U13973 (N_13973,N_12226,N_12454);
nor U13974 (N_13974,N_12974,N_12394);
nand U13975 (N_13975,N_12287,N_12486);
nor U13976 (N_13976,N_13314,N_12281);
nand U13977 (N_13977,N_12473,N_12895);
and U13978 (N_13978,N_12955,N_12207);
and U13979 (N_13979,N_12070,N_13305);
xnor U13980 (N_13980,N_13446,N_12621);
nand U13981 (N_13981,N_12601,N_13318);
nand U13982 (N_13982,N_12043,N_12347);
and U13983 (N_13983,N_12474,N_13153);
or U13984 (N_13984,N_12201,N_13095);
and U13985 (N_13985,N_13246,N_12397);
xnor U13986 (N_13986,N_12643,N_13388);
xor U13987 (N_13987,N_12563,N_13017);
or U13988 (N_13988,N_12380,N_12781);
and U13989 (N_13989,N_13278,N_12859);
nor U13990 (N_13990,N_13440,N_12294);
nor U13991 (N_13991,N_13164,N_12125);
nand U13992 (N_13992,N_12784,N_12622);
or U13993 (N_13993,N_12039,N_12634);
xnor U13994 (N_13994,N_12658,N_12773);
and U13995 (N_13995,N_13471,N_12553);
or U13996 (N_13996,N_13108,N_13106);
xnor U13997 (N_13997,N_12258,N_12184);
nand U13998 (N_13998,N_13383,N_12694);
nor U13999 (N_13999,N_12717,N_13315);
xor U14000 (N_14000,N_12218,N_12755);
or U14001 (N_14001,N_12815,N_13396);
nor U14002 (N_14002,N_13174,N_13352);
or U14003 (N_14003,N_12443,N_12855);
nor U14004 (N_14004,N_12103,N_12434);
nand U14005 (N_14005,N_12227,N_12489);
or U14006 (N_14006,N_13321,N_13405);
xnor U14007 (N_14007,N_12259,N_13275);
and U14008 (N_14008,N_12657,N_13252);
nor U14009 (N_14009,N_13124,N_12141);
and U14010 (N_14010,N_12588,N_13340);
or U14011 (N_14011,N_12063,N_13236);
nand U14012 (N_14012,N_13423,N_12329);
nor U14013 (N_14013,N_13439,N_13270);
and U14014 (N_14014,N_12345,N_13010);
and U14015 (N_14015,N_12038,N_12725);
and U14016 (N_14016,N_12395,N_13456);
and U14017 (N_14017,N_12629,N_12924);
nor U14018 (N_14018,N_13358,N_13167);
nand U14019 (N_14019,N_13284,N_12307);
nand U14020 (N_14020,N_12578,N_12610);
nand U14021 (N_14021,N_13331,N_12272);
or U14022 (N_14022,N_12887,N_13344);
xor U14023 (N_14023,N_12942,N_13341);
nor U14024 (N_14024,N_13387,N_13367);
xnor U14025 (N_14025,N_12010,N_12561);
or U14026 (N_14026,N_12649,N_12143);
xor U14027 (N_14027,N_12400,N_13371);
nand U14028 (N_14028,N_12687,N_12084);
xnor U14029 (N_14029,N_13000,N_13310);
xnor U14030 (N_14030,N_13101,N_12963);
nor U14031 (N_14031,N_12403,N_12798);
xnor U14032 (N_14032,N_12441,N_12936);
xnor U14033 (N_14033,N_12231,N_13448);
xor U14034 (N_14034,N_12790,N_12127);
and U14035 (N_14035,N_13301,N_12361);
xor U14036 (N_14036,N_13491,N_12165);
nor U14037 (N_14037,N_13019,N_12992);
nand U14038 (N_14038,N_13119,N_12585);
xor U14039 (N_14039,N_12847,N_12352);
nand U14040 (N_14040,N_13141,N_12827);
nand U14041 (N_14041,N_13201,N_12449);
nand U14042 (N_14042,N_12211,N_12480);
xor U14043 (N_14043,N_13286,N_12758);
nand U14044 (N_14044,N_13342,N_12548);
or U14045 (N_14045,N_12368,N_13374);
nand U14046 (N_14046,N_12713,N_12982);
nor U14047 (N_14047,N_12433,N_13210);
nor U14048 (N_14048,N_12339,N_13392);
xnor U14049 (N_14049,N_12689,N_12801);
and U14050 (N_14050,N_12064,N_12670);
nor U14051 (N_14051,N_13351,N_13410);
xor U14052 (N_14052,N_13335,N_13483);
nor U14053 (N_14053,N_12826,N_12178);
nand U14054 (N_14054,N_12047,N_12232);
xnor U14055 (N_14055,N_13251,N_12823);
or U14056 (N_14056,N_12931,N_12003);
nor U14057 (N_14057,N_12866,N_12284);
and U14058 (N_14058,N_12496,N_12699);
xnor U14059 (N_14059,N_12577,N_12504);
nor U14060 (N_14060,N_12613,N_13434);
nand U14061 (N_14061,N_13145,N_12840);
nand U14062 (N_14062,N_12478,N_12428);
nor U14063 (N_14063,N_12457,N_12158);
xnor U14064 (N_14064,N_12408,N_12257);
nor U14065 (N_14065,N_13063,N_12140);
and U14066 (N_14066,N_12952,N_12902);
or U14067 (N_14067,N_12079,N_13443);
or U14068 (N_14068,N_13319,N_12509);
nand U14069 (N_14069,N_13235,N_12335);
and U14070 (N_14070,N_13317,N_12814);
nor U14071 (N_14071,N_12122,N_12748);
xor U14072 (N_14072,N_13364,N_12404);
or U14073 (N_14073,N_12183,N_13306);
or U14074 (N_14074,N_12208,N_12278);
and U14075 (N_14075,N_13165,N_13274);
nor U14076 (N_14076,N_13239,N_12111);
or U14077 (N_14077,N_12910,N_13464);
and U14078 (N_14078,N_12436,N_12599);
xnor U14079 (N_14079,N_12176,N_13277);
or U14080 (N_14080,N_12221,N_13230);
nand U14081 (N_14081,N_12575,N_12282);
nand U14082 (N_14082,N_12315,N_12216);
or U14083 (N_14083,N_13261,N_12029);
xnor U14084 (N_14084,N_12742,N_12691);
and U14085 (N_14085,N_13175,N_13007);
xnor U14086 (N_14086,N_12323,N_12821);
xnor U14087 (N_14087,N_12469,N_12155);
nor U14088 (N_14088,N_12746,N_12157);
or U14089 (N_14089,N_13033,N_12721);
nand U14090 (N_14090,N_12754,N_13186);
and U14091 (N_14091,N_12633,N_12680);
or U14092 (N_14092,N_13398,N_13269);
or U14093 (N_14093,N_12240,N_12759);
xor U14094 (N_14094,N_13470,N_12289);
nor U14095 (N_14095,N_13132,N_13379);
and U14096 (N_14096,N_12695,N_13390);
and U14097 (N_14097,N_13460,N_12465);
and U14098 (N_14098,N_13053,N_13493);
nand U14099 (N_14099,N_12528,N_12065);
and U14100 (N_14100,N_12424,N_12080);
nor U14101 (N_14101,N_13242,N_13054);
and U14102 (N_14102,N_13255,N_12333);
nand U14103 (N_14103,N_12495,N_12537);
and U14104 (N_14104,N_13496,N_13313);
xnor U14105 (N_14105,N_12912,N_12597);
nand U14106 (N_14106,N_12508,N_12481);
and U14107 (N_14107,N_12115,N_12871);
nand U14108 (N_14108,N_12796,N_13067);
and U14109 (N_14109,N_13254,N_13279);
xnor U14110 (N_14110,N_12727,N_12251);
and U14111 (N_14111,N_12630,N_12332);
or U14112 (N_14112,N_12171,N_13389);
and U14113 (N_14113,N_13273,N_12538);
or U14114 (N_14114,N_12842,N_12935);
xnor U14115 (N_14115,N_12833,N_12681);
and U14116 (N_14116,N_12937,N_12914);
or U14117 (N_14117,N_12882,N_12056);
nand U14118 (N_14118,N_12617,N_12417);
nor U14119 (N_14119,N_13045,N_12305);
and U14120 (N_14120,N_12707,N_12965);
nand U14121 (N_14121,N_13412,N_12571);
nor U14122 (N_14122,N_13073,N_12402);
xnor U14123 (N_14123,N_13308,N_12566);
or U14124 (N_14124,N_12632,N_12098);
nand U14125 (N_14125,N_13029,N_13424);
and U14126 (N_14126,N_12559,N_12637);
nand U14127 (N_14127,N_12348,N_12523);
nor U14128 (N_14128,N_12684,N_12608);
nand U14129 (N_14129,N_12215,N_13332);
nor U14130 (N_14130,N_13071,N_12085);
and U14131 (N_14131,N_12179,N_12756);
nand U14132 (N_14132,N_13006,N_13151);
xnor U14133 (N_14133,N_13196,N_12997);
or U14134 (N_14134,N_12120,N_12852);
nand U14135 (N_14135,N_12181,N_12594);
nand U14136 (N_14136,N_12309,N_12551);
and U14137 (N_14137,N_12794,N_12607);
and U14138 (N_14138,N_12775,N_12894);
xnor U14139 (N_14139,N_12016,N_12984);
or U14140 (N_14140,N_12182,N_12214);
nor U14141 (N_14141,N_12835,N_13369);
nand U14142 (N_14142,N_12152,N_12926);
nor U14143 (N_14143,N_13077,N_13221);
and U14144 (N_14144,N_13482,N_12736);
and U14145 (N_14145,N_12572,N_12661);
nor U14146 (N_14146,N_12927,N_13327);
or U14147 (N_14147,N_12653,N_13414);
and U14148 (N_14148,N_12623,N_12139);
and U14149 (N_14149,N_13169,N_12267);
nor U14150 (N_14150,N_12192,N_12893);
or U14151 (N_14151,N_12088,N_12131);
and U14152 (N_14152,N_13028,N_13212);
or U14153 (N_14153,N_12609,N_13103);
or U14154 (N_14154,N_12734,N_12723);
and U14155 (N_14155,N_13042,N_12488);
nor U14156 (N_14156,N_13198,N_13475);
nor U14157 (N_14157,N_12467,N_13233);
nand U14158 (N_14158,N_12803,N_12904);
nand U14159 (N_14159,N_13442,N_12448);
and U14160 (N_14160,N_13227,N_12050);
nand U14161 (N_14161,N_12421,N_12475);
or U14162 (N_14162,N_12316,N_12497);
xor U14163 (N_14163,N_13072,N_13039);
nand U14164 (N_14164,N_12318,N_12458);
nor U14165 (N_14165,N_12059,N_13158);
nor U14166 (N_14166,N_13237,N_12612);
and U14167 (N_14167,N_12046,N_12364);
nor U14168 (N_14168,N_12320,N_12817);
or U14169 (N_14169,N_12648,N_12000);
and U14170 (N_14170,N_13049,N_12450);
or U14171 (N_14171,N_12967,N_12646);
nor U14172 (N_14172,N_12266,N_12180);
and U14173 (N_14173,N_13263,N_13127);
xnor U14174 (N_14174,N_12078,N_12398);
or U14175 (N_14175,N_12076,N_12788);
xor U14176 (N_14176,N_13403,N_12492);
or U14177 (N_14177,N_12108,N_13373);
and U14178 (N_14178,N_12800,N_13238);
nor U14179 (N_14179,N_12511,N_12860);
nand U14180 (N_14180,N_12190,N_12236);
nor U14181 (N_14181,N_12396,N_13411);
xor U14182 (N_14182,N_12837,N_12148);
xnor U14183 (N_14183,N_12263,N_12482);
and U14184 (N_14184,N_12810,N_13055);
and U14185 (N_14185,N_12512,N_13485);
nor U14186 (N_14186,N_12972,N_13171);
and U14187 (N_14187,N_13441,N_12737);
and U14188 (N_14188,N_13322,N_12562);
or U14189 (N_14189,N_12744,N_12146);
and U14190 (N_14190,N_13289,N_13093);
or U14191 (N_14191,N_12905,N_12916);
nor U14192 (N_14192,N_13330,N_12696);
or U14193 (N_14193,N_13268,N_13092);
nor U14194 (N_14194,N_13027,N_13435);
xnor U14195 (N_14195,N_13457,N_12539);
or U14196 (N_14196,N_12134,N_12913);
or U14197 (N_14197,N_12701,N_13262);
and U14198 (N_14198,N_13016,N_12435);
xnor U14199 (N_14199,N_13463,N_12948);
nand U14200 (N_14200,N_12502,N_12057);
or U14201 (N_14201,N_13142,N_13299);
or U14202 (N_14202,N_12576,N_12690);
xor U14203 (N_14203,N_13193,N_12845);
nor U14204 (N_14204,N_13495,N_12751);
nand U14205 (N_14205,N_12081,N_12920);
nand U14206 (N_14206,N_12210,N_12442);
or U14207 (N_14207,N_13256,N_12596);
nand U14208 (N_14208,N_12273,N_13377);
or U14209 (N_14209,N_12086,N_12745);
nand U14210 (N_14210,N_12464,N_12283);
xnor U14211 (N_14211,N_12541,N_12876);
xor U14212 (N_14212,N_12186,N_12580);
and U14213 (N_14213,N_12025,N_13391);
xnor U14214 (N_14214,N_13160,N_12960);
and U14215 (N_14215,N_12780,N_12353);
nor U14216 (N_14216,N_12799,N_12990);
nand U14217 (N_14217,N_12618,N_12807);
or U14218 (N_14218,N_13292,N_12995);
nor U14219 (N_14219,N_13034,N_13020);
and U14220 (N_14220,N_12651,N_13338);
and U14221 (N_14221,N_12747,N_13216);
nand U14222 (N_14222,N_12061,N_13120);
and U14223 (N_14223,N_13123,N_13217);
nand U14224 (N_14224,N_12243,N_12130);
xnor U14225 (N_14225,N_13044,N_13144);
or U14226 (N_14226,N_12170,N_13381);
or U14227 (N_14227,N_12336,N_12710);
and U14228 (N_14228,N_12094,N_12410);
nor U14229 (N_14229,N_12485,N_12416);
xnor U14230 (N_14230,N_13454,N_13129);
and U14231 (N_14231,N_13248,N_12560);
nor U14232 (N_14232,N_12943,N_12020);
xor U14233 (N_14233,N_12703,N_12941);
nor U14234 (N_14234,N_12750,N_13372);
or U14235 (N_14235,N_12234,N_13397);
or U14236 (N_14236,N_13429,N_13066);
or U14237 (N_14237,N_13140,N_12517);
nand U14238 (N_14238,N_12437,N_12792);
or U14239 (N_14239,N_13163,N_12235);
or U14240 (N_14240,N_12419,N_12521);
nor U14241 (N_14241,N_12595,N_12763);
nand U14242 (N_14242,N_12688,N_13050);
and U14243 (N_14243,N_13011,N_13004);
or U14244 (N_14244,N_12291,N_12077);
xor U14245 (N_14245,N_12626,N_12001);
or U14246 (N_14246,N_13182,N_12209);
xor U14247 (N_14247,N_12811,N_12923);
xnor U14248 (N_14248,N_12516,N_12040);
or U14249 (N_14249,N_13100,N_13087);
nor U14250 (N_14250,N_12704,N_12673);
nor U14251 (N_14251,N_12730,N_12196);
nor U14252 (N_14252,N_12240,N_13191);
or U14253 (N_14253,N_12571,N_12714);
nor U14254 (N_14254,N_13490,N_13031);
nor U14255 (N_14255,N_12040,N_13416);
xnor U14256 (N_14256,N_12267,N_12836);
or U14257 (N_14257,N_12234,N_13436);
or U14258 (N_14258,N_12356,N_12933);
nor U14259 (N_14259,N_12156,N_13312);
and U14260 (N_14260,N_13267,N_12045);
xnor U14261 (N_14261,N_12566,N_12141);
or U14262 (N_14262,N_12087,N_12805);
nand U14263 (N_14263,N_13385,N_13388);
or U14264 (N_14264,N_12975,N_13372);
or U14265 (N_14265,N_12543,N_12376);
xnor U14266 (N_14266,N_12867,N_12455);
xor U14267 (N_14267,N_12309,N_13126);
and U14268 (N_14268,N_12799,N_12124);
and U14269 (N_14269,N_13149,N_13214);
or U14270 (N_14270,N_12164,N_12404);
nand U14271 (N_14271,N_13431,N_12607);
and U14272 (N_14272,N_12525,N_12742);
or U14273 (N_14273,N_12856,N_12635);
or U14274 (N_14274,N_13494,N_13117);
and U14275 (N_14275,N_13326,N_13368);
xnor U14276 (N_14276,N_12415,N_13299);
nor U14277 (N_14277,N_13388,N_12779);
and U14278 (N_14278,N_13027,N_12997);
and U14279 (N_14279,N_13271,N_13267);
nand U14280 (N_14280,N_13365,N_12938);
nand U14281 (N_14281,N_12267,N_13132);
nand U14282 (N_14282,N_12701,N_12612);
xor U14283 (N_14283,N_12100,N_12540);
or U14284 (N_14284,N_13215,N_12969);
nor U14285 (N_14285,N_12264,N_13067);
or U14286 (N_14286,N_12928,N_12449);
or U14287 (N_14287,N_13256,N_12942);
xnor U14288 (N_14288,N_13471,N_13122);
nor U14289 (N_14289,N_12267,N_12997);
xnor U14290 (N_14290,N_12487,N_13177);
and U14291 (N_14291,N_13274,N_12267);
xor U14292 (N_14292,N_13400,N_12720);
nand U14293 (N_14293,N_12850,N_12124);
xnor U14294 (N_14294,N_12828,N_13143);
nor U14295 (N_14295,N_13414,N_12110);
and U14296 (N_14296,N_12056,N_13497);
and U14297 (N_14297,N_12213,N_12133);
xor U14298 (N_14298,N_12981,N_13390);
nor U14299 (N_14299,N_12197,N_12929);
nand U14300 (N_14300,N_12506,N_12200);
nor U14301 (N_14301,N_12168,N_13320);
xnor U14302 (N_14302,N_12349,N_12852);
and U14303 (N_14303,N_12198,N_12153);
or U14304 (N_14304,N_12913,N_12269);
and U14305 (N_14305,N_13291,N_12310);
or U14306 (N_14306,N_12854,N_13266);
nor U14307 (N_14307,N_13222,N_12030);
or U14308 (N_14308,N_12702,N_13449);
nand U14309 (N_14309,N_12124,N_13376);
and U14310 (N_14310,N_12196,N_12763);
nand U14311 (N_14311,N_13119,N_12660);
or U14312 (N_14312,N_12082,N_12908);
or U14313 (N_14313,N_12286,N_12092);
xor U14314 (N_14314,N_12267,N_12150);
or U14315 (N_14315,N_12700,N_13358);
xor U14316 (N_14316,N_12537,N_12517);
or U14317 (N_14317,N_12201,N_13066);
xor U14318 (N_14318,N_12792,N_12789);
nor U14319 (N_14319,N_12971,N_12693);
or U14320 (N_14320,N_12258,N_13252);
or U14321 (N_14321,N_12576,N_13033);
or U14322 (N_14322,N_12081,N_13295);
and U14323 (N_14323,N_12958,N_12268);
or U14324 (N_14324,N_13118,N_13039);
and U14325 (N_14325,N_12222,N_13372);
nor U14326 (N_14326,N_12489,N_13074);
and U14327 (N_14327,N_12686,N_12349);
and U14328 (N_14328,N_12073,N_13053);
nand U14329 (N_14329,N_12440,N_12114);
nor U14330 (N_14330,N_12926,N_12948);
and U14331 (N_14331,N_12976,N_13156);
xor U14332 (N_14332,N_12418,N_12542);
or U14333 (N_14333,N_12261,N_12527);
and U14334 (N_14334,N_12149,N_12350);
nor U14335 (N_14335,N_12656,N_13441);
nand U14336 (N_14336,N_12440,N_12038);
nor U14337 (N_14337,N_13064,N_12364);
or U14338 (N_14338,N_13156,N_12942);
nand U14339 (N_14339,N_12861,N_12209);
nand U14340 (N_14340,N_12663,N_12095);
and U14341 (N_14341,N_12778,N_13464);
nand U14342 (N_14342,N_12383,N_12540);
nand U14343 (N_14343,N_13308,N_13384);
nor U14344 (N_14344,N_12139,N_12253);
or U14345 (N_14345,N_12749,N_12247);
nand U14346 (N_14346,N_12525,N_12485);
nor U14347 (N_14347,N_12201,N_13491);
nand U14348 (N_14348,N_13301,N_13232);
and U14349 (N_14349,N_13272,N_12029);
and U14350 (N_14350,N_12432,N_12574);
nand U14351 (N_14351,N_13092,N_12163);
nor U14352 (N_14352,N_12223,N_12323);
nor U14353 (N_14353,N_13019,N_12760);
nor U14354 (N_14354,N_13482,N_12912);
or U14355 (N_14355,N_13056,N_13000);
and U14356 (N_14356,N_12609,N_12885);
xnor U14357 (N_14357,N_13242,N_13009);
nor U14358 (N_14358,N_12702,N_12172);
and U14359 (N_14359,N_12868,N_13333);
xor U14360 (N_14360,N_12105,N_12951);
xor U14361 (N_14361,N_13408,N_13255);
or U14362 (N_14362,N_13073,N_12994);
nand U14363 (N_14363,N_13450,N_13188);
nand U14364 (N_14364,N_12817,N_12319);
nor U14365 (N_14365,N_12477,N_12811);
xnor U14366 (N_14366,N_12934,N_13046);
nand U14367 (N_14367,N_12760,N_13154);
or U14368 (N_14368,N_13446,N_12315);
nand U14369 (N_14369,N_12189,N_12805);
xor U14370 (N_14370,N_12958,N_13075);
xor U14371 (N_14371,N_13402,N_12613);
nor U14372 (N_14372,N_13112,N_12267);
and U14373 (N_14373,N_13369,N_12133);
nor U14374 (N_14374,N_12467,N_13409);
nand U14375 (N_14375,N_13432,N_12844);
nand U14376 (N_14376,N_13471,N_12233);
nand U14377 (N_14377,N_13404,N_13015);
nor U14378 (N_14378,N_13164,N_12895);
nor U14379 (N_14379,N_13089,N_12823);
or U14380 (N_14380,N_12702,N_13026);
or U14381 (N_14381,N_13072,N_13416);
and U14382 (N_14382,N_12316,N_12939);
and U14383 (N_14383,N_12478,N_13490);
xnor U14384 (N_14384,N_12993,N_13449);
or U14385 (N_14385,N_12058,N_12202);
nand U14386 (N_14386,N_13114,N_12697);
or U14387 (N_14387,N_12174,N_12829);
xor U14388 (N_14388,N_12902,N_12951);
nand U14389 (N_14389,N_13298,N_13448);
nor U14390 (N_14390,N_12332,N_12265);
nor U14391 (N_14391,N_12958,N_12255);
xor U14392 (N_14392,N_13147,N_12024);
and U14393 (N_14393,N_12773,N_12017);
nand U14394 (N_14394,N_13221,N_12226);
nand U14395 (N_14395,N_12090,N_12218);
nor U14396 (N_14396,N_12273,N_12850);
nand U14397 (N_14397,N_13055,N_13432);
or U14398 (N_14398,N_13119,N_13180);
nor U14399 (N_14399,N_13488,N_12081);
xor U14400 (N_14400,N_12007,N_12133);
nand U14401 (N_14401,N_13377,N_12230);
and U14402 (N_14402,N_12743,N_13276);
nor U14403 (N_14403,N_12981,N_13461);
nand U14404 (N_14404,N_12401,N_13012);
nand U14405 (N_14405,N_13162,N_12114);
xnor U14406 (N_14406,N_13025,N_13416);
or U14407 (N_14407,N_12054,N_13138);
xnor U14408 (N_14408,N_12349,N_12400);
xnor U14409 (N_14409,N_12212,N_13029);
or U14410 (N_14410,N_12458,N_12862);
nor U14411 (N_14411,N_12823,N_12788);
xnor U14412 (N_14412,N_13071,N_13339);
or U14413 (N_14413,N_13076,N_13097);
xnor U14414 (N_14414,N_12433,N_13074);
and U14415 (N_14415,N_12132,N_12204);
and U14416 (N_14416,N_13439,N_13176);
or U14417 (N_14417,N_12666,N_13472);
nand U14418 (N_14418,N_12246,N_12573);
xnor U14419 (N_14419,N_12671,N_12898);
nand U14420 (N_14420,N_12806,N_12008);
or U14421 (N_14421,N_13207,N_13344);
and U14422 (N_14422,N_12214,N_12704);
nand U14423 (N_14423,N_12437,N_13150);
nand U14424 (N_14424,N_12710,N_13321);
xnor U14425 (N_14425,N_12266,N_13374);
or U14426 (N_14426,N_12825,N_13183);
nand U14427 (N_14427,N_12261,N_12595);
nand U14428 (N_14428,N_13030,N_13069);
nand U14429 (N_14429,N_13328,N_12117);
xor U14430 (N_14430,N_12172,N_13208);
xnor U14431 (N_14431,N_13397,N_13016);
nand U14432 (N_14432,N_12216,N_13360);
or U14433 (N_14433,N_12760,N_13126);
nor U14434 (N_14434,N_13456,N_12283);
nand U14435 (N_14435,N_12740,N_13068);
xnor U14436 (N_14436,N_13326,N_13101);
or U14437 (N_14437,N_12645,N_12459);
or U14438 (N_14438,N_13062,N_12636);
nand U14439 (N_14439,N_13046,N_13498);
or U14440 (N_14440,N_12020,N_12784);
nand U14441 (N_14441,N_12663,N_12426);
or U14442 (N_14442,N_13247,N_13101);
xnor U14443 (N_14443,N_13322,N_13188);
xor U14444 (N_14444,N_12678,N_13346);
xnor U14445 (N_14445,N_12084,N_12463);
xnor U14446 (N_14446,N_13348,N_12008);
nor U14447 (N_14447,N_12280,N_12594);
and U14448 (N_14448,N_12166,N_12010);
nor U14449 (N_14449,N_12083,N_13200);
nand U14450 (N_14450,N_12855,N_12485);
nand U14451 (N_14451,N_13353,N_12136);
xor U14452 (N_14452,N_12110,N_12739);
xnor U14453 (N_14453,N_12379,N_12863);
xor U14454 (N_14454,N_12503,N_13113);
nor U14455 (N_14455,N_12670,N_13099);
nand U14456 (N_14456,N_13484,N_13477);
and U14457 (N_14457,N_12356,N_12316);
xnor U14458 (N_14458,N_13354,N_13456);
xor U14459 (N_14459,N_12991,N_12515);
and U14460 (N_14460,N_12203,N_12584);
or U14461 (N_14461,N_12555,N_13402);
xor U14462 (N_14462,N_12422,N_12130);
and U14463 (N_14463,N_13290,N_12429);
and U14464 (N_14464,N_12661,N_12622);
nand U14465 (N_14465,N_12324,N_12649);
or U14466 (N_14466,N_13082,N_12737);
xor U14467 (N_14467,N_12603,N_12329);
and U14468 (N_14468,N_12770,N_12343);
nor U14469 (N_14469,N_12578,N_12123);
or U14470 (N_14470,N_12212,N_12319);
or U14471 (N_14471,N_12092,N_12073);
or U14472 (N_14472,N_12421,N_13334);
xnor U14473 (N_14473,N_12276,N_13080);
and U14474 (N_14474,N_12020,N_13045);
and U14475 (N_14475,N_13164,N_12315);
nor U14476 (N_14476,N_12905,N_13157);
xnor U14477 (N_14477,N_13056,N_13223);
nor U14478 (N_14478,N_13090,N_12400);
nor U14479 (N_14479,N_12954,N_13346);
xor U14480 (N_14480,N_12367,N_12190);
nor U14481 (N_14481,N_12925,N_12129);
nor U14482 (N_14482,N_13236,N_12245);
or U14483 (N_14483,N_12306,N_12920);
and U14484 (N_14484,N_13242,N_12254);
and U14485 (N_14485,N_12638,N_12864);
or U14486 (N_14486,N_12638,N_12778);
or U14487 (N_14487,N_12097,N_12248);
nor U14488 (N_14488,N_13107,N_13116);
xnor U14489 (N_14489,N_13144,N_12572);
xor U14490 (N_14490,N_13305,N_13459);
nand U14491 (N_14491,N_12689,N_12913);
nand U14492 (N_14492,N_13234,N_13416);
xnor U14493 (N_14493,N_13321,N_12582);
or U14494 (N_14494,N_12779,N_13130);
or U14495 (N_14495,N_12155,N_12591);
or U14496 (N_14496,N_12282,N_12179);
nand U14497 (N_14497,N_12583,N_12150);
or U14498 (N_14498,N_12129,N_12784);
xnor U14499 (N_14499,N_12390,N_12464);
nor U14500 (N_14500,N_12847,N_12200);
nor U14501 (N_14501,N_12740,N_12793);
and U14502 (N_14502,N_13410,N_13229);
xnor U14503 (N_14503,N_13384,N_13327);
nor U14504 (N_14504,N_12324,N_12860);
xnor U14505 (N_14505,N_12108,N_13206);
xor U14506 (N_14506,N_12033,N_12879);
nor U14507 (N_14507,N_12252,N_12011);
nor U14508 (N_14508,N_12021,N_12595);
xnor U14509 (N_14509,N_12054,N_12337);
xor U14510 (N_14510,N_13377,N_12546);
and U14511 (N_14511,N_13178,N_12715);
nor U14512 (N_14512,N_12857,N_12460);
and U14513 (N_14513,N_12731,N_12471);
nor U14514 (N_14514,N_13180,N_12051);
and U14515 (N_14515,N_13372,N_12512);
or U14516 (N_14516,N_12345,N_12647);
nor U14517 (N_14517,N_12608,N_12381);
xnor U14518 (N_14518,N_12354,N_13359);
xnor U14519 (N_14519,N_13091,N_13016);
nand U14520 (N_14520,N_13195,N_12139);
or U14521 (N_14521,N_13328,N_12456);
or U14522 (N_14522,N_13262,N_12261);
xnor U14523 (N_14523,N_12326,N_12388);
nor U14524 (N_14524,N_13128,N_13484);
and U14525 (N_14525,N_12246,N_12650);
nor U14526 (N_14526,N_13370,N_12575);
nor U14527 (N_14527,N_13377,N_12060);
nor U14528 (N_14528,N_13478,N_12686);
and U14529 (N_14529,N_12333,N_13320);
or U14530 (N_14530,N_12622,N_12497);
or U14531 (N_14531,N_12450,N_13447);
and U14532 (N_14532,N_12418,N_12937);
or U14533 (N_14533,N_13282,N_13484);
nor U14534 (N_14534,N_13072,N_12568);
nor U14535 (N_14535,N_13064,N_12799);
nor U14536 (N_14536,N_13144,N_13359);
xnor U14537 (N_14537,N_12245,N_12041);
or U14538 (N_14538,N_12157,N_13138);
nand U14539 (N_14539,N_12283,N_12801);
xnor U14540 (N_14540,N_12622,N_13361);
nor U14541 (N_14541,N_12359,N_13047);
or U14542 (N_14542,N_12202,N_13340);
nor U14543 (N_14543,N_13182,N_12953);
nor U14544 (N_14544,N_12443,N_12396);
nor U14545 (N_14545,N_12750,N_12456);
or U14546 (N_14546,N_13198,N_12912);
or U14547 (N_14547,N_12147,N_12609);
or U14548 (N_14548,N_12070,N_12610);
and U14549 (N_14549,N_12712,N_13228);
xor U14550 (N_14550,N_13210,N_13414);
or U14551 (N_14551,N_13378,N_12553);
nand U14552 (N_14552,N_12542,N_12189);
or U14553 (N_14553,N_13420,N_12485);
nor U14554 (N_14554,N_13484,N_12124);
and U14555 (N_14555,N_13128,N_12703);
xor U14556 (N_14556,N_12980,N_13288);
nor U14557 (N_14557,N_12558,N_12046);
and U14558 (N_14558,N_12347,N_13158);
nand U14559 (N_14559,N_12872,N_12830);
and U14560 (N_14560,N_12217,N_12411);
or U14561 (N_14561,N_12629,N_12158);
nor U14562 (N_14562,N_12692,N_12424);
nor U14563 (N_14563,N_12282,N_13364);
nor U14564 (N_14564,N_12607,N_13128);
nand U14565 (N_14565,N_12859,N_12981);
nand U14566 (N_14566,N_13052,N_12050);
xor U14567 (N_14567,N_12495,N_12375);
or U14568 (N_14568,N_13332,N_12971);
nor U14569 (N_14569,N_13251,N_13183);
nand U14570 (N_14570,N_12139,N_12173);
and U14571 (N_14571,N_12563,N_12136);
or U14572 (N_14572,N_12597,N_13047);
or U14573 (N_14573,N_12076,N_13375);
or U14574 (N_14574,N_12821,N_12527);
nor U14575 (N_14575,N_12282,N_12591);
nand U14576 (N_14576,N_13022,N_12143);
xnor U14577 (N_14577,N_12882,N_12467);
xor U14578 (N_14578,N_13443,N_13228);
nor U14579 (N_14579,N_13298,N_12362);
or U14580 (N_14580,N_12526,N_12297);
nor U14581 (N_14581,N_13433,N_13067);
xor U14582 (N_14582,N_12870,N_13180);
and U14583 (N_14583,N_13035,N_12356);
nand U14584 (N_14584,N_13458,N_12981);
or U14585 (N_14585,N_12031,N_13150);
or U14586 (N_14586,N_12870,N_13065);
and U14587 (N_14587,N_13477,N_12290);
and U14588 (N_14588,N_12006,N_12315);
or U14589 (N_14589,N_12867,N_12040);
or U14590 (N_14590,N_12308,N_13183);
nand U14591 (N_14591,N_12020,N_12495);
nand U14592 (N_14592,N_13136,N_13370);
xor U14593 (N_14593,N_12070,N_13330);
or U14594 (N_14594,N_12123,N_12174);
xor U14595 (N_14595,N_13412,N_12184);
nor U14596 (N_14596,N_13323,N_13371);
xnor U14597 (N_14597,N_12132,N_12393);
or U14598 (N_14598,N_12105,N_13353);
nor U14599 (N_14599,N_13039,N_12475);
xor U14600 (N_14600,N_12983,N_13475);
nand U14601 (N_14601,N_13211,N_13361);
nand U14602 (N_14602,N_13211,N_13039);
xnor U14603 (N_14603,N_12564,N_12645);
nor U14604 (N_14604,N_13010,N_12977);
nand U14605 (N_14605,N_12313,N_13320);
and U14606 (N_14606,N_13283,N_12405);
nand U14607 (N_14607,N_13191,N_13069);
nor U14608 (N_14608,N_12459,N_12637);
or U14609 (N_14609,N_12983,N_12689);
nand U14610 (N_14610,N_12243,N_12972);
and U14611 (N_14611,N_12808,N_12250);
xnor U14612 (N_14612,N_12065,N_12816);
nor U14613 (N_14613,N_13305,N_12479);
nor U14614 (N_14614,N_13326,N_12591);
xnor U14615 (N_14615,N_12838,N_12322);
nor U14616 (N_14616,N_13146,N_13313);
or U14617 (N_14617,N_12352,N_12152);
nand U14618 (N_14618,N_12334,N_12321);
or U14619 (N_14619,N_12606,N_12726);
or U14620 (N_14620,N_13050,N_12148);
and U14621 (N_14621,N_12306,N_12490);
nor U14622 (N_14622,N_12265,N_13496);
nand U14623 (N_14623,N_12016,N_13030);
nand U14624 (N_14624,N_13327,N_13228);
or U14625 (N_14625,N_13025,N_12248);
and U14626 (N_14626,N_13025,N_12290);
nor U14627 (N_14627,N_13226,N_12721);
nor U14628 (N_14628,N_12959,N_13461);
xnor U14629 (N_14629,N_12266,N_13081);
and U14630 (N_14630,N_12413,N_13121);
nor U14631 (N_14631,N_12599,N_12408);
or U14632 (N_14632,N_12500,N_13279);
or U14633 (N_14633,N_12693,N_12787);
xor U14634 (N_14634,N_12475,N_12313);
nand U14635 (N_14635,N_13313,N_12780);
xor U14636 (N_14636,N_12777,N_12773);
and U14637 (N_14637,N_13317,N_12110);
or U14638 (N_14638,N_12190,N_12434);
or U14639 (N_14639,N_12295,N_13313);
nand U14640 (N_14640,N_12438,N_12746);
or U14641 (N_14641,N_12567,N_12399);
nand U14642 (N_14642,N_12140,N_13244);
nor U14643 (N_14643,N_12531,N_12275);
and U14644 (N_14644,N_13051,N_12708);
and U14645 (N_14645,N_13417,N_12060);
xor U14646 (N_14646,N_12809,N_12878);
xor U14647 (N_14647,N_12252,N_12976);
or U14648 (N_14648,N_12541,N_12850);
or U14649 (N_14649,N_12018,N_12639);
or U14650 (N_14650,N_12790,N_12175);
xor U14651 (N_14651,N_12695,N_13223);
nor U14652 (N_14652,N_12335,N_13194);
or U14653 (N_14653,N_12685,N_13340);
nor U14654 (N_14654,N_12997,N_13337);
or U14655 (N_14655,N_12524,N_12985);
nor U14656 (N_14656,N_12791,N_12522);
xnor U14657 (N_14657,N_12572,N_13083);
nor U14658 (N_14658,N_12839,N_13491);
and U14659 (N_14659,N_13002,N_13271);
nor U14660 (N_14660,N_12347,N_12331);
or U14661 (N_14661,N_12749,N_12531);
nor U14662 (N_14662,N_13047,N_12183);
and U14663 (N_14663,N_12023,N_12624);
nor U14664 (N_14664,N_12809,N_12190);
or U14665 (N_14665,N_12556,N_13101);
xnor U14666 (N_14666,N_13351,N_12992);
or U14667 (N_14667,N_12452,N_12685);
nor U14668 (N_14668,N_12673,N_12067);
nand U14669 (N_14669,N_13457,N_13068);
or U14670 (N_14670,N_12384,N_12108);
nor U14671 (N_14671,N_12884,N_13210);
nand U14672 (N_14672,N_12337,N_13454);
and U14673 (N_14673,N_12742,N_13142);
nand U14674 (N_14674,N_12943,N_12295);
and U14675 (N_14675,N_12311,N_12230);
nand U14676 (N_14676,N_12133,N_12212);
or U14677 (N_14677,N_13137,N_12249);
and U14678 (N_14678,N_12170,N_12262);
nor U14679 (N_14679,N_12246,N_13031);
nand U14680 (N_14680,N_12888,N_13123);
or U14681 (N_14681,N_12727,N_12232);
nand U14682 (N_14682,N_12418,N_13134);
xor U14683 (N_14683,N_12751,N_12374);
nor U14684 (N_14684,N_12540,N_12236);
xor U14685 (N_14685,N_13242,N_12557);
and U14686 (N_14686,N_12363,N_13465);
xnor U14687 (N_14687,N_13161,N_12540);
nor U14688 (N_14688,N_12412,N_12228);
and U14689 (N_14689,N_13023,N_12220);
nor U14690 (N_14690,N_13345,N_12647);
nor U14691 (N_14691,N_12376,N_13295);
and U14692 (N_14692,N_13280,N_13236);
nand U14693 (N_14693,N_12358,N_12366);
nor U14694 (N_14694,N_12912,N_13444);
and U14695 (N_14695,N_13400,N_12487);
and U14696 (N_14696,N_12101,N_12718);
nand U14697 (N_14697,N_13372,N_12283);
nor U14698 (N_14698,N_13411,N_12950);
nand U14699 (N_14699,N_13018,N_12312);
and U14700 (N_14700,N_13215,N_13405);
or U14701 (N_14701,N_13260,N_12544);
xor U14702 (N_14702,N_13160,N_13382);
xnor U14703 (N_14703,N_13368,N_12179);
or U14704 (N_14704,N_13145,N_13189);
xnor U14705 (N_14705,N_12548,N_12279);
nand U14706 (N_14706,N_13385,N_12162);
xnor U14707 (N_14707,N_12276,N_13393);
nor U14708 (N_14708,N_12181,N_12630);
and U14709 (N_14709,N_12887,N_12794);
nor U14710 (N_14710,N_12929,N_12777);
xor U14711 (N_14711,N_13174,N_12185);
and U14712 (N_14712,N_12009,N_13039);
and U14713 (N_14713,N_12358,N_12844);
xnor U14714 (N_14714,N_12528,N_13003);
nor U14715 (N_14715,N_13224,N_12181);
or U14716 (N_14716,N_13373,N_12130);
nand U14717 (N_14717,N_12440,N_13258);
nand U14718 (N_14718,N_12564,N_12454);
nor U14719 (N_14719,N_12345,N_12949);
nor U14720 (N_14720,N_12368,N_13372);
nand U14721 (N_14721,N_12763,N_12327);
nor U14722 (N_14722,N_13117,N_12064);
nand U14723 (N_14723,N_13374,N_12077);
nor U14724 (N_14724,N_12811,N_13440);
nor U14725 (N_14725,N_12541,N_12240);
or U14726 (N_14726,N_12134,N_12060);
xnor U14727 (N_14727,N_12548,N_13460);
nand U14728 (N_14728,N_12712,N_12171);
and U14729 (N_14729,N_12318,N_12541);
or U14730 (N_14730,N_12982,N_13110);
or U14731 (N_14731,N_13347,N_12121);
or U14732 (N_14732,N_12309,N_12240);
nand U14733 (N_14733,N_13420,N_12413);
or U14734 (N_14734,N_12479,N_12319);
nor U14735 (N_14735,N_12392,N_12084);
nor U14736 (N_14736,N_12795,N_12477);
nand U14737 (N_14737,N_12935,N_12268);
nor U14738 (N_14738,N_12518,N_12638);
and U14739 (N_14739,N_13201,N_12793);
nand U14740 (N_14740,N_12746,N_13128);
nor U14741 (N_14741,N_12102,N_13299);
or U14742 (N_14742,N_13313,N_12806);
xnor U14743 (N_14743,N_12237,N_12692);
nor U14744 (N_14744,N_13248,N_13459);
nand U14745 (N_14745,N_13427,N_12967);
nor U14746 (N_14746,N_13315,N_12134);
nand U14747 (N_14747,N_13398,N_13203);
nor U14748 (N_14748,N_12571,N_12834);
xnor U14749 (N_14749,N_12352,N_12178);
xnor U14750 (N_14750,N_13251,N_13482);
nor U14751 (N_14751,N_13020,N_13060);
xor U14752 (N_14752,N_12446,N_13398);
or U14753 (N_14753,N_12248,N_13254);
and U14754 (N_14754,N_12048,N_13112);
or U14755 (N_14755,N_12072,N_12042);
xnor U14756 (N_14756,N_13176,N_12480);
or U14757 (N_14757,N_12656,N_12234);
xor U14758 (N_14758,N_13267,N_12410);
and U14759 (N_14759,N_12693,N_13390);
nand U14760 (N_14760,N_12663,N_13282);
nor U14761 (N_14761,N_13000,N_13464);
and U14762 (N_14762,N_12715,N_12784);
or U14763 (N_14763,N_13451,N_13171);
nor U14764 (N_14764,N_12328,N_12797);
or U14765 (N_14765,N_12261,N_12460);
nand U14766 (N_14766,N_13101,N_12663);
and U14767 (N_14767,N_12946,N_12175);
nor U14768 (N_14768,N_13199,N_12371);
xnor U14769 (N_14769,N_12960,N_13394);
xnor U14770 (N_14770,N_12546,N_12340);
xor U14771 (N_14771,N_12095,N_13497);
or U14772 (N_14772,N_13105,N_13420);
nand U14773 (N_14773,N_13065,N_12616);
and U14774 (N_14774,N_12573,N_12994);
nand U14775 (N_14775,N_12340,N_12106);
or U14776 (N_14776,N_13265,N_12233);
nand U14777 (N_14777,N_12674,N_12790);
nor U14778 (N_14778,N_13065,N_13383);
or U14779 (N_14779,N_12706,N_12900);
nand U14780 (N_14780,N_12393,N_12516);
or U14781 (N_14781,N_13357,N_12776);
nand U14782 (N_14782,N_12992,N_13096);
or U14783 (N_14783,N_12259,N_13164);
and U14784 (N_14784,N_12043,N_12362);
nand U14785 (N_14785,N_12463,N_12012);
nand U14786 (N_14786,N_13196,N_13043);
nand U14787 (N_14787,N_12467,N_12785);
or U14788 (N_14788,N_13284,N_13330);
and U14789 (N_14789,N_13396,N_12336);
nor U14790 (N_14790,N_12519,N_12725);
nor U14791 (N_14791,N_13296,N_13098);
or U14792 (N_14792,N_12858,N_12884);
or U14793 (N_14793,N_12537,N_13341);
xnor U14794 (N_14794,N_12955,N_13328);
and U14795 (N_14795,N_13495,N_12862);
and U14796 (N_14796,N_12770,N_13449);
or U14797 (N_14797,N_13201,N_13376);
xnor U14798 (N_14798,N_12759,N_12577);
nor U14799 (N_14799,N_13493,N_12040);
nor U14800 (N_14800,N_12895,N_12045);
and U14801 (N_14801,N_12864,N_13440);
nand U14802 (N_14802,N_12578,N_13225);
nand U14803 (N_14803,N_12665,N_13078);
nand U14804 (N_14804,N_13397,N_12443);
or U14805 (N_14805,N_12229,N_13342);
xor U14806 (N_14806,N_13241,N_12457);
nand U14807 (N_14807,N_12352,N_12212);
xor U14808 (N_14808,N_13340,N_12297);
nor U14809 (N_14809,N_12805,N_12696);
xnor U14810 (N_14810,N_12198,N_12767);
or U14811 (N_14811,N_12793,N_12472);
nand U14812 (N_14812,N_12280,N_12433);
or U14813 (N_14813,N_12077,N_13255);
and U14814 (N_14814,N_12868,N_12653);
xnor U14815 (N_14815,N_12945,N_12386);
or U14816 (N_14816,N_12545,N_12195);
and U14817 (N_14817,N_13438,N_13292);
or U14818 (N_14818,N_12280,N_12834);
nor U14819 (N_14819,N_13160,N_12985);
or U14820 (N_14820,N_13427,N_12762);
nor U14821 (N_14821,N_13086,N_12931);
nor U14822 (N_14822,N_12411,N_12402);
xor U14823 (N_14823,N_12503,N_12504);
and U14824 (N_14824,N_12178,N_13374);
nand U14825 (N_14825,N_12209,N_12331);
and U14826 (N_14826,N_12201,N_12641);
nor U14827 (N_14827,N_12884,N_12639);
and U14828 (N_14828,N_12501,N_12136);
nor U14829 (N_14829,N_12614,N_12729);
nand U14830 (N_14830,N_12130,N_13329);
and U14831 (N_14831,N_13297,N_13285);
nor U14832 (N_14832,N_12962,N_12565);
xor U14833 (N_14833,N_13431,N_13277);
or U14834 (N_14834,N_13316,N_12398);
xor U14835 (N_14835,N_12417,N_13227);
or U14836 (N_14836,N_12352,N_12683);
nor U14837 (N_14837,N_12726,N_13356);
nor U14838 (N_14838,N_12426,N_13248);
nor U14839 (N_14839,N_12219,N_12131);
and U14840 (N_14840,N_12963,N_12740);
nand U14841 (N_14841,N_12994,N_13122);
nand U14842 (N_14842,N_13235,N_13471);
xnor U14843 (N_14843,N_12410,N_13335);
and U14844 (N_14844,N_12113,N_13093);
or U14845 (N_14845,N_12564,N_12396);
nand U14846 (N_14846,N_13005,N_12716);
nor U14847 (N_14847,N_12080,N_12746);
nand U14848 (N_14848,N_12032,N_13219);
and U14849 (N_14849,N_13184,N_13223);
nor U14850 (N_14850,N_12512,N_12264);
nor U14851 (N_14851,N_13215,N_12617);
and U14852 (N_14852,N_12556,N_13031);
xor U14853 (N_14853,N_12125,N_13386);
nor U14854 (N_14854,N_12592,N_12269);
and U14855 (N_14855,N_13219,N_13117);
or U14856 (N_14856,N_12974,N_12496);
xor U14857 (N_14857,N_12904,N_12956);
nand U14858 (N_14858,N_12205,N_13422);
and U14859 (N_14859,N_13059,N_12528);
nand U14860 (N_14860,N_13174,N_12920);
xnor U14861 (N_14861,N_13072,N_13092);
nand U14862 (N_14862,N_12975,N_12038);
or U14863 (N_14863,N_13116,N_12585);
nor U14864 (N_14864,N_13416,N_13170);
xnor U14865 (N_14865,N_12588,N_12128);
or U14866 (N_14866,N_13239,N_12456);
and U14867 (N_14867,N_12453,N_12183);
or U14868 (N_14868,N_12783,N_13436);
nand U14869 (N_14869,N_12962,N_13232);
xnor U14870 (N_14870,N_12825,N_13464);
or U14871 (N_14871,N_13371,N_12067);
xnor U14872 (N_14872,N_12792,N_12652);
nor U14873 (N_14873,N_12952,N_12775);
and U14874 (N_14874,N_12666,N_13219);
nand U14875 (N_14875,N_12981,N_12378);
nand U14876 (N_14876,N_13239,N_12910);
xor U14877 (N_14877,N_13212,N_12771);
xor U14878 (N_14878,N_12322,N_12564);
nand U14879 (N_14879,N_12647,N_12407);
xnor U14880 (N_14880,N_12137,N_13012);
xor U14881 (N_14881,N_12801,N_13005);
or U14882 (N_14882,N_13285,N_12823);
nand U14883 (N_14883,N_12098,N_12147);
nor U14884 (N_14884,N_12910,N_12034);
or U14885 (N_14885,N_13048,N_12865);
and U14886 (N_14886,N_12200,N_12218);
or U14887 (N_14887,N_13007,N_13124);
xor U14888 (N_14888,N_12130,N_12872);
and U14889 (N_14889,N_12366,N_12460);
and U14890 (N_14890,N_13209,N_12075);
nand U14891 (N_14891,N_12389,N_13083);
xnor U14892 (N_14892,N_12156,N_12227);
nand U14893 (N_14893,N_12447,N_12672);
or U14894 (N_14894,N_13473,N_13047);
xor U14895 (N_14895,N_13425,N_13452);
and U14896 (N_14896,N_12528,N_12379);
xor U14897 (N_14897,N_12350,N_12948);
or U14898 (N_14898,N_12088,N_13179);
xor U14899 (N_14899,N_12314,N_12306);
and U14900 (N_14900,N_12889,N_13343);
or U14901 (N_14901,N_12950,N_12307);
nor U14902 (N_14902,N_13479,N_12243);
and U14903 (N_14903,N_12281,N_13262);
and U14904 (N_14904,N_12545,N_13326);
nor U14905 (N_14905,N_12046,N_13434);
nand U14906 (N_14906,N_13454,N_12755);
and U14907 (N_14907,N_13184,N_12517);
and U14908 (N_14908,N_12366,N_13080);
or U14909 (N_14909,N_12944,N_12561);
nand U14910 (N_14910,N_12165,N_12460);
nor U14911 (N_14911,N_12975,N_13406);
or U14912 (N_14912,N_12197,N_12992);
and U14913 (N_14913,N_12791,N_12776);
xor U14914 (N_14914,N_13321,N_13224);
xnor U14915 (N_14915,N_12962,N_12620);
nand U14916 (N_14916,N_12965,N_12096);
or U14917 (N_14917,N_12923,N_12859);
or U14918 (N_14918,N_12692,N_12119);
nor U14919 (N_14919,N_12329,N_13097);
xor U14920 (N_14920,N_13326,N_13182);
and U14921 (N_14921,N_13358,N_12084);
xor U14922 (N_14922,N_12779,N_12880);
nor U14923 (N_14923,N_12443,N_13403);
xor U14924 (N_14924,N_12204,N_12526);
or U14925 (N_14925,N_13432,N_13254);
nand U14926 (N_14926,N_12187,N_12393);
xnor U14927 (N_14927,N_12925,N_13315);
nor U14928 (N_14928,N_12657,N_12324);
nand U14929 (N_14929,N_12383,N_12001);
xnor U14930 (N_14930,N_12867,N_12381);
xnor U14931 (N_14931,N_12426,N_12270);
nand U14932 (N_14932,N_12930,N_12589);
or U14933 (N_14933,N_12547,N_13203);
xnor U14934 (N_14934,N_13392,N_12870);
nor U14935 (N_14935,N_12941,N_12603);
and U14936 (N_14936,N_12443,N_12814);
xor U14937 (N_14937,N_12723,N_12490);
nor U14938 (N_14938,N_13242,N_12051);
or U14939 (N_14939,N_12493,N_12540);
xnor U14940 (N_14940,N_12497,N_12252);
nor U14941 (N_14941,N_13388,N_12902);
nor U14942 (N_14942,N_12512,N_12035);
nand U14943 (N_14943,N_12934,N_12701);
and U14944 (N_14944,N_12607,N_12364);
or U14945 (N_14945,N_13424,N_12042);
or U14946 (N_14946,N_12258,N_12352);
and U14947 (N_14947,N_12743,N_13249);
nor U14948 (N_14948,N_13268,N_13149);
or U14949 (N_14949,N_13470,N_13186);
xor U14950 (N_14950,N_12722,N_12789);
nand U14951 (N_14951,N_12184,N_13208);
xor U14952 (N_14952,N_12626,N_12367);
nor U14953 (N_14953,N_12188,N_13446);
or U14954 (N_14954,N_13297,N_12718);
nand U14955 (N_14955,N_12809,N_12236);
nand U14956 (N_14956,N_12857,N_12880);
xor U14957 (N_14957,N_13359,N_12719);
xnor U14958 (N_14958,N_13396,N_13330);
nor U14959 (N_14959,N_12751,N_12197);
nor U14960 (N_14960,N_13062,N_12363);
xnor U14961 (N_14961,N_12087,N_12841);
nand U14962 (N_14962,N_12226,N_12430);
nand U14963 (N_14963,N_12316,N_12263);
nand U14964 (N_14964,N_12302,N_12161);
xnor U14965 (N_14965,N_12528,N_12709);
nor U14966 (N_14966,N_12098,N_12533);
nand U14967 (N_14967,N_13146,N_12421);
or U14968 (N_14968,N_12092,N_12742);
xor U14969 (N_14969,N_12034,N_12825);
and U14970 (N_14970,N_12372,N_13487);
and U14971 (N_14971,N_13475,N_13465);
nor U14972 (N_14972,N_13080,N_13401);
xnor U14973 (N_14973,N_12449,N_13193);
or U14974 (N_14974,N_13086,N_13076);
xnor U14975 (N_14975,N_12802,N_12585);
or U14976 (N_14976,N_12395,N_12655);
and U14977 (N_14977,N_13084,N_12050);
nor U14978 (N_14978,N_12993,N_13365);
xnor U14979 (N_14979,N_12429,N_13374);
xnor U14980 (N_14980,N_12305,N_13460);
or U14981 (N_14981,N_13404,N_12824);
and U14982 (N_14982,N_12250,N_12949);
and U14983 (N_14983,N_13081,N_12415);
nor U14984 (N_14984,N_12122,N_13048);
nor U14985 (N_14985,N_12818,N_12365);
nor U14986 (N_14986,N_12072,N_12844);
nor U14987 (N_14987,N_13231,N_12984);
or U14988 (N_14988,N_12457,N_13299);
nor U14989 (N_14989,N_12349,N_13026);
xnor U14990 (N_14990,N_12817,N_12006);
xor U14991 (N_14991,N_13176,N_12939);
or U14992 (N_14992,N_12334,N_12596);
nand U14993 (N_14993,N_12514,N_13470);
nor U14994 (N_14994,N_13021,N_12593);
xor U14995 (N_14995,N_13035,N_13124);
nand U14996 (N_14996,N_13325,N_12277);
nand U14997 (N_14997,N_13254,N_12471);
nor U14998 (N_14998,N_12645,N_13367);
nor U14999 (N_14999,N_13438,N_13249);
or U15000 (N_15000,N_14961,N_14851);
or U15001 (N_15001,N_13778,N_13535);
and U15002 (N_15002,N_14788,N_13624);
nor U15003 (N_15003,N_14958,N_13825);
and U15004 (N_15004,N_14755,N_14538);
or U15005 (N_15005,N_13544,N_14478);
and U15006 (N_15006,N_14456,N_13616);
and U15007 (N_15007,N_13645,N_13814);
or U15008 (N_15008,N_13972,N_14643);
nor U15009 (N_15009,N_14654,N_14989);
or U15010 (N_15010,N_14737,N_14226);
and U15011 (N_15011,N_14777,N_14563);
and U15012 (N_15012,N_14753,N_14114);
or U15013 (N_15013,N_14844,N_14276);
nand U15014 (N_15014,N_14768,N_14317);
xor U15015 (N_15015,N_14490,N_14818);
and U15016 (N_15016,N_14158,N_14612);
nand U15017 (N_15017,N_13986,N_13626);
nand U15018 (N_15018,N_14159,N_14202);
and U15019 (N_15019,N_14821,N_14319);
nor U15020 (N_15020,N_14133,N_13765);
nand U15021 (N_15021,N_14089,N_13822);
xor U15022 (N_15022,N_13963,N_14693);
nand U15023 (N_15023,N_13861,N_14959);
and U15024 (N_15024,N_13957,N_14942);
or U15025 (N_15025,N_14687,N_14901);
nand U15026 (N_15026,N_14894,N_14064);
nor U15027 (N_15027,N_14746,N_14832);
and U15028 (N_15028,N_13750,N_13643);
and U15029 (N_15029,N_14625,N_14730);
and U15030 (N_15030,N_13581,N_14173);
xor U15031 (N_15031,N_14546,N_14891);
or U15032 (N_15032,N_13826,N_13864);
nand U15033 (N_15033,N_14212,N_14077);
nor U15034 (N_15034,N_14984,N_13731);
xnor U15035 (N_15035,N_14008,N_13553);
nor U15036 (N_15036,N_14009,N_13910);
nor U15037 (N_15037,N_14751,N_13658);
and U15038 (N_15038,N_14448,N_13742);
nor U15039 (N_15039,N_14076,N_14154);
xor U15040 (N_15040,N_13894,N_14710);
nand U15041 (N_15041,N_13510,N_13813);
xnor U15042 (N_15042,N_14794,N_14667);
or U15043 (N_15043,N_14474,N_13599);
nor U15044 (N_15044,N_14447,N_13797);
and U15045 (N_15045,N_14201,N_14579);
xnor U15046 (N_15046,N_13831,N_13613);
nor U15047 (N_15047,N_14278,N_14800);
nand U15048 (N_15048,N_14219,N_14450);
and U15049 (N_15049,N_13646,N_14605);
nand U15050 (N_15050,N_13841,N_14039);
or U15051 (N_15051,N_13941,N_14198);
and U15052 (N_15052,N_14248,N_14912);
nand U15053 (N_15053,N_13533,N_13566);
nor U15054 (N_15054,N_14675,N_14137);
or U15055 (N_15055,N_13737,N_13523);
nor U15056 (N_15056,N_13876,N_14745);
nor U15057 (N_15057,N_14981,N_13890);
nand U15058 (N_15058,N_14398,N_14740);
and U15059 (N_15059,N_14081,N_13976);
or U15060 (N_15060,N_14203,N_14664);
xnor U15061 (N_15061,N_14444,N_14520);
nor U15062 (N_15062,N_14145,N_14528);
and U15063 (N_15063,N_14000,N_14140);
or U15064 (N_15064,N_14797,N_13611);
xor U15065 (N_15065,N_14555,N_14488);
nand U15066 (N_15066,N_13966,N_13816);
nand U15067 (N_15067,N_14998,N_14714);
or U15068 (N_15068,N_14518,N_14229);
and U15069 (N_15069,N_13653,N_13933);
nor U15070 (N_15070,N_14939,N_13904);
or U15071 (N_15071,N_13588,N_14500);
nand U15072 (N_15072,N_14952,N_13925);
xnor U15073 (N_15073,N_13579,N_14300);
or U15074 (N_15074,N_13732,N_14964);
xnor U15075 (N_15075,N_13843,N_14469);
xor U15076 (N_15076,N_14780,N_14749);
nand U15077 (N_15077,N_14434,N_14729);
xnor U15078 (N_15078,N_14014,N_14791);
nand U15079 (N_15079,N_14242,N_14858);
nand U15080 (N_15080,N_14193,N_13884);
xnor U15081 (N_15081,N_14040,N_14532);
nand U15082 (N_15082,N_14921,N_13929);
nor U15083 (N_15083,N_14302,N_14165);
nor U15084 (N_15084,N_13665,N_14757);
or U15085 (N_15085,N_14233,N_14351);
nor U15086 (N_15086,N_13952,N_13869);
or U15087 (N_15087,N_13980,N_14825);
and U15088 (N_15088,N_13744,N_13725);
nand U15089 (N_15089,N_14385,N_13766);
xor U15090 (N_15090,N_13949,N_14568);
nor U15091 (N_15091,N_14280,N_14170);
nor U15092 (N_15092,N_14421,N_14019);
and U15093 (N_15093,N_13714,N_13767);
nand U15094 (N_15094,N_14350,N_14222);
nor U15095 (N_15095,N_14069,N_14781);
nand U15096 (N_15096,N_14310,N_14423);
nor U15097 (N_15097,N_14815,N_13908);
nor U15098 (N_15098,N_14037,N_14656);
and U15099 (N_15099,N_14366,N_14752);
nand U15100 (N_15100,N_14570,N_14495);
nand U15101 (N_15101,N_14882,N_14100);
nor U15102 (N_15102,N_14264,N_14836);
nor U15103 (N_15103,N_14129,N_13607);
xor U15104 (N_15104,N_14718,N_14250);
or U15105 (N_15105,N_14839,N_14491);
nor U15106 (N_15106,N_14147,N_14621);
or U15107 (N_15107,N_14185,N_13691);
nor U15108 (N_15108,N_14281,N_14228);
and U15109 (N_15109,N_14188,N_14172);
xnor U15110 (N_15110,N_13503,N_14983);
nor U15111 (N_15111,N_14282,N_13569);
and U15112 (N_15112,N_13871,N_14134);
and U15113 (N_15113,N_14936,N_14196);
and U15114 (N_15114,N_14880,N_14686);
nand U15115 (N_15115,N_14445,N_14760);
and U15116 (N_15116,N_14871,N_13635);
and U15117 (N_15117,N_14006,N_13850);
nand U15118 (N_15118,N_14689,N_14820);
or U15119 (N_15119,N_14420,N_14412);
or U15120 (N_15120,N_13517,N_13558);
nand U15121 (N_15121,N_13804,N_14599);
xnor U15122 (N_15122,N_13991,N_14017);
nor U15123 (N_15123,N_13664,N_13760);
xnor U15124 (N_15124,N_14397,N_13522);
xor U15125 (N_15125,N_14462,N_13719);
xor U15126 (N_15126,N_14132,N_14722);
and U15127 (N_15127,N_13542,N_13838);
or U15128 (N_15128,N_13748,N_14523);
and U15129 (N_15129,N_14809,N_14956);
xor U15130 (N_15130,N_14988,N_13885);
or U15131 (N_15131,N_13504,N_14018);
nor U15132 (N_15132,N_14613,N_13552);
xor U15133 (N_15133,N_14769,N_14841);
or U15134 (N_15134,N_13902,N_14860);
and U15135 (N_15135,N_14123,N_13857);
nor U15136 (N_15136,N_14330,N_14050);
nor U15137 (N_15137,N_13514,N_14189);
and U15138 (N_15138,N_14504,N_14774);
or U15139 (N_15139,N_13708,N_13697);
and U15140 (N_15140,N_14245,N_14096);
nand U15141 (N_15141,N_14109,N_14094);
or U15142 (N_15142,N_14519,N_13911);
xor U15143 (N_15143,N_14510,N_14341);
or U15144 (N_15144,N_13571,N_14576);
or U15145 (N_15145,N_13649,N_14829);
xnor U15146 (N_15146,N_14063,N_14771);
or U15147 (N_15147,N_14015,N_14879);
nor U15148 (N_15148,N_14057,N_14526);
and U15149 (N_15149,N_13852,N_14151);
nand U15150 (N_15150,N_14442,N_14699);
xnor U15151 (N_15151,N_14890,N_13516);
nand U15152 (N_15152,N_14881,N_13680);
or U15153 (N_15153,N_14803,N_13543);
and U15154 (N_15154,N_13881,N_14443);
xor U15155 (N_15155,N_14941,N_14349);
nor U15156 (N_15156,N_14830,N_14802);
and U15157 (N_15157,N_14783,N_13576);
and U15158 (N_15158,N_14848,N_14003);
and U15159 (N_15159,N_14974,N_14235);
and U15160 (N_15160,N_13678,N_13805);
xnor U15161 (N_15161,N_14982,N_13992);
xor U15162 (N_15162,N_14726,N_13661);
or U15163 (N_15163,N_14082,N_13866);
nor U15164 (N_15164,N_14852,N_14262);
xor U15165 (N_15165,N_14937,N_13932);
and U15166 (N_15166,N_14150,N_13935);
nor U15167 (N_15167,N_13791,N_14176);
or U15168 (N_15168,N_13905,N_14918);
and U15169 (N_15169,N_14139,N_14241);
xnor U15170 (N_15170,N_13840,N_14609);
or U15171 (N_15171,N_14266,N_13741);
or U15172 (N_15172,N_13809,N_13886);
or U15173 (N_15173,N_14394,N_14466);
nand U15174 (N_15174,N_14208,N_14552);
xnor U15175 (N_15175,N_14935,N_14685);
xor U15176 (N_15176,N_13829,N_14766);
or U15177 (N_15177,N_14190,N_14376);
or U15178 (N_15178,N_14624,N_14298);
or U15179 (N_15179,N_13660,N_14712);
nor U15180 (N_15180,N_14425,N_13659);
nor U15181 (N_15181,N_14197,N_13743);
nand U15182 (N_15182,N_13855,N_14223);
and U15183 (N_15183,N_14590,N_13759);
and U15184 (N_15184,N_14738,N_14889);
xnor U15185 (N_15185,N_14143,N_13632);
and U15186 (N_15186,N_13548,N_14359);
and U15187 (N_15187,N_14976,N_14294);
or U15188 (N_15188,N_14915,N_14410);
nor U15189 (N_15189,N_13511,N_13573);
nor U15190 (N_15190,N_14217,N_13701);
xor U15191 (N_15191,N_13944,N_14325);
nand U15192 (N_15192,N_13700,N_14141);
and U15193 (N_15193,N_14405,N_14582);
or U15194 (N_15194,N_14790,N_13860);
xor U15195 (N_15195,N_14108,N_14782);
and U15196 (N_15196,N_14627,N_14786);
xnor U15197 (N_15197,N_13921,N_13705);
xnor U15198 (N_15198,N_14616,N_14011);
or U15199 (N_15199,N_14615,N_14822);
or U15200 (N_15200,N_13845,N_14418);
and U15201 (N_15201,N_14259,N_14292);
and U15202 (N_15202,N_14183,N_13836);
nor U15203 (N_15203,N_14042,N_14536);
or U15204 (N_15204,N_13679,N_14909);
and U15205 (N_15205,N_13739,N_14458);
xor U15206 (N_15206,N_13594,N_13720);
nand U15207 (N_15207,N_13648,N_14284);
nor U15208 (N_15208,N_14043,N_13936);
and U15209 (N_15209,N_14091,N_14269);
or U15210 (N_15210,N_14943,N_14494);
and U15211 (N_15211,N_14007,N_14638);
nand U15212 (N_15212,N_14911,N_14662);
and U15213 (N_15213,N_14713,N_14323);
nand U15214 (N_15214,N_13979,N_14097);
and U15215 (N_15215,N_14084,N_13612);
nand U15216 (N_15216,N_13781,N_14672);
and U15217 (N_15217,N_13554,N_13630);
or U15218 (N_15218,N_13993,N_14121);
and U15219 (N_15219,N_14066,N_14246);
xnor U15220 (N_15220,N_13668,N_14876);
nor U15221 (N_15221,N_14275,N_14467);
xor U15222 (N_15222,N_14953,N_14971);
and U15223 (N_15223,N_13536,N_14103);
nand U15224 (N_15224,N_13997,N_14034);
xnor U15225 (N_15225,N_14216,N_13519);
nor U15226 (N_15226,N_13983,N_14090);
xor U15227 (N_15227,N_14177,N_14869);
and U15228 (N_15228,N_14168,N_13790);
xnor U15229 (N_15229,N_14754,N_13785);
xor U15230 (N_15230,N_13682,N_14669);
or U15231 (N_15231,N_14016,N_14704);
nor U15232 (N_15232,N_14804,N_14473);
xnor U15233 (N_15233,N_13574,N_13789);
or U15234 (N_15234,N_13617,N_14736);
and U15235 (N_15235,N_14631,N_14358);
or U15236 (N_15236,N_13818,N_13923);
and U15237 (N_15237,N_13846,N_14299);
nand U15238 (N_15238,N_14905,N_13810);
xnor U15239 (N_15239,N_14853,N_14301);
or U15240 (N_15240,N_14079,N_13647);
nor U15241 (N_15241,N_13851,N_13507);
and U15242 (N_15242,N_13798,N_13508);
and U15243 (N_15243,N_14171,N_14061);
nor U15244 (N_15244,N_13513,N_14785);
nand U15245 (N_15245,N_14484,N_13951);
nor U15246 (N_15246,N_14928,N_14332);
or U15247 (N_15247,N_14169,N_14221);
nand U15248 (N_15248,N_13762,N_14338);
and U15249 (N_15249,N_13783,N_13589);
and U15250 (N_15250,N_14994,N_14556);
nor U15251 (N_15251,N_14424,N_14592);
nand U15252 (N_15252,N_14184,N_14966);
nor U15253 (N_15253,N_13967,N_14649);
nor U15254 (N_15254,N_14030,N_14949);
nand U15255 (N_15255,N_14130,N_13770);
and U15256 (N_15256,N_14864,N_14052);
xnor U15257 (N_15257,N_14254,N_13733);
nor U15258 (N_15258,N_13893,N_14348);
xor U15259 (N_15259,N_14382,N_14431);
nand U15260 (N_15260,N_13953,N_14578);
nor U15261 (N_15261,N_13696,N_14684);
xor U15262 (N_15262,N_13801,N_14544);
nor U15263 (N_15263,N_13891,N_13955);
nand U15264 (N_15264,N_13912,N_13954);
xnor U15265 (N_15265,N_14204,N_13915);
xor U15266 (N_15266,N_14062,N_13629);
and U15267 (N_15267,N_14303,N_13771);
or U15268 (N_15268,N_13694,N_13506);
or U15269 (N_15269,N_14875,N_14806);
nor U15270 (N_15270,N_14220,N_13878);
or U15271 (N_15271,N_14933,N_13833);
nand U15272 (N_15272,N_14762,N_14773);
nand U15273 (N_15273,N_14210,N_13977);
and U15274 (N_15274,N_13916,N_14162);
nor U15275 (N_15275,N_14496,N_14639);
nand U15276 (N_15276,N_13721,N_13591);
xnor U15277 (N_15277,N_14872,N_13650);
or U15278 (N_15278,N_14438,N_13776);
nand U15279 (N_15279,N_13882,N_13956);
or U15280 (N_15280,N_14427,N_14742);
or U15281 (N_15281,N_13920,N_14175);
xnor U15282 (N_15282,N_13639,N_14419);
nor U15283 (N_15283,N_14618,N_14868);
and U15284 (N_15284,N_14502,N_14148);
xor U15285 (N_15285,N_13978,N_14711);
nor U15286 (N_15286,N_14642,N_14522);
nand U15287 (N_15287,N_14483,N_14807);
or U15288 (N_15288,N_13560,N_14920);
nand U15289 (N_15289,N_13500,N_13572);
nand U15290 (N_15290,N_14411,N_13567);
nor U15291 (N_15291,N_14572,N_14731);
and U15292 (N_15292,N_14499,N_13652);
and U15293 (N_15293,N_14027,N_14842);
xor U15294 (N_15294,N_13928,N_14230);
or U15295 (N_15295,N_14614,N_13549);
or U15296 (N_15296,N_13625,N_13965);
nand U15297 (N_15297,N_14291,N_14827);
and U15298 (N_15298,N_14194,N_14873);
nand U15299 (N_15299,N_14346,N_14679);
nand U15300 (N_15300,N_14602,N_14065);
xor U15301 (N_15301,N_14367,N_13667);
nor U15302 (N_15302,N_13837,N_13848);
and U15303 (N_15303,N_14131,N_13620);
or U15304 (N_15304,N_14948,N_13559);
nand U15305 (N_15305,N_13969,N_14163);
nand U15306 (N_15306,N_13621,N_13862);
nand U15307 (N_15307,N_14646,N_14272);
and U15308 (N_15308,N_14663,N_14595);
nor U15309 (N_15309,N_14898,N_14877);
or U15310 (N_15310,N_14214,N_14593);
and U15311 (N_15311,N_14166,N_14485);
xnor U15312 (N_15312,N_13695,N_13931);
nor U15313 (N_15313,N_14102,N_13662);
nand U15314 (N_15314,N_13815,N_13873);
nor U15315 (N_15315,N_14354,N_13634);
nand U15316 (N_15316,N_14178,N_14309);
and U15317 (N_15317,N_13780,N_14051);
or U15318 (N_15318,N_14551,N_14534);
or U15319 (N_15319,N_13675,N_14925);
nand U15320 (N_15320,N_14290,N_14761);
nor U15321 (N_15321,N_14459,N_13819);
and U15322 (N_15322,N_14049,N_14985);
and U15323 (N_15323,N_13689,N_13686);
nor U15324 (N_15324,N_14471,N_14296);
or U15325 (N_15325,N_14914,N_14277);
nor U15326 (N_15326,N_13927,N_13619);
or U15327 (N_15327,N_14353,N_14694);
and U15328 (N_15328,N_14583,N_14573);
and U15329 (N_15329,N_13938,N_13764);
nand U15330 (N_15330,N_14048,N_14863);
or U15331 (N_15331,N_14564,N_13711);
nor U15332 (N_15332,N_14371,N_14831);
nand U15333 (N_15333,N_14088,N_14240);
nor U15334 (N_15334,N_14322,N_13609);
and U15335 (N_15335,N_14126,N_14940);
nor U15336 (N_15336,N_14112,N_13688);
and U15337 (N_15337,N_13671,N_13918);
xor U15338 (N_15338,N_13757,N_13999);
nand U15339 (N_15339,N_13706,N_14814);
or U15340 (N_15340,N_14792,N_14308);
xor U15341 (N_15341,N_13570,N_14938);
xor U15342 (N_15342,N_14020,N_14026);
nor U15343 (N_15343,N_14630,N_14452);
nor U15344 (N_15344,N_14924,N_14969);
nor U15345 (N_15345,N_14509,N_13557);
nand U15346 (N_15346,N_14598,N_14339);
nor U15347 (N_15347,N_13631,N_13520);
nand U15348 (N_15348,N_14747,N_14545);
nand U15349 (N_15349,N_13524,N_14327);
nand U15350 (N_15350,N_13755,N_14263);
xor U15351 (N_15351,N_14856,N_14334);
nand U15352 (N_15352,N_14934,N_14732);
xor U15353 (N_15353,N_13793,N_14960);
or U15354 (N_15354,N_14068,N_14659);
or U15355 (N_15355,N_14257,N_14415);
or U15356 (N_15356,N_14239,N_14489);
or U15357 (N_15357,N_13924,N_14874);
xnor U15358 (N_15358,N_14796,N_14629);
xnor U15359 (N_15359,N_13820,N_14023);
xor U15360 (N_15360,N_14373,N_13640);
nand U15361 (N_15361,N_14429,N_14288);
nor U15362 (N_15362,N_14946,N_13800);
or U15363 (N_15363,N_14293,N_14028);
nor U15364 (N_15364,N_14611,N_14507);
and U15365 (N_15365,N_13832,N_13761);
nand U15366 (N_15366,N_13666,N_13505);
and U15367 (N_15367,N_14253,N_14363);
nor U15368 (N_15368,N_14127,N_14333);
xnor U15369 (N_15369,N_13950,N_14913);
nand U15370 (N_15370,N_14798,N_13946);
nand U15371 (N_15371,N_13518,N_14623);
nor U15372 (N_15372,N_14980,N_14060);
xor U15373 (N_15373,N_14529,N_14756);
and U15374 (N_15374,N_14236,N_14561);
nand U15375 (N_15375,N_13606,N_13636);
nor U15376 (N_15376,N_14413,N_14521);
nor U15377 (N_15377,N_14417,N_14436);
nand U15378 (N_15378,N_14511,N_14368);
or U15379 (N_15379,N_14092,N_13703);
nand U15380 (N_15380,N_14917,N_14093);
and U15381 (N_15381,N_14384,N_14963);
xnor U15382 (N_15382,N_14977,N_14115);
and U15383 (N_15383,N_14929,N_14542);
xor U15384 (N_15384,N_14597,N_14892);
and U15385 (N_15385,N_14997,N_14304);
and U15386 (N_15386,N_14837,N_13930);
and U15387 (N_15387,N_14377,N_13875);
or U15388 (N_15388,N_13863,N_14978);
nand U15389 (N_15389,N_14734,N_14186);
or U15390 (N_15390,N_14036,N_14247);
and U15391 (N_15391,N_14947,N_14819);
nor U15392 (N_15392,N_14569,N_14965);
nand U15393 (N_15393,N_14074,N_13792);
nor U15394 (N_15394,N_14477,N_14101);
nor U15395 (N_15395,N_13718,N_14828);
or U15396 (N_15396,N_13998,N_14702);
and U15397 (N_15397,N_14224,N_14661);
or U15398 (N_15398,N_14717,N_14053);
nand U15399 (N_15399,N_13883,N_14640);
nor U15400 (N_15400,N_14380,N_14697);
or U15401 (N_15401,N_14787,N_14944);
nand U15402 (N_15402,N_14402,N_13515);
nand U15403 (N_15403,N_13868,N_13534);
nand U15404 (N_15404,N_14396,N_14311);
nor U15405 (N_15405,N_14668,N_13597);
nor U15406 (N_15406,N_14861,N_14047);
and U15407 (N_15407,N_14279,N_14735);
nor U15408 (N_15408,N_13988,N_13896);
xor U15409 (N_15409,N_13909,N_14390);
nand U15410 (N_15410,N_14446,N_14813);
nor U15411 (N_15411,N_14231,N_14655);
and U15412 (N_15412,N_14414,N_14372);
xnor U15413 (N_15413,N_14119,N_14073);
nand U15414 (N_15414,N_13537,N_14055);
xnor U15415 (N_15415,N_14182,N_14409);
nor U15416 (N_15416,N_14688,N_14087);
nor U15417 (N_15417,N_14498,N_14748);
and U15418 (N_15418,N_14690,N_13704);
nand U15419 (N_15419,N_14705,N_13958);
nor U15420 (N_15420,N_13879,N_13683);
xnor U15421 (N_15421,N_14811,N_13722);
xor U15422 (N_15422,N_13943,N_14560);
nor U15423 (N_15423,N_14801,N_14285);
and U15424 (N_15424,N_13964,N_14906);
or U15425 (N_15425,N_13975,N_14626);
nor U15426 (N_15426,N_14559,N_14464);
and U15427 (N_15427,N_14566,N_14306);
or U15428 (N_15428,N_14324,N_13512);
nand U15429 (N_15429,N_13545,N_14644);
and U15430 (N_15430,N_13577,N_14352);
nor U15431 (N_15431,N_14554,N_14199);
nor U15432 (N_15432,N_13595,N_14574);
and U15433 (N_15433,N_14548,N_14213);
xnor U15434 (N_15434,N_13787,N_13615);
xnor U15435 (N_15435,N_14764,N_14237);
and U15436 (N_15436,N_14657,N_14370);
nand U15437 (N_15437,N_14010,N_14975);
xnor U15438 (N_15438,N_14453,N_14987);
or U15439 (N_15439,N_13948,N_14955);
nor U15440 (N_15440,N_13669,N_13807);
and U15441 (N_15441,N_13602,N_14331);
nor U15442 (N_15442,N_14258,N_14388);
or U15443 (N_15443,N_13601,N_14897);
xnor U15444 (N_15444,N_13618,N_13758);
nor U15445 (N_15445,N_14849,N_14135);
nand U15446 (N_15446,N_14497,N_13940);
xnor U15447 (N_15447,N_14865,N_14588);
xor U15448 (N_15448,N_14085,N_14463);
xnor U15449 (N_15449,N_14926,N_14238);
or U15450 (N_15450,N_14041,N_13521);
nand U15451 (N_15451,N_13751,N_13777);
nand U15452 (N_15452,N_13555,N_13839);
and U15453 (N_15453,N_13580,N_13752);
nand U15454 (N_15454,N_14116,N_13586);
nand U15455 (N_15455,N_14273,N_14562);
nor U15456 (N_15456,N_13674,N_14122);
nor U15457 (N_15457,N_14763,N_14479);
and U15458 (N_15458,N_14772,N_14826);
or U15459 (N_15459,N_13530,N_14524);
nor U15460 (N_15460,N_13673,N_14181);
nor U15461 (N_15461,N_14750,N_14674);
nor U15462 (N_15462,N_14878,N_13578);
nor U15463 (N_15463,N_14886,N_14345);
or U15464 (N_15464,N_14180,N_14437);
or U15465 (N_15465,N_13657,N_14816);
nor U15466 (N_15466,N_13526,N_14632);
or U15467 (N_15467,N_13854,N_13598);
or U15468 (N_15468,N_13738,N_13945);
xor U15469 (N_15469,N_13702,N_13709);
xnor U15470 (N_15470,N_13587,N_14715);
nand U15471 (N_15471,N_14192,N_14209);
nand U15472 (N_15472,N_13913,N_14167);
and U15473 (N_15473,N_14610,N_14553);
or U15474 (N_15474,N_13973,N_14727);
and U15475 (N_15475,N_14441,N_14682);
xor U15476 (N_15476,N_13858,N_13769);
nand U15477 (N_15477,N_14812,N_14696);
xnor U15478 (N_15478,N_14843,N_14095);
and U15479 (N_15479,N_14329,N_14207);
nor U15480 (N_15480,N_14104,N_14086);
nand U15481 (N_15481,N_14287,N_14315);
nand U15482 (N_15482,N_13561,N_14707);
xor U15483 (N_15483,N_14706,N_14741);
and U15484 (N_15484,N_14503,N_13897);
and U15485 (N_15485,N_14342,N_13528);
and U15486 (N_15486,N_13663,N_14845);
nand U15487 (N_15487,N_14337,N_13692);
nor U15488 (N_15488,N_13982,N_14887);
xnor U15489 (N_15489,N_13914,N_13994);
or U15490 (N_15490,N_13726,N_13610);
or U15491 (N_15491,N_13907,N_14859);
or U15492 (N_15492,N_14885,N_14440);
and U15493 (N_15493,N_14283,N_14833);
xor U15494 (N_15494,N_14603,N_13736);
or U15495 (N_15495,N_14422,N_14779);
nor U15496 (N_15496,N_13926,N_13899);
xnor U15497 (N_15497,N_13590,N_14968);
nand U15498 (N_15498,N_14641,N_14647);
xor U15499 (N_15499,N_14305,N_14676);
nand U15500 (N_15500,N_13546,N_14487);
xnor U15501 (N_15501,N_14867,N_13735);
xnor U15502 (N_15502,N_14883,N_13981);
and U15503 (N_15503,N_13772,N_14365);
xnor U15504 (N_15504,N_14720,N_14307);
or U15505 (N_15505,N_14634,N_13638);
xnor U15506 (N_15506,N_13821,N_13729);
nor U15507 (N_15507,N_14716,N_14513);
nor U15508 (N_15508,N_14619,N_13723);
xnor U15509 (N_15509,N_13901,N_13962);
or U15510 (N_15510,N_14577,N_14587);
and U15511 (N_15511,N_14381,N_14550);
nand U15512 (N_15512,N_14002,N_13592);
nand U15513 (N_15513,N_13942,N_14468);
and U15514 (N_15514,N_14200,N_14004);
nor U15515 (N_15515,N_14635,N_14326);
xor U15516 (N_15516,N_14778,N_14695);
nor U15517 (N_15517,N_13717,N_14541);
and U15518 (N_15518,N_14701,N_14211);
or U15519 (N_15519,N_13608,N_14681);
xor U15520 (N_15520,N_14567,N_14703);
nand U15521 (N_15521,N_13786,N_14666);
xnor U15522 (N_15522,N_14401,N_13698);
and U15523 (N_15523,N_13880,N_14022);
or U15524 (N_15524,N_14999,N_13623);
xor U15525 (N_15525,N_14107,N_14355);
nand U15526 (N_15526,N_14045,N_14261);
xnor U15527 (N_15527,N_14361,N_13628);
xor U15528 (N_15528,N_14378,N_14033);
and U15529 (N_15529,N_14098,N_14075);
nor U15530 (N_15530,N_14161,N_13749);
nand U15531 (N_15531,N_13583,N_13775);
xor U15532 (N_15532,N_14653,N_14658);
nand U15533 (N_15533,N_13727,N_14950);
nand U15534 (N_15534,N_14482,N_14910);
xor U15535 (N_15535,N_14379,N_14799);
nor U15536 (N_15536,N_14492,N_13827);
nor U15537 (N_15537,N_14793,N_13811);
xor U15538 (N_15538,N_14724,N_14071);
or U15539 (N_15539,N_14072,N_13713);
nand U15540 (N_15540,N_13817,N_14144);
nand U15541 (N_15541,N_14460,N_13763);
or U15542 (N_15542,N_14633,N_14758);
nor U15543 (N_15543,N_14824,N_14530);
nand U15544 (N_15544,N_14347,N_14058);
xor U15545 (N_15545,N_14600,N_14840);
xnor U15546 (N_15546,N_13677,N_14234);
or U15547 (N_15547,N_14481,N_13870);
nor U15548 (N_15548,N_14700,N_13715);
xnor U15549 (N_15549,N_13582,N_14665);
nand U15550 (N_15550,N_14344,N_14904);
xor U15551 (N_15551,N_13971,N_14805);
or U15552 (N_15552,N_14340,N_13642);
nand U15553 (N_15553,N_14155,N_14032);
or U15554 (N_15554,N_14106,N_13895);
xor U15555 (N_15555,N_14031,N_13654);
xnor U15556 (N_15556,N_14493,N_13565);
or U15557 (N_15557,N_14451,N_14931);
or U15558 (N_15558,N_14357,N_14759);
nand U15559 (N_15559,N_13853,N_13823);
nand U15560 (N_15560,N_14916,N_13637);
xnor U15561 (N_15561,N_14117,N_13990);
nand U15562 (N_15562,N_13633,N_14501);
or U15563 (N_15563,N_13887,N_13812);
nand U15564 (N_15564,N_14895,N_14105);
nor U15565 (N_15565,N_14232,N_14286);
or U15566 (N_15566,N_14508,N_14038);
nand U15567 (N_15567,N_13538,N_14218);
xor U15568 (N_15568,N_13842,N_13774);
or U15569 (N_15569,N_14733,N_14585);
or U15570 (N_15570,N_13593,N_14991);
xor U15571 (N_15571,N_14589,N_14525);
and U15572 (N_15572,N_14903,N_13808);
xnor U15573 (N_15573,N_14515,N_14435);
nor U15574 (N_15574,N_14648,N_14919);
xnor U15575 (N_15575,N_13707,N_14320);
nand U15576 (N_15576,N_13922,N_13685);
xnor U15577 (N_15577,N_14215,N_14951);
nor U15578 (N_15578,N_14907,N_14930);
nor U15579 (N_15579,N_14118,N_14297);
and U15580 (N_15580,N_14547,N_14506);
or U15581 (N_15581,N_13734,N_13712);
nor U15582 (N_15582,N_14044,N_14328);
nor U15583 (N_15583,N_14683,N_14995);
nor U15584 (N_15584,N_14594,N_13830);
or U15585 (N_15585,N_14067,N_14392);
nor U15586 (N_15586,N_14516,N_14271);
xnor U15587 (N_15587,N_14680,N_14850);
nand U15588 (N_15588,N_14932,N_14608);
nand U15589 (N_15589,N_14628,N_13784);
nor U15590 (N_15590,N_14375,N_14517);
and U15591 (N_15591,N_13687,N_14620);
xor U15592 (N_15592,N_14013,N_14691);
or U15593 (N_15593,N_13799,N_14584);
and U15594 (N_15594,N_14855,N_14001);
xnor U15595 (N_15595,N_14249,N_13746);
nor U15596 (N_15596,N_14721,N_13984);
nor U15597 (N_15597,N_14725,N_13622);
nor U15598 (N_15598,N_14808,N_14847);
xor U15599 (N_15599,N_14775,N_14543);
nand U15600 (N_15600,N_14391,N_14992);
xor U15601 (N_15601,N_13603,N_14708);
and U15602 (N_15602,N_14834,N_14505);
nand U15603 (N_15603,N_14046,N_13754);
and U15604 (N_15604,N_14374,N_13568);
xnor U15605 (N_15605,N_14581,N_14795);
and U15606 (N_15606,N_14537,N_13564);
nand U15607 (N_15607,N_13551,N_14770);
or U15608 (N_15608,N_14896,N_14993);
or U15609 (N_15609,N_13877,N_13782);
nor U15610 (N_15610,N_14099,N_13995);
and U15611 (N_15611,N_13501,N_14670);
nand U15612 (N_15612,N_14596,N_13693);
and U15613 (N_15613,N_13906,N_14157);
nand U15614 (N_15614,N_13614,N_14364);
nor U15615 (N_15615,N_14967,N_14407);
nor U15616 (N_15616,N_14954,N_14406);
or U15617 (N_15617,N_13844,N_13989);
or U15618 (N_15618,N_14673,N_14539);
and U15619 (N_15619,N_13563,N_14404);
or U15620 (N_15620,N_13529,N_14268);
nand U15621 (N_15621,N_13604,N_14884);
and U15622 (N_15622,N_14433,N_13556);
or U15623 (N_15623,N_14645,N_13527);
xnor U15624 (N_15624,N_13985,N_14244);
nor U15625 (N_15625,N_14416,N_13670);
nand U15626 (N_15626,N_14179,N_14923);
nor U15627 (N_15627,N_14393,N_14270);
nor U15628 (N_15628,N_14191,N_13917);
or U15629 (N_15629,N_14486,N_14243);
nand U15630 (N_15630,N_14454,N_14838);
or U15631 (N_15631,N_13605,N_14153);
nand U15632 (N_15632,N_14070,N_13919);
nor U15633 (N_15633,N_13867,N_14979);
and U15634 (N_15634,N_14389,N_13540);
nor U15635 (N_15635,N_14252,N_14776);
xnor U15636 (N_15636,N_14900,N_13627);
nor U15637 (N_15637,N_13562,N_13960);
nand U15638 (N_15638,N_13690,N_14205);
nand U15639 (N_15639,N_14403,N_14866);
or U15640 (N_15640,N_14356,N_14617);
or U15641 (N_15641,N_13970,N_14336);
nand U15642 (N_15642,N_14149,N_14152);
and U15643 (N_15643,N_14719,N_13585);
nand U15644 (N_15644,N_14260,N_13974);
nand U15645 (N_15645,N_13888,N_14455);
and U15646 (N_15646,N_13745,N_14527);
nand U15647 (N_15647,N_14136,N_13641);
nand U15648 (N_15648,N_14160,N_13802);
nor U15649 (N_15649,N_13584,N_14902);
nor U15650 (N_15650,N_14142,N_14709);
nor U15651 (N_15651,N_13541,N_14225);
and U15652 (N_15652,N_13803,N_13724);
or U15653 (N_15653,N_14927,N_14124);
nor U15654 (N_15654,N_14156,N_14164);
and U15655 (N_15655,N_14810,N_14400);
xor U15656 (N_15656,N_13651,N_14465);
xnor U15657 (N_15657,N_14428,N_13655);
or U15658 (N_15658,N_14533,N_13753);
or U15659 (N_15659,N_13947,N_14314);
nor U15660 (N_15660,N_14476,N_14535);
and U15661 (N_15661,N_14187,N_14723);
or U15662 (N_15662,N_14514,N_14426);
or U15663 (N_15663,N_14312,N_14586);
nor U15664 (N_15664,N_14996,N_14698);
nor U15665 (N_15665,N_13872,N_14362);
xor U15666 (N_15666,N_14138,N_14399);
xnor U15667 (N_15667,N_14125,N_14789);
and U15668 (N_15668,N_14461,N_14558);
or U15669 (N_15669,N_14870,N_14025);
nor U15670 (N_15670,N_14056,N_13710);
and U15671 (N_15671,N_13934,N_14343);
or U15672 (N_15672,N_14957,N_14439);
or U15673 (N_15673,N_13889,N_14575);
or U15674 (N_15674,N_13959,N_13672);
and U15675 (N_15675,N_14512,N_14636);
nor U15676 (N_15676,N_13596,N_14565);
xor U15677 (N_15677,N_14990,N_14128);
nor U15678 (N_15678,N_14432,N_13531);
or U15679 (N_15679,N_13716,N_14360);
nand U15680 (N_15680,N_14601,N_14767);
or U15681 (N_15681,N_14475,N_14146);
or U15682 (N_15682,N_14835,N_14113);
and U15683 (N_15683,N_13779,N_14080);
nand U15684 (N_15684,N_14021,N_14078);
nand U15685 (N_15685,N_14765,N_14973);
and U15686 (N_15686,N_13699,N_14395);
nand U15687 (N_15687,N_13644,N_14862);
or U15688 (N_15688,N_14908,N_13898);
nand U15689 (N_15689,N_14607,N_14671);
xnor U15690 (N_15690,N_13806,N_14480);
nand U15691 (N_15691,N_14267,N_14660);
or U15692 (N_15692,N_14120,N_13794);
nor U15693 (N_15693,N_14945,N_13939);
and U15694 (N_15694,N_13796,N_14784);
nor U15695 (N_15695,N_14295,N_14651);
nand U15696 (N_15696,N_14251,N_13676);
nor U15697 (N_15697,N_13892,N_14677);
nor U15698 (N_15698,N_14531,N_14386);
and U15699 (N_15699,N_14823,N_14470);
xnor U15700 (N_15700,N_14744,N_14035);
xor U15701 (N_15701,N_13788,N_14321);
or U15702 (N_15702,N_14817,N_14739);
nand U15703 (N_15703,N_14888,N_13756);
and U15704 (N_15704,N_14893,N_13768);
or U15705 (N_15705,N_13996,N_14972);
nor U15706 (N_15706,N_14899,N_14743);
xor U15707 (N_15707,N_13600,N_14369);
and U15708 (N_15708,N_13849,N_14557);
nand U15709 (N_15709,N_13847,N_14029);
and U15710 (N_15710,N_14316,N_14289);
nand U15711 (N_15711,N_14580,N_13684);
or U15712 (N_15712,N_14255,N_13859);
or U15713 (N_15713,N_14005,N_14622);
nand U15714 (N_15714,N_14387,N_13968);
or U15715 (N_15715,N_14571,N_13539);
or U15716 (N_15716,N_14604,N_13773);
nand U15717 (N_15717,N_14335,N_13547);
and U15718 (N_15718,N_14054,N_13900);
nor U15719 (N_15719,N_14846,N_14606);
nor U15720 (N_15720,N_14854,N_14449);
xnor U15721 (N_15721,N_14265,N_13509);
and U15722 (N_15722,N_14457,N_14195);
xor U15723 (N_15723,N_14922,N_13835);
nand U15724 (N_15724,N_14637,N_13795);
nor U15725 (N_15725,N_13834,N_14012);
nor U15726 (N_15726,N_13681,N_13903);
xor U15727 (N_15727,N_14549,N_14256);
and U15728 (N_15728,N_13532,N_13740);
nor U15729 (N_15729,N_13856,N_13575);
xnor U15730 (N_15730,N_14206,N_13874);
xor U15731 (N_15731,N_14111,N_13728);
nand U15732 (N_15732,N_13987,N_14383);
nand U15733 (N_15733,N_14591,N_13937);
xor U15734 (N_15734,N_13730,N_14059);
and U15735 (N_15735,N_13502,N_13747);
xnor U15736 (N_15736,N_14540,N_13961);
nor U15737 (N_15737,N_13656,N_14318);
or U15738 (N_15738,N_14083,N_13525);
and U15739 (N_15739,N_14857,N_14652);
nor U15740 (N_15740,N_14110,N_14970);
and U15741 (N_15741,N_14650,N_14962);
and U15742 (N_15742,N_14174,N_14274);
and U15743 (N_15743,N_14728,N_14430);
or U15744 (N_15744,N_14472,N_14313);
and U15745 (N_15745,N_14986,N_13828);
nor U15746 (N_15746,N_14227,N_13865);
xnor U15747 (N_15747,N_14408,N_14024);
nand U15748 (N_15748,N_14678,N_14692);
xnor U15749 (N_15749,N_13550,N_13824);
and U15750 (N_15750,N_13908,N_13789);
and U15751 (N_15751,N_14334,N_13575);
xnor U15752 (N_15752,N_13757,N_14389);
or U15753 (N_15753,N_14154,N_13793);
nor U15754 (N_15754,N_13611,N_13740);
nand U15755 (N_15755,N_14026,N_13687);
and U15756 (N_15756,N_14319,N_14234);
and U15757 (N_15757,N_14217,N_14897);
and U15758 (N_15758,N_14670,N_13737);
or U15759 (N_15759,N_13552,N_13885);
and U15760 (N_15760,N_14187,N_13652);
and U15761 (N_15761,N_14443,N_14111);
xor U15762 (N_15762,N_13749,N_14368);
and U15763 (N_15763,N_14255,N_13753);
or U15764 (N_15764,N_14343,N_14581);
xor U15765 (N_15765,N_14579,N_13970);
nor U15766 (N_15766,N_14172,N_13727);
or U15767 (N_15767,N_14240,N_14652);
and U15768 (N_15768,N_14145,N_14261);
and U15769 (N_15769,N_13513,N_14027);
or U15770 (N_15770,N_13852,N_13641);
and U15771 (N_15771,N_13625,N_13973);
and U15772 (N_15772,N_14380,N_13799);
nor U15773 (N_15773,N_14059,N_14902);
xnor U15774 (N_15774,N_14302,N_13931);
or U15775 (N_15775,N_13641,N_13920);
or U15776 (N_15776,N_13539,N_14450);
nor U15777 (N_15777,N_13539,N_13909);
nor U15778 (N_15778,N_14389,N_13817);
nand U15779 (N_15779,N_14228,N_14634);
or U15780 (N_15780,N_14837,N_13881);
nor U15781 (N_15781,N_13807,N_14077);
xnor U15782 (N_15782,N_14883,N_14157);
xor U15783 (N_15783,N_14998,N_13818);
xnor U15784 (N_15784,N_13746,N_14745);
and U15785 (N_15785,N_13939,N_14039);
and U15786 (N_15786,N_14070,N_14882);
xnor U15787 (N_15787,N_13867,N_13725);
xnor U15788 (N_15788,N_14506,N_14856);
nand U15789 (N_15789,N_13852,N_13841);
xnor U15790 (N_15790,N_13888,N_14639);
xnor U15791 (N_15791,N_13635,N_14742);
xnor U15792 (N_15792,N_14655,N_14351);
nand U15793 (N_15793,N_14598,N_14526);
and U15794 (N_15794,N_14411,N_13998);
nor U15795 (N_15795,N_13763,N_14742);
nand U15796 (N_15796,N_14581,N_14255);
nand U15797 (N_15797,N_14579,N_13568);
nor U15798 (N_15798,N_13983,N_14138);
and U15799 (N_15799,N_14593,N_14763);
and U15800 (N_15800,N_14901,N_13629);
or U15801 (N_15801,N_14711,N_14692);
nor U15802 (N_15802,N_13596,N_13792);
nor U15803 (N_15803,N_14245,N_14411);
or U15804 (N_15804,N_14621,N_14879);
nor U15805 (N_15805,N_14768,N_14330);
or U15806 (N_15806,N_13754,N_14305);
or U15807 (N_15807,N_14180,N_14990);
xor U15808 (N_15808,N_14499,N_14455);
xor U15809 (N_15809,N_13710,N_13833);
nor U15810 (N_15810,N_14183,N_13656);
nor U15811 (N_15811,N_14152,N_14857);
or U15812 (N_15812,N_14414,N_14994);
or U15813 (N_15813,N_14767,N_14048);
nand U15814 (N_15814,N_14575,N_14794);
and U15815 (N_15815,N_14299,N_14922);
nand U15816 (N_15816,N_14128,N_14303);
nand U15817 (N_15817,N_14891,N_14556);
or U15818 (N_15818,N_14320,N_14877);
and U15819 (N_15819,N_14219,N_14141);
and U15820 (N_15820,N_14958,N_13964);
and U15821 (N_15821,N_13632,N_13606);
xnor U15822 (N_15822,N_14780,N_13913);
or U15823 (N_15823,N_14688,N_14329);
xnor U15824 (N_15824,N_14536,N_13747);
and U15825 (N_15825,N_13934,N_14817);
nor U15826 (N_15826,N_13933,N_13891);
or U15827 (N_15827,N_14425,N_14849);
nor U15828 (N_15828,N_13620,N_13531);
or U15829 (N_15829,N_13934,N_14807);
xnor U15830 (N_15830,N_14184,N_14567);
xor U15831 (N_15831,N_13650,N_14553);
nand U15832 (N_15832,N_14053,N_14126);
xor U15833 (N_15833,N_14374,N_13940);
and U15834 (N_15834,N_13554,N_14775);
and U15835 (N_15835,N_14189,N_14832);
or U15836 (N_15836,N_14416,N_13735);
nor U15837 (N_15837,N_14231,N_13512);
nand U15838 (N_15838,N_14381,N_14084);
xnor U15839 (N_15839,N_14306,N_13987);
nand U15840 (N_15840,N_13866,N_14455);
xnor U15841 (N_15841,N_14432,N_14747);
nand U15842 (N_15842,N_13551,N_13993);
xor U15843 (N_15843,N_14453,N_14711);
xor U15844 (N_15844,N_13884,N_14167);
and U15845 (N_15845,N_14622,N_14230);
nand U15846 (N_15846,N_13690,N_14523);
xnor U15847 (N_15847,N_14565,N_14318);
xnor U15848 (N_15848,N_13957,N_14828);
nand U15849 (N_15849,N_13876,N_14508);
nand U15850 (N_15850,N_13999,N_14857);
nor U15851 (N_15851,N_13565,N_14490);
xnor U15852 (N_15852,N_14883,N_14220);
or U15853 (N_15853,N_14167,N_13780);
xor U15854 (N_15854,N_14424,N_14758);
or U15855 (N_15855,N_13719,N_13984);
xor U15856 (N_15856,N_13919,N_14984);
or U15857 (N_15857,N_14283,N_14256);
nor U15858 (N_15858,N_14689,N_13632);
or U15859 (N_15859,N_13796,N_13743);
nand U15860 (N_15860,N_14415,N_14407);
xor U15861 (N_15861,N_14389,N_14338);
nor U15862 (N_15862,N_14066,N_13561);
nor U15863 (N_15863,N_14233,N_14615);
or U15864 (N_15864,N_14071,N_13709);
and U15865 (N_15865,N_13595,N_14291);
nor U15866 (N_15866,N_13623,N_13510);
nor U15867 (N_15867,N_14697,N_14595);
xnor U15868 (N_15868,N_13766,N_13927);
or U15869 (N_15869,N_14755,N_14418);
and U15870 (N_15870,N_14839,N_13871);
nor U15871 (N_15871,N_14326,N_13620);
nor U15872 (N_15872,N_14327,N_14429);
nor U15873 (N_15873,N_14297,N_13813);
and U15874 (N_15874,N_14346,N_14864);
nand U15875 (N_15875,N_14560,N_14423);
or U15876 (N_15876,N_13939,N_13959);
nand U15877 (N_15877,N_14005,N_14033);
nor U15878 (N_15878,N_14340,N_14166);
or U15879 (N_15879,N_13895,N_14481);
nand U15880 (N_15880,N_13983,N_14448);
or U15881 (N_15881,N_13932,N_14597);
or U15882 (N_15882,N_14320,N_14590);
nor U15883 (N_15883,N_14114,N_14278);
nor U15884 (N_15884,N_14482,N_14780);
xor U15885 (N_15885,N_14061,N_14862);
and U15886 (N_15886,N_14578,N_14721);
nor U15887 (N_15887,N_14472,N_14033);
xnor U15888 (N_15888,N_14640,N_14358);
or U15889 (N_15889,N_13673,N_14102);
nand U15890 (N_15890,N_14744,N_14528);
and U15891 (N_15891,N_13767,N_14859);
xor U15892 (N_15892,N_14502,N_14484);
nor U15893 (N_15893,N_14134,N_14155);
xor U15894 (N_15894,N_14588,N_14358);
nand U15895 (N_15895,N_13755,N_13955);
nor U15896 (N_15896,N_13620,N_14572);
nand U15897 (N_15897,N_13617,N_14559);
nor U15898 (N_15898,N_13785,N_14961);
or U15899 (N_15899,N_13840,N_13901);
xor U15900 (N_15900,N_13597,N_13556);
and U15901 (N_15901,N_13804,N_13626);
xor U15902 (N_15902,N_13777,N_14534);
xnor U15903 (N_15903,N_13845,N_14050);
nand U15904 (N_15904,N_14148,N_14006);
xnor U15905 (N_15905,N_14264,N_14517);
nand U15906 (N_15906,N_14756,N_14100);
or U15907 (N_15907,N_14548,N_14701);
or U15908 (N_15908,N_14585,N_14458);
xor U15909 (N_15909,N_14253,N_14702);
xnor U15910 (N_15910,N_14808,N_14630);
and U15911 (N_15911,N_13566,N_14484);
or U15912 (N_15912,N_14818,N_14267);
nand U15913 (N_15913,N_14699,N_14448);
nand U15914 (N_15914,N_14956,N_13841);
and U15915 (N_15915,N_13649,N_14589);
nor U15916 (N_15916,N_13685,N_14900);
xnor U15917 (N_15917,N_14990,N_13821);
and U15918 (N_15918,N_14570,N_13534);
nor U15919 (N_15919,N_14670,N_13718);
and U15920 (N_15920,N_14449,N_14508);
xnor U15921 (N_15921,N_13630,N_14412);
and U15922 (N_15922,N_14464,N_14465);
nand U15923 (N_15923,N_14300,N_13929);
nor U15924 (N_15924,N_14578,N_13651);
xnor U15925 (N_15925,N_13913,N_14941);
xnor U15926 (N_15926,N_14522,N_14326);
nor U15927 (N_15927,N_13705,N_14955);
and U15928 (N_15928,N_14514,N_13593);
xnor U15929 (N_15929,N_14017,N_14069);
nor U15930 (N_15930,N_13959,N_14082);
nand U15931 (N_15931,N_14011,N_14791);
nand U15932 (N_15932,N_14923,N_14343);
nand U15933 (N_15933,N_14918,N_13769);
nor U15934 (N_15934,N_13928,N_14653);
nand U15935 (N_15935,N_13783,N_13936);
and U15936 (N_15936,N_14827,N_13863);
and U15937 (N_15937,N_14170,N_14184);
nand U15938 (N_15938,N_14842,N_13653);
xnor U15939 (N_15939,N_14970,N_14260);
and U15940 (N_15940,N_13926,N_14479);
nor U15941 (N_15941,N_14167,N_14943);
or U15942 (N_15942,N_14780,N_14114);
and U15943 (N_15943,N_13623,N_14858);
or U15944 (N_15944,N_14269,N_14434);
nor U15945 (N_15945,N_13691,N_14714);
nand U15946 (N_15946,N_13792,N_14911);
nor U15947 (N_15947,N_14641,N_14526);
and U15948 (N_15948,N_14706,N_13892);
nor U15949 (N_15949,N_14651,N_13584);
or U15950 (N_15950,N_14582,N_13607);
and U15951 (N_15951,N_14343,N_14549);
and U15952 (N_15952,N_14956,N_14385);
xor U15953 (N_15953,N_14475,N_13653);
xor U15954 (N_15954,N_14199,N_14035);
and U15955 (N_15955,N_14017,N_14712);
and U15956 (N_15956,N_13674,N_14800);
nand U15957 (N_15957,N_13555,N_14806);
and U15958 (N_15958,N_14565,N_13551);
nor U15959 (N_15959,N_13769,N_14129);
nand U15960 (N_15960,N_14330,N_14294);
nor U15961 (N_15961,N_14178,N_14325);
nor U15962 (N_15962,N_14618,N_13802);
or U15963 (N_15963,N_14119,N_14195);
and U15964 (N_15964,N_14225,N_13873);
or U15965 (N_15965,N_13726,N_14231);
nand U15966 (N_15966,N_14705,N_13722);
or U15967 (N_15967,N_14038,N_13929);
nor U15968 (N_15968,N_14018,N_13956);
xor U15969 (N_15969,N_14610,N_14085);
or U15970 (N_15970,N_13558,N_14440);
and U15971 (N_15971,N_13687,N_13908);
xor U15972 (N_15972,N_14434,N_14234);
xnor U15973 (N_15973,N_14079,N_14091);
nand U15974 (N_15974,N_14881,N_14707);
and U15975 (N_15975,N_14886,N_13679);
and U15976 (N_15976,N_14821,N_13591);
or U15977 (N_15977,N_14120,N_14956);
or U15978 (N_15978,N_14191,N_14585);
nand U15979 (N_15979,N_14657,N_14197);
or U15980 (N_15980,N_14079,N_14524);
and U15981 (N_15981,N_14670,N_13525);
and U15982 (N_15982,N_14953,N_14146);
and U15983 (N_15983,N_14361,N_14259);
xor U15984 (N_15984,N_14818,N_14456);
or U15985 (N_15985,N_14857,N_13558);
or U15986 (N_15986,N_13878,N_14631);
nand U15987 (N_15987,N_14017,N_14317);
nand U15988 (N_15988,N_13758,N_13705);
and U15989 (N_15989,N_14609,N_13624);
nor U15990 (N_15990,N_13504,N_14475);
nand U15991 (N_15991,N_14764,N_14059);
and U15992 (N_15992,N_14312,N_14842);
nand U15993 (N_15993,N_14890,N_14842);
nand U15994 (N_15994,N_13579,N_14435);
or U15995 (N_15995,N_14396,N_14855);
xnor U15996 (N_15996,N_13653,N_13697);
xor U15997 (N_15997,N_14897,N_13590);
xor U15998 (N_15998,N_14022,N_14389);
xor U15999 (N_15999,N_13700,N_14247);
and U16000 (N_16000,N_14187,N_14952);
nand U16001 (N_16001,N_14512,N_13539);
nand U16002 (N_16002,N_14092,N_13960);
and U16003 (N_16003,N_14434,N_14266);
xnor U16004 (N_16004,N_14033,N_14949);
nor U16005 (N_16005,N_14212,N_14250);
nand U16006 (N_16006,N_13887,N_13748);
nor U16007 (N_16007,N_13515,N_14698);
or U16008 (N_16008,N_14546,N_13872);
xor U16009 (N_16009,N_14473,N_14199);
xor U16010 (N_16010,N_13940,N_14975);
xnor U16011 (N_16011,N_13685,N_14787);
and U16012 (N_16012,N_14570,N_14207);
xnor U16013 (N_16013,N_13719,N_13644);
nand U16014 (N_16014,N_13920,N_14233);
nand U16015 (N_16015,N_14051,N_14818);
xor U16016 (N_16016,N_14181,N_13553);
xnor U16017 (N_16017,N_13689,N_13855);
and U16018 (N_16018,N_14801,N_14985);
and U16019 (N_16019,N_14892,N_14956);
or U16020 (N_16020,N_14633,N_14938);
and U16021 (N_16021,N_14254,N_14988);
nor U16022 (N_16022,N_13519,N_13631);
xnor U16023 (N_16023,N_13770,N_13855);
nor U16024 (N_16024,N_14025,N_14253);
nor U16025 (N_16025,N_13868,N_14017);
xnor U16026 (N_16026,N_14271,N_14270);
nand U16027 (N_16027,N_14916,N_14632);
or U16028 (N_16028,N_14970,N_13699);
nand U16029 (N_16029,N_14156,N_13953);
nor U16030 (N_16030,N_13539,N_14962);
and U16031 (N_16031,N_14744,N_14151);
and U16032 (N_16032,N_14365,N_13755);
and U16033 (N_16033,N_14443,N_14653);
and U16034 (N_16034,N_14167,N_13790);
and U16035 (N_16035,N_14980,N_14480);
and U16036 (N_16036,N_14752,N_14938);
and U16037 (N_16037,N_14078,N_13630);
nand U16038 (N_16038,N_13574,N_14047);
nor U16039 (N_16039,N_14624,N_14161);
xor U16040 (N_16040,N_14345,N_13851);
or U16041 (N_16041,N_14364,N_13826);
nand U16042 (N_16042,N_14445,N_14930);
nand U16043 (N_16043,N_14962,N_13807);
xnor U16044 (N_16044,N_14167,N_13725);
and U16045 (N_16045,N_13988,N_14591);
xnor U16046 (N_16046,N_13906,N_14328);
or U16047 (N_16047,N_13511,N_14335);
or U16048 (N_16048,N_13600,N_14213);
and U16049 (N_16049,N_14961,N_14445);
or U16050 (N_16050,N_13991,N_13939);
xnor U16051 (N_16051,N_14751,N_14082);
xnor U16052 (N_16052,N_13825,N_13799);
and U16053 (N_16053,N_13521,N_13896);
nor U16054 (N_16054,N_13602,N_13766);
and U16055 (N_16055,N_14183,N_13532);
nor U16056 (N_16056,N_14912,N_14669);
or U16057 (N_16057,N_13726,N_14876);
nand U16058 (N_16058,N_14960,N_14276);
nor U16059 (N_16059,N_13838,N_13940);
or U16060 (N_16060,N_14264,N_14605);
or U16061 (N_16061,N_14363,N_14861);
and U16062 (N_16062,N_14130,N_13580);
and U16063 (N_16063,N_13532,N_14684);
nand U16064 (N_16064,N_14079,N_14897);
or U16065 (N_16065,N_14159,N_13999);
nor U16066 (N_16066,N_13920,N_13769);
nand U16067 (N_16067,N_14772,N_14967);
nand U16068 (N_16068,N_14476,N_14489);
nor U16069 (N_16069,N_14831,N_13862);
xnor U16070 (N_16070,N_14128,N_14961);
and U16071 (N_16071,N_14975,N_14188);
xnor U16072 (N_16072,N_13715,N_14042);
and U16073 (N_16073,N_13505,N_14401);
nand U16074 (N_16074,N_14295,N_13626);
and U16075 (N_16075,N_14066,N_14312);
nand U16076 (N_16076,N_14459,N_14056);
nand U16077 (N_16077,N_13710,N_14188);
or U16078 (N_16078,N_14690,N_13886);
xor U16079 (N_16079,N_14243,N_14197);
or U16080 (N_16080,N_13753,N_13923);
nor U16081 (N_16081,N_13643,N_14042);
and U16082 (N_16082,N_14617,N_14445);
and U16083 (N_16083,N_14542,N_14628);
xnor U16084 (N_16084,N_13874,N_14664);
nand U16085 (N_16085,N_13737,N_14252);
nand U16086 (N_16086,N_13809,N_14593);
and U16087 (N_16087,N_14739,N_14331);
nand U16088 (N_16088,N_14421,N_13861);
and U16089 (N_16089,N_14806,N_13893);
and U16090 (N_16090,N_14996,N_13507);
nand U16091 (N_16091,N_13535,N_14735);
nor U16092 (N_16092,N_14357,N_14648);
nor U16093 (N_16093,N_14159,N_14126);
nand U16094 (N_16094,N_14592,N_14185);
xor U16095 (N_16095,N_14959,N_14125);
and U16096 (N_16096,N_13723,N_14605);
nor U16097 (N_16097,N_14972,N_14387);
nand U16098 (N_16098,N_13538,N_14115);
and U16099 (N_16099,N_14393,N_13664);
xor U16100 (N_16100,N_13894,N_14229);
nor U16101 (N_16101,N_13686,N_14959);
xor U16102 (N_16102,N_14513,N_13615);
nand U16103 (N_16103,N_14890,N_13705);
xor U16104 (N_16104,N_14924,N_13822);
nand U16105 (N_16105,N_14009,N_14460);
and U16106 (N_16106,N_14464,N_13606);
or U16107 (N_16107,N_14884,N_13528);
nand U16108 (N_16108,N_14155,N_14649);
and U16109 (N_16109,N_13730,N_14224);
nand U16110 (N_16110,N_14990,N_13863);
xnor U16111 (N_16111,N_14435,N_13520);
nand U16112 (N_16112,N_14522,N_14253);
nand U16113 (N_16113,N_13773,N_13873);
nor U16114 (N_16114,N_14156,N_14010);
or U16115 (N_16115,N_14507,N_14642);
or U16116 (N_16116,N_13527,N_14386);
or U16117 (N_16117,N_14957,N_13557);
or U16118 (N_16118,N_14181,N_14629);
and U16119 (N_16119,N_13731,N_14953);
and U16120 (N_16120,N_14367,N_14362);
nand U16121 (N_16121,N_14145,N_14098);
nand U16122 (N_16122,N_13756,N_14279);
or U16123 (N_16123,N_14851,N_14083);
or U16124 (N_16124,N_14470,N_13717);
nor U16125 (N_16125,N_14212,N_14229);
nor U16126 (N_16126,N_13558,N_14964);
xnor U16127 (N_16127,N_13920,N_13658);
xnor U16128 (N_16128,N_14130,N_14834);
xor U16129 (N_16129,N_14402,N_13683);
nand U16130 (N_16130,N_13820,N_14145);
or U16131 (N_16131,N_14670,N_14889);
nor U16132 (N_16132,N_13648,N_13709);
nor U16133 (N_16133,N_14480,N_14644);
nor U16134 (N_16134,N_14707,N_13876);
xnor U16135 (N_16135,N_14129,N_14959);
and U16136 (N_16136,N_14277,N_13830);
or U16137 (N_16137,N_14439,N_14740);
or U16138 (N_16138,N_14887,N_14555);
nand U16139 (N_16139,N_13530,N_14722);
xor U16140 (N_16140,N_13608,N_14918);
nand U16141 (N_16141,N_14101,N_14308);
nand U16142 (N_16142,N_14433,N_14124);
and U16143 (N_16143,N_13772,N_14497);
and U16144 (N_16144,N_14084,N_13578);
xnor U16145 (N_16145,N_14251,N_14695);
and U16146 (N_16146,N_14935,N_13668);
nand U16147 (N_16147,N_14432,N_13523);
nor U16148 (N_16148,N_14220,N_13630);
xor U16149 (N_16149,N_14314,N_14449);
xnor U16150 (N_16150,N_13611,N_14686);
xor U16151 (N_16151,N_14519,N_14698);
and U16152 (N_16152,N_13580,N_13518);
xor U16153 (N_16153,N_14370,N_14842);
and U16154 (N_16154,N_14935,N_14897);
and U16155 (N_16155,N_13791,N_13969);
or U16156 (N_16156,N_13772,N_13919);
and U16157 (N_16157,N_14539,N_14909);
nand U16158 (N_16158,N_14898,N_13625);
or U16159 (N_16159,N_14876,N_14840);
xnor U16160 (N_16160,N_14123,N_13580);
nand U16161 (N_16161,N_13805,N_13669);
and U16162 (N_16162,N_14550,N_13641);
and U16163 (N_16163,N_14300,N_14014);
or U16164 (N_16164,N_13977,N_14384);
or U16165 (N_16165,N_13648,N_13952);
or U16166 (N_16166,N_13594,N_14932);
xnor U16167 (N_16167,N_14911,N_13970);
xor U16168 (N_16168,N_14668,N_14549);
and U16169 (N_16169,N_14231,N_13686);
nor U16170 (N_16170,N_14574,N_14970);
and U16171 (N_16171,N_14590,N_13870);
nor U16172 (N_16172,N_14385,N_13699);
or U16173 (N_16173,N_14183,N_14584);
nor U16174 (N_16174,N_14502,N_14041);
and U16175 (N_16175,N_13987,N_14580);
and U16176 (N_16176,N_14989,N_14195);
or U16177 (N_16177,N_14767,N_14482);
and U16178 (N_16178,N_13862,N_14564);
and U16179 (N_16179,N_13568,N_13758);
nor U16180 (N_16180,N_14161,N_14901);
nand U16181 (N_16181,N_14442,N_14449);
or U16182 (N_16182,N_13882,N_14913);
nor U16183 (N_16183,N_14437,N_13919);
nor U16184 (N_16184,N_14936,N_14154);
xor U16185 (N_16185,N_14655,N_14483);
xnor U16186 (N_16186,N_13500,N_14700);
and U16187 (N_16187,N_13613,N_13500);
or U16188 (N_16188,N_14080,N_14569);
xnor U16189 (N_16189,N_14510,N_14672);
nor U16190 (N_16190,N_13906,N_14545);
nor U16191 (N_16191,N_13698,N_14963);
nor U16192 (N_16192,N_14255,N_14752);
nand U16193 (N_16193,N_13769,N_14413);
nand U16194 (N_16194,N_13516,N_13968);
and U16195 (N_16195,N_14547,N_14988);
nor U16196 (N_16196,N_14980,N_14741);
and U16197 (N_16197,N_14702,N_13784);
xor U16198 (N_16198,N_14977,N_13942);
xor U16199 (N_16199,N_14887,N_13833);
xor U16200 (N_16200,N_13978,N_13844);
and U16201 (N_16201,N_14748,N_13669);
or U16202 (N_16202,N_14599,N_14767);
nor U16203 (N_16203,N_13865,N_14734);
nor U16204 (N_16204,N_14242,N_14765);
or U16205 (N_16205,N_14100,N_14598);
nor U16206 (N_16206,N_13739,N_14484);
nor U16207 (N_16207,N_14646,N_14267);
and U16208 (N_16208,N_14221,N_14027);
xnor U16209 (N_16209,N_14812,N_14286);
nand U16210 (N_16210,N_13685,N_14180);
and U16211 (N_16211,N_13977,N_14744);
nand U16212 (N_16212,N_14100,N_14026);
nand U16213 (N_16213,N_13586,N_14429);
xnor U16214 (N_16214,N_14018,N_13840);
and U16215 (N_16215,N_14342,N_13965);
nor U16216 (N_16216,N_14030,N_14041);
nand U16217 (N_16217,N_14270,N_14822);
xor U16218 (N_16218,N_14617,N_13753);
nor U16219 (N_16219,N_14555,N_14779);
nor U16220 (N_16220,N_14427,N_14964);
or U16221 (N_16221,N_14939,N_14768);
or U16222 (N_16222,N_13752,N_14794);
or U16223 (N_16223,N_14458,N_13554);
and U16224 (N_16224,N_13566,N_14979);
nand U16225 (N_16225,N_14314,N_14490);
and U16226 (N_16226,N_14529,N_13635);
or U16227 (N_16227,N_14003,N_14593);
or U16228 (N_16228,N_14869,N_14109);
and U16229 (N_16229,N_14083,N_13752);
and U16230 (N_16230,N_14169,N_13837);
nor U16231 (N_16231,N_14207,N_14367);
or U16232 (N_16232,N_13807,N_14426);
xnor U16233 (N_16233,N_14847,N_14980);
nand U16234 (N_16234,N_14251,N_14857);
and U16235 (N_16235,N_13674,N_14999);
nand U16236 (N_16236,N_14657,N_14130);
nand U16237 (N_16237,N_14982,N_13726);
nand U16238 (N_16238,N_14216,N_14140);
and U16239 (N_16239,N_14229,N_14405);
or U16240 (N_16240,N_13624,N_14622);
nand U16241 (N_16241,N_14970,N_13807);
xnor U16242 (N_16242,N_14757,N_14422);
xnor U16243 (N_16243,N_13565,N_14346);
or U16244 (N_16244,N_14425,N_14256);
or U16245 (N_16245,N_13938,N_14550);
and U16246 (N_16246,N_14797,N_14176);
or U16247 (N_16247,N_14487,N_13637);
nor U16248 (N_16248,N_13985,N_13784);
nor U16249 (N_16249,N_13977,N_13921);
or U16250 (N_16250,N_14863,N_14050);
nand U16251 (N_16251,N_14708,N_14897);
nor U16252 (N_16252,N_14657,N_13786);
nor U16253 (N_16253,N_13972,N_14630);
nor U16254 (N_16254,N_13701,N_13870);
xnor U16255 (N_16255,N_14019,N_14942);
xnor U16256 (N_16256,N_14649,N_14303);
xnor U16257 (N_16257,N_14171,N_14856);
xor U16258 (N_16258,N_14373,N_13819);
nand U16259 (N_16259,N_14411,N_13939);
nand U16260 (N_16260,N_14630,N_14393);
and U16261 (N_16261,N_14553,N_13693);
or U16262 (N_16262,N_14763,N_13595);
xnor U16263 (N_16263,N_13933,N_14501);
and U16264 (N_16264,N_13869,N_14125);
and U16265 (N_16265,N_13826,N_13559);
nor U16266 (N_16266,N_14201,N_14664);
nor U16267 (N_16267,N_14823,N_14988);
nor U16268 (N_16268,N_13791,N_14521);
nor U16269 (N_16269,N_14565,N_13897);
nor U16270 (N_16270,N_14802,N_14684);
and U16271 (N_16271,N_14140,N_14790);
xor U16272 (N_16272,N_14654,N_14075);
or U16273 (N_16273,N_13660,N_14800);
nor U16274 (N_16274,N_14990,N_13865);
xnor U16275 (N_16275,N_13700,N_13621);
nor U16276 (N_16276,N_14617,N_14241);
or U16277 (N_16277,N_14760,N_14244);
or U16278 (N_16278,N_13638,N_14309);
xor U16279 (N_16279,N_13910,N_14054);
nor U16280 (N_16280,N_13761,N_14915);
xnor U16281 (N_16281,N_14621,N_14640);
or U16282 (N_16282,N_14910,N_14389);
nor U16283 (N_16283,N_14319,N_14105);
and U16284 (N_16284,N_13920,N_13695);
nand U16285 (N_16285,N_14364,N_14045);
nand U16286 (N_16286,N_13585,N_14289);
xor U16287 (N_16287,N_13630,N_13694);
nand U16288 (N_16288,N_14898,N_13646);
or U16289 (N_16289,N_14288,N_14010);
nand U16290 (N_16290,N_14296,N_14231);
and U16291 (N_16291,N_13812,N_13711);
nor U16292 (N_16292,N_14915,N_13725);
xor U16293 (N_16293,N_14652,N_14952);
xor U16294 (N_16294,N_14799,N_14579);
or U16295 (N_16295,N_14018,N_14647);
and U16296 (N_16296,N_14066,N_14893);
nor U16297 (N_16297,N_14381,N_14302);
and U16298 (N_16298,N_14187,N_14563);
and U16299 (N_16299,N_14234,N_13985);
nor U16300 (N_16300,N_14554,N_13686);
and U16301 (N_16301,N_14851,N_14814);
and U16302 (N_16302,N_13959,N_14397);
nand U16303 (N_16303,N_14648,N_14166);
or U16304 (N_16304,N_14772,N_14376);
xor U16305 (N_16305,N_13930,N_13936);
and U16306 (N_16306,N_14978,N_14152);
or U16307 (N_16307,N_14186,N_14609);
nand U16308 (N_16308,N_14766,N_14955);
nor U16309 (N_16309,N_14433,N_14988);
xor U16310 (N_16310,N_13524,N_13747);
and U16311 (N_16311,N_14737,N_13868);
or U16312 (N_16312,N_14118,N_13952);
xor U16313 (N_16313,N_13747,N_14067);
or U16314 (N_16314,N_14906,N_14031);
or U16315 (N_16315,N_13635,N_14673);
xnor U16316 (N_16316,N_14496,N_14086);
nor U16317 (N_16317,N_14200,N_13631);
nand U16318 (N_16318,N_13804,N_13766);
nand U16319 (N_16319,N_14574,N_13654);
nor U16320 (N_16320,N_14897,N_14015);
xnor U16321 (N_16321,N_14208,N_13827);
nand U16322 (N_16322,N_14201,N_14417);
xor U16323 (N_16323,N_13995,N_14740);
nand U16324 (N_16324,N_14271,N_14071);
and U16325 (N_16325,N_14222,N_14383);
nor U16326 (N_16326,N_14747,N_14922);
nand U16327 (N_16327,N_13704,N_14210);
or U16328 (N_16328,N_14120,N_14305);
or U16329 (N_16329,N_14867,N_14299);
xnor U16330 (N_16330,N_14404,N_14919);
nand U16331 (N_16331,N_14905,N_14505);
nand U16332 (N_16332,N_13615,N_14254);
or U16333 (N_16333,N_13543,N_14398);
or U16334 (N_16334,N_14219,N_13582);
xnor U16335 (N_16335,N_14755,N_14332);
xor U16336 (N_16336,N_13550,N_14226);
and U16337 (N_16337,N_13621,N_14587);
and U16338 (N_16338,N_13899,N_13563);
or U16339 (N_16339,N_13919,N_14877);
nor U16340 (N_16340,N_14620,N_13627);
nor U16341 (N_16341,N_14915,N_13708);
nor U16342 (N_16342,N_14566,N_13991);
and U16343 (N_16343,N_13845,N_13907);
nor U16344 (N_16344,N_14570,N_14794);
nand U16345 (N_16345,N_13840,N_14368);
xor U16346 (N_16346,N_14319,N_14023);
or U16347 (N_16347,N_14348,N_14590);
xnor U16348 (N_16348,N_14328,N_14007);
xor U16349 (N_16349,N_14446,N_14295);
nand U16350 (N_16350,N_13714,N_13926);
nor U16351 (N_16351,N_14742,N_13702);
nand U16352 (N_16352,N_14115,N_14293);
nand U16353 (N_16353,N_14338,N_14989);
nor U16354 (N_16354,N_13926,N_13917);
or U16355 (N_16355,N_14673,N_13771);
nand U16356 (N_16356,N_14996,N_14900);
nor U16357 (N_16357,N_14068,N_13959);
or U16358 (N_16358,N_14311,N_14569);
and U16359 (N_16359,N_14014,N_14573);
nand U16360 (N_16360,N_14544,N_13586);
xor U16361 (N_16361,N_14085,N_14889);
nor U16362 (N_16362,N_14287,N_14519);
xor U16363 (N_16363,N_14197,N_14723);
and U16364 (N_16364,N_14658,N_14698);
or U16365 (N_16365,N_14016,N_14526);
nand U16366 (N_16366,N_14324,N_14874);
and U16367 (N_16367,N_14326,N_14751);
and U16368 (N_16368,N_14797,N_14682);
and U16369 (N_16369,N_14959,N_13514);
or U16370 (N_16370,N_13575,N_14084);
nand U16371 (N_16371,N_14574,N_14392);
or U16372 (N_16372,N_14443,N_13713);
or U16373 (N_16373,N_13900,N_14806);
nor U16374 (N_16374,N_14831,N_14465);
nor U16375 (N_16375,N_14348,N_13866);
and U16376 (N_16376,N_14977,N_14444);
or U16377 (N_16377,N_13564,N_14203);
xor U16378 (N_16378,N_13827,N_14080);
xnor U16379 (N_16379,N_14017,N_14565);
nor U16380 (N_16380,N_14934,N_14096);
xnor U16381 (N_16381,N_14897,N_14953);
nand U16382 (N_16382,N_13896,N_14807);
or U16383 (N_16383,N_14834,N_14447);
or U16384 (N_16384,N_14618,N_14521);
nor U16385 (N_16385,N_14334,N_14615);
or U16386 (N_16386,N_14664,N_13986);
and U16387 (N_16387,N_14831,N_14705);
or U16388 (N_16388,N_13892,N_14747);
nand U16389 (N_16389,N_14366,N_13931);
nor U16390 (N_16390,N_14648,N_14173);
nor U16391 (N_16391,N_14539,N_13688);
xor U16392 (N_16392,N_14448,N_14935);
or U16393 (N_16393,N_13866,N_14537);
nor U16394 (N_16394,N_14231,N_14957);
nor U16395 (N_16395,N_14009,N_13692);
nor U16396 (N_16396,N_14819,N_14010);
or U16397 (N_16397,N_13635,N_14546);
xnor U16398 (N_16398,N_13773,N_14214);
nor U16399 (N_16399,N_13815,N_14591);
and U16400 (N_16400,N_14952,N_14880);
nand U16401 (N_16401,N_14683,N_14749);
and U16402 (N_16402,N_14488,N_13671);
xnor U16403 (N_16403,N_13878,N_14768);
nand U16404 (N_16404,N_13626,N_14351);
xnor U16405 (N_16405,N_14069,N_14457);
or U16406 (N_16406,N_14445,N_13985);
nor U16407 (N_16407,N_14903,N_14111);
and U16408 (N_16408,N_13834,N_14050);
and U16409 (N_16409,N_13569,N_14683);
and U16410 (N_16410,N_14134,N_14816);
nand U16411 (N_16411,N_14480,N_13681);
nand U16412 (N_16412,N_13567,N_13820);
or U16413 (N_16413,N_13838,N_13887);
xnor U16414 (N_16414,N_14361,N_14896);
nor U16415 (N_16415,N_13540,N_14337);
nand U16416 (N_16416,N_14578,N_14337);
nor U16417 (N_16417,N_14121,N_13734);
xnor U16418 (N_16418,N_13573,N_14372);
or U16419 (N_16419,N_14797,N_13589);
nor U16420 (N_16420,N_14118,N_13823);
nand U16421 (N_16421,N_14909,N_14360);
xnor U16422 (N_16422,N_13505,N_14341);
nand U16423 (N_16423,N_13605,N_14187);
nand U16424 (N_16424,N_13722,N_14026);
nand U16425 (N_16425,N_14981,N_13968);
xnor U16426 (N_16426,N_14014,N_14851);
nor U16427 (N_16427,N_13520,N_14301);
nor U16428 (N_16428,N_14914,N_14919);
and U16429 (N_16429,N_14317,N_13939);
nor U16430 (N_16430,N_13905,N_14538);
or U16431 (N_16431,N_14666,N_14617);
nor U16432 (N_16432,N_14424,N_14019);
xnor U16433 (N_16433,N_14867,N_14054);
nor U16434 (N_16434,N_14512,N_14489);
nand U16435 (N_16435,N_14924,N_14964);
and U16436 (N_16436,N_13854,N_14668);
and U16437 (N_16437,N_14695,N_13552);
nor U16438 (N_16438,N_14561,N_13752);
nor U16439 (N_16439,N_14409,N_13831);
or U16440 (N_16440,N_14299,N_14538);
or U16441 (N_16441,N_14734,N_14247);
and U16442 (N_16442,N_14315,N_14549);
and U16443 (N_16443,N_13917,N_14003);
xnor U16444 (N_16444,N_13830,N_14121);
nor U16445 (N_16445,N_13860,N_13785);
xor U16446 (N_16446,N_13890,N_14872);
xnor U16447 (N_16447,N_14818,N_14207);
nand U16448 (N_16448,N_13826,N_13847);
xnor U16449 (N_16449,N_14777,N_13868);
nand U16450 (N_16450,N_14059,N_14044);
or U16451 (N_16451,N_14925,N_13920);
and U16452 (N_16452,N_13763,N_14315);
nand U16453 (N_16453,N_14914,N_14524);
nand U16454 (N_16454,N_14756,N_14388);
nor U16455 (N_16455,N_14400,N_14854);
nor U16456 (N_16456,N_13954,N_14368);
nand U16457 (N_16457,N_14151,N_14540);
nor U16458 (N_16458,N_14190,N_14854);
nand U16459 (N_16459,N_14976,N_14204);
and U16460 (N_16460,N_14947,N_14130);
and U16461 (N_16461,N_13786,N_13753);
nor U16462 (N_16462,N_14277,N_13905);
and U16463 (N_16463,N_14553,N_13568);
or U16464 (N_16464,N_13842,N_14416);
and U16465 (N_16465,N_14402,N_13860);
nor U16466 (N_16466,N_13698,N_14475);
nand U16467 (N_16467,N_14677,N_13513);
and U16468 (N_16468,N_14321,N_14835);
and U16469 (N_16469,N_14482,N_14774);
xor U16470 (N_16470,N_14045,N_14150);
or U16471 (N_16471,N_14078,N_14374);
nor U16472 (N_16472,N_14035,N_14718);
or U16473 (N_16473,N_14665,N_13641);
nand U16474 (N_16474,N_14892,N_14077);
and U16475 (N_16475,N_14331,N_14561);
nand U16476 (N_16476,N_14214,N_14561);
xnor U16477 (N_16477,N_13882,N_14297);
nor U16478 (N_16478,N_14733,N_14855);
nor U16479 (N_16479,N_14596,N_13657);
nor U16480 (N_16480,N_14429,N_14216);
nor U16481 (N_16481,N_14324,N_14177);
or U16482 (N_16482,N_14569,N_13828);
nor U16483 (N_16483,N_14429,N_14696);
xnor U16484 (N_16484,N_13995,N_14022);
nor U16485 (N_16485,N_14167,N_14143);
and U16486 (N_16486,N_14432,N_13735);
xor U16487 (N_16487,N_14773,N_14317);
nor U16488 (N_16488,N_14118,N_14823);
and U16489 (N_16489,N_13736,N_13528);
nand U16490 (N_16490,N_13804,N_14126);
nand U16491 (N_16491,N_14772,N_14479);
nor U16492 (N_16492,N_14202,N_13579);
nor U16493 (N_16493,N_14669,N_14314);
nand U16494 (N_16494,N_14388,N_13502);
xnor U16495 (N_16495,N_13698,N_14605);
nor U16496 (N_16496,N_14313,N_14183);
and U16497 (N_16497,N_14280,N_14394);
or U16498 (N_16498,N_14640,N_13644);
and U16499 (N_16499,N_13759,N_14253);
and U16500 (N_16500,N_15280,N_15987);
nor U16501 (N_16501,N_15402,N_15538);
xnor U16502 (N_16502,N_15419,N_15758);
or U16503 (N_16503,N_16122,N_15965);
nand U16504 (N_16504,N_15515,N_16482);
or U16505 (N_16505,N_15783,N_15213);
nor U16506 (N_16506,N_16466,N_15474);
nor U16507 (N_16507,N_15393,N_15675);
nor U16508 (N_16508,N_16095,N_16474);
and U16509 (N_16509,N_15053,N_16158);
and U16510 (N_16510,N_15547,N_16413);
or U16511 (N_16511,N_15268,N_15722);
and U16512 (N_16512,N_15631,N_15360);
nor U16513 (N_16513,N_15793,N_16327);
nand U16514 (N_16514,N_15037,N_15096);
nand U16515 (N_16515,N_15840,N_16308);
xnor U16516 (N_16516,N_15841,N_16355);
xor U16517 (N_16517,N_16395,N_16056);
nand U16518 (N_16518,N_15488,N_16354);
xor U16519 (N_16519,N_15262,N_16415);
or U16520 (N_16520,N_16377,N_15570);
nor U16521 (N_16521,N_15794,N_15322);
nor U16522 (N_16522,N_15774,N_16034);
and U16523 (N_16523,N_16256,N_15584);
and U16524 (N_16524,N_15316,N_15971);
xor U16525 (N_16525,N_15171,N_16182);
nor U16526 (N_16526,N_16003,N_15715);
nand U16527 (N_16527,N_15561,N_15478);
or U16528 (N_16528,N_15623,N_16352);
xor U16529 (N_16529,N_15852,N_15111);
and U16530 (N_16530,N_15896,N_16257);
or U16531 (N_16531,N_16362,N_16279);
or U16532 (N_16532,N_16453,N_16385);
or U16533 (N_16533,N_15523,N_15109);
or U16534 (N_16534,N_15389,N_15004);
or U16535 (N_16535,N_15269,N_15255);
and U16536 (N_16536,N_16037,N_15452);
or U16537 (N_16537,N_16269,N_16349);
xor U16538 (N_16538,N_16304,N_16188);
and U16539 (N_16539,N_16128,N_15778);
nor U16540 (N_16540,N_15988,N_16219);
nand U16541 (N_16541,N_15865,N_16195);
xor U16542 (N_16542,N_15916,N_15676);
xnor U16543 (N_16543,N_15796,N_16132);
and U16544 (N_16544,N_15301,N_15497);
or U16545 (N_16545,N_15242,N_15507);
or U16546 (N_16546,N_15953,N_15713);
nand U16547 (N_16547,N_16490,N_15358);
or U16548 (N_16548,N_15141,N_15076);
or U16549 (N_16549,N_15554,N_15510);
or U16550 (N_16550,N_15942,N_15278);
xnor U16551 (N_16551,N_15704,N_15336);
xnor U16552 (N_16552,N_15825,N_16163);
nand U16553 (N_16553,N_15996,N_15617);
or U16554 (N_16554,N_15308,N_16108);
and U16555 (N_16555,N_15589,N_15528);
or U16556 (N_16556,N_16222,N_16303);
xor U16557 (N_16557,N_15776,N_15600);
and U16558 (N_16558,N_15976,N_16330);
and U16559 (N_16559,N_16043,N_16042);
and U16560 (N_16560,N_16307,N_15388);
nor U16561 (N_16561,N_16293,N_15991);
and U16562 (N_16562,N_15525,N_15822);
or U16563 (N_16563,N_16210,N_15792);
nand U16564 (N_16564,N_15412,N_15010);
or U16565 (N_16565,N_15692,N_16129);
xor U16566 (N_16566,N_15798,N_15065);
nor U16567 (N_16567,N_16457,N_15231);
or U16568 (N_16568,N_15190,N_15216);
nor U16569 (N_16569,N_15626,N_16161);
or U16570 (N_16570,N_15870,N_15868);
xnor U16571 (N_16571,N_15445,N_15152);
nor U16572 (N_16572,N_16126,N_16053);
nand U16573 (N_16573,N_15031,N_16287);
nor U16574 (N_16574,N_15156,N_15804);
xor U16575 (N_16575,N_16370,N_15366);
or U16576 (N_16576,N_15657,N_16118);
xnor U16577 (N_16577,N_15457,N_15521);
or U16578 (N_16578,N_15112,N_15874);
xnor U16579 (N_16579,N_15305,N_15357);
nor U16580 (N_16580,N_15790,N_15009);
or U16581 (N_16581,N_16486,N_15335);
or U16582 (N_16582,N_15274,N_15451);
or U16583 (N_16583,N_16029,N_15977);
nor U16584 (N_16584,N_15502,N_15392);
xnor U16585 (N_16585,N_15831,N_16146);
nand U16586 (N_16586,N_16166,N_15655);
or U16587 (N_16587,N_15588,N_16398);
or U16588 (N_16588,N_15844,N_15967);
xor U16589 (N_16589,N_15479,N_15342);
or U16590 (N_16590,N_16365,N_16405);
nor U16591 (N_16591,N_16013,N_15081);
or U16592 (N_16592,N_16489,N_15481);
and U16593 (N_16593,N_16239,N_15805);
and U16594 (N_16594,N_15982,N_15134);
nand U16595 (N_16595,N_15292,N_16215);
xnor U16596 (N_16596,N_15957,N_15072);
or U16597 (N_16597,N_15661,N_16244);
nand U16598 (N_16598,N_15984,N_15816);
and U16599 (N_16599,N_16181,N_15299);
xor U16600 (N_16600,N_15233,N_15090);
or U16601 (N_16601,N_15283,N_16283);
xor U16602 (N_16602,N_16456,N_16258);
nand U16603 (N_16603,N_16030,N_15291);
or U16604 (N_16604,N_15490,N_16473);
or U16605 (N_16605,N_16424,N_15765);
nand U16606 (N_16606,N_15534,N_16484);
nor U16607 (N_16607,N_16455,N_15207);
and U16608 (N_16608,N_16315,N_16363);
nor U16609 (N_16609,N_15085,N_15245);
nor U16610 (N_16610,N_15239,N_15593);
nor U16611 (N_16611,N_16433,N_15106);
nor U16612 (N_16612,N_15116,N_15780);
and U16613 (N_16613,N_15416,N_15174);
xor U16614 (N_16614,N_16021,N_15801);
nor U16615 (N_16615,N_15887,N_16380);
and U16616 (N_16616,N_15968,N_15352);
and U16617 (N_16617,N_15341,N_15585);
nand U16618 (N_16618,N_16394,N_15082);
or U16619 (N_16619,N_15220,N_15737);
nand U16620 (N_16620,N_16452,N_16232);
xnor U16621 (N_16621,N_16241,N_15756);
xor U16622 (N_16622,N_15649,N_15959);
or U16623 (N_16623,N_16092,N_15423);
xor U16624 (N_16624,N_15215,N_15635);
and U16625 (N_16625,N_15634,N_15465);
nor U16626 (N_16626,N_15610,N_15048);
nor U16627 (N_16627,N_16091,N_16383);
nand U16628 (N_16628,N_15140,N_16052);
xor U16629 (N_16629,N_15818,N_15186);
nand U16630 (N_16630,N_15598,N_15855);
or U16631 (N_16631,N_15315,N_15817);
xnor U16632 (N_16632,N_15340,N_15736);
nor U16633 (N_16633,N_15154,N_15422);
xnor U16634 (N_16634,N_15093,N_16059);
nor U16635 (N_16635,N_15560,N_15836);
nor U16636 (N_16636,N_16321,N_15579);
nand U16637 (N_16637,N_16094,N_15363);
nand U16638 (N_16638,N_15732,N_15568);
xor U16639 (N_16639,N_15621,N_15222);
nand U16640 (N_16640,N_15952,N_15636);
xor U16641 (N_16641,N_15943,N_15477);
nor U16642 (N_16642,N_16298,N_15503);
nor U16643 (N_16643,N_16062,N_15845);
and U16644 (N_16644,N_16493,N_15842);
nand U16645 (N_16645,N_16375,N_15998);
xor U16646 (N_16646,N_16389,N_16427);
nand U16647 (N_16647,N_15074,N_15472);
nand U16648 (N_16648,N_15034,N_15056);
and U16649 (N_16649,N_16367,N_15068);
or U16650 (N_16650,N_15908,N_15620);
xnor U16651 (N_16651,N_15361,N_15903);
nand U16652 (N_16652,N_16294,N_15189);
or U16653 (N_16653,N_15411,N_16218);
nor U16654 (N_16654,N_16155,N_15716);
or U16655 (N_16655,N_16001,N_16420);
or U16656 (N_16656,N_15611,N_15974);
xor U16657 (N_16657,N_16265,N_15501);
xor U16658 (N_16658,N_15639,N_16458);
xnor U16659 (N_16659,N_16206,N_16150);
nand U16660 (N_16660,N_15045,N_15420);
nand U16661 (N_16661,N_16446,N_15992);
xnor U16662 (N_16662,N_15710,N_15766);
or U16663 (N_16663,N_15754,N_15223);
or U16664 (N_16664,N_16376,N_15829);
or U16665 (N_16665,N_15670,N_15548);
xnor U16666 (N_16666,N_15044,N_16419);
and U16667 (N_16667,N_16381,N_15489);
nand U16668 (N_16668,N_15442,N_16116);
xor U16669 (N_16669,N_15915,N_15520);
or U16670 (N_16670,N_15929,N_16319);
nor U16671 (N_16671,N_16470,N_16339);
and U16672 (N_16672,N_15815,N_15229);
nor U16673 (N_16673,N_16190,N_15695);
nor U16674 (N_16674,N_15181,N_15252);
and U16675 (N_16675,N_15294,N_16176);
nor U16676 (N_16676,N_15443,N_15764);
nor U16677 (N_16677,N_15257,N_15247);
nand U16678 (N_16678,N_16019,N_15356);
or U16679 (N_16679,N_15421,N_15517);
nor U16680 (N_16680,N_15260,N_15613);
nor U16681 (N_16681,N_15089,N_16164);
nor U16682 (N_16682,N_15033,N_15787);
or U16683 (N_16683,N_16491,N_16160);
nand U16684 (N_16684,N_15949,N_15185);
and U16685 (N_16685,N_15011,N_15003);
or U16686 (N_16686,N_16317,N_16282);
and U16687 (N_16687,N_15328,N_15265);
or U16688 (N_16688,N_16261,N_16478);
nor U16689 (N_16689,N_16302,N_15179);
and U16690 (N_16690,N_15772,N_16110);
or U16691 (N_16691,N_15781,N_15024);
nor U16692 (N_16692,N_15399,N_15729);
and U16693 (N_16693,N_16499,N_16088);
nor U16694 (N_16694,N_15436,N_15266);
xnor U16695 (N_16695,N_16007,N_16387);
or U16696 (N_16696,N_15348,N_15990);
nand U16697 (N_16697,N_15406,N_16255);
and U16698 (N_16698,N_16253,N_16310);
and U16699 (N_16699,N_15893,N_15103);
xor U16700 (N_16700,N_16072,N_16236);
or U16701 (N_16701,N_16173,N_15954);
nand U16702 (N_16702,N_15924,N_15046);
or U16703 (N_16703,N_15043,N_16425);
xor U16704 (N_16704,N_16076,N_16213);
and U16705 (N_16705,N_15197,N_16178);
nor U16706 (N_16706,N_15867,N_16494);
nand U16707 (N_16707,N_15051,N_15161);
nor U16708 (N_16708,N_15227,N_15725);
and U16709 (N_16709,N_16399,N_15755);
nor U16710 (N_16710,N_16038,N_15178);
xnor U16711 (N_16711,N_15110,N_16322);
or U16712 (N_16712,N_16048,N_16372);
or U16713 (N_16713,N_16171,N_15079);
nand U16714 (N_16714,N_16207,N_15448);
xor U16715 (N_16715,N_15157,N_16216);
and U16716 (N_16716,N_15484,N_15809);
and U16717 (N_16717,N_15938,N_15234);
nand U16718 (N_16718,N_15290,N_16196);
and U16719 (N_16719,N_15808,N_16475);
nand U16720 (N_16720,N_15877,N_15312);
xor U16721 (N_16721,N_15856,N_16252);
and U16722 (N_16722,N_15459,N_15373);
xnor U16723 (N_16723,N_15075,N_15061);
nor U16724 (N_16724,N_16378,N_15370);
and U16725 (N_16725,N_16454,N_16270);
xnor U16726 (N_16726,N_15683,N_15823);
xor U16727 (N_16727,N_16344,N_15820);
nand U16728 (N_16728,N_15961,N_16331);
and U16729 (N_16729,N_15450,N_15824);
nor U16730 (N_16730,N_16249,N_15062);
nand U16731 (N_16731,N_15426,N_15678);
or U16732 (N_16732,N_15115,N_15662);
xor U16733 (N_16733,N_15562,N_15875);
nor U16734 (N_16734,N_15017,N_15797);
or U16735 (N_16735,N_15738,N_16318);
or U16736 (N_16736,N_15496,N_16417);
or U16737 (N_16737,N_15993,N_16423);
or U16738 (N_16738,N_15254,N_15644);
or U16739 (N_16739,N_15843,N_16066);
and U16740 (N_16740,N_16393,N_15331);
or U16741 (N_16741,N_15762,N_15939);
or U16742 (N_16742,N_15691,N_16267);
or U16743 (N_16743,N_15830,N_15201);
or U16744 (N_16744,N_16471,N_15441);
nor U16745 (N_16745,N_15002,N_15860);
nor U16746 (N_16746,N_16100,N_15120);
and U16747 (N_16747,N_15752,N_15819);
nor U16748 (N_16748,N_15904,N_15175);
nand U16749 (N_16749,N_16280,N_15005);
and U16750 (N_16750,N_15279,N_16329);
xor U16751 (N_16751,N_16430,N_16187);
xnor U16752 (N_16752,N_15935,N_16063);
nand U16753 (N_16753,N_15616,N_15694);
or U16754 (N_16754,N_16106,N_15468);
nor U16755 (N_16755,N_15139,N_16462);
nand U16756 (N_16756,N_15559,N_15381);
nand U16757 (N_16757,N_15343,N_16245);
nand U16758 (N_16758,N_15487,N_16185);
nor U16759 (N_16759,N_15912,N_15828);
or U16760 (N_16760,N_15482,N_15891);
and U16761 (N_16761,N_15964,N_16358);
nor U16762 (N_16762,N_16000,N_15609);
nor U16763 (N_16763,N_15872,N_16151);
nor U16764 (N_16764,N_15576,N_15320);
and U16765 (N_16765,N_15169,N_15122);
nor U16766 (N_16766,N_15162,N_16492);
nor U16767 (N_16767,N_15272,N_16481);
nor U16768 (N_16768,N_15235,N_16004);
nor U16769 (N_16769,N_15835,N_15862);
xor U16770 (N_16770,N_15741,N_16198);
or U16771 (N_16771,N_16193,N_15196);
and U16772 (N_16772,N_16334,N_16006);
and U16773 (N_16773,N_15092,N_15369);
xor U16774 (N_16774,N_15379,N_16112);
or U16775 (N_16775,N_16123,N_16297);
nand U16776 (N_16776,N_15970,N_15923);
xor U16777 (N_16777,N_15105,N_15401);
or U16778 (N_16778,N_16276,N_15608);
xnor U16779 (N_16779,N_15720,N_16011);
nor U16780 (N_16780,N_15919,N_15512);
nand U16781 (N_16781,N_15126,N_15123);
or U16782 (N_16782,N_16268,N_16311);
xnor U16783 (N_16783,N_16046,N_15753);
nand U16784 (N_16784,N_15647,N_15454);
nand U16785 (N_16785,N_15067,N_15132);
xnor U16786 (N_16786,N_15446,N_16231);
xnor U16787 (N_16787,N_16031,N_15777);
and U16788 (N_16788,N_15371,N_16374);
nor U16789 (N_16789,N_15172,N_15858);
nor U16790 (N_16790,N_15637,N_16172);
and U16791 (N_16791,N_16469,N_15042);
nor U16792 (N_16792,N_16409,N_15837);
or U16793 (N_16793,N_16027,N_16058);
xor U16794 (N_16794,N_15095,N_16115);
nand U16795 (N_16795,N_15723,N_16071);
nor U16796 (N_16796,N_16049,N_15920);
xnor U16797 (N_16797,N_16104,N_15551);
nand U16798 (N_16798,N_15150,N_15296);
nand U16799 (N_16799,N_15565,N_16439);
nand U16800 (N_16800,N_15572,N_16266);
or U16801 (N_16801,N_15898,N_15873);
nand U16802 (N_16802,N_16217,N_16065);
and U16803 (N_16803,N_15311,N_16277);
xor U16804 (N_16804,N_15133,N_15368);
or U16805 (N_16805,N_15219,N_16356);
xor U16806 (N_16806,N_15098,N_15535);
xor U16807 (N_16807,N_16414,N_16403);
xor U16808 (N_16808,N_16246,N_15192);
nand U16809 (N_16809,N_15654,N_15211);
or U16810 (N_16810,N_16214,N_15099);
nand U16811 (N_16811,N_15881,N_15310);
xnor U16812 (N_16812,N_15078,N_16090);
and U16813 (N_16813,N_15376,N_16177);
nor U16814 (N_16814,N_15052,N_16229);
nand U16815 (N_16815,N_15149,N_15587);
and U16816 (N_16816,N_15183,N_16186);
or U16817 (N_16817,N_15909,N_15333);
or U16818 (N_16818,N_16488,N_16200);
or U16819 (N_16819,N_16361,N_15117);
nor U16820 (N_16820,N_15846,N_15289);
nand U16821 (N_16821,N_16098,N_16247);
xnor U16822 (N_16822,N_16295,N_15205);
xor U16823 (N_16823,N_16148,N_15251);
xnor U16824 (N_16824,N_15540,N_16026);
nand U16825 (N_16825,N_15253,N_15230);
or U16826 (N_16826,N_15086,N_16093);
or U16827 (N_16827,N_15345,N_16404);
or U16828 (N_16828,N_15417,N_15071);
nor U16829 (N_16829,N_15595,N_15667);
and U16830 (N_16830,N_15176,N_15771);
nor U16831 (N_16831,N_15407,N_15264);
xor U16832 (N_16832,N_16113,N_16301);
and U16833 (N_16833,N_16041,N_15890);
or U16834 (N_16834,N_15833,N_15131);
xor U16835 (N_16835,N_16199,N_15894);
nor U16836 (N_16836,N_15983,N_15799);
xor U16837 (N_16837,N_15769,N_16460);
nand U16838 (N_16838,N_15545,N_15466);
and U16839 (N_16839,N_15641,N_15885);
nor U16840 (N_16840,N_15386,N_16335);
or U16841 (N_16841,N_15979,N_15058);
xnor U16842 (N_16842,N_16134,N_15327);
nand U16843 (N_16843,N_15057,N_15329);
nor U16844 (N_16844,N_15925,N_15461);
nand U16845 (N_16845,N_16400,N_15326);
or U16846 (N_16846,N_16169,N_15748);
or U16847 (N_16847,N_15966,N_15138);
nand U16848 (N_16848,N_15458,N_15800);
and U16849 (N_16849,N_15849,N_15403);
nor U16850 (N_16850,N_16125,N_15351);
xor U16851 (N_16851,N_15372,N_15530);
nand U16852 (N_16852,N_15986,N_15226);
nand U16853 (N_16853,N_15951,N_16451);
nor U16854 (N_16854,N_15055,N_15094);
nand U16855 (N_16855,N_16240,N_15854);
and U16856 (N_16856,N_16416,N_15113);
and U16857 (N_16857,N_15643,N_15492);
nand U16858 (N_16858,N_15447,N_16472);
nand U16859 (N_16859,N_15449,N_16057);
nor U16860 (N_16860,N_15549,N_15869);
xor U16861 (N_16861,N_16289,N_15532);
or U16862 (N_16862,N_15006,N_15020);
xnor U16863 (N_16863,N_15785,N_15267);
nor U16864 (N_16864,N_16422,N_15439);
and U16865 (N_16865,N_16203,N_15581);
xnor U16866 (N_16866,N_16141,N_15153);
nor U16867 (N_16867,N_16067,N_15362);
xnor U16868 (N_16868,N_16159,N_15374);
and U16869 (N_16869,N_16073,N_15632);
xor U16870 (N_16870,N_15270,N_15127);
nand U16871 (N_16871,N_15603,N_16202);
or U16872 (N_16872,N_16306,N_15910);
or U16873 (N_16873,N_15339,N_16396);
nand U16874 (N_16874,N_15851,N_15184);
and U16875 (N_16875,N_16061,N_16124);
nor U16876 (N_16876,N_15546,N_16221);
and U16877 (N_16877,N_15651,N_16174);
or U16878 (N_16878,N_16254,N_16023);
or U16879 (N_16879,N_16450,N_16012);
or U16880 (N_16880,N_15658,N_15557);
or U16881 (N_16881,N_15526,N_15430);
and U16882 (N_16882,N_16291,N_15202);
or U16883 (N_16883,N_16175,N_15250);
or U16884 (N_16884,N_16170,N_15224);
xnor U16885 (N_16885,N_15317,N_16443);
nor U16886 (N_16886,N_15097,N_15170);
xnor U16887 (N_16887,N_15582,N_16426);
nand U16888 (N_16888,N_15701,N_16228);
and U16889 (N_16889,N_15509,N_15499);
and U16890 (N_16890,N_15880,N_16167);
nor U16891 (N_16891,N_15435,N_15905);
and U16892 (N_16892,N_15811,N_15876);
xnor U16893 (N_16893,N_15259,N_16184);
or U16894 (N_16894,N_15615,N_16341);
xnor U16895 (N_16895,N_16099,N_16153);
nor U16896 (N_16896,N_15604,N_15306);
xor U16897 (N_16897,N_15273,N_16305);
xnor U16898 (N_16898,N_15871,N_15015);
nand U16899 (N_16899,N_15030,N_15129);
nor U16900 (N_16900,N_15607,N_15091);
xnor U16901 (N_16901,N_15049,N_16431);
xnor U16902 (N_16902,N_15209,N_15404);
or U16903 (N_16903,N_15945,N_16064);
nand U16904 (N_16904,N_15646,N_15237);
and U16905 (N_16905,N_15980,N_15533);
xor U16906 (N_16906,N_15028,N_15907);
nand U16907 (N_16907,N_15995,N_15410);
xnor U16908 (N_16908,N_15775,N_16069);
xor U16909 (N_16909,N_16320,N_16314);
nor U16910 (N_16910,N_15969,N_15806);
xor U16911 (N_16911,N_15377,N_15200);
xnor U16912 (N_16912,N_15246,N_16441);
nor U16913 (N_16913,N_15628,N_15505);
nand U16914 (N_16914,N_16410,N_16024);
xnor U16915 (N_16915,N_15365,N_15295);
and U16916 (N_16916,N_15147,N_16495);
or U16917 (N_16917,N_15630,N_16237);
or U16918 (N_16918,N_16131,N_15070);
and U16919 (N_16919,N_15035,N_16434);
nor U16920 (N_16920,N_15325,N_15288);
nand U16921 (N_16921,N_16018,N_16262);
and U16922 (N_16922,N_15000,N_16197);
xor U16923 (N_16923,N_16101,N_16044);
nand U16924 (N_16924,N_15397,N_16144);
or U16925 (N_16925,N_15897,N_15687);
xnor U16926 (N_16926,N_15689,N_16045);
nand U16927 (N_16927,N_15191,N_15244);
and U16928 (N_16928,N_16086,N_16114);
nand U16929 (N_16929,N_15455,N_16233);
or U16930 (N_16930,N_15590,N_15396);
and U16931 (N_16931,N_16299,N_15763);
and U16932 (N_16932,N_15936,N_16224);
or U16933 (N_16933,N_15390,N_16447);
nor U16934 (N_16934,N_16209,N_15847);
xnor U16935 (N_16935,N_15696,N_16480);
and U16936 (N_16936,N_15434,N_15718);
and U16937 (N_16937,N_16017,N_15866);
nand U16938 (N_16938,N_16464,N_15937);
xnor U16939 (N_16939,N_15958,N_15650);
nand U16940 (N_16940,N_15779,N_15008);
xnor U16941 (N_16941,N_15879,N_16010);
nand U16942 (N_16942,N_15918,N_16168);
and U16943 (N_16943,N_16127,N_16278);
and U16944 (N_16944,N_15409,N_15944);
xnor U16945 (N_16945,N_16082,N_15210);
xnor U16946 (N_16946,N_15962,N_15975);
nand U16947 (N_16947,N_15271,N_16438);
and U16948 (N_16948,N_15791,N_16050);
xor U16949 (N_16949,N_16234,N_16497);
nor U16950 (N_16950,N_15606,N_16357);
or U16951 (N_16951,N_15660,N_16436);
nand U16952 (N_16952,N_15493,N_15387);
nor U16953 (N_16953,N_15414,N_15727);
xor U16954 (N_16954,N_15314,N_16461);
xor U16955 (N_16955,N_15124,N_15697);
nand U16956 (N_16956,N_15928,N_16364);
and U16957 (N_16957,N_15524,N_15803);
xnor U16958 (N_16958,N_15656,N_15432);
and U16959 (N_16959,N_15674,N_15575);
and U16960 (N_16960,N_16103,N_15088);
nor U16961 (N_16961,N_15145,N_16102);
and U16962 (N_16962,N_16015,N_15168);
and U16963 (N_16963,N_16467,N_15384);
nor U16964 (N_16964,N_16075,N_16487);
and U16965 (N_16965,N_15734,N_15114);
xnor U16966 (N_16966,N_15164,N_15659);
nor U16967 (N_16967,N_16350,N_15025);
nand U16968 (N_16968,N_16008,N_15059);
xor U16969 (N_16969,N_15119,N_16392);
xor U16970 (N_16970,N_15597,N_15542);
and U16971 (N_16971,N_15956,N_15321);
or U16972 (N_16972,N_16351,N_16296);
nor U16973 (N_16973,N_15155,N_16496);
xor U16974 (N_16974,N_16273,N_15475);
xnor U16975 (N_16975,N_16323,N_15125);
or U16976 (N_16976,N_15394,N_15940);
nand U16977 (N_16977,N_15243,N_15293);
or U16978 (N_16978,N_15188,N_15750);
or U16979 (N_16979,N_15889,N_16083);
nand U16980 (N_16980,N_16235,N_15281);
and U16981 (N_16981,N_15437,N_16035);
and U16982 (N_16982,N_15398,N_16368);
xnor U16983 (N_16983,N_15553,N_16371);
nand U16984 (N_16984,N_16040,N_15130);
and U16985 (N_16985,N_16373,N_15784);
nand U16986 (N_16986,N_15144,N_15552);
or U16987 (N_16987,N_16407,N_15495);
or U16988 (N_16988,N_16477,N_15693);
nand U16989 (N_16989,N_15955,N_16133);
nand U16990 (N_16990,N_16336,N_15413);
and U16991 (N_16991,N_16390,N_15782);
or U16992 (N_16992,N_16191,N_16442);
or U16993 (N_16993,N_16402,N_15927);
xor U16994 (N_16994,N_15848,N_15298);
nand U16995 (N_16995,N_16147,N_16440);
nand U16996 (N_16996,N_15878,N_15680);
and U16997 (N_16997,N_16194,N_15541);
xnor U16998 (N_16998,N_16353,N_15225);
or U16999 (N_16999,N_15640,N_15400);
nand U17000 (N_17000,N_15100,N_15917);
or U17001 (N_17001,N_15583,N_15313);
nor U17002 (N_17002,N_16087,N_15684);
nand U17003 (N_17003,N_16020,N_15702);
nand U17004 (N_17004,N_16028,N_15456);
and U17005 (N_17005,N_16136,N_15084);
and U17006 (N_17006,N_16211,N_15544);
xor U17007 (N_17007,N_15978,N_16259);
nor U17008 (N_17008,N_15364,N_16078);
xor U17009 (N_17009,N_16290,N_15663);
nand U17010 (N_17010,N_16397,N_15946);
and U17011 (N_17011,N_15911,N_15564);
nand U17012 (N_17012,N_16333,N_16281);
xor U17013 (N_17013,N_15483,N_15749);
xnor U17014 (N_17014,N_15947,N_15187);
nor U17015 (N_17015,N_15217,N_15733);
xnor U17016 (N_17016,N_15415,N_15338);
or U17017 (N_17017,N_15906,N_15240);
or U17018 (N_17018,N_15516,N_16060);
or U17019 (N_17019,N_15726,N_15931);
and U17020 (N_17020,N_15228,N_15638);
nand U17021 (N_17021,N_15864,N_15653);
or U17022 (N_17022,N_16347,N_15433);
nor U17023 (N_17023,N_15853,N_16033);
nor U17024 (N_17024,N_15768,N_15605);
and U17025 (N_17025,N_15204,N_16251);
xnor U17026 (N_17026,N_15166,N_15721);
xor U17027 (N_17027,N_16444,N_16412);
xnor U17028 (N_17028,N_16312,N_15813);
xnor U17029 (N_17029,N_16437,N_15063);
or U17030 (N_17030,N_16346,N_16432);
xor U17031 (N_17031,N_15504,N_15232);
or U17032 (N_17032,N_16248,N_15083);
and U17033 (N_17033,N_15485,N_15950);
xnor U17034 (N_17034,N_15263,N_16272);
or U17035 (N_17035,N_16435,N_16348);
and U17036 (N_17036,N_15193,N_15705);
or U17037 (N_17037,N_15380,N_15677);
or U17038 (N_17038,N_16369,N_16483);
nand U17039 (N_17039,N_15627,N_16300);
nand U17040 (N_17040,N_16382,N_15742);
or U17041 (N_17041,N_15814,N_16005);
or U17042 (N_17042,N_15926,N_15933);
and U17043 (N_17043,N_16250,N_15892);
or U17044 (N_17044,N_15453,N_16032);
xor U17045 (N_17045,N_16145,N_15556);
nor U17046 (N_17046,N_15309,N_15108);
nand U17047 (N_17047,N_15050,N_16192);
nand U17048 (N_17048,N_15241,N_15601);
or U17049 (N_17049,N_16337,N_15645);
nor U17050 (N_17050,N_15344,N_15355);
and U17051 (N_17051,N_15594,N_15307);
nor U17052 (N_17052,N_15165,N_15480);
and U17053 (N_17053,N_16016,N_15258);
nor U17054 (N_17054,N_15751,N_15728);
or U17055 (N_17055,N_15886,N_16201);
and U17056 (N_17056,N_15102,N_15519);
xnor U17057 (N_17057,N_15500,N_16068);
or U17058 (N_17058,N_15591,N_16079);
and U17059 (N_17059,N_15625,N_16119);
xor U17060 (N_17060,N_16014,N_15444);
xnor U17061 (N_17061,N_15973,N_15711);
nor U17062 (N_17062,N_16225,N_15863);
nand U17063 (N_17063,N_16022,N_15767);
or U17064 (N_17064,N_15679,N_16220);
xnor U17065 (N_17065,N_16485,N_16097);
nand U17066 (N_17066,N_15724,N_15332);
nand U17067 (N_17067,N_15027,N_15463);
and U17068 (N_17068,N_15900,N_15438);
nor U17069 (N_17069,N_15137,N_15285);
nor U17070 (N_17070,N_15198,N_15167);
and U17071 (N_17071,N_16468,N_16162);
nand U17072 (N_17072,N_15440,N_15699);
nor U17073 (N_17073,N_15014,N_15163);
or U17074 (N_17074,N_15429,N_16386);
nand U17075 (N_17075,N_15087,N_16313);
and U17076 (N_17076,N_15537,N_15812);
nor U17077 (N_17077,N_15238,N_15773);
nor U17078 (N_17078,N_15747,N_15743);
and U17079 (N_17079,N_15038,N_15602);
or U17080 (N_17080,N_16080,N_15731);
nor U17081 (N_17081,N_15574,N_15761);
nor U17082 (N_17082,N_15997,N_15236);
or U17083 (N_17083,N_16165,N_15032);
or U17084 (N_17084,N_15883,N_15060);
nor U17085 (N_17085,N_15019,N_15143);
or U17086 (N_17086,N_16343,N_15760);
xor U17087 (N_17087,N_15395,N_16379);
nand U17088 (N_17088,N_15382,N_16274);
nor U17089 (N_17089,N_15203,N_15558);
xor U17090 (N_17090,N_15029,N_15578);
or U17091 (N_17091,N_16316,N_15473);
nor U17092 (N_17092,N_15375,N_15688);
nand U17093 (N_17093,N_15476,N_15700);
and U17094 (N_17094,N_15902,N_16156);
xnor U17095 (N_17095,N_16286,N_15972);
or U17096 (N_17096,N_15899,N_15080);
xor U17097 (N_17097,N_15023,N_15346);
xnor U17098 (N_17098,N_15330,N_16384);
nand U17099 (N_17099,N_15941,N_15618);
nor U17100 (N_17100,N_16325,N_16292);
xnor U17101 (N_17101,N_15786,N_15681);
xor U17102 (N_17102,N_15664,N_16418);
nor U17103 (N_17103,N_15508,N_15026);
or U17104 (N_17104,N_16263,N_16138);
and U17105 (N_17105,N_16448,N_16328);
nand U17106 (N_17106,N_15464,N_16002);
nor U17107 (N_17107,N_16463,N_15334);
and U17108 (N_17108,N_15539,N_15648);
or U17109 (N_17109,N_15596,N_15666);
and U17110 (N_17110,N_15180,N_15104);
xnor U17111 (N_17111,N_15913,N_15832);
or U17112 (N_17112,N_15690,N_16077);
xnor U17113 (N_17113,N_16180,N_15555);
nand U17114 (N_17114,N_15018,N_16479);
nand U17115 (N_17115,N_15821,N_15022);
or U17116 (N_17116,N_15431,N_15286);
xor U17117 (N_17117,N_15531,N_15709);
or U17118 (N_17118,N_15857,N_15922);
and U17119 (N_17119,N_15016,N_15665);
xnor U17120 (N_17120,N_15624,N_16054);
and U17121 (N_17121,N_15599,N_15948);
xor U17122 (N_17122,N_15347,N_15550);
nor U17123 (N_17123,N_15571,N_15802);
or U17124 (N_17124,N_15177,N_15261);
xor U17125 (N_17125,N_15934,N_15303);
nand U17126 (N_17126,N_15712,N_15354);
or U17127 (N_17127,N_16036,N_15323);
or U17128 (N_17128,N_15218,N_15494);
xor U17129 (N_17129,N_15717,N_15248);
nand U17130 (N_17130,N_15302,N_16445);
nand U17131 (N_17131,N_15567,N_15619);
and U17132 (N_17132,N_16051,N_15981);
and U17133 (N_17133,N_15275,N_15622);
nor U17134 (N_17134,N_15160,N_15353);
xor U17135 (N_17135,N_16338,N_15807);
xor U17136 (N_17136,N_15746,N_16275);
xnor U17137 (N_17137,N_15039,N_15668);
xnor U17138 (N_17138,N_16047,N_15121);
and U17139 (N_17139,N_15673,N_16074);
xnor U17140 (N_17140,N_16183,N_16285);
or U17141 (N_17141,N_15319,N_16208);
nor U17142 (N_17142,N_16459,N_16340);
xnor U17143 (N_17143,N_15826,N_15740);
or U17144 (N_17144,N_15757,N_15040);
nor U17145 (N_17145,N_15629,N_16121);
nor U17146 (N_17146,N_15850,N_16189);
nor U17147 (N_17147,N_16271,N_15795);
nor U17148 (N_17148,N_15895,N_16391);
xnor U17149 (N_17149,N_15013,N_15349);
nand U17150 (N_17150,N_15427,N_15469);
nor U17151 (N_17151,N_15300,N_15708);
xnor U17152 (N_17152,N_16107,N_15514);
and U17153 (N_17153,N_16089,N_16264);
nor U17154 (N_17154,N_16309,N_15385);
nand U17155 (N_17155,N_16105,N_15707);
nand U17156 (N_17156,N_15810,N_16342);
and U17157 (N_17157,N_15212,N_15744);
nand U17158 (N_17158,N_15256,N_15580);
xnor U17159 (N_17159,N_15698,N_15543);
nor U17160 (N_17160,N_15101,N_16401);
xor U17161 (N_17161,N_15173,N_15367);
nor U17162 (N_17162,N_15424,N_15158);
or U17163 (N_17163,N_16084,N_15066);
xor U17164 (N_17164,N_15221,N_15827);
and U17165 (N_17165,N_16288,N_16332);
xnor U17166 (N_17166,N_16135,N_16142);
nand U17167 (N_17167,N_15989,N_15960);
and U17168 (N_17168,N_15682,N_15195);
or U17169 (N_17169,N_15383,N_16025);
or U17170 (N_17170,N_15378,N_16154);
xnor U17171 (N_17171,N_16085,N_16421);
or U17172 (N_17172,N_15730,N_15569);
xnor U17173 (N_17173,N_15001,N_15930);
nor U17174 (N_17174,N_15888,N_15007);
nor U17175 (N_17175,N_15839,N_15428);
and U17176 (N_17176,N_15706,N_16429);
xor U17177 (N_17177,N_16360,N_16428);
and U17178 (N_17178,N_15284,N_15884);
xnor U17179 (N_17179,N_15739,N_15182);
nand U17180 (N_17180,N_15276,N_16039);
nand U17181 (N_17181,N_15199,N_15498);
or U17182 (N_17182,N_15491,N_16204);
nor U17183 (N_17183,N_16284,N_16238);
nand U17184 (N_17184,N_15425,N_15214);
and U17185 (N_17185,N_15486,N_15159);
xor U17186 (N_17186,N_15021,N_16226);
nor U17187 (N_17187,N_15592,N_15054);
nand U17188 (N_17188,N_16243,N_15511);
nor U17189 (N_17189,N_15513,N_16366);
and U17190 (N_17190,N_15324,N_15206);
nor U17191 (N_17191,N_15012,N_16139);
or U17192 (N_17192,N_16406,N_15470);
or U17193 (N_17193,N_16326,N_15146);
or U17194 (N_17194,N_15685,N_15462);
and U17195 (N_17195,N_15041,N_15633);
and U17196 (N_17196,N_16179,N_15536);
xnor U17197 (N_17197,N_15135,N_15136);
xnor U17198 (N_17198,N_15882,N_15745);
xnor U17199 (N_17199,N_15148,N_15337);
xor U17200 (N_17200,N_15522,N_15999);
or U17201 (N_17201,N_15838,N_15566);
and U17202 (N_17202,N_15901,N_16223);
nor U17203 (N_17203,N_16408,N_16449);
nand U17204 (N_17204,N_15073,N_15249);
and U17205 (N_17205,N_15921,N_16212);
xnor U17206 (N_17206,N_16140,N_15142);
nor U17207 (N_17207,N_15277,N_15391);
nand U17208 (N_17208,N_15788,N_15297);
nor U17209 (N_17209,N_16096,N_15208);
or U17210 (N_17210,N_15506,N_16411);
or U17211 (N_17211,N_15151,N_15064);
and U17212 (N_17212,N_15467,N_15460);
xor U17213 (N_17213,N_15834,N_15118);
and U17214 (N_17214,N_15932,N_16070);
xnor U17215 (N_17215,N_15577,N_15350);
nor U17216 (N_17216,N_15719,N_15859);
nand U17217 (N_17217,N_15669,N_15471);
xor U17218 (N_17218,N_16498,N_16465);
and U17219 (N_17219,N_15642,N_15586);
xor U17220 (N_17220,N_15789,N_16230);
and U17221 (N_17221,N_15287,N_15671);
nor U17222 (N_17222,N_16055,N_16149);
nor U17223 (N_17223,N_15861,N_16227);
nor U17224 (N_17224,N_15304,N_16137);
xnor U17225 (N_17225,N_16345,N_15735);
xor U17226 (N_17226,N_15985,N_15405);
nand U17227 (N_17227,N_15282,N_16111);
nand U17228 (N_17228,N_15069,N_16130);
or U17229 (N_17229,N_15128,N_16205);
and U17230 (N_17230,N_15318,N_16324);
or U17231 (N_17231,N_15672,N_15612);
or U17232 (N_17232,N_15563,N_16109);
xor U17233 (N_17233,N_16117,N_16359);
or U17234 (N_17234,N_15914,N_15107);
or U17235 (N_17235,N_15714,N_15573);
nand U17236 (N_17236,N_15077,N_16242);
nand U17237 (N_17237,N_15770,N_15518);
xnor U17238 (N_17238,N_15686,N_16081);
or U17239 (N_17239,N_16143,N_16388);
nand U17240 (N_17240,N_15527,N_15652);
nor U17241 (N_17241,N_15994,N_15529);
and U17242 (N_17242,N_15963,N_16476);
xor U17243 (N_17243,N_15359,N_15614);
xnor U17244 (N_17244,N_16120,N_15703);
xnor U17245 (N_17245,N_16260,N_15036);
nand U17246 (N_17246,N_15047,N_15194);
nand U17247 (N_17247,N_16009,N_16152);
xor U17248 (N_17248,N_16157,N_15418);
and U17249 (N_17249,N_15408,N_15759);
nor U17250 (N_17250,N_16319,N_15903);
or U17251 (N_17251,N_15024,N_15983);
nand U17252 (N_17252,N_15289,N_16454);
or U17253 (N_17253,N_15025,N_15963);
nand U17254 (N_17254,N_16460,N_16275);
or U17255 (N_17255,N_15690,N_15315);
or U17256 (N_17256,N_16254,N_15399);
or U17257 (N_17257,N_15490,N_15686);
or U17258 (N_17258,N_15542,N_15909);
nand U17259 (N_17259,N_15446,N_15717);
nand U17260 (N_17260,N_16054,N_15467);
or U17261 (N_17261,N_15994,N_15280);
and U17262 (N_17262,N_15068,N_15921);
xor U17263 (N_17263,N_15959,N_15476);
or U17264 (N_17264,N_15749,N_15201);
xnor U17265 (N_17265,N_15735,N_16119);
nand U17266 (N_17266,N_16246,N_15990);
nand U17267 (N_17267,N_15799,N_15847);
xnor U17268 (N_17268,N_15305,N_15452);
and U17269 (N_17269,N_15494,N_15669);
and U17270 (N_17270,N_15670,N_15793);
nor U17271 (N_17271,N_15343,N_15716);
or U17272 (N_17272,N_15662,N_16253);
and U17273 (N_17273,N_15768,N_16279);
xor U17274 (N_17274,N_16431,N_15041);
or U17275 (N_17275,N_16431,N_15282);
nor U17276 (N_17276,N_15903,N_16265);
or U17277 (N_17277,N_15486,N_15568);
or U17278 (N_17278,N_15717,N_15898);
nor U17279 (N_17279,N_15579,N_16133);
nor U17280 (N_17280,N_15274,N_15083);
and U17281 (N_17281,N_15325,N_15280);
or U17282 (N_17282,N_16430,N_15292);
or U17283 (N_17283,N_16439,N_15048);
or U17284 (N_17284,N_15909,N_15876);
or U17285 (N_17285,N_16363,N_15989);
nor U17286 (N_17286,N_15406,N_15433);
nand U17287 (N_17287,N_15490,N_15538);
nand U17288 (N_17288,N_15347,N_15335);
and U17289 (N_17289,N_15752,N_15575);
or U17290 (N_17290,N_16151,N_16174);
and U17291 (N_17291,N_16093,N_16459);
nand U17292 (N_17292,N_16039,N_15156);
nand U17293 (N_17293,N_16267,N_15677);
xor U17294 (N_17294,N_16466,N_16446);
nor U17295 (N_17295,N_16090,N_15578);
nand U17296 (N_17296,N_15400,N_15755);
nand U17297 (N_17297,N_15552,N_15621);
xor U17298 (N_17298,N_16333,N_15849);
nor U17299 (N_17299,N_16033,N_16493);
nand U17300 (N_17300,N_15981,N_15542);
nand U17301 (N_17301,N_16482,N_15619);
and U17302 (N_17302,N_16324,N_15787);
nand U17303 (N_17303,N_16272,N_16105);
or U17304 (N_17304,N_15254,N_16435);
or U17305 (N_17305,N_15161,N_15853);
and U17306 (N_17306,N_16373,N_15444);
and U17307 (N_17307,N_15373,N_15897);
nand U17308 (N_17308,N_15260,N_16298);
xor U17309 (N_17309,N_15454,N_15160);
nand U17310 (N_17310,N_15848,N_16016);
xnor U17311 (N_17311,N_16474,N_16046);
or U17312 (N_17312,N_16391,N_15514);
or U17313 (N_17313,N_15793,N_15878);
xor U17314 (N_17314,N_15477,N_15431);
or U17315 (N_17315,N_15128,N_16396);
xnor U17316 (N_17316,N_15270,N_15225);
nor U17317 (N_17317,N_15163,N_15967);
xnor U17318 (N_17318,N_16468,N_15312);
xnor U17319 (N_17319,N_16330,N_15762);
or U17320 (N_17320,N_15524,N_16007);
nand U17321 (N_17321,N_16169,N_16301);
and U17322 (N_17322,N_15454,N_15376);
nand U17323 (N_17323,N_15005,N_16150);
nand U17324 (N_17324,N_15410,N_15601);
or U17325 (N_17325,N_16357,N_16445);
and U17326 (N_17326,N_15677,N_15832);
nor U17327 (N_17327,N_15485,N_16158);
or U17328 (N_17328,N_15622,N_15898);
nor U17329 (N_17329,N_15828,N_16456);
nor U17330 (N_17330,N_15874,N_16225);
or U17331 (N_17331,N_16238,N_16113);
xnor U17332 (N_17332,N_16230,N_15684);
nand U17333 (N_17333,N_16318,N_15600);
nor U17334 (N_17334,N_15698,N_15308);
nand U17335 (N_17335,N_16261,N_16438);
and U17336 (N_17336,N_15239,N_15576);
nor U17337 (N_17337,N_15919,N_16113);
nor U17338 (N_17338,N_15439,N_16363);
or U17339 (N_17339,N_16370,N_15094);
nor U17340 (N_17340,N_15961,N_15082);
and U17341 (N_17341,N_15921,N_16123);
nand U17342 (N_17342,N_15714,N_15472);
or U17343 (N_17343,N_16342,N_15940);
or U17344 (N_17344,N_15607,N_15223);
and U17345 (N_17345,N_16199,N_15943);
or U17346 (N_17346,N_16253,N_16400);
xor U17347 (N_17347,N_15811,N_15843);
or U17348 (N_17348,N_16494,N_16135);
nand U17349 (N_17349,N_16182,N_15985);
nor U17350 (N_17350,N_15918,N_15907);
nand U17351 (N_17351,N_16428,N_15044);
xor U17352 (N_17352,N_16038,N_15380);
and U17353 (N_17353,N_16142,N_15623);
nand U17354 (N_17354,N_16147,N_15993);
or U17355 (N_17355,N_16099,N_15830);
nand U17356 (N_17356,N_15453,N_15219);
and U17357 (N_17357,N_15777,N_15393);
nand U17358 (N_17358,N_15414,N_15121);
nor U17359 (N_17359,N_15839,N_15208);
nor U17360 (N_17360,N_15971,N_15348);
and U17361 (N_17361,N_16400,N_16256);
nand U17362 (N_17362,N_16151,N_15620);
or U17363 (N_17363,N_15804,N_15991);
nand U17364 (N_17364,N_15678,N_15331);
or U17365 (N_17365,N_15567,N_15391);
and U17366 (N_17366,N_15273,N_16047);
and U17367 (N_17367,N_15800,N_15968);
xnor U17368 (N_17368,N_15623,N_15377);
and U17369 (N_17369,N_16309,N_16041);
nor U17370 (N_17370,N_16196,N_16362);
or U17371 (N_17371,N_16083,N_16064);
and U17372 (N_17372,N_16142,N_16477);
and U17373 (N_17373,N_15556,N_16376);
nand U17374 (N_17374,N_16065,N_16082);
nand U17375 (N_17375,N_16174,N_15641);
nor U17376 (N_17376,N_16011,N_15746);
and U17377 (N_17377,N_15553,N_15328);
and U17378 (N_17378,N_16235,N_15839);
and U17379 (N_17379,N_15844,N_15778);
nor U17380 (N_17380,N_15325,N_16026);
nor U17381 (N_17381,N_15080,N_15688);
nor U17382 (N_17382,N_16247,N_16078);
xor U17383 (N_17383,N_15665,N_15074);
or U17384 (N_17384,N_15265,N_15948);
and U17385 (N_17385,N_16004,N_16144);
nor U17386 (N_17386,N_16477,N_15797);
or U17387 (N_17387,N_16387,N_15720);
xnor U17388 (N_17388,N_15834,N_15789);
or U17389 (N_17389,N_15615,N_15156);
nand U17390 (N_17390,N_15700,N_15934);
nand U17391 (N_17391,N_16365,N_15783);
xnor U17392 (N_17392,N_16075,N_16137);
xor U17393 (N_17393,N_16056,N_15307);
or U17394 (N_17394,N_15445,N_15146);
or U17395 (N_17395,N_15112,N_16000);
nand U17396 (N_17396,N_15047,N_16493);
nor U17397 (N_17397,N_15268,N_16331);
and U17398 (N_17398,N_16492,N_15284);
or U17399 (N_17399,N_15160,N_15608);
nand U17400 (N_17400,N_15946,N_16383);
nand U17401 (N_17401,N_16374,N_15189);
nor U17402 (N_17402,N_15219,N_15896);
and U17403 (N_17403,N_16471,N_16398);
or U17404 (N_17404,N_15671,N_15879);
nor U17405 (N_17405,N_16314,N_15824);
xnor U17406 (N_17406,N_15307,N_15803);
nand U17407 (N_17407,N_15539,N_16183);
or U17408 (N_17408,N_15588,N_16005);
nand U17409 (N_17409,N_15199,N_15913);
or U17410 (N_17410,N_16313,N_15541);
and U17411 (N_17411,N_15847,N_15779);
nor U17412 (N_17412,N_16123,N_16488);
nor U17413 (N_17413,N_15174,N_15566);
xor U17414 (N_17414,N_15902,N_15912);
and U17415 (N_17415,N_16256,N_16081);
nor U17416 (N_17416,N_15010,N_15540);
xnor U17417 (N_17417,N_15885,N_15986);
nor U17418 (N_17418,N_16246,N_15052);
xor U17419 (N_17419,N_15224,N_16239);
and U17420 (N_17420,N_15798,N_15768);
and U17421 (N_17421,N_15941,N_16291);
and U17422 (N_17422,N_15141,N_16078);
or U17423 (N_17423,N_15569,N_15397);
nand U17424 (N_17424,N_15422,N_15122);
or U17425 (N_17425,N_16124,N_16349);
xnor U17426 (N_17426,N_15015,N_15296);
xnor U17427 (N_17427,N_15636,N_16012);
and U17428 (N_17428,N_15179,N_15151);
and U17429 (N_17429,N_15476,N_15758);
xor U17430 (N_17430,N_15467,N_15977);
nor U17431 (N_17431,N_15613,N_15670);
xnor U17432 (N_17432,N_16334,N_15709);
nor U17433 (N_17433,N_16180,N_16066);
and U17434 (N_17434,N_15245,N_15421);
or U17435 (N_17435,N_15285,N_15923);
xor U17436 (N_17436,N_15311,N_16301);
xnor U17437 (N_17437,N_15734,N_16125);
nor U17438 (N_17438,N_16266,N_15839);
xnor U17439 (N_17439,N_15629,N_15043);
and U17440 (N_17440,N_16401,N_16001);
xor U17441 (N_17441,N_15235,N_15957);
nor U17442 (N_17442,N_15022,N_15909);
and U17443 (N_17443,N_16338,N_15575);
xnor U17444 (N_17444,N_15321,N_15880);
and U17445 (N_17445,N_16491,N_15583);
and U17446 (N_17446,N_16106,N_15719);
or U17447 (N_17447,N_15529,N_15267);
nor U17448 (N_17448,N_16269,N_16081);
nor U17449 (N_17449,N_16111,N_16068);
nand U17450 (N_17450,N_15484,N_15412);
and U17451 (N_17451,N_15475,N_15022);
nand U17452 (N_17452,N_15408,N_15341);
xor U17453 (N_17453,N_16092,N_16056);
xor U17454 (N_17454,N_16163,N_15462);
and U17455 (N_17455,N_15374,N_15231);
xnor U17456 (N_17456,N_16406,N_15583);
nand U17457 (N_17457,N_15192,N_15980);
or U17458 (N_17458,N_15882,N_16149);
nor U17459 (N_17459,N_15226,N_15412);
and U17460 (N_17460,N_15480,N_16452);
nor U17461 (N_17461,N_15997,N_15018);
and U17462 (N_17462,N_15467,N_16402);
and U17463 (N_17463,N_15237,N_15084);
or U17464 (N_17464,N_15431,N_15694);
xor U17465 (N_17465,N_15417,N_15386);
nand U17466 (N_17466,N_15086,N_16327);
nand U17467 (N_17467,N_15328,N_16416);
nor U17468 (N_17468,N_16120,N_15001);
or U17469 (N_17469,N_16034,N_15614);
nor U17470 (N_17470,N_15208,N_15711);
nand U17471 (N_17471,N_15245,N_16039);
or U17472 (N_17472,N_16030,N_16451);
nand U17473 (N_17473,N_16181,N_15297);
nand U17474 (N_17474,N_15438,N_15300);
and U17475 (N_17475,N_15307,N_15794);
or U17476 (N_17476,N_15843,N_15609);
xor U17477 (N_17477,N_15764,N_15181);
nand U17478 (N_17478,N_16462,N_15720);
nor U17479 (N_17479,N_15151,N_15425);
nor U17480 (N_17480,N_15560,N_15221);
nand U17481 (N_17481,N_15233,N_15664);
nand U17482 (N_17482,N_15177,N_15146);
xor U17483 (N_17483,N_15167,N_16293);
nor U17484 (N_17484,N_16078,N_15931);
and U17485 (N_17485,N_16103,N_15583);
and U17486 (N_17486,N_15865,N_15967);
and U17487 (N_17487,N_15662,N_15482);
xnor U17488 (N_17488,N_16140,N_15192);
nor U17489 (N_17489,N_15526,N_15110);
and U17490 (N_17490,N_15925,N_16318);
xnor U17491 (N_17491,N_15643,N_15444);
or U17492 (N_17492,N_15441,N_15552);
xnor U17493 (N_17493,N_16234,N_16208);
xor U17494 (N_17494,N_15599,N_15792);
nor U17495 (N_17495,N_16268,N_15909);
nor U17496 (N_17496,N_15540,N_15922);
and U17497 (N_17497,N_16353,N_15263);
nand U17498 (N_17498,N_16079,N_16260);
xor U17499 (N_17499,N_16376,N_16191);
xnor U17500 (N_17500,N_16128,N_16089);
or U17501 (N_17501,N_15593,N_16398);
nand U17502 (N_17502,N_16228,N_15801);
nand U17503 (N_17503,N_15217,N_15089);
xnor U17504 (N_17504,N_15675,N_16018);
or U17505 (N_17505,N_15418,N_15271);
nor U17506 (N_17506,N_15399,N_16223);
or U17507 (N_17507,N_15157,N_15113);
nand U17508 (N_17508,N_15337,N_15850);
xnor U17509 (N_17509,N_16119,N_16450);
nor U17510 (N_17510,N_15000,N_16045);
nor U17511 (N_17511,N_16313,N_15033);
and U17512 (N_17512,N_15468,N_15593);
or U17513 (N_17513,N_15354,N_15409);
nor U17514 (N_17514,N_15560,N_15429);
xnor U17515 (N_17515,N_15764,N_15451);
or U17516 (N_17516,N_16163,N_16327);
or U17517 (N_17517,N_16015,N_15212);
or U17518 (N_17518,N_15778,N_15563);
and U17519 (N_17519,N_15277,N_15841);
nor U17520 (N_17520,N_16221,N_15412);
xnor U17521 (N_17521,N_16399,N_15374);
nand U17522 (N_17522,N_16265,N_16235);
and U17523 (N_17523,N_16411,N_15267);
xnor U17524 (N_17524,N_15287,N_16376);
and U17525 (N_17525,N_15916,N_15784);
and U17526 (N_17526,N_15586,N_15851);
and U17527 (N_17527,N_16467,N_15392);
xnor U17528 (N_17528,N_15090,N_15771);
and U17529 (N_17529,N_15400,N_15745);
nor U17530 (N_17530,N_15692,N_16413);
xnor U17531 (N_17531,N_16374,N_16211);
nor U17532 (N_17532,N_16348,N_16170);
nand U17533 (N_17533,N_16038,N_16096);
or U17534 (N_17534,N_15216,N_15439);
nor U17535 (N_17535,N_16181,N_15536);
nor U17536 (N_17536,N_15389,N_15783);
xnor U17537 (N_17537,N_15865,N_16393);
xor U17538 (N_17538,N_16204,N_16421);
xor U17539 (N_17539,N_16356,N_16248);
or U17540 (N_17540,N_15913,N_15836);
and U17541 (N_17541,N_16383,N_15992);
xor U17542 (N_17542,N_15756,N_15779);
and U17543 (N_17543,N_16214,N_16476);
xor U17544 (N_17544,N_16249,N_16138);
nor U17545 (N_17545,N_15274,N_15398);
and U17546 (N_17546,N_15620,N_16100);
and U17547 (N_17547,N_15182,N_15657);
nor U17548 (N_17548,N_15527,N_15828);
nor U17549 (N_17549,N_16281,N_16410);
and U17550 (N_17550,N_15309,N_16045);
nand U17551 (N_17551,N_16277,N_15142);
nor U17552 (N_17552,N_16477,N_15232);
or U17553 (N_17553,N_16018,N_15056);
and U17554 (N_17554,N_16459,N_16200);
or U17555 (N_17555,N_15081,N_16168);
xnor U17556 (N_17556,N_16459,N_16235);
nand U17557 (N_17557,N_16163,N_16498);
nand U17558 (N_17558,N_15601,N_15803);
or U17559 (N_17559,N_16205,N_15811);
nor U17560 (N_17560,N_15931,N_15143);
and U17561 (N_17561,N_15935,N_15442);
or U17562 (N_17562,N_16370,N_15114);
nor U17563 (N_17563,N_15914,N_15745);
xor U17564 (N_17564,N_15670,N_16305);
nor U17565 (N_17565,N_16319,N_15606);
nand U17566 (N_17566,N_15668,N_15686);
nand U17567 (N_17567,N_15539,N_15284);
and U17568 (N_17568,N_15824,N_15169);
nand U17569 (N_17569,N_16438,N_15416);
nand U17570 (N_17570,N_16270,N_15655);
xor U17571 (N_17571,N_15403,N_15666);
nand U17572 (N_17572,N_15223,N_15833);
or U17573 (N_17573,N_15388,N_15527);
nand U17574 (N_17574,N_15487,N_15517);
and U17575 (N_17575,N_15438,N_15550);
nand U17576 (N_17576,N_16407,N_16329);
or U17577 (N_17577,N_15020,N_15398);
nand U17578 (N_17578,N_16038,N_15245);
xor U17579 (N_17579,N_15125,N_15684);
nand U17580 (N_17580,N_15901,N_15257);
nor U17581 (N_17581,N_15075,N_16272);
or U17582 (N_17582,N_15947,N_16394);
xnor U17583 (N_17583,N_15409,N_16379);
xnor U17584 (N_17584,N_16415,N_15563);
and U17585 (N_17585,N_16464,N_15428);
nor U17586 (N_17586,N_15811,N_16200);
xor U17587 (N_17587,N_15712,N_16416);
nand U17588 (N_17588,N_15887,N_15495);
nand U17589 (N_17589,N_16240,N_16221);
nor U17590 (N_17590,N_15383,N_16143);
or U17591 (N_17591,N_16134,N_15671);
and U17592 (N_17592,N_15176,N_15725);
nor U17593 (N_17593,N_15852,N_15164);
nor U17594 (N_17594,N_15665,N_15324);
xor U17595 (N_17595,N_15968,N_15847);
or U17596 (N_17596,N_15308,N_15934);
and U17597 (N_17597,N_15106,N_15719);
nor U17598 (N_17598,N_15403,N_15686);
or U17599 (N_17599,N_16152,N_15166);
nor U17600 (N_17600,N_15399,N_15955);
xor U17601 (N_17601,N_16351,N_15487);
xor U17602 (N_17602,N_15101,N_16321);
nor U17603 (N_17603,N_15506,N_15007);
and U17604 (N_17604,N_16426,N_16113);
nand U17605 (N_17605,N_15655,N_15719);
xor U17606 (N_17606,N_16088,N_15524);
nor U17607 (N_17607,N_15272,N_15566);
xor U17608 (N_17608,N_16329,N_16217);
nand U17609 (N_17609,N_15338,N_16410);
or U17610 (N_17610,N_16104,N_15081);
and U17611 (N_17611,N_15492,N_15253);
and U17612 (N_17612,N_15611,N_15804);
xor U17613 (N_17613,N_16374,N_16174);
xor U17614 (N_17614,N_16123,N_15147);
xor U17615 (N_17615,N_15141,N_15817);
xor U17616 (N_17616,N_16417,N_16354);
or U17617 (N_17617,N_15553,N_15418);
nor U17618 (N_17618,N_15466,N_16134);
and U17619 (N_17619,N_15126,N_15443);
xnor U17620 (N_17620,N_15889,N_16047);
xor U17621 (N_17621,N_15206,N_15537);
nand U17622 (N_17622,N_15163,N_15425);
xnor U17623 (N_17623,N_16167,N_15528);
nand U17624 (N_17624,N_15104,N_16425);
nor U17625 (N_17625,N_16467,N_15505);
xor U17626 (N_17626,N_15357,N_15782);
nand U17627 (N_17627,N_16093,N_15113);
or U17628 (N_17628,N_16451,N_15453);
nor U17629 (N_17629,N_15541,N_15609);
or U17630 (N_17630,N_16369,N_15045);
nor U17631 (N_17631,N_15731,N_16017);
nor U17632 (N_17632,N_15074,N_15211);
nand U17633 (N_17633,N_15842,N_16385);
nand U17634 (N_17634,N_15174,N_15062);
nand U17635 (N_17635,N_15913,N_15742);
and U17636 (N_17636,N_16166,N_16110);
or U17637 (N_17637,N_16044,N_16451);
or U17638 (N_17638,N_15836,N_15136);
xor U17639 (N_17639,N_16012,N_16123);
xor U17640 (N_17640,N_16396,N_15782);
xnor U17641 (N_17641,N_15165,N_15303);
nor U17642 (N_17642,N_15055,N_15654);
xnor U17643 (N_17643,N_15451,N_15546);
nor U17644 (N_17644,N_16183,N_16432);
and U17645 (N_17645,N_16406,N_16340);
nor U17646 (N_17646,N_15240,N_15271);
or U17647 (N_17647,N_15130,N_16116);
or U17648 (N_17648,N_15010,N_15309);
and U17649 (N_17649,N_15209,N_15575);
and U17650 (N_17650,N_16483,N_16115);
xor U17651 (N_17651,N_15875,N_16252);
nand U17652 (N_17652,N_16317,N_15653);
or U17653 (N_17653,N_15506,N_15499);
nand U17654 (N_17654,N_15576,N_16202);
xor U17655 (N_17655,N_15569,N_15561);
nand U17656 (N_17656,N_16434,N_15893);
and U17657 (N_17657,N_16108,N_16316);
nor U17658 (N_17658,N_15994,N_15410);
nor U17659 (N_17659,N_16357,N_16300);
nor U17660 (N_17660,N_16194,N_15626);
nand U17661 (N_17661,N_15409,N_16027);
xnor U17662 (N_17662,N_15111,N_16098);
and U17663 (N_17663,N_15574,N_15253);
xnor U17664 (N_17664,N_15094,N_15269);
or U17665 (N_17665,N_16118,N_15933);
xor U17666 (N_17666,N_16119,N_15830);
xnor U17667 (N_17667,N_16233,N_16028);
nand U17668 (N_17668,N_15762,N_15687);
nand U17669 (N_17669,N_16435,N_15862);
or U17670 (N_17670,N_15953,N_15450);
and U17671 (N_17671,N_15795,N_15738);
nor U17672 (N_17672,N_16027,N_15775);
xnor U17673 (N_17673,N_15970,N_15709);
or U17674 (N_17674,N_15762,N_15696);
xnor U17675 (N_17675,N_15194,N_16428);
nor U17676 (N_17676,N_15428,N_15324);
nor U17677 (N_17677,N_16414,N_15925);
nand U17678 (N_17678,N_15456,N_16469);
or U17679 (N_17679,N_15566,N_15882);
nor U17680 (N_17680,N_15511,N_15858);
and U17681 (N_17681,N_15015,N_15997);
or U17682 (N_17682,N_15633,N_15442);
nand U17683 (N_17683,N_16108,N_16437);
nand U17684 (N_17684,N_16035,N_15120);
xor U17685 (N_17685,N_15465,N_15521);
and U17686 (N_17686,N_16050,N_15964);
and U17687 (N_17687,N_15139,N_15878);
xnor U17688 (N_17688,N_15566,N_15037);
xor U17689 (N_17689,N_15545,N_15996);
xnor U17690 (N_17690,N_15312,N_16240);
or U17691 (N_17691,N_15787,N_15449);
nand U17692 (N_17692,N_15994,N_16388);
nor U17693 (N_17693,N_16078,N_16208);
or U17694 (N_17694,N_15248,N_16418);
or U17695 (N_17695,N_15190,N_16315);
or U17696 (N_17696,N_15566,N_15406);
nand U17697 (N_17697,N_15043,N_16124);
nor U17698 (N_17698,N_15289,N_15942);
xnor U17699 (N_17699,N_15621,N_15282);
nand U17700 (N_17700,N_15580,N_15573);
nor U17701 (N_17701,N_16041,N_15122);
nand U17702 (N_17702,N_15504,N_16332);
or U17703 (N_17703,N_15989,N_16060);
or U17704 (N_17704,N_16263,N_15624);
nor U17705 (N_17705,N_16047,N_15503);
xnor U17706 (N_17706,N_16263,N_15067);
nor U17707 (N_17707,N_15984,N_15690);
nor U17708 (N_17708,N_16183,N_16346);
and U17709 (N_17709,N_16108,N_15565);
nand U17710 (N_17710,N_15134,N_15822);
and U17711 (N_17711,N_15722,N_16164);
or U17712 (N_17712,N_15594,N_15770);
nand U17713 (N_17713,N_15615,N_15572);
and U17714 (N_17714,N_15567,N_15382);
nand U17715 (N_17715,N_16143,N_15472);
or U17716 (N_17716,N_15320,N_15257);
nand U17717 (N_17717,N_16472,N_15918);
or U17718 (N_17718,N_15813,N_16412);
and U17719 (N_17719,N_15037,N_16323);
nor U17720 (N_17720,N_15908,N_15868);
nor U17721 (N_17721,N_15455,N_15162);
nor U17722 (N_17722,N_15388,N_15148);
xor U17723 (N_17723,N_15345,N_16489);
nand U17724 (N_17724,N_15374,N_15829);
nor U17725 (N_17725,N_16215,N_15064);
xnor U17726 (N_17726,N_15187,N_15908);
and U17727 (N_17727,N_16172,N_15318);
xnor U17728 (N_17728,N_15388,N_15553);
and U17729 (N_17729,N_15334,N_15476);
nor U17730 (N_17730,N_15052,N_15648);
nand U17731 (N_17731,N_15813,N_16305);
nand U17732 (N_17732,N_15959,N_16214);
or U17733 (N_17733,N_15521,N_15366);
and U17734 (N_17734,N_15866,N_15527);
and U17735 (N_17735,N_15965,N_15350);
nand U17736 (N_17736,N_15175,N_15260);
or U17737 (N_17737,N_16472,N_15017);
or U17738 (N_17738,N_16387,N_15454);
nor U17739 (N_17739,N_16446,N_16423);
and U17740 (N_17740,N_16048,N_15853);
nor U17741 (N_17741,N_15992,N_15218);
nor U17742 (N_17742,N_15265,N_16242);
nor U17743 (N_17743,N_15841,N_15150);
xnor U17744 (N_17744,N_15184,N_15290);
and U17745 (N_17745,N_15572,N_16198);
or U17746 (N_17746,N_15290,N_16336);
xor U17747 (N_17747,N_15539,N_16360);
nor U17748 (N_17748,N_16476,N_16399);
nand U17749 (N_17749,N_15285,N_16270);
nor U17750 (N_17750,N_15165,N_16025);
and U17751 (N_17751,N_15454,N_15685);
nor U17752 (N_17752,N_15817,N_15380);
or U17753 (N_17753,N_16193,N_15685);
nor U17754 (N_17754,N_15089,N_15291);
xnor U17755 (N_17755,N_16028,N_15038);
or U17756 (N_17756,N_15990,N_15444);
or U17757 (N_17757,N_15744,N_16164);
nand U17758 (N_17758,N_16285,N_16295);
nand U17759 (N_17759,N_15264,N_16472);
nand U17760 (N_17760,N_15062,N_15443);
or U17761 (N_17761,N_15516,N_15552);
xnor U17762 (N_17762,N_16288,N_15255);
nand U17763 (N_17763,N_15566,N_16083);
nand U17764 (N_17764,N_15121,N_15301);
or U17765 (N_17765,N_15999,N_15509);
or U17766 (N_17766,N_15232,N_16489);
nand U17767 (N_17767,N_15307,N_15903);
nand U17768 (N_17768,N_15786,N_16388);
nand U17769 (N_17769,N_15582,N_15930);
nor U17770 (N_17770,N_16003,N_15836);
or U17771 (N_17771,N_15019,N_15074);
and U17772 (N_17772,N_15659,N_15298);
or U17773 (N_17773,N_15258,N_15752);
xnor U17774 (N_17774,N_15199,N_15969);
or U17775 (N_17775,N_16423,N_15042);
xnor U17776 (N_17776,N_15243,N_15695);
nor U17777 (N_17777,N_15934,N_15158);
or U17778 (N_17778,N_16018,N_15911);
nor U17779 (N_17779,N_15631,N_15528);
xor U17780 (N_17780,N_15254,N_16470);
xor U17781 (N_17781,N_16278,N_15890);
nand U17782 (N_17782,N_16314,N_16449);
and U17783 (N_17783,N_15673,N_16205);
and U17784 (N_17784,N_16055,N_15892);
nor U17785 (N_17785,N_15020,N_15140);
nor U17786 (N_17786,N_15194,N_15901);
nand U17787 (N_17787,N_15344,N_16088);
nor U17788 (N_17788,N_16293,N_15657);
xnor U17789 (N_17789,N_15820,N_16036);
nand U17790 (N_17790,N_16273,N_15427);
and U17791 (N_17791,N_16141,N_15139);
nor U17792 (N_17792,N_16231,N_15723);
and U17793 (N_17793,N_15027,N_16379);
xnor U17794 (N_17794,N_16356,N_15759);
nor U17795 (N_17795,N_16211,N_15828);
xor U17796 (N_17796,N_16267,N_15755);
nand U17797 (N_17797,N_15043,N_16029);
nand U17798 (N_17798,N_15153,N_15514);
xnor U17799 (N_17799,N_16406,N_16193);
nand U17800 (N_17800,N_15591,N_16184);
nand U17801 (N_17801,N_16488,N_15322);
and U17802 (N_17802,N_15688,N_15671);
and U17803 (N_17803,N_15482,N_15943);
and U17804 (N_17804,N_15786,N_16460);
nor U17805 (N_17805,N_15537,N_16146);
nand U17806 (N_17806,N_16076,N_16414);
nor U17807 (N_17807,N_16457,N_15440);
and U17808 (N_17808,N_15909,N_15275);
nand U17809 (N_17809,N_15565,N_15440);
or U17810 (N_17810,N_16324,N_15024);
and U17811 (N_17811,N_16207,N_15087);
or U17812 (N_17812,N_15506,N_15461);
xnor U17813 (N_17813,N_16129,N_15855);
and U17814 (N_17814,N_15688,N_16495);
nand U17815 (N_17815,N_15394,N_16164);
and U17816 (N_17816,N_16216,N_16366);
or U17817 (N_17817,N_15181,N_15747);
nor U17818 (N_17818,N_15121,N_15359);
nand U17819 (N_17819,N_15098,N_15625);
and U17820 (N_17820,N_15360,N_15629);
and U17821 (N_17821,N_15584,N_15137);
nand U17822 (N_17822,N_16088,N_15222);
nand U17823 (N_17823,N_15812,N_15964);
and U17824 (N_17824,N_15660,N_15265);
or U17825 (N_17825,N_16391,N_15231);
and U17826 (N_17826,N_15938,N_15740);
or U17827 (N_17827,N_16399,N_15249);
and U17828 (N_17828,N_15269,N_15702);
or U17829 (N_17829,N_16198,N_16051);
or U17830 (N_17830,N_15708,N_16174);
nand U17831 (N_17831,N_15514,N_15596);
and U17832 (N_17832,N_16073,N_15068);
or U17833 (N_17833,N_15823,N_15388);
nor U17834 (N_17834,N_15405,N_15155);
or U17835 (N_17835,N_16326,N_16179);
nand U17836 (N_17836,N_15330,N_15018);
xnor U17837 (N_17837,N_15102,N_15863);
and U17838 (N_17838,N_15670,N_16381);
nor U17839 (N_17839,N_16202,N_15102);
xor U17840 (N_17840,N_15545,N_15112);
nor U17841 (N_17841,N_15072,N_15802);
and U17842 (N_17842,N_15496,N_15105);
and U17843 (N_17843,N_15446,N_15629);
nor U17844 (N_17844,N_15369,N_15856);
or U17845 (N_17845,N_15814,N_16406);
xor U17846 (N_17846,N_16174,N_16236);
xnor U17847 (N_17847,N_16188,N_15305);
nand U17848 (N_17848,N_15590,N_16081);
nor U17849 (N_17849,N_16160,N_15613);
or U17850 (N_17850,N_15301,N_15201);
and U17851 (N_17851,N_15055,N_15399);
xnor U17852 (N_17852,N_15446,N_15946);
xor U17853 (N_17853,N_15500,N_16097);
nor U17854 (N_17854,N_15524,N_15664);
and U17855 (N_17855,N_15227,N_16217);
nor U17856 (N_17856,N_15192,N_15337);
nor U17857 (N_17857,N_15382,N_15405);
nor U17858 (N_17858,N_15898,N_15610);
and U17859 (N_17859,N_16106,N_15512);
and U17860 (N_17860,N_16402,N_15098);
xor U17861 (N_17861,N_16482,N_15075);
nor U17862 (N_17862,N_15434,N_15462);
or U17863 (N_17863,N_16344,N_16301);
nand U17864 (N_17864,N_16353,N_15587);
nand U17865 (N_17865,N_15124,N_15716);
and U17866 (N_17866,N_16335,N_16320);
and U17867 (N_17867,N_16363,N_15892);
or U17868 (N_17868,N_16349,N_15475);
or U17869 (N_17869,N_15296,N_16025);
nand U17870 (N_17870,N_16403,N_16270);
nor U17871 (N_17871,N_15515,N_15283);
and U17872 (N_17872,N_16164,N_15067);
and U17873 (N_17873,N_15654,N_15574);
nor U17874 (N_17874,N_16044,N_15949);
or U17875 (N_17875,N_15081,N_16281);
nand U17876 (N_17876,N_15949,N_16203);
nor U17877 (N_17877,N_15890,N_15448);
and U17878 (N_17878,N_16052,N_15022);
or U17879 (N_17879,N_16397,N_16244);
xnor U17880 (N_17880,N_15072,N_16190);
and U17881 (N_17881,N_15493,N_15126);
nand U17882 (N_17882,N_15101,N_16120);
and U17883 (N_17883,N_15926,N_15846);
nor U17884 (N_17884,N_16300,N_15964);
nor U17885 (N_17885,N_15751,N_16195);
nand U17886 (N_17886,N_15440,N_15049);
or U17887 (N_17887,N_15975,N_16109);
and U17888 (N_17888,N_15119,N_15595);
xor U17889 (N_17889,N_16477,N_15757);
xnor U17890 (N_17890,N_15325,N_16161);
or U17891 (N_17891,N_15886,N_15860);
xnor U17892 (N_17892,N_15827,N_15591);
xnor U17893 (N_17893,N_15010,N_15043);
or U17894 (N_17894,N_15106,N_15948);
nand U17895 (N_17895,N_16287,N_15740);
or U17896 (N_17896,N_15250,N_15400);
or U17897 (N_17897,N_15973,N_15701);
xor U17898 (N_17898,N_15151,N_15708);
xnor U17899 (N_17899,N_15494,N_16150);
or U17900 (N_17900,N_16449,N_16088);
or U17901 (N_17901,N_15136,N_15019);
and U17902 (N_17902,N_15257,N_16452);
nor U17903 (N_17903,N_15228,N_15899);
xnor U17904 (N_17904,N_16160,N_16004);
or U17905 (N_17905,N_15072,N_16295);
and U17906 (N_17906,N_15507,N_15614);
nand U17907 (N_17907,N_15300,N_15537);
nand U17908 (N_17908,N_15077,N_16170);
xnor U17909 (N_17909,N_15413,N_15030);
xor U17910 (N_17910,N_15835,N_16043);
nor U17911 (N_17911,N_15750,N_16114);
xnor U17912 (N_17912,N_15491,N_15545);
nand U17913 (N_17913,N_15538,N_15207);
and U17914 (N_17914,N_15248,N_16192);
xor U17915 (N_17915,N_15816,N_16129);
nand U17916 (N_17916,N_15647,N_16445);
or U17917 (N_17917,N_15669,N_16450);
xnor U17918 (N_17918,N_15710,N_15733);
xnor U17919 (N_17919,N_16068,N_15801);
nor U17920 (N_17920,N_15553,N_16012);
nand U17921 (N_17921,N_15469,N_15293);
or U17922 (N_17922,N_15218,N_15050);
and U17923 (N_17923,N_15611,N_15737);
nand U17924 (N_17924,N_15393,N_15526);
and U17925 (N_17925,N_16107,N_16099);
and U17926 (N_17926,N_16423,N_15178);
nand U17927 (N_17927,N_16074,N_15593);
and U17928 (N_17928,N_15108,N_15764);
nand U17929 (N_17929,N_15612,N_16337);
and U17930 (N_17930,N_15259,N_16434);
nand U17931 (N_17931,N_15647,N_16263);
or U17932 (N_17932,N_15647,N_15885);
or U17933 (N_17933,N_15720,N_15566);
xnor U17934 (N_17934,N_15208,N_15718);
xor U17935 (N_17935,N_16329,N_16467);
or U17936 (N_17936,N_15434,N_15994);
nor U17937 (N_17937,N_16353,N_15700);
and U17938 (N_17938,N_15768,N_16399);
or U17939 (N_17939,N_15690,N_15492);
nor U17940 (N_17940,N_15510,N_15677);
nand U17941 (N_17941,N_16212,N_16182);
or U17942 (N_17942,N_16294,N_15476);
nor U17943 (N_17943,N_16256,N_16445);
xor U17944 (N_17944,N_15954,N_15985);
and U17945 (N_17945,N_15782,N_15816);
and U17946 (N_17946,N_15420,N_16141);
xnor U17947 (N_17947,N_16018,N_15520);
xnor U17948 (N_17948,N_15138,N_16194);
nand U17949 (N_17949,N_15490,N_16145);
nor U17950 (N_17950,N_15311,N_16491);
xor U17951 (N_17951,N_16389,N_16253);
or U17952 (N_17952,N_15292,N_15765);
nand U17953 (N_17953,N_15483,N_15471);
and U17954 (N_17954,N_15052,N_15195);
xnor U17955 (N_17955,N_15463,N_15549);
or U17956 (N_17956,N_15260,N_15045);
nand U17957 (N_17957,N_15969,N_15054);
nor U17958 (N_17958,N_16087,N_15575);
nor U17959 (N_17959,N_16117,N_15896);
nor U17960 (N_17960,N_15308,N_15841);
and U17961 (N_17961,N_15169,N_15466);
nand U17962 (N_17962,N_16017,N_16309);
nor U17963 (N_17963,N_15797,N_15658);
or U17964 (N_17964,N_16429,N_16234);
nand U17965 (N_17965,N_15129,N_16016);
or U17966 (N_17966,N_15632,N_16208);
and U17967 (N_17967,N_15381,N_16049);
or U17968 (N_17968,N_16129,N_15564);
nand U17969 (N_17969,N_16375,N_16259);
or U17970 (N_17970,N_15280,N_15350);
xor U17971 (N_17971,N_15102,N_16457);
nor U17972 (N_17972,N_15203,N_15706);
nand U17973 (N_17973,N_16423,N_15732);
and U17974 (N_17974,N_16003,N_15726);
and U17975 (N_17975,N_15426,N_15853);
xor U17976 (N_17976,N_15355,N_15827);
xor U17977 (N_17977,N_15870,N_16362);
and U17978 (N_17978,N_16497,N_15266);
nor U17979 (N_17979,N_15147,N_15705);
and U17980 (N_17980,N_16319,N_16379);
nor U17981 (N_17981,N_15745,N_15603);
xor U17982 (N_17982,N_15385,N_16270);
nor U17983 (N_17983,N_15128,N_15779);
nand U17984 (N_17984,N_15798,N_15621);
nand U17985 (N_17985,N_15757,N_15931);
or U17986 (N_17986,N_15653,N_15649);
nor U17987 (N_17987,N_15335,N_16172);
or U17988 (N_17988,N_15773,N_16240);
and U17989 (N_17989,N_16059,N_15444);
nor U17990 (N_17990,N_16118,N_15693);
or U17991 (N_17991,N_15345,N_16441);
nand U17992 (N_17992,N_15753,N_16160);
nor U17993 (N_17993,N_15505,N_15344);
or U17994 (N_17994,N_16252,N_15427);
nand U17995 (N_17995,N_15188,N_15535);
or U17996 (N_17996,N_16283,N_16465);
nand U17997 (N_17997,N_15775,N_15671);
and U17998 (N_17998,N_15906,N_15666);
or U17999 (N_17999,N_15733,N_15338);
xnor U18000 (N_18000,N_17219,N_16991);
nor U18001 (N_18001,N_17885,N_16630);
or U18002 (N_18002,N_17036,N_17331);
nor U18003 (N_18003,N_17080,N_16934);
xnor U18004 (N_18004,N_17789,N_16806);
or U18005 (N_18005,N_16675,N_17960);
nand U18006 (N_18006,N_16732,N_16993);
nor U18007 (N_18007,N_16560,N_17049);
xor U18008 (N_18008,N_16725,N_16559);
or U18009 (N_18009,N_17500,N_17377);
or U18010 (N_18010,N_16664,N_17955);
xnor U18011 (N_18011,N_17570,N_17184);
nor U18012 (N_18012,N_17836,N_17233);
and U18013 (N_18013,N_17247,N_17461);
nor U18014 (N_18014,N_17590,N_17581);
xor U18015 (N_18015,N_17245,N_17828);
nor U18016 (N_18016,N_16743,N_17566);
xor U18017 (N_18017,N_17270,N_17772);
or U18018 (N_18018,N_17146,N_16670);
or U18019 (N_18019,N_16709,N_17416);
nor U18020 (N_18020,N_16573,N_17969);
nor U18021 (N_18021,N_17201,N_17453);
and U18022 (N_18022,N_16731,N_17639);
nor U18023 (N_18023,N_17425,N_17872);
nand U18024 (N_18024,N_17317,N_17356);
nor U18025 (N_18025,N_17095,N_17450);
nor U18026 (N_18026,N_17833,N_16811);
nor U18027 (N_18027,N_16584,N_17085);
xnor U18028 (N_18028,N_16947,N_17585);
nand U18029 (N_18029,N_17302,N_16884);
and U18030 (N_18030,N_17547,N_17602);
and U18031 (N_18031,N_17837,N_16631);
xnor U18032 (N_18032,N_16556,N_17409);
or U18033 (N_18033,N_17370,N_17978);
or U18034 (N_18034,N_16536,N_17522);
xnor U18035 (N_18035,N_16909,N_16507);
nor U18036 (N_18036,N_17740,N_17968);
nor U18037 (N_18037,N_16821,N_17708);
xnor U18038 (N_18038,N_17802,N_17880);
xnor U18039 (N_18039,N_17062,N_17505);
nand U18040 (N_18040,N_16707,N_16696);
xnor U18041 (N_18041,N_17207,N_17185);
and U18042 (N_18042,N_17156,N_16988);
nand U18043 (N_18043,N_17709,N_17166);
or U18044 (N_18044,N_17983,N_17520);
and U18045 (N_18045,N_16908,N_17335);
xor U18046 (N_18046,N_16916,N_17799);
nor U18047 (N_18047,N_17819,N_16962);
or U18048 (N_18048,N_17952,N_16865);
and U18049 (N_18049,N_17633,N_16766);
nor U18050 (N_18050,N_17455,N_17167);
or U18051 (N_18051,N_17527,N_17165);
nor U18052 (N_18052,N_17104,N_17869);
nor U18053 (N_18053,N_16983,N_17492);
and U18054 (N_18054,N_17072,N_17599);
and U18055 (N_18055,N_17624,N_17293);
or U18056 (N_18056,N_16537,N_16877);
nand U18057 (N_18057,N_17998,N_17329);
xnor U18058 (N_18058,N_17986,N_16936);
nor U18059 (N_18059,N_17260,N_17621);
nor U18060 (N_18060,N_17741,N_17313);
xor U18061 (N_18061,N_16797,N_16578);
xnor U18062 (N_18062,N_17660,N_17615);
and U18063 (N_18063,N_16717,N_17303);
xor U18064 (N_18064,N_16990,N_16981);
and U18065 (N_18065,N_17804,N_17205);
xor U18066 (N_18066,N_17683,N_17704);
and U18067 (N_18067,N_17060,N_16595);
nand U18068 (N_18068,N_16994,N_17163);
nand U18069 (N_18069,N_16885,N_17116);
xor U18070 (N_18070,N_17812,N_17160);
xor U18071 (N_18071,N_17820,N_17355);
and U18072 (N_18072,N_16554,N_16617);
nor U18073 (N_18073,N_17155,N_17651);
xor U18074 (N_18074,N_17738,N_17099);
or U18075 (N_18075,N_16856,N_16517);
or U18076 (N_18076,N_17857,N_17437);
and U18077 (N_18077,N_16579,N_17550);
nand U18078 (N_18078,N_16532,N_17090);
and U18079 (N_18079,N_17048,N_17171);
nor U18080 (N_18080,N_17491,N_16778);
nand U18081 (N_18081,N_16832,N_16810);
nor U18082 (N_18082,N_17702,N_17136);
nand U18083 (N_18083,N_17903,N_17078);
or U18084 (N_18084,N_17364,N_17597);
nand U18085 (N_18085,N_16921,N_16816);
nor U18086 (N_18086,N_17055,N_16757);
and U18087 (N_18087,N_17554,N_16645);
nand U18088 (N_18088,N_17056,N_16557);
nand U18089 (N_18089,N_16591,N_16683);
or U18090 (N_18090,N_16890,N_17315);
and U18091 (N_18091,N_16765,N_17618);
nand U18092 (N_18092,N_16752,N_16889);
or U18093 (N_18093,N_16639,N_16942);
nand U18094 (N_18094,N_17359,N_17324);
or U18095 (N_18095,N_16817,N_17284);
nor U18096 (N_18096,N_16929,N_17655);
or U18097 (N_18097,N_16710,N_17661);
nor U18098 (N_18098,N_16862,N_17577);
nor U18099 (N_18099,N_17002,N_17456);
or U18100 (N_18100,N_17130,N_16656);
or U18101 (N_18101,N_16924,N_17711);
xor U18102 (N_18102,N_17426,N_16657);
xor U18103 (N_18103,N_16615,N_17948);
xor U18104 (N_18104,N_17332,N_16602);
and U18105 (N_18105,N_16529,N_17699);
and U18106 (N_18106,N_17682,N_17557);
or U18107 (N_18107,N_17148,N_16860);
and U18108 (N_18108,N_17327,N_16576);
nand U18109 (N_18109,N_17912,N_16944);
and U18110 (N_18110,N_17796,N_16728);
or U18111 (N_18111,N_17764,N_17151);
xor U18112 (N_18112,N_17488,N_17777);
nand U18113 (N_18113,N_17606,N_16801);
nand U18114 (N_18114,N_17071,N_16999);
nor U18115 (N_18115,N_17419,N_16650);
nand U18116 (N_18116,N_17914,N_17949);
nand U18117 (N_18117,N_17962,N_17381);
or U18118 (N_18118,N_16516,N_16626);
nor U18119 (N_18119,N_17212,N_17045);
nor U18120 (N_18120,N_16963,N_16510);
nor U18121 (N_18121,N_16665,N_17743);
nand U18122 (N_18122,N_16967,N_17108);
nand U18123 (N_18123,N_17946,N_17530);
xnor U18124 (N_18124,N_16618,N_16718);
or U18125 (N_18125,N_17924,N_17712);
and U18126 (N_18126,N_16744,N_17813);
and U18127 (N_18127,N_17115,N_17287);
xor U18128 (N_18128,N_17288,N_16607);
xnor U18129 (N_18129,N_17626,N_17540);
nor U18130 (N_18130,N_16614,N_16610);
nor U18131 (N_18131,N_17497,N_16756);
nand U18132 (N_18132,N_16506,N_17169);
xor U18133 (N_18133,N_16629,N_17800);
or U18134 (N_18134,N_16694,N_17657);
nor U18135 (N_18135,N_17403,N_16899);
or U18136 (N_18136,N_16603,N_17997);
nor U18137 (N_18137,N_16634,N_17572);
or U18138 (N_18138,N_17395,N_16508);
or U18139 (N_18139,N_16918,N_17263);
nor U18140 (N_18140,N_16969,N_17209);
nor U18141 (N_18141,N_17418,N_17295);
or U18142 (N_18142,N_16850,N_17578);
and U18143 (N_18143,N_17121,N_17069);
or U18144 (N_18144,N_17620,N_17859);
xnor U18145 (N_18145,N_17579,N_16842);
or U18146 (N_18146,N_17018,N_17443);
nor U18147 (N_18147,N_17786,N_17162);
xor U18148 (N_18148,N_16601,N_17979);
nand U18149 (N_18149,N_17451,N_17571);
and U18150 (N_18150,N_17003,N_17230);
xor U18151 (N_18151,N_17725,N_17259);
nor U18152 (N_18152,N_16577,N_17464);
nor U18153 (N_18153,N_17784,N_16872);
nand U18154 (N_18154,N_16612,N_17498);
or U18155 (N_18155,N_17427,N_17797);
nor U18156 (N_18156,N_17243,N_16943);
or U18157 (N_18157,N_17235,N_17011);
and U18158 (N_18158,N_17452,N_17084);
nand U18159 (N_18159,N_17632,N_16653);
nor U18160 (N_18160,N_17719,N_17000);
or U18161 (N_18161,N_17686,N_17818);
or U18162 (N_18162,N_16830,N_17861);
nand U18163 (N_18163,N_17339,N_17191);
or U18164 (N_18164,N_17228,N_17371);
nor U18165 (N_18165,N_16809,N_16950);
and U18166 (N_18166,N_16940,N_16674);
and U18167 (N_18167,N_16592,N_17656);
or U18168 (N_18168,N_16875,N_16952);
xor U18169 (N_18169,N_17507,N_17584);
and U18170 (N_18170,N_16604,N_17417);
nand U18171 (N_18171,N_16677,N_17950);
nand U18172 (N_18172,N_17312,N_16863);
xor U18173 (N_18173,N_17325,N_17009);
nor U18174 (N_18174,N_16813,N_16997);
and U18175 (N_18175,N_17649,N_17052);
xor U18176 (N_18176,N_17470,N_17744);
or U18177 (N_18177,N_17523,N_17938);
nand U18178 (N_18178,N_17139,N_17546);
xnor U18179 (N_18179,N_17931,N_16682);
xor U18180 (N_18180,N_17753,N_17118);
nor U18181 (N_18181,N_17518,N_17053);
or U18182 (N_18182,N_16949,N_16825);
or U18183 (N_18183,N_17189,N_17598);
xnor U18184 (N_18184,N_17899,N_17714);
or U18185 (N_18185,N_17177,N_16763);
and U18186 (N_18186,N_17904,N_16686);
or U18187 (N_18187,N_16791,N_17311);
xor U18188 (N_18188,N_17376,N_17722);
and U18189 (N_18189,N_16805,N_17001);
and U18190 (N_18190,N_17441,N_17194);
nand U18191 (N_18191,N_17246,N_17888);
and U18192 (N_18192,N_16827,N_17771);
nor U18193 (N_18193,N_17856,N_17838);
xnor U18194 (N_18194,N_17769,N_16700);
xor U18195 (N_18195,N_17843,N_16910);
nand U18196 (N_18196,N_16742,N_17094);
or U18197 (N_18197,N_17272,N_17103);
nor U18198 (N_18198,N_16847,N_17958);
and U18199 (N_18199,N_16966,N_16666);
nand U18200 (N_18200,N_16965,N_17064);
xor U18201 (N_18201,N_17258,N_17877);
nand U18202 (N_18202,N_16741,N_16500);
or U18203 (N_18203,N_17398,N_17158);
nand U18204 (N_18204,N_17004,N_16530);
nand U18205 (N_18205,N_17558,N_16520);
or U18206 (N_18206,N_17746,N_17252);
and U18207 (N_18207,N_17951,N_17762);
xor U18208 (N_18208,N_17204,N_17675);
and U18209 (N_18209,N_16745,N_16844);
xor U18210 (N_18210,N_16628,N_17106);
or U18211 (N_18211,N_16734,N_16932);
nor U18212 (N_18212,N_17676,N_17143);
and U18213 (N_18213,N_17442,N_17536);
nor U18214 (N_18214,N_16786,N_17592);
xnor U18215 (N_18215,N_16894,N_16545);
nand U18216 (N_18216,N_17232,N_17641);
and U18217 (N_18217,N_17703,N_17752);
nand U18218 (N_18218,N_16688,N_17605);
xnor U18219 (N_18219,N_17568,N_17231);
xnor U18220 (N_18220,N_17250,N_17733);
nor U18221 (N_18221,N_17567,N_17411);
and U18222 (N_18222,N_17138,N_17369);
or U18223 (N_18223,N_16668,N_17855);
nor U18224 (N_18224,N_17925,N_16635);
nor U18225 (N_18225,N_17357,N_16678);
xor U18226 (N_18226,N_17509,N_17200);
xor U18227 (N_18227,N_16913,N_17975);
or U18228 (N_18228,N_16720,N_16526);
nor U18229 (N_18229,N_16722,N_17467);
xor U18230 (N_18230,N_17432,N_17829);
xor U18231 (N_18231,N_16689,N_17198);
nor U18232 (N_18232,N_17221,N_16960);
nor U18233 (N_18233,N_16712,N_17144);
and U18234 (N_18234,N_17468,N_17197);
xnor U18235 (N_18235,N_17465,N_17767);
xnor U18236 (N_18236,N_17534,N_17351);
xor U18237 (N_18237,N_17292,N_17765);
nor U18238 (N_18238,N_17864,N_17147);
and U18239 (N_18239,N_17511,N_17957);
or U18240 (N_18240,N_17236,N_16546);
or U18241 (N_18241,N_17689,N_17402);
or U18242 (N_18242,N_16833,N_16655);
nor U18243 (N_18243,N_17496,N_16853);
xor U18244 (N_18244,N_17239,N_16767);
nand U18245 (N_18245,N_16902,N_17956);
or U18246 (N_18246,N_16819,N_17024);
xor U18247 (N_18247,N_17430,N_17835);
or U18248 (N_18248,N_17129,N_17543);
nor U18249 (N_18249,N_16954,N_17512);
nand U18250 (N_18250,N_16726,N_17720);
nand U18251 (N_18251,N_17846,N_17029);
xnor U18252 (N_18252,N_17026,N_17379);
nand U18253 (N_18253,N_17273,N_17039);
xor U18254 (N_18254,N_17083,N_17054);
nand U18255 (N_18255,N_17360,N_17613);
nor U18256 (N_18256,N_17806,N_17493);
or U18257 (N_18257,N_16920,N_17695);
xor U18258 (N_18258,N_17612,N_17700);
or U18259 (N_18259,N_17556,N_17739);
nor U18260 (N_18260,N_17440,N_17279);
and U18261 (N_18261,N_17223,N_17323);
nand U18262 (N_18262,N_17349,N_16723);
nand U18263 (N_18263,N_16972,N_17933);
or U18264 (N_18264,N_16616,N_17735);
and U18265 (N_18265,N_17830,N_16669);
xor U18266 (N_18266,N_17017,N_16906);
and U18267 (N_18267,N_16661,N_16534);
nor U18268 (N_18268,N_16676,N_16719);
xor U18269 (N_18269,N_17603,N_17176);
nand U18270 (N_18270,N_17710,N_16880);
or U18271 (N_18271,N_17305,N_16845);
xnor U18272 (N_18272,N_16504,N_17319);
nand U18273 (N_18273,N_17928,N_17448);
nor U18274 (N_18274,N_17215,N_17101);
nor U18275 (N_18275,N_17113,N_17595);
or U18276 (N_18276,N_16690,N_16922);
nor U18277 (N_18277,N_16883,N_16846);
xor U18278 (N_18278,N_17947,N_16637);
nor U18279 (N_18279,N_16695,N_17945);
xor U18280 (N_18280,N_17891,N_17766);
xnor U18281 (N_18281,N_16774,N_16787);
or U18282 (N_18282,N_17199,N_17400);
nand U18283 (N_18283,N_16964,N_17153);
nor U18284 (N_18284,N_17826,N_16808);
nor U18285 (N_18285,N_17460,N_17718);
and U18286 (N_18286,N_17565,N_17611);
or U18287 (N_18287,N_17697,N_17976);
nor U18288 (N_18288,N_16822,N_17479);
nand U18289 (N_18289,N_17216,N_17894);
nor U18290 (N_18290,N_17435,N_17034);
nand U18291 (N_18291,N_17023,N_17886);
or U18292 (N_18292,N_17257,N_17734);
nor U18293 (N_18293,N_17524,N_17963);
and U18294 (N_18294,N_17934,N_17823);
nor U18295 (N_18295,N_17111,N_16945);
nand U18296 (N_18296,N_17299,N_17854);
xor U18297 (N_18297,N_17822,N_17730);
xor U18298 (N_18298,N_17269,N_17919);
and U18299 (N_18299,N_17253,N_16861);
xor U18300 (N_18300,N_16762,N_17466);
and U18301 (N_18301,N_16798,N_17990);
xnor U18302 (N_18302,N_17373,N_17878);
nor U18303 (N_18303,N_17973,N_17068);
xor U18304 (N_18304,N_17519,N_16681);
or U18305 (N_18305,N_16569,N_16973);
and U18306 (N_18306,N_17089,N_17076);
nand U18307 (N_18307,N_17634,N_17508);
and U18308 (N_18308,N_16502,N_17226);
nand U18309 (N_18309,N_17841,N_17617);
nand U18310 (N_18310,N_17482,N_17817);
or U18311 (N_18311,N_16859,N_17073);
xnor U18312 (N_18312,N_17042,N_17234);
xor U18313 (N_18313,N_17992,N_16571);
or U18314 (N_18314,N_17326,N_17642);
nor U18315 (N_18315,N_17525,N_17774);
nor U18316 (N_18316,N_16893,N_17614);
nor U18317 (N_18317,N_17724,N_17391);
xor U18318 (N_18318,N_17262,N_17428);
nand U18319 (N_18319,N_17296,N_17285);
nor U18320 (N_18320,N_17087,N_16996);
nand U18321 (N_18321,N_16761,N_17750);
xor U18322 (N_18322,N_17415,N_17690);
xor U18323 (N_18323,N_16998,N_17862);
and U18324 (N_18324,N_17607,N_16802);
nand U18325 (N_18325,N_17318,N_16840);
or U18326 (N_18326,N_16746,N_17681);
and U18327 (N_18327,N_16528,N_17643);
nand U18328 (N_18328,N_16748,N_17300);
or U18329 (N_18329,N_17057,N_17079);
and U18330 (N_18330,N_17283,N_17352);
nand U18331 (N_18331,N_17457,N_17170);
or U18332 (N_18332,N_17462,N_17141);
nor U18333 (N_18333,N_16549,N_16758);
xor U18334 (N_18334,N_17037,N_16551);
xor U18335 (N_18335,N_17149,N_17182);
xnor U18336 (N_18336,N_16769,N_16948);
xor U18337 (N_18337,N_16977,N_17668);
nand U18338 (N_18338,N_17588,N_16568);
or U18339 (N_18339,N_17237,N_16740);
xnor U18340 (N_18340,N_16620,N_16799);
nor U18341 (N_18341,N_17905,N_16512);
nor U18342 (N_18342,N_16593,N_16652);
xnor U18343 (N_18343,N_17123,N_17645);
nor U18344 (N_18344,N_16958,N_17399);
or U18345 (N_18345,N_17953,N_17206);
xnor U18346 (N_18346,N_16951,N_17911);
nor U18347 (N_18347,N_16982,N_16667);
xor U18348 (N_18348,N_16812,N_16826);
xnor U18349 (N_18349,N_17378,N_17559);
nor U18350 (N_18350,N_17808,N_17065);
and U18351 (N_18351,N_16575,N_17012);
xnor U18352 (N_18352,N_16687,N_16716);
xnor U18353 (N_18353,N_17161,N_17382);
xor U18354 (N_18354,N_16735,N_17706);
xnor U18355 (N_18355,N_16975,N_17555);
nor U18356 (N_18356,N_16978,N_17873);
and U18357 (N_18357,N_16933,N_17736);
xor U18358 (N_18358,N_17474,N_17413);
or U18359 (N_18359,N_17993,N_16881);
and U18360 (N_18360,N_16705,N_16895);
or U18361 (N_18361,N_16515,N_16649);
and U18362 (N_18362,N_16531,N_17715);
xnor U18363 (N_18363,N_17902,N_16702);
nor U18364 (N_18364,N_17574,N_17883);
nand U18365 (N_18365,N_16777,N_16772);
xor U18366 (N_18366,N_17157,N_17031);
nand U18367 (N_18367,N_16708,N_17770);
or U18368 (N_18368,N_16979,N_17780);
and U18369 (N_18369,N_17907,N_17429);
and U18370 (N_18370,N_16654,N_17210);
and U18371 (N_18371,N_17307,N_17619);
nor U18372 (N_18372,N_16660,N_16874);
nor U18373 (N_18373,N_17701,N_17940);
xor U18374 (N_18374,N_17896,N_17692);
nand U18375 (N_18375,N_17887,N_17995);
and U18376 (N_18376,N_17334,N_16814);
nor U18377 (N_18377,N_17046,N_17268);
nand U18378 (N_18378,N_16642,N_17889);
xnor U18379 (N_18379,N_17937,N_17345);
xnor U18380 (N_18380,N_16651,N_16585);
nand U18381 (N_18381,N_17663,N_16673);
and U18382 (N_18382,N_16588,N_17848);
nor U18383 (N_18383,N_17672,N_17696);
nor U18384 (N_18384,N_17168,N_17782);
nand U18385 (N_18385,N_16930,N_17688);
or U18386 (N_18386,N_17133,N_17870);
and U18387 (N_18387,N_17545,N_17637);
xor U18388 (N_18388,N_17320,N_16760);
nand U18389 (N_18389,N_16843,N_16698);
xor U18390 (N_18390,N_17791,N_17654);
and U18391 (N_18391,N_16961,N_17989);
nor U18392 (N_18392,N_17638,N_16541);
or U18393 (N_18393,N_16912,N_17890);
or U18394 (N_18394,N_16525,N_17291);
or U18395 (N_18395,N_16796,N_16956);
xnor U18396 (N_18396,N_17728,N_16858);
nor U18397 (N_18397,N_17222,N_17610);
or U18398 (N_18398,N_17539,N_16886);
xnor U18399 (N_18399,N_16503,N_17422);
nand U18400 (N_18400,N_16671,N_16823);
or U18401 (N_18401,N_17839,N_17261);
nand U18402 (N_18402,N_17987,N_16914);
nor U18403 (N_18403,N_16594,N_16563);
or U18404 (N_18404,N_17594,N_16538);
and U18405 (N_18405,N_16547,N_17208);
nand U18406 (N_18406,N_17982,N_17019);
and U18407 (N_18407,N_17255,N_16957);
nand U18408 (N_18408,N_17192,N_16784);
nor U18409 (N_18409,N_17516,N_17092);
nor U18410 (N_18410,N_17779,N_16931);
xnor U18411 (N_18411,N_17860,N_16509);
xnor U18412 (N_18412,N_17747,N_17276);
nand U18413 (N_18413,N_17622,N_17126);
or U18414 (N_18414,N_17020,N_17760);
nand U18415 (N_18415,N_16597,N_17694);
or U18416 (N_18416,N_16781,N_17788);
nor U18417 (N_18417,N_17898,N_17749);
nand U18418 (N_18418,N_17631,N_17495);
nand U18419 (N_18419,N_16623,N_17152);
xor U18420 (N_18420,N_17929,N_17795);
nand U18421 (N_18421,N_17271,N_16750);
or U18422 (N_18422,N_17366,N_17032);
nand U18423 (N_18423,N_16785,N_17977);
xor U18424 (N_18424,N_17447,N_17892);
and U18425 (N_18425,N_16857,N_17473);
or U18426 (N_18426,N_17297,N_16567);
nand U18427 (N_18427,N_16792,N_17050);
xor U18428 (N_18428,N_17397,N_17483);
nand U18429 (N_18429,N_16521,N_16704);
xnor U18430 (N_18430,N_17150,N_16927);
nor U18431 (N_18431,N_16866,N_17687);
nand U18432 (N_18432,N_17173,N_16621);
nand U18433 (N_18433,N_16938,N_17875);
nand U18434 (N_18434,N_17063,N_17266);
nor U18435 (N_18435,N_16768,N_17102);
and U18436 (N_18436,N_16782,N_17164);
or U18437 (N_18437,N_17363,N_17188);
or U18438 (N_18438,N_16878,N_17254);
and U18439 (N_18439,N_16751,N_17693);
and U18440 (N_18440,N_16776,N_17790);
or U18441 (N_18441,N_16627,N_17713);
nor U18442 (N_18442,N_17142,N_17984);
or U18443 (N_18443,N_16789,N_16523);
nand U18444 (N_18444,N_16848,N_16697);
nor U18445 (N_18445,N_16561,N_17781);
nor U18446 (N_18446,N_17727,N_17756);
or U18447 (N_18447,N_17514,N_17538);
xor U18448 (N_18448,N_17659,N_16555);
and U18449 (N_18449,N_17436,N_17122);
xnor U18450 (N_18450,N_16606,N_16613);
nand U18451 (N_18451,N_17421,N_17238);
xor U18452 (N_18452,N_17971,N_17203);
and U18453 (N_18453,N_17499,N_16736);
and U18454 (N_18454,N_17636,N_17183);
nor U18455 (N_18455,N_16692,N_17433);
or U18456 (N_18456,N_17107,N_17569);
and U18457 (N_18457,N_17480,N_17088);
nor U18458 (N_18458,N_17517,N_17591);
nand U18459 (N_18459,N_17314,N_17628);
xnor U18460 (N_18460,N_17186,N_17322);
or U18461 (N_18461,N_17134,N_16905);
or U18462 (N_18462,N_17717,N_17375);
nand U18463 (N_18463,N_17942,N_17810);
nand U18464 (N_18464,N_17691,N_17265);
xnor U18465 (N_18465,N_16837,N_17721);
or U18466 (N_18466,N_17077,N_16636);
nand U18467 (N_18467,N_17787,N_17393);
and U18468 (N_18468,N_17580,N_16733);
or U18469 (N_18469,N_17361,N_17458);
and U18470 (N_18470,N_16879,N_17586);
nor U18471 (N_18471,N_17097,N_17923);
xnor U18472 (N_18472,N_17671,N_16647);
and U18473 (N_18473,N_17290,N_16663);
xnor U18474 (N_18474,N_17469,N_17994);
nor U18475 (N_18475,N_16548,N_17286);
xor U18476 (N_18476,N_17181,N_17389);
nor U18477 (N_18477,N_17816,N_17666);
and U18478 (N_18478,N_17308,N_17966);
or U18479 (N_18479,N_17187,N_16544);
nor U18480 (N_18480,N_17867,N_16519);
nor U18481 (N_18481,N_17476,N_17600);
or U18482 (N_18482,N_17075,N_16854);
nor U18483 (N_18483,N_16928,N_16724);
and U18484 (N_18484,N_17785,N_16747);
or U18485 (N_18485,N_16946,N_16986);
xor U18486 (N_18486,N_17678,N_16711);
nand U18487 (N_18487,N_17340,N_17394);
and U18488 (N_18488,N_17941,N_17893);
or U18489 (N_18489,N_17040,N_16764);
and U18490 (N_18490,N_16565,N_17251);
nand U18491 (N_18491,N_17484,N_17967);
xnor U18492 (N_18492,N_17932,N_17445);
or U18493 (N_18493,N_16535,N_17685);
or U18494 (N_18494,N_17988,N_16898);
xor U18495 (N_18495,N_16514,N_17424);
nor U18496 (N_18496,N_16941,N_17882);
xor U18497 (N_18497,N_16882,N_16511);
nand U18498 (N_18498,N_17362,N_16835);
nor U18499 (N_18499,N_17475,N_17640);
nand U18500 (N_18500,N_17794,N_16590);
xor U18501 (N_18501,N_16923,N_17627);
nand U18502 (N_18502,N_17100,N_17532);
nor U18503 (N_18503,N_17723,N_16646);
or U18504 (N_18504,N_17404,N_17109);
nand U18505 (N_18505,N_17918,N_17913);
nand U18506 (N_18506,N_16773,N_17431);
xor U18507 (N_18507,N_17365,N_16589);
or U18508 (N_18508,N_17609,N_17535);
and U18509 (N_18509,N_17761,N_17876);
or U18510 (N_18510,N_17544,N_17844);
or U18511 (N_18511,N_17863,N_17321);
xor U18512 (N_18512,N_17179,N_17125);
xor U18513 (N_18513,N_17895,N_16562);
nor U18514 (N_18514,N_16552,N_17763);
or U18515 (N_18515,N_17027,N_16505);
or U18516 (N_18516,N_17647,N_17180);
and U18517 (N_18517,N_17653,N_17354);
xor U18518 (N_18518,N_17537,N_17338);
xnor U18519 (N_18519,N_17401,N_16640);
nor U18520 (N_18520,N_17635,N_17985);
nand U18521 (N_18521,N_17776,N_16648);
or U18522 (N_18522,N_16939,N_17745);
nor U18523 (N_18523,N_16907,N_16581);
nor U18524 (N_18524,N_17127,N_17350);
nor U18525 (N_18525,N_17825,N_16987);
and U18526 (N_18526,N_16976,N_17374);
nand U18527 (N_18527,N_16807,N_17793);
or U18528 (N_18528,N_17112,N_17677);
nand U18529 (N_18529,N_16953,N_17218);
or U18530 (N_18530,N_17005,N_16730);
nand U18531 (N_18531,N_16887,N_16794);
or U18532 (N_18532,N_16574,N_16713);
xor U18533 (N_18533,N_16901,N_16779);
and U18534 (N_18534,N_17030,N_17249);
or U18535 (N_18535,N_17096,N_17486);
and U18536 (N_18536,N_17330,N_16989);
xnor U18537 (N_18537,N_17390,N_17128);
or U18538 (N_18538,N_16518,N_16775);
xor U18539 (N_18539,N_17999,N_17070);
xnor U18540 (N_18540,N_16897,N_17202);
nor U18541 (N_18541,N_17757,N_17145);
nand U18542 (N_18542,N_17589,N_17408);
xor U18543 (N_18543,N_16714,N_17006);
or U18544 (N_18544,N_16992,N_16818);
xnor U18545 (N_18545,N_16737,N_17316);
xnor U18546 (N_18546,N_16800,N_17662);
and U18547 (N_18547,N_16572,N_17773);
and U18548 (N_18548,N_16770,N_16644);
nor U18549 (N_18549,N_16564,N_16550);
or U18550 (N_18550,N_17748,N_16917);
nand U18551 (N_18551,N_16790,N_16919);
nor U18552 (N_18552,N_17434,N_17016);
and U18553 (N_18553,N_17991,N_17384);
nand U18554 (N_18554,N_17501,N_17972);
or U18555 (N_18555,N_16638,N_16662);
nor U18556 (N_18556,N_17531,N_16566);
and U18557 (N_18557,N_16783,N_17159);
nand U18558 (N_18558,N_17705,N_17346);
nor U18559 (N_18559,N_17383,N_17807);
nand U18560 (N_18560,N_17277,N_16533);
nor U18561 (N_18561,N_17481,N_17616);
or U18562 (N_18562,N_17022,N_16828);
xnor U18563 (N_18563,N_17731,N_17552);
xnor U18564 (N_18564,N_17193,N_17601);
or U18565 (N_18565,N_17562,N_16849);
and U18566 (N_18566,N_16959,N_17137);
and U18567 (N_18567,N_17751,N_17066);
or U18568 (N_18568,N_17294,N_17560);
nand U18569 (N_18569,N_17775,N_16851);
nand U18570 (N_18570,N_17459,N_17646);
nor U18571 (N_18571,N_16839,N_17680);
or U18572 (N_18572,N_17974,N_17827);
or U18573 (N_18573,N_17405,N_17871);
nand U18574 (N_18574,N_16680,N_16824);
xnor U18575 (N_18575,N_17759,N_16524);
xor U18576 (N_18576,N_16780,N_16611);
nor U18577 (N_18577,N_17901,N_16582);
nor U18578 (N_18578,N_17368,N_17282);
xnor U18579 (N_18579,N_17665,N_16892);
and U18580 (N_18580,N_16968,N_17392);
nand U18581 (N_18581,N_17439,N_17140);
nand U18582 (N_18582,N_16852,N_17726);
or U18583 (N_18583,N_17241,N_17178);
xor U18584 (N_18584,N_17623,N_17850);
xor U18585 (N_18585,N_16729,N_17506);
xor U18586 (N_18586,N_17840,N_17135);
nor U18587 (N_18587,N_16699,N_17248);
xor U18588 (N_18588,N_17596,N_16608);
nand U18589 (N_18589,N_17067,N_17278);
nor U18590 (N_18590,N_16570,N_17306);
xor U18591 (N_18591,N_17098,N_17333);
xnor U18592 (N_18592,N_16804,N_17900);
xor U18593 (N_18593,N_17132,N_17674);
and U18594 (N_18594,N_17343,N_16815);
nand U18595 (N_18595,N_17964,N_17275);
and U18596 (N_18596,N_17093,N_17879);
nor U18597 (N_18597,N_17225,N_17423);
nor U18598 (N_18598,N_16721,N_17884);
and U18599 (N_18599,N_17959,N_17119);
nor U18600 (N_18600,N_17058,N_17783);
and U18601 (N_18601,N_17372,N_17658);
xnor U18602 (N_18602,N_16831,N_17337);
nand U18603 (N_18603,N_16820,N_17831);
xnor U18604 (N_18604,N_16841,N_16693);
and U18605 (N_18605,N_16609,N_16915);
xor U18606 (N_18606,N_17353,N_17120);
or U18607 (N_18607,N_17815,N_17582);
or U18608 (N_18608,N_17625,N_17669);
nor U18609 (N_18609,N_17110,N_17792);
xor U18610 (N_18610,N_17909,N_17449);
nand U18611 (N_18611,N_17814,N_17881);
and U18612 (N_18612,N_17175,N_16513);
or U18613 (N_18613,N_16904,N_17915);
xnor U18614 (N_18614,N_17920,N_17936);
and U18615 (N_18615,N_16605,N_17513);
xnor U18616 (N_18616,N_17471,N_17025);
nor U18617 (N_18617,N_17561,N_17980);
nor U18618 (N_18618,N_17244,N_17868);
nand U18619 (N_18619,N_17051,N_17494);
xor U18620 (N_18620,N_17242,N_17648);
or U18621 (N_18621,N_17114,N_17124);
nand U18622 (N_18622,N_17414,N_17038);
and U18623 (N_18623,N_17105,N_17490);
nand U18624 (N_18624,N_16685,N_16599);
nor U18625 (N_18625,N_16869,N_17811);
and U18626 (N_18626,N_17344,N_16727);
or U18627 (N_18627,N_16980,N_17117);
and U18628 (N_18628,N_17010,N_17803);
or U18629 (N_18629,N_17510,N_17768);
and U18630 (N_18630,N_17082,N_16971);
and U18631 (N_18631,N_17304,N_16955);
nand U18632 (N_18632,N_16624,N_17444);
xnor U18633 (N_18633,N_17679,N_17086);
xnor U18634 (N_18634,N_17015,N_17190);
and U18635 (N_18635,N_17673,N_17549);
nor U18636 (N_18636,N_17921,N_16684);
nand U18637 (N_18637,N_17195,N_16619);
and U18638 (N_18638,N_17407,N_17309);
and U18639 (N_18639,N_17310,N_17852);
nand U18640 (N_18640,N_17845,N_17438);
or U18641 (N_18641,N_16926,N_16622);
xor U18642 (N_18642,N_17301,N_16598);
nand U18643 (N_18643,N_16691,N_16771);
nand U18644 (N_18644,N_17380,N_17548);
or U18645 (N_18645,N_16632,N_17849);
and U18646 (N_18646,N_16583,N_16900);
and U18647 (N_18647,N_17576,N_17981);
nor U18648 (N_18648,N_17289,N_17939);
or U18649 (N_18649,N_16896,N_17961);
xnor U18650 (N_18650,N_16788,N_16527);
nand U18651 (N_18651,N_16864,N_17847);
or U18652 (N_18652,N_17388,N_16543);
xnor U18653 (N_18653,N_17174,N_16855);
nand U18654 (N_18654,N_17583,N_16868);
nand U18655 (N_18655,N_17091,N_17013);
xor U18656 (N_18656,N_17224,N_17211);
xnor U18657 (N_18657,N_17906,N_16795);
nor U18658 (N_18658,N_17754,N_17716);
nor U18659 (N_18659,N_17935,N_16522);
xnor U18660 (N_18660,N_17866,N_17778);
nand U18661 (N_18661,N_17264,N_17821);
and U18662 (N_18662,N_16870,N_16759);
nand U18663 (N_18663,N_17504,N_17348);
nand U18664 (N_18664,N_17396,N_17573);
xnor U18665 (N_18665,N_16838,N_17028);
xor U18666 (N_18666,N_17033,N_17832);
nor U18667 (N_18667,N_17533,N_16580);
or U18668 (N_18668,N_16935,N_17214);
or U18669 (N_18669,N_17541,N_16754);
nand U18670 (N_18670,N_17916,N_17587);
nand U18671 (N_18671,N_17801,N_17336);
or U18672 (N_18672,N_17412,N_16985);
and U18673 (N_18673,N_17742,N_17842);
nor U18674 (N_18674,N_17629,N_16873);
nand U18675 (N_18675,N_17575,N_17732);
or U18676 (N_18676,N_17367,N_17041);
nor U18677 (N_18677,N_17347,N_17489);
and U18678 (N_18678,N_17809,N_17944);
nand U18679 (N_18679,N_17858,N_17897);
nand U18680 (N_18680,N_17196,N_17463);
or U18681 (N_18681,N_17996,N_17564);
xor U18682 (N_18682,N_17503,N_16600);
nor U18683 (N_18683,N_17021,N_17798);
nor U18684 (N_18684,N_17927,N_17805);
nor U18685 (N_18685,N_17044,N_17485);
nand U18686 (N_18686,N_16834,N_17553);
xor U18687 (N_18687,N_17477,N_17446);
or U18688 (N_18688,N_16587,N_17074);
or U18689 (N_18689,N_17664,N_17652);
and U18690 (N_18690,N_17387,N_17834);
or U18691 (N_18691,N_17217,N_17954);
or U18692 (N_18692,N_17965,N_17502);
xnor U18693 (N_18693,N_17298,N_16558);
xor U18694 (N_18694,N_17698,N_17528);
nor U18695 (N_18695,N_16625,N_17229);
and U18696 (N_18696,N_17644,N_17737);
and U18697 (N_18697,N_16871,N_17281);
nor U18698 (N_18698,N_17563,N_17910);
and U18699 (N_18699,N_16888,N_17707);
nand U18700 (N_18700,N_17154,N_16542);
nor U18701 (N_18701,N_17035,N_16876);
xor U18702 (N_18702,N_16970,N_16715);
nand U18703 (N_18703,N_16803,N_17922);
nand U18704 (N_18704,N_16701,N_16679);
nand U18705 (N_18705,N_17047,N_17014);
and U18706 (N_18706,N_17454,N_17274);
or U18707 (N_18707,N_16891,N_16586);
or U18708 (N_18708,N_16995,N_16659);
or U18709 (N_18709,N_16974,N_16672);
xor U18710 (N_18710,N_17131,N_17172);
xnor U18711 (N_18711,N_17008,N_17943);
nand U18712 (N_18712,N_17227,N_17926);
nand U18713 (N_18713,N_17267,N_16706);
nor U18714 (N_18714,N_17043,N_17213);
or U18715 (N_18715,N_17280,N_16984);
nor U18716 (N_18716,N_17604,N_16641);
xor U18717 (N_18717,N_17478,N_16911);
xor U18718 (N_18718,N_17650,N_17007);
and U18719 (N_18719,N_17328,N_17081);
and U18720 (N_18720,N_16738,N_17853);
nor U18721 (N_18721,N_16829,N_16658);
xor U18722 (N_18722,N_16836,N_17930);
or U18723 (N_18723,N_16937,N_17529);
and U18724 (N_18724,N_17908,N_17874);
or U18725 (N_18725,N_17608,N_16703);
or U18726 (N_18726,N_17515,N_17542);
nand U18727 (N_18727,N_17667,N_17526);
or U18728 (N_18728,N_16501,N_17593);
and U18729 (N_18729,N_17061,N_17472);
nor U18730 (N_18730,N_17521,N_17729);
nor U18731 (N_18731,N_16925,N_17684);
or U18732 (N_18732,N_17420,N_17755);
or U18733 (N_18733,N_17059,N_16753);
nor U18734 (N_18734,N_17358,N_17406);
and U18735 (N_18735,N_17256,N_16643);
nand U18736 (N_18736,N_17865,N_17386);
nor U18737 (N_18737,N_16633,N_16749);
or U18738 (N_18738,N_17487,N_17341);
nor U18739 (N_18739,N_17551,N_16540);
xnor U18740 (N_18740,N_17917,N_17385);
nor U18741 (N_18741,N_17220,N_16903);
xor U18742 (N_18742,N_17758,N_16755);
and U18743 (N_18743,N_16539,N_16553);
or U18744 (N_18744,N_16793,N_16739);
nor U18745 (N_18745,N_17240,N_16596);
or U18746 (N_18746,N_17670,N_17970);
xnor U18747 (N_18747,N_16867,N_17410);
nor U18748 (N_18748,N_17630,N_17342);
nand U18749 (N_18749,N_17824,N_17851);
or U18750 (N_18750,N_16718,N_16745);
and U18751 (N_18751,N_17042,N_16844);
nand U18752 (N_18752,N_17123,N_17589);
and U18753 (N_18753,N_16789,N_17609);
or U18754 (N_18754,N_17005,N_17765);
nor U18755 (N_18755,N_17125,N_16692);
and U18756 (N_18756,N_16826,N_16668);
xor U18757 (N_18757,N_17045,N_16899);
and U18758 (N_18758,N_17669,N_17924);
nor U18759 (N_18759,N_16502,N_17863);
nand U18760 (N_18760,N_17248,N_17257);
nor U18761 (N_18761,N_17133,N_17144);
and U18762 (N_18762,N_16624,N_17234);
and U18763 (N_18763,N_17287,N_16816);
xnor U18764 (N_18764,N_16651,N_17981);
nand U18765 (N_18765,N_16812,N_16716);
nand U18766 (N_18766,N_17092,N_16964);
xnor U18767 (N_18767,N_17229,N_17809);
nand U18768 (N_18768,N_17217,N_17022);
or U18769 (N_18769,N_17746,N_16672);
xnor U18770 (N_18770,N_17832,N_17609);
nor U18771 (N_18771,N_16782,N_16962);
or U18772 (N_18772,N_17189,N_17945);
or U18773 (N_18773,N_16894,N_16886);
and U18774 (N_18774,N_17587,N_17149);
nor U18775 (N_18775,N_17621,N_17807);
nor U18776 (N_18776,N_17143,N_16984);
or U18777 (N_18777,N_17322,N_17827);
or U18778 (N_18778,N_17935,N_17732);
nand U18779 (N_18779,N_17230,N_16822);
nor U18780 (N_18780,N_17673,N_17059);
nor U18781 (N_18781,N_17814,N_16724);
or U18782 (N_18782,N_16926,N_17069);
nand U18783 (N_18783,N_17806,N_16789);
nor U18784 (N_18784,N_16725,N_17551);
nor U18785 (N_18785,N_17432,N_17764);
and U18786 (N_18786,N_17309,N_17862);
xor U18787 (N_18787,N_17203,N_17376);
and U18788 (N_18788,N_16573,N_16518);
nor U18789 (N_18789,N_16530,N_17735);
nand U18790 (N_18790,N_17920,N_17558);
xnor U18791 (N_18791,N_16588,N_16624);
or U18792 (N_18792,N_17739,N_17332);
nand U18793 (N_18793,N_17764,N_17690);
nor U18794 (N_18794,N_17709,N_16656);
and U18795 (N_18795,N_17833,N_16638);
or U18796 (N_18796,N_16634,N_16530);
or U18797 (N_18797,N_17426,N_16979);
xnor U18798 (N_18798,N_17424,N_17710);
nand U18799 (N_18799,N_16593,N_16600);
nor U18800 (N_18800,N_17205,N_16903);
or U18801 (N_18801,N_17021,N_16869);
or U18802 (N_18802,N_17115,N_16762);
xor U18803 (N_18803,N_17854,N_17830);
and U18804 (N_18804,N_16511,N_17969);
xor U18805 (N_18805,N_17319,N_17165);
xnor U18806 (N_18806,N_17814,N_17399);
nor U18807 (N_18807,N_17835,N_17284);
nor U18808 (N_18808,N_17574,N_17067);
nor U18809 (N_18809,N_16863,N_17351);
nor U18810 (N_18810,N_16797,N_17293);
xnor U18811 (N_18811,N_17565,N_16769);
nor U18812 (N_18812,N_16868,N_17663);
and U18813 (N_18813,N_17636,N_16905);
or U18814 (N_18814,N_17831,N_16897);
nor U18815 (N_18815,N_16548,N_17822);
or U18816 (N_18816,N_17022,N_17255);
or U18817 (N_18817,N_17907,N_17135);
xor U18818 (N_18818,N_17309,N_17471);
and U18819 (N_18819,N_17523,N_17883);
xnor U18820 (N_18820,N_17787,N_16745);
xnor U18821 (N_18821,N_16635,N_16678);
or U18822 (N_18822,N_17017,N_17947);
nor U18823 (N_18823,N_16589,N_17776);
and U18824 (N_18824,N_16753,N_16848);
and U18825 (N_18825,N_16862,N_16992);
xnor U18826 (N_18826,N_16686,N_17380);
xnor U18827 (N_18827,N_17689,N_17375);
nor U18828 (N_18828,N_16758,N_17541);
xnor U18829 (N_18829,N_17400,N_17145);
or U18830 (N_18830,N_16531,N_16707);
nand U18831 (N_18831,N_17078,N_16878);
nor U18832 (N_18832,N_16704,N_17307);
and U18833 (N_18833,N_16527,N_17234);
nor U18834 (N_18834,N_17202,N_17614);
nand U18835 (N_18835,N_16551,N_17952);
xor U18836 (N_18836,N_17089,N_16859);
nor U18837 (N_18837,N_16554,N_16987);
or U18838 (N_18838,N_17536,N_17727);
xor U18839 (N_18839,N_16619,N_17111);
nand U18840 (N_18840,N_17583,N_17709);
nor U18841 (N_18841,N_17722,N_17810);
xor U18842 (N_18842,N_17611,N_17431);
xnor U18843 (N_18843,N_16741,N_16613);
xor U18844 (N_18844,N_16677,N_17332);
nand U18845 (N_18845,N_16658,N_16929);
or U18846 (N_18846,N_16621,N_16755);
nand U18847 (N_18847,N_17551,N_17020);
nand U18848 (N_18848,N_16574,N_17193);
nand U18849 (N_18849,N_17292,N_17055);
xor U18850 (N_18850,N_17977,N_17859);
nor U18851 (N_18851,N_17279,N_17211);
nand U18852 (N_18852,N_17998,N_17764);
and U18853 (N_18853,N_17105,N_17748);
and U18854 (N_18854,N_17171,N_16868);
and U18855 (N_18855,N_16953,N_16902);
nand U18856 (N_18856,N_17106,N_17141);
and U18857 (N_18857,N_17783,N_17048);
xnor U18858 (N_18858,N_17106,N_17662);
nand U18859 (N_18859,N_17059,N_16507);
or U18860 (N_18860,N_17463,N_16503);
and U18861 (N_18861,N_17802,N_16759);
xnor U18862 (N_18862,N_17241,N_16658);
and U18863 (N_18863,N_16637,N_16690);
and U18864 (N_18864,N_17121,N_17442);
and U18865 (N_18865,N_16604,N_17497);
and U18866 (N_18866,N_17134,N_16593);
nand U18867 (N_18867,N_17345,N_17044);
and U18868 (N_18868,N_17825,N_17414);
and U18869 (N_18869,N_17555,N_16923);
xnor U18870 (N_18870,N_17638,N_17879);
nor U18871 (N_18871,N_17908,N_17976);
or U18872 (N_18872,N_17196,N_17026);
nor U18873 (N_18873,N_16588,N_17092);
nor U18874 (N_18874,N_17252,N_16883);
and U18875 (N_18875,N_17743,N_17197);
nor U18876 (N_18876,N_17213,N_16678);
or U18877 (N_18877,N_17682,N_16749);
and U18878 (N_18878,N_17674,N_17924);
or U18879 (N_18879,N_17017,N_16788);
or U18880 (N_18880,N_16529,N_16870);
and U18881 (N_18881,N_16740,N_16627);
nand U18882 (N_18882,N_16516,N_17564);
xnor U18883 (N_18883,N_17854,N_16528);
or U18884 (N_18884,N_17102,N_17988);
and U18885 (N_18885,N_17217,N_17613);
or U18886 (N_18886,N_17511,N_16835);
xnor U18887 (N_18887,N_17288,N_17430);
nand U18888 (N_18888,N_16501,N_16889);
nand U18889 (N_18889,N_16731,N_17032);
xnor U18890 (N_18890,N_17378,N_17414);
and U18891 (N_18891,N_17494,N_17783);
nand U18892 (N_18892,N_17247,N_17398);
xnor U18893 (N_18893,N_17071,N_17312);
nand U18894 (N_18894,N_17988,N_17843);
or U18895 (N_18895,N_17161,N_17179);
or U18896 (N_18896,N_16634,N_16569);
nand U18897 (N_18897,N_16898,N_17360);
nor U18898 (N_18898,N_17273,N_17339);
and U18899 (N_18899,N_16512,N_17891);
and U18900 (N_18900,N_16777,N_16838);
and U18901 (N_18901,N_17133,N_17865);
nor U18902 (N_18902,N_17449,N_17827);
or U18903 (N_18903,N_16876,N_16766);
nor U18904 (N_18904,N_17023,N_17013);
nor U18905 (N_18905,N_17689,N_17861);
nand U18906 (N_18906,N_17950,N_17523);
nor U18907 (N_18907,N_17566,N_16815);
and U18908 (N_18908,N_17454,N_17958);
and U18909 (N_18909,N_17116,N_16572);
and U18910 (N_18910,N_16642,N_17119);
nand U18911 (N_18911,N_16778,N_17888);
nor U18912 (N_18912,N_17848,N_17143);
nor U18913 (N_18913,N_17232,N_17302);
nor U18914 (N_18914,N_17634,N_17697);
and U18915 (N_18915,N_17625,N_17573);
nor U18916 (N_18916,N_16794,N_16911);
or U18917 (N_18917,N_16936,N_17090);
xor U18918 (N_18918,N_17098,N_16716);
xnor U18919 (N_18919,N_17122,N_16961);
and U18920 (N_18920,N_17456,N_17945);
xnor U18921 (N_18921,N_16905,N_17284);
nand U18922 (N_18922,N_16988,N_16583);
nor U18923 (N_18923,N_17832,N_17855);
xnor U18924 (N_18924,N_17528,N_17527);
nand U18925 (N_18925,N_16620,N_16885);
nor U18926 (N_18926,N_16628,N_17286);
nand U18927 (N_18927,N_17172,N_17540);
nand U18928 (N_18928,N_17080,N_17857);
xnor U18929 (N_18929,N_16818,N_17697);
nor U18930 (N_18930,N_17925,N_17039);
and U18931 (N_18931,N_17406,N_17942);
xor U18932 (N_18932,N_17058,N_17223);
or U18933 (N_18933,N_17497,N_17746);
nor U18934 (N_18934,N_17021,N_16691);
xnor U18935 (N_18935,N_17087,N_16692);
xnor U18936 (N_18936,N_16911,N_17570);
nand U18937 (N_18937,N_16628,N_17498);
nor U18938 (N_18938,N_17484,N_16770);
xnor U18939 (N_18939,N_17222,N_16659);
xnor U18940 (N_18940,N_17972,N_17159);
or U18941 (N_18941,N_17468,N_17584);
xnor U18942 (N_18942,N_17131,N_16626);
or U18943 (N_18943,N_16754,N_17124);
and U18944 (N_18944,N_17830,N_17639);
xor U18945 (N_18945,N_17633,N_17868);
and U18946 (N_18946,N_17867,N_17480);
and U18947 (N_18947,N_16649,N_17686);
nor U18948 (N_18948,N_17601,N_17238);
nand U18949 (N_18949,N_17991,N_17005);
and U18950 (N_18950,N_17728,N_17295);
nand U18951 (N_18951,N_16711,N_17478);
nor U18952 (N_18952,N_16518,N_16990);
nand U18953 (N_18953,N_16635,N_17134);
or U18954 (N_18954,N_17800,N_16598);
nor U18955 (N_18955,N_16659,N_16690);
xor U18956 (N_18956,N_17139,N_16710);
or U18957 (N_18957,N_17250,N_17777);
nand U18958 (N_18958,N_16985,N_17223);
xnor U18959 (N_18959,N_17204,N_17750);
xor U18960 (N_18960,N_16755,N_17330);
or U18961 (N_18961,N_17037,N_17104);
xnor U18962 (N_18962,N_16522,N_17726);
or U18963 (N_18963,N_17301,N_16872);
nor U18964 (N_18964,N_16658,N_16511);
xor U18965 (N_18965,N_17779,N_17556);
nor U18966 (N_18966,N_16834,N_17607);
xor U18967 (N_18967,N_16932,N_17165);
or U18968 (N_18968,N_17720,N_16989);
or U18969 (N_18969,N_16814,N_16856);
and U18970 (N_18970,N_16639,N_16645);
or U18971 (N_18971,N_16861,N_17299);
nor U18972 (N_18972,N_17174,N_17440);
nand U18973 (N_18973,N_16861,N_17466);
nand U18974 (N_18974,N_16753,N_17607);
nor U18975 (N_18975,N_17579,N_16853);
nand U18976 (N_18976,N_17759,N_17354);
and U18977 (N_18977,N_17201,N_17851);
and U18978 (N_18978,N_17095,N_17749);
xor U18979 (N_18979,N_17080,N_17099);
and U18980 (N_18980,N_17384,N_17649);
or U18981 (N_18981,N_17630,N_17042);
or U18982 (N_18982,N_17376,N_16634);
xor U18983 (N_18983,N_16977,N_16950);
and U18984 (N_18984,N_16964,N_17984);
and U18985 (N_18985,N_17611,N_16658);
and U18986 (N_18986,N_17447,N_17937);
nand U18987 (N_18987,N_17881,N_17414);
nor U18988 (N_18988,N_17480,N_17695);
nor U18989 (N_18989,N_17614,N_16940);
and U18990 (N_18990,N_17610,N_17715);
nand U18991 (N_18991,N_17660,N_17389);
or U18992 (N_18992,N_17344,N_16600);
nor U18993 (N_18993,N_17783,N_17789);
and U18994 (N_18994,N_17637,N_17643);
nand U18995 (N_18995,N_17832,N_17664);
or U18996 (N_18996,N_17394,N_17862);
or U18997 (N_18997,N_17098,N_17087);
xor U18998 (N_18998,N_17118,N_16819);
nor U18999 (N_18999,N_16998,N_17160);
xnor U19000 (N_19000,N_17848,N_17577);
xnor U19001 (N_19001,N_17507,N_16780);
or U19002 (N_19002,N_17545,N_17823);
or U19003 (N_19003,N_16572,N_17989);
and U19004 (N_19004,N_16794,N_17166);
xnor U19005 (N_19005,N_17769,N_17190);
nor U19006 (N_19006,N_16595,N_17213);
and U19007 (N_19007,N_17779,N_17480);
nand U19008 (N_19008,N_17700,N_16556);
nand U19009 (N_19009,N_17385,N_16909);
or U19010 (N_19010,N_17148,N_17640);
or U19011 (N_19011,N_17896,N_16643);
nor U19012 (N_19012,N_17352,N_16597);
xor U19013 (N_19013,N_16619,N_17378);
nand U19014 (N_19014,N_16713,N_17321);
nor U19015 (N_19015,N_16923,N_16688);
nor U19016 (N_19016,N_17962,N_17716);
and U19017 (N_19017,N_16588,N_16868);
and U19018 (N_19018,N_17934,N_17121);
or U19019 (N_19019,N_17160,N_16665);
and U19020 (N_19020,N_16914,N_16617);
xor U19021 (N_19021,N_17000,N_16746);
nor U19022 (N_19022,N_16603,N_16576);
and U19023 (N_19023,N_17008,N_16522);
or U19024 (N_19024,N_17464,N_17583);
nor U19025 (N_19025,N_16873,N_17823);
nor U19026 (N_19026,N_16560,N_16682);
nor U19027 (N_19027,N_17606,N_17933);
or U19028 (N_19028,N_16848,N_17579);
and U19029 (N_19029,N_17610,N_17594);
or U19030 (N_19030,N_17209,N_17798);
or U19031 (N_19031,N_16635,N_17730);
nand U19032 (N_19032,N_17665,N_17476);
and U19033 (N_19033,N_17414,N_17972);
xnor U19034 (N_19034,N_17665,N_16673);
nor U19035 (N_19035,N_16746,N_16716);
nor U19036 (N_19036,N_17431,N_17148);
nand U19037 (N_19037,N_16524,N_16952);
and U19038 (N_19038,N_16723,N_16706);
or U19039 (N_19039,N_17081,N_17298);
xnor U19040 (N_19040,N_16602,N_17820);
nand U19041 (N_19041,N_16603,N_17957);
nand U19042 (N_19042,N_17683,N_16626);
nor U19043 (N_19043,N_17468,N_17372);
or U19044 (N_19044,N_17005,N_17570);
and U19045 (N_19045,N_17633,N_16894);
and U19046 (N_19046,N_16606,N_16638);
nor U19047 (N_19047,N_17420,N_17178);
or U19048 (N_19048,N_17294,N_17220);
nand U19049 (N_19049,N_17223,N_17754);
or U19050 (N_19050,N_16786,N_17853);
nand U19051 (N_19051,N_17516,N_17322);
or U19052 (N_19052,N_17530,N_16691);
or U19053 (N_19053,N_16957,N_16718);
xor U19054 (N_19054,N_17504,N_17622);
and U19055 (N_19055,N_17775,N_16528);
xor U19056 (N_19056,N_17523,N_17391);
xor U19057 (N_19057,N_17755,N_17463);
or U19058 (N_19058,N_17089,N_16681);
and U19059 (N_19059,N_17683,N_16870);
or U19060 (N_19060,N_17080,N_17693);
xnor U19061 (N_19061,N_16744,N_16976);
and U19062 (N_19062,N_17653,N_16654);
nand U19063 (N_19063,N_16631,N_16990);
and U19064 (N_19064,N_17672,N_16755);
xnor U19065 (N_19065,N_16835,N_17846);
and U19066 (N_19066,N_17095,N_17561);
xnor U19067 (N_19067,N_17595,N_17582);
nand U19068 (N_19068,N_17615,N_17805);
or U19069 (N_19069,N_17911,N_16874);
nor U19070 (N_19070,N_17437,N_17310);
nand U19071 (N_19071,N_17463,N_17864);
or U19072 (N_19072,N_17375,N_16655);
xnor U19073 (N_19073,N_17075,N_16753);
or U19074 (N_19074,N_17018,N_16738);
or U19075 (N_19075,N_17694,N_16799);
and U19076 (N_19076,N_16964,N_17306);
nor U19077 (N_19077,N_17321,N_17645);
nor U19078 (N_19078,N_17032,N_17237);
xor U19079 (N_19079,N_17556,N_16701);
nand U19080 (N_19080,N_17012,N_17712);
nand U19081 (N_19081,N_16825,N_16656);
nor U19082 (N_19082,N_17641,N_17558);
and U19083 (N_19083,N_17562,N_16700);
nor U19084 (N_19084,N_17099,N_16824);
nor U19085 (N_19085,N_16606,N_17766);
and U19086 (N_19086,N_16658,N_17216);
nor U19087 (N_19087,N_17068,N_17217);
or U19088 (N_19088,N_16966,N_17920);
or U19089 (N_19089,N_17592,N_16798);
xor U19090 (N_19090,N_17514,N_16782);
nor U19091 (N_19091,N_16695,N_16623);
nor U19092 (N_19092,N_17491,N_17036);
nor U19093 (N_19093,N_17800,N_17521);
nor U19094 (N_19094,N_17989,N_17890);
nand U19095 (N_19095,N_17484,N_16728);
and U19096 (N_19096,N_17933,N_17712);
and U19097 (N_19097,N_17668,N_16528);
nor U19098 (N_19098,N_16990,N_17948);
nand U19099 (N_19099,N_17003,N_17155);
nand U19100 (N_19100,N_17154,N_17122);
or U19101 (N_19101,N_17261,N_17521);
xnor U19102 (N_19102,N_16983,N_17504);
and U19103 (N_19103,N_17839,N_17582);
and U19104 (N_19104,N_16686,N_17843);
or U19105 (N_19105,N_17618,N_17951);
or U19106 (N_19106,N_16873,N_17084);
xor U19107 (N_19107,N_17865,N_16541);
nand U19108 (N_19108,N_16699,N_16549);
nor U19109 (N_19109,N_17914,N_17493);
xnor U19110 (N_19110,N_17025,N_17130);
or U19111 (N_19111,N_17911,N_17360);
nand U19112 (N_19112,N_17780,N_17828);
nor U19113 (N_19113,N_16814,N_17642);
nand U19114 (N_19114,N_17289,N_17300);
xnor U19115 (N_19115,N_17429,N_16991);
nor U19116 (N_19116,N_16688,N_17053);
or U19117 (N_19117,N_17133,N_17466);
or U19118 (N_19118,N_16819,N_17069);
nand U19119 (N_19119,N_17258,N_17647);
or U19120 (N_19120,N_17502,N_17046);
nand U19121 (N_19121,N_16536,N_17425);
or U19122 (N_19122,N_16773,N_17694);
xor U19123 (N_19123,N_17057,N_17686);
nor U19124 (N_19124,N_17879,N_17138);
nand U19125 (N_19125,N_17062,N_17855);
nor U19126 (N_19126,N_17847,N_17520);
or U19127 (N_19127,N_16742,N_17163);
nor U19128 (N_19128,N_17506,N_17695);
or U19129 (N_19129,N_16918,N_16792);
or U19130 (N_19130,N_17967,N_17749);
and U19131 (N_19131,N_17815,N_17712);
nand U19132 (N_19132,N_17922,N_17448);
and U19133 (N_19133,N_17082,N_16601);
nor U19134 (N_19134,N_17063,N_17156);
and U19135 (N_19135,N_17080,N_16896);
nor U19136 (N_19136,N_16543,N_17396);
nand U19137 (N_19137,N_17813,N_17519);
or U19138 (N_19138,N_17650,N_17515);
and U19139 (N_19139,N_16773,N_17891);
xnor U19140 (N_19140,N_17270,N_17076);
xnor U19141 (N_19141,N_17574,N_17460);
or U19142 (N_19142,N_17294,N_17513);
or U19143 (N_19143,N_16928,N_17363);
or U19144 (N_19144,N_17624,N_16840);
xnor U19145 (N_19145,N_17239,N_17138);
and U19146 (N_19146,N_17547,N_16512);
and U19147 (N_19147,N_17127,N_17440);
nand U19148 (N_19148,N_17407,N_16980);
xor U19149 (N_19149,N_17876,N_16961);
xor U19150 (N_19150,N_17137,N_16586);
nand U19151 (N_19151,N_17274,N_17076);
or U19152 (N_19152,N_17995,N_16833);
xnor U19153 (N_19153,N_17891,N_16899);
xnor U19154 (N_19154,N_17755,N_17195);
nand U19155 (N_19155,N_17178,N_16793);
nor U19156 (N_19156,N_17641,N_17880);
nand U19157 (N_19157,N_17229,N_17489);
or U19158 (N_19158,N_17120,N_16665);
nor U19159 (N_19159,N_16795,N_17119);
or U19160 (N_19160,N_17224,N_17088);
and U19161 (N_19161,N_17055,N_17646);
and U19162 (N_19162,N_17817,N_16859);
and U19163 (N_19163,N_17378,N_16688);
xor U19164 (N_19164,N_17074,N_17990);
xor U19165 (N_19165,N_17494,N_17870);
and U19166 (N_19166,N_16699,N_17650);
nand U19167 (N_19167,N_17163,N_16512);
and U19168 (N_19168,N_17868,N_16598);
and U19169 (N_19169,N_16920,N_16654);
and U19170 (N_19170,N_17783,N_16591);
nor U19171 (N_19171,N_17563,N_17527);
or U19172 (N_19172,N_17079,N_17991);
or U19173 (N_19173,N_17642,N_16612);
nand U19174 (N_19174,N_16561,N_16718);
nor U19175 (N_19175,N_17969,N_17614);
or U19176 (N_19176,N_16895,N_17710);
nand U19177 (N_19177,N_17711,N_16849);
xnor U19178 (N_19178,N_17914,N_17531);
or U19179 (N_19179,N_17508,N_17696);
and U19180 (N_19180,N_17178,N_17072);
nand U19181 (N_19181,N_17634,N_16597);
nor U19182 (N_19182,N_17884,N_16810);
nand U19183 (N_19183,N_16838,N_17595);
xor U19184 (N_19184,N_16558,N_16814);
or U19185 (N_19185,N_16781,N_17626);
nand U19186 (N_19186,N_16947,N_16743);
or U19187 (N_19187,N_16569,N_17965);
nand U19188 (N_19188,N_17866,N_17863);
or U19189 (N_19189,N_16650,N_17264);
or U19190 (N_19190,N_17933,N_17614);
nand U19191 (N_19191,N_16656,N_17961);
xor U19192 (N_19192,N_17031,N_16699);
nor U19193 (N_19193,N_17518,N_17228);
or U19194 (N_19194,N_16710,N_17979);
nand U19195 (N_19195,N_16731,N_17181);
nor U19196 (N_19196,N_16698,N_17489);
xnor U19197 (N_19197,N_17193,N_17524);
xnor U19198 (N_19198,N_17148,N_17601);
or U19199 (N_19199,N_17277,N_16836);
xnor U19200 (N_19200,N_16922,N_17128);
nand U19201 (N_19201,N_17283,N_17832);
nor U19202 (N_19202,N_16677,N_17904);
or U19203 (N_19203,N_17555,N_16809);
xnor U19204 (N_19204,N_16974,N_17237);
and U19205 (N_19205,N_17711,N_16525);
or U19206 (N_19206,N_17126,N_17468);
xnor U19207 (N_19207,N_17235,N_17928);
and U19208 (N_19208,N_17486,N_17068);
and U19209 (N_19209,N_16628,N_17957);
or U19210 (N_19210,N_16719,N_17051);
nor U19211 (N_19211,N_17785,N_17754);
xnor U19212 (N_19212,N_17050,N_16760);
or U19213 (N_19213,N_17874,N_17536);
xnor U19214 (N_19214,N_16572,N_17421);
and U19215 (N_19215,N_16610,N_17631);
nand U19216 (N_19216,N_17866,N_16956);
nand U19217 (N_19217,N_17922,N_17773);
nand U19218 (N_19218,N_16737,N_16665);
and U19219 (N_19219,N_17870,N_17899);
or U19220 (N_19220,N_17220,N_17894);
and U19221 (N_19221,N_17793,N_16847);
and U19222 (N_19222,N_17075,N_17050);
nand U19223 (N_19223,N_16865,N_17154);
or U19224 (N_19224,N_16520,N_17922);
nand U19225 (N_19225,N_16895,N_16601);
nand U19226 (N_19226,N_17393,N_16510);
or U19227 (N_19227,N_17621,N_17523);
and U19228 (N_19228,N_16580,N_17282);
and U19229 (N_19229,N_17141,N_17670);
and U19230 (N_19230,N_17639,N_17995);
and U19231 (N_19231,N_16911,N_17969);
nor U19232 (N_19232,N_16634,N_17296);
or U19233 (N_19233,N_16803,N_16792);
nand U19234 (N_19234,N_16582,N_16567);
nor U19235 (N_19235,N_16910,N_17518);
nor U19236 (N_19236,N_17008,N_17875);
nand U19237 (N_19237,N_17225,N_17110);
nand U19238 (N_19238,N_17669,N_16845);
nand U19239 (N_19239,N_17995,N_17230);
xnor U19240 (N_19240,N_16976,N_16819);
xor U19241 (N_19241,N_16604,N_17435);
nand U19242 (N_19242,N_17249,N_16505);
xor U19243 (N_19243,N_17949,N_17620);
or U19244 (N_19244,N_16636,N_16955);
nor U19245 (N_19245,N_17158,N_16821);
nor U19246 (N_19246,N_16795,N_17896);
nor U19247 (N_19247,N_17140,N_16872);
nand U19248 (N_19248,N_16808,N_16524);
and U19249 (N_19249,N_17314,N_17134);
nand U19250 (N_19250,N_17912,N_17719);
and U19251 (N_19251,N_17856,N_17292);
or U19252 (N_19252,N_17475,N_16561);
or U19253 (N_19253,N_16560,N_17583);
nor U19254 (N_19254,N_17156,N_16536);
xor U19255 (N_19255,N_17329,N_17890);
nand U19256 (N_19256,N_17014,N_17775);
nor U19257 (N_19257,N_16550,N_17754);
xor U19258 (N_19258,N_17515,N_17366);
xor U19259 (N_19259,N_17965,N_16996);
and U19260 (N_19260,N_17114,N_17373);
nor U19261 (N_19261,N_17799,N_17599);
nand U19262 (N_19262,N_17465,N_16933);
xnor U19263 (N_19263,N_17021,N_16580);
xor U19264 (N_19264,N_16693,N_17812);
or U19265 (N_19265,N_17785,N_17907);
and U19266 (N_19266,N_16834,N_17601);
nand U19267 (N_19267,N_16899,N_17483);
nor U19268 (N_19268,N_16737,N_17637);
xnor U19269 (N_19269,N_17683,N_17540);
nor U19270 (N_19270,N_17315,N_17708);
and U19271 (N_19271,N_16933,N_17934);
and U19272 (N_19272,N_17595,N_17239);
nand U19273 (N_19273,N_17913,N_16811);
nand U19274 (N_19274,N_17675,N_16838);
xor U19275 (N_19275,N_16852,N_17684);
or U19276 (N_19276,N_17102,N_16974);
or U19277 (N_19277,N_17221,N_16648);
or U19278 (N_19278,N_16640,N_16796);
and U19279 (N_19279,N_16574,N_16769);
and U19280 (N_19280,N_17101,N_17116);
nand U19281 (N_19281,N_17906,N_17939);
xor U19282 (N_19282,N_17777,N_17894);
nor U19283 (N_19283,N_17979,N_17229);
and U19284 (N_19284,N_16672,N_16500);
nand U19285 (N_19285,N_17948,N_17685);
nand U19286 (N_19286,N_17396,N_17976);
nand U19287 (N_19287,N_16834,N_16600);
or U19288 (N_19288,N_17386,N_17623);
xnor U19289 (N_19289,N_17367,N_16756);
and U19290 (N_19290,N_16668,N_17980);
and U19291 (N_19291,N_17526,N_17799);
or U19292 (N_19292,N_17989,N_17533);
nor U19293 (N_19293,N_16935,N_16637);
xnor U19294 (N_19294,N_16933,N_16691);
or U19295 (N_19295,N_17094,N_16567);
xnor U19296 (N_19296,N_17452,N_16550);
and U19297 (N_19297,N_16816,N_17673);
nor U19298 (N_19298,N_17482,N_16693);
and U19299 (N_19299,N_16755,N_17647);
or U19300 (N_19300,N_17840,N_17699);
nand U19301 (N_19301,N_17287,N_17725);
and U19302 (N_19302,N_16598,N_17686);
nor U19303 (N_19303,N_16828,N_17361);
and U19304 (N_19304,N_17105,N_16964);
nor U19305 (N_19305,N_16677,N_17505);
nor U19306 (N_19306,N_16949,N_17710);
nand U19307 (N_19307,N_17152,N_16785);
and U19308 (N_19308,N_17986,N_16872);
xor U19309 (N_19309,N_16582,N_17401);
xnor U19310 (N_19310,N_17948,N_17833);
and U19311 (N_19311,N_16561,N_16770);
nor U19312 (N_19312,N_17910,N_17362);
or U19313 (N_19313,N_17905,N_17706);
and U19314 (N_19314,N_17126,N_17701);
and U19315 (N_19315,N_17785,N_16533);
or U19316 (N_19316,N_17121,N_16637);
nor U19317 (N_19317,N_17628,N_17133);
or U19318 (N_19318,N_17653,N_17587);
nor U19319 (N_19319,N_17681,N_17853);
and U19320 (N_19320,N_16552,N_17170);
nand U19321 (N_19321,N_17665,N_17509);
nand U19322 (N_19322,N_16793,N_17900);
nand U19323 (N_19323,N_17771,N_17508);
nand U19324 (N_19324,N_17226,N_17281);
nand U19325 (N_19325,N_17095,N_17431);
and U19326 (N_19326,N_16892,N_17325);
or U19327 (N_19327,N_17863,N_17516);
xor U19328 (N_19328,N_17687,N_17241);
xor U19329 (N_19329,N_17666,N_17198);
nor U19330 (N_19330,N_17405,N_17699);
xnor U19331 (N_19331,N_16755,N_17895);
nand U19332 (N_19332,N_17708,N_17108);
nand U19333 (N_19333,N_16547,N_16850);
and U19334 (N_19334,N_17182,N_17628);
or U19335 (N_19335,N_16608,N_17367);
or U19336 (N_19336,N_17045,N_17826);
and U19337 (N_19337,N_17864,N_17275);
xnor U19338 (N_19338,N_17477,N_16835);
nand U19339 (N_19339,N_17941,N_17547);
and U19340 (N_19340,N_16648,N_17083);
and U19341 (N_19341,N_16725,N_17890);
xor U19342 (N_19342,N_16778,N_17235);
and U19343 (N_19343,N_17783,N_16513);
nand U19344 (N_19344,N_17244,N_17041);
and U19345 (N_19345,N_17929,N_17757);
nand U19346 (N_19346,N_16600,N_17076);
and U19347 (N_19347,N_16900,N_16864);
or U19348 (N_19348,N_17813,N_17715);
nand U19349 (N_19349,N_16749,N_16716);
or U19350 (N_19350,N_17833,N_17697);
nor U19351 (N_19351,N_17583,N_17700);
or U19352 (N_19352,N_17820,N_16598);
xnor U19353 (N_19353,N_16938,N_17522);
or U19354 (N_19354,N_17032,N_17715);
nand U19355 (N_19355,N_16973,N_17485);
and U19356 (N_19356,N_16917,N_16682);
and U19357 (N_19357,N_17722,N_17252);
or U19358 (N_19358,N_17407,N_17956);
nor U19359 (N_19359,N_17681,N_17320);
and U19360 (N_19360,N_16635,N_16938);
nand U19361 (N_19361,N_16869,N_17630);
and U19362 (N_19362,N_17556,N_16958);
or U19363 (N_19363,N_17845,N_17294);
or U19364 (N_19364,N_17464,N_16529);
xor U19365 (N_19365,N_17810,N_16733);
xnor U19366 (N_19366,N_17528,N_17846);
or U19367 (N_19367,N_17316,N_17449);
nor U19368 (N_19368,N_16535,N_17018);
xnor U19369 (N_19369,N_17754,N_17231);
nand U19370 (N_19370,N_16517,N_17966);
and U19371 (N_19371,N_17924,N_17282);
nand U19372 (N_19372,N_16968,N_16553);
nand U19373 (N_19373,N_17463,N_16654);
nand U19374 (N_19374,N_17142,N_17125);
xnor U19375 (N_19375,N_16513,N_17919);
xor U19376 (N_19376,N_16819,N_17625);
and U19377 (N_19377,N_17500,N_17836);
and U19378 (N_19378,N_16514,N_17730);
xnor U19379 (N_19379,N_17073,N_16622);
or U19380 (N_19380,N_17234,N_17968);
and U19381 (N_19381,N_17380,N_17440);
nand U19382 (N_19382,N_16998,N_17684);
nand U19383 (N_19383,N_17458,N_16629);
nor U19384 (N_19384,N_17797,N_16563);
xnor U19385 (N_19385,N_17316,N_16690);
nor U19386 (N_19386,N_17042,N_17689);
nor U19387 (N_19387,N_17885,N_17817);
xor U19388 (N_19388,N_17969,N_16610);
nor U19389 (N_19389,N_16637,N_17848);
or U19390 (N_19390,N_17557,N_17798);
nor U19391 (N_19391,N_16606,N_17789);
xnor U19392 (N_19392,N_17717,N_17624);
or U19393 (N_19393,N_16507,N_17861);
or U19394 (N_19394,N_16820,N_16582);
or U19395 (N_19395,N_16859,N_16522);
or U19396 (N_19396,N_17367,N_16550);
xor U19397 (N_19397,N_17162,N_17574);
and U19398 (N_19398,N_17957,N_16908);
and U19399 (N_19399,N_17076,N_17433);
xnor U19400 (N_19400,N_17131,N_17735);
nand U19401 (N_19401,N_17665,N_16997);
or U19402 (N_19402,N_17361,N_17354);
xnor U19403 (N_19403,N_17448,N_17912);
nand U19404 (N_19404,N_17499,N_16999);
and U19405 (N_19405,N_17875,N_16828);
nor U19406 (N_19406,N_17654,N_16504);
xor U19407 (N_19407,N_16772,N_17534);
or U19408 (N_19408,N_17008,N_17453);
nor U19409 (N_19409,N_17024,N_16916);
or U19410 (N_19410,N_17441,N_16579);
xor U19411 (N_19411,N_17457,N_17191);
and U19412 (N_19412,N_17869,N_17578);
nor U19413 (N_19413,N_16944,N_17436);
xnor U19414 (N_19414,N_17673,N_17759);
or U19415 (N_19415,N_16524,N_16502);
and U19416 (N_19416,N_17985,N_17072);
xnor U19417 (N_19417,N_17329,N_17688);
nand U19418 (N_19418,N_17848,N_17614);
or U19419 (N_19419,N_17570,N_16769);
and U19420 (N_19420,N_17692,N_16721);
and U19421 (N_19421,N_17233,N_16975);
xnor U19422 (N_19422,N_16672,N_17205);
xnor U19423 (N_19423,N_17904,N_17752);
or U19424 (N_19424,N_17038,N_17774);
or U19425 (N_19425,N_16890,N_16788);
nor U19426 (N_19426,N_17973,N_17505);
xor U19427 (N_19427,N_17784,N_16839);
and U19428 (N_19428,N_17456,N_17903);
nand U19429 (N_19429,N_17212,N_16872);
or U19430 (N_19430,N_16620,N_17193);
and U19431 (N_19431,N_16941,N_17594);
xor U19432 (N_19432,N_16831,N_17094);
and U19433 (N_19433,N_17782,N_17522);
nor U19434 (N_19434,N_17484,N_17244);
xnor U19435 (N_19435,N_17601,N_16683);
nor U19436 (N_19436,N_17840,N_16986);
nor U19437 (N_19437,N_16784,N_17643);
nor U19438 (N_19438,N_17833,N_17658);
nor U19439 (N_19439,N_17838,N_16834);
and U19440 (N_19440,N_17693,N_16977);
nand U19441 (N_19441,N_16591,N_17699);
nand U19442 (N_19442,N_16898,N_17324);
and U19443 (N_19443,N_16768,N_17906);
xor U19444 (N_19444,N_16774,N_17976);
xor U19445 (N_19445,N_16595,N_16687);
xor U19446 (N_19446,N_16687,N_17726);
nor U19447 (N_19447,N_16746,N_17285);
or U19448 (N_19448,N_16545,N_17882);
and U19449 (N_19449,N_16866,N_16981);
nand U19450 (N_19450,N_17243,N_16837);
or U19451 (N_19451,N_17639,N_17856);
xor U19452 (N_19452,N_16566,N_17577);
and U19453 (N_19453,N_17484,N_17473);
nand U19454 (N_19454,N_17554,N_17066);
xnor U19455 (N_19455,N_17578,N_17637);
and U19456 (N_19456,N_17295,N_17492);
nor U19457 (N_19457,N_16599,N_16701);
xor U19458 (N_19458,N_17861,N_16809);
xor U19459 (N_19459,N_17756,N_17321);
and U19460 (N_19460,N_17171,N_16846);
nor U19461 (N_19461,N_17778,N_16879);
nand U19462 (N_19462,N_17334,N_17547);
or U19463 (N_19463,N_17528,N_17706);
nor U19464 (N_19464,N_17615,N_17526);
or U19465 (N_19465,N_16820,N_17434);
or U19466 (N_19466,N_17419,N_17016);
and U19467 (N_19467,N_17891,N_17224);
nor U19468 (N_19468,N_17424,N_16544);
nand U19469 (N_19469,N_17937,N_17017);
or U19470 (N_19470,N_17221,N_16547);
nor U19471 (N_19471,N_17262,N_16588);
or U19472 (N_19472,N_17137,N_17104);
xnor U19473 (N_19473,N_17787,N_17328);
or U19474 (N_19474,N_16853,N_17170);
or U19475 (N_19475,N_17259,N_17038);
or U19476 (N_19476,N_17507,N_16978);
or U19477 (N_19477,N_17986,N_17249);
nand U19478 (N_19478,N_16635,N_17117);
nor U19479 (N_19479,N_16516,N_16566);
or U19480 (N_19480,N_17190,N_17439);
or U19481 (N_19481,N_17537,N_16584);
or U19482 (N_19482,N_17055,N_17992);
nand U19483 (N_19483,N_17038,N_17751);
xor U19484 (N_19484,N_17145,N_17497);
nand U19485 (N_19485,N_16686,N_17477);
nor U19486 (N_19486,N_17131,N_16674);
xnor U19487 (N_19487,N_17352,N_16881);
xor U19488 (N_19488,N_17029,N_17322);
nor U19489 (N_19489,N_16750,N_16697);
nor U19490 (N_19490,N_16714,N_17399);
xnor U19491 (N_19491,N_17574,N_16939);
nand U19492 (N_19492,N_16928,N_16773);
xnor U19493 (N_19493,N_16777,N_16632);
or U19494 (N_19494,N_16911,N_16884);
or U19495 (N_19495,N_17010,N_16774);
nor U19496 (N_19496,N_17981,N_17810);
nor U19497 (N_19497,N_17418,N_17545);
nor U19498 (N_19498,N_16682,N_17782);
xor U19499 (N_19499,N_17387,N_17069);
or U19500 (N_19500,N_18693,N_18493);
or U19501 (N_19501,N_18454,N_18767);
nand U19502 (N_19502,N_19024,N_19477);
or U19503 (N_19503,N_18083,N_18045);
nor U19504 (N_19504,N_18340,N_18386);
and U19505 (N_19505,N_18319,N_19353);
nor U19506 (N_19506,N_18849,N_19136);
nor U19507 (N_19507,N_18635,N_19358);
nand U19508 (N_19508,N_18729,N_19314);
nor U19509 (N_19509,N_18309,N_18543);
nor U19510 (N_19510,N_18545,N_19365);
and U19511 (N_19511,N_18449,N_19191);
nor U19512 (N_19512,N_19349,N_19035);
or U19513 (N_19513,N_19258,N_19483);
or U19514 (N_19514,N_18660,N_18283);
nand U19515 (N_19515,N_18646,N_18297);
and U19516 (N_19516,N_18223,N_18916);
xnor U19517 (N_19517,N_19352,N_18005);
and U19518 (N_19518,N_19146,N_19327);
nor U19519 (N_19519,N_18194,N_18517);
nand U19520 (N_19520,N_19414,N_18908);
or U19521 (N_19521,N_18117,N_18534);
xor U19522 (N_19522,N_18164,N_18448);
and U19523 (N_19523,N_18671,N_18287);
or U19524 (N_19524,N_19206,N_19152);
nor U19525 (N_19525,N_19045,N_18930);
nor U19526 (N_19526,N_19490,N_18112);
xnor U19527 (N_19527,N_18709,N_19079);
or U19528 (N_19528,N_19217,N_18816);
nand U19529 (N_19529,N_18828,N_18688);
nand U19530 (N_19530,N_19297,N_18277);
nand U19531 (N_19531,N_18697,N_18648);
nor U19532 (N_19532,N_19244,N_18516);
nor U19533 (N_19533,N_19243,N_18855);
nand U19534 (N_19534,N_18244,N_18274);
xor U19535 (N_19535,N_18554,N_19169);
or U19536 (N_19536,N_18668,N_18644);
and U19537 (N_19537,N_19157,N_18181);
or U19538 (N_19538,N_18375,N_18626);
and U19539 (N_19539,N_19200,N_19451);
xor U19540 (N_19540,N_19446,N_18845);
nand U19541 (N_19541,N_18384,N_18861);
or U19542 (N_19542,N_19304,N_18048);
and U19543 (N_19543,N_19480,N_18102);
nand U19544 (N_19544,N_18457,N_18409);
xor U19545 (N_19545,N_18561,N_18848);
nor U19546 (N_19546,N_19094,N_18834);
nor U19547 (N_19547,N_18302,N_18445);
nor U19548 (N_19548,N_19404,N_18760);
or U19549 (N_19549,N_18461,N_18795);
nor U19550 (N_19550,N_19274,N_18405);
and U19551 (N_19551,N_18874,N_18503);
and U19552 (N_19552,N_18902,N_18242);
and U19553 (N_19553,N_18216,N_19050);
and U19554 (N_19554,N_19372,N_19322);
nand U19555 (N_19555,N_18433,N_18796);
and U19556 (N_19556,N_19034,N_18993);
nand U19557 (N_19557,N_19259,N_18326);
nor U19558 (N_19558,N_18490,N_18155);
and U19559 (N_19559,N_18969,N_18498);
xor U19560 (N_19560,N_18122,N_19474);
nand U19561 (N_19561,N_18583,N_18706);
xor U19562 (N_19562,N_18602,N_18723);
and U19563 (N_19563,N_18419,N_18803);
xor U19564 (N_19564,N_18379,N_18566);
nor U19565 (N_19565,N_18156,N_18754);
and U19566 (N_19566,N_18171,N_18264);
or U19567 (N_19567,N_19323,N_19091);
and U19568 (N_19568,N_18183,N_18530);
nand U19569 (N_19569,N_18696,N_18416);
and U19570 (N_19570,N_19184,N_19311);
and U19571 (N_19571,N_18794,N_18368);
or U19572 (N_19572,N_18486,N_19343);
xor U19573 (N_19573,N_18891,N_19456);
or U19574 (N_19574,N_19465,N_18841);
or U19575 (N_19575,N_18336,N_18019);
or U19576 (N_19576,N_18695,N_19129);
xnor U19577 (N_19577,N_18612,N_19292);
xnor U19578 (N_19578,N_18187,N_18506);
xnor U19579 (N_19579,N_18228,N_19239);
and U19580 (N_19580,N_18616,N_18995);
and U19581 (N_19581,N_18320,N_18768);
xor U19582 (N_19582,N_19484,N_18808);
nor U19583 (N_19583,N_18197,N_18650);
and U19584 (N_19584,N_18582,N_18331);
or U19585 (N_19585,N_18867,N_19100);
nor U19586 (N_19586,N_19105,N_19405);
or U19587 (N_19587,N_19312,N_19168);
and U19588 (N_19588,N_19076,N_19291);
nand U19589 (N_19589,N_18233,N_19084);
xnor U19590 (N_19590,N_18470,N_19262);
nor U19591 (N_19591,N_19143,N_18338);
nand U19592 (N_19592,N_18238,N_19166);
or U19593 (N_19593,N_18126,N_19495);
nor U19594 (N_19594,N_18741,N_18960);
and U19595 (N_19595,N_19163,N_18086);
xor U19596 (N_19596,N_19328,N_18017);
nor U19597 (N_19597,N_18676,N_18664);
and U19598 (N_19598,N_19317,N_18512);
and U19599 (N_19599,N_18686,N_18452);
nand U19600 (N_19600,N_18103,N_18492);
nor U19601 (N_19601,N_18414,N_19190);
xor U19602 (N_19602,N_18868,N_18275);
nor U19603 (N_19603,N_18429,N_19260);
or U19604 (N_19604,N_19072,N_19207);
xor U19605 (N_19605,N_18392,N_18897);
and U19606 (N_19606,N_18716,N_19131);
nor U19607 (N_19607,N_18356,N_19361);
and U19608 (N_19608,N_19144,N_19085);
nor U19609 (N_19609,N_18964,N_18608);
nor U19610 (N_19610,N_19121,N_18946);
and U19611 (N_19611,N_18026,N_18401);
xnor U19612 (N_19612,N_18888,N_18016);
nor U19613 (N_19613,N_18121,N_18611);
or U19614 (N_19614,N_19153,N_18988);
nand U19615 (N_19615,N_19102,N_18776);
or U19616 (N_19616,N_18489,N_18481);
or U19617 (N_19617,N_18549,N_18184);
and U19618 (N_19618,N_19042,N_18826);
and U19619 (N_19619,N_19038,N_19175);
and U19620 (N_19620,N_19266,N_19491);
and U19621 (N_19621,N_19057,N_18115);
or U19622 (N_19622,N_19473,N_18631);
or U19623 (N_19623,N_18865,N_18087);
nand U19624 (N_19624,N_19204,N_18621);
or U19625 (N_19625,N_18196,N_18278);
nand U19626 (N_19626,N_18797,N_18022);
or U19627 (N_19627,N_18259,N_18674);
nand U19628 (N_19628,N_19212,N_19338);
or U19629 (N_19629,N_19019,N_18496);
and U19630 (N_19630,N_18784,N_19160);
nand U19631 (N_19631,N_18685,N_19188);
nor U19632 (N_19632,N_18251,N_18509);
or U19633 (N_19633,N_18195,N_18254);
xnor U19634 (N_19634,N_18940,N_19049);
nor U19635 (N_19635,N_18010,N_18465);
xnor U19636 (N_19636,N_18243,N_18472);
xor U19637 (N_19637,N_18204,N_18292);
xnor U19638 (N_19638,N_18159,N_18950);
or U19639 (N_19639,N_19181,N_18589);
xor U19640 (N_19640,N_18057,N_19119);
nor U19641 (N_19641,N_19099,N_19060);
nor U19642 (N_19642,N_18847,N_18479);
or U19643 (N_19643,N_18476,N_19308);
nand U19644 (N_19644,N_18529,N_19296);
nand U19645 (N_19645,N_18771,N_18374);
nand U19646 (N_19646,N_18799,N_19108);
or U19647 (N_19647,N_18047,N_18176);
xnor U19648 (N_19648,N_18550,N_19123);
nor U19649 (N_19649,N_18381,N_18008);
nand U19650 (N_19650,N_18645,N_18820);
xnor U19651 (N_19651,N_18248,N_18373);
nand U19652 (N_19652,N_18630,N_18443);
xor U19653 (N_19653,N_18728,N_18200);
or U19654 (N_19654,N_19278,N_18748);
and U19655 (N_19655,N_18180,N_18221);
xnor U19656 (N_19656,N_18444,N_19230);
xnor U19657 (N_19657,N_18604,N_19013);
xnor U19658 (N_19658,N_18218,N_18568);
and U19659 (N_19659,N_19417,N_18012);
or U19660 (N_19660,N_19089,N_18442);
and U19661 (N_19661,N_18961,N_18640);
or U19662 (N_19662,N_18227,N_18347);
nand U19663 (N_19663,N_19329,N_18842);
and U19664 (N_19664,N_18835,N_19364);
or U19665 (N_19665,N_18641,N_19431);
nor U19666 (N_19666,N_18970,N_18974);
and U19667 (N_19667,N_19149,N_18118);
or U19668 (N_19668,N_18172,N_19186);
nand U19669 (N_19669,N_19211,N_19059);
nor U19670 (N_19670,N_18214,N_18323);
xor U19671 (N_19671,N_18252,N_18541);
nor U19672 (N_19672,N_18203,N_18025);
or U19673 (N_19673,N_18877,N_18034);
or U19674 (N_19674,N_18939,N_18355);
xnor U19675 (N_19675,N_18968,N_18286);
xnor U19676 (N_19676,N_19251,N_19133);
nor U19677 (N_19677,N_18864,N_18513);
and U19678 (N_19678,N_18889,N_18539);
or U19679 (N_19679,N_18963,N_18321);
and U19680 (N_19680,N_19093,N_18471);
xnor U19681 (N_19681,N_18191,N_18229);
and U19682 (N_19682,N_18410,N_19226);
nand U19683 (N_19683,N_18198,N_19137);
or U19684 (N_19684,N_19192,N_18138);
xnor U19685 (N_19685,N_18596,N_18033);
xnor U19686 (N_19686,N_18487,N_18436);
nand U19687 (N_19687,N_19039,N_19418);
nand U19688 (N_19688,N_18036,N_19003);
xnor U19689 (N_19689,N_19498,N_18819);
nor U19690 (N_19690,N_18982,N_19378);
or U19691 (N_19691,N_18898,N_18704);
and U19692 (N_19692,N_19098,N_18128);
and U19693 (N_19693,N_18058,N_18735);
xnor U19694 (N_19694,N_18967,N_19111);
nor U19695 (N_19695,N_18617,N_18189);
and U19696 (N_19696,N_18140,N_18722);
and U19697 (N_19697,N_18018,N_19124);
nor U19698 (N_19698,N_18193,N_18689);
or U19699 (N_19699,N_18300,N_18399);
nand U19700 (N_19700,N_18348,N_19159);
nand U19701 (N_19701,N_19265,N_18619);
or U19702 (N_19702,N_18120,N_19007);
or U19703 (N_19703,N_18468,N_18719);
xnor U19704 (N_19704,N_18753,N_18814);
nand U19705 (N_19705,N_19075,N_19242);
nand U19706 (N_19706,N_18623,N_18153);
nor U19707 (N_19707,N_18724,N_19028);
and U19708 (N_19708,N_18001,N_18170);
nor U19709 (N_19709,N_18850,N_19370);
nor U19710 (N_19710,N_19269,N_18605);
nand U19711 (N_19711,N_18677,N_18708);
or U19712 (N_19712,N_19032,N_18106);
and U19713 (N_19713,N_18592,N_18606);
and U19714 (N_19714,N_18294,N_18406);
xnor U19715 (N_19715,N_18084,N_18337);
xor U19716 (N_19716,N_18143,N_18522);
and U19717 (N_19717,N_18876,N_18966);
and U19718 (N_19718,N_18290,N_19344);
and U19719 (N_19719,N_19320,N_19205);
nor U19720 (N_19720,N_18772,N_18823);
nor U19721 (N_19721,N_19441,N_18114);
nor U19722 (N_19722,N_19330,N_19331);
or U19723 (N_19723,N_18839,N_19396);
nand U19724 (N_19724,N_19382,N_18332);
and U19725 (N_19725,N_18928,N_18261);
and U19726 (N_19726,N_19453,N_19310);
nor U19727 (N_19727,N_18149,N_18577);
nor U19728 (N_19728,N_18766,N_18901);
nor U19729 (N_19729,N_19415,N_19082);
xnor U19730 (N_19730,N_19257,N_18569);
nand U19731 (N_19731,N_18004,N_18109);
or U19732 (N_19732,N_19302,N_18060);
and U19733 (N_19733,N_19340,N_18832);
or U19734 (N_19734,N_19475,N_18413);
and U19735 (N_19735,N_19346,N_19041);
xor U19736 (N_19736,N_18127,N_19360);
nand U19737 (N_19737,N_18315,N_18307);
or U19738 (N_19738,N_19020,N_19234);
nor U19739 (N_19739,N_19301,N_18391);
nor U19740 (N_19740,N_19387,N_18024);
and U19741 (N_19741,N_18327,N_19288);
xor U19742 (N_19742,N_18777,N_19010);
and U19743 (N_19743,N_18711,N_18167);
and U19744 (N_19744,N_19359,N_18934);
and U19745 (N_19745,N_19454,N_18717);
nor U19746 (N_19746,N_18770,N_19012);
or U19747 (N_19747,N_18923,N_19196);
nor U19748 (N_19748,N_18871,N_19427);
nor U19749 (N_19749,N_18812,N_18279);
nand U19750 (N_19750,N_18725,N_18335);
xor U19751 (N_19751,N_18021,N_18459);
xor U19752 (N_19752,N_19351,N_18586);
nor U19753 (N_19753,N_18535,N_18484);
and U19754 (N_19754,N_18634,N_18032);
and U19755 (N_19755,N_18482,N_19276);
xor U19756 (N_19756,N_18978,N_19247);
or U19757 (N_19757,N_18973,N_19113);
xor U19758 (N_19758,N_18730,N_18791);
nor U19759 (N_19759,N_19088,N_18029);
nor U19760 (N_19760,N_19435,N_18380);
nor U19761 (N_19761,N_19332,N_18949);
xor U19762 (N_19762,N_18972,N_19017);
xnor U19763 (N_19763,N_18169,N_18639);
and U19764 (N_19764,N_19334,N_18069);
xnor U19765 (N_19765,N_18202,N_18752);
nor U19766 (N_19766,N_19367,N_19250);
nor U19767 (N_19767,N_18137,N_18986);
nor U19768 (N_19768,N_18291,N_18657);
nand U19769 (N_19769,N_18237,N_18378);
nand U19770 (N_19770,N_18312,N_19161);
nand U19771 (N_19771,N_18552,N_18937);
nand U19772 (N_19772,N_18093,N_18466);
nand U19773 (N_19773,N_18129,N_18130);
nor U19774 (N_19774,N_18737,N_18962);
or U19775 (N_19775,N_19101,N_18002);
or U19776 (N_19776,N_19097,N_18663);
xnor U19777 (N_19777,N_19164,N_18821);
and U19778 (N_19778,N_18316,N_19277);
nand U19779 (N_19779,N_19369,N_18996);
xor U19780 (N_19780,N_18288,N_19268);
or U19781 (N_19781,N_18351,N_18765);
or U19782 (N_19782,N_18975,N_18840);
nand U19783 (N_19783,N_18654,N_19392);
or U19784 (N_19784,N_19222,N_18370);
nand U19785 (N_19785,N_19120,N_18144);
xnor U19786 (N_19786,N_19033,N_18105);
nor U19787 (N_19787,N_18494,N_18330);
and U19788 (N_19788,N_18505,N_18070);
nand U19789 (N_19789,N_18843,N_19114);
or U19790 (N_19790,N_18670,N_18756);
xor U19791 (N_19791,N_18495,N_19496);
or U19792 (N_19792,N_18418,N_18232);
and U19793 (N_19793,N_18502,N_19235);
and U19794 (N_19794,N_19051,N_18651);
or U19795 (N_19795,N_18382,N_18064);
nor U19796 (N_19796,N_19363,N_18107);
nor U19797 (N_19797,N_19240,N_19064);
nor U19798 (N_19798,N_18111,N_18721);
nor U19799 (N_19799,N_18726,N_18041);
xor U19800 (N_19800,N_18104,N_19112);
or U19801 (N_19801,N_18357,N_19345);
or U19802 (N_19802,N_18562,N_18249);
xnor U19803 (N_19803,N_18636,N_18162);
or U19804 (N_19804,N_18584,N_18758);
nor U19805 (N_19805,N_18925,N_18225);
nor U19806 (N_19806,N_18396,N_18329);
or U19807 (N_19807,N_18455,N_18376);
nor U19808 (N_19808,N_19037,N_19444);
xor U19809 (N_19809,N_19214,N_18903);
and U19810 (N_19810,N_18751,N_18460);
and U19811 (N_19811,N_18652,N_19225);
nor U19812 (N_19812,N_18152,N_18628);
nand U19813 (N_19813,N_18510,N_18720);
or U19814 (N_19814,N_19104,N_19027);
and U19815 (N_19815,N_19021,N_18878);
and U19816 (N_19816,N_18453,N_18398);
xor U19817 (N_19817,N_19377,N_19249);
nor U19818 (N_19818,N_18407,N_19272);
nor U19819 (N_19819,N_18478,N_18295);
xor U19820 (N_19820,N_19397,N_19065);
xnor U19821 (N_19821,N_18071,N_18653);
nand U19822 (N_19822,N_18310,N_19463);
xor U19823 (N_19823,N_18718,N_19298);
or U19824 (N_19824,N_18833,N_18792);
and U19825 (N_19825,N_18591,N_18798);
xnor U19826 (N_19826,N_18423,N_18762);
xor U19827 (N_19827,N_18936,N_18918);
or U19828 (N_19828,N_19122,N_18136);
xnor U19829 (N_19829,N_19147,N_18343);
nor U19830 (N_19830,N_18304,N_19371);
xnor U19831 (N_19831,N_19455,N_18692);
nor U19832 (N_19832,N_18097,N_18615);
xor U19833 (N_19833,N_19096,N_19246);
xor U19834 (N_19834,N_18280,N_18428);
nand U19835 (N_19835,N_18558,N_18763);
and U19836 (N_19836,N_19255,N_19460);
nand U19837 (N_19837,N_19167,N_18055);
and U19838 (N_19838,N_19125,N_18257);
nor U19839 (N_19839,N_18388,N_18917);
xnor U19840 (N_19840,N_19466,N_19134);
nor U19841 (N_19841,N_18637,N_19031);
or U19842 (N_19842,N_19151,N_18145);
and U19843 (N_19843,N_18667,N_18345);
xnor U19844 (N_19844,N_18669,N_19380);
nor U19845 (N_19845,N_18914,N_18713);
and U19846 (N_19846,N_18077,N_18563);
nand U19847 (N_19847,N_19106,N_18383);
nand U19848 (N_19848,N_19450,N_19478);
and U19849 (N_19849,N_18125,N_18023);
nor U19850 (N_19850,N_18015,N_19178);
and U19851 (N_19851,N_18456,N_18234);
nor U19852 (N_19852,N_19406,N_18272);
nor U19853 (N_19853,N_18740,N_19410);
nor U19854 (N_19854,N_19400,N_19285);
nor U19855 (N_19855,N_18750,N_18020);
and U19856 (N_19856,N_19126,N_18464);
xnor U19857 (N_19857,N_18882,N_19081);
nand U19858 (N_19858,N_18096,N_19135);
nor U19859 (N_19859,N_18361,N_18743);
and U19860 (N_19860,N_18747,N_19236);
xor U19861 (N_19861,N_18235,N_19398);
xor U19862 (N_19862,N_19208,N_18824);
or U19863 (N_19863,N_18684,N_19472);
and U19864 (N_19864,N_18094,N_18553);
nor U19865 (N_19865,N_18907,N_18372);
and U19866 (N_19866,N_19103,N_19229);
nor U19867 (N_19867,N_18945,N_18879);
nand U19868 (N_19868,N_19118,N_19385);
or U19869 (N_19869,N_18009,N_19399);
xor U19870 (N_19870,N_18220,N_18014);
nor U19871 (N_19871,N_18177,N_18404);
nand U19872 (N_19872,N_19183,N_18095);
xnor U19873 (N_19873,N_18778,N_18303);
nor U19874 (N_19874,N_18926,N_19061);
and U19875 (N_19875,N_18518,N_18977);
or U19876 (N_19876,N_18857,N_18053);
or U19877 (N_19877,N_18941,N_19073);
nand U19878 (N_19878,N_19366,N_19368);
nand U19879 (N_19879,N_19290,N_19083);
xnor U19880 (N_19880,N_19248,N_19429);
or U19881 (N_19881,N_18655,N_18075);
nor U19882 (N_19882,N_19386,N_18201);
nand U19883 (N_19883,N_19138,N_18265);
and U19884 (N_19884,N_19139,N_18727);
nor U19885 (N_19885,N_18594,N_18825);
nor U19886 (N_19886,N_19279,N_18134);
nand U19887 (N_19887,N_18932,N_18691);
and U19888 (N_19888,N_18186,N_19150);
or U19889 (N_19889,N_19422,N_18827);
nor U19890 (N_19890,N_18862,N_18146);
or U19891 (N_19891,N_19018,N_19201);
or U19892 (N_19892,N_18869,N_19409);
nor U19893 (N_19893,N_18560,N_18567);
and U19894 (N_19894,N_19155,N_19256);
or U19895 (N_19895,N_19375,N_19005);
and U19896 (N_19896,N_19052,N_19030);
xnor U19897 (N_19897,N_18013,N_19174);
nand U19898 (N_19898,N_19305,N_18759);
or U19899 (N_19899,N_19437,N_18885);
nor U19900 (N_19900,N_18957,N_18595);
nand U19901 (N_19901,N_18074,N_18948);
and U19902 (N_19902,N_18698,N_18385);
nand U19903 (N_19903,N_18354,N_18301);
and U19904 (N_19904,N_19238,N_18955);
nor U19905 (N_19905,N_18369,N_18944);
or U19906 (N_19906,N_19336,N_18887);
nor U19907 (N_19907,N_18942,N_18205);
xor U19908 (N_19908,N_18813,N_19132);
nand U19909 (N_19909,N_18099,N_18090);
xor U19910 (N_19910,N_19165,N_18076);
xnor U19911 (N_19911,N_19390,N_18881);
nand U19912 (N_19912,N_18168,N_18421);
nand U19913 (N_19913,N_19179,N_18998);
nor U19914 (N_19914,N_18899,N_18933);
xnor U19915 (N_19915,N_18051,N_19185);
nand U19916 (N_19916,N_18514,N_19428);
or U19917 (N_19917,N_18904,N_18062);
xor U19918 (N_19918,N_19117,N_19048);
or U19919 (N_19919,N_18000,N_18206);
and U19920 (N_19920,N_19189,N_18638);
xnor U19921 (N_19921,N_19040,N_18629);
and U19922 (N_19922,N_18802,N_19215);
or U19923 (N_19923,N_18038,N_18811);
xor U19924 (N_19924,N_18987,N_18597);
or U19925 (N_19925,N_18700,N_19170);
nor U19926 (N_19926,N_18895,N_18893);
nor U19927 (N_19927,N_18426,N_19394);
nor U19928 (N_19928,N_18285,N_18538);
nand U19929 (N_19929,N_19252,N_18922);
nor U19930 (N_19930,N_18226,N_18165);
and U19931 (N_19931,N_18851,N_19086);
xnor U19932 (N_19932,N_18683,N_18714);
xnor U19933 (N_19933,N_18665,N_19202);
xor U19934 (N_19934,N_18800,N_18147);
and U19935 (N_19935,N_18483,N_19324);
nand U19936 (N_19936,N_18603,N_18788);
xor U19937 (N_19937,N_19182,N_18981);
nand U19938 (N_19938,N_19493,N_18931);
or U19939 (N_19939,N_19300,N_18324);
and U19940 (N_19940,N_18293,N_18523);
nand U19941 (N_19941,N_18035,N_18507);
or U19942 (N_19942,N_18157,N_18432);
or U19943 (N_19943,N_18625,N_19289);
and U19944 (N_19944,N_18992,N_18815);
or U19945 (N_19945,N_18953,N_19177);
nor U19946 (N_19946,N_18980,N_18705);
nor U19947 (N_19947,N_19321,N_18098);
nor U19948 (N_19948,N_18040,N_18927);
xor U19949 (N_19949,N_18052,N_19411);
nand U19950 (N_19950,N_18360,N_18417);
or U19951 (N_19951,N_19011,N_19492);
nand U19952 (N_19952,N_18031,N_18921);
nand U19953 (N_19953,N_18160,N_18593);
and U19954 (N_19954,N_18402,N_18462);
or U19955 (N_19955,N_18081,N_19194);
and U19956 (N_19956,N_18497,N_18469);
or U19957 (N_19957,N_19449,N_18647);
or U19958 (N_19958,N_18311,N_18527);
or U19959 (N_19959,N_19342,N_18439);
nor U19960 (N_19960,N_18804,N_18817);
or U19961 (N_19961,N_18999,N_18082);
nand U19962 (N_19962,N_18089,N_18614);
xor U19963 (N_19963,N_18480,N_18829);
nor U19964 (N_19964,N_18192,N_19293);
or U19965 (N_19965,N_18377,N_18943);
and U19966 (N_19966,N_19379,N_18158);
and U19967 (N_19967,N_18672,N_18662);
xor U19968 (N_19968,N_19068,N_18151);
or U19969 (N_19969,N_18182,N_18687);
or U19970 (N_19970,N_18458,N_18920);
and U19971 (N_19971,N_18546,N_18570);
or U19972 (N_19972,N_19044,N_18838);
nor U19973 (N_19973,N_19002,N_18131);
or U19974 (N_19974,N_18929,N_19471);
and U19975 (N_19975,N_19403,N_18209);
and U19976 (N_19976,N_19130,N_18954);
and U19977 (N_19977,N_18906,N_18175);
and U19978 (N_19978,N_18585,N_18148);
nor U19979 (N_19979,N_19376,N_18971);
nand U19980 (N_19980,N_18190,N_19221);
and U19981 (N_19981,N_18976,N_18352);
nor U19982 (N_19982,N_18707,N_19333);
nor U19983 (N_19983,N_19313,N_19462);
and U19984 (N_19984,N_18951,N_18306);
and U19985 (N_19985,N_18702,N_19487);
or U19986 (N_19986,N_19461,N_18736);
xor U19987 (N_19987,N_18178,N_18599);
and U19988 (N_19988,N_19128,N_18959);
and U19989 (N_19989,N_18427,N_18006);
nor U19990 (N_19990,N_18859,N_18011);
and U19991 (N_19991,N_18346,N_19419);
nor U19992 (N_19992,N_18536,N_18387);
xor U19993 (N_19993,N_18440,N_18618);
nand U19994 (N_19994,N_18984,N_18579);
xnor U19995 (N_19995,N_19267,N_18501);
nor U19996 (N_19996,N_19299,N_18079);
or U19997 (N_19997,N_19271,N_18547);
xor U19998 (N_19998,N_18296,N_18764);
xnor U19999 (N_19999,N_18912,N_18185);
xnor U20000 (N_20000,N_19341,N_18807);
nand U20001 (N_20001,N_18211,N_18135);
and U20002 (N_20002,N_18350,N_18322);
nor U20003 (N_20003,N_18990,N_18333);
nor U20004 (N_20004,N_18588,N_18213);
xnor U20005 (N_20005,N_19187,N_19499);
nand U20006 (N_20006,N_18210,N_19439);
nand U20007 (N_20007,N_18787,N_18699);
xnor U20008 (N_20008,N_18581,N_19090);
xor U20009 (N_20009,N_19384,N_19281);
and U20010 (N_20010,N_18199,N_19047);
nand U20011 (N_20011,N_18425,N_19115);
xor U20012 (N_20012,N_18837,N_18818);
or U20013 (N_20013,N_18952,N_19316);
and U20014 (N_20014,N_19231,N_18124);
xnor U20015 (N_20015,N_18900,N_18622);
nor U20016 (N_20016,N_18116,N_18499);
or U20017 (N_20017,N_18367,N_18779);
or U20018 (N_20018,N_19046,N_18854);
nand U20019 (N_20019,N_18555,N_18281);
or U20020 (N_20020,N_18793,N_18790);
nor U20021 (N_20021,N_19350,N_18810);
xor U20022 (N_20022,N_18991,N_18339);
xnor U20023 (N_20023,N_18113,N_19087);
xnor U20024 (N_20024,N_18110,N_18403);
or U20025 (N_20025,N_19430,N_18710);
nor U20026 (N_20026,N_19245,N_18263);
nand U20027 (N_20027,N_18166,N_19315);
and U20028 (N_20028,N_18508,N_18271);
and U20029 (N_20029,N_19162,N_18318);
or U20030 (N_20030,N_19148,N_18363);
nand U20031 (N_20031,N_18068,N_18883);
nor U20032 (N_20032,N_18245,N_18390);
nor U20033 (N_20033,N_19482,N_19176);
xor U20034 (N_20034,N_19339,N_18935);
and U20035 (N_20035,N_18852,N_18731);
and U20036 (N_20036,N_18738,N_18435);
and U20037 (N_20037,N_18276,N_19015);
nor U20038 (N_20038,N_18573,N_19053);
nor U20039 (N_20039,N_18694,N_18371);
or U20040 (N_20040,N_18600,N_18142);
nor U20041 (N_20041,N_19295,N_18732);
or U20042 (N_20042,N_18846,N_18042);
and U20043 (N_20043,N_19171,N_18544);
nor U20044 (N_20044,N_19055,N_18682);
nand U20045 (N_20045,N_18246,N_18441);
and U20046 (N_20046,N_19218,N_19457);
xor U20047 (N_20047,N_18773,N_19241);
nand U20048 (N_20048,N_18299,N_18715);
or U20049 (N_20049,N_18063,N_19432);
or U20050 (N_20050,N_18365,N_18774);
nor U20051 (N_20051,N_19420,N_18054);
nor U20052 (N_20052,N_18028,N_18132);
xor U20053 (N_20053,N_19347,N_19158);
nand U20054 (N_20054,N_18703,N_19172);
and U20055 (N_20055,N_19424,N_18872);
xor U20056 (N_20056,N_19016,N_19092);
nor U20057 (N_20057,N_18208,N_18870);
nor U20058 (N_20058,N_18911,N_18632);
xnor U20059 (N_20059,N_19286,N_18886);
nor U20060 (N_20060,N_18532,N_19067);
xor U20061 (N_20061,N_19443,N_18313);
and U20062 (N_20062,N_18072,N_18269);
nand U20063 (N_20063,N_18681,N_19209);
and U20064 (N_20064,N_18609,N_18389);
nand U20065 (N_20065,N_18359,N_18801);
and U20066 (N_20066,N_19008,N_18526);
nor U20067 (N_20067,N_19043,N_19283);
xor U20068 (N_20068,N_19001,N_19452);
and U20069 (N_20069,N_19391,N_18919);
nand U20070 (N_20070,N_18656,N_19280);
nor U20071 (N_20071,N_18043,N_19077);
nand U20072 (N_20072,N_18207,N_19335);
nand U20073 (N_20073,N_18450,N_19232);
or U20074 (N_20074,N_18633,N_18601);
nand U20075 (N_20075,N_19326,N_19210);
nand U20076 (N_20076,N_19408,N_19434);
or U20077 (N_20077,N_18624,N_18451);
xor U20078 (N_20078,N_19412,N_19253);
or U20079 (N_20079,N_18956,N_18781);
and U20080 (N_20080,N_19198,N_18431);
nor U20081 (N_20081,N_18393,N_18873);
nand U20082 (N_20082,N_19022,N_18521);
or U20083 (N_20083,N_18679,N_19036);
xor U20084 (N_20084,N_18091,N_19095);
nor U20085 (N_20085,N_18786,N_19109);
and U20086 (N_20086,N_18913,N_18438);
nor U20087 (N_20087,N_19389,N_18230);
and U20088 (N_20088,N_19436,N_18108);
nor U20089 (N_20089,N_19009,N_19354);
nand U20090 (N_20090,N_19142,N_19447);
or U20091 (N_20091,N_18412,N_18305);
xnor U20092 (N_20092,N_19402,N_18119);
xnor U20093 (N_20093,N_18892,N_19489);
xor U20094 (N_20094,N_18783,N_18349);
nand U20095 (N_20095,N_18531,N_18358);
xor U20096 (N_20096,N_18314,N_18548);
or U20097 (N_20097,N_19025,N_19071);
and U20098 (N_20098,N_18782,N_18649);
nor U20099 (N_20099,N_19180,N_18282);
and U20100 (N_20100,N_18905,N_18712);
or U20101 (N_20101,N_18485,N_19004);
nor U20102 (N_20102,N_18519,N_18217);
or U20103 (N_20103,N_19356,N_18092);
and U20104 (N_20104,N_18044,N_18989);
nor U20105 (N_20105,N_18733,N_18858);
nand U20106 (N_20106,N_19433,N_18173);
nor U20107 (N_20107,N_19141,N_18910);
xor U20108 (N_20108,N_19393,N_18806);
nor U20109 (N_20109,N_18580,N_19058);
xnor U20110 (N_20110,N_18154,N_18260);
and U20111 (N_20111,N_19494,N_19014);
nand U20112 (N_20112,N_18050,N_18039);
nor U20113 (N_20113,N_18610,N_18411);
and U20114 (N_20114,N_18924,N_18643);
xor U20115 (N_20115,N_18415,N_18270);
or U20116 (N_20116,N_18161,N_18066);
or U20117 (N_20117,N_19056,N_18742);
and U20118 (N_20118,N_18947,N_18575);
nor U20119 (N_20119,N_19154,N_18537);
nor U20120 (N_20120,N_18863,N_19228);
and U20121 (N_20121,N_18475,N_18078);
and U20122 (N_20122,N_19270,N_19140);
xnor U20123 (N_20123,N_18236,N_19306);
xnor U20124 (N_20124,N_18805,N_18620);
xor U20125 (N_20125,N_18325,N_18477);
and U20126 (N_20126,N_19173,N_18884);
or U20127 (N_20127,N_19374,N_18559);
nor U20128 (N_20128,N_18253,N_18215);
nor U20129 (N_20129,N_18262,N_19069);
nor U20130 (N_20130,N_19381,N_18434);
and U20131 (N_20131,N_19080,N_18446);
and U20132 (N_20132,N_18860,N_18150);
xor U20133 (N_20133,N_19107,N_18342);
or U20134 (N_20134,N_18734,N_18607);
nor U20135 (N_20135,N_19294,N_19263);
or U20136 (N_20136,N_18268,N_18661);
nand U20137 (N_20137,N_18100,N_18141);
nand U20138 (N_20138,N_18267,N_18328);
and U20139 (N_20139,N_18528,N_19216);
and U20140 (N_20140,N_18574,N_19318);
nor U20141 (N_20141,N_18500,N_18997);
nand U20142 (N_20142,N_19469,N_19476);
or U20143 (N_20143,N_18938,N_19127);
nor U20144 (N_20144,N_18394,N_18007);
xnor U20145 (N_20145,N_18853,N_19199);
nor U20146 (N_20146,N_18133,N_19348);
nand U20147 (N_20147,N_18447,N_19497);
nor U20148 (N_20148,N_18065,N_18785);
nor U20149 (N_20149,N_18769,N_18212);
nor U20150 (N_20150,N_18488,N_19373);
nand U20151 (N_20151,N_18344,N_19337);
and U20152 (N_20152,N_18701,N_19219);
or U20153 (N_20153,N_19442,N_18690);
nor U20154 (N_20154,N_18463,N_18049);
or U20155 (N_20155,N_18836,N_18341);
or U20156 (N_20156,N_19203,N_18780);
or U20157 (N_20157,N_18775,N_18744);
or U20158 (N_20158,N_19470,N_18353);
nor U20159 (N_20159,N_19481,N_18642);
xnor U20160 (N_20160,N_18658,N_18576);
nor U20161 (N_20161,N_18139,N_18675);
xor U20162 (N_20162,N_18958,N_18809);
nand U20163 (N_20163,N_19026,N_18179);
xor U20164 (N_20164,N_19287,N_19426);
xnor U20165 (N_20165,N_18163,N_18540);
nand U20166 (N_20166,N_18037,N_19223);
nand U20167 (N_20167,N_19062,N_18983);
nor U20168 (N_20168,N_19233,N_19488);
or U20169 (N_20169,N_19309,N_19227);
nand U20170 (N_20170,N_18761,N_18046);
and U20171 (N_20171,N_18003,N_19458);
nand U20172 (N_20172,N_18422,N_18587);
xnor U20173 (N_20173,N_18515,N_19213);
nand U20174 (N_20174,N_18822,N_19464);
xor U20175 (N_20175,N_18266,N_19303);
xnor U20176 (N_20176,N_19261,N_18362);
nor U20177 (N_20177,N_19116,N_19413);
nor U20178 (N_20178,N_19145,N_18059);
and U20179 (N_20179,N_19421,N_19066);
and U20180 (N_20180,N_19319,N_19074);
or U20181 (N_20181,N_19054,N_18364);
nand U20182 (N_20182,N_19425,N_19445);
nor U20183 (N_20183,N_18533,N_18188);
and U20184 (N_20184,N_18551,N_18239);
and U20185 (N_20185,N_18565,N_19156);
and U20186 (N_20186,N_18578,N_18395);
xor U20187 (N_20187,N_18088,N_19485);
nand U20188 (N_20188,N_19307,N_18890);
nor U20189 (N_20189,N_19063,N_18247);
or U20190 (N_20190,N_19467,N_18572);
xor U20191 (N_20191,N_18739,N_19468);
nand U20192 (N_20192,N_18525,N_18073);
xnor U20193 (N_20193,N_18424,N_18757);
xor U20194 (N_20194,N_18749,N_18896);
xor U20195 (N_20195,N_18856,N_18400);
and U20196 (N_20196,N_19362,N_19423);
nand U20197 (N_20197,N_19275,N_19273);
nor U20198 (N_20198,N_18256,N_19395);
or U20199 (N_20199,N_18680,N_19224);
or U20200 (N_20200,N_18894,N_19383);
and U20201 (N_20201,N_18298,N_18255);
or U20202 (N_20202,N_18556,N_19254);
nand U20203 (N_20203,N_18317,N_19006);
nand U20204 (N_20204,N_18231,N_18250);
and U20205 (N_20205,N_18994,N_18880);
xnor U20206 (N_20206,N_18027,N_19438);
or U20207 (N_20207,N_18222,N_19078);
or U20208 (N_20208,N_19110,N_18080);
xor U20209 (N_20209,N_18437,N_19197);
or U20210 (N_20210,N_18666,N_19357);
nand U20211 (N_20211,N_18524,N_18745);
and U20212 (N_20212,N_18511,N_18219);
nor U20213 (N_20213,N_18830,N_19479);
or U20214 (N_20214,N_18240,N_19407);
nand U20215 (N_20215,N_18985,N_18420);
nor U20216 (N_20216,N_18473,N_18030);
nor U20217 (N_20217,N_18085,N_18571);
or U20218 (N_20218,N_19264,N_18542);
nor U20219 (N_20219,N_18520,N_19195);
and U20220 (N_20220,N_18408,N_18289);
or U20221 (N_20221,N_19070,N_18866);
and U20222 (N_20222,N_19284,N_18056);
nand U20223 (N_20223,N_18123,N_18474);
and U20224 (N_20224,N_18504,N_18598);
or U20225 (N_20225,N_18101,N_18746);
xor U20226 (N_20226,N_19486,N_19401);
xnor U20227 (N_20227,N_18755,N_18430);
or U20228 (N_20228,N_19388,N_18673);
xnor U20229 (N_20229,N_18491,N_19282);
nor U20230 (N_20230,N_18174,N_18627);
and U20231 (N_20231,N_18564,N_18678);
nor U20232 (N_20232,N_18844,N_18067);
and U20233 (N_20233,N_18557,N_18334);
or U20234 (N_20234,N_18273,N_18965);
nor U20235 (N_20235,N_19448,N_19355);
nand U20236 (N_20236,N_19237,N_18789);
xnor U20237 (N_20237,N_18366,N_18659);
nor U20238 (N_20238,N_19220,N_18224);
or U20239 (N_20239,N_19325,N_18915);
and U20240 (N_20240,N_18909,N_18875);
or U20241 (N_20241,N_19000,N_18284);
xor U20242 (N_20242,N_18308,N_19193);
or U20243 (N_20243,N_18241,N_18397);
nor U20244 (N_20244,N_19023,N_19029);
nand U20245 (N_20245,N_18467,N_19459);
nand U20246 (N_20246,N_18831,N_19440);
nand U20247 (N_20247,N_18258,N_18979);
nor U20248 (N_20248,N_18590,N_18613);
and U20249 (N_20249,N_18061,N_19416);
nor U20250 (N_20250,N_19391,N_19035);
and U20251 (N_20251,N_18763,N_18228);
and U20252 (N_20252,N_19398,N_18808);
nor U20253 (N_20253,N_19252,N_18326);
and U20254 (N_20254,N_18718,N_19022);
xnor U20255 (N_20255,N_18993,N_18016);
or U20256 (N_20256,N_18211,N_18920);
or U20257 (N_20257,N_19177,N_18278);
nor U20258 (N_20258,N_19032,N_19413);
and U20259 (N_20259,N_18793,N_18087);
and U20260 (N_20260,N_18955,N_18075);
xor U20261 (N_20261,N_18389,N_18660);
nor U20262 (N_20262,N_19099,N_19186);
or U20263 (N_20263,N_18702,N_19193);
or U20264 (N_20264,N_19111,N_19044);
or U20265 (N_20265,N_18264,N_19132);
and U20266 (N_20266,N_19450,N_18406);
nor U20267 (N_20267,N_18500,N_18909);
nor U20268 (N_20268,N_19433,N_18870);
and U20269 (N_20269,N_19217,N_18403);
and U20270 (N_20270,N_18774,N_19331);
xor U20271 (N_20271,N_19496,N_18527);
or U20272 (N_20272,N_19022,N_19104);
xnor U20273 (N_20273,N_19400,N_18860);
and U20274 (N_20274,N_18434,N_19321);
xnor U20275 (N_20275,N_19023,N_19020);
or U20276 (N_20276,N_18759,N_18820);
or U20277 (N_20277,N_19290,N_18009);
xnor U20278 (N_20278,N_18023,N_19267);
nor U20279 (N_20279,N_19209,N_19093);
nand U20280 (N_20280,N_18075,N_18523);
or U20281 (N_20281,N_18542,N_18497);
nor U20282 (N_20282,N_18173,N_18372);
xnor U20283 (N_20283,N_18631,N_19132);
xnor U20284 (N_20284,N_18142,N_19175);
or U20285 (N_20285,N_19473,N_18452);
xor U20286 (N_20286,N_18886,N_19227);
nand U20287 (N_20287,N_19094,N_18083);
or U20288 (N_20288,N_19370,N_18711);
nand U20289 (N_20289,N_18107,N_18081);
or U20290 (N_20290,N_18416,N_19131);
nand U20291 (N_20291,N_19493,N_19065);
or U20292 (N_20292,N_18456,N_19060);
xor U20293 (N_20293,N_19072,N_18172);
xor U20294 (N_20294,N_18603,N_18623);
xnor U20295 (N_20295,N_19473,N_18319);
or U20296 (N_20296,N_18786,N_18688);
xor U20297 (N_20297,N_19193,N_19270);
or U20298 (N_20298,N_18319,N_18067);
or U20299 (N_20299,N_18725,N_18538);
and U20300 (N_20300,N_18703,N_19053);
and U20301 (N_20301,N_18836,N_19077);
or U20302 (N_20302,N_18318,N_18087);
or U20303 (N_20303,N_18626,N_18965);
and U20304 (N_20304,N_18925,N_18161);
nand U20305 (N_20305,N_18392,N_18378);
or U20306 (N_20306,N_18105,N_18684);
or U20307 (N_20307,N_18334,N_18918);
nand U20308 (N_20308,N_18187,N_18119);
nand U20309 (N_20309,N_19007,N_18932);
or U20310 (N_20310,N_18256,N_19420);
nor U20311 (N_20311,N_18606,N_18057);
nand U20312 (N_20312,N_18633,N_18379);
nor U20313 (N_20313,N_18569,N_18084);
and U20314 (N_20314,N_18333,N_18940);
or U20315 (N_20315,N_19046,N_18599);
nor U20316 (N_20316,N_19194,N_18236);
xor U20317 (N_20317,N_19014,N_18207);
and U20318 (N_20318,N_18237,N_19463);
and U20319 (N_20319,N_18740,N_19429);
nand U20320 (N_20320,N_19148,N_18322);
nor U20321 (N_20321,N_19468,N_18190);
xnor U20322 (N_20322,N_18817,N_18353);
nor U20323 (N_20323,N_18772,N_18461);
and U20324 (N_20324,N_18345,N_18876);
xor U20325 (N_20325,N_19008,N_19269);
and U20326 (N_20326,N_19140,N_19082);
xor U20327 (N_20327,N_19379,N_18519);
xnor U20328 (N_20328,N_18573,N_18546);
and U20329 (N_20329,N_18727,N_18199);
nor U20330 (N_20330,N_19327,N_19304);
and U20331 (N_20331,N_19264,N_18622);
nand U20332 (N_20332,N_19373,N_18777);
nor U20333 (N_20333,N_18861,N_18543);
xor U20334 (N_20334,N_18066,N_19098);
nor U20335 (N_20335,N_19330,N_18201);
nor U20336 (N_20336,N_18666,N_18296);
nor U20337 (N_20337,N_18495,N_18832);
nor U20338 (N_20338,N_19403,N_19057);
nand U20339 (N_20339,N_19049,N_19027);
nor U20340 (N_20340,N_18575,N_19470);
xor U20341 (N_20341,N_18979,N_18513);
xor U20342 (N_20342,N_18242,N_18498);
nor U20343 (N_20343,N_18029,N_19476);
nand U20344 (N_20344,N_18278,N_18939);
or U20345 (N_20345,N_18604,N_18152);
nor U20346 (N_20346,N_18734,N_18831);
or U20347 (N_20347,N_18410,N_18562);
xnor U20348 (N_20348,N_19077,N_18679);
nor U20349 (N_20349,N_19118,N_18723);
xor U20350 (N_20350,N_19186,N_19441);
and U20351 (N_20351,N_19414,N_18277);
or U20352 (N_20352,N_18149,N_18895);
and U20353 (N_20353,N_18833,N_19489);
xor U20354 (N_20354,N_18747,N_18489);
nor U20355 (N_20355,N_18646,N_18358);
xnor U20356 (N_20356,N_19142,N_19202);
nor U20357 (N_20357,N_18951,N_19297);
nand U20358 (N_20358,N_19256,N_19060);
and U20359 (N_20359,N_18558,N_19017);
or U20360 (N_20360,N_18321,N_19149);
xor U20361 (N_20361,N_19429,N_18605);
xor U20362 (N_20362,N_18779,N_19218);
nand U20363 (N_20363,N_19283,N_18742);
nor U20364 (N_20364,N_18856,N_18159);
nand U20365 (N_20365,N_19464,N_18511);
and U20366 (N_20366,N_18726,N_18276);
or U20367 (N_20367,N_18641,N_18177);
nor U20368 (N_20368,N_19448,N_18451);
and U20369 (N_20369,N_19032,N_18760);
xnor U20370 (N_20370,N_18444,N_18148);
nand U20371 (N_20371,N_19223,N_19274);
or U20372 (N_20372,N_18226,N_18961);
and U20373 (N_20373,N_19006,N_19220);
and U20374 (N_20374,N_18102,N_19340);
and U20375 (N_20375,N_18296,N_19489);
and U20376 (N_20376,N_19041,N_19090);
xnor U20377 (N_20377,N_18651,N_18853);
or U20378 (N_20378,N_18962,N_19073);
xor U20379 (N_20379,N_18617,N_18695);
and U20380 (N_20380,N_19090,N_19136);
or U20381 (N_20381,N_19315,N_18453);
xor U20382 (N_20382,N_18477,N_18580);
xor U20383 (N_20383,N_19002,N_19084);
nand U20384 (N_20384,N_18342,N_18339);
or U20385 (N_20385,N_19428,N_18599);
and U20386 (N_20386,N_18115,N_18500);
and U20387 (N_20387,N_18637,N_19044);
xor U20388 (N_20388,N_18489,N_18483);
and U20389 (N_20389,N_19155,N_18434);
and U20390 (N_20390,N_18893,N_18294);
nand U20391 (N_20391,N_18924,N_19211);
or U20392 (N_20392,N_18770,N_18923);
and U20393 (N_20393,N_19362,N_18646);
and U20394 (N_20394,N_18534,N_18126);
nor U20395 (N_20395,N_19055,N_18951);
and U20396 (N_20396,N_18052,N_19343);
or U20397 (N_20397,N_19094,N_18633);
xnor U20398 (N_20398,N_18716,N_18873);
nor U20399 (N_20399,N_18397,N_18815);
xor U20400 (N_20400,N_18469,N_19093);
and U20401 (N_20401,N_18546,N_18345);
or U20402 (N_20402,N_18354,N_18525);
or U20403 (N_20403,N_18243,N_18526);
xor U20404 (N_20404,N_18483,N_19125);
nor U20405 (N_20405,N_18288,N_19144);
nand U20406 (N_20406,N_18210,N_19402);
xor U20407 (N_20407,N_19033,N_19357);
nand U20408 (N_20408,N_18703,N_19267);
and U20409 (N_20409,N_18246,N_18168);
and U20410 (N_20410,N_19482,N_18942);
or U20411 (N_20411,N_18923,N_19032);
and U20412 (N_20412,N_19240,N_18689);
nand U20413 (N_20413,N_18375,N_18112);
or U20414 (N_20414,N_18668,N_19063);
and U20415 (N_20415,N_19418,N_18555);
and U20416 (N_20416,N_18439,N_18426);
and U20417 (N_20417,N_19445,N_18406);
nor U20418 (N_20418,N_18115,N_19460);
or U20419 (N_20419,N_19112,N_19141);
and U20420 (N_20420,N_18786,N_18938);
nand U20421 (N_20421,N_18626,N_19013);
and U20422 (N_20422,N_18458,N_19484);
xnor U20423 (N_20423,N_18156,N_18870);
or U20424 (N_20424,N_18309,N_18305);
nor U20425 (N_20425,N_19315,N_19011);
or U20426 (N_20426,N_18767,N_19399);
or U20427 (N_20427,N_19218,N_19250);
xor U20428 (N_20428,N_18887,N_18822);
xnor U20429 (N_20429,N_18476,N_18456);
and U20430 (N_20430,N_19462,N_18290);
nand U20431 (N_20431,N_18585,N_18075);
nor U20432 (N_20432,N_18286,N_18581);
and U20433 (N_20433,N_18042,N_18697);
nand U20434 (N_20434,N_18081,N_18574);
nor U20435 (N_20435,N_18401,N_18728);
or U20436 (N_20436,N_18997,N_18680);
nor U20437 (N_20437,N_18117,N_18601);
and U20438 (N_20438,N_19152,N_18664);
xor U20439 (N_20439,N_19453,N_19030);
nand U20440 (N_20440,N_19295,N_18845);
and U20441 (N_20441,N_18561,N_18099);
and U20442 (N_20442,N_18389,N_18371);
nand U20443 (N_20443,N_18364,N_19384);
nand U20444 (N_20444,N_18143,N_18373);
xor U20445 (N_20445,N_18461,N_18952);
or U20446 (N_20446,N_18178,N_18323);
and U20447 (N_20447,N_18436,N_18468);
nand U20448 (N_20448,N_18374,N_19242);
and U20449 (N_20449,N_19153,N_18718);
and U20450 (N_20450,N_19237,N_19383);
xor U20451 (N_20451,N_18266,N_18283);
nor U20452 (N_20452,N_18538,N_19194);
nor U20453 (N_20453,N_18190,N_18202);
or U20454 (N_20454,N_19116,N_18457);
nor U20455 (N_20455,N_18103,N_18238);
or U20456 (N_20456,N_18800,N_19423);
xor U20457 (N_20457,N_18916,N_18959);
or U20458 (N_20458,N_19081,N_18852);
and U20459 (N_20459,N_19051,N_18577);
and U20460 (N_20460,N_18710,N_19222);
xor U20461 (N_20461,N_18975,N_19366);
or U20462 (N_20462,N_18747,N_19451);
xor U20463 (N_20463,N_18149,N_18394);
or U20464 (N_20464,N_18414,N_19397);
nor U20465 (N_20465,N_19017,N_18463);
and U20466 (N_20466,N_18932,N_18033);
or U20467 (N_20467,N_19325,N_19476);
nand U20468 (N_20468,N_18483,N_18327);
nor U20469 (N_20469,N_18457,N_18820);
and U20470 (N_20470,N_19377,N_18156);
nor U20471 (N_20471,N_18181,N_18169);
xnor U20472 (N_20472,N_18665,N_18089);
or U20473 (N_20473,N_19228,N_18768);
nor U20474 (N_20474,N_18659,N_18714);
nor U20475 (N_20475,N_19346,N_19307);
nand U20476 (N_20476,N_18219,N_18834);
nor U20477 (N_20477,N_18377,N_18809);
or U20478 (N_20478,N_18750,N_18927);
and U20479 (N_20479,N_19108,N_19082);
nand U20480 (N_20480,N_18512,N_19126);
nand U20481 (N_20481,N_18716,N_18998);
nor U20482 (N_20482,N_18235,N_19373);
xnor U20483 (N_20483,N_18460,N_18511);
xnor U20484 (N_20484,N_18910,N_18915);
or U20485 (N_20485,N_18698,N_19431);
nand U20486 (N_20486,N_19316,N_19414);
or U20487 (N_20487,N_18462,N_18975);
xnor U20488 (N_20488,N_19274,N_18434);
nand U20489 (N_20489,N_18748,N_19388);
nand U20490 (N_20490,N_19337,N_18857);
and U20491 (N_20491,N_18137,N_18140);
nor U20492 (N_20492,N_18979,N_19245);
nand U20493 (N_20493,N_18681,N_19298);
and U20494 (N_20494,N_19134,N_19073);
nor U20495 (N_20495,N_19381,N_19067);
or U20496 (N_20496,N_18774,N_19432);
nor U20497 (N_20497,N_19231,N_19384);
nand U20498 (N_20498,N_18153,N_18019);
nor U20499 (N_20499,N_19056,N_18071);
and U20500 (N_20500,N_18307,N_18379);
nor U20501 (N_20501,N_19419,N_18127);
nand U20502 (N_20502,N_18892,N_18037);
xor U20503 (N_20503,N_18154,N_19182);
nand U20504 (N_20504,N_18330,N_19413);
nor U20505 (N_20505,N_18583,N_18075);
or U20506 (N_20506,N_19037,N_18393);
nor U20507 (N_20507,N_19035,N_18818);
nor U20508 (N_20508,N_19432,N_19382);
and U20509 (N_20509,N_18423,N_18738);
and U20510 (N_20510,N_18588,N_18296);
nor U20511 (N_20511,N_18255,N_18437);
or U20512 (N_20512,N_18787,N_18829);
or U20513 (N_20513,N_18732,N_18399);
xnor U20514 (N_20514,N_19404,N_18160);
nor U20515 (N_20515,N_18436,N_18214);
nor U20516 (N_20516,N_18256,N_18102);
nor U20517 (N_20517,N_19184,N_18719);
nor U20518 (N_20518,N_18359,N_18394);
or U20519 (N_20519,N_18733,N_18969);
xor U20520 (N_20520,N_18800,N_18280);
nor U20521 (N_20521,N_18337,N_18463);
nor U20522 (N_20522,N_18515,N_18703);
nand U20523 (N_20523,N_18774,N_18863);
and U20524 (N_20524,N_18863,N_18595);
nand U20525 (N_20525,N_19042,N_18420);
xor U20526 (N_20526,N_19350,N_19391);
nor U20527 (N_20527,N_19210,N_18670);
nand U20528 (N_20528,N_18685,N_18378);
or U20529 (N_20529,N_18388,N_18716);
and U20530 (N_20530,N_19242,N_18767);
nand U20531 (N_20531,N_18338,N_18234);
and U20532 (N_20532,N_18960,N_19075);
nand U20533 (N_20533,N_18403,N_18916);
or U20534 (N_20534,N_19163,N_18888);
or U20535 (N_20535,N_18733,N_19076);
xnor U20536 (N_20536,N_19065,N_18011);
nor U20537 (N_20537,N_18419,N_18728);
nand U20538 (N_20538,N_19284,N_18074);
and U20539 (N_20539,N_18174,N_18345);
nor U20540 (N_20540,N_18042,N_19185);
or U20541 (N_20541,N_19174,N_18099);
and U20542 (N_20542,N_18647,N_18283);
nand U20543 (N_20543,N_18250,N_18881);
nor U20544 (N_20544,N_18950,N_18324);
nand U20545 (N_20545,N_19343,N_19275);
nor U20546 (N_20546,N_18438,N_19089);
xor U20547 (N_20547,N_18878,N_18973);
or U20548 (N_20548,N_18420,N_19189);
or U20549 (N_20549,N_18726,N_18451);
xor U20550 (N_20550,N_19165,N_18595);
nand U20551 (N_20551,N_18218,N_19146);
nand U20552 (N_20552,N_19176,N_18984);
nand U20553 (N_20553,N_18646,N_19498);
or U20554 (N_20554,N_19186,N_18603);
and U20555 (N_20555,N_19444,N_19034);
xnor U20556 (N_20556,N_18064,N_19299);
or U20557 (N_20557,N_18865,N_19204);
nor U20558 (N_20558,N_18461,N_18904);
and U20559 (N_20559,N_18382,N_19026);
nor U20560 (N_20560,N_18910,N_19002);
nor U20561 (N_20561,N_18017,N_19003);
nor U20562 (N_20562,N_19403,N_18580);
nor U20563 (N_20563,N_18592,N_19254);
and U20564 (N_20564,N_18865,N_19282);
nand U20565 (N_20565,N_18418,N_19075);
xnor U20566 (N_20566,N_18108,N_18589);
or U20567 (N_20567,N_19378,N_19024);
nor U20568 (N_20568,N_19433,N_18506);
or U20569 (N_20569,N_19387,N_18088);
and U20570 (N_20570,N_18825,N_19449);
nor U20571 (N_20571,N_19199,N_18222);
nor U20572 (N_20572,N_19066,N_18485);
or U20573 (N_20573,N_18748,N_19292);
nor U20574 (N_20574,N_18495,N_18344);
nand U20575 (N_20575,N_18615,N_19269);
and U20576 (N_20576,N_18280,N_18817);
or U20577 (N_20577,N_18560,N_18704);
or U20578 (N_20578,N_19097,N_18435);
xnor U20579 (N_20579,N_18779,N_18878);
or U20580 (N_20580,N_18493,N_18499);
or U20581 (N_20581,N_18528,N_18907);
and U20582 (N_20582,N_18239,N_18856);
nand U20583 (N_20583,N_18030,N_18761);
and U20584 (N_20584,N_18247,N_18304);
and U20585 (N_20585,N_19418,N_19154);
xor U20586 (N_20586,N_19321,N_18140);
nand U20587 (N_20587,N_18106,N_19169);
and U20588 (N_20588,N_18940,N_18513);
and U20589 (N_20589,N_18006,N_18567);
nor U20590 (N_20590,N_18735,N_18413);
nand U20591 (N_20591,N_18355,N_19464);
or U20592 (N_20592,N_18651,N_19213);
nand U20593 (N_20593,N_18274,N_19470);
or U20594 (N_20594,N_18277,N_18265);
xor U20595 (N_20595,N_18167,N_18315);
and U20596 (N_20596,N_18998,N_18139);
nand U20597 (N_20597,N_18445,N_19205);
nand U20598 (N_20598,N_19117,N_18790);
and U20599 (N_20599,N_18722,N_18728);
and U20600 (N_20600,N_18425,N_19223);
or U20601 (N_20601,N_18150,N_18479);
xor U20602 (N_20602,N_18139,N_18292);
nand U20603 (N_20603,N_19176,N_19394);
or U20604 (N_20604,N_19084,N_19214);
and U20605 (N_20605,N_18153,N_18447);
and U20606 (N_20606,N_19031,N_18165);
xor U20607 (N_20607,N_19220,N_18799);
nor U20608 (N_20608,N_18367,N_18118);
nand U20609 (N_20609,N_19445,N_18269);
or U20610 (N_20610,N_18993,N_18918);
nor U20611 (N_20611,N_19203,N_18738);
nor U20612 (N_20612,N_19052,N_19492);
nor U20613 (N_20613,N_19031,N_19113);
nor U20614 (N_20614,N_18056,N_18609);
and U20615 (N_20615,N_18567,N_19361);
xnor U20616 (N_20616,N_18189,N_18007);
nor U20617 (N_20617,N_19293,N_18751);
nor U20618 (N_20618,N_18341,N_18251);
nor U20619 (N_20619,N_18750,N_18707);
nor U20620 (N_20620,N_18948,N_18931);
nor U20621 (N_20621,N_18059,N_19031);
nor U20622 (N_20622,N_18187,N_19079);
and U20623 (N_20623,N_18820,N_18523);
nor U20624 (N_20624,N_18113,N_18076);
and U20625 (N_20625,N_18660,N_18925);
and U20626 (N_20626,N_19247,N_19055);
and U20627 (N_20627,N_18762,N_18281);
and U20628 (N_20628,N_19487,N_18513);
or U20629 (N_20629,N_18942,N_19442);
nor U20630 (N_20630,N_18464,N_19187);
nor U20631 (N_20631,N_18267,N_18401);
nand U20632 (N_20632,N_18620,N_19499);
nand U20633 (N_20633,N_18272,N_18348);
or U20634 (N_20634,N_18275,N_19329);
nand U20635 (N_20635,N_18902,N_18320);
or U20636 (N_20636,N_19467,N_18709);
and U20637 (N_20637,N_19251,N_18104);
xnor U20638 (N_20638,N_18259,N_18565);
nand U20639 (N_20639,N_18239,N_18797);
or U20640 (N_20640,N_18799,N_18384);
and U20641 (N_20641,N_18485,N_18569);
nor U20642 (N_20642,N_19380,N_18889);
or U20643 (N_20643,N_18451,N_19146);
nand U20644 (N_20644,N_18863,N_18348);
xor U20645 (N_20645,N_19098,N_19056);
and U20646 (N_20646,N_18705,N_18647);
and U20647 (N_20647,N_18122,N_18766);
nand U20648 (N_20648,N_19288,N_18841);
or U20649 (N_20649,N_19421,N_18697);
nand U20650 (N_20650,N_18967,N_18652);
or U20651 (N_20651,N_18748,N_19483);
nor U20652 (N_20652,N_19248,N_18639);
nor U20653 (N_20653,N_18148,N_18166);
and U20654 (N_20654,N_19126,N_18589);
nand U20655 (N_20655,N_18635,N_18651);
and U20656 (N_20656,N_18383,N_18032);
and U20657 (N_20657,N_19189,N_18682);
or U20658 (N_20658,N_18497,N_19279);
or U20659 (N_20659,N_18372,N_18753);
nor U20660 (N_20660,N_19079,N_18229);
nand U20661 (N_20661,N_18831,N_19199);
xnor U20662 (N_20662,N_19260,N_19336);
nor U20663 (N_20663,N_18029,N_18986);
nor U20664 (N_20664,N_19020,N_18686);
nor U20665 (N_20665,N_18333,N_18789);
nand U20666 (N_20666,N_18679,N_18173);
or U20667 (N_20667,N_18212,N_18845);
xnor U20668 (N_20668,N_18661,N_18560);
nand U20669 (N_20669,N_18624,N_18580);
and U20670 (N_20670,N_19456,N_19312);
xor U20671 (N_20671,N_18444,N_18830);
and U20672 (N_20672,N_19198,N_18508);
nand U20673 (N_20673,N_19414,N_19470);
xnor U20674 (N_20674,N_19019,N_18768);
or U20675 (N_20675,N_18847,N_18057);
nor U20676 (N_20676,N_18822,N_18939);
or U20677 (N_20677,N_18341,N_18293);
nor U20678 (N_20678,N_18276,N_18172);
nand U20679 (N_20679,N_18941,N_19065);
and U20680 (N_20680,N_18200,N_18056);
nor U20681 (N_20681,N_18234,N_19210);
and U20682 (N_20682,N_18825,N_18004);
nand U20683 (N_20683,N_19229,N_18078);
nand U20684 (N_20684,N_19368,N_19121);
nand U20685 (N_20685,N_18920,N_18473);
and U20686 (N_20686,N_18968,N_18382);
nor U20687 (N_20687,N_19344,N_18582);
and U20688 (N_20688,N_19399,N_19342);
nor U20689 (N_20689,N_18376,N_18370);
xor U20690 (N_20690,N_19106,N_18944);
or U20691 (N_20691,N_18091,N_19397);
or U20692 (N_20692,N_18172,N_18604);
xnor U20693 (N_20693,N_18223,N_18969);
nand U20694 (N_20694,N_19000,N_19408);
xnor U20695 (N_20695,N_18429,N_19212);
nand U20696 (N_20696,N_19177,N_19072);
and U20697 (N_20697,N_19184,N_18353);
xor U20698 (N_20698,N_18451,N_18715);
or U20699 (N_20699,N_18823,N_18988);
nand U20700 (N_20700,N_18362,N_18399);
nor U20701 (N_20701,N_18828,N_18496);
nor U20702 (N_20702,N_18763,N_18695);
xor U20703 (N_20703,N_18870,N_19127);
nor U20704 (N_20704,N_18687,N_18770);
nor U20705 (N_20705,N_19173,N_18070);
nor U20706 (N_20706,N_18623,N_19077);
or U20707 (N_20707,N_19117,N_18939);
or U20708 (N_20708,N_19202,N_18546);
xor U20709 (N_20709,N_18120,N_19062);
nand U20710 (N_20710,N_18024,N_19118);
nand U20711 (N_20711,N_19016,N_19359);
nand U20712 (N_20712,N_18841,N_18455);
nor U20713 (N_20713,N_18038,N_19295);
xnor U20714 (N_20714,N_18474,N_18957);
nand U20715 (N_20715,N_18126,N_19057);
nor U20716 (N_20716,N_18079,N_18981);
nor U20717 (N_20717,N_18615,N_18652);
or U20718 (N_20718,N_18408,N_19328);
nor U20719 (N_20719,N_18373,N_19209);
nand U20720 (N_20720,N_18145,N_19082);
or U20721 (N_20721,N_18555,N_18111);
or U20722 (N_20722,N_18732,N_18253);
and U20723 (N_20723,N_18754,N_18657);
and U20724 (N_20724,N_18532,N_19177);
xnor U20725 (N_20725,N_18716,N_18914);
and U20726 (N_20726,N_18976,N_18958);
and U20727 (N_20727,N_18502,N_18574);
nand U20728 (N_20728,N_18149,N_18034);
or U20729 (N_20729,N_18248,N_18111);
xnor U20730 (N_20730,N_18872,N_18997);
and U20731 (N_20731,N_18643,N_18981);
nor U20732 (N_20732,N_18791,N_18439);
nand U20733 (N_20733,N_18775,N_19238);
or U20734 (N_20734,N_19018,N_19081);
nor U20735 (N_20735,N_19453,N_19386);
and U20736 (N_20736,N_19240,N_18788);
nor U20737 (N_20737,N_18505,N_18150);
nand U20738 (N_20738,N_18336,N_18767);
xor U20739 (N_20739,N_18313,N_18168);
xor U20740 (N_20740,N_18107,N_18193);
or U20741 (N_20741,N_19128,N_18307);
xnor U20742 (N_20742,N_18223,N_18503);
nand U20743 (N_20743,N_19375,N_19179);
and U20744 (N_20744,N_18498,N_18130);
or U20745 (N_20745,N_18495,N_19399);
or U20746 (N_20746,N_18726,N_19142);
or U20747 (N_20747,N_18412,N_18238);
xnor U20748 (N_20748,N_18236,N_18176);
xor U20749 (N_20749,N_18760,N_19232);
or U20750 (N_20750,N_18372,N_19235);
xnor U20751 (N_20751,N_19180,N_18872);
nand U20752 (N_20752,N_18303,N_19121);
and U20753 (N_20753,N_18968,N_18992);
nor U20754 (N_20754,N_19112,N_18925);
and U20755 (N_20755,N_18527,N_18446);
or U20756 (N_20756,N_18963,N_19225);
nor U20757 (N_20757,N_19113,N_19017);
and U20758 (N_20758,N_18502,N_19003);
xor U20759 (N_20759,N_18180,N_19485);
nor U20760 (N_20760,N_18976,N_18706);
nor U20761 (N_20761,N_18116,N_18504);
and U20762 (N_20762,N_19251,N_18621);
xnor U20763 (N_20763,N_19420,N_19276);
nand U20764 (N_20764,N_19137,N_18806);
or U20765 (N_20765,N_18291,N_19002);
and U20766 (N_20766,N_18172,N_18098);
xnor U20767 (N_20767,N_18628,N_18843);
xor U20768 (N_20768,N_18270,N_18451);
and U20769 (N_20769,N_19484,N_19377);
nand U20770 (N_20770,N_18951,N_18270);
and U20771 (N_20771,N_19494,N_19440);
nand U20772 (N_20772,N_18097,N_18301);
and U20773 (N_20773,N_19306,N_18934);
nand U20774 (N_20774,N_18096,N_19499);
and U20775 (N_20775,N_18853,N_18011);
and U20776 (N_20776,N_18277,N_18420);
xnor U20777 (N_20777,N_18251,N_19342);
and U20778 (N_20778,N_18863,N_18068);
and U20779 (N_20779,N_19300,N_18049);
and U20780 (N_20780,N_18826,N_18110);
xor U20781 (N_20781,N_19315,N_18854);
or U20782 (N_20782,N_19208,N_19450);
and U20783 (N_20783,N_19427,N_18093);
and U20784 (N_20784,N_18685,N_18151);
xor U20785 (N_20785,N_18703,N_18524);
or U20786 (N_20786,N_18335,N_18110);
or U20787 (N_20787,N_18431,N_19096);
xnor U20788 (N_20788,N_18730,N_19444);
or U20789 (N_20789,N_19446,N_18086);
and U20790 (N_20790,N_18266,N_19092);
or U20791 (N_20791,N_19060,N_19086);
nand U20792 (N_20792,N_18117,N_19224);
xor U20793 (N_20793,N_19473,N_18691);
xnor U20794 (N_20794,N_18879,N_18935);
and U20795 (N_20795,N_19034,N_18792);
nor U20796 (N_20796,N_18970,N_18574);
nand U20797 (N_20797,N_18704,N_18901);
or U20798 (N_20798,N_18055,N_19380);
and U20799 (N_20799,N_19382,N_18036);
or U20800 (N_20800,N_18570,N_18845);
or U20801 (N_20801,N_19116,N_18351);
or U20802 (N_20802,N_18435,N_18402);
and U20803 (N_20803,N_19003,N_18616);
or U20804 (N_20804,N_18521,N_19448);
nand U20805 (N_20805,N_18066,N_19377);
xor U20806 (N_20806,N_18173,N_19041);
or U20807 (N_20807,N_18732,N_18067);
and U20808 (N_20808,N_19306,N_18593);
nor U20809 (N_20809,N_19217,N_18041);
and U20810 (N_20810,N_18521,N_18993);
nand U20811 (N_20811,N_18188,N_18112);
xnor U20812 (N_20812,N_18184,N_19327);
xor U20813 (N_20813,N_18364,N_19366);
nand U20814 (N_20814,N_18028,N_18338);
nand U20815 (N_20815,N_18103,N_19191);
nor U20816 (N_20816,N_19353,N_18843);
nor U20817 (N_20817,N_18904,N_18561);
nand U20818 (N_20818,N_18888,N_18243);
or U20819 (N_20819,N_18967,N_19047);
or U20820 (N_20820,N_18661,N_18462);
nand U20821 (N_20821,N_18030,N_18211);
xnor U20822 (N_20822,N_18207,N_18674);
nor U20823 (N_20823,N_19126,N_18243);
xor U20824 (N_20824,N_18661,N_19173);
xor U20825 (N_20825,N_18505,N_18803);
or U20826 (N_20826,N_19058,N_19104);
and U20827 (N_20827,N_18853,N_18481);
nand U20828 (N_20828,N_19368,N_18946);
and U20829 (N_20829,N_18302,N_19150);
nor U20830 (N_20830,N_18177,N_18052);
and U20831 (N_20831,N_19046,N_18357);
nor U20832 (N_20832,N_19000,N_19303);
nand U20833 (N_20833,N_19395,N_19142);
or U20834 (N_20834,N_19328,N_18886);
and U20835 (N_20835,N_18783,N_19256);
or U20836 (N_20836,N_18955,N_18290);
nand U20837 (N_20837,N_18163,N_18274);
and U20838 (N_20838,N_18266,N_18896);
or U20839 (N_20839,N_19094,N_18168);
or U20840 (N_20840,N_18509,N_18807);
and U20841 (N_20841,N_19235,N_19374);
and U20842 (N_20842,N_18527,N_18053);
or U20843 (N_20843,N_18587,N_18631);
and U20844 (N_20844,N_18018,N_18249);
nor U20845 (N_20845,N_18886,N_19125);
nor U20846 (N_20846,N_19026,N_18892);
nor U20847 (N_20847,N_19227,N_19494);
or U20848 (N_20848,N_18252,N_18771);
or U20849 (N_20849,N_19353,N_18658);
xor U20850 (N_20850,N_19160,N_19123);
nor U20851 (N_20851,N_18990,N_18504);
and U20852 (N_20852,N_19466,N_18409);
nor U20853 (N_20853,N_18912,N_18263);
nand U20854 (N_20854,N_19496,N_18391);
xnor U20855 (N_20855,N_18158,N_18434);
nor U20856 (N_20856,N_18425,N_18845);
nand U20857 (N_20857,N_19289,N_18010);
nor U20858 (N_20858,N_18034,N_18602);
or U20859 (N_20859,N_19037,N_18431);
or U20860 (N_20860,N_18368,N_18393);
or U20861 (N_20861,N_18288,N_18231);
nor U20862 (N_20862,N_19388,N_18026);
and U20863 (N_20863,N_18243,N_18055);
nor U20864 (N_20864,N_18285,N_19012);
or U20865 (N_20865,N_19313,N_18571);
xor U20866 (N_20866,N_19454,N_18485);
or U20867 (N_20867,N_18405,N_18284);
xnor U20868 (N_20868,N_19281,N_18937);
and U20869 (N_20869,N_19182,N_19310);
nand U20870 (N_20870,N_19207,N_18443);
or U20871 (N_20871,N_19264,N_18690);
nand U20872 (N_20872,N_18153,N_18427);
nor U20873 (N_20873,N_19107,N_19220);
or U20874 (N_20874,N_18721,N_18141);
xor U20875 (N_20875,N_18606,N_19459);
nor U20876 (N_20876,N_19252,N_19257);
nor U20877 (N_20877,N_19245,N_18296);
xor U20878 (N_20878,N_18587,N_19224);
xor U20879 (N_20879,N_18863,N_18732);
xor U20880 (N_20880,N_18605,N_18640);
or U20881 (N_20881,N_19182,N_19027);
or U20882 (N_20882,N_19247,N_18342);
and U20883 (N_20883,N_18427,N_19124);
and U20884 (N_20884,N_18693,N_18119);
nand U20885 (N_20885,N_18978,N_18525);
nand U20886 (N_20886,N_18075,N_19282);
or U20887 (N_20887,N_18162,N_18036);
or U20888 (N_20888,N_19329,N_18357);
nand U20889 (N_20889,N_18051,N_18572);
nor U20890 (N_20890,N_19140,N_18839);
nor U20891 (N_20891,N_18502,N_18229);
nor U20892 (N_20892,N_19117,N_18090);
nand U20893 (N_20893,N_18677,N_18778);
nand U20894 (N_20894,N_19019,N_18522);
xnor U20895 (N_20895,N_18079,N_18326);
nand U20896 (N_20896,N_18197,N_19350);
nor U20897 (N_20897,N_18185,N_18278);
or U20898 (N_20898,N_19126,N_18165);
nor U20899 (N_20899,N_19258,N_18305);
nor U20900 (N_20900,N_19081,N_19073);
nand U20901 (N_20901,N_18816,N_18576);
and U20902 (N_20902,N_18970,N_19043);
nor U20903 (N_20903,N_18437,N_18724);
xnor U20904 (N_20904,N_19096,N_18085);
xnor U20905 (N_20905,N_18959,N_18118);
xor U20906 (N_20906,N_18659,N_18395);
or U20907 (N_20907,N_18973,N_19332);
nand U20908 (N_20908,N_18007,N_18863);
or U20909 (N_20909,N_18910,N_18120);
xnor U20910 (N_20910,N_18337,N_18333);
nand U20911 (N_20911,N_18880,N_18011);
xor U20912 (N_20912,N_18084,N_18272);
nor U20913 (N_20913,N_18052,N_18989);
nor U20914 (N_20914,N_19126,N_19282);
and U20915 (N_20915,N_18385,N_18706);
xnor U20916 (N_20916,N_18085,N_19145);
nor U20917 (N_20917,N_18870,N_18627);
nor U20918 (N_20918,N_18118,N_19188);
or U20919 (N_20919,N_18158,N_19497);
nor U20920 (N_20920,N_18505,N_19437);
nor U20921 (N_20921,N_18434,N_18557);
or U20922 (N_20922,N_18374,N_18700);
xnor U20923 (N_20923,N_18093,N_18815);
nor U20924 (N_20924,N_18496,N_18939);
nor U20925 (N_20925,N_18093,N_18899);
and U20926 (N_20926,N_19434,N_18449);
nand U20927 (N_20927,N_19243,N_18087);
nor U20928 (N_20928,N_18769,N_18360);
nand U20929 (N_20929,N_18148,N_19492);
nand U20930 (N_20930,N_18810,N_18654);
nand U20931 (N_20931,N_19011,N_19303);
nand U20932 (N_20932,N_18433,N_18473);
and U20933 (N_20933,N_18111,N_18521);
and U20934 (N_20934,N_18290,N_18989);
or U20935 (N_20935,N_19114,N_18822);
or U20936 (N_20936,N_18982,N_18732);
nor U20937 (N_20937,N_19076,N_18984);
or U20938 (N_20938,N_18763,N_18302);
and U20939 (N_20939,N_18007,N_18239);
nor U20940 (N_20940,N_18298,N_19254);
nand U20941 (N_20941,N_18515,N_18357);
nand U20942 (N_20942,N_19071,N_19192);
or U20943 (N_20943,N_18116,N_19038);
xnor U20944 (N_20944,N_18595,N_18111);
xor U20945 (N_20945,N_18778,N_18619);
and U20946 (N_20946,N_18407,N_19184);
or U20947 (N_20947,N_18360,N_18484);
nand U20948 (N_20948,N_18982,N_18929);
and U20949 (N_20949,N_18073,N_19141);
and U20950 (N_20950,N_18731,N_19133);
and U20951 (N_20951,N_19390,N_18669);
nor U20952 (N_20952,N_18484,N_18954);
xnor U20953 (N_20953,N_18228,N_18599);
and U20954 (N_20954,N_19405,N_18486);
nand U20955 (N_20955,N_19275,N_19123);
or U20956 (N_20956,N_18989,N_18510);
or U20957 (N_20957,N_18771,N_18266);
xor U20958 (N_20958,N_19353,N_18737);
or U20959 (N_20959,N_18517,N_18935);
nor U20960 (N_20960,N_19265,N_18112);
nor U20961 (N_20961,N_18708,N_18755);
or U20962 (N_20962,N_18526,N_18303);
nor U20963 (N_20963,N_18857,N_18968);
xor U20964 (N_20964,N_19005,N_19229);
and U20965 (N_20965,N_18974,N_18228);
nand U20966 (N_20966,N_18027,N_18357);
xor U20967 (N_20967,N_18721,N_19205);
and U20968 (N_20968,N_19011,N_18014);
nand U20969 (N_20969,N_18122,N_18878);
and U20970 (N_20970,N_19163,N_19125);
nor U20971 (N_20971,N_18734,N_18731);
and U20972 (N_20972,N_18193,N_18764);
and U20973 (N_20973,N_18334,N_19239);
xor U20974 (N_20974,N_19143,N_18687);
xor U20975 (N_20975,N_18962,N_18745);
and U20976 (N_20976,N_19188,N_18093);
nand U20977 (N_20977,N_18237,N_18861);
nor U20978 (N_20978,N_18440,N_18423);
or U20979 (N_20979,N_19072,N_19275);
and U20980 (N_20980,N_18024,N_18211);
nand U20981 (N_20981,N_18106,N_18979);
or U20982 (N_20982,N_18594,N_18616);
nor U20983 (N_20983,N_19134,N_19081);
or U20984 (N_20984,N_18818,N_18112);
nor U20985 (N_20985,N_19133,N_18624);
nand U20986 (N_20986,N_18336,N_18513);
nand U20987 (N_20987,N_18395,N_18061);
or U20988 (N_20988,N_19280,N_18116);
nand U20989 (N_20989,N_18794,N_19408);
and U20990 (N_20990,N_19426,N_18890);
and U20991 (N_20991,N_19367,N_18044);
nand U20992 (N_20992,N_18337,N_18559);
nor U20993 (N_20993,N_18352,N_19198);
or U20994 (N_20994,N_18030,N_18304);
or U20995 (N_20995,N_18271,N_19326);
and U20996 (N_20996,N_18644,N_19117);
xnor U20997 (N_20997,N_18982,N_18762);
or U20998 (N_20998,N_19452,N_18001);
nor U20999 (N_20999,N_18946,N_18598);
and U21000 (N_21000,N_20113,N_20044);
nand U21001 (N_21001,N_19652,N_20832);
nor U21002 (N_21002,N_19702,N_20345);
xnor U21003 (N_21003,N_20813,N_19798);
and U21004 (N_21004,N_19946,N_20790);
or U21005 (N_21005,N_19691,N_20673);
and U21006 (N_21006,N_20851,N_19500);
or U21007 (N_21007,N_20326,N_20491);
xnor U21008 (N_21008,N_20346,N_20939);
nand U21009 (N_21009,N_20074,N_20481);
nand U21010 (N_21010,N_19986,N_20511);
or U21011 (N_21011,N_20718,N_19918);
nand U21012 (N_21012,N_19952,N_20138);
or U21013 (N_21013,N_20947,N_20331);
or U21014 (N_21014,N_20150,N_20707);
nand U21015 (N_21015,N_20556,N_19516);
or U21016 (N_21016,N_20602,N_19988);
or U21017 (N_21017,N_20353,N_20770);
or U21018 (N_21018,N_20911,N_19842);
nand U21019 (N_21019,N_20065,N_19616);
or U21020 (N_21020,N_20985,N_20221);
or U21021 (N_21021,N_20862,N_20394);
and U21022 (N_21022,N_20266,N_19885);
nor U21023 (N_21023,N_20184,N_20217);
or U21024 (N_21024,N_20822,N_19751);
and U21025 (N_21025,N_20685,N_20139);
xnor U21026 (N_21026,N_20769,N_20493);
xnor U21027 (N_21027,N_20425,N_20523);
xnor U21028 (N_21028,N_19852,N_20350);
xnor U21029 (N_21029,N_20192,N_19588);
xor U21030 (N_21030,N_20216,N_19572);
nor U21031 (N_21031,N_20223,N_20143);
or U21032 (N_21032,N_20400,N_20245);
or U21033 (N_21033,N_19592,N_20046);
and U21034 (N_21034,N_19844,N_20432);
or U21035 (N_21035,N_20972,N_20103);
and U21036 (N_21036,N_20189,N_19941);
xnor U21037 (N_21037,N_20244,N_20118);
and U21038 (N_21038,N_19707,N_19875);
xnor U21039 (N_21039,N_20467,N_20666);
and U21040 (N_21040,N_19972,N_20355);
nand U21041 (N_21041,N_20909,N_20827);
or U21042 (N_21042,N_19843,N_20284);
xnor U21043 (N_21043,N_20681,N_20866);
xor U21044 (N_21044,N_20899,N_20323);
or U21045 (N_21045,N_20831,N_20030);
nand U21046 (N_21046,N_20413,N_20874);
nand U21047 (N_21047,N_20828,N_19512);
and U21048 (N_21048,N_20572,N_19673);
or U21049 (N_21049,N_20329,N_20258);
or U21050 (N_21050,N_20094,N_19502);
nor U21051 (N_21051,N_20895,N_19891);
nand U21052 (N_21052,N_20368,N_19510);
or U21053 (N_21053,N_20646,N_19936);
xnor U21054 (N_21054,N_20901,N_20754);
nand U21055 (N_21055,N_20659,N_20158);
nor U21056 (N_21056,N_19612,N_20239);
or U21057 (N_21057,N_19753,N_20104);
xor U21058 (N_21058,N_20234,N_19728);
nand U21059 (N_21059,N_20133,N_19676);
nand U21060 (N_21060,N_19987,N_19543);
xor U21061 (N_21061,N_20846,N_19504);
nor U21062 (N_21062,N_20648,N_19650);
nand U21063 (N_21063,N_20339,N_20297);
nor U21064 (N_21064,N_20004,N_20907);
or U21065 (N_21065,N_20296,N_20319);
nor U21066 (N_21066,N_20680,N_20075);
xnor U21067 (N_21067,N_19744,N_20971);
xnor U21068 (N_21068,N_20002,N_19723);
nor U21069 (N_21069,N_20797,N_19810);
nand U21070 (N_21070,N_20140,N_19834);
nor U21071 (N_21071,N_20238,N_20401);
and U21072 (N_21072,N_20931,N_20364);
nand U21073 (N_21073,N_19715,N_19640);
nand U21074 (N_21074,N_20338,N_20706);
nand U21075 (N_21075,N_20864,N_20460);
xnor U21076 (N_21076,N_20042,N_20810);
nor U21077 (N_21077,N_20398,N_19568);
xnor U21078 (N_21078,N_19882,N_20122);
and U21079 (N_21079,N_20102,N_20761);
nor U21080 (N_21080,N_19711,N_20960);
and U21081 (N_21081,N_19547,N_19587);
xor U21082 (N_21082,N_20913,N_20336);
nor U21083 (N_21083,N_19595,N_20464);
nor U21084 (N_21084,N_20496,N_20048);
nand U21085 (N_21085,N_19599,N_20387);
xnor U21086 (N_21086,N_19824,N_19506);
nand U21087 (N_21087,N_20019,N_20256);
and U21088 (N_21088,N_20624,N_20278);
xnor U21089 (N_21089,N_20363,N_20945);
xnor U21090 (N_21090,N_20585,N_20530);
and U21091 (N_21091,N_19726,N_20348);
nand U21092 (N_21092,N_20028,N_20752);
or U21093 (N_21093,N_20614,N_19670);
or U21094 (N_21094,N_19688,N_20154);
and U21095 (N_21095,N_19905,N_20396);
nor U21096 (N_21096,N_20578,N_19938);
or U21097 (N_21097,N_20069,N_20818);
and U21098 (N_21098,N_19737,N_20482);
or U21099 (N_21099,N_20001,N_19950);
xor U21100 (N_21100,N_20518,N_19749);
and U21101 (N_21101,N_20986,N_20384);
nand U21102 (N_21102,N_20593,N_20469);
nand U21103 (N_21103,N_20320,N_20224);
nor U21104 (N_21104,N_19927,N_20007);
nor U21105 (N_21105,N_20902,N_19994);
xnor U21106 (N_21106,N_20667,N_19878);
nor U21107 (N_21107,N_20881,N_20687);
nor U21108 (N_21108,N_20948,N_19575);
xnor U21109 (N_21109,N_19992,N_19755);
nand U21110 (N_21110,N_19783,N_20611);
nor U21111 (N_21111,N_20036,N_20183);
or U21112 (N_21112,N_19584,N_20748);
xnor U21113 (N_21113,N_20272,N_20105);
xnor U21114 (N_21114,N_19552,N_19618);
or U21115 (N_21115,N_19765,N_20737);
nand U21116 (N_21116,N_19872,N_19995);
and U21117 (N_21117,N_20974,N_19589);
and U21118 (N_21118,N_20382,N_19869);
xnor U21119 (N_21119,N_20175,N_20704);
and U21120 (N_21120,N_20807,N_20806);
xor U21121 (N_21121,N_20759,N_19619);
nand U21122 (N_21122,N_19615,N_19675);
or U21123 (N_21123,N_19971,N_19642);
and U21124 (N_21124,N_19780,N_20527);
nor U21125 (N_21125,N_19991,N_20962);
or U21126 (N_21126,N_20543,N_19509);
or U21127 (N_21127,N_19645,N_19793);
nor U21128 (N_21128,N_19910,N_20500);
nand U21129 (N_21129,N_19916,N_19597);
and U21130 (N_21130,N_20582,N_19563);
and U21131 (N_21131,N_20961,N_20542);
and U21132 (N_21132,N_19785,N_20892);
or U21133 (N_21133,N_20740,N_20416);
and U21134 (N_21134,N_20367,N_19635);
xnor U21135 (N_21135,N_20120,N_19591);
nand U21136 (N_21136,N_20424,N_20745);
xnor U21137 (N_21137,N_19606,N_20214);
nand U21138 (N_21138,N_19805,N_19919);
nand U21139 (N_21139,N_20494,N_20672);
xor U21140 (N_21140,N_20763,N_20640);
xor U21141 (N_21141,N_19583,N_20984);
nor U21142 (N_21142,N_19686,N_20005);
or U21143 (N_21143,N_20322,N_20210);
or U21144 (N_21144,N_20997,N_20734);
xor U21145 (N_21145,N_19800,N_20703);
and U21146 (N_21146,N_19840,N_20145);
nor U21147 (N_21147,N_20114,N_19685);
and U21148 (N_21148,N_20194,N_19790);
nor U21149 (N_21149,N_19848,N_20545);
xor U21150 (N_21150,N_20539,N_20723);
xor U21151 (N_21151,N_20503,N_19914);
nand U21152 (N_21152,N_19921,N_19763);
nand U21153 (N_21153,N_20466,N_20566);
xnor U21154 (N_21154,N_20242,N_20529);
xor U21155 (N_21155,N_20887,N_20237);
xor U21156 (N_21156,N_19935,N_20581);
nand U21157 (N_21157,N_20849,N_20124);
nand U21158 (N_21158,N_20567,N_19849);
nand U21159 (N_21159,N_20458,N_20535);
xor U21160 (N_21160,N_20983,N_20616);
and U21161 (N_21161,N_20372,N_20783);
nand U21162 (N_21162,N_20231,N_20405);
nand U21163 (N_21163,N_20845,N_20819);
nand U21164 (N_21164,N_20287,N_19970);
or U21165 (N_21165,N_20410,N_19863);
xor U21166 (N_21166,N_20442,N_20801);
or U21167 (N_21167,N_20600,N_19628);
nand U21168 (N_21168,N_19974,N_20923);
nor U21169 (N_21169,N_20097,N_19786);
or U21170 (N_21170,N_20248,N_20293);
or U21171 (N_21171,N_20483,N_19508);
and U21172 (N_21172,N_20484,N_20407);
nor U21173 (N_21173,N_20436,N_20032);
nor U21174 (N_21174,N_20531,N_20383);
xor U21175 (N_21175,N_20357,N_19578);
xor U21176 (N_21176,N_19717,N_20975);
xor U21177 (N_21177,N_20497,N_19963);
nand U21178 (N_21178,N_20839,N_20084);
nand U21179 (N_21179,N_20476,N_20299);
nand U21180 (N_21180,N_19920,N_19807);
xnor U21181 (N_21181,N_19625,N_20422);
nor U21182 (N_21182,N_20385,N_20990);
and U21183 (N_21183,N_20033,N_19948);
and U21184 (N_21184,N_19955,N_19672);
nand U21185 (N_21185,N_20771,N_19764);
or U21186 (N_21186,N_20713,N_20589);
nand U21187 (N_21187,N_20817,N_20843);
or U21188 (N_21188,N_20399,N_20487);
or U21189 (N_21189,N_20583,N_20314);
and U21190 (N_21190,N_20716,N_20789);
and U21191 (N_21191,N_20804,N_20608);
xor U21192 (N_21192,N_20291,N_20760);
nor U21193 (N_21193,N_20419,N_20579);
nor U21194 (N_21194,N_20684,N_20017);
nand U21195 (N_21195,N_20190,N_19689);
or U21196 (N_21196,N_20668,N_20841);
nor U21197 (N_21197,N_19854,N_20273);
xor U21198 (N_21198,N_20811,N_19890);
and U21199 (N_21199,N_19735,N_20860);
or U21200 (N_21200,N_20222,N_19904);
xnor U21201 (N_21201,N_20625,N_19624);
and U21202 (N_21202,N_19958,N_20853);
xnor U21203 (N_21203,N_20325,N_20128);
and U21204 (N_21204,N_20262,N_20049);
nand U21205 (N_21205,N_20996,N_19602);
nand U21206 (N_21206,N_20719,N_20730);
or U21207 (N_21207,N_19906,N_19832);
or U21208 (N_21208,N_20309,N_20773);
xor U21209 (N_21209,N_19536,N_20115);
and U21210 (N_21210,N_19733,N_19725);
xnor U21211 (N_21211,N_19556,N_20279);
nor U21212 (N_21212,N_19788,N_19996);
xor U21213 (N_21213,N_20934,N_20848);
xnor U21214 (N_21214,N_20863,N_19697);
nor U21215 (N_21215,N_20623,N_20587);
xnor U21216 (N_21216,N_20604,N_20316);
nand U21217 (N_21217,N_19542,N_20209);
nor U21218 (N_21218,N_20289,N_20762);
xnor U21219 (N_21219,N_20428,N_19682);
and U21220 (N_21220,N_20930,N_20080);
and U21221 (N_21221,N_19839,N_19975);
xnor U21222 (N_21222,N_20219,N_20937);
nand U21223 (N_21223,N_20433,N_20977);
or U21224 (N_21224,N_20177,N_20510);
or U21225 (N_21225,N_20047,N_20506);
nand U21226 (N_21226,N_20559,N_20144);
nor U21227 (N_21227,N_19695,N_19865);
nor U21228 (N_21228,N_20129,N_20081);
xor U21229 (N_21229,N_20315,N_20896);
nor U21230 (N_21230,N_19656,N_20477);
and U21231 (N_21231,N_20307,N_20898);
nand U21232 (N_21232,N_19739,N_20448);
nor U21233 (N_21233,N_20010,N_20588);
and U21234 (N_21234,N_20944,N_19626);
or U21235 (N_21235,N_19850,N_20093);
nor U21236 (N_21236,N_19664,N_20963);
nand U21237 (N_21237,N_20838,N_20031);
xnor U21238 (N_21238,N_20645,N_19957);
xnor U21239 (N_21239,N_20456,N_20781);
nand U21240 (N_21240,N_20083,N_19620);
or U21241 (N_21241,N_20142,N_19570);
or U21242 (N_21242,N_19838,N_19956);
or U21243 (N_21243,N_19915,N_19911);
and U21244 (N_21244,N_19870,N_19644);
or U21245 (N_21245,N_19989,N_20270);
nand U21246 (N_21246,N_20702,N_19548);
xnor U21247 (N_21247,N_20502,N_20018);
nor U21248 (N_21248,N_19973,N_20584);
nor U21249 (N_21249,N_19774,N_20774);
and U21250 (N_21250,N_19678,N_20199);
nand U21251 (N_21251,N_19893,N_19775);
nand U21252 (N_21252,N_19883,N_20228);
and U21253 (N_21253,N_20912,N_20815);
nor U21254 (N_21254,N_20446,N_20203);
and U21255 (N_21255,N_20161,N_20855);
nand U21256 (N_21256,N_19634,N_20117);
nand U21257 (N_21257,N_20548,N_20686);
nand U21258 (N_21258,N_19703,N_20360);
xnor U21259 (N_21259,N_20966,N_20859);
xnor U21260 (N_21260,N_19933,N_19637);
and U21261 (N_21261,N_20461,N_20858);
or U21262 (N_21262,N_20550,N_19738);
or U21263 (N_21263,N_20431,N_19757);
xnor U21264 (N_21264,N_20474,N_20765);
xnor U21265 (N_21265,N_20897,N_20301);
xnor U21266 (N_21266,N_20823,N_20649);
or U21267 (N_21267,N_20099,N_20178);
xor U21268 (N_21268,N_19687,N_19953);
or U21269 (N_21269,N_20330,N_20925);
xor U21270 (N_21270,N_20731,N_20091);
nor U21271 (N_21271,N_20250,N_19555);
or U21272 (N_21272,N_20919,N_20756);
and U21273 (N_21273,N_20027,N_19818);
nand U21274 (N_21274,N_20568,N_19968);
nand U21275 (N_21275,N_19982,N_19621);
nor U21276 (N_21276,N_20562,N_20772);
and U21277 (N_21277,N_19517,N_20900);
nor U21278 (N_21278,N_20024,N_19837);
and U21279 (N_21279,N_20890,N_20854);
nor U21280 (N_21280,N_20626,N_20109);
and U21281 (N_21281,N_20799,N_20800);
nor U21282 (N_21282,N_19665,N_20110);
nand U21283 (N_21283,N_20193,N_19831);
or U21284 (N_21284,N_20021,N_20269);
or U21285 (N_21285,N_19633,N_20969);
nor U21286 (N_21286,N_20286,N_20313);
nor U21287 (N_21287,N_19902,N_20844);
and U21288 (N_21288,N_20886,N_20308);
xnor U21289 (N_21289,N_20630,N_19627);
and U21290 (N_21290,N_20359,N_19551);
or U21291 (N_21291,N_20764,N_20463);
or U21292 (N_21292,N_20173,N_20455);
or U21293 (N_21293,N_20417,N_19845);
and U21294 (N_21294,N_20073,N_19758);
nor U21295 (N_21295,N_20029,N_19629);
nor U21296 (N_21296,N_20054,N_20546);
nor U21297 (N_21297,N_20664,N_19661);
or U21298 (N_21298,N_19666,N_20180);
nand U21299 (N_21299,N_19704,N_20016);
and U21300 (N_21300,N_19718,N_19586);
xor U21301 (N_21301,N_20657,N_20515);
nand U21302 (N_21302,N_19525,N_20200);
nand U21303 (N_21303,N_20067,N_20514);
nand U21304 (N_21304,N_20970,N_20921);
nor U21305 (N_21305,N_20427,N_19828);
nor U21306 (N_21306,N_20776,N_19590);
nor U21307 (N_21307,N_20560,N_20915);
or U21308 (N_21308,N_19750,N_20932);
nand U21309 (N_21309,N_19754,N_19929);
or U21310 (N_21310,N_19544,N_20471);
nor U21311 (N_21311,N_20092,N_20634);
nand U21312 (N_21312,N_20820,N_19527);
nor U21313 (N_21313,N_20775,N_20796);
nor U21314 (N_21314,N_20498,N_20628);
nor U21315 (N_21315,N_20968,N_20825);
xor U21316 (N_21316,N_19814,N_20592);
or U21317 (N_21317,N_19846,N_20670);
nand U21318 (N_21318,N_20480,N_20064);
nor U21319 (N_21319,N_20617,N_19823);
xnor U21320 (N_21320,N_20620,N_20876);
nor U21321 (N_21321,N_20333,N_19748);
or U21322 (N_21322,N_20728,N_20188);
nor U21323 (N_21323,N_20705,N_20285);
nand U21324 (N_21324,N_19534,N_19794);
nand U21325 (N_21325,N_19752,N_19960);
nand U21326 (N_21326,N_19978,N_20744);
and U21327 (N_21327,N_20955,N_19535);
and U21328 (N_21328,N_20711,N_20867);
nand U21329 (N_21329,N_20981,N_19817);
or U21330 (N_21330,N_20644,N_20337);
or U21331 (N_21331,N_20119,N_20198);
nand U21332 (N_21332,N_19520,N_19641);
xor U21333 (N_21333,N_20650,N_20386);
and U21334 (N_21334,N_19990,N_19879);
xnor U21335 (N_21335,N_19734,N_19600);
or U21336 (N_21336,N_20596,N_20488);
nand U21337 (N_21337,N_20652,N_20089);
or U21338 (N_21338,N_19897,N_20167);
and U21339 (N_21339,N_19917,N_20207);
or U21340 (N_21340,N_19965,N_20479);
nand U21341 (N_21341,N_19771,N_20980);
and U21342 (N_21342,N_20682,N_20470);
and U21343 (N_21343,N_19855,N_20647);
and U21344 (N_21344,N_20549,N_19856);
and U21345 (N_21345,N_19643,N_20295);
nand U21346 (N_21346,N_20465,N_20112);
and U21347 (N_21347,N_19576,N_20688);
or U21348 (N_21348,N_20720,N_20077);
xnor U21349 (N_21349,N_20824,N_19847);
xnor U21350 (N_21350,N_19709,N_19773);
nand U21351 (N_21351,N_20786,N_20777);
and U21352 (N_21352,N_20651,N_20735);
and U21353 (N_21353,N_20127,N_20495);
and U21354 (N_21354,N_20717,N_20061);
or U21355 (N_21355,N_20429,N_19770);
and U21356 (N_21356,N_20513,N_19822);
nand U21357 (N_21357,N_19529,N_19611);
and U21358 (N_21358,N_19694,N_19660);
nand U21359 (N_21359,N_19769,N_19873);
nand U21360 (N_21360,N_20710,N_19696);
or U21361 (N_21361,N_20918,N_20159);
nand U21362 (N_21362,N_20440,N_20791);
xnor U21363 (N_21363,N_20926,N_20743);
and U21364 (N_21364,N_20533,N_19913);
and U21365 (N_21365,N_19900,N_20613);
or U21366 (N_21366,N_20840,N_20976);
nand U21367 (N_21367,N_20232,N_20342);
nand U21368 (N_21368,N_20792,N_19884);
nor U21369 (N_21369,N_20052,N_20908);
nand U21370 (N_21370,N_19825,N_20402);
and U21371 (N_21371,N_19928,N_20871);
nand U21372 (N_21372,N_20212,N_19518);
nor U21373 (N_21373,N_19659,N_20537);
xor U21374 (N_21374,N_20565,N_19530);
nor U21375 (N_21375,N_20903,N_19614);
nand U21376 (N_21376,N_19761,N_20950);
nand U21377 (N_21377,N_20332,N_20692);
or U21378 (N_21378,N_19819,N_20747);
nand U21379 (N_21379,N_20344,N_19545);
and U21380 (N_21380,N_20837,N_20766);
nand U21381 (N_21381,N_20618,N_20501);
and U21382 (N_21382,N_19699,N_20938);
and U21383 (N_21383,N_20437,N_19713);
xnor U21384 (N_21384,N_19522,N_19967);
or U21385 (N_21385,N_19966,N_20987);
nor U21386 (N_21386,N_20988,N_20246);
nand U21387 (N_21387,N_20310,N_19712);
xor U21388 (N_21388,N_19903,N_20978);
and U21389 (N_21389,N_20430,N_20758);
xnor U21390 (N_21390,N_20187,N_20904);
xnor U21391 (N_21391,N_20780,N_20675);
and U21392 (N_21392,N_20186,N_20563);
xor U21393 (N_21393,N_20882,N_20327);
xnor U21394 (N_21394,N_20564,N_19820);
and U21395 (N_21395,N_20201,N_20633);
nand U21396 (N_21396,N_20555,N_20421);
nor U21397 (N_21397,N_19719,N_20056);
nor U21398 (N_21398,N_20107,N_20964);
nand U21399 (N_21399,N_20263,N_20249);
and U21400 (N_21400,N_20126,N_19647);
nand U21401 (N_21401,N_19605,N_20283);
nor U21402 (N_21402,N_20078,N_20090);
xor U21403 (N_21403,N_19782,N_19806);
and U21404 (N_21404,N_19851,N_20300);
nor U21405 (N_21405,N_19684,N_20473);
nand U21406 (N_21406,N_19922,N_19671);
and U21407 (N_21407,N_19768,N_20595);
xor U21408 (N_21408,N_20035,N_20395);
and U21409 (N_21409,N_20733,N_19874);
xnor U21410 (N_21410,N_20008,N_20132);
nor U21411 (N_21411,N_20660,N_20101);
nor U21412 (N_21412,N_20812,N_20022);
nor U21413 (N_21413,N_20519,N_20445);
and U21414 (N_21414,N_20532,N_20577);
nand U21415 (N_21415,N_20544,N_19571);
or U21416 (N_21416,N_20347,N_20009);
xor U21417 (N_21417,N_20516,N_20725);
or U21418 (N_21418,N_20162,N_20302);
or U21419 (N_21419,N_19925,N_20696);
nor U21420 (N_21420,N_20489,N_19797);
or U21421 (N_21421,N_20674,N_19803);
nor U21422 (N_21422,N_20629,N_19776);
nor U21423 (N_21423,N_20375,N_20251);
nand U21424 (N_21424,N_19674,N_20700);
nor U21425 (N_21425,N_20942,N_19610);
and U21426 (N_21426,N_20610,N_20197);
or U21427 (N_21427,N_20169,N_19836);
nand U21428 (N_21428,N_19663,N_20079);
xnor U21429 (N_21429,N_20534,N_20742);
nor U21430 (N_21430,N_20454,N_19947);
or U21431 (N_21431,N_19521,N_20936);
nand U21432 (N_21432,N_20965,N_20779);
or U21433 (N_21433,N_20785,N_19864);
xnor U21434 (N_21434,N_20040,N_19745);
and U21435 (N_21435,N_20362,N_20746);
nor U21436 (N_21436,N_20906,N_20371);
xnor U21437 (N_21437,N_19896,N_19731);
nor U21438 (N_21438,N_19809,N_20693);
or U21439 (N_21439,N_20096,N_20643);
nand U21440 (N_21440,N_20195,N_20225);
and U21441 (N_21441,N_20220,N_20953);
nand U21442 (N_21442,N_19899,N_19505);
nor U21443 (N_21443,N_20155,N_20176);
xor U21444 (N_21444,N_19976,N_20505);
or U21445 (N_21445,N_20958,N_20995);
or U21446 (N_21446,N_19924,N_19772);
nand U21447 (N_21447,N_20590,N_20478);
or U21448 (N_21448,N_19951,N_20768);
nand U21449 (N_21449,N_19876,N_20755);
nor U21450 (N_21450,N_20875,N_20973);
or U21451 (N_21451,N_19513,N_19894);
or U21452 (N_21452,N_19562,N_20050);
and U21453 (N_21453,N_20541,N_20449);
nor U21454 (N_21454,N_20388,N_20916);
or U21455 (N_21455,N_20808,N_20757);
and U21456 (N_21456,N_20317,N_19558);
nor U21457 (N_21457,N_20994,N_19714);
nand U21458 (N_21458,N_20485,N_20181);
xnor U21459 (N_21459,N_20750,N_19741);
nand U21460 (N_21460,N_20929,N_19705);
nor U21461 (N_21461,N_19743,N_20164);
xnor U21462 (N_21462,N_19742,N_20136);
nor U21463 (N_21463,N_19557,N_19657);
nor U21464 (N_21464,N_20282,N_20053);
or U21465 (N_21465,N_20861,N_20922);
nor U21466 (N_21466,N_20946,N_20037);
nand U21467 (N_21467,N_20732,N_19826);
xnor U21468 (N_21468,N_20941,N_19531);
nand U21469 (N_21469,N_19706,N_19777);
or U21470 (N_21470,N_20163,N_20202);
nand U21471 (N_21471,N_20782,N_20993);
and U21472 (N_21472,N_20956,N_20259);
or U21473 (N_21473,N_19932,N_20134);
nor U21474 (N_21474,N_20857,N_20444);
nor U21475 (N_21475,N_20951,N_19553);
and U21476 (N_21476,N_20689,N_20125);
and U21477 (N_21477,N_19593,N_19887);
nor U21478 (N_21478,N_20443,N_20168);
nor U21479 (N_21479,N_20023,N_20227);
nor U21480 (N_21480,N_20369,N_19944);
nor U21481 (N_21481,N_20914,N_20343);
xnor U21482 (N_21482,N_20522,N_20185);
nor U21483 (N_21483,N_19601,N_19931);
nor U21484 (N_21484,N_20475,N_19604);
or U21485 (N_21485,N_20457,N_19582);
or U21486 (N_21486,N_19984,N_19766);
or U21487 (N_21487,N_20294,N_20298);
xnor U21488 (N_21488,N_19937,N_20524);
xnor U21489 (N_21489,N_20253,N_19909);
nand U21490 (N_21490,N_20020,N_20156);
xnor U21491 (N_21491,N_20709,N_20636);
or U21492 (N_21492,N_20607,N_20172);
xnor U21493 (N_21493,N_20472,N_20041);
nand U21494 (N_21494,N_20137,N_20170);
xor U21495 (N_21495,N_20379,N_20521);
nand U21496 (N_21496,N_20509,N_20598);
and U21497 (N_21497,N_19617,N_20575);
and U21498 (N_21498,N_20609,N_19613);
nor U21499 (N_21499,N_20252,N_19821);
xor U21500 (N_21500,N_19511,N_20328);
and U21501 (N_21501,N_20570,N_20952);
xnor U21502 (N_21502,N_20835,N_19784);
xor U21503 (N_21503,N_19609,N_19669);
or U21504 (N_21504,N_20034,N_19730);
and U21505 (N_21505,N_20795,N_19564);
xnor U21506 (N_21506,N_20793,N_19532);
nor U21507 (N_21507,N_20213,N_20160);
or U21508 (N_21508,N_19943,N_20597);
or U21509 (N_21509,N_20468,N_20574);
xor U21510 (N_21510,N_20205,N_20635);
nand U21511 (N_21511,N_20254,N_19708);
xnor U21512 (N_21512,N_20580,N_19740);
nor U21513 (N_21513,N_20715,N_20490);
xnor U21514 (N_21514,N_19962,N_20641);
xnor U21515 (N_21515,N_19981,N_20441);
xor U21516 (N_21516,N_20147,N_20979);
and U21517 (N_21517,N_20277,N_19853);
xor U21518 (N_21518,N_20694,N_19528);
xor U21519 (N_21519,N_19801,N_20243);
or U21520 (N_21520,N_20698,N_19813);
xnor U21521 (N_21521,N_20809,N_20275);
nand U21522 (N_21522,N_20108,N_20235);
and U21523 (N_21523,N_20569,N_20374);
xnor U21524 (N_21524,N_19787,N_20615);
and U21525 (N_21525,N_19683,N_19539);
nand U21526 (N_21526,N_19679,N_19833);
nand U21527 (N_21527,N_20152,N_20257);
nand U21528 (N_21528,N_20940,N_20957);
xnor U21529 (N_21529,N_20058,N_19632);
nand U21530 (N_21530,N_19861,N_20072);
xor U21531 (N_21531,N_19540,N_20517);
xor U21532 (N_21532,N_19779,N_20662);
and U21533 (N_21533,N_20039,N_20599);
nor U21534 (N_21534,N_20240,N_20992);
xnor U21535 (N_21535,N_20591,N_20447);
or U21536 (N_21536,N_20894,N_20554);
or U21537 (N_21537,N_20459,N_20998);
and U21538 (N_21538,N_20605,N_20586);
or U21539 (N_21539,N_19732,N_20699);
nor U21540 (N_21540,N_19680,N_19811);
nor U21541 (N_21541,N_19596,N_20803);
nand U21542 (N_21542,N_19580,N_20230);
or U21543 (N_21543,N_20917,N_19789);
nor U21544 (N_21544,N_19959,N_20012);
xnor U21545 (N_21545,N_19523,N_20218);
or U21546 (N_21546,N_20340,N_20695);
and U21547 (N_21547,N_20943,N_20179);
xnor U21548 (N_21548,N_20380,N_19607);
nand U21549 (N_21549,N_20165,N_20408);
and U21550 (N_21550,N_20106,N_19778);
nor U21551 (N_21551,N_20868,N_20933);
nor U21552 (N_21552,N_20528,N_19898);
or U21553 (N_21553,N_20438,N_20280);
and U21554 (N_21554,N_20905,N_20352);
xnor U21555 (N_21555,N_20814,N_20678);
and U21556 (N_21556,N_19934,N_19651);
or U21557 (N_21557,N_20788,N_19561);
and U21558 (N_21558,N_20697,N_19662);
xor U21559 (N_21559,N_20085,N_20935);
xnor U21560 (N_21560,N_20116,N_19524);
nand U21561 (N_21561,N_20724,N_19942);
nand U21562 (N_21562,N_20051,N_19829);
nand U21563 (N_21563,N_20870,N_19871);
nor U21564 (N_21564,N_20661,N_20059);
or U21565 (N_21565,N_19945,N_19926);
nand U21566 (N_21566,N_20850,N_20753);
or U21567 (N_21567,N_20525,N_19636);
xor U21568 (N_21568,N_20335,N_19866);
nor U21569 (N_21569,N_19997,N_20351);
nand U21570 (N_21570,N_19888,N_20274);
or U21571 (N_21571,N_20880,N_19507);
xnor U21572 (N_21572,N_20434,N_19554);
xor U21573 (N_21573,N_20070,N_19598);
or U21574 (N_21574,N_20226,N_20426);
nor U21575 (N_21575,N_19546,N_20642);
or U21576 (N_21576,N_19881,N_20453);
or U21577 (N_21577,N_20211,N_20989);
nand U21578 (N_21578,N_20206,N_19720);
xnor U21579 (N_21579,N_19623,N_20389);
nor U21580 (N_21580,N_20055,N_20011);
and U21581 (N_21581,N_20833,N_19892);
xnor U21582 (N_21582,N_19969,N_19608);
nor U21583 (N_21583,N_20677,N_20376);
nor U21584 (N_21584,N_19907,N_20146);
or U21585 (N_21585,N_19692,N_20450);
nand U21586 (N_21586,N_20712,N_20370);
nor U21587 (N_21587,N_20520,N_20679);
nand U21588 (N_21588,N_20767,N_20166);
or U21589 (N_21589,N_20304,N_20358);
or U21590 (N_21590,N_20727,N_19646);
xnor U21591 (N_21591,N_20393,N_20014);
and U21592 (N_21592,N_20229,N_20749);
or U21593 (N_21593,N_20999,N_20174);
nor U21594 (N_21594,N_19762,N_20303);
nand U21595 (N_21595,N_20276,N_20547);
nand U21596 (N_21596,N_19923,N_20622);
nor U21597 (N_21597,N_20721,N_19721);
xnor U21598 (N_21598,N_20722,N_20098);
or U21599 (N_21599,N_19815,N_20507);
and U21600 (N_21600,N_19759,N_20281);
nand U21601 (N_21601,N_20638,N_19880);
and U21602 (N_21602,N_20991,N_20508);
and U21603 (N_21603,N_20411,N_20182);
nand U21604 (N_21604,N_20561,N_19912);
xor U21605 (N_21605,N_20415,N_20842);
nand U21606 (N_21606,N_20601,N_20452);
xor U21607 (N_21607,N_20373,N_20026);
nor U21608 (N_21608,N_20639,N_20910);
xnor U21609 (N_21609,N_20045,N_19799);
or U21610 (N_21610,N_20071,N_19722);
nor U21611 (N_21611,N_19514,N_20062);
or U21612 (N_21612,N_20391,N_19541);
nor U21613 (N_21613,N_19729,N_20121);
and U21614 (N_21614,N_19549,N_19841);
or U21615 (N_21615,N_19980,N_19716);
xnor U21616 (N_21616,N_19862,N_20312);
xor U21617 (N_21617,N_20361,N_20271);
or U21618 (N_21618,N_19827,N_19886);
or U21619 (N_21619,N_20082,N_19964);
nand U21620 (N_21620,N_20893,N_19867);
and U21621 (N_21621,N_20538,N_19649);
and U21622 (N_21622,N_20261,N_20111);
xnor U21623 (N_21623,N_20057,N_20068);
xnor U21624 (N_21624,N_19638,N_20879);
and U21625 (N_21625,N_20409,N_20654);
xor U21626 (N_21626,N_19977,N_20954);
nand U21627 (N_21627,N_19804,N_19700);
nor U21628 (N_21628,N_20265,N_20366);
nand U21629 (N_21629,N_20013,N_19901);
and U21630 (N_21630,N_19653,N_20131);
or U21631 (N_21631,N_19569,N_19581);
xnor U21632 (N_21632,N_20236,N_20135);
nand U21633 (N_21633,N_20439,N_20690);
xor U21634 (N_21634,N_20208,N_19908);
nor U21635 (N_21635,N_19698,N_20191);
nor U21636 (N_21636,N_20006,N_20873);
nand U21637 (N_21637,N_20852,N_19767);
or U21638 (N_21638,N_20404,N_19727);
nand U21639 (N_21639,N_19574,N_20123);
xor U21640 (N_21640,N_19603,N_20655);
nand U21641 (N_21641,N_19677,N_20865);
xnor U21642 (N_21642,N_20676,N_19567);
nand U21643 (N_21643,N_20247,N_20341);
and U21644 (N_21644,N_20888,N_19859);
xor U21645 (N_21645,N_20891,N_19630);
and U21646 (N_21646,N_20292,N_20834);
and U21647 (N_21647,N_20982,N_20403);
xnor U21648 (N_21648,N_20043,N_20486);
or U21649 (N_21649,N_20153,N_20927);
or U21650 (N_21650,N_20805,N_19746);
xor U21651 (N_21651,N_20215,N_20377);
nand U21652 (N_21652,N_20798,N_20816);
xnor U21653 (N_21653,N_20573,N_20924);
nor U21654 (N_21654,N_20321,N_20354);
xnor U21655 (N_21655,N_19756,N_19577);
and U21656 (N_21656,N_19503,N_19526);
xor U21657 (N_21657,N_19979,N_20665);
xnor U21658 (N_21658,N_20558,N_19812);
and U21659 (N_21659,N_20241,N_20392);
xnor U21660 (N_21660,N_20632,N_20268);
xor U21661 (N_21661,N_20671,N_20653);
nor U21662 (N_21662,N_20390,N_19690);
and U21663 (N_21663,N_19796,N_20451);
and U21664 (N_21664,N_20884,N_19985);
and U21665 (N_21665,N_19895,N_20149);
nor U21666 (N_21666,N_20612,N_20378);
nor U21667 (N_21667,N_20290,N_19736);
nand U21668 (N_21668,N_20196,N_20306);
xnor U21669 (N_21669,N_19791,N_19877);
and U21670 (N_21670,N_20729,N_19501);
nand U21671 (N_21671,N_19594,N_20397);
or U21672 (N_21672,N_20086,N_19830);
xnor U21673 (N_21673,N_19747,N_20060);
nand U21674 (N_21674,N_19566,N_20691);
nor U21675 (N_21675,N_20856,N_20412);
or U21676 (N_21676,N_19999,N_19538);
xnor U21677 (N_21677,N_20435,N_19792);
xnor U21678 (N_21678,N_20171,N_19954);
nor U21679 (N_21679,N_19681,N_20260);
or U21680 (N_21680,N_20714,N_20552);
xnor U21681 (N_21681,N_19639,N_20802);
xor U21682 (N_21682,N_20778,N_20499);
xor U21683 (N_21683,N_20920,N_20365);
or U21684 (N_21684,N_20959,N_20726);
nor U21685 (N_21685,N_19533,N_19724);
or U21686 (N_21686,N_20414,N_20594);
nor U21687 (N_21687,N_20829,N_20967);
nand U21688 (N_21688,N_20462,N_20621);
nand U21689 (N_21689,N_19655,N_20324);
and U21690 (N_21690,N_19795,N_20088);
and U21691 (N_21691,N_20504,N_19579);
xor U21692 (N_21692,N_19550,N_20751);
nand U21693 (N_21693,N_20741,N_20836);
xor U21694 (N_21694,N_19816,N_19781);
nor U21695 (N_21695,N_19537,N_20536);
and U21696 (N_21696,N_19560,N_19857);
nor U21697 (N_21697,N_19860,N_19961);
and U21698 (N_21698,N_19658,N_19515);
xnor U21699 (N_21699,N_20000,N_20076);
nor U21700 (N_21700,N_19998,N_19868);
and U21701 (N_21701,N_20663,N_19802);
and U21702 (N_21702,N_20826,N_20264);
and U21703 (N_21703,N_20334,N_20512);
or U21704 (N_21704,N_20571,N_20738);
or U21705 (N_21705,N_19693,N_20087);
nor U21706 (N_21706,N_20883,N_20631);
nor U21707 (N_21707,N_19631,N_20025);
and U21708 (N_21708,N_19808,N_20708);
and U21709 (N_21709,N_20637,N_20619);
nand U21710 (N_21710,N_20095,N_20356);
nor U21711 (N_21711,N_20821,N_19648);
and U21712 (N_21712,N_20318,N_20553);
or U21713 (N_21713,N_20151,N_20233);
xnor U21714 (N_21714,N_20669,N_20492);
xor U21715 (N_21715,N_19983,N_20928);
or U21716 (N_21716,N_20311,N_20830);
nand U21717 (N_21717,N_19667,N_20878);
nand U21718 (N_21718,N_20576,N_20038);
nor U21719 (N_21719,N_19710,N_19940);
and U21720 (N_21720,N_20015,N_20701);
or U21721 (N_21721,N_20148,N_20406);
nor U21722 (N_21722,N_20420,N_19519);
nand U21723 (N_21723,N_20204,N_20847);
or U21724 (N_21724,N_19654,N_20736);
xnor U21725 (N_21725,N_20889,N_20381);
nand U21726 (N_21726,N_20794,N_19559);
or U21727 (N_21727,N_20869,N_20526);
or U21728 (N_21728,N_20100,N_20305);
or U21729 (N_21729,N_20349,N_20872);
or U21730 (N_21730,N_19573,N_20557);
and U21731 (N_21731,N_20157,N_20784);
or U21732 (N_21732,N_19760,N_20787);
nor U21733 (N_21733,N_20739,N_20130);
nor U21734 (N_21734,N_20683,N_20540);
and U21735 (N_21735,N_20418,N_19993);
xnor U21736 (N_21736,N_19565,N_20656);
xnor U21737 (N_21737,N_20885,N_20658);
nor U21738 (N_21738,N_20423,N_20949);
or U21739 (N_21739,N_20603,N_19585);
or U21740 (N_21740,N_20003,N_19701);
xor U21741 (N_21741,N_20627,N_20551);
xor U21742 (N_21742,N_20141,N_19930);
or U21743 (N_21743,N_19858,N_19939);
and U21744 (N_21744,N_19835,N_20255);
nand U21745 (N_21745,N_20606,N_20288);
nor U21746 (N_21746,N_20267,N_20877);
and U21747 (N_21747,N_20063,N_19949);
nand U21748 (N_21748,N_19668,N_19622);
and U21749 (N_21749,N_20066,N_19889);
or U21750 (N_21750,N_20065,N_20861);
xor U21751 (N_21751,N_20067,N_20147);
nor U21752 (N_21752,N_20987,N_19507);
nor U21753 (N_21753,N_20670,N_20089);
nand U21754 (N_21754,N_19807,N_19928);
xnor U21755 (N_21755,N_20039,N_20988);
xnor U21756 (N_21756,N_20283,N_20968);
and U21757 (N_21757,N_19630,N_20415);
and U21758 (N_21758,N_19830,N_19823);
or U21759 (N_21759,N_20791,N_20455);
and U21760 (N_21760,N_20718,N_20097);
or U21761 (N_21761,N_20855,N_20276);
and U21762 (N_21762,N_20021,N_19826);
nor U21763 (N_21763,N_19796,N_20963);
nor U21764 (N_21764,N_19957,N_20229);
and U21765 (N_21765,N_20322,N_20054);
and U21766 (N_21766,N_20993,N_20921);
nand U21767 (N_21767,N_20574,N_20549);
nor U21768 (N_21768,N_20378,N_19711);
xor U21769 (N_21769,N_20326,N_20434);
nand U21770 (N_21770,N_19922,N_19727);
xor U21771 (N_21771,N_20498,N_20822);
and U21772 (N_21772,N_19561,N_20423);
and U21773 (N_21773,N_20868,N_20358);
xor U21774 (N_21774,N_20385,N_20135);
xnor U21775 (N_21775,N_20948,N_20870);
xor U21776 (N_21776,N_20671,N_20074);
or U21777 (N_21777,N_19575,N_20882);
nor U21778 (N_21778,N_19647,N_19680);
xor U21779 (N_21779,N_20897,N_19545);
nor U21780 (N_21780,N_20925,N_20546);
xnor U21781 (N_21781,N_19770,N_20373);
and U21782 (N_21782,N_19824,N_20907);
xor U21783 (N_21783,N_20054,N_20654);
nor U21784 (N_21784,N_20735,N_20774);
nand U21785 (N_21785,N_19586,N_20094);
or U21786 (N_21786,N_20093,N_19537);
or U21787 (N_21787,N_20634,N_19775);
nor U21788 (N_21788,N_20859,N_20662);
nand U21789 (N_21789,N_20302,N_20983);
nor U21790 (N_21790,N_19731,N_19658);
and U21791 (N_21791,N_20512,N_19599);
or U21792 (N_21792,N_20343,N_20504);
or U21793 (N_21793,N_20566,N_19661);
and U21794 (N_21794,N_20365,N_20760);
or U21795 (N_21795,N_19615,N_20507);
nor U21796 (N_21796,N_20792,N_19546);
xor U21797 (N_21797,N_20181,N_20762);
xor U21798 (N_21798,N_19751,N_20677);
or U21799 (N_21799,N_20938,N_20643);
xor U21800 (N_21800,N_19516,N_19810);
or U21801 (N_21801,N_19624,N_20501);
and U21802 (N_21802,N_20430,N_19836);
nor U21803 (N_21803,N_20651,N_19565);
or U21804 (N_21804,N_19749,N_19852);
and U21805 (N_21805,N_19604,N_19950);
and U21806 (N_21806,N_20692,N_19780);
nand U21807 (N_21807,N_20545,N_20205);
nand U21808 (N_21808,N_19662,N_20277);
or U21809 (N_21809,N_20216,N_20806);
and U21810 (N_21810,N_19942,N_20662);
and U21811 (N_21811,N_20064,N_19800);
nand U21812 (N_21812,N_20087,N_20608);
and U21813 (N_21813,N_20456,N_19939);
or U21814 (N_21814,N_19563,N_20202);
and U21815 (N_21815,N_20447,N_20621);
and U21816 (N_21816,N_19529,N_20130);
nor U21817 (N_21817,N_20036,N_19805);
nand U21818 (N_21818,N_20529,N_20424);
nand U21819 (N_21819,N_19598,N_20892);
and U21820 (N_21820,N_20837,N_20426);
nand U21821 (N_21821,N_20557,N_20202);
or U21822 (N_21822,N_20945,N_20751);
and U21823 (N_21823,N_20358,N_20459);
or U21824 (N_21824,N_19810,N_19513);
nor U21825 (N_21825,N_20803,N_20808);
or U21826 (N_21826,N_19533,N_20691);
nor U21827 (N_21827,N_20169,N_20680);
xnor U21828 (N_21828,N_19711,N_20739);
xor U21829 (N_21829,N_19839,N_19748);
xnor U21830 (N_21830,N_19996,N_19566);
nand U21831 (N_21831,N_20892,N_19798);
xnor U21832 (N_21832,N_20645,N_20843);
or U21833 (N_21833,N_20951,N_20556);
nand U21834 (N_21834,N_19905,N_20150);
xnor U21835 (N_21835,N_20340,N_20762);
and U21836 (N_21836,N_20971,N_19584);
and U21837 (N_21837,N_20085,N_20618);
nor U21838 (N_21838,N_20737,N_19657);
and U21839 (N_21839,N_20416,N_20684);
nand U21840 (N_21840,N_20003,N_19572);
nor U21841 (N_21841,N_20383,N_20863);
and U21842 (N_21842,N_20879,N_20885);
or U21843 (N_21843,N_19995,N_20513);
or U21844 (N_21844,N_20644,N_19906);
or U21845 (N_21845,N_20692,N_20434);
nand U21846 (N_21846,N_20953,N_19593);
nand U21847 (N_21847,N_19701,N_20503);
xnor U21848 (N_21848,N_20124,N_19580);
nand U21849 (N_21849,N_19635,N_19902);
nor U21850 (N_21850,N_20957,N_20058);
nor U21851 (N_21851,N_20666,N_20717);
nand U21852 (N_21852,N_19810,N_20197);
nor U21853 (N_21853,N_20315,N_19908);
nand U21854 (N_21854,N_20667,N_19580);
or U21855 (N_21855,N_19968,N_20421);
nor U21856 (N_21856,N_19983,N_20261);
or U21857 (N_21857,N_19869,N_19662);
xnor U21858 (N_21858,N_20231,N_20363);
nor U21859 (N_21859,N_20313,N_19552);
xnor U21860 (N_21860,N_20585,N_19970);
and U21861 (N_21861,N_20261,N_20405);
or U21862 (N_21862,N_20070,N_20717);
xor U21863 (N_21863,N_20442,N_20800);
or U21864 (N_21864,N_20415,N_20734);
nor U21865 (N_21865,N_20765,N_20714);
nand U21866 (N_21866,N_19532,N_20939);
or U21867 (N_21867,N_20318,N_19678);
and U21868 (N_21868,N_20514,N_19926);
nand U21869 (N_21869,N_19765,N_19697);
or U21870 (N_21870,N_19967,N_20518);
or U21871 (N_21871,N_20223,N_20403);
and U21872 (N_21872,N_20031,N_20072);
nand U21873 (N_21873,N_20593,N_20963);
or U21874 (N_21874,N_19581,N_20871);
nand U21875 (N_21875,N_20831,N_20065);
or U21876 (N_21876,N_20533,N_20576);
nor U21877 (N_21877,N_19912,N_20559);
and U21878 (N_21878,N_20414,N_20279);
xnor U21879 (N_21879,N_20522,N_20934);
xor U21880 (N_21880,N_19576,N_20329);
xor U21881 (N_21881,N_19544,N_20699);
or U21882 (N_21882,N_19661,N_20528);
nor U21883 (N_21883,N_20506,N_20834);
nand U21884 (N_21884,N_20971,N_20960);
nand U21885 (N_21885,N_20734,N_20637);
or U21886 (N_21886,N_20747,N_20786);
nor U21887 (N_21887,N_20598,N_20134);
and U21888 (N_21888,N_20758,N_19928);
nor U21889 (N_21889,N_20277,N_19882);
or U21890 (N_21890,N_20661,N_19561);
and U21891 (N_21891,N_19635,N_20606);
nand U21892 (N_21892,N_19806,N_19631);
xnor U21893 (N_21893,N_19736,N_20651);
xor U21894 (N_21894,N_20378,N_20281);
xor U21895 (N_21895,N_20937,N_20387);
nand U21896 (N_21896,N_19893,N_19648);
xor U21897 (N_21897,N_20063,N_19865);
nor U21898 (N_21898,N_19874,N_20509);
and U21899 (N_21899,N_20644,N_20102);
nor U21900 (N_21900,N_20286,N_19683);
nor U21901 (N_21901,N_20623,N_20255);
or U21902 (N_21902,N_19598,N_20224);
or U21903 (N_21903,N_20039,N_19507);
or U21904 (N_21904,N_20987,N_19935);
nand U21905 (N_21905,N_19826,N_20812);
nor U21906 (N_21906,N_19506,N_20569);
nor U21907 (N_21907,N_20507,N_20495);
nor U21908 (N_21908,N_19500,N_19772);
or U21909 (N_21909,N_20810,N_20635);
nor U21910 (N_21910,N_19796,N_20184);
nor U21911 (N_21911,N_20728,N_19595);
nand U21912 (N_21912,N_19702,N_20766);
nand U21913 (N_21913,N_19613,N_20965);
or U21914 (N_21914,N_19984,N_19540);
and U21915 (N_21915,N_19870,N_20333);
xor U21916 (N_21916,N_20730,N_19529);
xor U21917 (N_21917,N_20248,N_20219);
nor U21918 (N_21918,N_20118,N_20766);
and U21919 (N_21919,N_20737,N_20693);
or U21920 (N_21920,N_20099,N_19691);
xnor U21921 (N_21921,N_19970,N_19973);
nor U21922 (N_21922,N_20739,N_20052);
and U21923 (N_21923,N_19645,N_20770);
xor U21924 (N_21924,N_20583,N_20001);
xnor U21925 (N_21925,N_20823,N_20523);
nand U21926 (N_21926,N_20087,N_20118);
xnor U21927 (N_21927,N_20149,N_20507);
nor U21928 (N_21928,N_20234,N_20143);
nor U21929 (N_21929,N_20300,N_20336);
xor U21930 (N_21930,N_20998,N_20771);
nand U21931 (N_21931,N_20004,N_20391);
or U21932 (N_21932,N_20865,N_19620);
nand U21933 (N_21933,N_20072,N_20850);
and U21934 (N_21934,N_19514,N_20139);
nor U21935 (N_21935,N_20422,N_20205);
or U21936 (N_21936,N_20181,N_20603);
and U21937 (N_21937,N_19514,N_19969);
nand U21938 (N_21938,N_20720,N_20068);
xnor U21939 (N_21939,N_20384,N_19832);
nor U21940 (N_21940,N_20459,N_19584);
nand U21941 (N_21941,N_19630,N_20429);
xor U21942 (N_21942,N_20538,N_20636);
nor U21943 (N_21943,N_20964,N_20266);
nor U21944 (N_21944,N_19909,N_20767);
xor U21945 (N_21945,N_19534,N_19821);
nand U21946 (N_21946,N_19731,N_20442);
or U21947 (N_21947,N_19751,N_20023);
and U21948 (N_21948,N_20117,N_20963);
nand U21949 (N_21949,N_19644,N_20232);
nor U21950 (N_21950,N_20164,N_20979);
xnor U21951 (N_21951,N_19957,N_20615);
or U21952 (N_21952,N_19571,N_20060);
or U21953 (N_21953,N_19548,N_20852);
xnor U21954 (N_21954,N_19607,N_20822);
nand U21955 (N_21955,N_19634,N_20106);
and U21956 (N_21956,N_19705,N_19504);
xor U21957 (N_21957,N_19671,N_20805);
and U21958 (N_21958,N_20520,N_20082);
nor U21959 (N_21959,N_20163,N_20461);
or U21960 (N_21960,N_19751,N_20216);
nand U21961 (N_21961,N_19744,N_20961);
or U21962 (N_21962,N_20014,N_19904);
xor U21963 (N_21963,N_20107,N_19913);
and U21964 (N_21964,N_19896,N_20230);
xor U21965 (N_21965,N_19769,N_20000);
nor U21966 (N_21966,N_19845,N_19836);
or U21967 (N_21967,N_19746,N_20062);
xor U21968 (N_21968,N_20321,N_20425);
nand U21969 (N_21969,N_20900,N_19931);
xnor U21970 (N_21970,N_20198,N_19897);
and U21971 (N_21971,N_20430,N_19705);
or U21972 (N_21972,N_20956,N_19666);
nor U21973 (N_21973,N_20570,N_20554);
xor U21974 (N_21974,N_20180,N_20772);
or U21975 (N_21975,N_20546,N_20223);
nand U21976 (N_21976,N_19985,N_20116);
nand U21977 (N_21977,N_20704,N_20035);
or U21978 (N_21978,N_19582,N_20380);
xor U21979 (N_21979,N_19789,N_20197);
or U21980 (N_21980,N_19757,N_20846);
xor U21981 (N_21981,N_19961,N_20671);
nand U21982 (N_21982,N_20114,N_20247);
nand U21983 (N_21983,N_19911,N_20761);
xor U21984 (N_21984,N_19996,N_19943);
or U21985 (N_21985,N_20925,N_20261);
nand U21986 (N_21986,N_20091,N_20585);
xor U21987 (N_21987,N_20415,N_19722);
and U21988 (N_21988,N_19553,N_20282);
and U21989 (N_21989,N_20617,N_20505);
nor U21990 (N_21990,N_19755,N_20714);
xnor U21991 (N_21991,N_19687,N_20095);
or U21992 (N_21992,N_19572,N_20736);
nand U21993 (N_21993,N_19613,N_19816);
and U21994 (N_21994,N_20250,N_19632);
xor U21995 (N_21995,N_20408,N_20907);
nand U21996 (N_21996,N_20364,N_20360);
or U21997 (N_21997,N_20581,N_19864);
xnor U21998 (N_21998,N_20252,N_19804);
nand U21999 (N_21999,N_20613,N_20684);
and U22000 (N_22000,N_20873,N_19924);
nor U22001 (N_22001,N_20997,N_20360);
nor U22002 (N_22002,N_20049,N_20992);
and U22003 (N_22003,N_19623,N_20080);
nand U22004 (N_22004,N_19547,N_20315);
or U22005 (N_22005,N_20275,N_20670);
or U22006 (N_22006,N_20065,N_20995);
and U22007 (N_22007,N_19944,N_19945);
xor U22008 (N_22008,N_20019,N_19939);
xor U22009 (N_22009,N_19716,N_20274);
nand U22010 (N_22010,N_20471,N_20186);
nor U22011 (N_22011,N_20230,N_20580);
xnor U22012 (N_22012,N_19735,N_20172);
nand U22013 (N_22013,N_19800,N_19591);
and U22014 (N_22014,N_19647,N_20463);
xor U22015 (N_22015,N_20012,N_20683);
or U22016 (N_22016,N_20285,N_20972);
or U22017 (N_22017,N_20978,N_20489);
or U22018 (N_22018,N_19939,N_20029);
or U22019 (N_22019,N_19587,N_20206);
and U22020 (N_22020,N_20685,N_20219);
nor U22021 (N_22021,N_20814,N_20800);
or U22022 (N_22022,N_20614,N_20958);
and U22023 (N_22023,N_19590,N_19585);
and U22024 (N_22024,N_20537,N_20908);
xor U22025 (N_22025,N_20532,N_19506);
nand U22026 (N_22026,N_19843,N_20792);
or U22027 (N_22027,N_19520,N_20461);
nand U22028 (N_22028,N_19574,N_20349);
xnor U22029 (N_22029,N_20287,N_20721);
and U22030 (N_22030,N_19523,N_19926);
and U22031 (N_22031,N_20761,N_20483);
nand U22032 (N_22032,N_19876,N_20508);
xnor U22033 (N_22033,N_19538,N_20071);
xor U22034 (N_22034,N_19505,N_20321);
and U22035 (N_22035,N_20800,N_20843);
nand U22036 (N_22036,N_19648,N_20885);
and U22037 (N_22037,N_20506,N_20901);
xnor U22038 (N_22038,N_20946,N_19607);
xnor U22039 (N_22039,N_20859,N_19887);
nor U22040 (N_22040,N_20919,N_19756);
nand U22041 (N_22041,N_20027,N_19903);
and U22042 (N_22042,N_19727,N_19921);
nand U22043 (N_22043,N_19953,N_19735);
nand U22044 (N_22044,N_20945,N_19715);
or U22045 (N_22045,N_20098,N_20486);
or U22046 (N_22046,N_20350,N_20214);
or U22047 (N_22047,N_20545,N_20670);
or U22048 (N_22048,N_19805,N_20931);
nand U22049 (N_22049,N_20683,N_20880);
or U22050 (N_22050,N_20022,N_19789);
and U22051 (N_22051,N_19715,N_19864);
or U22052 (N_22052,N_20517,N_20344);
nor U22053 (N_22053,N_19628,N_19583);
nand U22054 (N_22054,N_19743,N_20698);
or U22055 (N_22055,N_19812,N_20926);
nor U22056 (N_22056,N_19987,N_19866);
and U22057 (N_22057,N_19997,N_20732);
nor U22058 (N_22058,N_20965,N_19816);
nor U22059 (N_22059,N_20419,N_20643);
or U22060 (N_22060,N_19797,N_20071);
or U22061 (N_22061,N_20838,N_19785);
xnor U22062 (N_22062,N_19676,N_19736);
and U22063 (N_22063,N_20370,N_20699);
xnor U22064 (N_22064,N_20147,N_19803);
or U22065 (N_22065,N_19969,N_20243);
nand U22066 (N_22066,N_20008,N_20303);
nand U22067 (N_22067,N_19555,N_20019);
nor U22068 (N_22068,N_19841,N_20440);
nor U22069 (N_22069,N_20388,N_20889);
or U22070 (N_22070,N_19940,N_20388);
nor U22071 (N_22071,N_19582,N_20598);
nor U22072 (N_22072,N_20185,N_19517);
xnor U22073 (N_22073,N_19828,N_20490);
xor U22074 (N_22074,N_20758,N_19519);
nand U22075 (N_22075,N_20453,N_19518);
nor U22076 (N_22076,N_19640,N_20343);
or U22077 (N_22077,N_19817,N_19910);
xor U22078 (N_22078,N_20838,N_20961);
or U22079 (N_22079,N_20616,N_20838);
and U22080 (N_22080,N_19828,N_20637);
or U22081 (N_22081,N_20794,N_19966);
nand U22082 (N_22082,N_19692,N_20031);
and U22083 (N_22083,N_19649,N_20828);
and U22084 (N_22084,N_20793,N_20088);
and U22085 (N_22085,N_20761,N_20259);
nor U22086 (N_22086,N_20299,N_19732);
nand U22087 (N_22087,N_20792,N_20576);
and U22088 (N_22088,N_20377,N_19759);
and U22089 (N_22089,N_19574,N_20140);
xnor U22090 (N_22090,N_20827,N_20706);
xnor U22091 (N_22091,N_19966,N_20236);
xnor U22092 (N_22092,N_19700,N_19743);
and U22093 (N_22093,N_20909,N_20695);
nor U22094 (N_22094,N_20331,N_20103);
nor U22095 (N_22095,N_20446,N_20265);
nor U22096 (N_22096,N_19800,N_20741);
and U22097 (N_22097,N_20731,N_20557);
nor U22098 (N_22098,N_19574,N_19650);
xor U22099 (N_22099,N_20297,N_20731);
nor U22100 (N_22100,N_20780,N_19906);
nand U22101 (N_22101,N_20416,N_20616);
and U22102 (N_22102,N_20721,N_19991);
and U22103 (N_22103,N_19513,N_20367);
nand U22104 (N_22104,N_19656,N_20194);
xnor U22105 (N_22105,N_19705,N_20367);
or U22106 (N_22106,N_20288,N_20964);
nand U22107 (N_22107,N_20668,N_20565);
nand U22108 (N_22108,N_20087,N_19706);
xor U22109 (N_22109,N_20608,N_20217);
nor U22110 (N_22110,N_20822,N_20652);
xnor U22111 (N_22111,N_19559,N_20611);
nor U22112 (N_22112,N_19586,N_19846);
nor U22113 (N_22113,N_20859,N_20983);
nand U22114 (N_22114,N_20696,N_20032);
nand U22115 (N_22115,N_20905,N_20944);
xor U22116 (N_22116,N_19918,N_19569);
nor U22117 (N_22117,N_19623,N_19584);
nor U22118 (N_22118,N_20080,N_19526);
and U22119 (N_22119,N_20390,N_20001);
xor U22120 (N_22120,N_19644,N_19945);
nand U22121 (N_22121,N_19869,N_20258);
nand U22122 (N_22122,N_20138,N_19614);
and U22123 (N_22123,N_19860,N_19998);
or U22124 (N_22124,N_20374,N_20168);
nor U22125 (N_22125,N_20282,N_20018);
xor U22126 (N_22126,N_19731,N_19952);
nor U22127 (N_22127,N_20197,N_20793);
nand U22128 (N_22128,N_20556,N_19629);
nand U22129 (N_22129,N_20320,N_20537);
or U22130 (N_22130,N_20027,N_20540);
xnor U22131 (N_22131,N_20793,N_20639);
nand U22132 (N_22132,N_19677,N_20772);
nor U22133 (N_22133,N_20743,N_20878);
nand U22134 (N_22134,N_20961,N_20964);
and U22135 (N_22135,N_19866,N_20489);
nand U22136 (N_22136,N_20175,N_19855);
nor U22137 (N_22137,N_19965,N_20159);
nor U22138 (N_22138,N_20030,N_19653);
nand U22139 (N_22139,N_19608,N_19589);
or U22140 (N_22140,N_20773,N_20402);
or U22141 (N_22141,N_19502,N_20484);
and U22142 (N_22142,N_19720,N_20919);
or U22143 (N_22143,N_20579,N_20517);
xnor U22144 (N_22144,N_20628,N_19759);
and U22145 (N_22145,N_19909,N_19698);
or U22146 (N_22146,N_20958,N_20225);
nor U22147 (N_22147,N_20196,N_20869);
and U22148 (N_22148,N_20295,N_19512);
and U22149 (N_22149,N_19779,N_19683);
and U22150 (N_22150,N_20388,N_19968);
or U22151 (N_22151,N_20601,N_20708);
and U22152 (N_22152,N_20889,N_20899);
xnor U22153 (N_22153,N_20245,N_19561);
nor U22154 (N_22154,N_20044,N_19630);
nor U22155 (N_22155,N_20177,N_19687);
and U22156 (N_22156,N_19838,N_20497);
nor U22157 (N_22157,N_20362,N_20972);
nor U22158 (N_22158,N_19680,N_19605);
nor U22159 (N_22159,N_20471,N_20738);
and U22160 (N_22160,N_19574,N_19522);
nor U22161 (N_22161,N_20507,N_20623);
xnor U22162 (N_22162,N_20543,N_20902);
nand U22163 (N_22163,N_19994,N_20150);
or U22164 (N_22164,N_20214,N_20450);
xnor U22165 (N_22165,N_20330,N_20613);
or U22166 (N_22166,N_19859,N_19903);
and U22167 (N_22167,N_19714,N_20871);
nor U22168 (N_22168,N_19623,N_20055);
or U22169 (N_22169,N_20330,N_19908);
nor U22170 (N_22170,N_19888,N_19668);
nor U22171 (N_22171,N_20520,N_20286);
xnor U22172 (N_22172,N_20276,N_20145);
nand U22173 (N_22173,N_19719,N_20292);
and U22174 (N_22174,N_20774,N_20822);
nor U22175 (N_22175,N_19943,N_20794);
xnor U22176 (N_22176,N_20785,N_19799);
nand U22177 (N_22177,N_20714,N_19524);
nand U22178 (N_22178,N_19820,N_20975);
nor U22179 (N_22179,N_19544,N_20939);
xor U22180 (N_22180,N_19964,N_20290);
nor U22181 (N_22181,N_20069,N_20185);
nand U22182 (N_22182,N_20050,N_20024);
and U22183 (N_22183,N_20489,N_19547);
nor U22184 (N_22184,N_20417,N_19881);
xnor U22185 (N_22185,N_19684,N_20678);
nand U22186 (N_22186,N_20795,N_20543);
nand U22187 (N_22187,N_19561,N_20648);
and U22188 (N_22188,N_20501,N_20275);
and U22189 (N_22189,N_20781,N_20473);
nand U22190 (N_22190,N_20199,N_20230);
and U22191 (N_22191,N_20966,N_20309);
xnor U22192 (N_22192,N_19648,N_20294);
or U22193 (N_22193,N_19796,N_20150);
nand U22194 (N_22194,N_20622,N_20886);
xor U22195 (N_22195,N_20430,N_20747);
xor U22196 (N_22196,N_20612,N_19728);
or U22197 (N_22197,N_20442,N_20906);
nor U22198 (N_22198,N_20964,N_20779);
or U22199 (N_22199,N_19776,N_20085);
and U22200 (N_22200,N_20332,N_20029);
nand U22201 (N_22201,N_19596,N_20285);
or U22202 (N_22202,N_20091,N_20338);
and U22203 (N_22203,N_20072,N_20206);
xnor U22204 (N_22204,N_20236,N_20206);
nor U22205 (N_22205,N_20704,N_19836);
and U22206 (N_22206,N_20644,N_20026);
or U22207 (N_22207,N_19919,N_20355);
and U22208 (N_22208,N_20646,N_19536);
xnor U22209 (N_22209,N_20632,N_19937);
xor U22210 (N_22210,N_19660,N_20449);
nand U22211 (N_22211,N_19667,N_20852);
or U22212 (N_22212,N_20749,N_20328);
or U22213 (N_22213,N_20127,N_20852);
or U22214 (N_22214,N_19569,N_20368);
xor U22215 (N_22215,N_20235,N_19981);
xnor U22216 (N_22216,N_20620,N_20661);
xnor U22217 (N_22217,N_19952,N_19932);
and U22218 (N_22218,N_19688,N_19820);
or U22219 (N_22219,N_20346,N_20841);
and U22220 (N_22220,N_19680,N_20596);
nor U22221 (N_22221,N_19552,N_20235);
or U22222 (N_22222,N_19814,N_20116);
and U22223 (N_22223,N_20885,N_20505);
xor U22224 (N_22224,N_20593,N_19814);
nand U22225 (N_22225,N_19814,N_19583);
nand U22226 (N_22226,N_20554,N_20579);
nand U22227 (N_22227,N_20193,N_20116);
or U22228 (N_22228,N_20517,N_20979);
nor U22229 (N_22229,N_20994,N_19866);
xnor U22230 (N_22230,N_20271,N_20684);
nand U22231 (N_22231,N_19651,N_20990);
or U22232 (N_22232,N_20786,N_19875);
nor U22233 (N_22233,N_20715,N_19621);
or U22234 (N_22234,N_20992,N_19835);
nand U22235 (N_22235,N_19549,N_20739);
nand U22236 (N_22236,N_20806,N_20265);
xor U22237 (N_22237,N_20854,N_19576);
xnor U22238 (N_22238,N_20709,N_20121);
or U22239 (N_22239,N_20036,N_20858);
nor U22240 (N_22240,N_20294,N_19549);
or U22241 (N_22241,N_19897,N_20320);
xor U22242 (N_22242,N_19796,N_19851);
and U22243 (N_22243,N_19806,N_20860);
or U22244 (N_22244,N_20865,N_20857);
and U22245 (N_22245,N_19593,N_19934);
xor U22246 (N_22246,N_19582,N_19741);
nor U22247 (N_22247,N_19755,N_20351);
nor U22248 (N_22248,N_19841,N_19960);
xor U22249 (N_22249,N_20289,N_20325);
or U22250 (N_22250,N_20272,N_19842);
nand U22251 (N_22251,N_20076,N_19965);
xor U22252 (N_22252,N_19824,N_20740);
or U22253 (N_22253,N_20935,N_20151);
nor U22254 (N_22254,N_19886,N_19948);
nand U22255 (N_22255,N_20733,N_20844);
or U22256 (N_22256,N_20835,N_20562);
and U22257 (N_22257,N_19505,N_20606);
or U22258 (N_22258,N_20451,N_20220);
xor U22259 (N_22259,N_20210,N_19714);
and U22260 (N_22260,N_20927,N_20736);
nand U22261 (N_22261,N_20612,N_20748);
nand U22262 (N_22262,N_20424,N_20292);
and U22263 (N_22263,N_20774,N_20390);
or U22264 (N_22264,N_20459,N_20380);
xnor U22265 (N_22265,N_20325,N_20082);
xnor U22266 (N_22266,N_19880,N_20327);
or U22267 (N_22267,N_20272,N_19545);
xor U22268 (N_22268,N_20438,N_20372);
nand U22269 (N_22269,N_20452,N_20704);
or U22270 (N_22270,N_19625,N_20496);
and U22271 (N_22271,N_20067,N_19832);
nand U22272 (N_22272,N_20956,N_19617);
xnor U22273 (N_22273,N_19610,N_20033);
xnor U22274 (N_22274,N_19785,N_20389);
xnor U22275 (N_22275,N_20177,N_20158);
nor U22276 (N_22276,N_20773,N_20376);
nor U22277 (N_22277,N_19605,N_20220);
nand U22278 (N_22278,N_20180,N_19571);
and U22279 (N_22279,N_20037,N_19760);
or U22280 (N_22280,N_19561,N_19766);
nand U22281 (N_22281,N_19974,N_20315);
nand U22282 (N_22282,N_20347,N_19909);
or U22283 (N_22283,N_20081,N_20824);
nand U22284 (N_22284,N_19804,N_19923);
and U22285 (N_22285,N_20256,N_19700);
nor U22286 (N_22286,N_20955,N_20564);
nand U22287 (N_22287,N_20313,N_20812);
or U22288 (N_22288,N_19880,N_19702);
nor U22289 (N_22289,N_20012,N_19700);
nor U22290 (N_22290,N_20127,N_20441);
or U22291 (N_22291,N_20698,N_20706);
xnor U22292 (N_22292,N_20567,N_20191);
xor U22293 (N_22293,N_20775,N_20142);
nor U22294 (N_22294,N_19787,N_19611);
nor U22295 (N_22295,N_19648,N_20748);
and U22296 (N_22296,N_20290,N_19577);
or U22297 (N_22297,N_20964,N_20080);
nor U22298 (N_22298,N_20917,N_20462);
or U22299 (N_22299,N_20057,N_19668);
and U22300 (N_22300,N_20589,N_20023);
nor U22301 (N_22301,N_19983,N_20366);
nor U22302 (N_22302,N_20356,N_19580);
nand U22303 (N_22303,N_20263,N_19623);
nor U22304 (N_22304,N_19778,N_20212);
or U22305 (N_22305,N_20614,N_19896);
or U22306 (N_22306,N_20215,N_20093);
or U22307 (N_22307,N_20867,N_20963);
xnor U22308 (N_22308,N_19738,N_20924);
xor U22309 (N_22309,N_19576,N_19517);
nand U22310 (N_22310,N_20099,N_20749);
and U22311 (N_22311,N_20877,N_20797);
nand U22312 (N_22312,N_20504,N_19551);
nand U22313 (N_22313,N_19973,N_20495);
nand U22314 (N_22314,N_20368,N_19913);
and U22315 (N_22315,N_19931,N_20263);
nor U22316 (N_22316,N_20580,N_19604);
nand U22317 (N_22317,N_20105,N_19871);
or U22318 (N_22318,N_19630,N_19677);
or U22319 (N_22319,N_20695,N_19855);
and U22320 (N_22320,N_19994,N_20340);
nand U22321 (N_22321,N_20592,N_20152);
nor U22322 (N_22322,N_20899,N_20022);
nand U22323 (N_22323,N_20379,N_20127);
nand U22324 (N_22324,N_20451,N_20394);
or U22325 (N_22325,N_19828,N_20124);
nor U22326 (N_22326,N_20284,N_20147);
or U22327 (N_22327,N_19792,N_20112);
nand U22328 (N_22328,N_20785,N_20581);
or U22329 (N_22329,N_20401,N_20912);
nor U22330 (N_22330,N_20304,N_20002);
or U22331 (N_22331,N_20797,N_20296);
nand U22332 (N_22332,N_20696,N_20034);
xor U22333 (N_22333,N_20268,N_19988);
nand U22334 (N_22334,N_19633,N_20833);
nand U22335 (N_22335,N_20681,N_20672);
nand U22336 (N_22336,N_20203,N_19678);
or U22337 (N_22337,N_20125,N_20730);
nand U22338 (N_22338,N_19838,N_20931);
or U22339 (N_22339,N_20845,N_19716);
xnor U22340 (N_22340,N_19731,N_20226);
or U22341 (N_22341,N_20441,N_20219);
xnor U22342 (N_22342,N_20890,N_19580);
xor U22343 (N_22343,N_19742,N_19739);
or U22344 (N_22344,N_20160,N_20007);
nand U22345 (N_22345,N_20615,N_20991);
nor U22346 (N_22346,N_20595,N_20426);
or U22347 (N_22347,N_20928,N_19629);
or U22348 (N_22348,N_19923,N_19672);
or U22349 (N_22349,N_20067,N_20502);
nor U22350 (N_22350,N_20568,N_20972);
xnor U22351 (N_22351,N_20059,N_19994);
xor U22352 (N_22352,N_20717,N_20123);
nor U22353 (N_22353,N_19869,N_20205);
xnor U22354 (N_22354,N_19861,N_19947);
xnor U22355 (N_22355,N_19796,N_20526);
nor U22356 (N_22356,N_20228,N_20159);
nor U22357 (N_22357,N_19988,N_19994);
or U22358 (N_22358,N_19636,N_19834);
xnor U22359 (N_22359,N_20650,N_20355);
and U22360 (N_22360,N_20621,N_20288);
and U22361 (N_22361,N_20353,N_20486);
nand U22362 (N_22362,N_20381,N_19912);
and U22363 (N_22363,N_20599,N_19881);
nand U22364 (N_22364,N_19627,N_20209);
or U22365 (N_22365,N_20105,N_20856);
nand U22366 (N_22366,N_20681,N_20043);
xor U22367 (N_22367,N_20357,N_19879);
xnor U22368 (N_22368,N_20276,N_19533);
nor U22369 (N_22369,N_20376,N_20137);
or U22370 (N_22370,N_20512,N_19527);
nand U22371 (N_22371,N_19644,N_20079);
and U22372 (N_22372,N_19776,N_20963);
nor U22373 (N_22373,N_20257,N_20138);
nor U22374 (N_22374,N_20129,N_19904);
nor U22375 (N_22375,N_19588,N_20234);
nand U22376 (N_22376,N_20405,N_20944);
xnor U22377 (N_22377,N_19774,N_19973);
nand U22378 (N_22378,N_19560,N_20495);
xor U22379 (N_22379,N_20408,N_20697);
or U22380 (N_22380,N_20254,N_20011);
or U22381 (N_22381,N_20017,N_19860);
nand U22382 (N_22382,N_19834,N_19852);
or U22383 (N_22383,N_19997,N_20540);
nor U22384 (N_22384,N_20023,N_20116);
or U22385 (N_22385,N_20463,N_20541);
or U22386 (N_22386,N_19525,N_19626);
nor U22387 (N_22387,N_20749,N_20774);
or U22388 (N_22388,N_20489,N_19601);
or U22389 (N_22389,N_19553,N_20907);
nand U22390 (N_22390,N_19579,N_19999);
xnor U22391 (N_22391,N_19648,N_20708);
nor U22392 (N_22392,N_19550,N_19855);
and U22393 (N_22393,N_19924,N_19695);
xor U22394 (N_22394,N_20182,N_19680);
nor U22395 (N_22395,N_19755,N_19922);
nand U22396 (N_22396,N_19625,N_19982);
and U22397 (N_22397,N_20783,N_20130);
nand U22398 (N_22398,N_20089,N_20641);
nand U22399 (N_22399,N_19697,N_20145);
nand U22400 (N_22400,N_20751,N_19688);
and U22401 (N_22401,N_19710,N_20176);
xor U22402 (N_22402,N_20362,N_20153);
and U22403 (N_22403,N_20215,N_19947);
nor U22404 (N_22404,N_20448,N_19983);
xnor U22405 (N_22405,N_20015,N_19734);
and U22406 (N_22406,N_19854,N_20462);
and U22407 (N_22407,N_19920,N_20282);
nand U22408 (N_22408,N_20127,N_19771);
xor U22409 (N_22409,N_20611,N_20600);
nor U22410 (N_22410,N_20943,N_20304);
xnor U22411 (N_22411,N_20188,N_20145);
and U22412 (N_22412,N_19961,N_20774);
nand U22413 (N_22413,N_19625,N_19757);
and U22414 (N_22414,N_19938,N_20439);
nand U22415 (N_22415,N_19973,N_20670);
nor U22416 (N_22416,N_20041,N_20741);
and U22417 (N_22417,N_20720,N_19808);
nand U22418 (N_22418,N_20680,N_20326);
xor U22419 (N_22419,N_20715,N_20030);
and U22420 (N_22420,N_20112,N_19580);
nand U22421 (N_22421,N_20575,N_19679);
nand U22422 (N_22422,N_20708,N_20794);
nand U22423 (N_22423,N_20173,N_20745);
nor U22424 (N_22424,N_20070,N_20596);
nand U22425 (N_22425,N_19991,N_20041);
nand U22426 (N_22426,N_20098,N_19978);
nor U22427 (N_22427,N_19727,N_20425);
or U22428 (N_22428,N_20006,N_20597);
nor U22429 (N_22429,N_19770,N_19535);
and U22430 (N_22430,N_19715,N_20648);
xor U22431 (N_22431,N_19505,N_20167);
xnor U22432 (N_22432,N_19539,N_19966);
or U22433 (N_22433,N_19927,N_19503);
xnor U22434 (N_22434,N_19823,N_20913);
nor U22435 (N_22435,N_20553,N_20727);
and U22436 (N_22436,N_19701,N_20132);
or U22437 (N_22437,N_20292,N_20940);
or U22438 (N_22438,N_20846,N_20709);
nand U22439 (N_22439,N_20856,N_19883);
nand U22440 (N_22440,N_19978,N_20272);
nand U22441 (N_22441,N_20383,N_20142);
and U22442 (N_22442,N_20094,N_20664);
and U22443 (N_22443,N_20535,N_20460);
or U22444 (N_22444,N_20108,N_20023);
xor U22445 (N_22445,N_20416,N_20375);
xnor U22446 (N_22446,N_20142,N_19883);
nand U22447 (N_22447,N_19876,N_20413);
nor U22448 (N_22448,N_20057,N_20265);
or U22449 (N_22449,N_20191,N_20473);
nand U22450 (N_22450,N_19812,N_20207);
nand U22451 (N_22451,N_20134,N_20628);
and U22452 (N_22452,N_19530,N_20876);
xnor U22453 (N_22453,N_20440,N_19816);
nor U22454 (N_22454,N_19571,N_20991);
nor U22455 (N_22455,N_19575,N_20206);
or U22456 (N_22456,N_20687,N_19965);
xnor U22457 (N_22457,N_19903,N_20746);
and U22458 (N_22458,N_20812,N_20153);
nand U22459 (N_22459,N_20561,N_20067);
xor U22460 (N_22460,N_19722,N_19681);
xor U22461 (N_22461,N_20093,N_19619);
and U22462 (N_22462,N_20196,N_20718);
nand U22463 (N_22463,N_19645,N_20716);
xor U22464 (N_22464,N_20581,N_20770);
or U22465 (N_22465,N_19992,N_20430);
and U22466 (N_22466,N_20762,N_20386);
and U22467 (N_22467,N_19502,N_20997);
or U22468 (N_22468,N_19735,N_20386);
nor U22469 (N_22469,N_20579,N_20432);
xnor U22470 (N_22470,N_19709,N_19915);
and U22471 (N_22471,N_19681,N_20686);
nor U22472 (N_22472,N_19619,N_19704);
nand U22473 (N_22473,N_20222,N_20814);
nand U22474 (N_22474,N_20965,N_19971);
xor U22475 (N_22475,N_20963,N_19996);
xnor U22476 (N_22476,N_20635,N_19535);
or U22477 (N_22477,N_20139,N_20169);
and U22478 (N_22478,N_19580,N_20354);
nand U22479 (N_22479,N_20119,N_20813);
and U22480 (N_22480,N_20289,N_20588);
xor U22481 (N_22481,N_20228,N_19763);
nand U22482 (N_22482,N_20460,N_19975);
nor U22483 (N_22483,N_20533,N_20386);
nand U22484 (N_22484,N_20543,N_20962);
or U22485 (N_22485,N_20456,N_20629);
nand U22486 (N_22486,N_19512,N_20089);
or U22487 (N_22487,N_20516,N_20095);
and U22488 (N_22488,N_19681,N_20942);
or U22489 (N_22489,N_20400,N_20544);
xnor U22490 (N_22490,N_19544,N_20955);
or U22491 (N_22491,N_20080,N_20392);
xnor U22492 (N_22492,N_19618,N_20948);
xnor U22493 (N_22493,N_20487,N_20243);
and U22494 (N_22494,N_19569,N_20358);
nor U22495 (N_22495,N_20827,N_20481);
xor U22496 (N_22496,N_20433,N_19844);
xnor U22497 (N_22497,N_19801,N_20411);
xor U22498 (N_22498,N_19568,N_19633);
or U22499 (N_22499,N_20865,N_19810);
or U22500 (N_22500,N_21983,N_21261);
xor U22501 (N_22501,N_21147,N_22111);
and U22502 (N_22502,N_22179,N_21195);
nor U22503 (N_22503,N_22182,N_21306);
or U22504 (N_22504,N_22354,N_21839);
nor U22505 (N_22505,N_21146,N_22462);
nand U22506 (N_22506,N_22107,N_21116);
nor U22507 (N_22507,N_21810,N_21965);
xor U22508 (N_22508,N_21605,N_21363);
nor U22509 (N_22509,N_21454,N_22408);
or U22510 (N_22510,N_21703,N_21968);
nand U22511 (N_22511,N_22250,N_21148);
nand U22512 (N_22512,N_21291,N_22460);
nand U22513 (N_22513,N_21027,N_21155);
or U22514 (N_22514,N_21964,N_21044);
or U22515 (N_22515,N_21534,N_21949);
nand U22516 (N_22516,N_21866,N_21446);
or U22517 (N_22517,N_22450,N_21380);
xor U22518 (N_22518,N_21565,N_21159);
and U22519 (N_22519,N_21936,N_22007);
nor U22520 (N_22520,N_21880,N_22225);
xnor U22521 (N_22521,N_22164,N_22289);
nor U22522 (N_22522,N_22132,N_21741);
nor U22523 (N_22523,N_21466,N_21327);
or U22524 (N_22524,N_21761,N_21873);
xnor U22525 (N_22525,N_21742,N_22487);
nor U22526 (N_22526,N_21387,N_21416);
or U22527 (N_22527,N_21900,N_22196);
nor U22528 (N_22528,N_21394,N_21831);
xnor U22529 (N_22529,N_22171,N_21995);
xnor U22530 (N_22530,N_22029,N_21141);
or U22531 (N_22531,N_21897,N_21135);
and U22532 (N_22532,N_21039,N_21067);
nor U22533 (N_22533,N_21792,N_22037);
or U22534 (N_22534,N_21802,N_21302);
and U22535 (N_22535,N_22229,N_21206);
or U22536 (N_22536,N_22168,N_21844);
or U22537 (N_22537,N_21209,N_21314);
or U22538 (N_22538,N_21561,N_21865);
nor U22539 (N_22539,N_22180,N_21511);
xnor U22540 (N_22540,N_22078,N_22358);
nor U22541 (N_22541,N_22451,N_21988);
or U22542 (N_22542,N_22165,N_21033);
and U22543 (N_22543,N_21715,N_21684);
or U22544 (N_22544,N_21568,N_21485);
xnor U22545 (N_22545,N_21219,N_21053);
nand U22546 (N_22546,N_21932,N_22334);
and U22547 (N_22547,N_21422,N_21819);
or U22548 (N_22548,N_22436,N_22474);
nand U22549 (N_22549,N_21107,N_21836);
nand U22550 (N_22550,N_21309,N_22255);
xor U22551 (N_22551,N_21590,N_22243);
nor U22552 (N_22552,N_21137,N_21992);
or U22553 (N_22553,N_21971,N_21688);
nand U22554 (N_22554,N_21961,N_22060);
xnor U22555 (N_22555,N_21267,N_21718);
or U22556 (N_22556,N_22300,N_21097);
nor U22557 (N_22557,N_21073,N_22323);
or U22558 (N_22558,N_21700,N_22430);
xnor U22559 (N_22559,N_21056,N_21922);
nor U22560 (N_22560,N_21878,N_22001);
xor U22561 (N_22561,N_22072,N_22293);
and U22562 (N_22562,N_21627,N_22195);
nand U22563 (N_22563,N_21734,N_21243);
nand U22564 (N_22564,N_22062,N_22480);
nor U22565 (N_22565,N_21987,N_22011);
and U22566 (N_22566,N_21164,N_21042);
or U22567 (N_22567,N_21224,N_22110);
nand U22568 (N_22568,N_21917,N_21772);
or U22569 (N_22569,N_21007,N_21708);
xor U22570 (N_22570,N_21910,N_21052);
xor U22571 (N_22571,N_21115,N_21445);
xnor U22572 (N_22572,N_22096,N_22493);
nor U22573 (N_22573,N_21066,N_21040);
or U22574 (N_22574,N_21307,N_22264);
nand U22575 (N_22575,N_21528,N_21239);
nor U22576 (N_22576,N_21990,N_22076);
and U22577 (N_22577,N_21533,N_21925);
or U22578 (N_22578,N_21664,N_22377);
nor U22579 (N_22579,N_21048,N_21784);
or U22580 (N_22580,N_21730,N_21208);
xor U22581 (N_22581,N_22280,N_21101);
xor U22582 (N_22582,N_22237,N_22105);
and U22583 (N_22583,N_22321,N_21808);
xnor U22584 (N_22584,N_22461,N_22283);
or U22585 (N_22585,N_21109,N_22442);
or U22586 (N_22586,N_21414,N_22476);
xnor U22587 (N_22587,N_22342,N_21942);
or U22588 (N_22588,N_22371,N_21420);
nand U22589 (N_22589,N_21202,N_22205);
nand U22590 (N_22590,N_21524,N_21439);
nand U22591 (N_22591,N_22120,N_21061);
nand U22592 (N_22592,N_21547,N_21737);
and U22593 (N_22593,N_21712,N_21694);
and U22594 (N_22594,N_21399,N_22138);
nand U22595 (N_22595,N_21670,N_21330);
nor U22596 (N_22596,N_21038,N_21832);
xnor U22597 (N_22597,N_21080,N_21704);
nand U22598 (N_22598,N_21283,N_21723);
and U22599 (N_22599,N_21889,N_21129);
or U22600 (N_22600,N_22005,N_22221);
xor U22601 (N_22601,N_21525,N_21360);
nor U22602 (N_22602,N_21699,N_22348);
xor U22603 (N_22603,N_21523,N_21957);
xor U22604 (N_22604,N_21319,N_21478);
nor U22605 (N_22605,N_21138,N_22340);
nand U22606 (N_22606,N_21111,N_21530);
nor U22607 (N_22607,N_21002,N_22343);
or U22608 (N_22608,N_21941,N_21368);
nand U22609 (N_22609,N_22475,N_21361);
and U22610 (N_22610,N_21709,N_21848);
and U22611 (N_22611,N_22213,N_21672);
or U22612 (N_22612,N_22421,N_21725);
nor U22613 (N_22613,N_21595,N_21176);
nand U22614 (N_22614,N_21807,N_21816);
xnor U22615 (N_22615,N_21482,N_21496);
nor U22616 (N_22616,N_22071,N_21133);
nand U22617 (N_22617,N_21170,N_22208);
nor U22618 (N_22618,N_21321,N_21365);
xnor U22619 (N_22619,N_21008,N_21434);
and U22620 (N_22620,N_21218,N_22291);
nand U22621 (N_22621,N_21271,N_21674);
or U22622 (N_22622,N_21915,N_21163);
nand U22623 (N_22623,N_21788,N_22484);
nor U22624 (N_22624,N_22330,N_21213);
or U22625 (N_22625,N_21787,N_21877);
or U22626 (N_22626,N_22329,N_21275);
nand U22627 (N_22627,N_21721,N_22028);
nor U22628 (N_22628,N_22080,N_22376);
nor U22629 (N_22629,N_21642,N_22126);
or U22630 (N_22630,N_21151,N_22178);
nand U22631 (N_22631,N_21102,N_21671);
nor U22632 (N_22632,N_22081,N_22274);
or U22633 (N_22633,N_22425,N_21356);
or U22634 (N_22634,N_22315,N_22337);
nand U22635 (N_22635,N_21564,N_22392);
nand U22636 (N_22636,N_22458,N_21079);
xor U22637 (N_22637,N_22279,N_21789);
and U22638 (N_22638,N_22419,N_21333);
or U22639 (N_22639,N_21953,N_21045);
or U22640 (N_22640,N_21967,N_21397);
xnor U22641 (N_22641,N_21405,N_21841);
or U22642 (N_22642,N_21276,N_21935);
xnor U22643 (N_22643,N_21894,N_22322);
nand U22644 (N_22644,N_21659,N_22478);
and U22645 (N_22645,N_21903,N_22135);
or U22646 (N_22646,N_22372,N_21475);
and U22647 (N_22647,N_22440,N_21887);
or U22648 (N_22648,N_22370,N_21367);
nand U22649 (N_22649,N_21090,N_22079);
nor U22650 (N_22650,N_21049,N_21654);
nand U22651 (N_22651,N_21775,N_22252);
nand U22652 (N_22652,N_21152,N_22035);
and U22653 (N_22653,N_22150,N_21635);
or U22654 (N_22654,N_21824,N_21046);
nor U22655 (N_22655,N_21803,N_21606);
xnor U22656 (N_22656,N_22361,N_21277);
xor U22657 (N_22657,N_22085,N_21875);
and U22658 (N_22658,N_21255,N_21054);
or U22659 (N_22659,N_21926,N_22021);
or U22660 (N_22660,N_21172,N_21187);
xnor U22661 (N_22661,N_21300,N_21881);
or U22662 (N_22662,N_21489,N_21041);
or U22663 (N_22663,N_21329,N_21753);
xor U22664 (N_22664,N_21411,N_21144);
xnor U22665 (N_22665,N_22015,N_21854);
nand U22666 (N_22666,N_22006,N_21354);
nor U22667 (N_22667,N_22346,N_21604);
xor U22668 (N_22668,N_22134,N_21641);
xor U22669 (N_22669,N_22039,N_21242);
and U22670 (N_22670,N_21668,N_21452);
nor U22671 (N_22671,N_21216,N_21117);
nor U22672 (N_22672,N_22122,N_22384);
xor U22673 (N_22673,N_21143,N_22486);
and U22674 (N_22674,N_22143,N_21015);
xor U22675 (N_22675,N_21252,N_21826);
and U22676 (N_22676,N_21843,N_22103);
nor U22677 (N_22677,N_22404,N_21149);
nand U22678 (N_22678,N_21016,N_21795);
nand U22679 (N_22679,N_21566,N_21643);
nor U22680 (N_22680,N_22292,N_22317);
and U22681 (N_22681,N_21059,N_22194);
and U22682 (N_22682,N_21316,N_21701);
xor U22683 (N_22683,N_21132,N_22275);
nor U22684 (N_22684,N_21532,N_21522);
nor U22685 (N_22685,N_22148,N_21058);
nand U22686 (N_22686,N_21929,N_22251);
nand U22687 (N_22687,N_22163,N_21513);
nor U22688 (N_22688,N_21351,N_21274);
nand U22689 (N_22689,N_21459,N_21230);
nor U22690 (N_22690,N_21562,N_21696);
nand U22691 (N_22691,N_21933,N_21462);
xnor U22692 (N_22692,N_22124,N_21473);
or U22693 (N_22693,N_21771,N_21982);
xnor U22694 (N_22694,N_22417,N_21505);
and U22695 (N_22695,N_21140,N_22227);
and U22696 (N_22696,N_22333,N_21621);
and U22697 (N_22697,N_22091,N_21337);
nor U22698 (N_22698,N_21636,N_21376);
nor U22699 (N_22699,N_21428,N_22248);
nor U22700 (N_22700,N_21483,N_21818);
and U22701 (N_22701,N_22448,N_22181);
and U22702 (N_22702,N_21339,N_21853);
and U22703 (N_22703,N_21755,N_21966);
nand U22704 (N_22704,N_21322,N_21287);
and U22705 (N_22705,N_21024,N_21396);
nor U22706 (N_22706,N_21427,N_21124);
and U22707 (N_22707,N_21259,N_22100);
nor U22708 (N_22708,N_21520,N_22063);
or U22709 (N_22709,N_21179,N_21759);
or U22710 (N_22710,N_21999,N_22199);
or U22711 (N_22711,N_21254,N_21006);
or U22712 (N_22712,N_21594,N_21245);
and U22713 (N_22713,N_21096,N_21728);
nor U22714 (N_22714,N_21804,N_22118);
or U22715 (N_22715,N_22309,N_21783);
nor U22716 (N_22716,N_22265,N_21945);
or U22717 (N_22717,N_22396,N_21260);
or U22718 (N_22718,N_21290,N_21297);
nor U22719 (N_22719,N_21774,N_21729);
xnor U22720 (N_22720,N_21000,N_22158);
and U22721 (N_22721,N_22287,N_21212);
and U22722 (N_22722,N_21269,N_22220);
and U22723 (N_22723,N_21619,N_22121);
nor U22724 (N_22724,N_22016,N_21499);
and U22725 (N_22725,N_22153,N_22355);
or U22726 (N_22726,N_22273,N_21182);
nor U22727 (N_22727,N_21913,N_21573);
or U22728 (N_22728,N_21705,N_21253);
xnor U22729 (N_22729,N_22187,N_21438);
and U22730 (N_22730,N_21504,N_21676);
nand U22731 (N_22731,N_21205,N_21185);
or U22732 (N_22732,N_21960,N_21622);
and U22733 (N_22733,N_22497,N_21592);
nand U22734 (N_22734,N_21764,N_21448);
and U22735 (N_22735,N_21324,N_22232);
nor U22736 (N_22736,N_21345,N_21588);
and U22737 (N_22737,N_21312,N_22380);
nand U22738 (N_22738,N_22098,N_21584);
nor U22739 (N_22739,N_21472,N_22328);
and U22740 (N_22740,N_21194,N_21196);
and U22741 (N_22741,N_22052,N_21480);
nor U22742 (N_22742,N_21994,N_21211);
nand U22743 (N_22743,N_21201,N_21927);
nand U22744 (N_22744,N_22444,N_21872);
or U22745 (N_22745,N_22498,N_21257);
nor U22746 (N_22746,N_21131,N_21418);
nand U22747 (N_22747,N_21022,N_21229);
or U22748 (N_22748,N_21481,N_21738);
nor U22749 (N_22749,N_21374,N_21436);
nor U22750 (N_22750,N_22261,N_21154);
nor U22751 (N_22751,N_21349,N_22061);
nor U22752 (N_22752,N_21369,N_22316);
nor U22753 (N_22753,N_21630,N_22432);
nand U22754 (N_22754,N_22472,N_22259);
or U22755 (N_22755,N_22285,N_22188);
and U22756 (N_22756,N_21542,N_22010);
and U22757 (N_22757,N_22192,N_22344);
xnor U22758 (N_22758,N_21089,N_22299);
and U22759 (N_22759,N_22075,N_22364);
nand U22760 (N_22760,N_21247,N_21153);
and U22761 (N_22761,N_22041,N_22422);
xnor U22762 (N_22762,N_21423,N_22236);
nor U22763 (N_22763,N_22073,N_21785);
nor U22764 (N_22764,N_22018,N_21318);
xnor U22765 (N_22765,N_22152,N_21251);
xor U22766 (N_22766,N_21711,N_22239);
nor U22767 (N_22767,N_22169,N_21099);
and U22768 (N_22768,N_21461,N_21150);
nand U22769 (N_22769,N_21845,N_21050);
and U22770 (N_22770,N_22104,N_21282);
nand U22771 (N_22771,N_22145,N_22186);
nand U22772 (N_22772,N_22288,N_21495);
and U22773 (N_22773,N_22055,N_21714);
and U22774 (N_22774,N_21227,N_21572);
and U22775 (N_22775,N_22147,N_22211);
nor U22776 (N_22776,N_21092,N_21686);
nand U22777 (N_22777,N_21426,N_21863);
or U22778 (N_22778,N_22172,N_21012);
nand U22779 (N_22779,N_21649,N_21552);
nand U22780 (N_22780,N_21395,N_21838);
and U22781 (N_22781,N_21431,N_22067);
or U22782 (N_22782,N_21756,N_21827);
nor U22783 (N_22783,N_22203,N_21019);
and U22784 (N_22784,N_22185,N_21453);
xnor U22785 (N_22785,N_21221,N_22156);
nand U22786 (N_22786,N_21571,N_21441);
nor U22787 (N_22787,N_21996,N_22406);
or U22788 (N_22788,N_22395,N_21487);
nand U22789 (N_22789,N_21717,N_22151);
nand U22790 (N_22790,N_22426,N_21527);
nor U22791 (N_22791,N_21557,N_21560);
xor U22792 (N_22792,N_21444,N_21346);
xnor U22793 (N_22793,N_21871,N_22209);
nand U22794 (N_22794,N_21550,N_22362);
and U22795 (N_22795,N_21105,N_21128);
nand U22796 (N_22796,N_21234,N_21026);
xor U22797 (N_22797,N_21490,N_21930);
and U22798 (N_22798,N_21861,N_21952);
xnor U22799 (N_22799,N_22271,N_21805);
or U22800 (N_22800,N_21432,N_21407);
nor U22801 (N_22801,N_21786,N_21722);
and U22802 (N_22802,N_21435,N_21943);
xnor U22803 (N_22803,N_21806,N_21001);
nor U22804 (N_22804,N_22234,N_21912);
and U22805 (N_22805,N_21799,N_21165);
xnor U22806 (N_22806,N_21471,N_22428);
nor U22807 (N_22807,N_21739,N_22004);
or U22808 (N_22808,N_22385,N_21813);
xor U22809 (N_22809,N_22009,N_21727);
or U22810 (N_22810,N_21359,N_21401);
or U22811 (N_22811,N_21569,N_21984);
nand U22812 (N_22812,N_22218,N_22381);
nor U22813 (N_22813,N_21545,N_21860);
and U22814 (N_22814,N_22352,N_21162);
and U22815 (N_22815,N_21158,N_22324);
nand U22816 (N_22816,N_21693,N_21655);
nand U22817 (N_22817,N_21136,N_21749);
or U22818 (N_22818,N_21546,N_21579);
and U22819 (N_22819,N_21521,N_22210);
nor U22820 (N_22820,N_21713,N_21313);
xor U22821 (N_22821,N_21458,N_22382);
xnor U22822 (N_22822,N_21508,N_22154);
nand U22823 (N_22823,N_21597,N_21398);
xnor U22824 (N_22824,N_22258,N_21973);
or U22825 (N_22825,N_21651,N_21575);
and U22826 (N_22826,N_21548,N_22379);
xor U22827 (N_22827,N_22032,N_22268);
nand U22828 (N_22828,N_22242,N_21862);
nor U22829 (N_22829,N_22008,N_21197);
nor U22830 (N_22830,N_21304,N_22413);
nor U22831 (N_22831,N_22435,N_22115);
and U22832 (N_22832,N_21256,N_21653);
or U22833 (N_22833,N_22254,N_22349);
xor U22834 (N_22834,N_21625,N_22245);
nand U22835 (N_22835,N_21334,N_21660);
xnor U22836 (N_22836,N_21650,N_21815);
or U22837 (N_22837,N_21393,N_21859);
or U22838 (N_22838,N_21326,N_21119);
nand U22839 (N_22839,N_22434,N_21869);
xnor U22840 (N_22840,N_22094,N_22481);
nand U22841 (N_22841,N_21905,N_21959);
or U22842 (N_22842,N_21637,N_21631);
nand U22843 (N_22843,N_21032,N_22391);
xor U22844 (N_22844,N_22375,N_21685);
or U22845 (N_22845,N_21474,N_21633);
and U22846 (N_22846,N_22183,N_21944);
and U22847 (N_22847,N_21955,N_21191);
and U22848 (N_22848,N_21767,N_21570);
xnor U22849 (N_22849,N_21268,N_22167);
nor U22850 (N_22850,N_21989,N_21343);
or U22851 (N_22851,N_22070,N_21134);
and U22852 (N_22852,N_21011,N_21248);
xnor U22853 (N_22853,N_21626,N_22184);
xnor U22854 (N_22854,N_21094,N_22042);
nor U22855 (N_22855,N_21358,N_21874);
nor U22856 (N_22856,N_21781,N_22137);
xnor U22857 (N_22857,N_22198,N_21325);
and U22858 (N_22858,N_21232,N_21126);
nand U22859 (N_22859,N_21214,N_21113);
xnor U22860 (N_22860,N_21486,N_21336);
nor U22861 (N_22861,N_21451,N_22224);
or U22862 (N_22862,N_22051,N_22013);
or U22863 (N_22863,N_21879,N_21081);
or U22864 (N_22864,N_22363,N_21956);
xnor U22865 (N_22865,N_21745,N_21004);
nand U22866 (N_22866,N_22197,N_22040);
or U22867 (N_22867,N_21183,N_21634);
nand U22868 (N_22868,N_21009,N_22469);
nand U22869 (N_22869,N_21666,N_22114);
or U22870 (N_22870,N_21616,N_21997);
or U22871 (N_22871,N_21577,N_21578);
nand U22872 (N_22872,N_21777,N_21084);
nand U22873 (N_22873,N_21931,N_22311);
xnor U22874 (N_22874,N_21980,N_21516);
or U22875 (N_22875,N_21840,N_21383);
xnor U22876 (N_22876,N_22420,N_22389);
or U22877 (N_22877,N_21352,N_21847);
xor U22878 (N_22878,N_22284,N_21920);
nor U22879 (N_22879,N_21125,N_22014);
nor U22880 (N_22880,N_22113,N_21112);
nand U22881 (N_22881,N_21823,N_21433);
nor U22882 (N_22882,N_21751,N_22141);
nand U22883 (N_22883,N_22222,N_22207);
and U22884 (N_22884,N_21591,N_21598);
and U22885 (N_22885,N_21100,N_22360);
and U22886 (N_22886,N_21576,N_21406);
nor U22887 (N_22887,N_21586,N_21954);
nand U22888 (N_22888,N_21223,N_22339);
nor U22889 (N_22889,N_22108,N_22095);
xor U22890 (N_22890,N_22367,N_22369);
nor U22891 (N_22891,N_21766,N_22059);
xor U22892 (N_22892,N_21262,N_21430);
xnor U22893 (N_22893,N_22054,N_21065);
or U22894 (N_22894,N_21294,N_21914);
nand U22895 (N_22895,N_21602,N_22048);
nand U22896 (N_22896,N_22002,N_21301);
nand U22897 (N_22897,N_21876,N_21122);
or U22898 (N_22898,N_22437,N_21014);
and U22899 (N_22899,N_21702,N_21901);
nor U22900 (N_22900,N_21733,N_21834);
or U22901 (N_22901,N_21348,N_21724);
and U22902 (N_22902,N_21335,N_21178);
nand U22903 (N_22903,N_22125,N_21850);
or U22904 (N_22904,N_21902,N_21895);
or U22905 (N_22905,N_21510,N_21890);
or U22906 (N_22906,N_21037,N_22446);
nor U22907 (N_22907,N_21184,N_21580);
nand U22908 (N_22908,N_22093,N_21662);
and U22909 (N_22909,N_22106,N_22160);
nand U22910 (N_22910,N_22025,N_21071);
and U22911 (N_22911,N_21768,N_22407);
or U22912 (N_22912,N_21856,N_21656);
nand U22913 (N_22913,N_22102,N_21226);
nand U22914 (N_22914,N_21793,N_21034);
or U22915 (N_22915,N_22495,N_21601);
nor U22916 (N_22916,N_22443,N_22269);
nand U22917 (N_22917,N_21043,N_22368);
or U22918 (N_22918,N_21951,N_21190);
or U22919 (N_22919,N_22429,N_22438);
and U22920 (N_22920,N_22022,N_21303);
and U22921 (N_22921,N_21500,N_21540);
and U22922 (N_22922,N_22202,N_21222);
or U22923 (N_22923,N_22351,N_21829);
or U22924 (N_22924,N_21344,N_21975);
nand U22925 (N_22925,N_21280,N_22084);
nand U22926 (N_22926,N_21403,N_22297);
nor U22927 (N_22927,N_22353,N_22318);
nand U22928 (N_22928,N_22112,N_21687);
nor U22929 (N_22929,N_21904,N_21225);
xnor U22930 (N_22930,N_21171,N_21391);
and U22931 (N_22931,N_22286,N_22412);
xnor U22932 (N_22932,N_21517,N_21790);
or U22933 (N_22933,N_21249,N_21614);
nand U22934 (N_22934,N_21776,N_21647);
xor U22935 (N_22935,N_21295,N_21246);
or U22936 (N_22936,N_21736,N_21028);
and U22937 (N_22937,N_22466,N_21948);
nor U22938 (N_22938,N_22492,N_21456);
or U22939 (N_22939,N_21258,N_21317);
nor U22940 (N_22940,N_21518,N_22023);
and U22941 (N_22941,N_21064,N_21720);
and U22942 (N_22942,N_22046,N_21817);
or U22943 (N_22943,N_21305,N_22482);
and U22944 (N_22944,N_21706,N_21308);
and U22945 (N_22945,N_21192,N_21589);
xnor U22946 (N_22946,N_22418,N_22090);
nand U22947 (N_22947,N_22235,N_22454);
and U22948 (N_22948,N_21507,N_22393);
or U22949 (N_22949,N_21526,N_21574);
nand U22950 (N_22950,N_22131,N_22057);
xnor U22951 (N_22951,N_22173,N_21091);
or U22952 (N_22952,N_22136,N_22415);
nand U22953 (N_22953,N_21867,N_21130);
xor U22954 (N_22954,N_22244,N_21814);
nor U22955 (N_22955,N_21266,N_21265);
and U22956 (N_22956,N_22452,N_21559);
nand U22957 (N_22957,N_21169,N_21939);
or U22958 (N_22958,N_21556,N_22290);
nand U22959 (N_22959,N_21492,N_21969);
nand U22960 (N_22960,N_22485,N_22200);
nand U22961 (N_22961,N_21379,N_22499);
nand U22962 (N_22962,N_21075,N_21613);
nor U22963 (N_22963,N_22431,N_21189);
nor U22964 (N_22964,N_21549,N_21181);
xnor U22965 (N_22965,N_22301,N_22175);
or U22966 (N_22966,N_21998,N_22086);
nor U22967 (N_22967,N_21665,N_22439);
nor U22968 (N_22968,N_21893,N_21108);
nor U22969 (N_22969,N_21429,N_21744);
xor U22970 (N_22970,N_21934,N_22277);
and U22971 (N_22971,N_21864,N_22471);
nand U22972 (N_22972,N_21425,N_21285);
nand U22973 (N_22973,N_22445,N_22116);
xor U22974 (N_22974,N_21600,N_22246);
and U22975 (N_22975,N_21388,N_21923);
or U22976 (N_22976,N_22336,N_21801);
nand U22977 (N_22977,N_21264,N_21110);
xor U22978 (N_22978,N_21467,N_21536);
nor U22979 (N_22979,N_22003,N_21123);
xor U22980 (N_22980,N_22082,N_21278);
nor U22981 (N_22981,N_22483,N_22044);
or U22982 (N_22982,N_21068,N_21553);
and U22983 (N_22983,N_22455,N_22341);
or U22984 (N_22984,N_21005,N_22026);
xnor U22985 (N_22985,N_21652,N_21644);
nand U22986 (N_22986,N_22189,N_21103);
and U22987 (N_22987,N_21991,N_21402);
xor U22988 (N_22988,N_22414,N_21608);
or U22989 (N_22989,N_21972,N_21615);
nand U22990 (N_22990,N_21928,N_21347);
nor U22991 (N_22991,N_21921,N_21691);
nand U22992 (N_22992,N_21638,N_21378);
xnor U22993 (N_22993,N_21371,N_21238);
or U22994 (N_22994,N_21442,N_21884);
or U22995 (N_22995,N_21618,N_21629);
and U22996 (N_22996,N_22473,N_21978);
nand U22997 (N_22997,N_21076,N_21535);
nand U22998 (N_22998,N_21870,N_21241);
xor U22999 (N_22999,N_21778,N_22101);
and U23000 (N_23000,N_22304,N_21299);
and U23001 (N_23001,N_21281,N_21404);
xnor U23002 (N_23002,N_21228,N_21413);
nand U23003 (N_23003,N_21353,N_21740);
nor U23004 (N_23004,N_21120,N_22020);
nor U23005 (N_23005,N_21494,N_21362);
or U23006 (N_23006,N_21692,N_21469);
nor U23007 (N_23007,N_21648,N_21624);
xnor U23008 (N_23008,N_21798,N_21350);
nor U23009 (N_23009,N_22083,N_22256);
nand U23010 (N_23010,N_21640,N_21544);
nand U23011 (N_23011,N_21970,N_21193);
nor U23012 (N_23012,N_21770,N_21315);
and U23013 (N_23013,N_21493,N_21509);
nand U23014 (N_23014,N_21235,N_21087);
or U23015 (N_23015,N_21200,N_21609);
and U23016 (N_23016,N_21479,N_21796);
nor U23017 (N_23017,N_21911,N_22038);
and U23018 (N_23018,N_21320,N_22088);
or U23019 (N_23019,N_21377,N_22331);
or U23020 (N_23020,N_21673,N_22398);
or U23021 (N_23021,N_22441,N_21993);
nor U23022 (N_23022,N_21563,N_22423);
xnor U23023 (N_23023,N_21118,N_21782);
nand U23024 (N_23024,N_21963,N_22087);
or U23025 (N_23025,N_21415,N_21139);
nor U23026 (N_23026,N_21658,N_21498);
nor U23027 (N_23027,N_21822,N_22350);
nand U23028 (N_23028,N_21323,N_21852);
nor U23029 (N_23029,N_21791,N_22278);
nand U23030 (N_23030,N_21667,N_21679);
or U23031 (N_23031,N_22449,N_21908);
nor U23032 (N_23032,N_21017,N_21981);
and U23033 (N_23033,N_21063,N_21400);
xnor U23034 (N_23034,N_22390,N_22128);
nand U23035 (N_23035,N_21289,N_21800);
xor U23036 (N_23036,N_21919,N_21976);
nand U23037 (N_23037,N_21175,N_21204);
or U23038 (N_23038,N_21677,N_22130);
xor U23039 (N_23039,N_22109,N_21419);
nor U23040 (N_23040,N_22017,N_22295);
and U23041 (N_23041,N_21891,N_21506);
nand U23042 (N_23042,N_22424,N_22212);
or U23043 (N_23043,N_21062,N_21055);
and U23044 (N_23044,N_21082,N_22266);
or U23045 (N_23045,N_21669,N_22190);
nor U23046 (N_23046,N_22117,N_22459);
or U23047 (N_23047,N_21690,N_22281);
xnor U23048 (N_23048,N_21074,N_21773);
or U23049 (N_23049,N_21539,N_22253);
nor U23050 (N_23050,N_21909,N_22241);
and U23051 (N_23051,N_22024,N_22347);
xor U23052 (N_23052,N_22308,N_21047);
nor U23053 (N_23053,N_22066,N_21437);
xor U23054 (N_23054,N_22496,N_22386);
xor U23055 (N_23055,N_21681,N_21167);
nor U23056 (N_23056,N_22411,N_21512);
or U23057 (N_23057,N_22047,N_21455);
and U23058 (N_23058,N_22335,N_21639);
nand U23059 (N_23059,N_21514,N_21166);
nor U23060 (N_23060,N_21078,N_21938);
nor U23061 (N_23061,N_22365,N_21979);
or U23062 (N_23062,N_21583,N_22276);
nor U23063 (N_23063,N_21695,N_22247);
or U23064 (N_23064,N_22031,N_21596);
and U23065 (N_23065,N_21440,N_21661);
xnor U23066 (N_23066,N_21581,N_21410);
nand U23067 (N_23067,N_21233,N_21515);
and U23068 (N_23068,N_21477,N_21585);
nand U23069 (N_23069,N_21199,N_22260);
and U23070 (N_23070,N_22089,N_21645);
or U23071 (N_23071,N_21907,N_22399);
nand U23072 (N_23072,N_22272,N_21408);
xnor U23073 (N_23073,N_22314,N_22394);
xor U23074 (N_23074,N_21328,N_22325);
xnor U23075 (N_23075,N_21476,N_21168);
or U23076 (N_23076,N_22405,N_22456);
nor U23077 (N_23077,N_22097,N_21077);
xor U23078 (N_23078,N_21443,N_21828);
or U23079 (N_23079,N_21088,N_22064);
nor U23080 (N_23080,N_21342,N_22133);
nor U23081 (N_23081,N_21023,N_21070);
nand U23082 (N_23082,N_21623,N_22373);
and U23083 (N_23083,N_21160,N_21501);
nand U23084 (N_23084,N_21837,N_21292);
nor U23085 (N_23085,N_21215,N_21036);
xnor U23086 (N_23086,N_22257,N_21710);
xnor U23087 (N_23087,N_22077,N_21762);
or U23088 (N_23088,N_21392,N_21628);
nor U23089 (N_23089,N_21338,N_22157);
xor U23090 (N_23090,N_22217,N_22326);
and U23091 (N_23091,N_22053,N_21370);
nand U23092 (N_23092,N_22416,N_21332);
nand U23093 (N_23093,N_21029,N_21203);
nand U23094 (N_23094,N_21985,N_21611);
or U23095 (N_23095,N_21031,N_21003);
xor U23096 (N_23096,N_21057,N_21886);
and U23097 (N_23097,N_21888,N_22065);
and U23098 (N_23098,N_22453,N_21809);
or U23099 (N_23099,N_22176,N_21757);
nand U23100 (N_23100,N_21279,N_21298);
xnor U23101 (N_23101,N_21746,N_21537);
and U23102 (N_23102,N_21060,N_21240);
nor U23103 (N_23103,N_21025,N_21698);
xnor U23104 (N_23104,N_21632,N_21754);
nor U23105 (N_23105,N_21743,N_22488);
xor U23106 (N_23106,N_21697,N_22238);
and U23107 (N_23107,N_22049,N_22489);
and U23108 (N_23108,N_22119,N_21842);
or U23109 (N_23109,N_22410,N_22201);
or U23110 (N_23110,N_21719,N_21263);
nor U23111 (N_23111,N_21607,N_21846);
xor U23112 (N_23112,N_21555,N_22228);
and U23113 (N_23113,N_21250,N_22467);
nor U23114 (N_23114,N_21083,N_21286);
or U23115 (N_23115,N_21551,N_22033);
xnor U23116 (N_23116,N_21341,N_22433);
nor U23117 (N_23117,N_21962,N_22140);
and U23118 (N_23118,N_21127,N_22312);
nand U23119 (N_23119,N_21340,N_21896);
nor U23120 (N_23120,N_22223,N_21373);
nand U23121 (N_23121,N_22215,N_21465);
nor U23122 (N_23122,N_21689,N_21599);
or U23123 (N_23123,N_21177,N_21821);
xnor U23124 (N_23124,N_21390,N_21797);
and U23125 (N_23125,N_21758,N_22155);
nand U23126 (N_23126,N_21567,N_21231);
and U23127 (N_23127,N_22397,N_21885);
or U23128 (N_23128,N_21947,N_21538);
xnor U23129 (N_23129,N_21610,N_21765);
nor U23130 (N_23130,N_22296,N_21620);
nand U23131 (N_23131,N_21311,N_22491);
or U23132 (N_23132,N_22457,N_21502);
or U23133 (N_23133,N_21883,N_21497);
and U23134 (N_23134,N_21950,N_21529);
or U23135 (N_23135,N_22216,N_21554);
and U23136 (N_23136,N_22191,N_21779);
nor U23137 (N_23137,N_21663,N_21104);
or U23138 (N_23138,N_21491,N_21519);
or U23139 (N_23139,N_22226,N_21186);
nor U23140 (N_23140,N_21543,N_22193);
xnor U23141 (N_23141,N_22069,N_21825);
and U23142 (N_23142,N_21617,N_22303);
nor U23143 (N_23143,N_22327,N_22357);
nor U23144 (N_23144,N_21716,N_21683);
and U23145 (N_23145,N_21731,N_21820);
or U23146 (N_23146,N_22262,N_21812);
xnor U23147 (N_23147,N_22294,N_21769);
or U23148 (N_23148,N_21830,N_22034);
or U23149 (N_23149,N_22387,N_21217);
nand U23150 (N_23150,N_22214,N_21899);
nor U23151 (N_23151,N_22490,N_22092);
or U23152 (N_23152,N_21357,N_21558);
nor U23153 (N_23153,N_22409,N_21180);
and U23154 (N_23154,N_21582,N_21735);
xor U23155 (N_23155,N_22027,N_21450);
or U23156 (N_23156,N_21293,N_21752);
or U23157 (N_23157,N_21750,N_21210);
and U23158 (N_23158,N_22159,N_21272);
or U23159 (N_23159,N_21384,N_22050);
nand U23160 (N_23160,N_21449,N_22074);
and U23161 (N_23161,N_22170,N_21484);
nor U23162 (N_23162,N_21531,N_22465);
nand U23163 (N_23163,N_21157,N_21855);
and U23164 (N_23164,N_22464,N_21463);
nor U23165 (N_23165,N_22319,N_21977);
or U23166 (N_23166,N_21020,N_21121);
nand U23167 (N_23167,N_22233,N_21173);
and U23168 (N_23168,N_22447,N_22302);
and U23169 (N_23169,N_21460,N_21093);
or U23170 (N_23170,N_22479,N_21364);
or U23171 (N_23171,N_22345,N_22463);
nand U23172 (N_23172,N_21021,N_22388);
and U23173 (N_23173,N_22306,N_21035);
and U23174 (N_23174,N_21244,N_21220);
nand U23175 (N_23175,N_22177,N_22470);
xnor U23176 (N_23176,N_22249,N_22401);
and U23177 (N_23177,N_21937,N_21678);
xnor U23178 (N_23178,N_22240,N_21156);
xor U23179 (N_23179,N_22494,N_21273);
and U23180 (N_23180,N_21868,N_22400);
nor U23181 (N_23181,N_21675,N_22012);
xnor U23182 (N_23182,N_22099,N_21906);
xor U23183 (N_23183,N_21188,N_21898);
nand U23184 (N_23184,N_22263,N_22383);
nor U23185 (N_23185,N_21270,N_21835);
and U23186 (N_23186,N_21085,N_21069);
xnor U23187 (N_23187,N_21355,N_22043);
nor U23188 (N_23188,N_22366,N_21447);
xnor U23189 (N_23189,N_21375,N_21726);
nand U23190 (N_23190,N_21986,N_21366);
or U23191 (N_23191,N_22166,N_21763);
nand U23192 (N_23192,N_21198,N_21603);
nand U23193 (N_23193,N_21207,N_22123);
or U23194 (N_23194,N_22378,N_22332);
and U23195 (N_23195,N_22146,N_22310);
xnor U23196 (N_23196,N_21424,N_21833);
xnor U23197 (N_23197,N_21030,N_22144);
or U23198 (N_23198,N_22162,N_21288);
nor U23199 (N_23199,N_21488,N_22045);
or U23200 (N_23200,N_21412,N_21385);
or U23201 (N_23201,N_21386,N_22298);
nor U23202 (N_23202,N_21457,N_22305);
nand U23203 (N_23203,N_21174,N_22149);
or U23204 (N_23204,N_21857,N_21946);
nor U23205 (N_23205,N_21682,N_21780);
and U23206 (N_23206,N_21409,N_22030);
nor U23207 (N_23207,N_21940,N_21760);
and U23208 (N_23208,N_21811,N_22356);
nand U23209 (N_23209,N_22313,N_22231);
or U23210 (N_23210,N_21051,N_21086);
nor U23211 (N_23211,N_22206,N_21114);
nor U23212 (N_23212,N_22036,N_22230);
xnor U23213 (N_23213,N_22142,N_21018);
xnor U23214 (N_23214,N_21858,N_21417);
xnor U23215 (N_23215,N_21680,N_21732);
xor U23216 (N_23216,N_21849,N_22338);
nand U23217 (N_23217,N_21612,N_21098);
xnor U23218 (N_23218,N_21236,N_21237);
xor U23219 (N_23219,N_21587,N_22282);
and U23220 (N_23220,N_21381,N_21389);
and U23221 (N_23221,N_21916,N_22058);
nor U23222 (N_23222,N_21748,N_21593);
or U23223 (N_23223,N_22204,N_22139);
and U23224 (N_23224,N_22127,N_21145);
nand U23225 (N_23225,N_22374,N_22129);
nor U23226 (N_23226,N_21851,N_21924);
and U23227 (N_23227,N_22219,N_21161);
nor U23228 (N_23228,N_22468,N_22019);
or U23229 (N_23229,N_22402,N_21421);
or U23230 (N_23230,N_22161,N_22427);
nor U23231 (N_23231,N_21106,N_21892);
nor U23232 (N_23232,N_21464,N_21010);
nand U23233 (N_23233,N_22000,N_21541);
nor U23234 (N_23234,N_21882,N_22320);
nand U23235 (N_23235,N_22307,N_21095);
or U23236 (N_23236,N_22068,N_21646);
nand U23237 (N_23237,N_22403,N_22359);
or U23238 (N_23238,N_21310,N_21372);
xor U23239 (N_23239,N_21382,N_22267);
or U23240 (N_23240,N_21072,N_21142);
nor U23241 (N_23241,N_22056,N_21794);
nor U23242 (N_23242,N_22174,N_21657);
or U23243 (N_23243,N_21331,N_22270);
and U23244 (N_23244,N_21707,N_21974);
or U23245 (N_23245,N_21284,N_22477);
nor U23246 (N_23246,N_21958,N_21747);
or U23247 (N_23247,N_21468,N_21918);
and U23248 (N_23248,N_21503,N_21013);
xnor U23249 (N_23249,N_21296,N_21470);
nor U23250 (N_23250,N_21570,N_21356);
or U23251 (N_23251,N_21601,N_22238);
xnor U23252 (N_23252,N_22400,N_21330);
or U23253 (N_23253,N_21373,N_22264);
or U23254 (N_23254,N_21355,N_22088);
nor U23255 (N_23255,N_22006,N_21218);
xnor U23256 (N_23256,N_21508,N_22291);
or U23257 (N_23257,N_21767,N_21558);
or U23258 (N_23258,N_21611,N_21359);
xor U23259 (N_23259,N_21348,N_21980);
nor U23260 (N_23260,N_21225,N_21499);
xor U23261 (N_23261,N_22070,N_22376);
nand U23262 (N_23262,N_22481,N_21459);
nand U23263 (N_23263,N_21151,N_22210);
and U23264 (N_23264,N_21661,N_22188);
or U23265 (N_23265,N_22134,N_21314);
nand U23266 (N_23266,N_21563,N_21790);
nor U23267 (N_23267,N_22169,N_21322);
xor U23268 (N_23268,N_21025,N_21838);
xnor U23269 (N_23269,N_21690,N_22312);
nor U23270 (N_23270,N_21784,N_21545);
xor U23271 (N_23271,N_21769,N_21199);
and U23272 (N_23272,N_21435,N_22495);
nand U23273 (N_23273,N_21975,N_21222);
nor U23274 (N_23274,N_21208,N_21405);
nand U23275 (N_23275,N_22340,N_22429);
and U23276 (N_23276,N_22001,N_22309);
or U23277 (N_23277,N_22285,N_21082);
nand U23278 (N_23278,N_21788,N_21500);
nor U23279 (N_23279,N_21425,N_22421);
and U23280 (N_23280,N_22243,N_21011);
nor U23281 (N_23281,N_21335,N_21479);
nand U23282 (N_23282,N_21399,N_22052);
and U23283 (N_23283,N_21207,N_21859);
xnor U23284 (N_23284,N_21642,N_21036);
nor U23285 (N_23285,N_22254,N_21892);
or U23286 (N_23286,N_21708,N_22138);
nor U23287 (N_23287,N_21885,N_22074);
or U23288 (N_23288,N_22064,N_22110);
xnor U23289 (N_23289,N_22063,N_21151);
and U23290 (N_23290,N_22265,N_22337);
or U23291 (N_23291,N_21390,N_21689);
or U23292 (N_23292,N_21321,N_21481);
or U23293 (N_23293,N_21526,N_21140);
and U23294 (N_23294,N_21203,N_22493);
or U23295 (N_23295,N_22355,N_21136);
xor U23296 (N_23296,N_21114,N_21766);
or U23297 (N_23297,N_21556,N_22010);
xor U23298 (N_23298,N_21757,N_22165);
and U23299 (N_23299,N_21200,N_21628);
and U23300 (N_23300,N_21580,N_21346);
and U23301 (N_23301,N_22005,N_21589);
nor U23302 (N_23302,N_21107,N_21361);
and U23303 (N_23303,N_21883,N_22123);
nand U23304 (N_23304,N_21910,N_21105);
xor U23305 (N_23305,N_22161,N_22146);
or U23306 (N_23306,N_21726,N_22321);
nor U23307 (N_23307,N_21889,N_21303);
nand U23308 (N_23308,N_22173,N_21253);
or U23309 (N_23309,N_21462,N_21510);
nand U23310 (N_23310,N_21525,N_21594);
xor U23311 (N_23311,N_21649,N_21975);
or U23312 (N_23312,N_21463,N_21317);
nand U23313 (N_23313,N_21734,N_21637);
xnor U23314 (N_23314,N_21828,N_21254);
or U23315 (N_23315,N_21844,N_21512);
xor U23316 (N_23316,N_21788,N_21510);
nand U23317 (N_23317,N_21334,N_21170);
nand U23318 (N_23318,N_22175,N_22163);
nor U23319 (N_23319,N_21157,N_22448);
xor U23320 (N_23320,N_21202,N_22320);
xnor U23321 (N_23321,N_21456,N_22140);
xor U23322 (N_23322,N_21555,N_21136);
and U23323 (N_23323,N_21145,N_21367);
xnor U23324 (N_23324,N_21162,N_21000);
xnor U23325 (N_23325,N_22080,N_21848);
nand U23326 (N_23326,N_21366,N_22110);
nand U23327 (N_23327,N_21676,N_21528);
and U23328 (N_23328,N_21444,N_21482);
nor U23329 (N_23329,N_21192,N_21884);
nor U23330 (N_23330,N_22210,N_21183);
nand U23331 (N_23331,N_21457,N_22094);
or U23332 (N_23332,N_21578,N_21605);
nand U23333 (N_23333,N_21153,N_21985);
and U23334 (N_23334,N_22161,N_21594);
or U23335 (N_23335,N_22120,N_21471);
or U23336 (N_23336,N_21874,N_21586);
nand U23337 (N_23337,N_21312,N_22142);
nand U23338 (N_23338,N_22125,N_22247);
xnor U23339 (N_23339,N_21512,N_21278);
or U23340 (N_23340,N_21021,N_21520);
nor U23341 (N_23341,N_22278,N_22019);
xnor U23342 (N_23342,N_21298,N_22381);
nor U23343 (N_23343,N_21129,N_21786);
and U23344 (N_23344,N_22050,N_21789);
and U23345 (N_23345,N_22378,N_22429);
nor U23346 (N_23346,N_22381,N_21224);
or U23347 (N_23347,N_21641,N_21154);
and U23348 (N_23348,N_22427,N_22138);
nor U23349 (N_23349,N_21673,N_22015);
nand U23350 (N_23350,N_22442,N_21289);
or U23351 (N_23351,N_21094,N_21434);
nor U23352 (N_23352,N_22440,N_22360);
nor U23353 (N_23353,N_21690,N_21927);
nand U23354 (N_23354,N_21989,N_22422);
xor U23355 (N_23355,N_21950,N_22156);
and U23356 (N_23356,N_21723,N_21428);
or U23357 (N_23357,N_21509,N_21540);
nor U23358 (N_23358,N_21804,N_22053);
nor U23359 (N_23359,N_22366,N_22435);
nor U23360 (N_23360,N_22127,N_21503);
nand U23361 (N_23361,N_22024,N_21962);
nor U23362 (N_23362,N_21683,N_21221);
nor U23363 (N_23363,N_22143,N_22153);
nand U23364 (N_23364,N_21664,N_21204);
xor U23365 (N_23365,N_21733,N_22413);
nand U23366 (N_23366,N_21617,N_21286);
nand U23367 (N_23367,N_22139,N_21130);
nand U23368 (N_23368,N_21336,N_22350);
nand U23369 (N_23369,N_21332,N_22449);
nor U23370 (N_23370,N_21189,N_21433);
nand U23371 (N_23371,N_21304,N_22029);
xor U23372 (N_23372,N_22381,N_21504);
and U23373 (N_23373,N_21857,N_21088);
or U23374 (N_23374,N_22340,N_21033);
xnor U23375 (N_23375,N_22444,N_21510);
xor U23376 (N_23376,N_21706,N_22440);
nand U23377 (N_23377,N_22278,N_21764);
nand U23378 (N_23378,N_22334,N_21874);
nand U23379 (N_23379,N_22283,N_21624);
nor U23380 (N_23380,N_21532,N_21221);
or U23381 (N_23381,N_21260,N_21057);
xnor U23382 (N_23382,N_21872,N_21296);
xnor U23383 (N_23383,N_22406,N_21164);
nor U23384 (N_23384,N_21531,N_21387);
and U23385 (N_23385,N_21700,N_21873);
xnor U23386 (N_23386,N_21315,N_21577);
nand U23387 (N_23387,N_21935,N_22081);
and U23388 (N_23388,N_21803,N_22443);
and U23389 (N_23389,N_22167,N_22019);
and U23390 (N_23390,N_22026,N_21197);
xnor U23391 (N_23391,N_21179,N_22485);
nor U23392 (N_23392,N_22262,N_22488);
and U23393 (N_23393,N_21278,N_22479);
xor U23394 (N_23394,N_21109,N_21226);
and U23395 (N_23395,N_22332,N_21602);
xnor U23396 (N_23396,N_21721,N_21090);
nor U23397 (N_23397,N_22276,N_22492);
nor U23398 (N_23398,N_22477,N_22471);
and U23399 (N_23399,N_21560,N_21893);
xnor U23400 (N_23400,N_21976,N_22028);
nand U23401 (N_23401,N_21575,N_21813);
xor U23402 (N_23402,N_21148,N_21558);
nand U23403 (N_23403,N_21609,N_21446);
xnor U23404 (N_23404,N_21855,N_21502);
and U23405 (N_23405,N_22111,N_21643);
nand U23406 (N_23406,N_21407,N_21306);
nand U23407 (N_23407,N_21081,N_21846);
nor U23408 (N_23408,N_22341,N_21274);
and U23409 (N_23409,N_21360,N_21008);
nor U23410 (N_23410,N_21291,N_21946);
or U23411 (N_23411,N_21180,N_22426);
nand U23412 (N_23412,N_21884,N_21003);
and U23413 (N_23413,N_21261,N_21344);
nand U23414 (N_23414,N_22440,N_21937);
xor U23415 (N_23415,N_21408,N_21641);
or U23416 (N_23416,N_22103,N_21195);
or U23417 (N_23417,N_21003,N_21944);
nor U23418 (N_23418,N_21313,N_21863);
or U23419 (N_23419,N_21180,N_21243);
nor U23420 (N_23420,N_21996,N_21018);
xor U23421 (N_23421,N_21270,N_21913);
nand U23422 (N_23422,N_22135,N_21435);
xnor U23423 (N_23423,N_21526,N_21325);
and U23424 (N_23424,N_22052,N_21404);
or U23425 (N_23425,N_22221,N_21854);
nand U23426 (N_23426,N_21568,N_21729);
nand U23427 (N_23427,N_21060,N_22382);
nand U23428 (N_23428,N_21309,N_22470);
or U23429 (N_23429,N_22174,N_22177);
and U23430 (N_23430,N_22454,N_21683);
nand U23431 (N_23431,N_22362,N_21392);
nand U23432 (N_23432,N_22498,N_21961);
and U23433 (N_23433,N_21698,N_21902);
nor U23434 (N_23434,N_21073,N_21584);
xor U23435 (N_23435,N_21020,N_22475);
nor U23436 (N_23436,N_21571,N_21797);
nor U23437 (N_23437,N_21455,N_21772);
and U23438 (N_23438,N_21669,N_21838);
nor U23439 (N_23439,N_21179,N_22065);
and U23440 (N_23440,N_21137,N_21815);
nor U23441 (N_23441,N_22036,N_21245);
xnor U23442 (N_23442,N_21914,N_21966);
and U23443 (N_23443,N_21050,N_21741);
or U23444 (N_23444,N_21589,N_22470);
xnor U23445 (N_23445,N_22110,N_21664);
nand U23446 (N_23446,N_22456,N_22301);
nand U23447 (N_23447,N_21586,N_21768);
or U23448 (N_23448,N_21369,N_21631);
nand U23449 (N_23449,N_21035,N_21043);
and U23450 (N_23450,N_21280,N_22119);
nand U23451 (N_23451,N_22047,N_22001);
xor U23452 (N_23452,N_21351,N_22376);
xor U23453 (N_23453,N_21922,N_21041);
nor U23454 (N_23454,N_21677,N_22305);
nand U23455 (N_23455,N_22385,N_22073);
xnor U23456 (N_23456,N_21840,N_21246);
nand U23457 (N_23457,N_22330,N_21139);
nand U23458 (N_23458,N_21253,N_21468);
or U23459 (N_23459,N_22160,N_22274);
and U23460 (N_23460,N_21112,N_22197);
or U23461 (N_23461,N_22380,N_22337);
and U23462 (N_23462,N_21645,N_22252);
or U23463 (N_23463,N_21493,N_22363);
xor U23464 (N_23464,N_21518,N_22244);
or U23465 (N_23465,N_22430,N_21280);
and U23466 (N_23466,N_21078,N_22316);
xor U23467 (N_23467,N_21619,N_21691);
nor U23468 (N_23468,N_21844,N_21252);
nand U23469 (N_23469,N_21921,N_21755);
or U23470 (N_23470,N_21467,N_21385);
nand U23471 (N_23471,N_21194,N_22446);
nand U23472 (N_23472,N_21528,N_21405);
xnor U23473 (N_23473,N_21892,N_22266);
or U23474 (N_23474,N_22260,N_21853);
and U23475 (N_23475,N_22003,N_22439);
and U23476 (N_23476,N_21149,N_21408);
nand U23477 (N_23477,N_21163,N_21316);
nand U23478 (N_23478,N_21090,N_22068);
xnor U23479 (N_23479,N_21767,N_21394);
and U23480 (N_23480,N_22284,N_22187);
or U23481 (N_23481,N_21932,N_21591);
nand U23482 (N_23482,N_22356,N_21315);
xnor U23483 (N_23483,N_22112,N_21040);
xor U23484 (N_23484,N_21153,N_21478);
or U23485 (N_23485,N_21427,N_21535);
and U23486 (N_23486,N_21690,N_21182);
or U23487 (N_23487,N_21893,N_22117);
xnor U23488 (N_23488,N_22054,N_22113);
and U23489 (N_23489,N_21813,N_21321);
nand U23490 (N_23490,N_21526,N_22309);
or U23491 (N_23491,N_22201,N_22270);
nor U23492 (N_23492,N_21773,N_21603);
or U23493 (N_23493,N_21836,N_22293);
and U23494 (N_23494,N_21337,N_21816);
nor U23495 (N_23495,N_21655,N_21423);
or U23496 (N_23496,N_21224,N_22010);
xnor U23497 (N_23497,N_21277,N_21571);
nand U23498 (N_23498,N_22179,N_22426);
nand U23499 (N_23499,N_21495,N_21661);
xnor U23500 (N_23500,N_22214,N_22420);
nand U23501 (N_23501,N_21980,N_21815);
and U23502 (N_23502,N_21442,N_22285);
or U23503 (N_23503,N_21841,N_22327);
nand U23504 (N_23504,N_21516,N_21672);
and U23505 (N_23505,N_21161,N_22446);
or U23506 (N_23506,N_21003,N_21568);
or U23507 (N_23507,N_21249,N_21673);
and U23508 (N_23508,N_22227,N_22345);
xnor U23509 (N_23509,N_21387,N_21702);
nand U23510 (N_23510,N_21597,N_21074);
nor U23511 (N_23511,N_21505,N_22306);
nand U23512 (N_23512,N_22339,N_22084);
nor U23513 (N_23513,N_21404,N_22093);
xnor U23514 (N_23514,N_21684,N_21301);
and U23515 (N_23515,N_22285,N_21092);
nor U23516 (N_23516,N_22070,N_21641);
xnor U23517 (N_23517,N_21134,N_21227);
and U23518 (N_23518,N_21510,N_22487);
nand U23519 (N_23519,N_21636,N_21891);
xnor U23520 (N_23520,N_22136,N_21071);
xnor U23521 (N_23521,N_22123,N_22284);
or U23522 (N_23522,N_22480,N_21538);
and U23523 (N_23523,N_21779,N_21975);
or U23524 (N_23524,N_22010,N_21832);
nand U23525 (N_23525,N_21462,N_21467);
nor U23526 (N_23526,N_22086,N_21702);
nand U23527 (N_23527,N_21990,N_22179);
or U23528 (N_23528,N_21857,N_21231);
and U23529 (N_23529,N_22079,N_21385);
xnor U23530 (N_23530,N_21963,N_22470);
nand U23531 (N_23531,N_22413,N_21032);
nand U23532 (N_23532,N_22018,N_22132);
nor U23533 (N_23533,N_22036,N_22138);
and U23534 (N_23534,N_21633,N_21851);
and U23535 (N_23535,N_22189,N_21007);
or U23536 (N_23536,N_22078,N_21116);
and U23537 (N_23537,N_22073,N_21628);
or U23538 (N_23538,N_22290,N_21350);
xor U23539 (N_23539,N_21937,N_21656);
and U23540 (N_23540,N_21629,N_21572);
or U23541 (N_23541,N_21874,N_22205);
xor U23542 (N_23542,N_21426,N_21833);
nand U23543 (N_23543,N_21198,N_21696);
nand U23544 (N_23544,N_21178,N_21272);
nor U23545 (N_23545,N_21669,N_21167);
or U23546 (N_23546,N_22176,N_21426);
xnor U23547 (N_23547,N_22169,N_21328);
and U23548 (N_23548,N_21212,N_22281);
or U23549 (N_23549,N_22325,N_22343);
nor U23550 (N_23550,N_21357,N_21127);
xor U23551 (N_23551,N_21101,N_22256);
nor U23552 (N_23552,N_22391,N_22407);
xor U23553 (N_23553,N_21303,N_21766);
or U23554 (N_23554,N_21970,N_21377);
and U23555 (N_23555,N_21655,N_22351);
or U23556 (N_23556,N_21151,N_21297);
nor U23557 (N_23557,N_22119,N_22051);
nand U23558 (N_23558,N_22431,N_21264);
nor U23559 (N_23559,N_21178,N_22119);
and U23560 (N_23560,N_21031,N_21380);
xnor U23561 (N_23561,N_22089,N_21714);
nand U23562 (N_23562,N_22026,N_22489);
nand U23563 (N_23563,N_21812,N_22313);
and U23564 (N_23564,N_21994,N_22322);
nand U23565 (N_23565,N_21549,N_22163);
xnor U23566 (N_23566,N_21440,N_21553);
or U23567 (N_23567,N_21751,N_22446);
and U23568 (N_23568,N_21703,N_21875);
nor U23569 (N_23569,N_22486,N_22045);
and U23570 (N_23570,N_22325,N_22441);
and U23571 (N_23571,N_21162,N_21338);
and U23572 (N_23572,N_22483,N_21480);
nor U23573 (N_23573,N_21938,N_21566);
nor U23574 (N_23574,N_21620,N_21801);
and U23575 (N_23575,N_22387,N_21806);
or U23576 (N_23576,N_21875,N_22381);
nand U23577 (N_23577,N_22144,N_22079);
xor U23578 (N_23578,N_21121,N_22433);
nor U23579 (N_23579,N_21896,N_21125);
nor U23580 (N_23580,N_21259,N_21763);
or U23581 (N_23581,N_21218,N_21534);
nand U23582 (N_23582,N_22433,N_22207);
xnor U23583 (N_23583,N_21486,N_21682);
nor U23584 (N_23584,N_21596,N_21156);
nor U23585 (N_23585,N_22243,N_21354);
or U23586 (N_23586,N_22474,N_21428);
xor U23587 (N_23587,N_22403,N_21610);
nor U23588 (N_23588,N_21187,N_22225);
xnor U23589 (N_23589,N_21569,N_21458);
or U23590 (N_23590,N_22310,N_22004);
or U23591 (N_23591,N_21050,N_22026);
nor U23592 (N_23592,N_21031,N_21022);
or U23593 (N_23593,N_22074,N_21104);
or U23594 (N_23594,N_21192,N_22071);
nand U23595 (N_23595,N_22179,N_21913);
nand U23596 (N_23596,N_22325,N_21496);
xnor U23597 (N_23597,N_21754,N_21062);
or U23598 (N_23598,N_21387,N_21438);
nor U23599 (N_23599,N_22176,N_21974);
nor U23600 (N_23600,N_21225,N_21632);
nor U23601 (N_23601,N_22317,N_21696);
or U23602 (N_23602,N_21074,N_21959);
nor U23603 (N_23603,N_21416,N_22219);
and U23604 (N_23604,N_22162,N_21387);
nand U23605 (N_23605,N_21240,N_22015);
or U23606 (N_23606,N_21947,N_21004);
xnor U23607 (N_23607,N_21143,N_21253);
or U23608 (N_23608,N_22306,N_21341);
nand U23609 (N_23609,N_21342,N_21403);
nand U23610 (N_23610,N_22219,N_22021);
nand U23611 (N_23611,N_21776,N_21762);
and U23612 (N_23612,N_21134,N_21132);
xnor U23613 (N_23613,N_21913,N_22159);
nand U23614 (N_23614,N_22252,N_21786);
xnor U23615 (N_23615,N_22268,N_22007);
xor U23616 (N_23616,N_22454,N_21795);
nor U23617 (N_23617,N_22294,N_21067);
nor U23618 (N_23618,N_22417,N_21944);
nand U23619 (N_23619,N_22237,N_21698);
nand U23620 (N_23620,N_22449,N_21750);
or U23621 (N_23621,N_22091,N_22118);
nand U23622 (N_23622,N_21152,N_22347);
and U23623 (N_23623,N_22311,N_21862);
and U23624 (N_23624,N_22038,N_21151);
or U23625 (N_23625,N_21834,N_22377);
xnor U23626 (N_23626,N_21072,N_21724);
nor U23627 (N_23627,N_21296,N_21092);
xor U23628 (N_23628,N_21932,N_21356);
nor U23629 (N_23629,N_22296,N_21485);
or U23630 (N_23630,N_21544,N_21117);
xnor U23631 (N_23631,N_22292,N_21318);
xor U23632 (N_23632,N_21726,N_21183);
or U23633 (N_23633,N_21724,N_21678);
or U23634 (N_23634,N_22320,N_22487);
nand U23635 (N_23635,N_22454,N_22226);
or U23636 (N_23636,N_21353,N_22397);
nand U23637 (N_23637,N_21929,N_21366);
or U23638 (N_23638,N_22032,N_21017);
or U23639 (N_23639,N_21388,N_21381);
nand U23640 (N_23640,N_22190,N_21509);
and U23641 (N_23641,N_21823,N_21036);
xor U23642 (N_23642,N_22499,N_21647);
and U23643 (N_23643,N_21364,N_22019);
xnor U23644 (N_23644,N_21536,N_22283);
nand U23645 (N_23645,N_22343,N_21938);
nor U23646 (N_23646,N_22111,N_21598);
nor U23647 (N_23647,N_21221,N_21678);
nor U23648 (N_23648,N_21628,N_21323);
xnor U23649 (N_23649,N_21419,N_21306);
and U23650 (N_23650,N_21469,N_21108);
and U23651 (N_23651,N_22325,N_21108);
nand U23652 (N_23652,N_21535,N_22327);
and U23653 (N_23653,N_21512,N_21343);
nor U23654 (N_23654,N_21322,N_22379);
xor U23655 (N_23655,N_21660,N_21915);
or U23656 (N_23656,N_21242,N_21459);
nor U23657 (N_23657,N_21989,N_21005);
nor U23658 (N_23658,N_21745,N_22107);
nor U23659 (N_23659,N_21368,N_21699);
or U23660 (N_23660,N_21422,N_22387);
and U23661 (N_23661,N_21608,N_21420);
xor U23662 (N_23662,N_21744,N_22317);
xnor U23663 (N_23663,N_21488,N_21183);
xor U23664 (N_23664,N_21664,N_21769);
nor U23665 (N_23665,N_21827,N_21267);
xor U23666 (N_23666,N_21393,N_22436);
or U23667 (N_23667,N_21899,N_21232);
nand U23668 (N_23668,N_21484,N_21196);
nand U23669 (N_23669,N_22122,N_22172);
or U23670 (N_23670,N_21905,N_22127);
and U23671 (N_23671,N_22082,N_21991);
or U23672 (N_23672,N_21752,N_21942);
nor U23673 (N_23673,N_21886,N_22321);
and U23674 (N_23674,N_22015,N_22435);
nor U23675 (N_23675,N_22170,N_22117);
and U23676 (N_23676,N_22149,N_22154);
or U23677 (N_23677,N_21102,N_21388);
nand U23678 (N_23678,N_21974,N_21414);
or U23679 (N_23679,N_22404,N_22208);
nand U23680 (N_23680,N_21076,N_21398);
or U23681 (N_23681,N_22368,N_22123);
or U23682 (N_23682,N_21950,N_21876);
and U23683 (N_23683,N_21354,N_21693);
and U23684 (N_23684,N_22262,N_21607);
nor U23685 (N_23685,N_21239,N_21204);
nor U23686 (N_23686,N_22253,N_21090);
xor U23687 (N_23687,N_21139,N_22138);
or U23688 (N_23688,N_22445,N_22139);
and U23689 (N_23689,N_21147,N_21815);
xnor U23690 (N_23690,N_22453,N_21905);
and U23691 (N_23691,N_21168,N_22217);
or U23692 (N_23692,N_21581,N_22299);
or U23693 (N_23693,N_22469,N_21994);
or U23694 (N_23694,N_21653,N_21194);
nand U23695 (N_23695,N_21610,N_21530);
and U23696 (N_23696,N_21018,N_22189);
and U23697 (N_23697,N_22469,N_21481);
nand U23698 (N_23698,N_22104,N_21018);
nand U23699 (N_23699,N_22347,N_21548);
nand U23700 (N_23700,N_21829,N_21461);
or U23701 (N_23701,N_21425,N_21487);
or U23702 (N_23702,N_21359,N_21504);
and U23703 (N_23703,N_22431,N_21710);
and U23704 (N_23704,N_21968,N_21626);
or U23705 (N_23705,N_21311,N_22368);
and U23706 (N_23706,N_22020,N_21785);
nor U23707 (N_23707,N_21911,N_21592);
nand U23708 (N_23708,N_21177,N_22272);
nor U23709 (N_23709,N_21885,N_21345);
xor U23710 (N_23710,N_21821,N_22413);
xor U23711 (N_23711,N_22443,N_21776);
xor U23712 (N_23712,N_21925,N_22394);
or U23713 (N_23713,N_21270,N_21171);
xnor U23714 (N_23714,N_21070,N_21499);
or U23715 (N_23715,N_21935,N_21590);
or U23716 (N_23716,N_21059,N_22306);
nor U23717 (N_23717,N_21246,N_21865);
and U23718 (N_23718,N_21334,N_22204);
nand U23719 (N_23719,N_21496,N_21133);
nand U23720 (N_23720,N_21108,N_21474);
or U23721 (N_23721,N_21148,N_21875);
or U23722 (N_23722,N_22201,N_22019);
nand U23723 (N_23723,N_22386,N_22315);
and U23724 (N_23724,N_21894,N_21691);
nand U23725 (N_23725,N_21547,N_22309);
or U23726 (N_23726,N_21790,N_21987);
nand U23727 (N_23727,N_22104,N_22450);
xnor U23728 (N_23728,N_21727,N_21567);
or U23729 (N_23729,N_22141,N_21359);
xor U23730 (N_23730,N_22403,N_21213);
and U23731 (N_23731,N_21505,N_21062);
and U23732 (N_23732,N_21605,N_22032);
nor U23733 (N_23733,N_21651,N_22405);
or U23734 (N_23734,N_21707,N_21677);
nand U23735 (N_23735,N_21038,N_21569);
or U23736 (N_23736,N_22252,N_22420);
and U23737 (N_23737,N_21666,N_21451);
nor U23738 (N_23738,N_22405,N_22053);
or U23739 (N_23739,N_21113,N_21590);
xnor U23740 (N_23740,N_22289,N_22262);
and U23741 (N_23741,N_21593,N_22236);
or U23742 (N_23742,N_22251,N_21410);
nor U23743 (N_23743,N_22111,N_21934);
or U23744 (N_23744,N_21134,N_21365);
and U23745 (N_23745,N_21684,N_21401);
nor U23746 (N_23746,N_22423,N_21732);
nor U23747 (N_23747,N_22098,N_21235);
nand U23748 (N_23748,N_22487,N_21828);
nor U23749 (N_23749,N_21183,N_21277);
or U23750 (N_23750,N_21309,N_21885);
nand U23751 (N_23751,N_22288,N_21372);
nand U23752 (N_23752,N_22169,N_21504);
nand U23753 (N_23753,N_21031,N_22004);
or U23754 (N_23754,N_21481,N_21407);
and U23755 (N_23755,N_21967,N_21046);
nand U23756 (N_23756,N_21461,N_22474);
nand U23757 (N_23757,N_22134,N_21893);
xor U23758 (N_23758,N_21236,N_22222);
nor U23759 (N_23759,N_21800,N_22281);
xnor U23760 (N_23760,N_21329,N_22003);
nand U23761 (N_23761,N_21551,N_22275);
nor U23762 (N_23762,N_21829,N_21419);
and U23763 (N_23763,N_21955,N_22358);
or U23764 (N_23764,N_21582,N_22139);
nand U23765 (N_23765,N_22219,N_22023);
or U23766 (N_23766,N_21658,N_22226);
or U23767 (N_23767,N_21473,N_21147);
nor U23768 (N_23768,N_21796,N_21339);
and U23769 (N_23769,N_21475,N_22363);
or U23770 (N_23770,N_21720,N_21184);
nand U23771 (N_23771,N_22355,N_22409);
and U23772 (N_23772,N_21859,N_21133);
or U23773 (N_23773,N_22048,N_22301);
nand U23774 (N_23774,N_22437,N_22293);
nor U23775 (N_23775,N_21614,N_21396);
and U23776 (N_23776,N_21237,N_21888);
or U23777 (N_23777,N_21843,N_21309);
nand U23778 (N_23778,N_21051,N_22343);
nand U23779 (N_23779,N_21877,N_22130);
nand U23780 (N_23780,N_22285,N_21038);
nor U23781 (N_23781,N_21040,N_21207);
or U23782 (N_23782,N_22333,N_21838);
nor U23783 (N_23783,N_22377,N_21784);
nand U23784 (N_23784,N_21188,N_21763);
and U23785 (N_23785,N_21894,N_21500);
xor U23786 (N_23786,N_21384,N_21391);
nor U23787 (N_23787,N_21701,N_21602);
nor U23788 (N_23788,N_22376,N_21496);
nand U23789 (N_23789,N_21941,N_21667);
xor U23790 (N_23790,N_22100,N_22417);
and U23791 (N_23791,N_22413,N_21827);
and U23792 (N_23792,N_21234,N_21077);
and U23793 (N_23793,N_21021,N_22252);
or U23794 (N_23794,N_21354,N_22038);
nor U23795 (N_23795,N_22323,N_22469);
nor U23796 (N_23796,N_22413,N_22010);
xnor U23797 (N_23797,N_21245,N_21187);
or U23798 (N_23798,N_21214,N_22387);
xor U23799 (N_23799,N_21716,N_22486);
xnor U23800 (N_23800,N_21057,N_21221);
and U23801 (N_23801,N_21836,N_21319);
or U23802 (N_23802,N_22341,N_21889);
and U23803 (N_23803,N_22068,N_21942);
nand U23804 (N_23804,N_22123,N_21906);
nor U23805 (N_23805,N_21141,N_21673);
and U23806 (N_23806,N_21167,N_21345);
nor U23807 (N_23807,N_22325,N_21116);
and U23808 (N_23808,N_22428,N_22461);
nor U23809 (N_23809,N_22067,N_22056);
xor U23810 (N_23810,N_21193,N_21273);
nand U23811 (N_23811,N_22409,N_22489);
nor U23812 (N_23812,N_21379,N_21437);
or U23813 (N_23813,N_21152,N_21569);
nor U23814 (N_23814,N_21048,N_22307);
nand U23815 (N_23815,N_21284,N_21191);
nor U23816 (N_23816,N_21329,N_22195);
nand U23817 (N_23817,N_21926,N_21549);
xor U23818 (N_23818,N_21299,N_21177);
and U23819 (N_23819,N_21228,N_21726);
nor U23820 (N_23820,N_22182,N_21620);
or U23821 (N_23821,N_21117,N_22456);
xnor U23822 (N_23822,N_21408,N_21713);
and U23823 (N_23823,N_21513,N_22435);
or U23824 (N_23824,N_21654,N_21727);
and U23825 (N_23825,N_22249,N_22438);
xnor U23826 (N_23826,N_21845,N_21049);
nor U23827 (N_23827,N_22307,N_21387);
and U23828 (N_23828,N_21005,N_21137);
and U23829 (N_23829,N_21482,N_21508);
xor U23830 (N_23830,N_21860,N_21799);
xor U23831 (N_23831,N_21514,N_21593);
and U23832 (N_23832,N_21935,N_21392);
nor U23833 (N_23833,N_21349,N_21664);
or U23834 (N_23834,N_22309,N_22288);
and U23835 (N_23835,N_21692,N_21843);
or U23836 (N_23836,N_21100,N_21447);
or U23837 (N_23837,N_21273,N_22232);
or U23838 (N_23838,N_21956,N_21127);
and U23839 (N_23839,N_21443,N_21643);
xor U23840 (N_23840,N_22083,N_21385);
nand U23841 (N_23841,N_22097,N_22044);
nor U23842 (N_23842,N_21048,N_21695);
and U23843 (N_23843,N_21421,N_21854);
nor U23844 (N_23844,N_22494,N_21967);
nor U23845 (N_23845,N_22433,N_21280);
xor U23846 (N_23846,N_22035,N_21650);
or U23847 (N_23847,N_21767,N_22293);
and U23848 (N_23848,N_21274,N_22303);
nand U23849 (N_23849,N_22128,N_21958);
nand U23850 (N_23850,N_21072,N_21308);
nand U23851 (N_23851,N_21022,N_21603);
nor U23852 (N_23852,N_21781,N_21192);
xor U23853 (N_23853,N_22188,N_21232);
or U23854 (N_23854,N_21754,N_22212);
and U23855 (N_23855,N_21503,N_21228);
or U23856 (N_23856,N_22050,N_21173);
and U23857 (N_23857,N_21150,N_21358);
xor U23858 (N_23858,N_21355,N_21519);
or U23859 (N_23859,N_22135,N_21110);
and U23860 (N_23860,N_21391,N_21101);
xnor U23861 (N_23861,N_22363,N_21418);
nand U23862 (N_23862,N_22376,N_21254);
nor U23863 (N_23863,N_21709,N_22173);
or U23864 (N_23864,N_21868,N_22420);
xor U23865 (N_23865,N_22242,N_21134);
or U23866 (N_23866,N_21069,N_22496);
xor U23867 (N_23867,N_22371,N_21671);
nor U23868 (N_23868,N_22494,N_22478);
xor U23869 (N_23869,N_21748,N_22250);
xor U23870 (N_23870,N_22143,N_21168);
xor U23871 (N_23871,N_22127,N_21995);
nor U23872 (N_23872,N_22185,N_22266);
or U23873 (N_23873,N_22159,N_22349);
nand U23874 (N_23874,N_22224,N_21470);
nand U23875 (N_23875,N_21204,N_22154);
and U23876 (N_23876,N_22137,N_21867);
or U23877 (N_23877,N_21588,N_21636);
and U23878 (N_23878,N_21964,N_22482);
nand U23879 (N_23879,N_21445,N_21829);
and U23880 (N_23880,N_22449,N_22225);
and U23881 (N_23881,N_21050,N_21228);
and U23882 (N_23882,N_22402,N_21154);
nor U23883 (N_23883,N_21042,N_22487);
and U23884 (N_23884,N_21011,N_21750);
or U23885 (N_23885,N_21358,N_21947);
nand U23886 (N_23886,N_21320,N_21319);
nand U23887 (N_23887,N_22354,N_21702);
or U23888 (N_23888,N_22080,N_22259);
xnor U23889 (N_23889,N_22404,N_21729);
or U23890 (N_23890,N_21923,N_22496);
nor U23891 (N_23891,N_22074,N_21108);
or U23892 (N_23892,N_21654,N_21133);
nor U23893 (N_23893,N_22285,N_21185);
or U23894 (N_23894,N_21186,N_21263);
nor U23895 (N_23895,N_21924,N_22378);
xor U23896 (N_23896,N_21192,N_21797);
nand U23897 (N_23897,N_21292,N_21379);
nor U23898 (N_23898,N_22478,N_21279);
or U23899 (N_23899,N_21499,N_21078);
nand U23900 (N_23900,N_21521,N_22038);
nand U23901 (N_23901,N_22352,N_21683);
xnor U23902 (N_23902,N_21045,N_22214);
or U23903 (N_23903,N_22259,N_21500);
xor U23904 (N_23904,N_21947,N_21562);
and U23905 (N_23905,N_21278,N_21793);
or U23906 (N_23906,N_21267,N_21570);
xor U23907 (N_23907,N_21016,N_21891);
nand U23908 (N_23908,N_21280,N_21777);
and U23909 (N_23909,N_22489,N_21102);
and U23910 (N_23910,N_22375,N_21652);
nor U23911 (N_23911,N_21629,N_21916);
and U23912 (N_23912,N_21368,N_22250);
nor U23913 (N_23913,N_21843,N_22247);
and U23914 (N_23914,N_22464,N_21250);
nor U23915 (N_23915,N_21159,N_22121);
nor U23916 (N_23916,N_22444,N_21257);
and U23917 (N_23917,N_22386,N_22493);
and U23918 (N_23918,N_21771,N_21623);
xnor U23919 (N_23919,N_22379,N_21514);
or U23920 (N_23920,N_21601,N_22189);
xnor U23921 (N_23921,N_21196,N_21853);
xnor U23922 (N_23922,N_21388,N_22436);
and U23923 (N_23923,N_21672,N_22314);
or U23924 (N_23924,N_22244,N_21679);
or U23925 (N_23925,N_21687,N_21450);
nand U23926 (N_23926,N_22487,N_21340);
and U23927 (N_23927,N_21897,N_22358);
and U23928 (N_23928,N_22182,N_21661);
and U23929 (N_23929,N_21856,N_22476);
nor U23930 (N_23930,N_21633,N_21089);
xnor U23931 (N_23931,N_22339,N_21082);
nand U23932 (N_23932,N_21011,N_22340);
and U23933 (N_23933,N_21122,N_21063);
nor U23934 (N_23934,N_21045,N_21453);
xor U23935 (N_23935,N_21327,N_21936);
xnor U23936 (N_23936,N_21000,N_22171);
xor U23937 (N_23937,N_21637,N_21763);
xnor U23938 (N_23938,N_22250,N_21654);
and U23939 (N_23939,N_21789,N_21716);
or U23940 (N_23940,N_21806,N_21197);
xor U23941 (N_23941,N_22343,N_22045);
nor U23942 (N_23942,N_22217,N_21389);
nor U23943 (N_23943,N_21413,N_22144);
nand U23944 (N_23944,N_22493,N_22001);
or U23945 (N_23945,N_21642,N_22103);
nor U23946 (N_23946,N_22250,N_21715);
and U23947 (N_23947,N_22008,N_21065);
or U23948 (N_23948,N_21291,N_21737);
or U23949 (N_23949,N_21100,N_22110);
or U23950 (N_23950,N_21581,N_21167);
or U23951 (N_23951,N_21763,N_22459);
nor U23952 (N_23952,N_21922,N_22217);
and U23953 (N_23953,N_22476,N_21945);
nand U23954 (N_23954,N_21079,N_21058);
and U23955 (N_23955,N_21870,N_22017);
and U23956 (N_23956,N_22420,N_21174);
and U23957 (N_23957,N_21287,N_21188);
and U23958 (N_23958,N_21840,N_21123);
or U23959 (N_23959,N_22423,N_21929);
nor U23960 (N_23960,N_22242,N_21128);
nand U23961 (N_23961,N_21449,N_21713);
or U23962 (N_23962,N_22197,N_21409);
and U23963 (N_23963,N_21694,N_21692);
nor U23964 (N_23964,N_21827,N_22218);
nor U23965 (N_23965,N_22330,N_21426);
and U23966 (N_23966,N_21340,N_22144);
xor U23967 (N_23967,N_22197,N_21052);
nand U23968 (N_23968,N_21910,N_22429);
xor U23969 (N_23969,N_21245,N_22100);
xnor U23970 (N_23970,N_21428,N_21568);
xor U23971 (N_23971,N_21292,N_21662);
nand U23972 (N_23972,N_21868,N_22046);
and U23973 (N_23973,N_21216,N_22164);
xor U23974 (N_23974,N_21161,N_21289);
xnor U23975 (N_23975,N_22400,N_22092);
or U23976 (N_23976,N_22081,N_21740);
xor U23977 (N_23977,N_22364,N_22212);
and U23978 (N_23978,N_22163,N_21987);
or U23979 (N_23979,N_22022,N_21552);
and U23980 (N_23980,N_21985,N_21718);
xor U23981 (N_23981,N_21384,N_22013);
xor U23982 (N_23982,N_21595,N_22157);
xor U23983 (N_23983,N_21998,N_21314);
nor U23984 (N_23984,N_21566,N_21907);
nor U23985 (N_23985,N_21086,N_22263);
or U23986 (N_23986,N_21372,N_21163);
and U23987 (N_23987,N_21253,N_21000);
nor U23988 (N_23988,N_21584,N_21813);
and U23989 (N_23989,N_22059,N_21782);
nor U23990 (N_23990,N_21060,N_21600);
and U23991 (N_23991,N_21635,N_21222);
or U23992 (N_23992,N_21033,N_21316);
and U23993 (N_23993,N_21753,N_21963);
or U23994 (N_23994,N_21967,N_21234);
nand U23995 (N_23995,N_22032,N_22132);
or U23996 (N_23996,N_21760,N_21537);
or U23997 (N_23997,N_21351,N_22317);
or U23998 (N_23998,N_22099,N_21952);
nor U23999 (N_23999,N_21480,N_22384);
nor U24000 (N_24000,N_22745,N_22818);
nor U24001 (N_24001,N_23434,N_23762);
nor U24002 (N_24002,N_23484,N_22506);
xor U24003 (N_24003,N_22791,N_23346);
and U24004 (N_24004,N_23756,N_23715);
xor U24005 (N_24005,N_23776,N_23724);
and U24006 (N_24006,N_23148,N_23304);
nand U24007 (N_24007,N_23009,N_23576);
nor U24008 (N_24008,N_23183,N_23510);
or U24009 (N_24009,N_23508,N_23401);
nand U24010 (N_24010,N_23769,N_22652);
xor U24011 (N_24011,N_22517,N_22642);
and U24012 (N_24012,N_23624,N_23109);
or U24013 (N_24013,N_23774,N_22696);
or U24014 (N_24014,N_22737,N_23988);
or U24015 (N_24015,N_23651,N_23477);
xor U24016 (N_24016,N_23034,N_23515);
or U24017 (N_24017,N_23259,N_22631);
and U24018 (N_24018,N_22741,N_23619);
nand U24019 (N_24019,N_23408,N_22606);
xor U24020 (N_24020,N_22688,N_23425);
and U24021 (N_24021,N_23823,N_23439);
nor U24022 (N_24022,N_23302,N_23656);
or U24023 (N_24023,N_23683,N_23893);
xnor U24024 (N_24024,N_22985,N_23303);
xnor U24025 (N_24025,N_23815,N_23443);
nand U24026 (N_24026,N_23940,N_23523);
or U24027 (N_24027,N_22984,N_23432);
and U24028 (N_24028,N_22601,N_22739);
xor U24029 (N_24029,N_23696,N_23778);
nand U24030 (N_24030,N_23031,N_22844);
nor U24031 (N_24031,N_22882,N_22880);
xor U24032 (N_24032,N_23305,N_22525);
or U24033 (N_24033,N_22563,N_23190);
nand U24034 (N_24034,N_23121,N_22596);
xnor U24035 (N_24035,N_23688,N_22807);
or U24036 (N_24036,N_22928,N_23060);
nand U24037 (N_24037,N_23344,N_22616);
nand U24038 (N_24038,N_23935,N_22997);
xnor U24039 (N_24039,N_23565,N_22521);
or U24040 (N_24040,N_23603,N_23937);
xnor U24041 (N_24041,N_22780,N_22542);
or U24042 (N_24042,N_23520,N_23705);
or U24043 (N_24043,N_23637,N_23743);
nand U24044 (N_24044,N_23597,N_22982);
nor U24045 (N_24045,N_22874,N_23197);
xor U24046 (N_24046,N_23525,N_22862);
and U24047 (N_24047,N_23822,N_22940);
nand U24048 (N_24048,N_23154,N_23051);
and U24049 (N_24049,N_22678,N_23793);
nand U24050 (N_24050,N_23518,N_23755);
or U24051 (N_24051,N_23638,N_22813);
xor U24052 (N_24052,N_23287,N_22715);
xnor U24053 (N_24053,N_23693,N_23005);
or U24054 (N_24054,N_23646,N_23699);
nand U24055 (N_24055,N_23248,N_23065);
or U24056 (N_24056,N_22538,N_23224);
or U24057 (N_24057,N_23332,N_22593);
nor U24058 (N_24058,N_22574,N_22812);
xor U24059 (N_24059,N_22788,N_22580);
nand U24060 (N_24060,N_22838,N_22733);
nand U24061 (N_24061,N_22988,N_23045);
nor U24062 (N_24062,N_23751,N_23772);
nand U24063 (N_24063,N_23609,N_23904);
or U24064 (N_24064,N_22981,N_22938);
or U24065 (N_24065,N_23560,N_23278);
and U24066 (N_24066,N_22720,N_22529);
or U24067 (N_24067,N_23113,N_22568);
and U24068 (N_24068,N_22846,N_23294);
xor U24069 (N_24069,N_22775,N_23008);
xnor U24070 (N_24070,N_23285,N_23410);
nor U24071 (N_24071,N_22700,N_23843);
and U24072 (N_24072,N_23440,N_22948);
nand U24073 (N_24073,N_23268,N_22570);
or U24074 (N_24074,N_22600,N_23633);
nand U24075 (N_24075,N_23747,N_23883);
or U24076 (N_24076,N_23878,N_23276);
nor U24077 (N_24077,N_23959,N_22833);
nand U24078 (N_24078,N_22528,N_23036);
nor U24079 (N_24079,N_22725,N_23295);
nand U24080 (N_24080,N_22522,N_22539);
xor U24081 (N_24081,N_23068,N_23389);
and U24082 (N_24082,N_23375,N_22835);
xor U24083 (N_24083,N_22668,N_23986);
nor U24084 (N_24084,N_23577,N_23249);
xor U24085 (N_24085,N_22625,N_22577);
or U24086 (N_24086,N_23029,N_23606);
or U24087 (N_24087,N_22787,N_23236);
and U24088 (N_24088,N_23385,N_22967);
xnor U24089 (N_24089,N_23451,N_22507);
and U24090 (N_24090,N_23899,N_23067);
or U24091 (N_24091,N_23080,N_22943);
xnor U24092 (N_24092,N_23101,N_23469);
xnor U24093 (N_24093,N_22626,N_23813);
nor U24094 (N_24094,N_23483,N_22659);
and U24095 (N_24095,N_22935,N_23417);
or U24096 (N_24096,N_23460,N_23164);
or U24097 (N_24097,N_22890,N_23003);
or U24098 (N_24098,N_22803,N_23157);
or U24099 (N_24099,N_23966,N_23313);
xnor U24100 (N_24100,N_23501,N_23330);
and U24101 (N_24101,N_23889,N_23876);
or U24102 (N_24102,N_23455,N_23915);
xnor U24103 (N_24103,N_22591,N_23342);
nand U24104 (N_24104,N_22508,N_22530);
or U24105 (N_24105,N_23012,N_23186);
or U24106 (N_24106,N_23253,N_23407);
nand U24107 (N_24107,N_23674,N_23396);
and U24108 (N_24108,N_23569,N_23108);
nand U24109 (N_24109,N_23139,N_23409);
nand U24110 (N_24110,N_22930,N_23886);
nor U24111 (N_24111,N_22698,N_23329);
nand U24112 (N_24112,N_22755,N_23226);
and U24113 (N_24113,N_22744,N_22964);
or U24114 (N_24114,N_23708,N_23559);
or U24115 (N_24115,N_22876,N_23445);
and U24116 (N_24116,N_23710,N_23522);
nor U24117 (N_24117,N_22918,N_23640);
nor U24118 (N_24118,N_23777,N_22808);
nor U24119 (N_24119,N_22996,N_23496);
nor U24120 (N_24120,N_22629,N_22978);
nand U24121 (N_24121,N_22947,N_22977);
nor U24122 (N_24122,N_23561,N_22735);
xnor U24123 (N_24123,N_22848,N_22802);
and U24124 (N_24124,N_23430,N_23908);
nand U24125 (N_24125,N_23262,N_23393);
or U24126 (N_24126,N_23798,N_22841);
nand U24127 (N_24127,N_22965,N_22792);
xor U24128 (N_24128,N_23703,N_23614);
nand U24129 (N_24129,N_23931,N_23392);
or U24130 (N_24130,N_22630,N_23079);
and U24131 (N_24131,N_22582,N_22853);
or U24132 (N_24132,N_22878,N_22676);
xnor U24133 (N_24133,N_23568,N_22576);
and U24134 (N_24134,N_23978,N_23814);
or U24135 (N_24135,N_23837,N_23394);
nor U24136 (N_24136,N_23310,N_22702);
nor U24137 (N_24137,N_22915,N_23205);
xnor U24138 (N_24138,N_23037,N_22781);
xor U24139 (N_24139,N_23807,N_23076);
nand U24140 (N_24140,N_22681,N_23449);
or U24141 (N_24141,N_22974,N_23070);
xor U24142 (N_24142,N_22973,N_23676);
xor U24143 (N_24143,N_23232,N_23691);
xor U24144 (N_24144,N_22860,N_23082);
nor U24145 (N_24145,N_23879,N_23943);
and U24146 (N_24146,N_23073,N_23675);
or U24147 (N_24147,N_23093,N_22502);
and U24148 (N_24148,N_23869,N_22881);
nand U24149 (N_24149,N_23855,N_23120);
or U24150 (N_24150,N_22815,N_23307);
or U24151 (N_24151,N_23198,N_22583);
nand U24152 (N_24152,N_23549,N_22597);
and U24153 (N_24153,N_22913,N_23605);
xor U24154 (N_24154,N_23413,N_22857);
and U24155 (N_24155,N_23433,N_23763);
xor U24156 (N_24156,N_22959,N_23150);
nor U24157 (N_24157,N_23088,N_23907);
or U24158 (N_24158,N_23384,N_23880);
or U24159 (N_24159,N_22885,N_23103);
and U24160 (N_24160,N_22843,N_22799);
and U24161 (N_24161,N_23898,N_23402);
nor U24162 (N_24162,N_23970,N_22670);
nor U24163 (N_24163,N_22758,N_23475);
nor U24164 (N_24164,N_23511,N_23352);
or U24165 (N_24165,N_22581,N_23492);
and U24166 (N_24166,N_23997,N_23206);
nor U24167 (N_24167,N_23348,N_22557);
xor U24168 (N_24168,N_23136,N_23507);
or U24169 (N_24169,N_23246,N_22760);
xnor U24170 (N_24170,N_23336,N_22872);
nor U24171 (N_24171,N_23438,N_23854);
and U24172 (N_24172,N_23465,N_23601);
or U24173 (N_24173,N_23064,N_23053);
xnor U24174 (N_24174,N_23398,N_23238);
and U24175 (N_24175,N_22695,N_23494);
nand U24176 (N_24176,N_23579,N_23820);
xor U24177 (N_24177,N_22692,N_22953);
nand U24178 (N_24178,N_23290,N_23578);
nand U24179 (N_24179,N_23766,N_23144);
nand U24180 (N_24180,N_22518,N_23547);
or U24181 (N_24181,N_22786,N_23953);
xnor U24182 (N_24182,N_23191,N_22510);
nand U24183 (N_24183,N_23868,N_22889);
nand U24184 (N_24184,N_23337,N_23370);
or U24185 (N_24185,N_22613,N_22536);
and U24186 (N_24186,N_22635,N_22732);
or U24187 (N_24187,N_22794,N_22654);
and U24188 (N_24188,N_22908,N_23939);
nand U24189 (N_24189,N_23857,N_22699);
nor U24190 (N_24190,N_22620,N_23063);
and U24191 (N_24191,N_23944,N_22736);
nand U24192 (N_24192,N_23240,N_23308);
xnor U24193 (N_24193,N_23821,N_23237);
or U24194 (N_24194,N_23200,N_23096);
xor U24195 (N_24195,N_23277,N_23531);
xor U24196 (N_24196,N_23870,N_22810);
or U24197 (N_24197,N_22672,N_22968);
or U24198 (N_24198,N_23718,N_23553);
nor U24199 (N_24199,N_23324,N_22936);
and U24200 (N_24200,N_22774,N_23618);
nor U24201 (N_24201,N_23833,N_23583);
xnor U24202 (N_24202,N_23626,N_22979);
and U24203 (N_24203,N_23851,N_23671);
and U24204 (N_24204,N_23625,N_22541);
nor U24205 (N_24205,N_22624,N_22571);
nand U24206 (N_24206,N_23506,N_23901);
nor U24207 (N_24207,N_23266,N_22925);
and U24208 (N_24208,N_23975,N_23830);
or U24209 (N_24209,N_23875,N_23172);
or U24210 (N_24210,N_22500,N_22865);
or U24211 (N_24211,N_22648,N_23419);
or U24212 (N_24212,N_23351,N_22893);
or U24213 (N_24213,N_23958,N_23156);
nor U24214 (N_24214,N_23802,N_23846);
nand U24215 (N_24215,N_22937,N_23229);
or U24216 (N_24216,N_23087,N_22638);
xnor U24217 (N_24217,N_23590,N_22734);
nor U24218 (N_24218,N_22859,N_23428);
xnor U24219 (N_24219,N_22868,N_23215);
xnor U24220 (N_24220,N_22640,N_23620);
or U24221 (N_24221,N_22962,N_22592);
xnor U24222 (N_24222,N_23949,N_23900);
and U24223 (N_24223,N_23784,N_23025);
xor U24224 (N_24224,N_23530,N_23887);
nand U24225 (N_24225,N_23829,N_23994);
or U24226 (N_24226,N_23098,N_23104);
and U24227 (N_24227,N_22759,N_23357);
and U24228 (N_24228,N_23414,N_23733);
and U24229 (N_24229,N_23890,N_22867);
xnor U24230 (N_24230,N_23759,N_23704);
nand U24231 (N_24231,N_23669,N_23977);
nand U24232 (N_24232,N_22817,N_23049);
nand U24233 (N_24233,N_23859,N_23922);
nor U24234 (N_24234,N_23202,N_22708);
and U24235 (N_24235,N_23527,N_22726);
nand U24236 (N_24236,N_23666,N_23380);
xnor U24237 (N_24237,N_23126,N_22513);
nor U24238 (N_24238,N_23074,N_23368);
or U24239 (N_24239,N_23946,N_23378);
nand U24240 (N_24240,N_23300,N_23423);
xor U24241 (N_24241,N_23453,N_23461);
or U24242 (N_24242,N_22680,N_23111);
nand U24243 (N_24243,N_22628,N_23149);
nor U24244 (N_24244,N_23916,N_23657);
nor U24245 (N_24245,N_23291,N_23299);
and U24246 (N_24246,N_22686,N_23686);
and U24247 (N_24247,N_23968,N_23081);
nor U24248 (N_24248,N_23957,N_23424);
and U24249 (N_24249,N_23347,N_23474);
and U24250 (N_24250,N_23914,N_23002);
and U24251 (N_24251,N_22797,N_23399);
nand U24252 (N_24252,N_23083,N_23539);
nor U24253 (N_24253,N_23631,N_22611);
or U24254 (N_24254,N_23697,N_23545);
nand U24255 (N_24255,N_23600,N_23207);
xnor U24256 (N_24256,N_23932,N_23091);
xor U24257 (N_24257,N_23589,N_22963);
and U24258 (N_24258,N_23193,N_23827);
or U24259 (N_24259,N_22907,N_23864);
nor U24260 (N_24260,N_22669,N_22801);
xnor U24261 (N_24261,N_23279,N_23143);
xnor U24262 (N_24262,N_22607,N_23538);
nor U24263 (N_24263,N_23418,N_22924);
xor U24264 (N_24264,N_23487,N_23613);
nor U24265 (N_24265,N_22748,N_23790);
and U24266 (N_24266,N_23905,N_23644);
xnor U24267 (N_24267,N_23698,N_23526);
and U24268 (N_24268,N_23092,N_22995);
or U24269 (N_24269,N_22809,N_23209);
xor U24270 (N_24270,N_22746,N_23714);
and U24271 (N_24271,N_23142,N_22683);
nand U24272 (N_24272,N_23188,N_23540);
or U24273 (N_24273,N_23220,N_22713);
and U24274 (N_24274,N_23885,N_23086);
nand U24275 (N_24275,N_23273,N_22667);
or U24276 (N_24276,N_23667,N_22831);
or U24277 (N_24277,N_22604,N_23095);
nand U24278 (N_24278,N_23834,N_23804);
nand U24279 (N_24279,N_23261,N_23680);
nand U24280 (N_24280,N_23764,N_22863);
nor U24281 (N_24281,N_23996,N_23405);
nor U24282 (N_24282,N_22641,N_22605);
or U24283 (N_24283,N_23653,N_22795);
xor U24284 (N_24284,N_22850,N_23479);
nand U24285 (N_24285,N_23773,N_22891);
or U24286 (N_24286,N_23865,N_23873);
nand U24287 (N_24287,N_23591,N_23860);
nand U24288 (N_24288,N_23493,N_22989);
nor U24289 (N_24289,N_23789,N_23061);
nand U24290 (N_24290,N_22697,N_23811);
xor U24291 (N_24291,N_22703,N_23296);
nor U24292 (N_24292,N_22911,N_23754);
xnor U24293 (N_24293,N_22598,N_23967);
nor U24294 (N_24294,N_23364,N_23588);
nor U24295 (N_24295,N_22821,N_23203);
xor U24296 (N_24296,N_22599,N_23806);
and U24297 (N_24297,N_23623,N_23331);
xnor U24298 (N_24298,N_23367,N_23557);
nor U24299 (N_24299,N_23738,N_22694);
or U24300 (N_24300,N_22728,N_23000);
xor U24301 (N_24301,N_23020,N_22994);
or U24302 (N_24302,N_22951,N_22722);
xnor U24303 (N_24303,N_23952,N_23217);
nor U24304 (N_24304,N_22705,N_23670);
xor U24305 (N_24305,N_23519,N_23488);
xnor U24306 (N_24306,N_23356,N_23628);
nor U24307 (N_24307,N_22960,N_23562);
xnor U24308 (N_24308,N_23403,N_23159);
nand U24309 (N_24309,N_23228,N_23742);
or U24310 (N_24310,N_23251,N_22840);
or U24311 (N_24311,N_23318,N_23981);
and U24312 (N_24312,N_23912,N_23586);
nor U24313 (N_24313,N_22990,N_23884);
xor U24314 (N_24314,N_23643,N_22800);
nor U24315 (N_24315,N_22651,N_22939);
xor U24316 (N_24316,N_23016,N_23011);
and U24317 (N_24317,N_23223,N_23818);
xnor U24318 (N_24318,N_22742,N_23819);
xnor U24319 (N_24319,N_23976,N_22776);
or U24320 (N_24320,N_22905,N_22917);
nor U24321 (N_24321,N_22552,N_23701);
and U24322 (N_24322,N_22553,N_23642);
xor U24323 (N_24323,N_22828,N_22569);
nor U24324 (N_24324,N_23750,N_23564);
xnor U24325 (N_24325,N_23436,N_23335);
nor U24326 (N_24326,N_22766,N_23963);
or U24327 (N_24327,N_22969,N_22712);
or U24328 (N_24328,N_23309,N_23993);
xnor U24329 (N_24329,N_23635,N_23138);
nand U24330 (N_24330,N_23711,N_22826);
nor U24331 (N_24331,N_22645,N_22639);
or U24332 (N_24332,N_22887,N_23544);
or U24333 (N_24333,N_23482,N_22509);
or U24334 (N_24334,N_22816,N_22608);
nand U24335 (N_24335,N_23171,N_23141);
nor U24336 (N_24336,N_23166,N_23298);
nor U24337 (N_24337,N_23555,N_22782);
and U24338 (N_24338,N_23316,N_22723);
xnor U24339 (N_24339,N_22926,N_22655);
or U24340 (N_24340,N_23566,N_23546);
and U24341 (N_24341,N_22901,N_22514);
and U24342 (N_24342,N_22886,N_23684);
and U24343 (N_24343,N_23616,N_23489);
nand U24344 (N_24344,N_22549,N_23575);
and U24345 (N_24345,N_23604,N_23416);
xor U24346 (N_24346,N_22866,N_22796);
and U24347 (N_24347,N_23354,N_22614);
nor U24348 (N_24348,N_22830,N_23896);
nor U24349 (N_24349,N_23582,N_23964);
nand U24350 (N_24350,N_22677,N_22823);
or U24351 (N_24351,N_23119,N_23690);
xor U24352 (N_24352,N_23892,N_23841);
nor U24353 (N_24353,N_22658,N_23805);
xor U24354 (N_24354,N_22559,N_22869);
xnor U24355 (N_24355,N_22798,N_23731);
nor U24356 (N_24356,N_23785,N_22532);
nand U24357 (N_24357,N_22661,N_23945);
nor U24358 (N_24358,N_23168,N_23258);
or U24359 (N_24359,N_23874,N_23381);
xor U24360 (N_24360,N_23383,N_22535);
xnor U24361 (N_24361,N_23788,N_23938);
xor U24362 (N_24362,N_23481,N_22785);
xor U24363 (N_24363,N_23881,N_22949);
nor U24364 (N_24364,N_22546,N_23219);
and U24365 (N_24365,N_22855,N_23151);
nand U24366 (N_24366,N_22916,N_23412);
nand U24367 (N_24367,N_22912,N_23225);
and U24368 (N_24368,N_22660,N_23021);
or U24369 (N_24369,N_23809,N_23973);
nor U24370 (N_24370,N_22545,N_23326);
nand U24371 (N_24371,N_23077,N_23752);
xnor U24372 (N_24372,N_23388,N_23235);
xnor U24373 (N_24373,N_23127,N_23283);
nand U24374 (N_24374,N_23639,N_23222);
xor U24375 (N_24375,N_23694,N_22665);
xor U24376 (N_24376,N_23230,N_23182);
xor U24377 (N_24377,N_23786,N_22673);
xnor U24378 (N_24378,N_23252,N_22523);
or U24379 (N_24379,N_23180,N_22684);
nand U24380 (N_24380,N_23075,N_22729);
nand U24381 (N_24381,N_23196,N_22738);
or U24382 (N_24382,N_23122,N_23594);
or U24383 (N_24383,N_23926,N_23660);
nand U24384 (N_24384,N_23599,N_23286);
and U24385 (N_24385,N_23343,N_22675);
or U24386 (N_24386,N_23800,N_22870);
xor U24387 (N_24387,N_22527,N_23374);
or U24388 (N_24388,N_23214,N_23779);
nand U24389 (N_24389,N_23395,N_22824);
xnor U24390 (N_24390,N_22589,N_23695);
or U24391 (N_24391,N_23132,N_23333);
or U24392 (N_24392,N_23028,N_22743);
nor U24393 (N_24393,N_22556,N_22691);
xor U24394 (N_24394,N_23231,N_23850);
xnor U24395 (N_24395,N_23706,N_22615);
nor U24396 (N_24396,N_23289,N_22664);
and U24397 (N_24397,N_23737,N_23001);
and U24398 (N_24398,N_22501,N_23450);
and U24399 (N_24399,N_23580,N_23170);
nor U24400 (N_24400,N_22879,N_22537);
and U24401 (N_24401,N_22544,N_22922);
xnor U24402 (N_24402,N_23467,N_23882);
nand U24403 (N_24403,N_23210,N_23543);
and U24404 (N_24404,N_23421,N_23117);
or U24405 (N_24405,N_23462,N_23221);
nor U24406 (N_24406,N_23971,N_23145);
and U24407 (N_24407,N_22554,N_23845);
nor U24408 (N_24408,N_23794,N_22612);
nand U24409 (N_24409,N_23853,N_23528);
or U24410 (N_24410,N_23542,N_22883);
and U24411 (N_24411,N_22561,N_22933);
and U24412 (N_24412,N_23504,N_22820);
and U24413 (N_24413,N_23247,N_23116);
and U24414 (N_24414,N_23816,N_23019);
or U24415 (N_24415,N_23133,N_22632);
or U24416 (N_24416,N_22772,N_23140);
nand U24417 (N_24417,N_22573,N_23571);
xor U24418 (N_24418,N_23740,N_23371);
nor U24419 (N_24419,N_23022,N_22590);
nor U24420 (N_24420,N_23535,N_22849);
or U24421 (N_24421,N_23292,N_23288);
or U24422 (N_24422,N_23721,N_23529);
xor U24423 (N_24423,N_23563,N_23181);
xor U24424 (N_24424,N_22927,N_22971);
and U24425 (N_24425,N_23204,N_23801);
and U24426 (N_24426,N_22649,N_22836);
xor U24427 (N_24427,N_23062,N_23263);
and U24428 (N_24428,N_22618,N_23100);
nand U24429 (N_24429,N_23505,N_23930);
xnor U24430 (N_24430,N_23315,N_23741);
or U24431 (N_24431,N_23573,N_22839);
xnor U24432 (N_24432,N_23345,N_23652);
nor U24433 (N_24433,N_23498,N_23163);
xor U24434 (N_24434,N_22534,N_23934);
xnor U24435 (N_24435,N_22769,N_23612);
nand U24436 (N_24436,N_23645,N_23720);
nand U24437 (N_24437,N_23610,N_23856);
or U24438 (N_24438,N_23534,N_23334);
or U24439 (N_24439,N_23458,N_22627);
nand U24440 (N_24440,N_22762,N_23135);
nor U24441 (N_24441,N_23495,N_23089);
nor U24442 (N_24442,N_23727,N_23010);
and U24443 (N_24443,N_22656,N_22966);
nand U24444 (N_24444,N_23211,N_22992);
xnor U24445 (N_24445,N_23463,N_23570);
nand U24446 (N_24446,N_23152,N_23679);
nor U24447 (N_24447,N_22643,N_22942);
nor U24448 (N_24448,N_22650,N_23057);
nand U24449 (N_24449,N_23924,N_23312);
xnor U24450 (N_24450,N_23602,N_23466);
nor U24451 (N_24451,N_23218,N_23947);
and U24452 (N_24452,N_23105,N_22647);
nor U24453 (N_24453,N_22690,N_23941);
xor U24454 (N_24454,N_23004,N_22829);
xnor U24455 (N_24455,N_23473,N_22934);
nand U24456 (N_24456,N_22904,N_23194);
nor U24457 (N_24457,N_23376,N_22771);
and U24458 (N_24458,N_23838,N_23014);
or U24459 (N_24459,N_22610,N_22920);
or U24460 (N_24460,N_22636,N_23340);
nand U24461 (N_24461,N_23744,N_23842);
xnor U24462 (N_24462,N_22819,N_22991);
and U24463 (N_24463,N_23983,N_22856);
nand U24464 (N_24464,N_22619,N_23867);
or U24465 (N_24465,N_23244,N_22531);
nand U24466 (N_24466,N_23866,N_23390);
and U24467 (N_24467,N_23621,N_23084);
nor U24468 (N_24468,N_23275,N_23491);
xnor U24469 (N_24469,N_23179,N_23212);
nor U24470 (N_24470,N_23353,N_23464);
nand U24471 (N_24471,N_23713,N_23007);
nand U24472 (N_24472,N_23245,N_22790);
nand U24473 (N_24473,N_23046,N_23685);
and U24474 (N_24474,N_23596,N_23707);
xnor U24475 (N_24475,N_23783,N_22644);
or U24476 (N_24476,N_23677,N_22754);
and U24477 (N_24477,N_23611,N_23655);
and U24478 (N_24478,N_23849,N_23189);
and U24479 (N_24479,N_22749,N_23533);
or U24480 (N_24480,N_22761,N_23114);
nand U24481 (N_24481,N_23749,N_23863);
or U24482 (N_24482,N_22701,N_23782);
or U24483 (N_24483,N_22789,N_23629);
xor U24484 (N_24484,N_22747,N_23270);
nor U24485 (N_24485,N_22567,N_23282);
nand U24486 (N_24486,N_22950,N_23745);
or U24487 (N_24487,N_23636,N_23961);
and U24488 (N_24488,N_23593,N_22842);
xor U24489 (N_24489,N_23293,N_22814);
nand U24490 (N_24490,N_23765,N_23895);
and U24491 (N_24491,N_23584,N_23592);
or U24492 (N_24492,N_23072,N_22609);
xor U24493 (N_24493,N_23928,N_22986);
or U24494 (N_24494,N_23227,N_22674);
or U24495 (N_24495,N_23648,N_22623);
xor U24496 (N_24496,N_23341,N_23269);
and U24497 (N_24497,N_23585,N_23317);
and U24498 (N_24498,N_23391,N_22919);
nor U24499 (N_24499,N_23955,N_22634);
or U24500 (N_24500,N_23942,N_23426);
xor U24501 (N_24501,N_23826,N_23195);
xor U24502 (N_24502,N_22983,N_23722);
nor U24503 (N_24503,N_23897,N_23129);
xnor U24504 (N_24504,N_23906,N_22515);
nand U24505 (N_24505,N_23835,N_22822);
or U24506 (N_24506,N_22520,N_23954);
nand U24507 (N_24507,N_23689,N_23558);
xor U24508 (N_24508,N_22564,N_23572);
or U24509 (N_24509,N_22767,N_23243);
and U24510 (N_24510,N_22566,N_22779);
or U24511 (N_24511,N_22730,N_23369);
nor U24512 (N_24512,N_22827,N_23681);
and U24513 (N_24513,N_23716,N_22903);
or U24514 (N_24514,N_23687,N_23536);
and U24515 (N_24515,N_23732,N_23918);
nand U24516 (N_24516,N_23411,N_22896);
xor U24517 (N_24517,N_23662,N_23476);
or U24518 (N_24518,N_22718,N_22679);
nand U24519 (N_24519,N_22714,N_23987);
xnor U24520 (N_24520,N_22717,N_23052);
xnor U24521 (N_24521,N_22533,N_23658);
nor U24522 (N_24522,N_22946,N_23349);
or U24523 (N_24523,N_23760,N_23775);
nor U24524 (N_24524,N_23272,N_23023);
and U24525 (N_24525,N_23516,N_23808);
or U24526 (N_24526,N_23128,N_23260);
or U24527 (N_24527,N_22871,N_22551);
xnor U24528 (N_24528,N_23951,N_23692);
nor U24529 (N_24529,N_23124,N_23950);
xor U24530 (N_24530,N_23264,N_22633);
nand U24531 (N_24531,N_23162,N_23567);
or U24532 (N_24532,N_22897,N_22858);
or U24533 (N_24533,N_22671,N_23615);
nand U24534 (N_24534,N_23991,N_23902);
nor U24535 (N_24535,N_22864,N_23982);
and U24536 (N_24536,N_23017,N_23948);
and U24537 (N_24537,N_22540,N_23472);
nor U24538 (N_24538,N_23137,N_23118);
and U24539 (N_24539,N_23574,N_22764);
xnor U24540 (N_24540,N_22768,N_23131);
or U24541 (N_24541,N_23106,N_23709);
and U24542 (N_24542,N_22902,N_23791);
and U24543 (N_24543,N_22503,N_22961);
nor U24544 (N_24544,N_23406,N_23847);
nand U24545 (N_24545,N_22765,N_23085);
or U24546 (N_24546,N_23598,N_23123);
nor U24547 (N_24547,N_23267,N_22892);
nand U24548 (N_24548,N_23632,N_22832);
nand U24549 (N_24549,N_23832,N_23537);
xor U24550 (N_24550,N_22877,N_22751);
xnor U24551 (N_24551,N_23386,N_22910);
or U24552 (N_24552,N_22783,N_23725);
or U24553 (N_24553,N_23158,N_23055);
nor U24554 (N_24554,N_22572,N_22516);
nand U24555 (N_24555,N_22716,N_23446);
nand U24556 (N_24556,N_22952,N_23812);
nor U24557 (N_24557,N_23470,N_23497);
nor U24558 (N_24558,N_23927,N_23254);
or U24559 (N_24559,N_23297,N_22875);
and U24560 (N_24560,N_23739,N_23174);
or U24561 (N_24561,N_23415,N_23962);
nor U24562 (N_24562,N_22972,N_23355);
nand U24563 (N_24563,N_23173,N_22757);
xor U24564 (N_24564,N_23444,N_23723);
or U24565 (N_24565,N_23678,N_22756);
nand U24566 (N_24566,N_23490,N_23250);
nand U24567 (N_24567,N_23771,N_23255);
nor U24568 (N_24568,N_22899,N_22663);
or U24569 (N_24569,N_23256,N_22519);
nor U24570 (N_24570,N_22511,N_23071);
nor U24571 (N_24571,N_23115,N_22944);
or U24572 (N_24572,N_22894,N_23780);
and U24573 (N_24573,N_23130,N_22957);
and U24574 (N_24574,N_23110,N_23066);
and U24575 (N_24575,N_23925,N_23216);
and U24576 (N_24576,N_23454,N_23420);
nor U24577 (N_24577,N_22621,N_23184);
nor U24578 (N_24578,N_22993,N_23852);
or U24579 (N_24579,N_23107,N_23422);
xor U24580 (N_24580,N_23936,N_23366);
or U24581 (N_24581,N_23058,N_23972);
or U24582 (N_24582,N_23437,N_23825);
nand U24583 (N_24583,N_23844,N_23478);
nand U24584 (N_24584,N_22646,N_22685);
nand U24585 (N_24585,N_23320,N_23933);
and U24586 (N_24586,N_23984,N_23659);
xor U24587 (N_24587,N_23030,N_23672);
nand U24588 (N_24588,N_23169,N_23327);
nor U24589 (N_24589,N_22584,N_22931);
and U24590 (N_24590,N_23358,N_23035);
nand U24591 (N_24591,N_22793,N_22706);
nor U24592 (N_24592,N_23485,N_22851);
and U24593 (N_24593,N_23920,N_22588);
or U24594 (N_24594,N_23239,N_23913);
nand U24595 (N_24595,N_23241,N_23550);
or U24596 (N_24596,N_23176,N_22721);
or U24597 (N_24597,N_22773,N_22565);
or U24598 (N_24598,N_23094,N_23323);
nand U24599 (N_24599,N_22637,N_23921);
nor U24600 (N_24600,N_22845,N_23306);
or U24601 (N_24601,N_23541,N_23903);
and U24602 (N_24602,N_22662,N_22958);
nor U24603 (N_24603,N_23185,N_22975);
and U24604 (N_24604,N_22548,N_23042);
nand U24605 (N_24605,N_23552,N_23796);
nor U24606 (N_24606,N_23909,N_23155);
nor U24607 (N_24607,N_22587,N_22900);
nor U24608 (N_24608,N_22884,N_23233);
or U24609 (N_24609,N_23910,N_23363);
or U24610 (N_24610,N_23069,N_23700);
and U24611 (N_24611,N_23026,N_23201);
or U24612 (N_24612,N_22602,N_22666);
nor U24613 (N_24613,N_22710,N_22560);
or U24614 (N_24614,N_23457,N_22777);
nand U24615 (N_24615,N_23872,N_23753);
xnor U24616 (N_24616,N_23650,N_23024);
and U24617 (N_24617,N_23015,N_22861);
xor U24618 (N_24618,N_23595,N_22750);
nand U24619 (N_24619,N_23719,N_23828);
nand U24620 (N_24620,N_23767,N_23797);
nand U24621 (N_24621,N_23877,N_23208);
nand U24622 (N_24622,N_22753,N_23960);
nor U24623 (N_24623,N_23362,N_23848);
nor U24624 (N_24624,N_23321,N_23929);
or U24625 (N_24625,N_23213,N_23770);
nand U24626 (N_24626,N_23734,N_23271);
and U24627 (N_24627,N_22941,N_23956);
xnor U24628 (N_24628,N_23125,N_22505);
nand U24629 (N_24629,N_22512,N_23989);
xnor U24630 (N_24630,N_23441,N_23810);
nor U24631 (N_24631,N_22954,N_23513);
xor U24632 (N_24632,N_22932,N_22929);
nand U24633 (N_24633,N_22709,N_22847);
xor U24634 (N_24634,N_23861,N_23781);
or U24635 (N_24635,N_23817,N_22825);
and U24636 (N_24636,N_22724,N_23480);
or U24637 (N_24637,N_22898,N_23894);
nor U24638 (N_24638,N_22707,N_23757);
xor U24639 (N_24639,N_23365,N_22687);
or U24640 (N_24640,N_23649,N_23839);
or U24641 (N_24641,N_23735,N_23521);
nor U24642 (N_24642,N_23018,N_23097);
nor U24643 (N_24643,N_23379,N_22731);
or U24644 (N_24644,N_23548,N_23647);
and U24645 (N_24645,N_22727,N_22980);
nand U24646 (N_24646,N_23452,N_23382);
nand U24647 (N_24647,N_22524,N_23630);
xnor U24648 (N_24648,N_22657,N_23325);
nand U24649 (N_24649,N_23990,N_23985);
and U24650 (N_24650,N_23502,N_23339);
nand U24651 (N_24651,N_23556,N_23514);
nor U24652 (N_24652,N_23102,N_23486);
xnor U24653 (N_24653,N_23146,N_23459);
xnor U24654 (N_24654,N_23165,N_23554);
nor U24655 (N_24655,N_23634,N_22504);
or U24656 (N_24656,N_22956,N_22711);
nor U24657 (N_24657,N_23134,N_23265);
xnor U24658 (N_24658,N_22873,N_23175);
xor U24659 (N_24659,N_22778,N_23281);
or U24660 (N_24660,N_23979,N_23917);
nor U24661 (N_24661,N_23448,N_23761);
nand U24662 (N_24662,N_23242,N_23047);
and U24663 (N_24663,N_23361,N_23442);
or U24664 (N_24664,N_23147,N_23969);
xor U24665 (N_24665,N_23199,N_23328);
nor U24666 (N_24666,N_23372,N_23923);
and U24667 (N_24667,N_23840,N_22945);
and U24668 (N_24668,N_23280,N_23112);
or U24669 (N_24669,N_23995,N_23888);
or U24670 (N_24670,N_23161,N_23319);
nand U24671 (N_24671,N_23027,N_22970);
nor U24672 (N_24672,N_23919,N_23673);
and U24673 (N_24673,N_23160,N_23360);
or U24674 (N_24674,N_22585,N_23456);
and U24675 (N_24675,N_23729,N_23301);
nand U24676 (N_24676,N_23048,N_22763);
nor U24677 (N_24677,N_23871,N_23862);
nand U24678 (N_24678,N_22594,N_23468);
nand U24679 (N_24679,N_22558,N_22914);
xnor U24680 (N_24680,N_23056,N_22834);
or U24681 (N_24681,N_22579,N_23581);
or U24682 (N_24682,N_23787,N_23187);
xor U24683 (N_24683,N_23974,N_22895);
nand U24684 (N_24684,N_23447,N_23032);
nand U24685 (N_24685,N_23748,N_22526);
or U24686 (N_24686,N_23587,N_23768);
nand U24687 (N_24687,N_22586,N_23359);
nor U24688 (N_24688,N_22740,N_22550);
xor U24689 (N_24689,N_23999,N_22921);
nand U24690 (N_24690,N_22682,N_23746);
nor U24691 (N_24691,N_23654,N_23435);
and U24692 (N_24692,N_23284,N_22752);
xnor U24693 (N_24693,N_22693,N_23665);
nand U24694 (N_24694,N_23397,N_23387);
or U24695 (N_24695,N_23702,N_23499);
and U24696 (N_24696,N_22987,N_23471);
nor U24697 (N_24697,N_23059,N_22955);
xnor U24698 (N_24698,N_23377,N_23712);
and U24699 (N_24699,N_22806,N_22543);
nand U24700 (N_24700,N_23795,N_23033);
nor U24701 (N_24701,N_22804,N_23006);
xnor U24702 (N_24702,N_23178,N_23799);
or U24703 (N_24703,N_23257,N_22562);
nand U24704 (N_24704,N_23661,N_23664);
nor U24705 (N_24705,N_23792,N_22784);
nand U24706 (N_24706,N_23668,N_23726);
nor U24707 (N_24707,N_23153,N_23311);
and U24708 (N_24708,N_23980,N_23831);
nor U24709 (N_24709,N_22854,N_22852);
nor U24710 (N_24710,N_22719,N_23758);
nand U24711 (N_24711,N_23551,N_22906);
and U24712 (N_24712,N_23532,N_23192);
nand U24713 (N_24713,N_23641,N_23858);
nand U24714 (N_24714,N_22595,N_22888);
or U24715 (N_24715,N_23622,N_23617);
and U24716 (N_24716,N_23041,N_23429);
xnor U24717 (N_24717,N_23099,N_23274);
nand U24718 (N_24718,N_22575,N_22704);
nor U24719 (N_24719,N_23350,N_23503);
or U24720 (N_24720,N_22689,N_23431);
nor U24721 (N_24721,N_23608,N_23627);
nand U24722 (N_24722,N_23038,N_23338);
or U24723 (N_24723,N_23400,N_22622);
xnor U24724 (N_24724,N_22999,N_23427);
or U24725 (N_24725,N_23911,N_23039);
xor U24726 (N_24726,N_22976,N_23404);
xor U24727 (N_24727,N_22805,N_23314);
or U24728 (N_24728,N_22923,N_22653);
nor U24729 (N_24729,N_23013,N_22578);
xor U24730 (N_24730,N_23512,N_22909);
and U24731 (N_24731,N_22811,N_23234);
nor U24732 (N_24732,N_23992,N_22555);
and U24733 (N_24733,N_23824,N_23500);
nand U24734 (N_24734,N_23040,N_22547);
nor U24735 (N_24735,N_23322,N_22617);
xor U24736 (N_24736,N_23891,N_23167);
nor U24737 (N_24737,N_22998,N_23803);
or U24738 (N_24738,N_23078,N_23607);
nand U24739 (N_24739,N_23524,N_23054);
and U24740 (N_24740,N_23373,N_22770);
xnor U24741 (N_24741,N_23044,N_23728);
nor U24742 (N_24742,N_23043,N_23517);
nand U24743 (N_24743,N_23509,N_22837);
or U24744 (N_24744,N_23663,N_23736);
and U24745 (N_24745,N_23965,N_23682);
or U24746 (N_24746,N_23730,N_23050);
nand U24747 (N_24747,N_23717,N_23177);
or U24748 (N_24748,N_23998,N_22603);
nor U24749 (N_24749,N_23090,N_23836);
xnor U24750 (N_24750,N_23714,N_22663);
xor U24751 (N_24751,N_23395,N_23788);
or U24752 (N_24752,N_23946,N_23473);
and U24753 (N_24753,N_23203,N_23788);
or U24754 (N_24754,N_22998,N_22824);
or U24755 (N_24755,N_23854,N_23029);
and U24756 (N_24756,N_23123,N_23552);
xor U24757 (N_24757,N_22747,N_23238);
and U24758 (N_24758,N_23146,N_23794);
and U24759 (N_24759,N_23535,N_23175);
xnor U24760 (N_24760,N_23106,N_22887);
nand U24761 (N_24761,N_22837,N_22571);
nor U24762 (N_24762,N_22791,N_22960);
xor U24763 (N_24763,N_22742,N_22729);
and U24764 (N_24764,N_22509,N_22600);
nor U24765 (N_24765,N_22913,N_23712);
and U24766 (N_24766,N_23315,N_23968);
nand U24767 (N_24767,N_22883,N_22580);
nand U24768 (N_24768,N_22635,N_23731);
nor U24769 (N_24769,N_23808,N_22937);
nand U24770 (N_24770,N_23395,N_23990);
xor U24771 (N_24771,N_23521,N_23700);
and U24772 (N_24772,N_22765,N_22728);
nand U24773 (N_24773,N_23618,N_23949);
xnor U24774 (N_24774,N_23764,N_23570);
nand U24775 (N_24775,N_23666,N_23126);
and U24776 (N_24776,N_22925,N_23589);
xnor U24777 (N_24777,N_23917,N_23603);
nand U24778 (N_24778,N_23933,N_23884);
xnor U24779 (N_24779,N_23785,N_22540);
nand U24780 (N_24780,N_22915,N_23885);
nand U24781 (N_24781,N_23352,N_23440);
nand U24782 (N_24782,N_23695,N_23832);
nor U24783 (N_24783,N_23255,N_23476);
and U24784 (N_24784,N_23441,N_23499);
xnor U24785 (N_24785,N_23875,N_23055);
nor U24786 (N_24786,N_22869,N_22873);
or U24787 (N_24787,N_23496,N_23003);
or U24788 (N_24788,N_23234,N_23646);
nor U24789 (N_24789,N_22797,N_23968);
xnor U24790 (N_24790,N_22953,N_22856);
or U24791 (N_24791,N_23433,N_23631);
and U24792 (N_24792,N_23605,N_23317);
and U24793 (N_24793,N_22646,N_23098);
xnor U24794 (N_24794,N_23391,N_22511);
nor U24795 (N_24795,N_23015,N_23378);
nand U24796 (N_24796,N_23874,N_23468);
nor U24797 (N_24797,N_23124,N_23617);
nand U24798 (N_24798,N_23993,N_23000);
xor U24799 (N_24799,N_22857,N_22688);
xor U24800 (N_24800,N_23819,N_23010);
or U24801 (N_24801,N_23982,N_23810);
and U24802 (N_24802,N_22714,N_22805);
and U24803 (N_24803,N_23739,N_23592);
and U24804 (N_24804,N_23879,N_23001);
nand U24805 (N_24805,N_23732,N_23316);
or U24806 (N_24806,N_22810,N_22794);
nand U24807 (N_24807,N_23684,N_23788);
nand U24808 (N_24808,N_23652,N_23066);
and U24809 (N_24809,N_22585,N_23613);
and U24810 (N_24810,N_22960,N_23518);
or U24811 (N_24811,N_23154,N_22863);
or U24812 (N_24812,N_23039,N_23487);
and U24813 (N_24813,N_23319,N_23965);
xnor U24814 (N_24814,N_22702,N_22873);
xor U24815 (N_24815,N_23591,N_22924);
or U24816 (N_24816,N_23256,N_22544);
xor U24817 (N_24817,N_22907,N_22788);
or U24818 (N_24818,N_23855,N_23806);
nor U24819 (N_24819,N_22546,N_23611);
or U24820 (N_24820,N_23349,N_22789);
nand U24821 (N_24821,N_22508,N_23811);
nand U24822 (N_24822,N_22999,N_22733);
xor U24823 (N_24823,N_23835,N_23099);
or U24824 (N_24824,N_23775,N_22964);
nor U24825 (N_24825,N_23124,N_22993);
and U24826 (N_24826,N_23004,N_22995);
nor U24827 (N_24827,N_23137,N_23098);
or U24828 (N_24828,N_23675,N_23298);
xor U24829 (N_24829,N_23829,N_23644);
and U24830 (N_24830,N_23205,N_22976);
or U24831 (N_24831,N_23792,N_23920);
nand U24832 (N_24832,N_22557,N_23778);
xor U24833 (N_24833,N_22534,N_23350);
xnor U24834 (N_24834,N_22502,N_22751);
or U24835 (N_24835,N_23861,N_23461);
and U24836 (N_24836,N_23478,N_22829);
xor U24837 (N_24837,N_23224,N_23695);
and U24838 (N_24838,N_22721,N_23172);
xnor U24839 (N_24839,N_22961,N_23122);
nor U24840 (N_24840,N_22774,N_23540);
or U24841 (N_24841,N_23935,N_22567);
and U24842 (N_24842,N_22950,N_23793);
nand U24843 (N_24843,N_22506,N_23912);
nand U24844 (N_24844,N_23384,N_23324);
xor U24845 (N_24845,N_22974,N_22608);
and U24846 (N_24846,N_23818,N_22734);
nor U24847 (N_24847,N_23280,N_22941);
or U24848 (N_24848,N_23999,N_22797);
and U24849 (N_24849,N_23452,N_22646);
and U24850 (N_24850,N_23034,N_23957);
xnor U24851 (N_24851,N_23125,N_23451);
nor U24852 (N_24852,N_23049,N_23644);
and U24853 (N_24853,N_23529,N_22944);
xnor U24854 (N_24854,N_23485,N_23204);
nand U24855 (N_24855,N_23204,N_23816);
xor U24856 (N_24856,N_23768,N_22656);
nor U24857 (N_24857,N_23682,N_23653);
or U24858 (N_24858,N_22530,N_23722);
nor U24859 (N_24859,N_22713,N_23800);
nand U24860 (N_24860,N_22975,N_23152);
and U24861 (N_24861,N_22757,N_22602);
or U24862 (N_24862,N_22889,N_23588);
nor U24863 (N_24863,N_23364,N_23564);
xnor U24864 (N_24864,N_22900,N_23776);
xnor U24865 (N_24865,N_23701,N_23399);
nand U24866 (N_24866,N_22927,N_23244);
and U24867 (N_24867,N_23249,N_23536);
and U24868 (N_24868,N_22795,N_23771);
or U24869 (N_24869,N_23614,N_23071);
nor U24870 (N_24870,N_23414,N_23563);
nor U24871 (N_24871,N_23859,N_23255);
xnor U24872 (N_24872,N_23369,N_23359);
xnor U24873 (N_24873,N_23717,N_23720);
nand U24874 (N_24874,N_23809,N_23877);
nand U24875 (N_24875,N_23881,N_22955);
and U24876 (N_24876,N_23122,N_22635);
nand U24877 (N_24877,N_23347,N_23776);
nand U24878 (N_24878,N_23481,N_23917);
nand U24879 (N_24879,N_23197,N_23909);
xnor U24880 (N_24880,N_22597,N_22533);
xor U24881 (N_24881,N_23995,N_23761);
and U24882 (N_24882,N_23390,N_22656);
nor U24883 (N_24883,N_22565,N_22794);
and U24884 (N_24884,N_23123,N_23467);
nor U24885 (N_24885,N_23160,N_22840);
or U24886 (N_24886,N_23241,N_23946);
xnor U24887 (N_24887,N_22558,N_22508);
nand U24888 (N_24888,N_23895,N_23457);
xor U24889 (N_24889,N_23335,N_22920);
xor U24890 (N_24890,N_23219,N_23178);
or U24891 (N_24891,N_23844,N_23949);
xor U24892 (N_24892,N_22946,N_23511);
nand U24893 (N_24893,N_23225,N_23220);
or U24894 (N_24894,N_23798,N_22930);
xor U24895 (N_24895,N_22896,N_23740);
nor U24896 (N_24896,N_23567,N_23830);
xor U24897 (N_24897,N_23075,N_23433);
nand U24898 (N_24898,N_23462,N_23398);
and U24899 (N_24899,N_23964,N_23097);
nand U24900 (N_24900,N_23391,N_22968);
or U24901 (N_24901,N_23100,N_23367);
xnor U24902 (N_24902,N_23557,N_22711);
or U24903 (N_24903,N_22574,N_22892);
nand U24904 (N_24904,N_23150,N_22640);
and U24905 (N_24905,N_23592,N_23832);
and U24906 (N_24906,N_23609,N_23004);
nand U24907 (N_24907,N_22895,N_22577);
nor U24908 (N_24908,N_23818,N_23522);
xnor U24909 (N_24909,N_22791,N_23138);
nand U24910 (N_24910,N_22750,N_23040);
or U24911 (N_24911,N_23893,N_23295);
xnor U24912 (N_24912,N_23670,N_23010);
nand U24913 (N_24913,N_23454,N_23191);
and U24914 (N_24914,N_22797,N_22866);
xnor U24915 (N_24915,N_22716,N_22586);
or U24916 (N_24916,N_23577,N_23761);
or U24917 (N_24917,N_23450,N_23188);
nor U24918 (N_24918,N_23624,N_23139);
nor U24919 (N_24919,N_23924,N_23921);
xnor U24920 (N_24920,N_23868,N_23591);
nand U24921 (N_24921,N_23152,N_22999);
xor U24922 (N_24922,N_23928,N_22900);
nand U24923 (N_24923,N_22742,N_22653);
xor U24924 (N_24924,N_23915,N_23397);
and U24925 (N_24925,N_23505,N_23007);
nand U24926 (N_24926,N_23184,N_23087);
or U24927 (N_24927,N_23827,N_23825);
nand U24928 (N_24928,N_23288,N_23175);
nand U24929 (N_24929,N_23292,N_22802);
and U24930 (N_24930,N_23250,N_23995);
nor U24931 (N_24931,N_22704,N_22955);
xnor U24932 (N_24932,N_22526,N_23509);
nand U24933 (N_24933,N_23533,N_23589);
nand U24934 (N_24934,N_22835,N_22564);
nand U24935 (N_24935,N_22617,N_22928);
or U24936 (N_24936,N_23087,N_23961);
nand U24937 (N_24937,N_22535,N_22509);
nor U24938 (N_24938,N_22886,N_23649);
nand U24939 (N_24939,N_22950,N_22937);
xnor U24940 (N_24940,N_23203,N_23748);
xor U24941 (N_24941,N_23377,N_23008);
nand U24942 (N_24942,N_23967,N_23090);
and U24943 (N_24943,N_22936,N_23102);
and U24944 (N_24944,N_23270,N_23559);
xnor U24945 (N_24945,N_23232,N_23668);
nand U24946 (N_24946,N_22712,N_23357);
xor U24947 (N_24947,N_23594,N_23537);
or U24948 (N_24948,N_22631,N_23854);
nor U24949 (N_24949,N_22525,N_22573);
nand U24950 (N_24950,N_23511,N_22670);
nand U24951 (N_24951,N_23214,N_23347);
nor U24952 (N_24952,N_22826,N_22774);
xor U24953 (N_24953,N_23347,N_22861);
nor U24954 (N_24954,N_23855,N_23158);
and U24955 (N_24955,N_23591,N_22831);
xor U24956 (N_24956,N_23510,N_23945);
and U24957 (N_24957,N_23687,N_23011);
or U24958 (N_24958,N_22592,N_23574);
xnor U24959 (N_24959,N_23572,N_23436);
nor U24960 (N_24960,N_22739,N_22589);
nand U24961 (N_24961,N_23933,N_23292);
and U24962 (N_24962,N_23908,N_23965);
or U24963 (N_24963,N_22973,N_23692);
and U24964 (N_24964,N_23173,N_23515);
nor U24965 (N_24965,N_23394,N_23443);
nor U24966 (N_24966,N_23374,N_22537);
xor U24967 (N_24967,N_23152,N_22826);
nand U24968 (N_24968,N_23440,N_22624);
nand U24969 (N_24969,N_23367,N_23611);
or U24970 (N_24970,N_23521,N_22808);
and U24971 (N_24971,N_23612,N_22558);
xnor U24972 (N_24972,N_23001,N_22897);
nand U24973 (N_24973,N_23270,N_22822);
and U24974 (N_24974,N_22769,N_23717);
nor U24975 (N_24975,N_23749,N_23335);
and U24976 (N_24976,N_23371,N_22503);
and U24977 (N_24977,N_22666,N_23696);
or U24978 (N_24978,N_22543,N_23130);
xor U24979 (N_24979,N_22920,N_22940);
nor U24980 (N_24980,N_22996,N_23852);
and U24981 (N_24981,N_22672,N_22932);
xor U24982 (N_24982,N_23753,N_22576);
nor U24983 (N_24983,N_22964,N_23157);
xnor U24984 (N_24984,N_23805,N_23205);
nor U24985 (N_24985,N_23182,N_23190);
xor U24986 (N_24986,N_22543,N_23885);
xnor U24987 (N_24987,N_22579,N_23348);
or U24988 (N_24988,N_23854,N_23537);
or U24989 (N_24989,N_23864,N_23654);
xor U24990 (N_24990,N_23714,N_23483);
and U24991 (N_24991,N_23766,N_22559);
nor U24992 (N_24992,N_22821,N_22832);
and U24993 (N_24993,N_23678,N_22868);
xor U24994 (N_24994,N_23274,N_23610);
nand U24995 (N_24995,N_23860,N_22534);
and U24996 (N_24996,N_23895,N_22980);
and U24997 (N_24997,N_22507,N_22910);
xor U24998 (N_24998,N_23505,N_23726);
nor U24999 (N_24999,N_23973,N_23069);
xor U25000 (N_25000,N_22713,N_23856);
or U25001 (N_25001,N_22867,N_22875);
nand U25002 (N_25002,N_23978,N_23910);
and U25003 (N_25003,N_23263,N_22575);
nor U25004 (N_25004,N_23450,N_23643);
nand U25005 (N_25005,N_23535,N_22843);
or U25006 (N_25006,N_23297,N_23280);
nor U25007 (N_25007,N_23668,N_23296);
nand U25008 (N_25008,N_23307,N_23782);
and U25009 (N_25009,N_22672,N_22575);
and U25010 (N_25010,N_23322,N_22629);
nor U25011 (N_25011,N_22815,N_23641);
xor U25012 (N_25012,N_23594,N_23374);
and U25013 (N_25013,N_23260,N_22580);
or U25014 (N_25014,N_23987,N_23102);
nor U25015 (N_25015,N_22929,N_23709);
xnor U25016 (N_25016,N_22677,N_23468);
nor U25017 (N_25017,N_23297,N_23660);
nor U25018 (N_25018,N_23221,N_22718);
nand U25019 (N_25019,N_23656,N_23629);
and U25020 (N_25020,N_23292,N_23703);
xnor U25021 (N_25021,N_23688,N_23203);
xor U25022 (N_25022,N_22905,N_23887);
nor U25023 (N_25023,N_23063,N_23655);
or U25024 (N_25024,N_23405,N_22629);
nor U25025 (N_25025,N_23140,N_23891);
nor U25026 (N_25026,N_23532,N_23913);
and U25027 (N_25027,N_23531,N_23006);
xor U25028 (N_25028,N_22584,N_22917);
and U25029 (N_25029,N_23754,N_23175);
and U25030 (N_25030,N_23182,N_23409);
and U25031 (N_25031,N_23138,N_23560);
nor U25032 (N_25032,N_22585,N_23466);
nor U25033 (N_25033,N_23233,N_23083);
and U25034 (N_25034,N_23038,N_22546);
or U25035 (N_25035,N_22722,N_23035);
nand U25036 (N_25036,N_23714,N_23249);
xnor U25037 (N_25037,N_23616,N_22769);
nand U25038 (N_25038,N_23971,N_23463);
xnor U25039 (N_25039,N_23119,N_22922);
nor U25040 (N_25040,N_22889,N_23403);
or U25041 (N_25041,N_23391,N_22927);
or U25042 (N_25042,N_22807,N_23285);
nand U25043 (N_25043,N_22558,N_22594);
nand U25044 (N_25044,N_22596,N_22900);
or U25045 (N_25045,N_22686,N_23739);
nand U25046 (N_25046,N_23994,N_23419);
nor U25047 (N_25047,N_22977,N_23508);
and U25048 (N_25048,N_23836,N_23670);
and U25049 (N_25049,N_23691,N_22985);
nand U25050 (N_25050,N_23994,N_23022);
nand U25051 (N_25051,N_22635,N_23791);
nor U25052 (N_25052,N_23569,N_22571);
and U25053 (N_25053,N_22984,N_23999);
nor U25054 (N_25054,N_23861,N_22742);
or U25055 (N_25055,N_23983,N_23640);
nor U25056 (N_25056,N_22626,N_23409);
nor U25057 (N_25057,N_23131,N_22923);
nor U25058 (N_25058,N_23266,N_23855);
xor U25059 (N_25059,N_22684,N_23476);
or U25060 (N_25060,N_23904,N_23639);
and U25061 (N_25061,N_23026,N_23304);
xor U25062 (N_25062,N_23075,N_23897);
or U25063 (N_25063,N_22569,N_22538);
nor U25064 (N_25064,N_23848,N_23344);
nor U25065 (N_25065,N_22912,N_23607);
nor U25066 (N_25066,N_22775,N_23739);
or U25067 (N_25067,N_23376,N_23808);
or U25068 (N_25068,N_22962,N_23725);
xnor U25069 (N_25069,N_23728,N_23893);
xor U25070 (N_25070,N_23102,N_22877);
nor U25071 (N_25071,N_22742,N_22916);
nand U25072 (N_25072,N_23561,N_23365);
or U25073 (N_25073,N_23798,N_22608);
and U25074 (N_25074,N_22562,N_23081);
nor U25075 (N_25075,N_23727,N_23978);
and U25076 (N_25076,N_22856,N_22893);
nor U25077 (N_25077,N_23315,N_23673);
xor U25078 (N_25078,N_22944,N_23020);
nand U25079 (N_25079,N_23098,N_23162);
or U25080 (N_25080,N_23889,N_23667);
xnor U25081 (N_25081,N_22877,N_22714);
nor U25082 (N_25082,N_23307,N_23196);
and U25083 (N_25083,N_23701,N_23891);
or U25084 (N_25084,N_23555,N_23876);
or U25085 (N_25085,N_23035,N_22739);
nand U25086 (N_25086,N_23417,N_22664);
nor U25087 (N_25087,N_22720,N_23849);
or U25088 (N_25088,N_22827,N_22819);
nor U25089 (N_25089,N_23334,N_23236);
nor U25090 (N_25090,N_23219,N_23994);
nand U25091 (N_25091,N_23773,N_23939);
nand U25092 (N_25092,N_23000,N_23439);
and U25093 (N_25093,N_22774,N_22981);
or U25094 (N_25094,N_23637,N_22793);
nand U25095 (N_25095,N_23965,N_22631);
nor U25096 (N_25096,N_23664,N_23976);
xor U25097 (N_25097,N_22973,N_23066);
nand U25098 (N_25098,N_23088,N_23944);
xor U25099 (N_25099,N_22796,N_23450);
nor U25100 (N_25100,N_22934,N_23306);
and U25101 (N_25101,N_23289,N_22734);
and U25102 (N_25102,N_22530,N_22686);
xor U25103 (N_25103,N_23363,N_23773);
and U25104 (N_25104,N_22869,N_23720);
nand U25105 (N_25105,N_22633,N_23477);
xor U25106 (N_25106,N_23551,N_23044);
or U25107 (N_25107,N_23008,N_23158);
xnor U25108 (N_25108,N_23398,N_23758);
or U25109 (N_25109,N_23237,N_23122);
and U25110 (N_25110,N_23166,N_22796);
or U25111 (N_25111,N_22886,N_22608);
and U25112 (N_25112,N_22638,N_23828);
nor U25113 (N_25113,N_23897,N_23664);
nand U25114 (N_25114,N_22970,N_22996);
nand U25115 (N_25115,N_22701,N_23401);
and U25116 (N_25116,N_22862,N_22531);
xor U25117 (N_25117,N_23335,N_23183);
nand U25118 (N_25118,N_23947,N_23378);
nor U25119 (N_25119,N_22856,N_22584);
or U25120 (N_25120,N_22525,N_22617);
or U25121 (N_25121,N_22963,N_22940);
nand U25122 (N_25122,N_23603,N_22666);
and U25123 (N_25123,N_23897,N_23461);
and U25124 (N_25124,N_22769,N_23894);
nand U25125 (N_25125,N_23773,N_23657);
or U25126 (N_25126,N_23118,N_23877);
and U25127 (N_25127,N_23734,N_23547);
nand U25128 (N_25128,N_23904,N_23715);
xnor U25129 (N_25129,N_22665,N_22948);
or U25130 (N_25130,N_22828,N_23333);
and U25131 (N_25131,N_23942,N_22511);
or U25132 (N_25132,N_23125,N_23392);
or U25133 (N_25133,N_23056,N_22583);
nand U25134 (N_25134,N_23211,N_23238);
or U25135 (N_25135,N_23003,N_22516);
and U25136 (N_25136,N_23508,N_22833);
and U25137 (N_25137,N_23544,N_23726);
nand U25138 (N_25138,N_23881,N_22943);
nand U25139 (N_25139,N_23028,N_22755);
or U25140 (N_25140,N_22595,N_23868);
xnor U25141 (N_25141,N_23733,N_23523);
and U25142 (N_25142,N_23171,N_23729);
nor U25143 (N_25143,N_23637,N_23037);
nor U25144 (N_25144,N_22853,N_22522);
nand U25145 (N_25145,N_23886,N_23517);
nand U25146 (N_25146,N_23827,N_23136);
nand U25147 (N_25147,N_22673,N_22895);
nor U25148 (N_25148,N_23740,N_23925);
nor U25149 (N_25149,N_23638,N_23038);
nor U25150 (N_25150,N_22749,N_23003);
nand U25151 (N_25151,N_22797,N_22815);
xnor U25152 (N_25152,N_23224,N_23427);
nor U25153 (N_25153,N_23587,N_23859);
or U25154 (N_25154,N_22976,N_23954);
nand U25155 (N_25155,N_23248,N_22639);
or U25156 (N_25156,N_22783,N_22507);
or U25157 (N_25157,N_22677,N_23042);
xnor U25158 (N_25158,N_23305,N_23337);
and U25159 (N_25159,N_22906,N_23834);
or U25160 (N_25160,N_23107,N_22509);
or U25161 (N_25161,N_23337,N_22554);
nor U25162 (N_25162,N_23221,N_23126);
nor U25163 (N_25163,N_23440,N_23381);
or U25164 (N_25164,N_23716,N_23201);
xnor U25165 (N_25165,N_23901,N_23561);
or U25166 (N_25166,N_23367,N_22639);
and U25167 (N_25167,N_23834,N_23201);
xor U25168 (N_25168,N_23915,N_22548);
or U25169 (N_25169,N_23870,N_22797);
nor U25170 (N_25170,N_23431,N_22589);
nand U25171 (N_25171,N_23279,N_23666);
nand U25172 (N_25172,N_22829,N_22842);
xnor U25173 (N_25173,N_23101,N_23625);
nand U25174 (N_25174,N_23484,N_23308);
nand U25175 (N_25175,N_23258,N_22858);
xnor U25176 (N_25176,N_23324,N_22784);
or U25177 (N_25177,N_23295,N_23911);
xnor U25178 (N_25178,N_22996,N_22559);
nor U25179 (N_25179,N_22620,N_22801);
or U25180 (N_25180,N_22748,N_23939);
xor U25181 (N_25181,N_23318,N_22954);
nand U25182 (N_25182,N_23719,N_22664);
xnor U25183 (N_25183,N_22745,N_23788);
nor U25184 (N_25184,N_23677,N_23221);
nor U25185 (N_25185,N_23677,N_22720);
nand U25186 (N_25186,N_22511,N_23727);
or U25187 (N_25187,N_23695,N_23072);
xor U25188 (N_25188,N_22787,N_23550);
and U25189 (N_25189,N_23942,N_23308);
nor U25190 (N_25190,N_22987,N_22986);
and U25191 (N_25191,N_22692,N_23963);
nand U25192 (N_25192,N_23653,N_23503);
and U25193 (N_25193,N_23455,N_22675);
or U25194 (N_25194,N_23523,N_23921);
nor U25195 (N_25195,N_22921,N_23833);
nand U25196 (N_25196,N_23084,N_22931);
or U25197 (N_25197,N_22677,N_23370);
nand U25198 (N_25198,N_23087,N_23016);
nand U25199 (N_25199,N_23598,N_22739);
or U25200 (N_25200,N_22970,N_22628);
nand U25201 (N_25201,N_22601,N_22768);
xor U25202 (N_25202,N_22930,N_22687);
nor U25203 (N_25203,N_23749,N_22761);
and U25204 (N_25204,N_22923,N_22875);
and U25205 (N_25205,N_23552,N_22545);
nor U25206 (N_25206,N_23967,N_22560);
nor U25207 (N_25207,N_23377,N_23600);
nand U25208 (N_25208,N_23317,N_22673);
nand U25209 (N_25209,N_23498,N_23867);
or U25210 (N_25210,N_23862,N_23037);
xor U25211 (N_25211,N_23235,N_23939);
and U25212 (N_25212,N_22849,N_23884);
nor U25213 (N_25213,N_23115,N_23196);
nand U25214 (N_25214,N_23887,N_23292);
nor U25215 (N_25215,N_23583,N_22669);
nand U25216 (N_25216,N_23995,N_23180);
and U25217 (N_25217,N_23272,N_23753);
nand U25218 (N_25218,N_22921,N_23338);
xnor U25219 (N_25219,N_22941,N_23819);
nor U25220 (N_25220,N_23995,N_23666);
xnor U25221 (N_25221,N_22835,N_23961);
nand U25222 (N_25222,N_23190,N_22827);
xor U25223 (N_25223,N_22776,N_23091);
xor U25224 (N_25224,N_23429,N_23288);
xnor U25225 (N_25225,N_23078,N_23643);
or U25226 (N_25226,N_23630,N_23945);
nand U25227 (N_25227,N_23097,N_23546);
and U25228 (N_25228,N_23904,N_23690);
nand U25229 (N_25229,N_22814,N_22863);
xor U25230 (N_25230,N_23803,N_22635);
xor U25231 (N_25231,N_23331,N_23242);
nand U25232 (N_25232,N_22898,N_23133);
or U25233 (N_25233,N_22986,N_23077);
nor U25234 (N_25234,N_22514,N_23491);
or U25235 (N_25235,N_23203,N_23626);
and U25236 (N_25236,N_23655,N_23041);
nor U25237 (N_25237,N_23925,N_23241);
or U25238 (N_25238,N_23627,N_23605);
nand U25239 (N_25239,N_23678,N_22542);
and U25240 (N_25240,N_23948,N_23144);
or U25241 (N_25241,N_23131,N_22730);
nor U25242 (N_25242,N_22679,N_23515);
and U25243 (N_25243,N_22614,N_23582);
or U25244 (N_25244,N_23486,N_23876);
xor U25245 (N_25245,N_23591,N_22818);
or U25246 (N_25246,N_23578,N_23079);
nor U25247 (N_25247,N_23477,N_23901);
and U25248 (N_25248,N_22545,N_23618);
or U25249 (N_25249,N_23964,N_22767);
nor U25250 (N_25250,N_23169,N_23925);
nand U25251 (N_25251,N_22686,N_23652);
nand U25252 (N_25252,N_22842,N_22881);
nand U25253 (N_25253,N_23434,N_22521);
nor U25254 (N_25254,N_23597,N_22806);
nand U25255 (N_25255,N_23381,N_23156);
or U25256 (N_25256,N_22680,N_23215);
or U25257 (N_25257,N_22740,N_23947);
or U25258 (N_25258,N_22613,N_22627);
nor U25259 (N_25259,N_23647,N_23479);
nor U25260 (N_25260,N_23403,N_23831);
nand U25261 (N_25261,N_22675,N_23087);
nor U25262 (N_25262,N_22776,N_23144);
xor U25263 (N_25263,N_23462,N_23671);
and U25264 (N_25264,N_23576,N_22690);
nand U25265 (N_25265,N_23559,N_23457);
xnor U25266 (N_25266,N_22942,N_23978);
or U25267 (N_25267,N_23787,N_22995);
and U25268 (N_25268,N_22955,N_23893);
xor U25269 (N_25269,N_22565,N_22975);
nor U25270 (N_25270,N_23886,N_22615);
nor U25271 (N_25271,N_22972,N_23089);
nor U25272 (N_25272,N_23847,N_22971);
nor U25273 (N_25273,N_23984,N_22542);
and U25274 (N_25274,N_22511,N_22932);
and U25275 (N_25275,N_23408,N_22927);
xnor U25276 (N_25276,N_23632,N_23225);
xnor U25277 (N_25277,N_23321,N_23233);
nand U25278 (N_25278,N_23802,N_22713);
and U25279 (N_25279,N_23580,N_22533);
and U25280 (N_25280,N_22925,N_23518);
xor U25281 (N_25281,N_23831,N_23603);
or U25282 (N_25282,N_23972,N_23033);
or U25283 (N_25283,N_23767,N_22797);
and U25284 (N_25284,N_22755,N_22756);
nor U25285 (N_25285,N_22611,N_22664);
nor U25286 (N_25286,N_22787,N_23991);
nor U25287 (N_25287,N_23853,N_23955);
and U25288 (N_25288,N_23690,N_23168);
nand U25289 (N_25289,N_22956,N_22594);
nand U25290 (N_25290,N_23196,N_22958);
or U25291 (N_25291,N_23677,N_23857);
nand U25292 (N_25292,N_23547,N_23900);
xor U25293 (N_25293,N_22806,N_22628);
nor U25294 (N_25294,N_23519,N_23708);
and U25295 (N_25295,N_23867,N_23057);
nand U25296 (N_25296,N_22587,N_23685);
nand U25297 (N_25297,N_22557,N_23379);
xor U25298 (N_25298,N_23739,N_23871);
nor U25299 (N_25299,N_23781,N_23687);
nand U25300 (N_25300,N_23437,N_23649);
or U25301 (N_25301,N_23807,N_22604);
nand U25302 (N_25302,N_23938,N_22768);
nor U25303 (N_25303,N_22523,N_22545);
and U25304 (N_25304,N_22648,N_23353);
or U25305 (N_25305,N_22716,N_23968);
nand U25306 (N_25306,N_23890,N_22809);
xor U25307 (N_25307,N_23816,N_23845);
xor U25308 (N_25308,N_22548,N_23743);
and U25309 (N_25309,N_23189,N_23645);
xnor U25310 (N_25310,N_23300,N_22986);
nand U25311 (N_25311,N_23765,N_23645);
nand U25312 (N_25312,N_22956,N_23932);
nor U25313 (N_25313,N_23335,N_22649);
nor U25314 (N_25314,N_22616,N_23806);
nand U25315 (N_25315,N_23689,N_22735);
and U25316 (N_25316,N_22661,N_23901);
nor U25317 (N_25317,N_22969,N_23416);
nand U25318 (N_25318,N_23274,N_23511);
nor U25319 (N_25319,N_22926,N_22707);
and U25320 (N_25320,N_22925,N_23927);
nand U25321 (N_25321,N_23125,N_22727);
or U25322 (N_25322,N_22634,N_22724);
or U25323 (N_25323,N_23211,N_23070);
nand U25324 (N_25324,N_22527,N_23673);
nand U25325 (N_25325,N_23683,N_23684);
xnor U25326 (N_25326,N_23577,N_22717);
or U25327 (N_25327,N_23622,N_23832);
nand U25328 (N_25328,N_22529,N_23141);
or U25329 (N_25329,N_22527,N_23475);
nor U25330 (N_25330,N_22909,N_23839);
xor U25331 (N_25331,N_23494,N_23602);
nand U25332 (N_25332,N_22547,N_22574);
xnor U25333 (N_25333,N_22729,N_23604);
xor U25334 (N_25334,N_23494,N_23666);
nor U25335 (N_25335,N_23191,N_22584);
and U25336 (N_25336,N_23031,N_23815);
or U25337 (N_25337,N_22602,N_23118);
nor U25338 (N_25338,N_23523,N_22617);
nand U25339 (N_25339,N_22705,N_23403);
or U25340 (N_25340,N_22941,N_23634);
or U25341 (N_25341,N_22506,N_22742);
and U25342 (N_25342,N_22910,N_23663);
nor U25343 (N_25343,N_23463,N_23721);
nor U25344 (N_25344,N_23532,N_22748);
nor U25345 (N_25345,N_23260,N_23277);
nor U25346 (N_25346,N_23187,N_23267);
or U25347 (N_25347,N_22652,N_22552);
or U25348 (N_25348,N_23527,N_22881);
and U25349 (N_25349,N_22904,N_23514);
xnor U25350 (N_25350,N_22827,N_23982);
xnor U25351 (N_25351,N_22968,N_22766);
xor U25352 (N_25352,N_23692,N_23793);
nand U25353 (N_25353,N_23812,N_23709);
nand U25354 (N_25354,N_23446,N_22948);
nand U25355 (N_25355,N_23650,N_23795);
nand U25356 (N_25356,N_23533,N_22898);
or U25357 (N_25357,N_23724,N_23302);
and U25358 (N_25358,N_22731,N_23024);
or U25359 (N_25359,N_22709,N_22581);
nand U25360 (N_25360,N_22680,N_23484);
xor U25361 (N_25361,N_23911,N_23721);
nand U25362 (N_25362,N_22669,N_22955);
and U25363 (N_25363,N_22670,N_22754);
or U25364 (N_25364,N_23654,N_23123);
nor U25365 (N_25365,N_23134,N_23188);
nand U25366 (N_25366,N_22818,N_23351);
or U25367 (N_25367,N_23756,N_23939);
xor U25368 (N_25368,N_22990,N_23108);
nand U25369 (N_25369,N_22559,N_23503);
nor U25370 (N_25370,N_23063,N_23966);
or U25371 (N_25371,N_23661,N_23414);
nand U25372 (N_25372,N_22892,N_23330);
and U25373 (N_25373,N_22966,N_22524);
and U25374 (N_25374,N_22880,N_22580);
xnor U25375 (N_25375,N_23467,N_22708);
or U25376 (N_25376,N_22573,N_22837);
nor U25377 (N_25377,N_23920,N_23554);
and U25378 (N_25378,N_22877,N_23412);
nor U25379 (N_25379,N_23960,N_22972);
xnor U25380 (N_25380,N_22646,N_22767);
nor U25381 (N_25381,N_22775,N_23805);
nand U25382 (N_25382,N_23202,N_22974);
nand U25383 (N_25383,N_23465,N_22627);
or U25384 (N_25384,N_23317,N_23225);
xor U25385 (N_25385,N_23290,N_23568);
xor U25386 (N_25386,N_23092,N_22958);
or U25387 (N_25387,N_22655,N_23312);
and U25388 (N_25388,N_22761,N_22987);
and U25389 (N_25389,N_22518,N_22897);
or U25390 (N_25390,N_23259,N_23356);
nor U25391 (N_25391,N_23654,N_22775);
nor U25392 (N_25392,N_23849,N_23374);
xor U25393 (N_25393,N_22799,N_23059);
and U25394 (N_25394,N_23725,N_22507);
nor U25395 (N_25395,N_23534,N_22577);
xor U25396 (N_25396,N_22669,N_23639);
nand U25397 (N_25397,N_22724,N_23902);
and U25398 (N_25398,N_22952,N_23320);
nor U25399 (N_25399,N_23186,N_23820);
xor U25400 (N_25400,N_22528,N_23234);
nand U25401 (N_25401,N_22681,N_23397);
or U25402 (N_25402,N_23961,N_22897);
or U25403 (N_25403,N_22642,N_22639);
nor U25404 (N_25404,N_22953,N_23489);
or U25405 (N_25405,N_23989,N_22874);
nand U25406 (N_25406,N_22909,N_22877);
nand U25407 (N_25407,N_23998,N_23854);
or U25408 (N_25408,N_23819,N_22840);
and U25409 (N_25409,N_22973,N_23029);
nor U25410 (N_25410,N_22961,N_23487);
xor U25411 (N_25411,N_23456,N_23987);
and U25412 (N_25412,N_22830,N_22944);
or U25413 (N_25413,N_23730,N_23161);
nand U25414 (N_25414,N_23131,N_23783);
and U25415 (N_25415,N_22840,N_23298);
and U25416 (N_25416,N_23086,N_22986);
or U25417 (N_25417,N_23851,N_23923);
nand U25418 (N_25418,N_23982,N_22531);
nor U25419 (N_25419,N_22934,N_22841);
or U25420 (N_25420,N_23122,N_23750);
nor U25421 (N_25421,N_23701,N_23824);
xnor U25422 (N_25422,N_23162,N_23537);
and U25423 (N_25423,N_22516,N_22843);
or U25424 (N_25424,N_23977,N_22911);
or U25425 (N_25425,N_23719,N_22746);
and U25426 (N_25426,N_22689,N_23895);
nand U25427 (N_25427,N_22795,N_22675);
xnor U25428 (N_25428,N_23817,N_23610);
nor U25429 (N_25429,N_22567,N_23930);
xnor U25430 (N_25430,N_22789,N_22632);
and U25431 (N_25431,N_23802,N_22536);
or U25432 (N_25432,N_22688,N_23565);
or U25433 (N_25433,N_23801,N_23363);
and U25434 (N_25434,N_23790,N_22721);
or U25435 (N_25435,N_23956,N_22668);
and U25436 (N_25436,N_23673,N_23539);
nand U25437 (N_25437,N_23911,N_23873);
and U25438 (N_25438,N_23382,N_23934);
nor U25439 (N_25439,N_22627,N_23555);
nand U25440 (N_25440,N_23180,N_22856);
xor U25441 (N_25441,N_23126,N_22831);
and U25442 (N_25442,N_22901,N_22643);
or U25443 (N_25443,N_22988,N_22806);
or U25444 (N_25444,N_23585,N_22539);
nor U25445 (N_25445,N_23009,N_23227);
or U25446 (N_25446,N_22721,N_23512);
and U25447 (N_25447,N_23202,N_23828);
or U25448 (N_25448,N_23229,N_23082);
or U25449 (N_25449,N_22583,N_22971);
or U25450 (N_25450,N_23266,N_22717);
and U25451 (N_25451,N_22927,N_22679);
and U25452 (N_25452,N_23614,N_23294);
nor U25453 (N_25453,N_22984,N_22849);
and U25454 (N_25454,N_22685,N_23652);
and U25455 (N_25455,N_22750,N_23786);
nand U25456 (N_25456,N_23705,N_23684);
and U25457 (N_25457,N_22782,N_23265);
nand U25458 (N_25458,N_23585,N_22846);
and U25459 (N_25459,N_22576,N_22685);
or U25460 (N_25460,N_23450,N_23163);
xor U25461 (N_25461,N_23984,N_23219);
and U25462 (N_25462,N_22857,N_23996);
nor U25463 (N_25463,N_23653,N_23860);
and U25464 (N_25464,N_23812,N_22755);
or U25465 (N_25465,N_23349,N_23549);
xor U25466 (N_25466,N_22873,N_23509);
and U25467 (N_25467,N_22928,N_22740);
nand U25468 (N_25468,N_22619,N_22776);
nor U25469 (N_25469,N_23933,N_23555);
and U25470 (N_25470,N_23977,N_22646);
xnor U25471 (N_25471,N_23782,N_23141);
nand U25472 (N_25472,N_22731,N_23946);
nand U25473 (N_25473,N_23487,N_23646);
and U25474 (N_25474,N_23712,N_23397);
xor U25475 (N_25475,N_22749,N_23553);
xor U25476 (N_25476,N_23934,N_23544);
and U25477 (N_25477,N_22995,N_23250);
or U25478 (N_25478,N_23706,N_23198);
nand U25479 (N_25479,N_23695,N_22500);
nand U25480 (N_25480,N_23497,N_23824);
nand U25481 (N_25481,N_22737,N_23239);
and U25482 (N_25482,N_22767,N_23229);
nand U25483 (N_25483,N_22561,N_22550);
or U25484 (N_25484,N_23796,N_23132);
nand U25485 (N_25485,N_23166,N_23792);
xnor U25486 (N_25486,N_23725,N_22503);
or U25487 (N_25487,N_23629,N_23517);
and U25488 (N_25488,N_23375,N_22703);
and U25489 (N_25489,N_23926,N_23913);
nand U25490 (N_25490,N_23942,N_23887);
nand U25491 (N_25491,N_23120,N_22925);
and U25492 (N_25492,N_23336,N_22601);
nand U25493 (N_25493,N_23465,N_22749);
nor U25494 (N_25494,N_23554,N_23769);
xor U25495 (N_25495,N_23178,N_23460);
nand U25496 (N_25496,N_22875,N_23806);
and U25497 (N_25497,N_23274,N_23100);
nor U25498 (N_25498,N_23633,N_23844);
xnor U25499 (N_25499,N_23235,N_22817);
and U25500 (N_25500,N_25203,N_24571);
or U25501 (N_25501,N_24802,N_25280);
nand U25502 (N_25502,N_24504,N_25436);
and U25503 (N_25503,N_24039,N_25062);
nor U25504 (N_25504,N_25355,N_25098);
and U25505 (N_25505,N_25399,N_24219);
or U25506 (N_25506,N_24756,N_24115);
xnor U25507 (N_25507,N_25193,N_25104);
or U25508 (N_25508,N_24528,N_24805);
xnor U25509 (N_25509,N_24598,N_25414);
and U25510 (N_25510,N_24468,N_24263);
nor U25511 (N_25511,N_24976,N_24878);
or U25512 (N_25512,N_24070,N_24259);
xor U25513 (N_25513,N_24635,N_24673);
nor U25514 (N_25514,N_25151,N_24617);
and U25515 (N_25515,N_25293,N_24602);
or U25516 (N_25516,N_24241,N_24315);
nand U25517 (N_25517,N_25069,N_24725);
or U25518 (N_25518,N_24205,N_24909);
nor U25519 (N_25519,N_24233,N_25469);
and U25520 (N_25520,N_24535,N_24652);
or U25521 (N_25521,N_24511,N_25157);
nand U25522 (N_25522,N_24587,N_24250);
and U25523 (N_25523,N_25146,N_25400);
xor U25524 (N_25524,N_24564,N_25457);
and U25525 (N_25525,N_24732,N_24918);
nor U25526 (N_25526,N_24236,N_25106);
nor U25527 (N_25527,N_25370,N_24414);
nor U25528 (N_25528,N_25264,N_24765);
xor U25529 (N_25529,N_24611,N_24033);
and U25530 (N_25530,N_25216,N_25390);
nand U25531 (N_25531,N_24580,N_24268);
nor U25532 (N_25532,N_24684,N_24514);
nand U25533 (N_25533,N_24405,N_25415);
xnor U25534 (N_25534,N_24006,N_24188);
or U25535 (N_25535,N_25347,N_24620);
or U25536 (N_25536,N_25211,N_25341);
nor U25537 (N_25537,N_25350,N_24842);
and U25538 (N_25538,N_25006,N_24973);
and U25539 (N_25539,N_25140,N_25054);
nor U25540 (N_25540,N_24054,N_25017);
and U25541 (N_25541,N_25316,N_24690);
xor U25542 (N_25542,N_24440,N_24492);
nand U25543 (N_25543,N_25074,N_24694);
or U25544 (N_25544,N_24478,N_24410);
xnor U25545 (N_25545,N_24829,N_24955);
nand U25546 (N_25546,N_24630,N_25161);
and U25547 (N_25547,N_25463,N_24256);
xor U25548 (N_25548,N_25032,N_24416);
or U25549 (N_25549,N_24914,N_25085);
nor U25550 (N_25550,N_25425,N_24109);
or U25551 (N_25551,N_24851,N_24940);
or U25552 (N_25552,N_24828,N_24246);
or U25553 (N_25553,N_25498,N_24105);
nand U25554 (N_25554,N_24874,N_25486);
or U25555 (N_25555,N_25308,N_24755);
or U25556 (N_25556,N_25395,N_25099);
xor U25557 (N_25557,N_24360,N_24476);
nor U25558 (N_25558,N_24668,N_24121);
and U25559 (N_25559,N_24938,N_24191);
xnor U25560 (N_25560,N_24852,N_24685);
xnor U25561 (N_25561,N_25291,N_25070);
and U25562 (N_25562,N_24037,N_24713);
nor U25563 (N_25563,N_24333,N_24597);
and U25564 (N_25564,N_24444,N_25337);
and U25565 (N_25565,N_25214,N_25255);
nor U25566 (N_25566,N_25016,N_25172);
nor U25567 (N_25567,N_24723,N_25028);
and U25568 (N_25568,N_24375,N_24599);
and U25569 (N_25569,N_24279,N_24386);
and U25570 (N_25570,N_25179,N_24783);
xor U25571 (N_25571,N_24174,N_24436);
nand U25572 (N_25572,N_24996,N_25010);
and U25573 (N_25573,N_24482,N_24563);
nor U25574 (N_25574,N_24549,N_24750);
nor U25575 (N_25575,N_25305,N_24882);
nor U25576 (N_25576,N_24005,N_24569);
xnor U25577 (N_25577,N_24650,N_24752);
and U25578 (N_25578,N_24902,N_25134);
nor U25579 (N_25579,N_24212,N_24001);
xor U25580 (N_25580,N_24226,N_24434);
nand U25581 (N_25581,N_24056,N_24303);
nand U25582 (N_25582,N_24097,N_24203);
nor U25583 (N_25583,N_25475,N_24149);
and U25584 (N_25584,N_24074,N_25324);
nor U25585 (N_25585,N_24510,N_25294);
and U25586 (N_25586,N_25411,N_25353);
or U25587 (N_25587,N_24509,N_25493);
or U25588 (N_25588,N_24340,N_25409);
nor U25589 (N_25589,N_25336,N_24449);
xnor U25590 (N_25590,N_25015,N_25278);
or U25591 (N_25591,N_24168,N_24898);
and U25592 (N_25592,N_24746,N_24531);
and U25593 (N_25593,N_25103,N_25218);
and U25594 (N_25594,N_25205,N_24151);
or U25595 (N_25595,N_24181,N_24180);
nor U25596 (N_25596,N_24832,N_25426);
nor U25597 (N_25597,N_24223,N_25335);
nor U25598 (N_25598,N_24541,N_24773);
or U25599 (N_25599,N_24915,N_24779);
nand U25600 (N_25600,N_25227,N_25012);
or U25601 (N_25601,N_24472,N_25221);
or U25602 (N_25602,N_24102,N_24888);
or U25603 (N_25603,N_24911,N_24692);
nor U25604 (N_25604,N_24679,N_25267);
and U25605 (N_25605,N_24807,N_24719);
or U25606 (N_25606,N_25364,N_24077);
and U25607 (N_25607,N_24084,N_24895);
nor U25608 (N_25608,N_24066,N_25471);
nor U25609 (N_25609,N_24220,N_24524);
nand U25610 (N_25610,N_25259,N_24607);
or U25611 (N_25611,N_24099,N_25332);
nor U25612 (N_25612,N_25287,N_24264);
nor U25613 (N_25613,N_24002,N_25086);
xnor U25614 (N_25614,N_25290,N_24273);
and U25615 (N_25615,N_25046,N_25257);
nand U25616 (N_25616,N_24873,N_24604);
nor U25617 (N_25617,N_24301,N_24496);
and U25618 (N_25618,N_25217,N_24804);
and U25619 (N_25619,N_24024,N_24213);
xor U25620 (N_25620,N_24753,N_24701);
nor U25621 (N_25621,N_24869,N_24556);
and U25622 (N_25622,N_24332,N_25173);
nand U25623 (N_25623,N_24565,N_25049);
and U25624 (N_25624,N_25111,N_25389);
nand U25625 (N_25625,N_24495,N_24425);
and U25626 (N_25626,N_25368,N_25472);
and U25627 (N_25627,N_24560,N_24784);
or U25628 (N_25628,N_24396,N_24224);
xor U25629 (N_25629,N_24031,N_25147);
and U25630 (N_25630,N_24678,N_25077);
nand U25631 (N_25631,N_25063,N_24485);
nor U25632 (N_25632,N_24321,N_24886);
nand U25633 (N_25633,N_24349,N_25485);
or U25634 (N_25634,N_25029,N_24450);
or U25635 (N_25635,N_24285,N_24816);
or U25636 (N_25636,N_24809,N_24900);
and U25637 (N_25637,N_24818,N_24395);
nor U25638 (N_25638,N_25182,N_24658);
xnor U25639 (N_25639,N_24372,N_25265);
nor U25640 (N_25640,N_24262,N_24454);
nor U25641 (N_25641,N_25230,N_24076);
nor U25642 (N_25642,N_24218,N_24848);
xor U25643 (N_25643,N_25199,N_24331);
xor U25644 (N_25644,N_25481,N_25301);
and U25645 (N_25645,N_24664,N_24391);
xor U25646 (N_25646,N_24439,N_24570);
nand U25647 (N_25647,N_24982,N_24126);
nand U25648 (N_25648,N_24728,N_25158);
xor U25649 (N_25649,N_24374,N_24930);
or U25650 (N_25650,N_25040,N_25196);
nand U25651 (N_25651,N_24574,N_24239);
and U25652 (N_25652,N_24924,N_24286);
or U25653 (N_25653,N_25170,N_25138);
nand U25654 (N_25654,N_25351,N_24408);
nor U25655 (N_25655,N_24884,N_25256);
nand U25656 (N_25656,N_25285,N_25432);
xor U25657 (N_25657,N_24759,N_24781);
nand U25658 (N_25658,N_24101,N_24634);
nor U25659 (N_25659,N_24428,N_24370);
nand U25660 (N_25660,N_24163,N_24619);
and U25661 (N_25661,N_25470,N_24615);
and U25662 (N_25662,N_25131,N_24065);
xor U25663 (N_25663,N_25339,N_24993);
or U25664 (N_25664,N_25494,N_24871);
nand U25665 (N_25665,N_24743,N_24278);
and U25666 (N_25666,N_24917,N_24612);
xnor U25667 (N_25667,N_24269,N_24545);
xnor U25668 (N_25668,N_25283,N_24782);
nor U25669 (N_25669,N_24614,N_25478);
and U25670 (N_25670,N_24653,N_24355);
nand U25671 (N_25671,N_24398,N_24124);
xor U25672 (N_25672,N_24584,N_24985);
nor U25673 (N_25673,N_25094,N_24698);
xnor U25674 (N_25674,N_25456,N_24277);
nor U25675 (N_25675,N_24422,N_24092);
and U25676 (N_25676,N_24605,N_24307);
and U25677 (N_25677,N_24159,N_24792);
xor U25678 (N_25678,N_24361,N_25109);
and U25679 (N_25679,N_24629,N_24382);
xnor U25680 (N_25680,N_24883,N_25300);
nand U25681 (N_25681,N_24933,N_24855);
or U25682 (N_25682,N_24061,N_24081);
nor U25683 (N_25683,N_24306,N_25021);
xor U25684 (N_25684,N_25295,N_24093);
nand U25685 (N_25685,N_24748,N_25178);
nand U25686 (N_25686,N_24276,N_25174);
nand U25687 (N_25687,N_24953,N_25082);
xnor U25688 (N_25688,N_24242,N_24316);
nand U25689 (N_25689,N_24550,N_25465);
xnor U25690 (N_25690,N_25123,N_24974);
nor U25691 (N_25691,N_24800,N_25223);
nor U25692 (N_25692,N_24196,N_25358);
xor U25693 (N_25693,N_24125,N_25027);
and U25694 (N_25694,N_24029,N_24548);
nor U25695 (N_25695,N_25410,N_25297);
xnor U25696 (N_25696,N_25299,N_25059);
and U25697 (N_25697,N_24090,N_24661);
xor U25698 (N_25698,N_24158,N_24173);
nor U25699 (N_25699,N_24362,N_24339);
or U25700 (N_25700,N_24868,N_25317);
nand U25701 (N_25701,N_24260,N_24992);
nor U25702 (N_25702,N_24537,N_24026);
and U25703 (N_25703,N_25483,N_24193);
nor U25704 (N_25704,N_24216,N_25165);
xnor U25705 (N_25705,N_24711,N_25144);
and U25706 (N_25706,N_25378,N_25365);
xor U25707 (N_25707,N_24790,N_24864);
nand U25708 (N_25708,N_25458,N_24027);
nor U25709 (N_25709,N_24460,N_24210);
nand U25710 (N_25710,N_25459,N_25228);
nand U25711 (N_25711,N_24532,N_24704);
and U25712 (N_25712,N_25405,N_24770);
or U25713 (N_25713,N_24381,N_24437);
nand U25714 (N_25714,N_24887,N_24538);
nand U25715 (N_25715,N_25473,N_24860);
nand U25716 (N_25716,N_25268,N_25124);
and U25717 (N_25717,N_24075,N_24356);
or U25718 (N_25718,N_25330,N_25304);
or U25719 (N_25719,N_24847,N_24899);
xnor U25720 (N_25720,N_24967,N_24108);
nand U25721 (N_25721,N_24910,N_25443);
or U25722 (N_25722,N_25314,N_24787);
and U25723 (N_25723,N_25377,N_24506);
and U25724 (N_25724,N_24129,N_24956);
xnor U25725 (N_25725,N_24834,N_25089);
xor U25726 (N_25726,N_24544,N_24591);
and U25727 (N_25727,N_24192,N_24946);
nor U25728 (N_25728,N_24572,N_24494);
and U25729 (N_25729,N_24359,N_24707);
nor U25730 (N_25730,N_24096,N_25428);
and U25731 (N_25731,N_25344,N_24813);
xnor U25732 (N_25732,N_24794,N_25420);
nand U25733 (N_25733,N_25447,N_25435);
and U25734 (N_25734,N_24880,N_24778);
nand U25735 (N_25735,N_24222,N_25288);
or U25736 (N_25736,N_25119,N_25439);
xnor U25737 (N_25737,N_25204,N_25148);
nor U25738 (N_25738,N_25164,N_24867);
xor U25739 (N_25739,N_24417,N_24823);
nor U25740 (N_25740,N_24551,N_24589);
nand U25741 (N_25741,N_24747,N_25326);
nand U25742 (N_25742,N_25137,N_24473);
xor U25743 (N_25743,N_24811,N_24486);
or U25744 (N_25744,N_25133,N_24032);
nand U25745 (N_25745,N_24722,N_25242);
xnor U25746 (N_25746,N_24997,N_24963);
xnor U25747 (N_25747,N_24691,N_24407);
and U25748 (N_25748,N_25302,N_25118);
and U25749 (N_25749,N_25495,N_25396);
xnor U25750 (N_25750,N_24237,N_24209);
xor U25751 (N_25751,N_24048,N_24905);
xor U25752 (N_25752,N_25236,N_24826);
or U25753 (N_25753,N_24948,N_24189);
and U25754 (N_25754,N_25359,N_24385);
or U25755 (N_25755,N_24302,N_24194);
xnor U25756 (N_25756,N_25277,N_25421);
or U25757 (N_25757,N_25129,N_25424);
and U25758 (N_25758,N_24161,N_24042);
nand U25759 (N_25759,N_24866,N_24009);
xor U25760 (N_25760,N_25220,N_24643);
xnor U25761 (N_25761,N_25321,N_25446);
nor U25762 (N_25762,N_24720,N_24153);
or U25763 (N_25763,N_24513,N_24505);
xor U25764 (N_25764,N_24474,N_24377);
or U25765 (N_25765,N_24272,N_24043);
xor U25766 (N_25766,N_24775,N_24111);
and U25767 (N_25767,N_24319,N_24676);
and U25768 (N_25768,N_25487,N_24215);
and U25769 (N_25769,N_24919,N_24353);
nand U25770 (N_25770,N_24502,N_24517);
nor U25771 (N_25771,N_25113,N_24774);
and U25772 (N_25772,N_24730,N_24364);
and U25773 (N_25773,N_24702,N_24705);
nand U25774 (N_25774,N_24089,N_24925);
xor U25775 (N_25775,N_24490,N_24830);
nand U25776 (N_25776,N_24312,N_25194);
or U25777 (N_25777,N_24341,N_24347);
or U25778 (N_25778,N_24631,N_24791);
or U25779 (N_25779,N_24889,N_24935);
or U25780 (N_25780,N_24808,N_24558);
nand U25781 (N_25781,N_25269,N_24641);
or U25782 (N_25782,N_25202,N_24461);
or U25783 (N_25783,N_24683,N_25052);
or U25784 (N_25784,N_24363,N_25184);
nand U25785 (N_25785,N_25163,N_25219);
xor U25786 (N_25786,N_25404,N_25452);
nor U25787 (N_25787,N_24234,N_24164);
or U25788 (N_25788,N_25333,N_24104);
nand U25789 (N_25789,N_25056,N_24843);
and U25790 (N_25790,N_24145,N_25169);
and U25791 (N_25791,N_24309,N_24799);
nor U25792 (N_25792,N_24771,N_24471);
or U25793 (N_25793,N_25002,N_25212);
or U25794 (N_25794,N_25100,N_24367);
nor U25795 (N_25795,N_24069,N_24764);
nand U25796 (N_25796,N_24432,N_24606);
and U25797 (N_25797,N_24950,N_25438);
nor U25798 (N_25798,N_25388,N_24632);
and U25799 (N_25799,N_24766,N_24835);
xnor U25800 (N_25800,N_24696,N_24959);
and U25801 (N_25801,N_24304,N_25253);
and U25802 (N_25802,N_25372,N_25116);
or U25803 (N_25803,N_24579,N_24175);
and U25804 (N_25804,N_25231,N_24710);
and U25805 (N_25805,N_24585,N_25423);
nand U25806 (N_25806,N_24185,N_25306);
nor U25807 (N_25807,N_25071,N_24839);
nand U25808 (N_25808,N_25386,N_24981);
or U25809 (N_25809,N_25051,N_24738);
nand U25810 (N_25810,N_25298,N_24357);
and U25811 (N_25811,N_24515,N_24618);
or U25812 (N_25812,N_25266,N_24964);
or U25813 (N_25813,N_24609,N_25431);
nor U25814 (N_25814,N_25261,N_24477);
and U25815 (N_25815,N_24621,N_24378);
nand U25816 (N_25816,N_24318,N_25477);
or U25817 (N_25817,N_24610,N_25079);
and U25818 (N_25818,N_24846,N_25433);
or U25819 (N_25819,N_25057,N_25289);
and U25820 (N_25820,N_25488,N_24392);
nand U25821 (N_25821,N_24525,N_25043);
xnor U25822 (N_25822,N_24561,N_24299);
nand U25823 (N_25823,N_25121,N_25108);
xnor U25824 (N_25824,N_25407,N_25391);
and U25825 (N_25825,N_25026,N_24252);
or U25826 (N_25826,N_25361,N_24709);
xnor U25827 (N_25827,N_24559,N_24943);
nand U25828 (N_25828,N_24429,N_24801);
nand U25829 (N_25829,N_25023,N_24231);
or U25830 (N_25830,N_24712,N_24942);
nor U25831 (N_25831,N_25047,N_25024);
nand U25832 (N_25832,N_25429,N_24156);
nor U25833 (N_25833,N_25454,N_24393);
xor U25834 (N_25834,N_24297,N_25461);
nor U25835 (N_25835,N_24825,N_25375);
and U25836 (N_25836,N_24007,N_24994);
nor U25837 (N_25837,N_24403,N_24110);
nor U25838 (N_25838,N_24073,N_24131);
or U25839 (N_25839,N_25105,N_24539);
and U25840 (N_25840,N_25360,N_24588);
and U25841 (N_25841,N_24795,N_24885);
or U25842 (N_25842,N_25484,N_24965);
and U25843 (N_25843,N_24282,N_24453);
nand U25844 (N_25844,N_24672,N_24063);
nand U25845 (N_25845,N_25035,N_25346);
nand U25846 (N_25846,N_24856,N_25050);
and U25847 (N_25847,N_24071,N_25307);
or U25848 (N_25848,N_25352,N_25284);
or U25849 (N_25849,N_24675,N_24369);
nand U25850 (N_25850,N_24399,N_24803);
nand U25851 (N_25851,N_25087,N_24921);
and U25852 (N_25852,N_24445,N_24814);
or U25853 (N_25853,N_24430,N_24734);
xnor U25854 (N_25854,N_24136,N_25160);
xor U25855 (N_25855,N_24133,N_24697);
or U25856 (N_25856,N_24366,N_24271);
and U25857 (N_25857,N_24972,N_24228);
or U25858 (N_25858,N_25011,N_24291);
nand U25859 (N_25859,N_24499,N_24815);
or U25860 (N_25860,N_25499,N_24821);
or U25861 (N_25861,N_24441,N_25455);
and U25862 (N_25862,N_24595,N_24833);
or U25863 (N_25863,N_25225,N_24741);
xnor U25864 (N_25864,N_24334,N_24198);
nor U25865 (N_25865,N_24463,N_24881);
nand U25866 (N_25866,N_24098,N_24051);
or U25867 (N_25867,N_25496,N_24908);
or U25868 (N_25868,N_24642,N_24283);
xnor U25869 (N_25869,N_25076,N_25482);
nor U25870 (N_25870,N_24023,N_24777);
xor U25871 (N_25871,N_24944,N_24443);
or U25872 (N_25872,N_24916,N_24527);
nor U25873 (N_25873,N_24893,N_24677);
xor U25874 (N_25874,N_25251,N_24623);
or U25875 (N_25875,N_24901,N_24155);
or U25876 (N_25876,N_24979,N_24238);
nor U25877 (N_25877,N_24796,N_24526);
nor U25878 (N_25878,N_24822,N_24716);
xnor U25879 (N_25879,N_25000,N_24507);
nand U25880 (N_25880,N_24128,N_25383);
or U25881 (N_25881,N_24030,N_25345);
or U25882 (N_25882,N_25093,N_25191);
and U25883 (N_25883,N_25045,N_24421);
nand U25884 (N_25884,N_24785,N_24613);
and U25885 (N_25885,N_25480,N_24183);
and U25886 (N_25886,N_24969,N_25393);
and U25887 (N_25887,N_24208,N_24251);
xor U25888 (N_25888,N_25362,N_24862);
nand U25889 (N_25889,N_24763,N_24966);
or U25890 (N_25890,N_24715,N_24831);
or U25891 (N_25891,N_25394,N_25209);
or U25892 (N_25892,N_24654,N_24446);
nor U25893 (N_25893,N_24127,N_25038);
or U25894 (N_25894,N_24330,N_24433);
or U25895 (N_25895,N_24214,N_25247);
nor U25896 (N_25896,N_25083,N_24424);
nand U25897 (N_25897,N_24257,N_24512);
nand U25898 (N_25898,N_24975,N_24352);
nor U25899 (N_25899,N_24624,N_24529);
xor U25900 (N_25900,N_24418,N_24566);
and U25901 (N_25901,N_24265,N_24055);
xor U25902 (N_25902,N_24957,N_25249);
and U25903 (N_25903,N_24518,N_24891);
nand U25904 (N_25904,N_24977,N_24397);
xnor U25905 (N_25905,N_25309,N_24960);
xnor U25906 (N_25906,N_24480,N_25490);
xor U25907 (N_25907,N_25112,N_25371);
and U25908 (N_25908,N_24258,N_24522);
xnor U25909 (N_25909,N_24058,N_25126);
nor U25910 (N_25910,N_25175,N_24991);
nand U25911 (N_25911,N_24797,N_24376);
and U25912 (N_25912,N_24336,N_24420);
xor U25913 (N_25913,N_24247,N_24423);
nand U25914 (N_25914,N_24249,N_24295);
or U25915 (N_25915,N_25198,N_24567);
nand U25916 (N_25916,N_24988,N_24687);
nand U25917 (N_25917,N_24068,N_24229);
and U25918 (N_25918,N_24300,N_25025);
nor U25919 (N_25919,N_24406,N_25296);
xnor U25920 (N_25920,N_24036,N_25241);
and U25921 (N_25921,N_24986,N_24447);
or U25922 (N_25922,N_25380,N_24186);
or U25923 (N_25923,N_25244,N_24594);
or U25924 (N_25924,N_24827,N_25460);
nor U25925 (N_25925,N_25328,N_24281);
or U25926 (N_25926,N_24458,N_24254);
nor U25927 (N_25927,N_25096,N_25319);
or U25928 (N_25928,N_24195,N_25382);
nor U25929 (N_25929,N_24655,N_24451);
xor U25930 (N_25930,N_24949,N_24789);
and U25931 (N_25931,N_24922,N_24798);
and U25932 (N_25932,N_24926,N_25376);
or U25933 (N_25933,N_24990,N_24178);
nor U25934 (N_25934,N_25366,N_25462);
xor U25935 (N_25935,N_24543,N_24000);
nand U25936 (N_25936,N_25379,N_24487);
nand U25937 (N_25937,N_24388,N_24958);
and U25938 (N_25938,N_24731,N_24086);
and U25939 (N_25939,N_24622,N_24894);
nand U25940 (N_25940,N_24503,N_25222);
nor U25941 (N_25941,N_25413,N_25450);
and U25942 (N_25942,N_24590,N_25215);
and U25943 (N_25943,N_25467,N_24941);
xnor U25944 (N_25944,N_25479,N_25381);
xnor U25945 (N_25945,N_25197,N_24931);
or U25946 (N_25946,N_24172,N_25088);
or U25947 (N_25947,N_25342,N_24442);
xnor U25948 (N_25948,N_24328,N_24095);
xor U25949 (N_25949,N_25186,N_24394);
xor U25950 (N_25950,N_24409,N_24904);
nor U25951 (N_25951,N_24721,N_25048);
nor U25952 (N_25952,N_24426,N_24872);
nand U25953 (N_25953,N_24844,N_24470);
nor U25954 (N_25954,N_24912,N_25136);
nand U25955 (N_25955,N_24401,N_24100);
xnor U25956 (N_25956,N_24592,N_24140);
xor U25957 (N_25957,N_24368,N_24718);
or U25958 (N_25958,N_24983,N_24044);
and U25959 (N_25959,N_25260,N_24467);
xnor U25960 (N_25960,N_25206,N_24865);
nor U25961 (N_25961,N_25067,N_24670);
or U25962 (N_25962,N_24040,N_25444);
and U25963 (N_25963,N_25279,N_24135);
or U25964 (N_25964,N_24736,N_24601);
and U25965 (N_25965,N_24817,N_25022);
nor U25966 (N_25966,N_24729,N_24989);
xor U25967 (N_25967,N_25232,N_25037);
nand U25968 (N_25968,N_24274,N_24581);
or U25969 (N_25969,N_24176,N_25181);
and U25970 (N_25970,N_25125,N_24768);
and U25971 (N_25971,N_24937,N_24221);
nor U25972 (N_25972,N_24980,N_24600);
nor U25973 (N_25973,N_24358,N_24555);
nor U25974 (N_25974,N_24608,N_25320);
or U25975 (N_25975,N_25210,N_24003);
or U25976 (N_25976,N_24547,N_24112);
xnor U25977 (N_25977,N_25313,N_24681);
nand U25978 (N_25978,N_24365,N_25020);
and U25979 (N_25979,N_25142,N_24780);
or U25980 (N_25980,N_24671,N_24523);
and U25981 (N_25981,N_25252,N_25058);
and U25982 (N_25982,N_24190,N_24230);
and U25983 (N_25983,N_24861,N_24737);
or U25984 (N_25984,N_25234,N_25392);
xor U25985 (N_25985,N_25274,N_24324);
and U25986 (N_25986,N_24041,N_24059);
and U25987 (N_25987,N_24141,N_25187);
xnor U25988 (N_25988,N_24961,N_25387);
nor U25989 (N_25989,N_24936,N_25132);
and U25990 (N_25990,N_24636,N_24849);
and U25991 (N_25991,N_24275,N_24335);
nand U25992 (N_25992,N_24501,N_24462);
nand U25993 (N_25993,N_24735,N_24962);
xnor U25994 (N_25994,N_24015,N_25406);
nor U25995 (N_25995,N_24008,N_25448);
xor U25996 (N_25996,N_24651,N_24498);
or U25997 (N_25997,N_24907,N_24087);
and U25998 (N_25998,N_25449,N_24516);
and U25999 (N_25999,N_24038,N_24647);
or U26000 (N_26000,N_25117,N_24928);
xor U26001 (N_26001,N_25081,N_25007);
xnor U26002 (N_26002,N_24287,N_24952);
nor U26003 (N_26003,N_25271,N_24745);
nor U26004 (N_26004,N_24947,N_25356);
xor U26005 (N_26005,N_24402,N_25168);
or U26006 (N_26006,N_24464,N_24665);
nor U26007 (N_26007,N_25003,N_25282);
nor U26008 (N_26008,N_24317,N_24118);
nand U26009 (N_26009,N_24179,N_24680);
or U26010 (N_26010,N_24227,N_24999);
or U26011 (N_26011,N_25189,N_24520);
nor U26012 (N_26012,N_24625,N_25363);
or U26013 (N_26013,N_24019,N_25343);
and U26014 (N_26014,N_24786,N_25412);
or U26015 (N_26015,N_25176,N_24863);
xor U26016 (N_26016,N_24200,N_24667);
nor U26017 (N_26017,N_24327,N_24708);
or U26018 (N_26018,N_24130,N_24383);
or U26019 (N_26019,N_24456,N_24479);
or U26020 (N_26020,N_24727,N_24659);
and U26021 (N_26021,N_25042,N_24666);
nand U26022 (N_26022,N_25369,N_24182);
xor U26023 (N_26023,N_24207,N_24345);
and U26024 (N_26024,N_24984,N_25240);
or U26025 (N_26025,N_24806,N_24326);
nand U26026 (N_26026,N_25195,N_25120);
or U26027 (N_26027,N_24767,N_24859);
nor U26028 (N_26028,N_24157,N_25009);
or U26029 (N_26029,N_24266,N_24014);
and U26030 (N_26030,N_24998,N_24144);
nand U26031 (N_26031,N_25374,N_24308);
or U26032 (N_26032,N_25033,N_24660);
nor U26033 (N_26033,N_24744,N_24626);
nor U26034 (N_26034,N_25233,N_24107);
nand U26035 (N_26035,N_24776,N_24267);
and U26036 (N_26036,N_24289,N_25292);
and U26037 (N_26037,N_24106,N_24546);
and U26038 (N_26038,N_24586,N_24337);
and U26039 (N_26039,N_24138,N_25440);
xnor U26040 (N_26040,N_25213,N_24793);
nand U26041 (N_26041,N_24897,N_25323);
nor U26042 (N_26042,N_24010,N_24255);
and U26043 (N_26043,N_24020,N_25075);
nor U26044 (N_26044,N_24165,N_25403);
and U26045 (N_26045,N_25466,N_24117);
nand U26046 (N_26046,N_24348,N_24740);
xnor U26047 (N_26047,N_24248,N_24243);
and U26048 (N_26048,N_24245,N_24013);
or U26049 (N_26049,N_25402,N_24870);
and U26050 (N_26050,N_24419,N_24343);
xor U26051 (N_26051,N_24838,N_25239);
or U26052 (N_26052,N_25263,N_24968);
nand U26053 (N_26053,N_24296,N_24469);
nor U26054 (N_26054,N_24628,N_25250);
and U26055 (N_26055,N_25357,N_24540);
xnor U26056 (N_26056,N_24148,N_25180);
xnor U26057 (N_26057,N_24298,N_25329);
or U26058 (N_26058,N_24699,N_25229);
xnor U26059 (N_26059,N_25464,N_25072);
xnor U26060 (N_26060,N_25427,N_24582);
xor U26061 (N_26061,N_25226,N_24879);
and U26062 (N_26062,N_24103,N_25065);
or U26063 (N_26063,N_24412,N_25334);
nand U26064 (N_26064,N_25066,N_25060);
or U26065 (N_26065,N_25030,N_24292);
xnor U26066 (N_26066,N_24466,N_24232);
nor U26067 (N_26067,N_24167,N_24305);
nand U26068 (N_26068,N_25101,N_24519);
and U26069 (N_26069,N_24578,N_24384);
nor U26070 (N_26070,N_24491,N_25185);
or U26071 (N_26071,N_24329,N_24583);
or U26072 (N_26072,N_24577,N_25401);
or U26073 (N_26073,N_25200,N_25080);
xor U26074 (N_26074,N_24739,N_24603);
or U26075 (N_26075,N_24554,N_25145);
or U26076 (N_26076,N_24530,N_25441);
and U26077 (N_26077,N_24187,N_24812);
xnor U26078 (N_26078,N_25018,N_24971);
xor U26079 (N_26079,N_24875,N_24576);
nand U26080 (N_26080,N_24022,N_24920);
and U26081 (N_26081,N_25073,N_24211);
and U26082 (N_26082,N_24284,N_25153);
nand U26083 (N_26083,N_24113,N_25237);
nor U26084 (N_26084,N_25171,N_25453);
or U26085 (N_26085,N_24072,N_24703);
xnor U26086 (N_26086,N_24322,N_24052);
and U26087 (N_26087,N_24146,N_24154);
nand U26088 (N_26088,N_24270,N_24749);
and U26089 (N_26089,N_25245,N_24674);
and U26090 (N_26090,N_24342,N_24018);
nor U26091 (N_26091,N_24177,N_25192);
nand U26092 (N_26092,N_25036,N_25053);
nor U26093 (N_26093,N_25468,N_24841);
and U26094 (N_26094,N_24639,N_24954);
or U26095 (N_26095,N_24083,N_25122);
nand U26096 (N_26096,N_24533,N_25272);
nor U26097 (N_26097,N_24235,N_25064);
nand U26098 (N_26098,N_25318,N_24411);
xnor U26099 (N_26099,N_24627,N_24662);
nor U26100 (N_26100,N_24371,N_24404);
and U26101 (N_26101,N_25188,N_24028);
nor U26102 (N_26102,N_25031,N_25130);
xor U26103 (N_26103,N_24047,N_25155);
and U26104 (N_26104,N_24310,N_25183);
nand U26105 (N_26105,N_24616,N_25004);
nand U26106 (N_26106,N_25005,N_25258);
or U26107 (N_26107,N_24757,N_24754);
nor U26108 (N_26108,N_25419,N_25340);
xnor U26109 (N_26109,N_24049,N_25338);
nand U26110 (N_26110,N_25491,N_25430);
and U26111 (N_26111,N_24903,N_24134);
and U26112 (N_26112,N_25270,N_24923);
or U26113 (N_26113,N_24079,N_24457);
xor U26114 (N_26114,N_25159,N_24082);
or U26115 (N_26115,N_24311,N_25281);
and U26116 (N_26116,N_25208,N_25442);
nor U26117 (N_26117,N_25019,N_24649);
xnor U26118 (N_26118,N_25090,N_24481);
or U26119 (N_26119,N_24646,N_24890);
or U26120 (N_26120,N_24088,N_25084);
xnor U26121 (N_26121,N_25044,N_24896);
xor U26122 (N_26122,N_24455,N_24021);
xor U26123 (N_26123,N_25327,N_24534);
nor U26124 (N_26124,N_25008,N_24147);
and U26125 (N_26125,N_25110,N_24142);
and U26126 (N_26126,N_24204,N_25078);
or U26127 (N_26127,N_24483,N_25254);
xnor U26128 (N_26128,N_24119,N_24724);
nor U26129 (N_26129,N_25474,N_24488);
nor U26130 (N_26130,N_25398,N_25497);
nand U26131 (N_26131,N_24199,N_24017);
and U26132 (N_26132,N_25384,N_24448);
nand U26133 (N_26133,N_24170,N_24351);
nand U26134 (N_26134,N_24810,N_24927);
xor U26135 (N_26135,N_24225,N_25354);
nor U26136 (N_26136,N_24689,N_25489);
nor U26137 (N_26137,N_24820,N_24379);
and U26138 (N_26138,N_24150,N_24536);
nand U26139 (N_26139,N_24568,N_25311);
or U26140 (N_26140,N_25167,N_24593);
xor U26141 (N_26141,N_24772,N_25224);
nand U26142 (N_26142,N_24338,N_24080);
nor U26143 (N_26143,N_24116,N_25149);
or U26144 (N_26144,N_24160,N_25349);
xnor U26145 (N_26145,N_24995,N_24389);
nor U26146 (N_26146,N_24769,N_25315);
or U26147 (N_26147,N_24120,N_25102);
and U26148 (N_26148,N_25385,N_24913);
or U26149 (N_26149,N_24078,N_24035);
or U26150 (N_26150,N_24663,N_25107);
nor U26151 (N_26151,N_24313,N_25154);
and U26152 (N_26152,N_24034,N_24637);
nand U26153 (N_26153,N_25092,N_25162);
or U26154 (N_26154,N_24459,N_24325);
nor U26155 (N_26155,N_24760,N_24114);
or U26156 (N_26156,N_24493,N_25418);
or U26157 (N_26157,N_24714,N_24850);
xor U26158 (N_26158,N_24644,N_24573);
nand U26159 (N_26159,N_25061,N_24892);
nor U26160 (N_26160,N_25408,N_24122);
xnor U26161 (N_26161,N_24682,N_24280);
or U26162 (N_26162,N_24004,N_25143);
or U26163 (N_26163,N_24553,N_24261);
nor U26164 (N_26164,N_25201,N_25331);
nor U26165 (N_26165,N_24293,N_25166);
and U26166 (N_26166,N_25150,N_24244);
and U26167 (N_26167,N_25422,N_25445);
nand U26168 (N_26168,N_25348,N_24762);
or U26169 (N_26169,N_25310,N_24046);
xor U26170 (N_26170,N_25416,N_24091);
nor U26171 (N_26171,N_24945,N_24011);
or U26172 (N_26172,N_24413,N_24640);
or U26173 (N_26173,N_24645,N_24726);
xor U26174 (N_26174,N_24521,N_24067);
nand U26175 (N_26175,N_24987,N_24452);
xnor U26176 (N_26176,N_24706,N_25039);
nand U26177 (N_26177,N_25246,N_24350);
nor U26178 (N_26178,N_24288,N_24085);
nor U26179 (N_26179,N_24475,N_24123);
or U26180 (N_26180,N_24344,N_24438);
or U26181 (N_26181,N_25238,N_24197);
xor U26182 (N_26182,N_25322,N_25235);
or U26183 (N_26183,N_24500,N_24557);
and U26184 (N_26184,N_25275,N_24489);
nand U26185 (N_26185,N_24427,N_24053);
or U26186 (N_26186,N_24431,N_24137);
and U26187 (N_26187,N_24184,N_24854);
xor U26188 (N_26188,N_24837,N_24314);
nor U26189 (N_26189,N_24845,N_24970);
xor U26190 (N_26190,N_24162,N_24508);
and U26191 (N_26191,N_25303,N_25001);
nor U26192 (N_26192,N_24877,N_24686);
nand U26193 (N_26193,N_24139,N_25013);
xor U26194 (N_26194,N_24788,N_25397);
nand U26195 (N_26195,N_24542,N_25312);
and U26196 (N_26196,N_24050,N_24202);
xnor U26197 (N_26197,N_24761,N_24253);
nand U26198 (N_26198,N_25014,N_25034);
and U26199 (N_26199,N_24323,N_24094);
or U26200 (N_26200,N_24016,N_24929);
and U26201 (N_26201,N_24733,N_25492);
nand U26202 (N_26202,N_25434,N_24387);
nor U26203 (N_26203,N_24853,N_24951);
and U26204 (N_26204,N_24836,N_24169);
nor U26205 (N_26205,N_25190,N_24906);
or U26206 (N_26206,N_24633,N_24978);
and U26207 (N_26207,N_24857,N_24669);
or U26208 (N_26208,N_24057,N_24693);
and U26209 (N_26209,N_25127,N_25114);
or U26210 (N_26210,N_24217,N_24171);
or U26211 (N_26211,N_24320,N_24045);
and U26212 (N_26212,N_24290,N_25091);
and U26213 (N_26213,N_24354,N_24380);
or U26214 (N_26214,N_24201,N_24758);
or U26215 (N_26215,N_25139,N_25262);
or U26216 (N_26216,N_24596,N_25177);
nor U26217 (N_26217,N_24152,N_24840);
nor U26218 (N_26218,N_25207,N_24934);
or U26219 (N_26219,N_24656,N_24435);
xnor U26220 (N_26220,N_24400,N_25417);
nand U26221 (N_26221,N_24876,N_25097);
xnor U26222 (N_26222,N_24062,N_25128);
xor U26223 (N_26223,N_24390,N_24688);
nand U26224 (N_26224,N_25041,N_25156);
nor U26225 (N_26225,N_24932,N_24206);
and U26226 (N_26226,N_24060,N_24700);
nor U26227 (N_26227,N_24012,N_25276);
nor U26228 (N_26228,N_24143,N_24025);
xor U26229 (N_26229,N_25141,N_24166);
and U26230 (N_26230,N_24552,N_24819);
or U26231 (N_26231,N_24751,N_24240);
and U26232 (N_26232,N_24638,N_24346);
xnor U26233 (N_26233,N_24064,N_25325);
nor U26234 (N_26234,N_25135,N_24484);
xnor U26235 (N_26235,N_24294,N_24858);
and U26236 (N_26236,N_24695,N_25286);
nand U26237 (N_26237,N_24939,N_24415);
nor U26238 (N_26238,N_25095,N_24373);
or U26239 (N_26239,N_24648,N_24742);
xnor U26240 (N_26240,N_24465,N_25273);
nor U26241 (N_26241,N_24132,N_25068);
and U26242 (N_26242,N_25243,N_24824);
nor U26243 (N_26243,N_25476,N_24657);
xnor U26244 (N_26244,N_25152,N_25367);
nand U26245 (N_26245,N_25055,N_24562);
xnor U26246 (N_26246,N_25437,N_25373);
and U26247 (N_26247,N_25451,N_24717);
or U26248 (N_26248,N_24575,N_25248);
nor U26249 (N_26249,N_25115,N_24497);
nand U26250 (N_26250,N_24045,N_25382);
nor U26251 (N_26251,N_24257,N_24615);
and U26252 (N_26252,N_25432,N_24214);
xor U26253 (N_26253,N_24545,N_24098);
or U26254 (N_26254,N_25208,N_24098);
nor U26255 (N_26255,N_24486,N_24908);
nand U26256 (N_26256,N_24270,N_25348);
and U26257 (N_26257,N_24867,N_24014);
or U26258 (N_26258,N_25268,N_24020);
xor U26259 (N_26259,N_24998,N_24985);
nand U26260 (N_26260,N_25100,N_24413);
or U26261 (N_26261,N_24331,N_24153);
nand U26262 (N_26262,N_24243,N_25124);
nor U26263 (N_26263,N_25188,N_25194);
nand U26264 (N_26264,N_25329,N_25339);
nor U26265 (N_26265,N_24732,N_24647);
xor U26266 (N_26266,N_24523,N_25397);
and U26267 (N_26267,N_24511,N_24571);
nand U26268 (N_26268,N_24503,N_24443);
nor U26269 (N_26269,N_24618,N_24273);
nor U26270 (N_26270,N_25162,N_24984);
nor U26271 (N_26271,N_25419,N_25184);
xnor U26272 (N_26272,N_24633,N_24338);
nor U26273 (N_26273,N_24191,N_25137);
and U26274 (N_26274,N_24390,N_24161);
and U26275 (N_26275,N_24865,N_25126);
xnor U26276 (N_26276,N_24023,N_25047);
nand U26277 (N_26277,N_24027,N_24950);
nor U26278 (N_26278,N_24123,N_24506);
nand U26279 (N_26279,N_24472,N_24065);
nor U26280 (N_26280,N_24307,N_25338);
nor U26281 (N_26281,N_24720,N_25183);
nand U26282 (N_26282,N_25128,N_24684);
xor U26283 (N_26283,N_25330,N_25030);
nand U26284 (N_26284,N_24159,N_24568);
nand U26285 (N_26285,N_25075,N_24011);
xor U26286 (N_26286,N_24233,N_25461);
and U26287 (N_26287,N_24352,N_24766);
xnor U26288 (N_26288,N_25174,N_25153);
nor U26289 (N_26289,N_25345,N_24155);
nor U26290 (N_26290,N_25446,N_25180);
nand U26291 (N_26291,N_24540,N_24815);
nand U26292 (N_26292,N_24629,N_24253);
nor U26293 (N_26293,N_25434,N_25408);
xor U26294 (N_26294,N_25215,N_25085);
nand U26295 (N_26295,N_24647,N_25366);
xor U26296 (N_26296,N_24637,N_25391);
or U26297 (N_26297,N_24133,N_24601);
or U26298 (N_26298,N_24230,N_24572);
nor U26299 (N_26299,N_25189,N_24260);
and U26300 (N_26300,N_25130,N_25149);
nor U26301 (N_26301,N_24404,N_24112);
and U26302 (N_26302,N_24715,N_24621);
nand U26303 (N_26303,N_25125,N_24535);
xnor U26304 (N_26304,N_25489,N_25118);
and U26305 (N_26305,N_25082,N_25193);
nand U26306 (N_26306,N_25420,N_24666);
nor U26307 (N_26307,N_24290,N_25351);
nand U26308 (N_26308,N_25492,N_24814);
xnor U26309 (N_26309,N_25221,N_24185);
xor U26310 (N_26310,N_24273,N_24639);
nand U26311 (N_26311,N_24224,N_24383);
or U26312 (N_26312,N_25128,N_24224);
xor U26313 (N_26313,N_24857,N_24641);
xor U26314 (N_26314,N_24252,N_25247);
or U26315 (N_26315,N_25011,N_24084);
xor U26316 (N_26316,N_25331,N_24426);
nand U26317 (N_26317,N_25430,N_25107);
nor U26318 (N_26318,N_24373,N_25396);
and U26319 (N_26319,N_24287,N_24224);
or U26320 (N_26320,N_25156,N_25409);
and U26321 (N_26321,N_25046,N_24999);
or U26322 (N_26322,N_25489,N_24223);
and U26323 (N_26323,N_24499,N_24900);
nor U26324 (N_26324,N_24171,N_25002);
and U26325 (N_26325,N_24224,N_25444);
and U26326 (N_26326,N_24678,N_24438);
xor U26327 (N_26327,N_25009,N_24360);
nand U26328 (N_26328,N_24781,N_24989);
nor U26329 (N_26329,N_24198,N_25331);
and U26330 (N_26330,N_24474,N_24403);
or U26331 (N_26331,N_24737,N_25246);
nand U26332 (N_26332,N_24935,N_24003);
nand U26333 (N_26333,N_24667,N_25125);
and U26334 (N_26334,N_25392,N_24805);
nand U26335 (N_26335,N_25248,N_24178);
nor U26336 (N_26336,N_24190,N_24597);
nand U26337 (N_26337,N_24699,N_24260);
and U26338 (N_26338,N_24465,N_25428);
or U26339 (N_26339,N_24328,N_24407);
nor U26340 (N_26340,N_25363,N_24538);
nand U26341 (N_26341,N_24127,N_24070);
and U26342 (N_26342,N_25372,N_25429);
or U26343 (N_26343,N_24550,N_24782);
xnor U26344 (N_26344,N_24227,N_25022);
and U26345 (N_26345,N_25371,N_24247);
or U26346 (N_26346,N_25149,N_24860);
nand U26347 (N_26347,N_25399,N_24995);
xnor U26348 (N_26348,N_24465,N_25458);
and U26349 (N_26349,N_24747,N_24190);
or U26350 (N_26350,N_25458,N_25293);
xnor U26351 (N_26351,N_25087,N_24208);
nor U26352 (N_26352,N_24533,N_25372);
xor U26353 (N_26353,N_25435,N_24594);
nor U26354 (N_26354,N_25188,N_25477);
and U26355 (N_26355,N_24214,N_24429);
xnor U26356 (N_26356,N_24685,N_24667);
and U26357 (N_26357,N_24519,N_24164);
xor U26358 (N_26358,N_25206,N_25301);
xor U26359 (N_26359,N_25320,N_25129);
and U26360 (N_26360,N_25360,N_25250);
or U26361 (N_26361,N_24897,N_24194);
and U26362 (N_26362,N_24097,N_24979);
xnor U26363 (N_26363,N_24763,N_24923);
xnor U26364 (N_26364,N_24209,N_24009);
nor U26365 (N_26365,N_25307,N_24519);
nor U26366 (N_26366,N_25434,N_25239);
or U26367 (N_26367,N_24067,N_24615);
and U26368 (N_26368,N_24184,N_24719);
and U26369 (N_26369,N_24557,N_24204);
nand U26370 (N_26370,N_25460,N_24773);
or U26371 (N_26371,N_24407,N_25040);
nor U26372 (N_26372,N_25125,N_25422);
or U26373 (N_26373,N_24595,N_24665);
and U26374 (N_26374,N_24403,N_24725);
or U26375 (N_26375,N_24496,N_24541);
nand U26376 (N_26376,N_24361,N_25135);
nor U26377 (N_26377,N_25251,N_24286);
and U26378 (N_26378,N_24858,N_24731);
nor U26379 (N_26379,N_24618,N_24775);
or U26380 (N_26380,N_25090,N_25180);
nand U26381 (N_26381,N_24010,N_25085);
xor U26382 (N_26382,N_24536,N_24102);
xor U26383 (N_26383,N_24201,N_25499);
xor U26384 (N_26384,N_24970,N_25388);
nand U26385 (N_26385,N_24022,N_25024);
nand U26386 (N_26386,N_24221,N_24327);
nand U26387 (N_26387,N_24761,N_25121);
nor U26388 (N_26388,N_25168,N_24663);
and U26389 (N_26389,N_25312,N_24856);
and U26390 (N_26390,N_24463,N_25475);
or U26391 (N_26391,N_25453,N_24106);
or U26392 (N_26392,N_25110,N_25023);
and U26393 (N_26393,N_25022,N_24485);
xor U26394 (N_26394,N_24726,N_24786);
and U26395 (N_26395,N_25293,N_24728);
nand U26396 (N_26396,N_25208,N_24719);
and U26397 (N_26397,N_25285,N_25078);
or U26398 (N_26398,N_24996,N_24300);
xnor U26399 (N_26399,N_24549,N_25430);
nand U26400 (N_26400,N_24505,N_24310);
or U26401 (N_26401,N_25428,N_24496);
or U26402 (N_26402,N_24962,N_24903);
or U26403 (N_26403,N_24850,N_24492);
nand U26404 (N_26404,N_24530,N_24160);
nor U26405 (N_26405,N_25096,N_24216);
and U26406 (N_26406,N_24213,N_24868);
and U26407 (N_26407,N_24148,N_25262);
nand U26408 (N_26408,N_25206,N_25452);
nand U26409 (N_26409,N_25404,N_25052);
nor U26410 (N_26410,N_25240,N_24799);
and U26411 (N_26411,N_24008,N_24628);
nand U26412 (N_26412,N_25011,N_24941);
nor U26413 (N_26413,N_24325,N_24684);
nor U26414 (N_26414,N_24606,N_24631);
or U26415 (N_26415,N_24324,N_25384);
xnor U26416 (N_26416,N_24701,N_25283);
nor U26417 (N_26417,N_24302,N_24640);
or U26418 (N_26418,N_25011,N_25116);
xor U26419 (N_26419,N_24737,N_24173);
and U26420 (N_26420,N_24658,N_24143);
nand U26421 (N_26421,N_24944,N_24922);
nand U26422 (N_26422,N_24634,N_25000);
or U26423 (N_26423,N_24851,N_24368);
and U26424 (N_26424,N_24667,N_24459);
or U26425 (N_26425,N_25005,N_24585);
nor U26426 (N_26426,N_25209,N_24750);
and U26427 (N_26427,N_24674,N_24753);
or U26428 (N_26428,N_24126,N_24695);
nor U26429 (N_26429,N_24186,N_24556);
nand U26430 (N_26430,N_24894,N_24913);
nand U26431 (N_26431,N_25329,N_25084);
nor U26432 (N_26432,N_24809,N_24732);
xnor U26433 (N_26433,N_24262,N_24753);
nand U26434 (N_26434,N_24277,N_25369);
and U26435 (N_26435,N_24756,N_25168);
xor U26436 (N_26436,N_24640,N_25363);
nor U26437 (N_26437,N_24064,N_25052);
or U26438 (N_26438,N_24195,N_24576);
and U26439 (N_26439,N_24093,N_25308);
or U26440 (N_26440,N_24122,N_24878);
and U26441 (N_26441,N_24249,N_24459);
or U26442 (N_26442,N_24406,N_24569);
xor U26443 (N_26443,N_24716,N_24820);
and U26444 (N_26444,N_25077,N_25247);
or U26445 (N_26445,N_25093,N_24970);
nor U26446 (N_26446,N_24158,N_25194);
or U26447 (N_26447,N_24459,N_24434);
or U26448 (N_26448,N_24883,N_24072);
xnor U26449 (N_26449,N_25350,N_24794);
or U26450 (N_26450,N_25312,N_24208);
xnor U26451 (N_26451,N_24006,N_24073);
nor U26452 (N_26452,N_24643,N_24090);
nand U26453 (N_26453,N_24770,N_24116);
xnor U26454 (N_26454,N_24390,N_24149);
nand U26455 (N_26455,N_24435,N_24864);
nand U26456 (N_26456,N_24087,N_24597);
or U26457 (N_26457,N_25149,N_24716);
or U26458 (N_26458,N_25363,N_25018);
nand U26459 (N_26459,N_24588,N_24319);
and U26460 (N_26460,N_25386,N_25410);
xor U26461 (N_26461,N_24735,N_24823);
or U26462 (N_26462,N_24820,N_24714);
and U26463 (N_26463,N_24441,N_24033);
nand U26464 (N_26464,N_24253,N_24801);
nand U26465 (N_26465,N_24557,N_24138);
nor U26466 (N_26466,N_24856,N_24039);
xor U26467 (N_26467,N_24483,N_25343);
nor U26468 (N_26468,N_24200,N_24184);
nor U26469 (N_26469,N_24386,N_25192);
and U26470 (N_26470,N_25260,N_25218);
xnor U26471 (N_26471,N_24731,N_24802);
and U26472 (N_26472,N_24448,N_25131);
nor U26473 (N_26473,N_24929,N_24574);
nand U26474 (N_26474,N_24330,N_25082);
and U26475 (N_26475,N_24586,N_25137);
nor U26476 (N_26476,N_24623,N_24006);
or U26477 (N_26477,N_24562,N_24181);
and U26478 (N_26478,N_24318,N_25326);
nor U26479 (N_26479,N_24597,N_25431);
or U26480 (N_26480,N_24629,N_24041);
nor U26481 (N_26481,N_24127,N_24010);
xor U26482 (N_26482,N_25393,N_24062);
nand U26483 (N_26483,N_25391,N_24712);
and U26484 (N_26484,N_24034,N_24022);
xnor U26485 (N_26485,N_25279,N_24459);
or U26486 (N_26486,N_24214,N_25191);
xor U26487 (N_26487,N_24604,N_24992);
and U26488 (N_26488,N_24534,N_24239);
nor U26489 (N_26489,N_24638,N_24116);
or U26490 (N_26490,N_25370,N_24891);
nor U26491 (N_26491,N_24660,N_25124);
nand U26492 (N_26492,N_25179,N_25264);
nand U26493 (N_26493,N_25038,N_25232);
xor U26494 (N_26494,N_25471,N_24346);
or U26495 (N_26495,N_24324,N_25326);
and U26496 (N_26496,N_24524,N_24015);
and U26497 (N_26497,N_24395,N_25232);
nor U26498 (N_26498,N_25306,N_24648);
nor U26499 (N_26499,N_24198,N_24850);
xor U26500 (N_26500,N_24272,N_24855);
nor U26501 (N_26501,N_24056,N_25096);
xor U26502 (N_26502,N_24041,N_25013);
nand U26503 (N_26503,N_24428,N_25129);
xor U26504 (N_26504,N_24035,N_24642);
nand U26505 (N_26505,N_24622,N_25312);
nand U26506 (N_26506,N_24213,N_24709);
and U26507 (N_26507,N_24129,N_24058);
or U26508 (N_26508,N_24818,N_24365);
xor U26509 (N_26509,N_24256,N_24436);
and U26510 (N_26510,N_24469,N_24754);
nand U26511 (N_26511,N_24931,N_24469);
and U26512 (N_26512,N_24894,N_25066);
xnor U26513 (N_26513,N_25214,N_24391);
nor U26514 (N_26514,N_24734,N_25263);
and U26515 (N_26515,N_24535,N_24062);
and U26516 (N_26516,N_24850,N_25260);
and U26517 (N_26517,N_25057,N_24730);
and U26518 (N_26518,N_24421,N_25048);
xnor U26519 (N_26519,N_24372,N_25053);
nor U26520 (N_26520,N_25327,N_25132);
nand U26521 (N_26521,N_25175,N_24919);
or U26522 (N_26522,N_24806,N_25101);
xor U26523 (N_26523,N_24859,N_25287);
xor U26524 (N_26524,N_24936,N_24913);
or U26525 (N_26525,N_24383,N_25449);
nand U26526 (N_26526,N_24834,N_24013);
and U26527 (N_26527,N_24574,N_24289);
or U26528 (N_26528,N_25371,N_24957);
and U26529 (N_26529,N_24060,N_24706);
xor U26530 (N_26530,N_24383,N_24016);
or U26531 (N_26531,N_24541,N_25095);
nor U26532 (N_26532,N_24503,N_25157);
nor U26533 (N_26533,N_24885,N_24424);
and U26534 (N_26534,N_25067,N_24194);
nand U26535 (N_26535,N_24675,N_24140);
nand U26536 (N_26536,N_25142,N_24590);
and U26537 (N_26537,N_25435,N_24207);
and U26538 (N_26538,N_24115,N_25461);
xor U26539 (N_26539,N_24051,N_25492);
nand U26540 (N_26540,N_25286,N_25371);
nand U26541 (N_26541,N_25353,N_24845);
or U26542 (N_26542,N_24635,N_25205);
nand U26543 (N_26543,N_24540,N_24065);
nand U26544 (N_26544,N_25177,N_25367);
nand U26545 (N_26545,N_25103,N_24113);
nand U26546 (N_26546,N_24080,N_24335);
or U26547 (N_26547,N_24223,N_25316);
nand U26548 (N_26548,N_24157,N_24662);
or U26549 (N_26549,N_24555,N_25415);
nor U26550 (N_26550,N_24472,N_24556);
nor U26551 (N_26551,N_25349,N_24999);
or U26552 (N_26552,N_24880,N_24581);
or U26553 (N_26553,N_24701,N_25413);
nand U26554 (N_26554,N_25304,N_24813);
and U26555 (N_26555,N_25098,N_24599);
and U26556 (N_26556,N_24182,N_24100);
xor U26557 (N_26557,N_24468,N_24399);
and U26558 (N_26558,N_24034,N_25402);
xor U26559 (N_26559,N_25068,N_24291);
xnor U26560 (N_26560,N_25032,N_25393);
xnor U26561 (N_26561,N_24020,N_25123);
nand U26562 (N_26562,N_24393,N_25105);
and U26563 (N_26563,N_25119,N_24236);
nor U26564 (N_26564,N_24039,N_25165);
and U26565 (N_26565,N_24523,N_25495);
nor U26566 (N_26566,N_24397,N_25226);
nor U26567 (N_26567,N_24995,N_24065);
nand U26568 (N_26568,N_24048,N_25271);
nor U26569 (N_26569,N_24188,N_24083);
and U26570 (N_26570,N_25106,N_24032);
nor U26571 (N_26571,N_25415,N_24734);
xor U26572 (N_26572,N_25458,N_25161);
or U26573 (N_26573,N_24978,N_24184);
or U26574 (N_26574,N_24425,N_25164);
nor U26575 (N_26575,N_24180,N_25168);
and U26576 (N_26576,N_24971,N_25316);
or U26577 (N_26577,N_24170,N_24093);
and U26578 (N_26578,N_24672,N_25021);
or U26579 (N_26579,N_24315,N_25052);
nor U26580 (N_26580,N_25317,N_25103);
nor U26581 (N_26581,N_24929,N_25184);
xnor U26582 (N_26582,N_25335,N_24454);
nor U26583 (N_26583,N_24855,N_24355);
or U26584 (N_26584,N_24810,N_24393);
nand U26585 (N_26585,N_24123,N_25388);
xor U26586 (N_26586,N_24784,N_24263);
xor U26587 (N_26587,N_25281,N_24651);
xor U26588 (N_26588,N_24033,N_24169);
or U26589 (N_26589,N_24914,N_24094);
or U26590 (N_26590,N_25451,N_24041);
and U26591 (N_26591,N_24933,N_24672);
and U26592 (N_26592,N_25197,N_24965);
or U26593 (N_26593,N_24698,N_24257);
xor U26594 (N_26594,N_24591,N_25038);
or U26595 (N_26595,N_24480,N_24130);
and U26596 (N_26596,N_25378,N_25468);
and U26597 (N_26597,N_25345,N_25405);
nor U26598 (N_26598,N_25396,N_25392);
and U26599 (N_26599,N_25092,N_25282);
nand U26600 (N_26600,N_25237,N_24714);
nand U26601 (N_26601,N_25133,N_25241);
or U26602 (N_26602,N_25467,N_24956);
and U26603 (N_26603,N_24962,N_24620);
or U26604 (N_26604,N_24107,N_24335);
nand U26605 (N_26605,N_24888,N_24821);
and U26606 (N_26606,N_24637,N_24425);
nor U26607 (N_26607,N_24963,N_25220);
and U26608 (N_26608,N_25172,N_24072);
or U26609 (N_26609,N_24215,N_25172);
nor U26610 (N_26610,N_24947,N_24733);
xor U26611 (N_26611,N_24705,N_24406);
xnor U26612 (N_26612,N_25171,N_25287);
or U26613 (N_26613,N_24055,N_24013);
or U26614 (N_26614,N_25079,N_24967);
xor U26615 (N_26615,N_25282,N_25041);
nor U26616 (N_26616,N_25448,N_24034);
nand U26617 (N_26617,N_24893,N_25006);
or U26618 (N_26618,N_24512,N_25013);
or U26619 (N_26619,N_25196,N_25407);
xnor U26620 (N_26620,N_25136,N_24909);
and U26621 (N_26621,N_24070,N_24266);
nor U26622 (N_26622,N_24614,N_24843);
and U26623 (N_26623,N_24122,N_25472);
or U26624 (N_26624,N_24540,N_25161);
and U26625 (N_26625,N_24874,N_24480);
or U26626 (N_26626,N_24902,N_24019);
and U26627 (N_26627,N_24663,N_24053);
nor U26628 (N_26628,N_24222,N_25108);
nor U26629 (N_26629,N_24925,N_24842);
xnor U26630 (N_26630,N_24699,N_24341);
and U26631 (N_26631,N_25144,N_24261);
nand U26632 (N_26632,N_24102,N_25318);
or U26633 (N_26633,N_25314,N_25239);
nor U26634 (N_26634,N_24227,N_24191);
or U26635 (N_26635,N_24394,N_24354);
nand U26636 (N_26636,N_24483,N_24456);
xor U26637 (N_26637,N_24105,N_24602);
nor U26638 (N_26638,N_24921,N_24746);
or U26639 (N_26639,N_25465,N_25366);
nand U26640 (N_26640,N_24939,N_24162);
or U26641 (N_26641,N_24881,N_25227);
nor U26642 (N_26642,N_25068,N_24807);
nor U26643 (N_26643,N_24334,N_24467);
and U26644 (N_26644,N_24176,N_24515);
xnor U26645 (N_26645,N_24300,N_25193);
or U26646 (N_26646,N_25420,N_25363);
xor U26647 (N_26647,N_24018,N_24416);
nor U26648 (N_26648,N_24180,N_24392);
xor U26649 (N_26649,N_25299,N_24414);
nand U26650 (N_26650,N_24585,N_25260);
or U26651 (N_26651,N_24337,N_24220);
nand U26652 (N_26652,N_24849,N_25394);
or U26653 (N_26653,N_25162,N_24065);
and U26654 (N_26654,N_24984,N_24952);
or U26655 (N_26655,N_24954,N_24428);
xor U26656 (N_26656,N_24519,N_24778);
and U26657 (N_26657,N_24432,N_24912);
nand U26658 (N_26658,N_24929,N_24483);
nand U26659 (N_26659,N_24567,N_25037);
and U26660 (N_26660,N_25147,N_25453);
nand U26661 (N_26661,N_25289,N_25472);
nor U26662 (N_26662,N_24227,N_24529);
nand U26663 (N_26663,N_25149,N_24379);
or U26664 (N_26664,N_25490,N_24367);
xnor U26665 (N_26665,N_25311,N_24558);
and U26666 (N_26666,N_25483,N_24106);
xnor U26667 (N_26667,N_24326,N_25218);
or U26668 (N_26668,N_25236,N_24489);
nand U26669 (N_26669,N_24298,N_24306);
xnor U26670 (N_26670,N_24833,N_25188);
nor U26671 (N_26671,N_24023,N_25455);
or U26672 (N_26672,N_24091,N_24778);
nor U26673 (N_26673,N_24023,N_25383);
nand U26674 (N_26674,N_24686,N_25027);
xnor U26675 (N_26675,N_25496,N_25484);
nor U26676 (N_26676,N_24918,N_24748);
nor U26677 (N_26677,N_25433,N_24982);
xor U26678 (N_26678,N_24250,N_25057);
nor U26679 (N_26679,N_24878,N_24146);
xnor U26680 (N_26680,N_24550,N_24482);
and U26681 (N_26681,N_24185,N_24480);
xnor U26682 (N_26682,N_24341,N_25247);
xnor U26683 (N_26683,N_25485,N_25176);
or U26684 (N_26684,N_25398,N_24297);
xnor U26685 (N_26685,N_25344,N_25268);
nor U26686 (N_26686,N_24500,N_25159);
nand U26687 (N_26687,N_24712,N_25083);
nor U26688 (N_26688,N_24877,N_25186);
and U26689 (N_26689,N_25065,N_24484);
nand U26690 (N_26690,N_25170,N_24723);
xnor U26691 (N_26691,N_24515,N_24377);
xor U26692 (N_26692,N_25053,N_25088);
nand U26693 (N_26693,N_24589,N_24383);
nand U26694 (N_26694,N_25310,N_25247);
nand U26695 (N_26695,N_24791,N_25097);
nand U26696 (N_26696,N_24273,N_24522);
nand U26697 (N_26697,N_24049,N_25190);
nand U26698 (N_26698,N_25386,N_25473);
nor U26699 (N_26699,N_24817,N_25483);
and U26700 (N_26700,N_25347,N_25046);
and U26701 (N_26701,N_25167,N_24500);
or U26702 (N_26702,N_25164,N_25250);
and U26703 (N_26703,N_25037,N_24877);
nor U26704 (N_26704,N_24500,N_25208);
nor U26705 (N_26705,N_24511,N_24262);
or U26706 (N_26706,N_25120,N_24966);
and U26707 (N_26707,N_24319,N_24693);
xor U26708 (N_26708,N_24880,N_25267);
nor U26709 (N_26709,N_25490,N_25333);
or U26710 (N_26710,N_24230,N_24433);
xor U26711 (N_26711,N_24985,N_24553);
nor U26712 (N_26712,N_24806,N_24486);
nand U26713 (N_26713,N_24721,N_25384);
nor U26714 (N_26714,N_25355,N_25468);
xor U26715 (N_26715,N_24365,N_24371);
or U26716 (N_26716,N_25188,N_24763);
and U26717 (N_26717,N_24297,N_25251);
nor U26718 (N_26718,N_24652,N_25295);
and U26719 (N_26719,N_24942,N_24153);
and U26720 (N_26720,N_25126,N_24434);
and U26721 (N_26721,N_24800,N_24843);
nor U26722 (N_26722,N_24899,N_25193);
or U26723 (N_26723,N_25209,N_24718);
nor U26724 (N_26724,N_24854,N_24303);
xor U26725 (N_26725,N_24902,N_24783);
and U26726 (N_26726,N_24583,N_24578);
nand U26727 (N_26727,N_25287,N_24132);
and U26728 (N_26728,N_24923,N_24957);
and U26729 (N_26729,N_24331,N_24048);
or U26730 (N_26730,N_25097,N_24120);
xor U26731 (N_26731,N_24484,N_24821);
nor U26732 (N_26732,N_25309,N_25052);
or U26733 (N_26733,N_24106,N_24097);
nand U26734 (N_26734,N_25099,N_24202);
or U26735 (N_26735,N_25214,N_24660);
nor U26736 (N_26736,N_25475,N_24078);
and U26737 (N_26737,N_24193,N_24711);
xor U26738 (N_26738,N_24486,N_24316);
xnor U26739 (N_26739,N_25126,N_24946);
nor U26740 (N_26740,N_24801,N_24138);
or U26741 (N_26741,N_24658,N_25442);
xor U26742 (N_26742,N_25267,N_25191);
or U26743 (N_26743,N_24865,N_24509);
or U26744 (N_26744,N_25160,N_24258);
and U26745 (N_26745,N_25220,N_25059);
or U26746 (N_26746,N_25272,N_25367);
nand U26747 (N_26747,N_25364,N_25398);
nand U26748 (N_26748,N_24451,N_24155);
and U26749 (N_26749,N_24213,N_24001);
nand U26750 (N_26750,N_25387,N_25157);
nor U26751 (N_26751,N_24618,N_25086);
and U26752 (N_26752,N_24890,N_25005);
nor U26753 (N_26753,N_24378,N_25055);
or U26754 (N_26754,N_25428,N_24321);
xor U26755 (N_26755,N_24952,N_25013);
or U26756 (N_26756,N_24027,N_25348);
nand U26757 (N_26757,N_24223,N_25494);
nand U26758 (N_26758,N_24159,N_24621);
nand U26759 (N_26759,N_24799,N_24701);
nor U26760 (N_26760,N_24493,N_24995);
and U26761 (N_26761,N_24168,N_24741);
xnor U26762 (N_26762,N_25326,N_24027);
nand U26763 (N_26763,N_24027,N_24489);
xor U26764 (N_26764,N_24251,N_25041);
and U26765 (N_26765,N_25031,N_25203);
or U26766 (N_26766,N_25057,N_25116);
xor U26767 (N_26767,N_24003,N_25461);
nand U26768 (N_26768,N_24085,N_24219);
and U26769 (N_26769,N_24728,N_25109);
or U26770 (N_26770,N_25345,N_24890);
nand U26771 (N_26771,N_24824,N_24535);
nor U26772 (N_26772,N_25226,N_25326);
and U26773 (N_26773,N_25379,N_24550);
nor U26774 (N_26774,N_24864,N_24982);
or U26775 (N_26775,N_24498,N_25483);
nand U26776 (N_26776,N_24657,N_24154);
nor U26777 (N_26777,N_25000,N_24931);
nor U26778 (N_26778,N_24053,N_25460);
nor U26779 (N_26779,N_24537,N_25242);
xor U26780 (N_26780,N_24841,N_24037);
and U26781 (N_26781,N_24702,N_24791);
xnor U26782 (N_26782,N_25423,N_24289);
nand U26783 (N_26783,N_24705,N_25483);
xnor U26784 (N_26784,N_24669,N_24600);
nor U26785 (N_26785,N_24505,N_24511);
and U26786 (N_26786,N_24880,N_24809);
xnor U26787 (N_26787,N_25144,N_24870);
nor U26788 (N_26788,N_25375,N_25381);
and U26789 (N_26789,N_24968,N_24213);
xor U26790 (N_26790,N_24538,N_24635);
nor U26791 (N_26791,N_24328,N_24215);
xor U26792 (N_26792,N_24471,N_24873);
nor U26793 (N_26793,N_24345,N_24697);
nand U26794 (N_26794,N_24179,N_24550);
and U26795 (N_26795,N_25365,N_25372);
or U26796 (N_26796,N_24727,N_25496);
xnor U26797 (N_26797,N_24273,N_25045);
or U26798 (N_26798,N_24339,N_24890);
or U26799 (N_26799,N_24768,N_25065);
nand U26800 (N_26800,N_24807,N_24829);
nor U26801 (N_26801,N_24417,N_24464);
or U26802 (N_26802,N_24655,N_25075);
xnor U26803 (N_26803,N_25355,N_24345);
or U26804 (N_26804,N_24214,N_24478);
nor U26805 (N_26805,N_25064,N_24568);
xnor U26806 (N_26806,N_24386,N_24978);
or U26807 (N_26807,N_24606,N_25312);
xnor U26808 (N_26808,N_24972,N_24008);
or U26809 (N_26809,N_24398,N_25173);
and U26810 (N_26810,N_24417,N_24209);
and U26811 (N_26811,N_24241,N_25233);
and U26812 (N_26812,N_24348,N_25090);
and U26813 (N_26813,N_24446,N_24948);
nor U26814 (N_26814,N_24893,N_24372);
nand U26815 (N_26815,N_25336,N_25125);
nor U26816 (N_26816,N_25407,N_24304);
xor U26817 (N_26817,N_24691,N_24830);
or U26818 (N_26818,N_24214,N_25272);
xnor U26819 (N_26819,N_25020,N_24911);
nand U26820 (N_26820,N_25139,N_25331);
and U26821 (N_26821,N_24267,N_25374);
xor U26822 (N_26822,N_24566,N_24984);
nor U26823 (N_26823,N_24982,N_24788);
nand U26824 (N_26824,N_24172,N_24641);
or U26825 (N_26825,N_24919,N_24529);
and U26826 (N_26826,N_24729,N_24642);
and U26827 (N_26827,N_25150,N_24082);
nor U26828 (N_26828,N_24794,N_25407);
and U26829 (N_26829,N_24542,N_24942);
nand U26830 (N_26830,N_24514,N_24296);
or U26831 (N_26831,N_24610,N_25112);
and U26832 (N_26832,N_24731,N_24738);
or U26833 (N_26833,N_25142,N_24810);
or U26834 (N_26834,N_25059,N_24788);
nor U26835 (N_26835,N_24706,N_25277);
or U26836 (N_26836,N_24053,N_24346);
or U26837 (N_26837,N_24322,N_24175);
nor U26838 (N_26838,N_24238,N_25476);
and U26839 (N_26839,N_24396,N_24430);
xor U26840 (N_26840,N_24160,N_25192);
nor U26841 (N_26841,N_25439,N_24799);
or U26842 (N_26842,N_25152,N_25392);
or U26843 (N_26843,N_25234,N_24944);
nand U26844 (N_26844,N_25288,N_24370);
or U26845 (N_26845,N_25300,N_24560);
nor U26846 (N_26846,N_24243,N_25106);
xnor U26847 (N_26847,N_24323,N_24813);
nor U26848 (N_26848,N_25486,N_24922);
or U26849 (N_26849,N_24466,N_25220);
and U26850 (N_26850,N_24942,N_24603);
and U26851 (N_26851,N_24333,N_24859);
and U26852 (N_26852,N_24891,N_24427);
nand U26853 (N_26853,N_24880,N_25328);
nand U26854 (N_26854,N_25015,N_24585);
xnor U26855 (N_26855,N_25221,N_24366);
and U26856 (N_26856,N_24839,N_24720);
and U26857 (N_26857,N_25352,N_24546);
and U26858 (N_26858,N_24983,N_24585);
and U26859 (N_26859,N_25042,N_24761);
nor U26860 (N_26860,N_25216,N_24902);
nand U26861 (N_26861,N_24591,N_24276);
or U26862 (N_26862,N_24394,N_25221);
nand U26863 (N_26863,N_24149,N_25454);
and U26864 (N_26864,N_24865,N_24852);
nor U26865 (N_26865,N_24526,N_24106);
and U26866 (N_26866,N_25067,N_24259);
or U26867 (N_26867,N_25008,N_24632);
and U26868 (N_26868,N_25028,N_24030);
nor U26869 (N_26869,N_24234,N_24835);
nor U26870 (N_26870,N_24987,N_24165);
and U26871 (N_26871,N_24576,N_24798);
xor U26872 (N_26872,N_24458,N_24624);
xnor U26873 (N_26873,N_24028,N_25486);
and U26874 (N_26874,N_24786,N_25491);
and U26875 (N_26875,N_25135,N_25203);
or U26876 (N_26876,N_25014,N_25323);
nand U26877 (N_26877,N_24318,N_24562);
or U26878 (N_26878,N_24762,N_25139);
and U26879 (N_26879,N_24204,N_24521);
and U26880 (N_26880,N_25145,N_25278);
xnor U26881 (N_26881,N_24177,N_24268);
and U26882 (N_26882,N_25377,N_24578);
nand U26883 (N_26883,N_24849,N_25470);
nor U26884 (N_26884,N_25416,N_25231);
xnor U26885 (N_26885,N_25006,N_25425);
nand U26886 (N_26886,N_25082,N_24259);
nand U26887 (N_26887,N_25255,N_24413);
xnor U26888 (N_26888,N_25339,N_24895);
or U26889 (N_26889,N_24488,N_24360);
nor U26890 (N_26890,N_24709,N_24593);
nand U26891 (N_26891,N_24526,N_24584);
or U26892 (N_26892,N_24951,N_24915);
and U26893 (N_26893,N_24840,N_25103);
xnor U26894 (N_26894,N_25194,N_24340);
nor U26895 (N_26895,N_24283,N_24829);
xnor U26896 (N_26896,N_24120,N_24421);
xnor U26897 (N_26897,N_24762,N_24838);
nor U26898 (N_26898,N_25119,N_25150);
and U26899 (N_26899,N_25322,N_24384);
and U26900 (N_26900,N_24370,N_24539);
nor U26901 (N_26901,N_24089,N_24856);
nand U26902 (N_26902,N_25239,N_24440);
xnor U26903 (N_26903,N_25200,N_25172);
and U26904 (N_26904,N_24475,N_24027);
or U26905 (N_26905,N_24712,N_24335);
nand U26906 (N_26906,N_24789,N_25378);
xor U26907 (N_26907,N_25476,N_24569);
nor U26908 (N_26908,N_25171,N_24507);
xor U26909 (N_26909,N_24168,N_24643);
or U26910 (N_26910,N_25386,N_24280);
nor U26911 (N_26911,N_24207,N_25033);
or U26912 (N_26912,N_24734,N_24255);
and U26913 (N_26913,N_24040,N_24036);
or U26914 (N_26914,N_24344,N_24439);
and U26915 (N_26915,N_25453,N_24310);
nand U26916 (N_26916,N_25343,N_25069);
or U26917 (N_26917,N_24986,N_24133);
nor U26918 (N_26918,N_25268,N_25226);
and U26919 (N_26919,N_24987,N_25124);
xnor U26920 (N_26920,N_25257,N_24561);
and U26921 (N_26921,N_24981,N_24083);
and U26922 (N_26922,N_24014,N_24862);
nand U26923 (N_26923,N_24448,N_24590);
nor U26924 (N_26924,N_24859,N_24688);
xor U26925 (N_26925,N_24214,N_25013);
nand U26926 (N_26926,N_24002,N_24228);
nand U26927 (N_26927,N_25425,N_24931);
nand U26928 (N_26928,N_24111,N_24113);
xnor U26929 (N_26929,N_24131,N_25402);
nand U26930 (N_26930,N_25118,N_25457);
or U26931 (N_26931,N_24873,N_24360);
nor U26932 (N_26932,N_25008,N_24421);
nand U26933 (N_26933,N_25250,N_24333);
and U26934 (N_26934,N_25450,N_24317);
and U26935 (N_26935,N_24456,N_24492);
nand U26936 (N_26936,N_25154,N_24053);
nand U26937 (N_26937,N_24937,N_24641);
nand U26938 (N_26938,N_24283,N_24149);
or U26939 (N_26939,N_24799,N_25266);
nand U26940 (N_26940,N_25371,N_24410);
nor U26941 (N_26941,N_24114,N_25272);
and U26942 (N_26942,N_24406,N_24504);
nor U26943 (N_26943,N_24284,N_25180);
or U26944 (N_26944,N_25158,N_24449);
nor U26945 (N_26945,N_24775,N_24491);
xor U26946 (N_26946,N_24261,N_25048);
xor U26947 (N_26947,N_25181,N_25339);
nor U26948 (N_26948,N_24471,N_24156);
nand U26949 (N_26949,N_24928,N_24441);
or U26950 (N_26950,N_24620,N_25006);
nand U26951 (N_26951,N_24113,N_24513);
and U26952 (N_26952,N_24657,N_25074);
nor U26953 (N_26953,N_24894,N_24895);
xnor U26954 (N_26954,N_24531,N_25280);
nand U26955 (N_26955,N_24928,N_24636);
and U26956 (N_26956,N_24811,N_24500);
and U26957 (N_26957,N_24125,N_25484);
and U26958 (N_26958,N_25187,N_24799);
and U26959 (N_26959,N_24346,N_25045);
and U26960 (N_26960,N_24522,N_24203);
nand U26961 (N_26961,N_24146,N_24355);
and U26962 (N_26962,N_24162,N_24741);
or U26963 (N_26963,N_24487,N_25120);
and U26964 (N_26964,N_24735,N_24744);
xnor U26965 (N_26965,N_24948,N_25326);
or U26966 (N_26966,N_25306,N_24744);
and U26967 (N_26967,N_24323,N_24175);
nand U26968 (N_26968,N_25294,N_24405);
nor U26969 (N_26969,N_24398,N_24601);
or U26970 (N_26970,N_25241,N_24144);
and U26971 (N_26971,N_24369,N_24057);
or U26972 (N_26972,N_24900,N_24091);
xor U26973 (N_26973,N_24724,N_24363);
and U26974 (N_26974,N_24746,N_25147);
nor U26975 (N_26975,N_24526,N_24966);
nand U26976 (N_26976,N_25072,N_24075);
nor U26977 (N_26977,N_24074,N_25366);
xnor U26978 (N_26978,N_25083,N_24263);
and U26979 (N_26979,N_25129,N_25325);
nand U26980 (N_26980,N_25240,N_24350);
xor U26981 (N_26981,N_25467,N_25329);
nand U26982 (N_26982,N_25152,N_24225);
nand U26983 (N_26983,N_24153,N_24831);
nand U26984 (N_26984,N_25346,N_24281);
nand U26985 (N_26985,N_25131,N_24754);
nand U26986 (N_26986,N_25133,N_24868);
nor U26987 (N_26987,N_24596,N_24063);
or U26988 (N_26988,N_24440,N_25097);
nand U26989 (N_26989,N_24470,N_24414);
nand U26990 (N_26990,N_24082,N_25193);
and U26991 (N_26991,N_24617,N_24142);
or U26992 (N_26992,N_25219,N_25087);
nor U26993 (N_26993,N_24553,N_24909);
nor U26994 (N_26994,N_24038,N_24693);
and U26995 (N_26995,N_24887,N_24177);
nor U26996 (N_26996,N_25371,N_25023);
and U26997 (N_26997,N_24346,N_24785);
nor U26998 (N_26998,N_24638,N_25159);
xor U26999 (N_26999,N_24641,N_25162);
and U27000 (N_27000,N_26863,N_26773);
xor U27001 (N_27001,N_26961,N_26458);
nor U27002 (N_27002,N_26512,N_26790);
nand U27003 (N_27003,N_26627,N_26808);
and U27004 (N_27004,N_26155,N_26399);
and U27005 (N_27005,N_25541,N_26066);
nand U27006 (N_27006,N_26491,N_26717);
or U27007 (N_27007,N_26482,N_26084);
nor U27008 (N_27008,N_26533,N_25721);
or U27009 (N_27009,N_25895,N_26093);
or U27010 (N_27010,N_26036,N_26164);
xnor U27011 (N_27011,N_25738,N_26621);
or U27012 (N_27012,N_25967,N_25976);
nor U27013 (N_27013,N_26161,N_26200);
xor U27014 (N_27014,N_26017,N_26337);
nand U27015 (N_27015,N_25821,N_25787);
or U27016 (N_27016,N_25733,N_26962);
and U27017 (N_27017,N_25992,N_26438);
nor U27018 (N_27018,N_26645,N_26068);
and U27019 (N_27019,N_26283,N_26519);
or U27020 (N_27020,N_25988,N_26543);
nor U27021 (N_27021,N_26819,N_26062);
nand U27022 (N_27022,N_25605,N_25990);
or U27023 (N_27023,N_26074,N_26174);
or U27024 (N_27024,N_26460,N_26065);
nand U27025 (N_27025,N_26432,N_26010);
xor U27026 (N_27026,N_26871,N_25994);
and U27027 (N_27027,N_26671,N_25526);
and U27028 (N_27028,N_26565,N_25513);
nand U27029 (N_27029,N_25973,N_26481);
nor U27030 (N_27030,N_26631,N_26130);
and U27031 (N_27031,N_26058,N_26247);
or U27032 (N_27032,N_26329,N_25851);
or U27033 (N_27033,N_26106,N_26461);
nor U27034 (N_27034,N_26550,N_25810);
nand U27035 (N_27035,N_26159,N_26226);
nor U27036 (N_27036,N_25584,N_25841);
or U27037 (N_27037,N_26239,N_26063);
nor U27038 (N_27038,N_26797,N_26782);
xnor U27039 (N_27039,N_25722,N_26508);
or U27040 (N_27040,N_26588,N_26404);
nand U27041 (N_27041,N_26560,N_26876);
xnor U27042 (N_27042,N_25806,N_26464);
and U27043 (N_27043,N_26196,N_26448);
and U27044 (N_27044,N_25545,N_26330);
or U27045 (N_27045,N_26986,N_26589);
nor U27046 (N_27046,N_26860,N_25788);
or U27047 (N_27047,N_26783,N_26480);
nor U27048 (N_27048,N_25752,N_26103);
or U27049 (N_27049,N_25843,N_26682);
or U27050 (N_27050,N_26271,N_26555);
or U27051 (N_27051,N_26557,N_26647);
nand U27052 (N_27052,N_26234,N_26622);
nand U27053 (N_27053,N_26223,N_26493);
nor U27054 (N_27054,N_25944,N_26218);
and U27055 (N_27055,N_25812,N_25708);
nor U27056 (N_27056,N_25522,N_25766);
xnor U27057 (N_27057,N_26840,N_26443);
and U27058 (N_27058,N_25888,N_25585);
nand U27059 (N_27059,N_26075,N_26187);
xnor U27060 (N_27060,N_26211,N_26850);
and U27061 (N_27061,N_26978,N_25739);
and U27062 (N_27062,N_26514,N_25671);
and U27063 (N_27063,N_26657,N_25934);
nand U27064 (N_27064,N_26474,N_26920);
nand U27065 (N_27065,N_25508,N_25601);
or U27066 (N_27066,N_25996,N_26270);
nand U27067 (N_27067,N_25887,N_26381);
xnor U27068 (N_27068,N_26230,N_26427);
or U27069 (N_27069,N_26041,N_25500);
nor U27070 (N_27070,N_26050,N_26167);
nand U27071 (N_27071,N_26890,N_25679);
nand U27072 (N_27072,N_26308,N_26559);
and U27073 (N_27073,N_26343,N_26774);
or U27074 (N_27074,N_25616,N_26634);
or U27075 (N_27075,N_26294,N_25893);
and U27076 (N_27076,N_26713,N_25701);
nor U27077 (N_27077,N_25564,N_26426);
or U27078 (N_27078,N_26997,N_26269);
or U27079 (N_27079,N_26140,N_25998);
xor U27080 (N_27080,N_26886,N_26618);
nand U27081 (N_27081,N_26019,N_26915);
and U27082 (N_27082,N_26542,N_26317);
nor U27083 (N_27083,N_26959,N_25657);
nor U27084 (N_27084,N_26433,N_26864);
and U27085 (N_27085,N_25754,N_26047);
nor U27086 (N_27086,N_26410,N_26267);
or U27087 (N_27087,N_25724,N_25637);
nor U27088 (N_27088,N_25875,N_26880);
nor U27089 (N_27089,N_25795,N_26984);
nor U27090 (N_27090,N_26449,N_26829);
or U27091 (N_27091,N_25838,N_26566);
nand U27092 (N_27092,N_25598,N_25702);
and U27093 (N_27093,N_25784,N_26833);
nor U27094 (N_27094,N_26729,N_26654);
or U27095 (N_27095,N_26168,N_25751);
or U27096 (N_27096,N_26600,N_26029);
and U27097 (N_27097,N_26788,N_25932);
xnor U27098 (N_27098,N_25727,N_26584);
nor U27099 (N_27099,N_25799,N_26420);
and U27100 (N_27100,N_26328,N_26652);
nor U27101 (N_27101,N_26158,N_26938);
nor U27102 (N_27102,N_25693,N_26994);
and U27103 (N_27103,N_25803,N_26007);
or U27104 (N_27104,N_26692,N_25868);
or U27105 (N_27105,N_26490,N_26623);
or U27106 (N_27106,N_25879,N_26563);
nor U27107 (N_27107,N_26082,N_26693);
nor U27108 (N_27108,N_25547,N_26506);
or U27109 (N_27109,N_26384,N_25749);
and U27110 (N_27110,N_25544,N_26614);
nand U27111 (N_27111,N_26757,N_26478);
and U27112 (N_27112,N_26660,N_26263);
and U27113 (N_27113,N_25614,N_26435);
and U27114 (N_27114,N_26043,N_26897);
and U27115 (N_27115,N_26815,N_26502);
nand U27116 (N_27116,N_26227,N_25781);
xor U27117 (N_27117,N_26677,N_26535);
or U27118 (N_27118,N_26577,N_26603);
nand U27119 (N_27119,N_26094,N_25758);
nor U27120 (N_27120,N_26455,N_25641);
or U27121 (N_27121,N_26500,N_25984);
nor U27122 (N_27122,N_26977,N_25955);
nand U27123 (N_27123,N_26666,N_26472);
nor U27124 (N_27124,N_26031,N_26607);
xor U27125 (N_27125,N_26248,N_26368);
nand U27126 (N_27126,N_25677,N_26881);
xnor U27127 (N_27127,N_26644,N_26295);
xor U27128 (N_27128,N_26112,N_26698);
and U27129 (N_27129,N_25570,N_26796);
nand U27130 (N_27130,N_25549,N_26250);
nor U27131 (N_27131,N_25891,N_26910);
or U27132 (N_27132,N_25878,N_26291);
nor U27133 (N_27133,N_25873,N_26213);
nand U27134 (N_27134,N_26090,N_26347);
nor U27135 (N_27135,N_26471,N_26628);
xnor U27136 (N_27136,N_25501,N_26632);
nor U27137 (N_27137,N_25673,N_26759);
nor U27138 (N_27138,N_25509,N_26590);
nor U27139 (N_27139,N_26616,N_25573);
xnor U27140 (N_27140,N_26470,N_26606);
and U27141 (N_27141,N_26111,N_25989);
nand U27142 (N_27142,N_25719,N_26971);
or U27143 (N_27143,N_25874,N_26691);
nand U27144 (N_27144,N_25777,N_26816);
and U27145 (N_27145,N_26516,N_26037);
or U27146 (N_27146,N_26894,N_25825);
or U27147 (N_27147,N_25774,N_25950);
nor U27148 (N_27148,N_26637,N_25577);
xor U27149 (N_27149,N_26053,N_25642);
nor U27150 (N_27150,N_25931,N_26278);
and U27151 (N_27151,N_26342,N_25904);
xnor U27152 (N_27152,N_25816,N_26099);
and U27153 (N_27153,N_26518,N_26462);
xor U27154 (N_27154,N_26624,N_26222);
or U27155 (N_27155,N_25589,N_26306);
nand U27156 (N_27156,N_25772,N_26129);
nand U27157 (N_27157,N_26497,N_26730);
nand U27158 (N_27158,N_26414,N_26353);
and U27159 (N_27159,N_26486,N_26954);
xnor U27160 (N_27160,N_25780,N_26803);
xor U27161 (N_27161,N_26804,N_26763);
nor U27162 (N_27162,N_26992,N_25889);
and U27163 (N_27163,N_26033,N_26113);
or U27164 (N_27164,N_25921,N_25713);
nand U27165 (N_27165,N_26081,N_25796);
and U27166 (N_27166,N_25668,N_26760);
and U27167 (N_27167,N_26630,N_26725);
or U27168 (N_27168,N_26909,N_25839);
xor U27169 (N_27169,N_25567,N_26030);
nor U27170 (N_27170,N_26356,N_26552);
xnor U27171 (N_27171,N_26604,N_26290);
nand U27172 (N_27172,N_26967,N_25938);
and U27173 (N_27173,N_26571,N_26018);
xor U27174 (N_27174,N_26320,N_25809);
nor U27175 (N_27175,N_25986,N_25649);
nand U27176 (N_27176,N_25746,N_26902);
and U27177 (N_27177,N_26667,N_25715);
xor U27178 (N_27178,N_25909,N_26743);
or U27179 (N_27179,N_25556,N_26219);
or U27180 (N_27180,N_25937,N_25791);
and U27181 (N_27181,N_25761,N_25652);
xor U27182 (N_27182,N_26363,N_26859);
nand U27183 (N_27183,N_26747,N_26659);
xor U27184 (N_27184,N_26020,N_26258);
xor U27185 (N_27185,N_26195,N_25995);
nand U27186 (N_27186,N_26903,N_26423);
and U27187 (N_27187,N_25737,N_26612);
xnor U27188 (N_27188,N_26649,N_26891);
or U27189 (N_27189,N_26289,N_26224);
nor U27190 (N_27190,N_26731,N_26045);
or U27191 (N_27191,N_26709,N_25852);
and U27192 (N_27192,N_26832,N_25849);
or U27193 (N_27193,N_26349,N_26704);
and U27194 (N_27194,N_26197,N_26925);
nand U27195 (N_27195,N_25854,N_26252);
or U27196 (N_27196,N_26193,N_26238);
or U27197 (N_27197,N_26888,N_26143);
nand U27198 (N_27198,N_26198,N_26051);
and U27199 (N_27199,N_26489,N_25837);
or U27200 (N_27200,N_26246,N_25593);
nand U27201 (N_27201,N_26052,N_25999);
xor U27202 (N_27202,N_26683,N_26307);
xnor U27203 (N_27203,N_26855,N_26390);
nor U27204 (N_27204,N_26408,N_26769);
nor U27205 (N_27205,N_26454,N_26153);
and U27206 (N_27206,N_26981,N_26642);
nand U27207 (N_27207,N_26044,N_25604);
xor U27208 (N_27208,N_25591,N_26078);
or U27209 (N_27209,N_25865,N_26318);
and U27210 (N_27210,N_25956,N_26596);
or U27211 (N_27211,N_26901,N_26488);
and U27212 (N_27212,N_26723,N_25606);
xor U27213 (N_27213,N_26277,N_26949);
nand U27214 (N_27214,N_26573,N_26396);
or U27215 (N_27215,N_25540,N_26753);
nor U27216 (N_27216,N_26989,N_26733);
nand U27217 (N_27217,N_25853,N_26171);
nand U27218 (N_27218,N_25624,N_26182);
and U27219 (N_27219,N_25689,N_26825);
xnor U27220 (N_27220,N_26707,N_25655);
nand U27221 (N_27221,N_26366,N_26998);
nor U27222 (N_27222,N_26067,N_25716);
xor U27223 (N_27223,N_26201,N_26857);
nand U27224 (N_27224,N_26939,N_26236);
xor U27225 (N_27225,N_26123,N_26597);
nand U27226 (N_27226,N_26787,N_25857);
xor U27227 (N_27227,N_25928,N_26706);
and U27228 (N_27228,N_25793,N_26119);
xnor U27229 (N_27229,N_26973,N_26359);
xor U27230 (N_27230,N_26749,N_26694);
or U27231 (N_27231,N_26186,N_25822);
xnor U27232 (N_27232,N_26225,N_25817);
nor U27233 (N_27233,N_26245,N_26726);
and U27234 (N_27234,N_26003,N_26549);
and U27235 (N_27235,N_26276,N_26879);
xnor U27236 (N_27236,N_26152,N_26766);
xnor U27237 (N_27237,N_26424,N_25906);
and U27238 (N_27238,N_26581,N_26385);
or U27239 (N_27239,N_26024,N_26554);
nor U27240 (N_27240,N_26892,N_26822);
nor U27241 (N_27241,N_25767,N_26340);
nand U27242 (N_27242,N_26466,N_26662);
nor U27243 (N_27243,N_26374,N_26737);
and U27244 (N_27244,N_26601,N_25523);
and U27245 (N_27245,N_25987,N_26281);
xnor U27246 (N_27246,N_26280,N_25694);
nor U27247 (N_27247,N_25610,N_25551);
nor U27248 (N_27248,N_26689,N_26511);
or U27249 (N_27249,N_26485,N_25947);
nor U27250 (N_27250,N_26180,N_25506);
xnor U27251 (N_27251,N_26445,N_25645);
and U27252 (N_27252,N_25687,N_25962);
and U27253 (N_27253,N_25706,N_26005);
xor U27254 (N_27254,N_25881,N_25820);
or U27255 (N_27255,N_26951,N_25528);
and U27256 (N_27256,N_25759,N_26847);
xnor U27257 (N_27257,N_25897,N_26015);
or U27258 (N_27258,N_26212,N_25623);
nor U27259 (N_27259,N_25900,N_26640);
nor U27260 (N_27260,N_25902,N_25804);
or U27261 (N_27261,N_25983,N_25705);
xor U27262 (N_27262,N_26137,N_26710);
nand U27263 (N_27263,N_25933,N_26653);
and U27264 (N_27264,N_25818,N_25783);
or U27265 (N_27265,N_25617,N_26964);
nor U27266 (N_27266,N_26300,N_26751);
or U27267 (N_27267,N_26836,N_26004);
nor U27268 (N_27268,N_25847,N_26096);
nand U27269 (N_27269,N_26771,N_25676);
xor U27270 (N_27270,N_25836,N_25674);
and U27271 (N_27271,N_25765,N_26389);
xor U27272 (N_27272,N_26873,N_26205);
or U27273 (N_27273,N_26952,N_26282);
and U27274 (N_27274,N_25794,N_25587);
and U27275 (N_27275,N_25845,N_25517);
or U27276 (N_27276,N_26135,N_26372);
nand U27277 (N_27277,N_26440,N_26208);
nand U27278 (N_27278,N_26673,N_25725);
and U27279 (N_27279,N_26217,N_25941);
nor U27280 (N_27280,N_26522,N_26332);
or U27281 (N_27281,N_25583,N_25621);
or U27282 (N_27282,N_26023,N_26629);
and U27283 (N_27283,N_26001,N_26398);
nor U27284 (N_27284,N_26229,N_26450);
nand U27285 (N_27285,N_26288,N_26820);
and U27286 (N_27286,N_26418,N_25886);
nor U27287 (N_27287,N_26484,N_26442);
xor U27288 (N_27288,N_25524,N_26022);
or U27289 (N_27289,N_25626,N_25916);
nand U27290 (N_27290,N_25529,N_26861);
nand U27291 (N_27291,N_26856,N_25704);
or U27292 (N_27292,N_25699,N_25553);
nand U27293 (N_27293,N_25808,N_26297);
xor U27294 (N_27294,N_26546,N_26100);
or U27295 (N_27295,N_26237,N_26403);
nor U27296 (N_27296,N_26678,N_26061);
nor U27297 (N_27297,N_25968,N_26688);
xor U27298 (N_27298,N_26166,N_26341);
nor U27299 (N_27299,N_25537,N_26108);
or U27300 (N_27300,N_26070,N_26823);
and U27301 (N_27301,N_25586,N_25964);
xor U27302 (N_27302,N_26173,N_25731);
nand U27303 (N_27303,N_25561,N_26999);
xor U27304 (N_27304,N_25557,N_26578);
or U27305 (N_27305,N_25555,N_26446);
nor U27306 (N_27306,N_25634,N_26401);
nor U27307 (N_27307,N_26179,N_25579);
and U27308 (N_27308,N_25898,N_26170);
nor U27309 (N_27309,N_25858,N_26333);
xor U27310 (N_27310,N_25832,N_26532);
xnor U27311 (N_27311,N_26987,N_25630);
or U27312 (N_27312,N_25943,N_25920);
nand U27313 (N_27313,N_26091,N_25613);
and U27314 (N_27314,N_26483,N_26839);
nand U27315 (N_27315,N_26344,N_26947);
xor U27316 (N_27316,N_26383,N_26473);
nand U27317 (N_27317,N_25978,N_26304);
xor U27318 (N_27318,N_26646,N_26206);
and U27319 (N_27319,N_26551,N_26371);
nor U27320 (N_27320,N_26346,N_25682);
or U27321 (N_27321,N_26256,N_25985);
nor U27322 (N_27322,N_25919,N_26101);
xor U27323 (N_27323,N_25778,N_26548);
or U27324 (N_27324,N_25678,N_26993);
and U27325 (N_27325,N_26088,N_25753);
nand U27326 (N_27326,N_25743,N_26085);
or U27327 (N_27327,N_26049,N_26658);
xor U27328 (N_27328,N_26807,N_25646);
or U27329 (N_27329,N_26244,N_26388);
or U27330 (N_27330,N_25681,N_26405);
and U27331 (N_27331,N_26274,N_26937);
or U27332 (N_27332,N_25571,N_26865);
nand U27333 (N_27333,N_26121,N_25504);
xnor U27334 (N_27334,N_25710,N_26927);
and U27335 (N_27335,N_26955,N_26501);
nor U27336 (N_27336,N_26800,N_26035);
nand U27337 (N_27337,N_26114,N_26918);
nor U27338 (N_27338,N_26755,N_25667);
and U27339 (N_27339,N_26721,N_26853);
and U27340 (N_27340,N_26564,N_26908);
nor U27341 (N_27341,N_26228,N_26467);
and U27342 (N_27342,N_26315,N_26866);
and U27343 (N_27343,N_26375,N_26505);
and U27344 (N_27344,N_26945,N_25882);
or U27345 (N_27345,N_26609,N_26586);
or U27346 (N_27346,N_25952,N_25647);
xor U27347 (N_27347,N_25734,N_25639);
xnor U27348 (N_27348,N_26150,N_26580);
or U27349 (N_27349,N_26625,N_25763);
or U27350 (N_27350,N_25692,N_26996);
or U27351 (N_27351,N_26459,N_26127);
nand U27352 (N_27352,N_25911,N_26702);
xnor U27353 (N_27353,N_25776,N_26812);
nor U27354 (N_27354,N_26963,N_25607);
and U27355 (N_27355,N_26917,N_26750);
xor U27356 (N_27356,N_26331,N_26313);
xor U27357 (N_27357,N_26525,N_25914);
xor U27358 (N_27358,N_26011,N_25627);
xnor U27359 (N_27359,N_26160,N_25756);
or U27360 (N_27360,N_26469,N_26188);
nor U27361 (N_27361,N_26380,N_26770);
or U27362 (N_27362,N_26190,N_25855);
xnor U27363 (N_27363,N_26727,N_25519);
nand U27364 (N_27364,N_26758,N_25558);
and U27365 (N_27365,N_26793,N_26008);
xnor U27366 (N_27366,N_26715,N_26303);
or U27367 (N_27367,N_26293,N_25927);
nor U27368 (N_27368,N_26817,N_26744);
xor U27369 (N_27369,N_26038,N_25801);
and U27370 (N_27370,N_26496,N_25939);
xor U27371 (N_27371,N_26568,N_26779);
or U27372 (N_27372,N_25636,N_26844);
xor U27373 (N_27373,N_26794,N_25867);
and U27374 (N_27374,N_26570,N_26145);
nand U27375 (N_27375,N_26422,N_25755);
and U27376 (N_27376,N_26437,N_26386);
and U27377 (N_27377,N_26379,N_26921);
and U27378 (N_27378,N_25594,N_26738);
nand U27379 (N_27379,N_26169,N_25930);
nand U27380 (N_27380,N_26620,N_26456);
and U27381 (N_27381,N_26933,N_26275);
nand U27382 (N_27382,N_26444,N_25535);
and U27383 (N_27383,N_25883,N_25741);
nor U27384 (N_27384,N_25521,N_26569);
and U27385 (N_27385,N_26765,N_26089);
nand U27386 (N_27386,N_26305,N_25814);
or U27387 (N_27387,N_26686,N_26358);
nor U27388 (N_27388,N_25953,N_26762);
and U27389 (N_27389,N_26463,N_26072);
nand U27390 (N_27390,N_25805,N_26394);
and U27391 (N_27391,N_25894,N_26656);
nand U27392 (N_27392,N_26064,N_25936);
nor U27393 (N_27393,N_26869,N_25569);
nand U27394 (N_27394,N_25903,N_25792);
and U27395 (N_27395,N_25745,N_26465);
xnor U27396 (N_27396,N_26830,N_25546);
nor U27397 (N_27397,N_26811,N_25518);
xnor U27398 (N_27398,N_26336,N_26536);
nand U27399 (N_27399,N_25660,N_26574);
nand U27400 (N_27400,N_26599,N_25856);
nand U27401 (N_27401,N_25982,N_26348);
and U27402 (N_27402,N_26835,N_25663);
xor U27403 (N_27403,N_26781,N_26468);
or U27404 (N_27404,N_26255,N_25760);
nand U27405 (N_27405,N_25729,N_25797);
nand U27406 (N_27406,N_26273,N_25884);
nor U27407 (N_27407,N_26364,N_26287);
and U27408 (N_27408,N_26314,N_26665);
or U27409 (N_27409,N_26360,N_26818);
nand U27410 (N_27410,N_26447,N_26395);
nor U27411 (N_27411,N_26675,N_26932);
xor U27412 (N_27412,N_25935,N_26350);
and U27413 (N_27413,N_26935,N_25538);
xnor U27414 (N_27414,N_26133,N_26365);
nand U27415 (N_27415,N_26705,N_25568);
xor U27416 (N_27416,N_25644,N_26409);
xnor U27417 (N_27417,N_26400,N_25951);
nand U27418 (N_27418,N_26016,N_26587);
and U27419 (N_27419,N_25785,N_26428);
or U27420 (N_27420,N_25876,N_26777);
and U27421 (N_27421,N_25665,N_26235);
xor U27422 (N_27422,N_25769,N_25807);
and U27423 (N_27423,N_26028,N_26210);
xor U27424 (N_27424,N_26528,N_26583);
and U27425 (N_27425,N_26392,N_26724);
and U27426 (N_27426,N_25740,N_25516);
and U27427 (N_27427,N_26824,N_26610);
xnor U27428 (N_27428,N_26434,N_26185);
xnor U27429 (N_27429,N_25732,N_26714);
xnor U27430 (N_27430,N_26792,N_26681);
or U27431 (N_27431,N_26872,N_26527);
nor U27432 (N_27432,N_26887,N_26849);
or U27433 (N_27433,N_26547,N_26509);
nor U27434 (N_27434,N_26006,N_26115);
xor U27435 (N_27435,N_25707,N_26175);
nor U27436 (N_27436,N_26026,N_26151);
nand U27437 (N_27437,N_26700,N_26699);
and U27438 (N_27438,N_25861,N_26253);
nand U27439 (N_27439,N_25625,N_26785);
nand U27440 (N_27440,N_26896,N_26057);
xor U27441 (N_27441,N_26407,N_26838);
xor U27442 (N_27442,N_26608,N_25828);
and U27443 (N_27443,N_25975,N_25515);
xor U27444 (N_27444,N_26795,N_25844);
xnor U27445 (N_27445,N_26079,N_26870);
xor U27446 (N_27446,N_26900,N_26696);
and U27447 (N_27447,N_26761,N_26852);
nor U27448 (N_27448,N_25829,N_26821);
xor U27449 (N_27449,N_26541,N_26635);
nand U27450 (N_27450,N_25550,N_26641);
or U27451 (N_27451,N_26284,N_25714);
or U27452 (N_27452,N_26882,N_25831);
xnor U27453 (N_27453,N_26183,N_26943);
nor U27454 (N_27454,N_26097,N_26056);
nand U27455 (N_27455,N_26534,N_25654);
nor U27456 (N_27456,N_26837,N_26980);
and U27457 (N_27457,N_26791,N_26138);
xor U27458 (N_27458,N_26338,N_26039);
nor U27459 (N_27459,N_25723,N_25862);
xor U27460 (N_27460,N_26524,N_26054);
nor U27461 (N_27461,N_25698,N_26266);
xnor U27462 (N_27462,N_25747,N_26249);
and U27463 (N_27463,N_25826,N_26867);
or U27464 (N_27464,N_26476,N_26638);
or U27465 (N_27465,N_26286,N_26012);
nor U27466 (N_27466,N_26736,N_25926);
or U27467 (N_27467,N_26452,N_25672);
and U27468 (N_27468,N_26076,N_25802);
nor U27469 (N_27469,N_25533,N_26576);
or U27470 (N_27470,N_26327,N_26177);
or U27471 (N_27471,N_26260,N_25525);
xnor U27472 (N_27472,N_26789,N_25859);
nor U27473 (N_27473,N_25910,N_25590);
or U27474 (N_27474,N_25790,N_26369);
and U27475 (N_27475,N_26352,N_26953);
or U27476 (N_27476,N_26846,N_25742);
nor U27477 (N_27477,N_26778,N_26391);
xor U27478 (N_27478,N_26968,N_26194);
and U27479 (N_27479,N_26421,N_26265);
or U27480 (N_27480,N_25581,N_26719);
xor U27481 (N_27481,N_25997,N_26430);
or U27482 (N_27482,N_26134,N_25991);
xor U27483 (N_27483,N_26802,N_26132);
nand U27484 (N_27484,N_26301,N_25680);
nor U27485 (N_27485,N_25896,N_25924);
xnor U27486 (N_27486,N_26916,N_26988);
nand U27487 (N_27487,N_26745,N_26436);
nor U27488 (N_27488,N_26475,N_26602);
nor U27489 (N_27489,N_26156,N_26148);
nand U27490 (N_27490,N_26655,N_26595);
nand U27491 (N_27491,N_25726,N_26221);
nor U27492 (N_27492,N_25736,N_26189);
xor U27493 (N_27493,N_25675,N_26545);
nand U27494 (N_27494,N_26663,N_26122);
nor U27495 (N_27495,N_25744,N_26083);
or U27496 (N_27496,N_25664,N_26387);
nor U27497 (N_27497,N_26685,N_26095);
and U27498 (N_27498,N_26191,N_26510);
and U27499 (N_27499,N_26172,N_25503);
xor U27500 (N_27500,N_26046,N_26069);
nor U27501 (N_27501,N_25915,N_26739);
and U27502 (N_27502,N_25596,N_25912);
and U27503 (N_27503,N_25942,N_26339);
nor U27504 (N_27504,N_26826,N_25728);
or U27505 (N_27505,N_26009,N_25768);
or U27506 (N_27506,N_26411,N_26639);
nand U27507 (N_27507,N_26862,N_26799);
xnor U27508 (N_27508,N_26141,N_26325);
xnor U27509 (N_27509,N_25574,N_26254);
xnor U27510 (N_27510,N_25566,N_26136);
nand U27511 (N_27511,N_26507,N_26711);
nand U27512 (N_27512,N_26854,N_26615);
nand U27513 (N_27513,N_26124,N_25971);
nand U27514 (N_27514,N_25830,N_26810);
xnor U27515 (N_27515,N_25863,N_25824);
nand U27516 (N_27516,N_26354,N_25612);
or U27517 (N_27517,N_25977,N_25658);
xnor U27518 (N_27518,N_25542,N_26257);
nor U27519 (N_27519,N_26128,N_26165);
and U27520 (N_27520,N_26941,N_25530);
or U27521 (N_27521,N_26319,N_25548);
or U27522 (N_27522,N_26928,N_26684);
or U27523 (N_27523,N_26285,N_26526);
nand U27524 (N_27524,N_25502,N_26242);
xor U27525 (N_27525,N_25922,N_26415);
or U27526 (N_27526,N_26416,N_26633);
and U27527 (N_27527,N_25963,N_25835);
xor U27528 (N_27528,N_26537,N_26268);
nand U27529 (N_27529,N_26334,N_26441);
or U27530 (N_27530,N_26157,N_26429);
or U27531 (N_27531,N_26930,N_26716);
xor U27532 (N_27532,N_26674,N_25543);
xor U27533 (N_27533,N_26431,N_25560);
nand U27534 (N_27534,N_26740,N_26178);
nor U27535 (N_27535,N_25779,N_25592);
and U27536 (N_27536,N_26784,N_25615);
xor U27537 (N_27537,N_26889,N_26139);
xnor U27538 (N_27538,N_26969,N_26021);
nand U27539 (N_27539,N_26000,N_26617);
nand U27540 (N_27540,N_26377,N_26233);
nor U27541 (N_27541,N_25510,N_26302);
nand U27542 (N_27542,N_26071,N_26042);
or U27543 (N_27543,N_25718,N_26417);
nand U27544 (N_27544,N_26561,N_26335);
nand U27545 (N_27545,N_26923,N_25532);
or U27546 (N_27546,N_26110,N_26858);
nor U27547 (N_27547,N_26934,N_26643);
nor U27548 (N_27548,N_26664,N_26105);
and U27549 (N_27549,N_25929,N_26752);
nor U27550 (N_27550,N_25575,N_26979);
and U27551 (N_27551,N_25949,N_26048);
nor U27552 (N_27552,N_26439,N_26912);
or U27553 (N_27553,N_26402,N_25552);
and U27554 (N_27554,N_26697,N_25842);
nand U27555 (N_27555,N_25913,N_26966);
nor U27556 (N_27556,N_25582,N_26118);
nand U27557 (N_27557,N_26517,N_26741);
and U27558 (N_27558,N_26492,N_26911);
and U27559 (N_27559,N_26776,N_25599);
or U27560 (N_27560,N_26523,N_25860);
nand U27561 (N_27561,N_26885,N_26220);
and U27562 (N_27562,N_25730,N_26529);
and U27563 (N_27563,N_25823,N_25981);
nand U27564 (N_27564,N_26243,N_25620);
nor U27565 (N_27565,N_25534,N_25846);
nor U27566 (N_27566,N_25762,N_26544);
xor U27567 (N_27567,N_25632,N_26530);
nor U27568 (N_27568,N_26868,N_26669);
nor U27569 (N_27569,N_25650,N_25940);
and U27570 (N_27570,N_26376,N_25628);
nor U27571 (N_27571,N_26619,N_25735);
and U27572 (N_27572,N_26585,N_25640);
nand U27573 (N_27573,N_26990,N_25597);
or U27574 (N_27574,N_26690,N_26922);
xnor U27575 (N_27575,N_26251,N_25562);
xnor U27576 (N_27576,N_25565,N_26592);
nand U27577 (N_27577,N_25771,N_25685);
nor U27578 (N_27578,N_25611,N_26775);
and U27579 (N_27579,N_25960,N_25866);
nor U27580 (N_27580,N_25869,N_26742);
nor U27581 (N_27581,N_25833,N_26264);
nor U27582 (N_27582,N_26214,N_25789);
or U27583 (N_27583,N_26960,N_26362);
nand U27584 (N_27584,N_26893,N_25595);
xnor U27585 (N_27585,N_26014,N_25864);
and U27586 (N_27586,N_26991,N_25905);
and U27587 (N_27587,N_26087,N_26513);
nand U27588 (N_27588,N_26926,N_26034);
nand U27589 (N_27589,N_26184,N_26809);
xor U27590 (N_27590,N_25661,N_26131);
xor U27591 (N_27591,N_26919,N_26805);
nor U27592 (N_27592,N_26668,N_26983);
or U27593 (N_27593,N_26451,N_25505);
nor U27594 (N_27594,N_25653,N_26754);
nand U27595 (N_27595,N_25899,N_26125);
xnor U27596 (N_27596,N_26950,N_26648);
nand U27597 (N_27597,N_25656,N_26357);
xor U27598 (N_27598,N_25850,N_26748);
nor U27599 (N_27599,N_26322,N_26708);
nor U27600 (N_27600,N_26240,N_25827);
xnor U27601 (N_27601,N_26806,N_25619);
nor U27602 (N_27602,N_26878,N_26831);
and U27603 (N_27603,N_26843,N_26553);
xor U27604 (N_27604,N_25923,N_25559);
or U27605 (N_27605,N_25834,N_26453);
or U27606 (N_27606,N_25918,N_26216);
or U27607 (N_27607,N_25697,N_26494);
nor U27608 (N_27608,N_26680,N_26572);
nor U27609 (N_27609,N_26279,N_26126);
nor U27610 (N_27610,N_26558,N_26904);
nor U27611 (N_27611,N_26055,N_26098);
nor U27612 (N_27612,N_26974,N_26147);
and U27613 (N_27613,N_26813,N_26734);
nor U27614 (N_27614,N_25507,N_26232);
nand U27615 (N_27615,N_26732,N_26636);
or U27616 (N_27616,N_26701,N_26413);
or U27617 (N_27617,N_26370,N_25819);
xnor U27618 (N_27618,N_26695,N_25871);
nor U27619 (N_27619,N_26845,N_26102);
nor U27620 (N_27620,N_26531,N_26499);
xnor U27621 (N_27621,N_25958,N_26323);
xor U27622 (N_27622,N_25800,N_25974);
or U27623 (N_27623,N_25690,N_26582);
or U27624 (N_27624,N_26940,N_26116);
nor U27625 (N_27625,N_25946,N_26798);
or U27626 (N_27626,N_26907,N_25603);
or U27627 (N_27627,N_25782,N_26828);
xnor U27628 (N_27628,N_25638,N_26146);
nor U27629 (N_27629,N_25578,N_26109);
xor U27630 (N_27630,N_26670,N_25892);
and U27631 (N_27631,N_25662,N_25972);
and U27632 (N_27632,N_25954,N_26942);
or U27633 (N_27633,N_26722,N_26746);
or U27634 (N_27634,N_26931,N_26027);
or U27635 (N_27635,N_26367,N_26120);
xnor U27636 (N_27636,N_26965,N_26487);
and U27637 (N_27637,N_26594,N_26672);
xnor U27638 (N_27638,N_26593,N_25907);
or U27639 (N_27639,N_26884,N_26906);
nor U27640 (N_27640,N_25980,N_26204);
or U27641 (N_27641,N_26520,N_26479);
xor U27642 (N_27642,N_25748,N_25683);
nand U27643 (N_27643,N_26355,N_26199);
or U27644 (N_27644,N_25651,N_26877);
nor U27645 (N_27645,N_26958,N_26162);
xnor U27646 (N_27646,N_25877,N_26786);
nand U27647 (N_27647,N_26948,N_26207);
or U27648 (N_27648,N_26539,N_26149);
and U27649 (N_27649,N_26834,N_25720);
xor U27650 (N_27650,N_26025,N_25688);
nand U27651 (N_27651,N_26827,N_25959);
and U27652 (N_27652,N_26687,N_26540);
nor U27653 (N_27653,N_26626,N_25512);
nor U27654 (N_27654,N_26425,N_26324);
or U27655 (N_27655,N_26202,N_25608);
nand U27656 (N_27656,N_26203,N_26875);
nand U27657 (N_27657,N_25712,N_26077);
nand U27658 (N_27658,N_25629,N_26905);
or U27659 (N_27659,N_26598,N_26914);
and U27660 (N_27660,N_26326,N_25890);
nand U27661 (N_27661,N_25580,N_26259);
nor U27662 (N_27662,N_25703,N_26117);
nand U27663 (N_27663,N_26261,N_25917);
or U27664 (N_27664,N_25514,N_26567);
nand U27665 (N_27665,N_26515,N_26215);
and U27666 (N_27666,N_25643,N_26144);
and U27667 (N_27667,N_26913,N_26312);
or U27668 (N_27668,N_26676,N_25750);
nand U27669 (N_27669,N_26382,N_25993);
nor U27670 (N_27670,N_26929,N_26412);
xor U27671 (N_27671,N_26316,N_25901);
nand U27672 (N_27672,N_26092,N_26720);
nand U27673 (N_27673,N_26104,N_26899);
and U27674 (N_27674,N_25670,N_26457);
or U27675 (N_27675,N_26651,N_25609);
or U27676 (N_27676,N_26995,N_26107);
and U27677 (N_27677,N_26764,N_26477);
or U27678 (N_27678,N_26562,N_25957);
nand U27679 (N_27679,N_25848,N_26898);
and U27680 (N_27680,N_26851,N_25631);
xnor U27681 (N_27681,N_26296,N_26591);
nand U27682 (N_27682,N_26060,N_26361);
nor U27683 (N_27683,N_26503,N_26406);
xor U27684 (N_27684,N_25572,N_26613);
nand U27685 (N_27685,N_26397,N_26373);
or U27686 (N_27686,N_25717,N_26002);
or U27687 (N_27687,N_26073,N_26801);
nand U27688 (N_27688,N_25511,N_26605);
nand U27689 (N_27689,N_25669,N_26780);
nand U27690 (N_27690,N_26814,N_25798);
or U27691 (N_27691,N_25945,N_26756);
and U27692 (N_27692,N_26735,N_26956);
xnor U27693 (N_27693,N_26298,N_26946);
nand U27694 (N_27694,N_26728,N_26718);
xor U27695 (N_27695,N_26504,N_26086);
nor U27696 (N_27696,N_26985,N_26378);
nor U27697 (N_27697,N_26059,N_26498);
nand U27698 (N_27698,N_26679,N_26351);
nand U27699 (N_27699,N_26768,N_26772);
nor U27700 (N_27700,N_26703,N_25786);
nor U27701 (N_27701,N_25635,N_26040);
nand U27702 (N_27702,N_25840,N_26241);
nor U27703 (N_27703,N_26538,N_26848);
nor U27704 (N_27704,N_26311,N_26176);
or U27705 (N_27705,N_25961,N_25588);
or U27706 (N_27706,N_25666,N_26192);
and U27707 (N_27707,N_26767,N_25554);
or U27708 (N_27708,N_26976,N_26982);
nor U27709 (N_27709,N_25539,N_26924);
or U27710 (N_27710,N_25602,N_25618);
xnor U27711 (N_27711,N_26841,N_25686);
or U27712 (N_27712,N_25691,N_26321);
nor U27713 (N_27713,N_25966,N_26895);
nor U27714 (N_27714,N_26299,N_26393);
nand U27715 (N_27715,N_26661,N_26495);
and U27716 (N_27716,N_25969,N_25520);
and U27717 (N_27717,N_26310,N_25885);
nor U27718 (N_27718,N_26975,N_26874);
and U27719 (N_27719,N_25757,N_26309);
and U27720 (N_27720,N_25813,N_25925);
nor U27721 (N_27721,N_25536,N_26154);
xor U27722 (N_27722,N_25870,N_25908);
and U27723 (N_27723,N_25648,N_25711);
xor U27724 (N_27724,N_26957,N_25696);
and U27725 (N_27725,N_26575,N_25948);
and U27726 (N_27726,N_25563,N_25576);
xor U27727 (N_27727,N_25770,N_25622);
xor U27728 (N_27728,N_26883,N_26611);
and U27729 (N_27729,N_26080,N_26013);
nor U27730 (N_27730,N_26032,N_26944);
and U27731 (N_27731,N_25775,N_25633);
and U27732 (N_27732,N_26209,N_26972);
nand U27733 (N_27733,N_26521,N_26142);
nor U27734 (N_27734,N_26579,N_25880);
or U27735 (N_27735,N_25527,N_25709);
xor U27736 (N_27736,N_25815,N_26272);
xor U27737 (N_27737,N_26712,N_26345);
nor U27738 (N_27738,N_25979,N_26556);
xor U27739 (N_27739,N_26419,N_25764);
xor U27740 (N_27740,N_25773,N_25695);
and U27741 (N_27741,N_26650,N_26181);
nand U27742 (N_27742,N_26262,N_25700);
nand U27743 (N_27743,N_25684,N_26163);
or U27744 (N_27744,N_26292,N_25872);
or U27745 (N_27745,N_26936,N_25659);
and U27746 (N_27746,N_25965,N_25600);
and U27747 (N_27747,N_26231,N_25970);
nor U27748 (N_27748,N_26842,N_25531);
xnor U27749 (N_27749,N_25811,N_26970);
and U27750 (N_27750,N_25859,N_26324);
xor U27751 (N_27751,N_26235,N_26905);
and U27752 (N_27752,N_26271,N_26095);
nand U27753 (N_27753,N_26696,N_26015);
or U27754 (N_27754,N_25808,N_26835);
xor U27755 (N_27755,N_25559,N_26940);
or U27756 (N_27756,N_26320,N_26097);
and U27757 (N_27757,N_26516,N_26669);
nand U27758 (N_27758,N_26179,N_25616);
or U27759 (N_27759,N_26307,N_26733);
xnor U27760 (N_27760,N_25652,N_26383);
nand U27761 (N_27761,N_26311,N_26128);
or U27762 (N_27762,N_26456,N_26668);
xor U27763 (N_27763,N_25765,N_25611);
nor U27764 (N_27764,N_26143,N_26785);
nor U27765 (N_27765,N_25720,N_25813);
nand U27766 (N_27766,N_25725,N_26542);
xor U27767 (N_27767,N_26058,N_26841);
xnor U27768 (N_27768,N_26560,N_26520);
or U27769 (N_27769,N_26652,N_25602);
xor U27770 (N_27770,N_26411,N_26486);
nor U27771 (N_27771,N_26261,N_26367);
nor U27772 (N_27772,N_25910,N_25634);
xnor U27773 (N_27773,N_26657,N_26380);
nand U27774 (N_27774,N_26582,N_26786);
nor U27775 (N_27775,N_26738,N_26417);
nand U27776 (N_27776,N_26904,N_26456);
nand U27777 (N_27777,N_25757,N_26136);
or U27778 (N_27778,N_26568,N_26523);
xor U27779 (N_27779,N_26901,N_26717);
nand U27780 (N_27780,N_26972,N_26179);
nand U27781 (N_27781,N_25887,N_25878);
nand U27782 (N_27782,N_25526,N_26038);
or U27783 (N_27783,N_26962,N_26947);
xnor U27784 (N_27784,N_25805,N_26995);
xor U27785 (N_27785,N_26517,N_26721);
nand U27786 (N_27786,N_26739,N_26342);
xnor U27787 (N_27787,N_26966,N_26618);
or U27788 (N_27788,N_25869,N_26368);
and U27789 (N_27789,N_26878,N_26294);
or U27790 (N_27790,N_26920,N_26478);
nand U27791 (N_27791,N_25666,N_26634);
xnor U27792 (N_27792,N_25837,N_26244);
and U27793 (N_27793,N_26693,N_26969);
and U27794 (N_27794,N_25524,N_26815);
nor U27795 (N_27795,N_26773,N_26388);
or U27796 (N_27796,N_26624,N_26288);
nor U27797 (N_27797,N_25797,N_25662);
nand U27798 (N_27798,N_26305,N_26811);
xnor U27799 (N_27799,N_26167,N_26193);
nor U27800 (N_27800,N_25663,N_26328);
nor U27801 (N_27801,N_26657,N_26155);
nand U27802 (N_27802,N_26166,N_25836);
or U27803 (N_27803,N_26046,N_26862);
nor U27804 (N_27804,N_26900,N_26258);
and U27805 (N_27805,N_26736,N_25518);
nand U27806 (N_27806,N_25636,N_26037);
and U27807 (N_27807,N_26388,N_26827);
nor U27808 (N_27808,N_26052,N_25765);
or U27809 (N_27809,N_25853,N_25502);
or U27810 (N_27810,N_26245,N_26531);
nor U27811 (N_27811,N_26777,N_26907);
and U27812 (N_27812,N_26049,N_26030);
nor U27813 (N_27813,N_26371,N_26115);
and U27814 (N_27814,N_26609,N_25829);
xor U27815 (N_27815,N_26721,N_26501);
nor U27816 (N_27816,N_26197,N_26905);
xor U27817 (N_27817,N_26308,N_26896);
and U27818 (N_27818,N_26123,N_26677);
nand U27819 (N_27819,N_26971,N_25944);
xor U27820 (N_27820,N_26614,N_26876);
and U27821 (N_27821,N_26626,N_26712);
and U27822 (N_27822,N_26543,N_25592);
and U27823 (N_27823,N_26790,N_25999);
and U27824 (N_27824,N_25765,N_26095);
nand U27825 (N_27825,N_26714,N_26009);
or U27826 (N_27826,N_25992,N_26973);
xnor U27827 (N_27827,N_25943,N_25818);
xor U27828 (N_27828,N_26302,N_26251);
xnor U27829 (N_27829,N_25674,N_26137);
or U27830 (N_27830,N_26687,N_26785);
xnor U27831 (N_27831,N_25566,N_26058);
nand U27832 (N_27832,N_25895,N_25675);
nand U27833 (N_27833,N_26061,N_26151);
or U27834 (N_27834,N_26771,N_25692);
or U27835 (N_27835,N_25520,N_25883);
nor U27836 (N_27836,N_26017,N_26696);
nand U27837 (N_27837,N_25924,N_26015);
and U27838 (N_27838,N_26698,N_26273);
and U27839 (N_27839,N_26193,N_26405);
or U27840 (N_27840,N_26325,N_26584);
or U27841 (N_27841,N_26526,N_26947);
xor U27842 (N_27842,N_26267,N_26764);
and U27843 (N_27843,N_25615,N_25992);
nand U27844 (N_27844,N_26953,N_25863);
and U27845 (N_27845,N_26104,N_25694);
and U27846 (N_27846,N_26606,N_26212);
nor U27847 (N_27847,N_26788,N_26415);
and U27848 (N_27848,N_26807,N_26645);
or U27849 (N_27849,N_25819,N_25968);
and U27850 (N_27850,N_25778,N_25766);
or U27851 (N_27851,N_25719,N_25791);
nor U27852 (N_27852,N_26889,N_26325);
nand U27853 (N_27853,N_26068,N_25842);
nor U27854 (N_27854,N_26636,N_26635);
or U27855 (N_27855,N_26196,N_26302);
or U27856 (N_27856,N_26928,N_25505);
xor U27857 (N_27857,N_25500,N_26158);
or U27858 (N_27858,N_26911,N_26083);
xnor U27859 (N_27859,N_26659,N_26654);
and U27860 (N_27860,N_26716,N_25765);
or U27861 (N_27861,N_26554,N_26972);
nor U27862 (N_27862,N_25877,N_26634);
xor U27863 (N_27863,N_26160,N_26858);
and U27864 (N_27864,N_26028,N_25734);
xnor U27865 (N_27865,N_25762,N_26105);
and U27866 (N_27866,N_25822,N_25856);
or U27867 (N_27867,N_26614,N_26470);
or U27868 (N_27868,N_26542,N_26801);
nand U27869 (N_27869,N_26608,N_26712);
and U27870 (N_27870,N_26444,N_26966);
xnor U27871 (N_27871,N_25802,N_26897);
xor U27872 (N_27872,N_25837,N_25993);
or U27873 (N_27873,N_26800,N_25997);
nand U27874 (N_27874,N_25998,N_26874);
xnor U27875 (N_27875,N_25555,N_26904);
xnor U27876 (N_27876,N_26872,N_25554);
xor U27877 (N_27877,N_26738,N_26196);
nand U27878 (N_27878,N_26853,N_25769);
nand U27879 (N_27879,N_26563,N_26606);
xnor U27880 (N_27880,N_26810,N_25630);
xnor U27881 (N_27881,N_25872,N_26265);
and U27882 (N_27882,N_26883,N_26654);
nor U27883 (N_27883,N_26802,N_25748);
nand U27884 (N_27884,N_25675,N_26998);
nand U27885 (N_27885,N_25914,N_26971);
or U27886 (N_27886,N_26798,N_26143);
nor U27887 (N_27887,N_26790,N_25549);
nand U27888 (N_27888,N_25788,N_26352);
and U27889 (N_27889,N_26243,N_25971);
xor U27890 (N_27890,N_26472,N_25760);
or U27891 (N_27891,N_25935,N_26649);
xnor U27892 (N_27892,N_26714,N_26405);
or U27893 (N_27893,N_25780,N_25892);
or U27894 (N_27894,N_26922,N_26594);
nand U27895 (N_27895,N_25959,N_25883);
or U27896 (N_27896,N_26078,N_25783);
or U27897 (N_27897,N_26551,N_26262);
or U27898 (N_27898,N_25768,N_26323);
nand U27899 (N_27899,N_26270,N_26554);
and U27900 (N_27900,N_26981,N_25804);
nor U27901 (N_27901,N_26921,N_26246);
xnor U27902 (N_27902,N_25838,N_25826);
and U27903 (N_27903,N_26152,N_26052);
nor U27904 (N_27904,N_26143,N_25757);
xnor U27905 (N_27905,N_26545,N_26749);
xnor U27906 (N_27906,N_25729,N_26749);
or U27907 (N_27907,N_25525,N_25568);
nor U27908 (N_27908,N_25557,N_25636);
nand U27909 (N_27909,N_25833,N_26098);
or U27910 (N_27910,N_25631,N_26574);
and U27911 (N_27911,N_25653,N_26384);
or U27912 (N_27912,N_26394,N_26645);
or U27913 (N_27913,N_25748,N_26722);
or U27914 (N_27914,N_26436,N_26792);
or U27915 (N_27915,N_26648,N_26982);
nor U27916 (N_27916,N_26412,N_26330);
nor U27917 (N_27917,N_26300,N_25602);
nor U27918 (N_27918,N_26141,N_25783);
nor U27919 (N_27919,N_26640,N_25676);
and U27920 (N_27920,N_26881,N_26491);
or U27921 (N_27921,N_26339,N_26828);
and U27922 (N_27922,N_26060,N_26624);
and U27923 (N_27923,N_26873,N_25563);
nor U27924 (N_27924,N_26527,N_26542);
and U27925 (N_27925,N_26879,N_25597);
and U27926 (N_27926,N_26780,N_26696);
xnor U27927 (N_27927,N_26821,N_26276);
nor U27928 (N_27928,N_26707,N_26650);
nand U27929 (N_27929,N_25989,N_26513);
or U27930 (N_27930,N_26825,N_26017);
nand U27931 (N_27931,N_26083,N_26617);
nand U27932 (N_27932,N_25979,N_25665);
xnor U27933 (N_27933,N_26446,N_26103);
or U27934 (N_27934,N_25890,N_26563);
nand U27935 (N_27935,N_25966,N_26719);
and U27936 (N_27936,N_26415,N_25923);
or U27937 (N_27937,N_26091,N_25545);
nand U27938 (N_27938,N_26440,N_26275);
nor U27939 (N_27939,N_25747,N_25749);
xor U27940 (N_27940,N_25519,N_25626);
nand U27941 (N_27941,N_26646,N_25981);
xor U27942 (N_27942,N_25564,N_25933);
nor U27943 (N_27943,N_25816,N_25691);
nor U27944 (N_27944,N_25739,N_25651);
nand U27945 (N_27945,N_26404,N_25978);
or U27946 (N_27946,N_25645,N_26425);
or U27947 (N_27947,N_26331,N_26354);
or U27948 (N_27948,N_25774,N_25670);
xnor U27949 (N_27949,N_26814,N_26083);
and U27950 (N_27950,N_26896,N_26746);
and U27951 (N_27951,N_25694,N_26246);
nor U27952 (N_27952,N_26898,N_25554);
and U27953 (N_27953,N_26773,N_26648);
nand U27954 (N_27954,N_26835,N_26923);
nand U27955 (N_27955,N_26519,N_25536);
or U27956 (N_27956,N_25837,N_26617);
nand U27957 (N_27957,N_26231,N_26349);
and U27958 (N_27958,N_26105,N_26394);
nand U27959 (N_27959,N_26459,N_26091);
and U27960 (N_27960,N_26896,N_26865);
and U27961 (N_27961,N_26026,N_25520);
nand U27962 (N_27962,N_26219,N_25888);
nor U27963 (N_27963,N_26492,N_26294);
xor U27964 (N_27964,N_26557,N_26232);
nand U27965 (N_27965,N_25547,N_26806);
nor U27966 (N_27966,N_26605,N_26277);
nand U27967 (N_27967,N_26707,N_26439);
and U27968 (N_27968,N_26378,N_25506);
xnor U27969 (N_27969,N_25585,N_25500);
or U27970 (N_27970,N_26205,N_25598);
or U27971 (N_27971,N_26286,N_26607);
or U27972 (N_27972,N_25505,N_25756);
xnor U27973 (N_27973,N_26485,N_26613);
nand U27974 (N_27974,N_26560,N_26273);
or U27975 (N_27975,N_26022,N_25844);
xor U27976 (N_27976,N_26554,N_25500);
or U27977 (N_27977,N_26101,N_26392);
and U27978 (N_27978,N_26772,N_26919);
nor U27979 (N_27979,N_26201,N_26835);
nand U27980 (N_27980,N_25805,N_26607);
nand U27981 (N_27981,N_25805,N_26668);
xnor U27982 (N_27982,N_25809,N_26020);
xor U27983 (N_27983,N_26218,N_26395);
xor U27984 (N_27984,N_26307,N_26570);
nor U27985 (N_27985,N_25747,N_26245);
nand U27986 (N_27986,N_26530,N_26616);
or U27987 (N_27987,N_26634,N_26992);
or U27988 (N_27988,N_26382,N_26449);
nor U27989 (N_27989,N_26424,N_26959);
or U27990 (N_27990,N_26906,N_25631);
or U27991 (N_27991,N_25943,N_25667);
and U27992 (N_27992,N_26804,N_26109);
nand U27993 (N_27993,N_26196,N_26093);
nand U27994 (N_27994,N_25793,N_25763);
or U27995 (N_27995,N_25865,N_25861);
xnor U27996 (N_27996,N_25718,N_26032);
xnor U27997 (N_27997,N_26651,N_26337);
nand U27998 (N_27998,N_25761,N_26411);
or U27999 (N_27999,N_26442,N_26098);
nor U28000 (N_28000,N_25654,N_26653);
and U28001 (N_28001,N_26160,N_26562);
and U28002 (N_28002,N_25985,N_25708);
xor U28003 (N_28003,N_25624,N_26721);
or U28004 (N_28004,N_26976,N_26888);
or U28005 (N_28005,N_26679,N_26058);
or U28006 (N_28006,N_26145,N_26494);
xnor U28007 (N_28007,N_25844,N_25693);
and U28008 (N_28008,N_26248,N_25628);
nor U28009 (N_28009,N_26739,N_26484);
and U28010 (N_28010,N_26473,N_26504);
or U28011 (N_28011,N_25712,N_26742);
or U28012 (N_28012,N_26302,N_26390);
and U28013 (N_28013,N_25774,N_26866);
nand U28014 (N_28014,N_26518,N_25913);
nand U28015 (N_28015,N_25638,N_26221);
xor U28016 (N_28016,N_25724,N_26845);
and U28017 (N_28017,N_26561,N_26708);
nand U28018 (N_28018,N_26804,N_26323);
nor U28019 (N_28019,N_26298,N_26584);
and U28020 (N_28020,N_26884,N_26535);
nor U28021 (N_28021,N_26089,N_26006);
nand U28022 (N_28022,N_26348,N_25627);
nand U28023 (N_28023,N_26142,N_25930);
or U28024 (N_28024,N_26442,N_26524);
nand U28025 (N_28025,N_25595,N_25599);
nor U28026 (N_28026,N_25709,N_26183);
and U28027 (N_28027,N_25781,N_26224);
nor U28028 (N_28028,N_26415,N_26327);
nor U28029 (N_28029,N_26744,N_26516);
and U28030 (N_28030,N_26703,N_26695);
xnor U28031 (N_28031,N_26811,N_25917);
nand U28032 (N_28032,N_26366,N_26261);
or U28033 (N_28033,N_25889,N_26435);
nand U28034 (N_28034,N_26010,N_26773);
xor U28035 (N_28035,N_25876,N_26280);
and U28036 (N_28036,N_26715,N_26922);
nand U28037 (N_28037,N_25530,N_25701);
nor U28038 (N_28038,N_26592,N_25519);
xnor U28039 (N_28039,N_25504,N_25735);
and U28040 (N_28040,N_26463,N_26586);
nor U28041 (N_28041,N_25629,N_26740);
nand U28042 (N_28042,N_26092,N_26962);
nor U28043 (N_28043,N_26530,N_26367);
nor U28044 (N_28044,N_26659,N_26373);
nor U28045 (N_28045,N_25945,N_25740);
nand U28046 (N_28046,N_25715,N_26799);
nor U28047 (N_28047,N_25733,N_25573);
nor U28048 (N_28048,N_26720,N_26427);
nor U28049 (N_28049,N_25529,N_26830);
nand U28050 (N_28050,N_26336,N_26631);
nor U28051 (N_28051,N_26963,N_25732);
or U28052 (N_28052,N_26345,N_25883);
xor U28053 (N_28053,N_25731,N_26315);
xnor U28054 (N_28054,N_26221,N_26826);
nand U28055 (N_28055,N_26412,N_26434);
nand U28056 (N_28056,N_26044,N_25879);
nor U28057 (N_28057,N_26237,N_26751);
nand U28058 (N_28058,N_26068,N_26908);
nand U28059 (N_28059,N_26713,N_25978);
nor U28060 (N_28060,N_25844,N_26614);
and U28061 (N_28061,N_26062,N_25779);
nand U28062 (N_28062,N_25710,N_26276);
nand U28063 (N_28063,N_26593,N_25500);
nor U28064 (N_28064,N_26312,N_26874);
xor U28065 (N_28065,N_26135,N_25770);
and U28066 (N_28066,N_25908,N_26554);
and U28067 (N_28067,N_26316,N_26040);
nor U28068 (N_28068,N_26986,N_25631);
nor U28069 (N_28069,N_25933,N_26798);
nor U28070 (N_28070,N_26016,N_26722);
nand U28071 (N_28071,N_26938,N_26312);
nand U28072 (N_28072,N_26216,N_26011);
xor U28073 (N_28073,N_26953,N_26334);
xor U28074 (N_28074,N_25992,N_26919);
xnor U28075 (N_28075,N_26813,N_25851);
or U28076 (N_28076,N_25929,N_25605);
nor U28077 (N_28077,N_26898,N_26660);
xnor U28078 (N_28078,N_26759,N_26758);
or U28079 (N_28079,N_25946,N_26496);
or U28080 (N_28080,N_25869,N_26829);
nor U28081 (N_28081,N_25719,N_26539);
and U28082 (N_28082,N_25976,N_26508);
and U28083 (N_28083,N_25822,N_26858);
nand U28084 (N_28084,N_26649,N_25831);
and U28085 (N_28085,N_26229,N_26151);
and U28086 (N_28086,N_26486,N_26838);
nand U28087 (N_28087,N_26706,N_26286);
nand U28088 (N_28088,N_26325,N_26644);
nand U28089 (N_28089,N_26869,N_26881);
nand U28090 (N_28090,N_26490,N_25815);
xnor U28091 (N_28091,N_26524,N_26610);
and U28092 (N_28092,N_25877,N_25734);
nand U28093 (N_28093,N_25714,N_26875);
xnor U28094 (N_28094,N_26862,N_26783);
xor U28095 (N_28095,N_25840,N_26875);
nor U28096 (N_28096,N_26026,N_26175);
nand U28097 (N_28097,N_25991,N_26291);
xnor U28098 (N_28098,N_25849,N_26955);
xor U28099 (N_28099,N_25501,N_25823);
and U28100 (N_28100,N_25535,N_25533);
or U28101 (N_28101,N_25537,N_26006);
and U28102 (N_28102,N_25819,N_26086);
nor U28103 (N_28103,N_26122,N_26443);
nand U28104 (N_28104,N_26186,N_26083);
nand U28105 (N_28105,N_26980,N_25547);
nand U28106 (N_28106,N_26503,N_26418);
and U28107 (N_28107,N_26962,N_26451);
nand U28108 (N_28108,N_25694,N_25976);
or U28109 (N_28109,N_26815,N_26063);
or U28110 (N_28110,N_26219,N_26751);
nand U28111 (N_28111,N_25977,N_25898);
nand U28112 (N_28112,N_26748,N_26576);
and U28113 (N_28113,N_26140,N_26875);
or U28114 (N_28114,N_26204,N_26034);
or U28115 (N_28115,N_25970,N_25531);
or U28116 (N_28116,N_26206,N_25923);
xor U28117 (N_28117,N_26469,N_26141);
nor U28118 (N_28118,N_26308,N_26006);
nor U28119 (N_28119,N_26635,N_26230);
and U28120 (N_28120,N_26138,N_26120);
nand U28121 (N_28121,N_25606,N_26816);
nand U28122 (N_28122,N_26034,N_26661);
xor U28123 (N_28123,N_26442,N_26363);
nand U28124 (N_28124,N_26893,N_25720);
nor U28125 (N_28125,N_26981,N_25730);
xnor U28126 (N_28126,N_26523,N_26355);
nand U28127 (N_28127,N_25550,N_25872);
nand U28128 (N_28128,N_26612,N_26695);
and U28129 (N_28129,N_25640,N_26080);
or U28130 (N_28130,N_26093,N_25761);
nand U28131 (N_28131,N_26956,N_25613);
or U28132 (N_28132,N_26453,N_25597);
or U28133 (N_28133,N_25842,N_25554);
nor U28134 (N_28134,N_25991,N_25747);
xnor U28135 (N_28135,N_26365,N_25723);
or U28136 (N_28136,N_25785,N_25538);
nand U28137 (N_28137,N_25598,N_26457);
nand U28138 (N_28138,N_26212,N_25580);
xnor U28139 (N_28139,N_25923,N_26438);
nand U28140 (N_28140,N_26260,N_26213);
nand U28141 (N_28141,N_26859,N_26604);
nor U28142 (N_28142,N_26993,N_26617);
nand U28143 (N_28143,N_26099,N_26576);
xor U28144 (N_28144,N_26850,N_25827);
and U28145 (N_28145,N_26838,N_25784);
xnor U28146 (N_28146,N_26847,N_25681);
nand U28147 (N_28147,N_26426,N_26327);
nand U28148 (N_28148,N_26876,N_26654);
nand U28149 (N_28149,N_26248,N_25889);
nor U28150 (N_28150,N_26614,N_26555);
nand U28151 (N_28151,N_26258,N_26116);
nand U28152 (N_28152,N_26916,N_26190);
nor U28153 (N_28153,N_25620,N_25838);
nor U28154 (N_28154,N_25687,N_25683);
and U28155 (N_28155,N_26070,N_25653);
nand U28156 (N_28156,N_25784,N_26038);
nor U28157 (N_28157,N_26602,N_26515);
xnor U28158 (N_28158,N_26180,N_26298);
or U28159 (N_28159,N_26645,N_25664);
nor U28160 (N_28160,N_26060,N_25991);
nand U28161 (N_28161,N_26722,N_26405);
nand U28162 (N_28162,N_26861,N_26599);
nor U28163 (N_28163,N_26371,N_25561);
nand U28164 (N_28164,N_25804,N_26438);
or U28165 (N_28165,N_26640,N_25738);
nand U28166 (N_28166,N_25977,N_26784);
xor U28167 (N_28167,N_26466,N_26069);
nand U28168 (N_28168,N_26658,N_25721);
nor U28169 (N_28169,N_26956,N_25655);
xor U28170 (N_28170,N_25736,N_26659);
or U28171 (N_28171,N_25878,N_26553);
xnor U28172 (N_28172,N_26565,N_26654);
nor U28173 (N_28173,N_26962,N_25619);
nor U28174 (N_28174,N_26022,N_25698);
and U28175 (N_28175,N_26439,N_26666);
or U28176 (N_28176,N_26364,N_25613);
and U28177 (N_28177,N_26466,N_26192);
nor U28178 (N_28178,N_25775,N_25823);
or U28179 (N_28179,N_26687,N_26483);
xor U28180 (N_28180,N_26338,N_25628);
nand U28181 (N_28181,N_25876,N_26323);
nand U28182 (N_28182,N_25515,N_26561);
or U28183 (N_28183,N_25530,N_26304);
xnor U28184 (N_28184,N_26953,N_26106);
xnor U28185 (N_28185,N_25815,N_26118);
xnor U28186 (N_28186,N_26932,N_26549);
nor U28187 (N_28187,N_26366,N_26270);
nor U28188 (N_28188,N_26750,N_25545);
xor U28189 (N_28189,N_26870,N_26196);
nor U28190 (N_28190,N_26820,N_25830);
and U28191 (N_28191,N_26344,N_26072);
xor U28192 (N_28192,N_26140,N_26337);
nand U28193 (N_28193,N_25703,N_25862);
and U28194 (N_28194,N_25723,N_26503);
xor U28195 (N_28195,N_26867,N_26001);
or U28196 (N_28196,N_26819,N_25751);
nand U28197 (N_28197,N_26680,N_25706);
and U28198 (N_28198,N_26506,N_25790);
xor U28199 (N_28199,N_26796,N_26235);
and U28200 (N_28200,N_26758,N_26927);
nor U28201 (N_28201,N_25857,N_26676);
and U28202 (N_28202,N_25583,N_26734);
nand U28203 (N_28203,N_25819,N_26339);
and U28204 (N_28204,N_26300,N_25878);
or U28205 (N_28205,N_26138,N_25752);
or U28206 (N_28206,N_26392,N_26488);
or U28207 (N_28207,N_26350,N_25994);
and U28208 (N_28208,N_25805,N_26391);
nand U28209 (N_28209,N_26202,N_26056);
or U28210 (N_28210,N_26610,N_26473);
nor U28211 (N_28211,N_25818,N_26381);
xor U28212 (N_28212,N_25938,N_25704);
or U28213 (N_28213,N_26257,N_25988);
nand U28214 (N_28214,N_26589,N_25958);
nor U28215 (N_28215,N_26967,N_25911);
or U28216 (N_28216,N_26014,N_25997);
and U28217 (N_28217,N_26959,N_25772);
and U28218 (N_28218,N_26892,N_26122);
nor U28219 (N_28219,N_25879,N_26747);
nand U28220 (N_28220,N_25569,N_26510);
nand U28221 (N_28221,N_26504,N_25737);
nand U28222 (N_28222,N_25942,N_26225);
or U28223 (N_28223,N_26852,N_26049);
nand U28224 (N_28224,N_26411,N_25857);
nand U28225 (N_28225,N_26448,N_26431);
nand U28226 (N_28226,N_26839,N_25833);
xor U28227 (N_28227,N_25716,N_25920);
xor U28228 (N_28228,N_26879,N_26126);
and U28229 (N_28229,N_25672,N_26879);
nand U28230 (N_28230,N_26155,N_25503);
and U28231 (N_28231,N_26332,N_26717);
xor U28232 (N_28232,N_26516,N_26372);
xnor U28233 (N_28233,N_26829,N_26744);
or U28234 (N_28234,N_26157,N_25603);
and U28235 (N_28235,N_26881,N_26658);
nand U28236 (N_28236,N_26560,N_25792);
or U28237 (N_28237,N_26886,N_25571);
xnor U28238 (N_28238,N_26277,N_25849);
nor U28239 (N_28239,N_25676,N_26127);
or U28240 (N_28240,N_26254,N_25845);
nand U28241 (N_28241,N_25962,N_26334);
or U28242 (N_28242,N_26539,N_26867);
nand U28243 (N_28243,N_25676,N_26165);
nor U28244 (N_28244,N_25584,N_26078);
nor U28245 (N_28245,N_26065,N_25655);
or U28246 (N_28246,N_25880,N_25952);
nor U28247 (N_28247,N_26144,N_26693);
nand U28248 (N_28248,N_26197,N_25803);
nor U28249 (N_28249,N_25875,N_26874);
nor U28250 (N_28250,N_25657,N_26233);
xor U28251 (N_28251,N_26853,N_26542);
or U28252 (N_28252,N_26451,N_26227);
nand U28253 (N_28253,N_25686,N_25525);
and U28254 (N_28254,N_26138,N_26801);
nor U28255 (N_28255,N_26014,N_26745);
and U28256 (N_28256,N_26850,N_26121);
and U28257 (N_28257,N_26103,N_26337);
nor U28258 (N_28258,N_26137,N_26276);
or U28259 (N_28259,N_26247,N_26599);
and U28260 (N_28260,N_26803,N_26806);
and U28261 (N_28261,N_26268,N_25915);
and U28262 (N_28262,N_26724,N_26420);
and U28263 (N_28263,N_26932,N_26341);
and U28264 (N_28264,N_25937,N_26734);
or U28265 (N_28265,N_26205,N_26353);
or U28266 (N_28266,N_26380,N_26253);
or U28267 (N_28267,N_26593,N_25835);
or U28268 (N_28268,N_26751,N_25951);
nor U28269 (N_28269,N_26423,N_26260);
or U28270 (N_28270,N_26589,N_26403);
nand U28271 (N_28271,N_26637,N_26489);
xnor U28272 (N_28272,N_25698,N_26097);
nor U28273 (N_28273,N_25913,N_26628);
nand U28274 (N_28274,N_25992,N_26165);
and U28275 (N_28275,N_26585,N_26594);
xor U28276 (N_28276,N_25819,N_25793);
or U28277 (N_28277,N_26074,N_25911);
and U28278 (N_28278,N_25757,N_26788);
nor U28279 (N_28279,N_26794,N_26471);
or U28280 (N_28280,N_26542,N_25662);
or U28281 (N_28281,N_25623,N_25831);
nand U28282 (N_28282,N_25897,N_26541);
and U28283 (N_28283,N_26290,N_25868);
xnor U28284 (N_28284,N_25743,N_26632);
and U28285 (N_28285,N_26524,N_26219);
xnor U28286 (N_28286,N_26778,N_26719);
or U28287 (N_28287,N_25618,N_26292);
nand U28288 (N_28288,N_26621,N_26741);
or U28289 (N_28289,N_26267,N_26661);
nor U28290 (N_28290,N_26573,N_25809);
and U28291 (N_28291,N_26925,N_26808);
xor U28292 (N_28292,N_25551,N_26975);
nor U28293 (N_28293,N_26172,N_26257);
or U28294 (N_28294,N_26943,N_25562);
nand U28295 (N_28295,N_26734,N_25943);
and U28296 (N_28296,N_26344,N_26144);
nor U28297 (N_28297,N_26844,N_25852);
or U28298 (N_28298,N_25525,N_25664);
or U28299 (N_28299,N_26076,N_26639);
nor U28300 (N_28300,N_26190,N_25692);
and U28301 (N_28301,N_26591,N_26353);
or U28302 (N_28302,N_25576,N_25825);
xnor U28303 (N_28303,N_26542,N_26236);
nor U28304 (N_28304,N_25926,N_26634);
nor U28305 (N_28305,N_26749,N_26001);
nor U28306 (N_28306,N_26512,N_26218);
nor U28307 (N_28307,N_26110,N_26529);
or U28308 (N_28308,N_26828,N_26019);
or U28309 (N_28309,N_25642,N_26214);
nand U28310 (N_28310,N_26179,N_26564);
xnor U28311 (N_28311,N_26512,N_26179);
nand U28312 (N_28312,N_26314,N_26691);
or U28313 (N_28313,N_26398,N_25772);
or U28314 (N_28314,N_26657,N_25880);
xor U28315 (N_28315,N_26593,N_26261);
and U28316 (N_28316,N_26026,N_26782);
nor U28317 (N_28317,N_25594,N_26902);
nand U28318 (N_28318,N_26952,N_25530);
nand U28319 (N_28319,N_26170,N_25598);
nor U28320 (N_28320,N_26428,N_25670);
nand U28321 (N_28321,N_25582,N_26904);
nand U28322 (N_28322,N_26150,N_26810);
nand U28323 (N_28323,N_25690,N_26910);
or U28324 (N_28324,N_26224,N_25815);
and U28325 (N_28325,N_26837,N_26529);
or U28326 (N_28326,N_26237,N_25667);
and U28327 (N_28327,N_26037,N_25957);
xor U28328 (N_28328,N_26253,N_26968);
and U28329 (N_28329,N_25698,N_25838);
nand U28330 (N_28330,N_26603,N_26619);
nor U28331 (N_28331,N_26330,N_26366);
and U28332 (N_28332,N_26467,N_25913);
and U28333 (N_28333,N_26706,N_26925);
xnor U28334 (N_28334,N_26346,N_25978);
and U28335 (N_28335,N_26507,N_25839);
nor U28336 (N_28336,N_25711,N_26009);
and U28337 (N_28337,N_26336,N_25516);
or U28338 (N_28338,N_26995,N_26295);
and U28339 (N_28339,N_25983,N_25999);
or U28340 (N_28340,N_25978,N_26639);
nand U28341 (N_28341,N_26281,N_26170);
and U28342 (N_28342,N_26220,N_26080);
xnor U28343 (N_28343,N_26191,N_25640);
nand U28344 (N_28344,N_25993,N_25513);
or U28345 (N_28345,N_26842,N_25714);
xnor U28346 (N_28346,N_25725,N_26423);
or U28347 (N_28347,N_25906,N_26596);
nand U28348 (N_28348,N_26609,N_26369);
xnor U28349 (N_28349,N_25837,N_25506);
xnor U28350 (N_28350,N_25666,N_25890);
nand U28351 (N_28351,N_26994,N_26163);
and U28352 (N_28352,N_26189,N_26172);
or U28353 (N_28353,N_25782,N_25589);
or U28354 (N_28354,N_26692,N_25947);
and U28355 (N_28355,N_26779,N_26035);
nand U28356 (N_28356,N_26199,N_25804);
nand U28357 (N_28357,N_26634,N_26275);
nor U28358 (N_28358,N_26600,N_25904);
nand U28359 (N_28359,N_26325,N_26982);
xnor U28360 (N_28360,N_25579,N_26128);
nand U28361 (N_28361,N_25654,N_26463);
nand U28362 (N_28362,N_25990,N_25615);
nand U28363 (N_28363,N_26346,N_25539);
and U28364 (N_28364,N_26868,N_25624);
nand U28365 (N_28365,N_25659,N_26098);
nor U28366 (N_28366,N_26517,N_26963);
nor U28367 (N_28367,N_25994,N_26706);
or U28368 (N_28368,N_26148,N_26539);
nand U28369 (N_28369,N_26591,N_25771);
nand U28370 (N_28370,N_25729,N_25738);
nor U28371 (N_28371,N_26303,N_26913);
or U28372 (N_28372,N_25718,N_25560);
or U28373 (N_28373,N_25835,N_25530);
nor U28374 (N_28374,N_25866,N_25586);
nand U28375 (N_28375,N_26969,N_25861);
nor U28376 (N_28376,N_26177,N_26224);
or U28377 (N_28377,N_26083,N_25778);
nor U28378 (N_28378,N_26197,N_26155);
nand U28379 (N_28379,N_25574,N_26999);
nand U28380 (N_28380,N_26492,N_25828);
and U28381 (N_28381,N_26809,N_25693);
nand U28382 (N_28382,N_25782,N_25521);
nor U28383 (N_28383,N_26004,N_26954);
and U28384 (N_28384,N_26242,N_25631);
and U28385 (N_28385,N_26936,N_26015);
xor U28386 (N_28386,N_25504,N_26283);
nand U28387 (N_28387,N_25956,N_26591);
nand U28388 (N_28388,N_26265,N_26322);
and U28389 (N_28389,N_26099,N_26489);
xnor U28390 (N_28390,N_25963,N_26478);
and U28391 (N_28391,N_26388,N_26998);
and U28392 (N_28392,N_26088,N_25842);
xor U28393 (N_28393,N_26636,N_26022);
nand U28394 (N_28394,N_26098,N_25557);
or U28395 (N_28395,N_26456,N_26467);
xor U28396 (N_28396,N_26588,N_26410);
nand U28397 (N_28397,N_25802,N_25869);
or U28398 (N_28398,N_25746,N_26106);
or U28399 (N_28399,N_26792,N_26884);
xor U28400 (N_28400,N_26297,N_25681);
nand U28401 (N_28401,N_25956,N_26706);
and U28402 (N_28402,N_26570,N_26499);
xnor U28403 (N_28403,N_25980,N_25919);
or U28404 (N_28404,N_26359,N_26006);
or U28405 (N_28405,N_26247,N_26140);
xnor U28406 (N_28406,N_25676,N_25922);
xor U28407 (N_28407,N_26553,N_26084);
xnor U28408 (N_28408,N_26809,N_26845);
xnor U28409 (N_28409,N_26334,N_26244);
nor U28410 (N_28410,N_25792,N_26017);
and U28411 (N_28411,N_25933,N_25581);
nand U28412 (N_28412,N_26279,N_26671);
xnor U28413 (N_28413,N_26219,N_26424);
nor U28414 (N_28414,N_25914,N_26819);
nor U28415 (N_28415,N_26057,N_25999);
and U28416 (N_28416,N_26753,N_26371);
xor U28417 (N_28417,N_26614,N_26236);
nand U28418 (N_28418,N_26523,N_25735);
and U28419 (N_28419,N_26718,N_25640);
nor U28420 (N_28420,N_25604,N_25690);
and U28421 (N_28421,N_26609,N_26582);
xnor U28422 (N_28422,N_26447,N_25725);
nor U28423 (N_28423,N_26433,N_25577);
or U28424 (N_28424,N_26019,N_25683);
and U28425 (N_28425,N_26900,N_25873);
xnor U28426 (N_28426,N_25973,N_26101);
nor U28427 (N_28427,N_25870,N_26884);
xor U28428 (N_28428,N_26134,N_26391);
xor U28429 (N_28429,N_26725,N_26042);
nor U28430 (N_28430,N_26000,N_26605);
and U28431 (N_28431,N_26804,N_26099);
xnor U28432 (N_28432,N_26298,N_26712);
and U28433 (N_28433,N_26663,N_25877);
nor U28434 (N_28434,N_26195,N_26946);
nand U28435 (N_28435,N_26034,N_26686);
and U28436 (N_28436,N_26744,N_26625);
nand U28437 (N_28437,N_25900,N_26869);
xor U28438 (N_28438,N_26467,N_25765);
xnor U28439 (N_28439,N_26781,N_26632);
nand U28440 (N_28440,N_26181,N_26397);
and U28441 (N_28441,N_26969,N_25971);
or U28442 (N_28442,N_26310,N_26811);
and U28443 (N_28443,N_26009,N_26832);
or U28444 (N_28444,N_25948,N_25551);
xnor U28445 (N_28445,N_26112,N_26385);
and U28446 (N_28446,N_26867,N_25895);
nand U28447 (N_28447,N_25522,N_26841);
nor U28448 (N_28448,N_26174,N_25929);
or U28449 (N_28449,N_25598,N_25893);
xnor U28450 (N_28450,N_26782,N_26640);
and U28451 (N_28451,N_26865,N_25805);
xor U28452 (N_28452,N_25984,N_26203);
xnor U28453 (N_28453,N_26949,N_26384);
nor U28454 (N_28454,N_26687,N_26317);
or U28455 (N_28455,N_25627,N_26525);
nor U28456 (N_28456,N_25812,N_26319);
xor U28457 (N_28457,N_26063,N_25820);
and U28458 (N_28458,N_26726,N_26903);
xor U28459 (N_28459,N_26905,N_26620);
xor U28460 (N_28460,N_25866,N_25609);
or U28461 (N_28461,N_26540,N_25567);
nor U28462 (N_28462,N_26958,N_25720);
or U28463 (N_28463,N_26016,N_26910);
or U28464 (N_28464,N_26200,N_26196);
and U28465 (N_28465,N_26581,N_25923);
nand U28466 (N_28466,N_26857,N_25628);
or U28467 (N_28467,N_26855,N_25596);
xor U28468 (N_28468,N_26262,N_25985);
and U28469 (N_28469,N_25557,N_25753);
and U28470 (N_28470,N_25740,N_25803);
and U28471 (N_28471,N_25536,N_26149);
and U28472 (N_28472,N_26504,N_26047);
or U28473 (N_28473,N_26416,N_25510);
xor U28474 (N_28474,N_26250,N_25722);
or U28475 (N_28475,N_25759,N_25532);
or U28476 (N_28476,N_26470,N_26890);
and U28477 (N_28477,N_26113,N_25874);
and U28478 (N_28478,N_26888,N_26046);
and U28479 (N_28479,N_26814,N_25698);
xnor U28480 (N_28480,N_25503,N_26536);
or U28481 (N_28481,N_25777,N_25954);
nand U28482 (N_28482,N_26716,N_25919);
or U28483 (N_28483,N_25876,N_26322);
nor U28484 (N_28484,N_25620,N_26682);
and U28485 (N_28485,N_26253,N_25516);
and U28486 (N_28486,N_25582,N_25938);
xnor U28487 (N_28487,N_26898,N_26582);
nand U28488 (N_28488,N_26579,N_26858);
nor U28489 (N_28489,N_26209,N_25641);
nand U28490 (N_28490,N_26494,N_26458);
or U28491 (N_28491,N_26363,N_25662);
or U28492 (N_28492,N_26568,N_25755);
or U28493 (N_28493,N_26049,N_25826);
and U28494 (N_28494,N_26478,N_26403);
nor U28495 (N_28495,N_25614,N_26813);
nand U28496 (N_28496,N_26201,N_26561);
nor U28497 (N_28497,N_25952,N_26326);
and U28498 (N_28498,N_26359,N_26535);
and U28499 (N_28499,N_26608,N_26533);
nand U28500 (N_28500,N_27774,N_27832);
and U28501 (N_28501,N_27050,N_27688);
or U28502 (N_28502,N_27247,N_27376);
nor U28503 (N_28503,N_28257,N_27638);
xor U28504 (N_28504,N_27130,N_28438);
and U28505 (N_28505,N_28376,N_27422);
xor U28506 (N_28506,N_27118,N_28450);
or U28507 (N_28507,N_27812,N_27049);
nand U28508 (N_28508,N_27484,N_27886);
nor U28509 (N_28509,N_27252,N_27485);
xnor U28510 (N_28510,N_28305,N_28269);
and U28511 (N_28511,N_27302,N_27365);
or U28512 (N_28512,N_27428,N_27319);
xnor U28513 (N_28513,N_28379,N_27132);
or U28514 (N_28514,N_27855,N_27299);
nand U28515 (N_28515,N_27462,N_28444);
and U28516 (N_28516,N_27227,N_27902);
xnor U28517 (N_28517,N_27841,N_27408);
nand U28518 (N_28518,N_27268,N_28171);
xnor U28519 (N_28519,N_28299,N_27248);
nand U28520 (N_28520,N_28074,N_27294);
nand U28521 (N_28521,N_27303,N_27188);
or U28522 (N_28522,N_28119,N_28015);
and U28523 (N_28523,N_27581,N_27766);
nor U28524 (N_28524,N_27906,N_27684);
and U28525 (N_28525,N_27004,N_27487);
nor U28526 (N_28526,N_27585,N_27880);
nor U28527 (N_28527,N_27963,N_28273);
xor U28528 (N_28528,N_27259,N_27583);
nor U28529 (N_28529,N_27021,N_27289);
nor U28530 (N_28530,N_28236,N_27596);
xor U28531 (N_28531,N_28222,N_27957);
or U28532 (N_28532,N_27134,N_28064);
and U28533 (N_28533,N_27033,N_27123);
nand U28534 (N_28534,N_28398,N_27994);
nor U28535 (N_28535,N_28090,N_27269);
nand U28536 (N_28536,N_27213,N_28146);
and U28537 (N_28537,N_27680,N_27710);
and U28538 (N_28538,N_27988,N_27477);
or U28539 (N_28539,N_27073,N_28293);
xnor U28540 (N_28540,N_28012,N_27787);
and U28541 (N_28541,N_28336,N_27324);
or U28542 (N_28542,N_27052,N_27557);
or U28543 (N_28543,N_27386,N_27790);
and U28544 (N_28544,N_27367,N_27037);
or U28545 (N_28545,N_28075,N_27821);
or U28546 (N_28546,N_28041,N_27579);
xor U28547 (N_28547,N_27076,N_27899);
and U28548 (N_28548,N_28499,N_27340);
and U28549 (N_28549,N_27005,N_27475);
xnor U28550 (N_28550,N_27537,N_27858);
or U28551 (N_28551,N_28202,N_28322);
xnor U28552 (N_28552,N_27186,N_27452);
nor U28553 (N_28553,N_27115,N_27629);
nand U28554 (N_28554,N_27893,N_27610);
and U28555 (N_28555,N_28161,N_27410);
or U28556 (N_28556,N_27960,N_28410);
nor U28557 (N_28557,N_27089,N_27000);
and U28558 (N_28558,N_27335,N_27962);
nor U28559 (N_28559,N_27580,N_27479);
or U28560 (N_28560,N_27257,N_27167);
and U28561 (N_28561,N_28114,N_27469);
xnor U28562 (N_28562,N_27313,N_28429);
nor U28563 (N_28563,N_27421,N_27308);
or U28564 (N_28564,N_27124,N_28439);
nor U28565 (N_28565,N_27322,N_27430);
and U28566 (N_28566,N_28489,N_28203);
and U28567 (N_28567,N_27008,N_27200);
nand U28568 (N_28568,N_27657,N_27728);
nand U28569 (N_28569,N_27862,N_27330);
xor U28570 (N_28570,N_27418,N_28488);
xor U28571 (N_28571,N_27178,N_27206);
xor U28572 (N_28572,N_27652,N_27411);
nor U28573 (N_28573,N_27511,N_28413);
nor U28574 (N_28574,N_28158,N_28253);
nor U28575 (N_28575,N_28474,N_28352);
xnor U28576 (N_28576,N_27744,N_27375);
nand U28577 (N_28577,N_27575,N_27195);
nor U28578 (N_28578,N_27378,N_28251);
xnor U28579 (N_28579,N_28003,N_28033);
xnor U28580 (N_28580,N_27498,N_27509);
nor U28581 (N_28581,N_28343,N_27329);
or U28582 (N_28582,N_28229,N_27772);
nand U28583 (N_28583,N_27990,N_27518);
or U28584 (N_28584,N_27292,N_27887);
nor U28585 (N_28585,N_27937,N_27516);
or U28586 (N_28586,N_27474,N_27729);
or U28587 (N_28587,N_28362,N_27871);
nor U28588 (N_28588,N_27122,N_27587);
nor U28589 (N_28589,N_27136,N_27077);
nand U28590 (N_28590,N_27951,N_27342);
nor U28591 (N_28591,N_27320,N_27120);
xor U28592 (N_28592,N_27226,N_27718);
nand U28593 (N_28593,N_28148,N_27189);
and U28594 (N_28594,N_28492,N_27746);
nand U28595 (N_28595,N_27819,N_27187);
nand U28596 (N_28596,N_28479,N_28463);
xor U28597 (N_28597,N_27471,N_28260);
nand U28598 (N_28598,N_27641,N_27529);
and U28599 (N_28599,N_27085,N_27045);
or U28600 (N_28600,N_27336,N_28081);
and U28601 (N_28601,N_27524,N_28340);
and U28602 (N_28602,N_27467,N_27443);
xor U28603 (N_28603,N_27755,N_27797);
and U28604 (N_28604,N_27568,N_28195);
nand U28605 (N_28605,N_28028,N_28278);
nor U28606 (N_28606,N_27080,N_27267);
xor U28607 (N_28607,N_27013,N_28310);
and U28608 (N_28608,N_28226,N_27611);
or U28609 (N_28609,N_27846,N_27553);
xor U28610 (N_28610,N_27423,N_27700);
nor U28611 (N_28611,N_28483,N_27091);
nand U28612 (N_28612,N_27141,N_28136);
nor U28613 (N_28613,N_27799,N_28454);
nand U28614 (N_28614,N_27170,N_28065);
or U28615 (N_28615,N_28349,N_27977);
nor U28616 (N_28616,N_27952,N_27672);
nor U28617 (N_28617,N_28001,N_28459);
nor U28618 (N_28618,N_27041,N_28211);
nand U28619 (N_28619,N_28159,N_27043);
or U28620 (N_28620,N_27626,N_28453);
nor U28621 (N_28621,N_28373,N_27505);
or U28622 (N_28622,N_27722,N_28032);
and U28623 (N_28623,N_28476,N_28217);
or U28624 (N_28624,N_27415,N_27876);
nand U28625 (N_28625,N_27143,N_27119);
xor U28626 (N_28626,N_28268,N_28049);
and U28627 (N_28627,N_27555,N_27765);
nor U28628 (N_28628,N_27621,N_27732);
nand U28629 (N_28629,N_28281,N_27642);
xnor U28630 (N_28630,N_28381,N_27613);
or U28631 (N_28631,N_28311,N_27792);
nor U28632 (N_28632,N_27543,N_27196);
and U28633 (N_28633,N_27798,N_27762);
xnor U28634 (N_28634,N_27117,N_28177);
xor U28635 (N_28635,N_28408,N_28233);
or U28636 (N_28636,N_27215,N_27780);
and U28637 (N_28637,N_27333,N_28404);
xor U28638 (N_28638,N_27157,N_27889);
nand U28639 (N_28639,N_28180,N_27873);
xnor U28640 (N_28640,N_27346,N_28153);
xor U28641 (N_28641,N_27959,N_27087);
or U28642 (N_28642,N_27857,N_27923);
xor U28643 (N_28643,N_27293,N_28187);
nand U28644 (N_28644,N_27872,N_28369);
and U28645 (N_28645,N_27493,N_27218);
or U28646 (N_28646,N_27689,N_27653);
nand U28647 (N_28647,N_28042,N_28484);
or U28648 (N_28648,N_27417,N_28017);
xor U28649 (N_28649,N_28416,N_28143);
xnor U28650 (N_28650,N_28319,N_27190);
and U28651 (N_28651,N_27995,N_27769);
nand U28652 (N_28652,N_27369,N_27907);
and U28653 (N_28653,N_27687,N_28462);
nor U28654 (N_28654,N_27788,N_28421);
and U28655 (N_28655,N_28289,N_27864);
nand U28656 (N_28656,N_27881,N_28024);
nor U28657 (N_28657,N_28068,N_27607);
nor U28658 (N_28658,N_27823,N_28250);
xnor U28659 (N_28659,N_27817,N_28447);
xor U28660 (N_28660,N_28393,N_27752);
or U28661 (N_28661,N_27933,N_27738);
nand U28662 (N_28662,N_28098,N_28051);
nand U28663 (N_28663,N_28286,N_28204);
xor U28664 (N_28664,N_27010,N_27260);
nand U28665 (N_28665,N_28035,N_28231);
nand U28666 (N_28666,N_27090,N_27332);
and U28667 (N_28667,N_28004,N_28296);
xnor U28668 (N_28668,N_28436,N_27448);
or U28669 (N_28669,N_28384,N_27096);
nand U28670 (N_28670,N_28411,N_27290);
and U28671 (N_28671,N_27343,N_28209);
and U28672 (N_28672,N_27840,N_27446);
nand U28673 (N_28673,N_27399,N_27701);
nor U28674 (N_28674,N_27915,N_28168);
nand U28675 (N_28675,N_27197,N_27104);
xnor U28676 (N_28676,N_27686,N_27595);
xnor U28677 (N_28677,N_27121,N_28294);
xor U28678 (N_28678,N_28259,N_27549);
xnor U28679 (N_28679,N_27300,N_27255);
and U28680 (N_28680,N_27985,N_27162);
and U28681 (N_28681,N_27225,N_27605);
nand U28682 (N_28682,N_28131,N_27497);
xnor U28683 (N_28683,N_27402,N_28247);
nand U28684 (N_28684,N_28058,N_27295);
and U28685 (N_28685,N_27879,N_27747);
nor U28686 (N_28686,N_27639,N_28298);
nand U28687 (N_28687,N_28256,N_27285);
or U28688 (N_28688,N_27166,N_28297);
or U28689 (N_28689,N_28277,N_28280);
and U28690 (N_28690,N_27814,N_28060);
nand U28691 (N_28691,N_27109,N_28368);
and U28692 (N_28692,N_28077,N_27412);
and U28693 (N_28693,N_28040,N_27387);
and U28694 (N_28694,N_27699,N_28225);
nand U28695 (N_28695,N_27550,N_27997);
xor U28696 (N_28696,N_27753,N_27724);
nor U28697 (N_28697,N_27586,N_27665);
nand U28698 (N_28698,N_27608,N_27420);
xor U28699 (N_28699,N_27949,N_28082);
xor U28700 (N_28700,N_28435,N_27370);
nor U28701 (N_28701,N_28219,N_28216);
and U28702 (N_28702,N_27251,N_28312);
nor U28703 (N_28703,N_27107,N_27964);
nor U28704 (N_28704,N_28071,N_27459);
nor U28705 (N_28705,N_28262,N_27110);
or U28706 (N_28706,N_27069,N_28053);
nand U28707 (N_28707,N_27203,N_27897);
xor U28708 (N_28708,N_27311,N_27092);
xnor U28709 (N_28709,N_27507,N_27741);
and U28710 (N_28710,N_28224,N_27204);
or U28711 (N_28711,N_27305,N_27736);
xnor U28712 (N_28712,N_28045,N_27882);
or U28713 (N_28713,N_27079,N_27145);
or U28714 (N_28714,N_27253,N_27974);
and U28715 (N_28715,N_28440,N_27455);
and U28716 (N_28716,N_27827,N_27914);
and U28717 (N_28717,N_28050,N_27159);
and U28718 (N_28718,N_28457,N_27433);
and U28719 (N_28719,N_27640,N_27270);
xnor U28720 (N_28720,N_27835,N_28481);
and U28721 (N_28721,N_27192,N_28495);
and U28722 (N_28722,N_27184,N_28498);
xnor U28723 (N_28723,N_28324,N_27643);
and U28724 (N_28724,N_28473,N_27989);
nand U28725 (N_28725,N_27707,N_28170);
nor U28726 (N_28726,N_27379,N_27174);
xor U28727 (N_28727,N_27044,N_27712);
xor U28728 (N_28728,N_27784,N_27669);
nand U28729 (N_28729,N_27150,N_28383);
xor U28730 (N_28730,N_28016,N_28487);
xor U28731 (N_28731,N_28140,N_27185);
nor U28732 (N_28732,N_27648,N_28283);
and U28733 (N_28733,N_27725,N_27490);
nand U28734 (N_28734,N_28401,N_27698);
or U28735 (N_28735,N_27539,N_27463);
nand U28736 (N_28736,N_27590,N_27212);
xnor U28737 (N_28737,N_27315,N_27768);
xnor U28738 (N_28738,N_27849,N_28232);
or U28739 (N_28739,N_28307,N_28160);
and U28740 (N_28740,N_28417,N_27046);
and U28741 (N_28741,N_27970,N_28107);
or U28742 (N_28742,N_28265,N_27165);
nor U28743 (N_28743,N_27967,N_28109);
nor U28744 (N_28744,N_27360,N_27249);
or U28745 (N_28745,N_27279,N_27274);
nand U28746 (N_28746,N_27848,N_28104);
or U28747 (N_28747,N_28069,N_27619);
xor U28748 (N_28748,N_27602,N_27936);
nand U28749 (N_28749,N_27314,N_28422);
nand U28750 (N_28750,N_27114,N_27663);
nor U28751 (N_28751,N_27235,N_28385);
nand U28752 (N_28752,N_28261,N_28342);
and U28753 (N_28753,N_28423,N_27675);
or U28754 (N_28754,N_28134,N_28207);
xor U28755 (N_28755,N_27504,N_28263);
and U28756 (N_28756,N_28333,N_27065);
and U28757 (N_28757,N_27198,N_27647);
xnor U28758 (N_28758,N_28184,N_27221);
nor U28759 (N_28759,N_28094,N_27476);
nor U28760 (N_28760,N_27829,N_28306);
and U28761 (N_28761,N_27926,N_27025);
or U28762 (N_28762,N_27931,N_27238);
nor U28763 (N_28763,N_27540,N_27796);
nor U28764 (N_28764,N_27811,N_27261);
xor U28765 (N_28765,N_27371,N_27615);
xnor U28766 (N_28766,N_27128,N_27526);
xnor U28767 (N_28767,N_28034,N_27522);
xor U28768 (N_28768,N_28095,N_27012);
nand U28769 (N_28769,N_28471,N_27097);
nor U28770 (N_28770,N_27824,N_28317);
xor U28771 (N_28771,N_27865,N_27655);
and U28772 (N_28772,N_27106,N_27658);
nand U28773 (N_28773,N_28292,N_27362);
and U28774 (N_28774,N_28152,N_27828);
xor U28775 (N_28775,N_27217,N_27870);
nand U28776 (N_28776,N_27742,N_27427);
and U28777 (N_28777,N_27023,N_28173);
nand U28778 (N_28778,N_28097,N_27620);
xor U28779 (N_28779,N_28288,N_27017);
nor U28780 (N_28780,N_27534,N_27572);
and U28781 (N_28781,N_28361,N_28270);
xor U28782 (N_28782,N_27465,N_27491);
nand U28783 (N_28783,N_27804,N_27966);
nor U28784 (N_28784,N_27339,N_28382);
or U28785 (N_28785,N_27527,N_27131);
nand U28786 (N_28786,N_27086,N_28192);
nand U28787 (N_28787,N_27554,N_27517);
or U28788 (N_28788,N_28164,N_27598);
nor U28789 (N_28789,N_28026,N_27383);
xor U28790 (N_28790,N_28360,N_27057);
and U28791 (N_28791,N_27545,N_27400);
or U28792 (N_28792,N_27681,N_28006);
xnor U28793 (N_28793,N_28355,N_27098);
and U28794 (N_28794,N_27390,N_28139);
xor U28795 (N_28795,N_27567,N_28111);
or U28796 (N_28796,N_27355,N_28201);
or U28797 (N_28797,N_27382,N_27327);
and U28798 (N_28798,N_27307,N_27909);
or U28799 (N_28799,N_28128,N_28047);
nand U28800 (N_28800,N_28027,N_28010);
and U28801 (N_28801,N_27194,N_28420);
or U28802 (N_28802,N_28234,N_27135);
or U28803 (N_28803,N_27565,N_28276);
nor U28804 (N_28804,N_28405,N_27214);
nand U28805 (N_28805,N_27070,N_27241);
xnor U28806 (N_28806,N_27345,N_27802);
and U28807 (N_28807,N_28044,N_27246);
nor U28808 (N_28808,N_28000,N_27499);
and U28809 (N_28809,N_27898,N_28358);
nor U28810 (N_28810,N_28415,N_28066);
nand U28811 (N_28811,N_27547,N_27054);
xnor U28812 (N_28812,N_27291,N_27789);
nand U28813 (N_28813,N_27494,N_27156);
nor U28814 (N_28814,N_28274,N_28364);
or U28815 (N_28815,N_28338,N_27969);
xnor U28816 (N_28816,N_28301,N_27818);
xnor U28817 (N_28817,N_28442,N_27296);
xnor U28818 (N_28818,N_28169,N_27786);
nand U28819 (N_28819,N_27453,N_27171);
xnor U28820 (N_28820,N_27393,N_27304);
nand U28821 (N_28821,N_27263,N_28185);
nor U28822 (N_28822,N_28093,N_27042);
and U28823 (N_28823,N_28287,N_27473);
nand U28824 (N_28824,N_27414,N_27468);
or U28825 (N_28825,N_28331,N_28179);
nand U28826 (N_28826,N_28387,N_27634);
nor U28827 (N_28827,N_27265,N_27208);
xor U28828 (N_28828,N_27466,N_27301);
nand U28829 (N_28829,N_28452,N_28388);
nand U28830 (N_28830,N_28374,N_28316);
xor U28831 (N_28831,N_27254,N_27904);
and U28832 (N_28832,N_28334,N_27694);
xor U28833 (N_28833,N_28264,N_28021);
xnor U28834 (N_28834,N_27894,N_28118);
and U28835 (N_28835,N_27730,N_28403);
nand U28836 (N_28836,N_27434,N_27791);
xnor U28837 (N_28837,N_27432,N_27978);
or U28838 (N_28838,N_28302,N_27357);
nor U28839 (N_28839,N_27622,N_27100);
nor U28840 (N_28840,N_28455,N_28282);
and U28841 (N_28841,N_28380,N_27794);
nand U28842 (N_28842,N_27404,N_27372);
nor U28843 (N_28843,N_27591,N_28099);
and U28844 (N_28844,N_27928,N_27071);
nand U28845 (N_28845,N_27094,N_27721);
nand U28846 (N_28846,N_27972,N_28088);
or U28847 (N_28847,N_27939,N_28356);
and U28848 (N_28848,N_27759,N_27696);
xor U28849 (N_28849,N_27760,N_28129);
xor U28850 (N_28850,N_27693,N_28396);
nand U28851 (N_28851,N_27703,N_28434);
or U28852 (N_28852,N_28431,N_27403);
nor U28853 (N_28853,N_28245,N_27885);
xnor U28854 (N_28854,N_28091,N_28314);
nor U28855 (N_28855,N_28328,N_28011);
nand U28856 (N_28856,N_27775,N_27083);
xor U28857 (N_28857,N_27440,N_27503);
or U28858 (N_28858,N_27278,N_27297);
or U28859 (N_28859,N_27852,N_27144);
nand U28860 (N_28860,N_27650,N_28165);
nor U28861 (N_28861,N_27510,N_27584);
nand U28862 (N_28862,N_27726,N_27435);
xor U28863 (N_28863,N_27112,N_27234);
or U28864 (N_28864,N_27078,N_27180);
or U28865 (N_28865,N_27661,N_27055);
nand U28866 (N_28866,N_27851,N_27088);
nand U28867 (N_28867,N_28448,N_27793);
or U28868 (N_28868,N_28472,N_27064);
nand U28869 (N_28869,N_28080,N_28318);
nand U28870 (N_28870,N_27582,N_27168);
or U28871 (N_28871,N_28391,N_27478);
xnor U28872 (N_28872,N_27930,N_28190);
nor U28873 (N_28873,N_27878,N_28105);
or U28874 (N_28874,N_27975,N_28428);
nor U28875 (N_28875,N_27938,N_27922);
and U28876 (N_28876,N_27523,N_27483);
nor U28877 (N_28877,N_27659,N_27003);
xor U28878 (N_28878,N_27442,N_27101);
or U28879 (N_28879,N_27202,N_27337);
or U28880 (N_28880,N_27843,N_27457);
xnor U28881 (N_28881,N_28437,N_28130);
xnor U28882 (N_28882,N_28389,N_27232);
or U28883 (N_28883,N_27201,N_28424);
or U28884 (N_28884,N_28375,N_27809);
or U28885 (N_28885,N_27623,N_27918);
or U28886 (N_28886,N_28432,N_27908);
and U28887 (N_28887,N_27674,N_27306);
nand U28888 (N_28888,N_27562,N_27325);
nor U28889 (N_28889,N_28295,N_27697);
nor U28890 (N_28890,N_27986,N_27060);
or U28891 (N_28891,N_28020,N_27495);
and U28892 (N_28892,N_27860,N_27636);
nand U28893 (N_28893,N_27531,N_28426);
or U28894 (N_28894,N_27544,N_27589);
or U28895 (N_28895,N_27139,N_28057);
and U28896 (N_28896,N_27389,N_27979);
and U28897 (N_28897,N_28078,N_28249);
and U28898 (N_28898,N_27058,N_27530);
or U28899 (N_28899,N_28491,N_28315);
or U28900 (N_28900,N_27500,N_28430);
nand U28901 (N_28901,N_28056,N_27644);
and U28902 (N_28902,N_28371,N_27014);
nor U28903 (N_28903,N_27075,N_27481);
xnor U28904 (N_28904,N_27018,N_27781);
nand U28905 (N_28905,N_28290,N_27321);
nand U28906 (N_28906,N_28341,N_27020);
xor U28907 (N_28907,N_27932,N_28377);
nor U28908 (N_28908,N_28189,N_27773);
or U28909 (N_28909,N_27616,N_27676);
and U28910 (N_28910,N_27934,N_27711);
nor U28911 (N_28911,N_27950,N_27713);
or U28912 (N_28912,N_27646,N_27053);
and U28913 (N_28913,N_27148,N_27891);
or U28914 (N_28914,N_27351,N_27924);
or U28915 (N_28915,N_27910,N_27679);
nand U28916 (N_28916,N_27556,N_28451);
nor U28917 (N_28917,N_28446,N_27275);
or U28918 (N_28918,N_27318,N_28323);
xnor U28919 (N_28919,N_28036,N_27633);
and U28920 (N_28920,N_27778,N_27971);
nand U28921 (N_28921,N_27231,N_28043);
xor U28922 (N_28922,N_28359,N_27153);
nand U28923 (N_28923,N_28397,N_27604);
or U28924 (N_28924,N_27999,N_27905);
xnor U28925 (N_28925,N_27287,N_28102);
and U28926 (N_28926,N_28174,N_27955);
and U28927 (N_28927,N_27776,N_27875);
and U28928 (N_28928,N_27095,N_27649);
nor U28929 (N_28929,N_27074,N_28200);
nor U28930 (N_28930,N_27401,N_27323);
nor U28931 (N_28931,N_27533,N_27734);
or U28932 (N_28932,N_27929,N_28237);
nor U28933 (N_28933,N_28335,N_28354);
nor U28934 (N_28934,N_27250,N_27716);
xnor U28935 (N_28935,N_27348,N_27108);
nor U28936 (N_28936,N_27667,N_27594);
nand U28937 (N_28937,N_27039,N_27551);
or U28938 (N_28938,N_27838,N_28329);
nor U28939 (N_28939,N_28121,N_28230);
xnor U28940 (N_28940,N_28480,N_27284);
xor U28941 (N_28941,N_27282,N_28073);
and U28942 (N_28942,N_27883,N_28466);
nand U28943 (N_28943,N_27488,N_28126);
and U28944 (N_28944,N_27771,N_27176);
or U28945 (N_28945,N_27702,N_27831);
and U28946 (N_28946,N_27482,N_27751);
xnor U28947 (N_28947,N_27264,N_27245);
nand U28948 (N_28948,N_28197,N_28054);
xor U28949 (N_28949,N_27384,N_27193);
nand U28950 (N_28950,N_27763,N_27991);
or U28951 (N_28951,N_27614,N_27945);
and U28952 (N_28952,N_27748,N_28223);
nand U28953 (N_28953,N_28156,N_27982);
nor U28954 (N_28954,N_27800,N_27438);
nand U28955 (N_28955,N_27016,N_27358);
or U28956 (N_28956,N_27364,N_27782);
or U28957 (N_28957,N_28208,N_28258);
or U28958 (N_28958,N_27558,N_28133);
nand U28959 (N_28959,N_28425,N_27683);
or U28960 (N_28960,N_28023,N_27160);
and U28961 (N_28961,N_27884,N_27954);
or U28962 (N_28962,N_27056,N_27419);
or U28963 (N_28963,N_27125,N_28124);
nor U28964 (N_28964,N_28101,N_27158);
nand U28965 (N_28965,N_28242,N_27177);
nor U28966 (N_28966,N_28252,N_28330);
nand U28967 (N_28967,N_28188,N_28477);
or U28968 (N_28968,N_27385,N_27958);
nand U28969 (N_28969,N_27381,N_28456);
nand U28970 (N_28970,N_27354,N_27965);
and U28971 (N_28971,N_28132,N_28067);
or U28972 (N_28972,N_28149,N_27845);
nand U28973 (N_28973,N_27731,N_28176);
nor U28974 (N_28974,N_28059,N_28254);
or U28975 (N_28975,N_27133,N_27082);
and U28976 (N_28976,N_27155,N_27612);
nand U28977 (N_28977,N_28186,N_28291);
xor U28978 (N_28978,N_27205,N_27352);
or U28979 (N_28979,N_28092,N_27941);
xnor U28980 (N_28980,N_27854,N_28072);
nor U28981 (N_28981,N_27361,N_28365);
or U28982 (N_28982,N_27146,N_28150);
nand U28983 (N_28983,N_27630,N_28493);
and U28984 (N_28984,N_28497,N_27976);
or U28985 (N_28985,N_27508,N_27061);
nor U28986 (N_28986,N_28025,N_27183);
or U28987 (N_28987,N_28038,N_28194);
and U28988 (N_28988,N_27563,N_27837);
xnor U28989 (N_28989,N_28409,N_28089);
xnor U28990 (N_28990,N_28019,N_27874);
or U28991 (N_28991,N_27801,N_27528);
xor U28992 (N_28992,N_27031,N_28272);
xor U28993 (N_28993,N_27256,N_27576);
and U28994 (N_28994,N_27066,N_27635);
nand U28995 (N_28995,N_27807,N_27113);
or U28996 (N_28996,N_28412,N_27968);
nand U28997 (N_28997,N_27380,N_27191);
and U28998 (N_28998,N_27397,N_27601);
xnor U28999 (N_28999,N_27216,N_27027);
nand U29000 (N_29000,N_27678,N_27298);
or U29001 (N_29001,N_28485,N_27515);
xnor U29002 (N_29002,N_28321,N_27593);
nor U29003 (N_29003,N_27743,N_27723);
or U29004 (N_29004,N_27210,N_28304);
nor U29005 (N_29005,N_27309,N_27472);
or U29006 (N_29006,N_28357,N_27283);
nand U29007 (N_29007,N_27993,N_27149);
xnor U29008 (N_29008,N_27677,N_27022);
or U29009 (N_29009,N_28125,N_27592);
nor U29010 (N_29010,N_28284,N_28332);
or U29011 (N_29011,N_28266,N_27161);
xor U29012 (N_29012,N_27271,N_28467);
or U29013 (N_29013,N_27735,N_27142);
nand U29014 (N_29014,N_28244,N_27035);
nand U29015 (N_29015,N_27312,N_27223);
nand U29016 (N_29016,N_28445,N_27588);
or U29017 (N_29017,N_28303,N_27152);
xor U29018 (N_29018,N_27242,N_28198);
or U29019 (N_29019,N_28220,N_27239);
and U29020 (N_29020,N_28181,N_27172);
nor U29021 (N_29021,N_27561,N_27426);
and U29022 (N_29022,N_27288,N_28337);
xnor U29023 (N_29023,N_28351,N_27869);
and U29024 (N_29024,N_27405,N_27750);
xor U29025 (N_29025,N_27925,N_27051);
xor U29026 (N_29026,N_27489,N_28309);
xnor U29027 (N_29027,N_27770,N_27597);
xor U29028 (N_29028,N_27029,N_27129);
and U29029 (N_29029,N_27391,N_27163);
or U29030 (N_29030,N_28441,N_27625);
nor U29031 (N_29031,N_27892,N_27179);
nor U29032 (N_29032,N_27445,N_28478);
or U29033 (N_29033,N_27138,N_28029);
nor U29034 (N_29034,N_27273,N_27631);
xnor U29035 (N_29035,N_28395,N_27777);
and U29036 (N_29036,N_28172,N_27356);
xor U29037 (N_29037,N_27233,N_28037);
or U29038 (N_29038,N_28048,N_27783);
or U29039 (N_29039,N_28363,N_27998);
xnor U29040 (N_29040,N_28449,N_28496);
nand U29041 (N_29041,N_28475,N_28271);
or U29042 (N_29042,N_27169,N_27040);
nor U29043 (N_29043,N_27541,N_28214);
nand U29044 (N_29044,N_28002,N_27570);
or U29045 (N_29045,N_28327,N_27946);
nand U29046 (N_29046,N_28063,N_28110);
and U29047 (N_29047,N_27406,N_28141);
and U29048 (N_29048,N_28183,N_27310);
nand U29049 (N_29049,N_27953,N_27609);
xor U29050 (N_29050,N_27501,N_27431);
xnor U29051 (N_29051,N_28320,N_27377);
or U29052 (N_29052,N_27714,N_27353);
nor U29053 (N_29053,N_27888,N_27810);
nor U29054 (N_29054,N_27956,N_27236);
nand U29055 (N_29055,N_28113,N_27836);
or U29056 (N_29056,N_27181,N_27280);
and U29057 (N_29057,N_27532,N_27038);
and U29058 (N_29058,N_27749,N_27164);
nand U29059 (N_29059,N_28427,N_28070);
nor U29060 (N_29060,N_27825,N_27673);
nor U29061 (N_29061,N_28347,N_27015);
and U29062 (N_29062,N_27853,N_27373);
xor U29063 (N_29063,N_27173,N_28079);
xnor U29064 (N_29064,N_27316,N_27912);
xor U29065 (N_29065,N_27341,N_28086);
xnor U29066 (N_29066,N_27047,N_27103);
and U29067 (N_29067,N_27535,N_28494);
and U29068 (N_29068,N_27105,N_27492);
or U29069 (N_29069,N_27394,N_27542);
nand U29070 (N_29070,N_27779,N_28370);
nand U29071 (N_29071,N_28112,N_28255);
and U29072 (N_29072,N_27569,N_27277);
xor U29073 (N_29073,N_28157,N_27506);
nor U29074 (N_29074,N_27244,N_28239);
nor U29075 (N_29075,N_28240,N_28039);
and U29076 (N_29076,N_28199,N_27839);
or U29077 (N_29077,N_27019,N_27651);
and U29078 (N_29078,N_27859,N_27948);
nor U29079 (N_29079,N_27266,N_27059);
or U29080 (N_29080,N_28344,N_27441);
xor U29081 (N_29081,N_28138,N_27662);
nand U29082 (N_29082,N_27850,N_27276);
or U29083 (N_29083,N_28366,N_27992);
nand U29084 (N_29084,N_28142,N_28279);
nand U29085 (N_29085,N_27175,N_28392);
xor U29086 (N_29086,N_27660,N_27826);
and U29087 (N_29087,N_28052,N_28443);
xnor U29088 (N_29088,N_28135,N_27258);
xor U29089 (N_29089,N_27834,N_27733);
or U29090 (N_29090,N_27374,N_28419);
nand U29091 (N_29091,N_28085,N_27536);
and U29092 (N_29092,N_27331,N_27856);
or U29093 (N_29093,N_28350,N_27973);
or U29094 (N_29094,N_27392,N_27692);
and U29095 (N_29095,N_27599,N_28123);
xnor U29096 (N_29096,N_27437,N_27617);
nor U29097 (N_29097,N_27666,N_28137);
or U29098 (N_29098,N_27007,N_27359);
and U29099 (N_29099,N_27116,N_27127);
nand U29100 (N_29100,N_27632,N_27228);
xnor U29101 (N_29101,N_27207,N_28386);
and U29102 (N_29102,N_27036,N_27436);
and U29103 (N_29103,N_27900,N_27219);
xnor U29104 (N_29104,N_28390,N_27230);
and U29105 (N_29105,N_27447,N_28215);
xnor U29106 (N_29106,N_27460,N_27705);
or U29107 (N_29107,N_27220,N_27901);
and U29108 (N_29108,N_27691,N_27820);
xnor U29109 (N_29109,N_27521,N_27030);
nand U29110 (N_29110,N_28106,N_27833);
nor U29111 (N_29111,N_27338,N_27458);
and U29112 (N_29112,N_28433,N_27983);
nand U29113 (N_29113,N_28367,N_27943);
and U29114 (N_29114,N_28490,N_27668);
and U29115 (N_29115,N_27895,N_27350);
and U29116 (N_29116,N_27564,N_27719);
nor U29117 (N_29117,N_28406,N_27618);
nand U29118 (N_29118,N_28007,N_27761);
nor U29119 (N_29119,N_28008,N_27844);
xnor U29120 (N_29120,N_27727,N_27764);
nor U29121 (N_29121,N_27451,N_28147);
and U29122 (N_29122,N_27863,N_27756);
xnor U29123 (N_29123,N_27429,N_28100);
xnor U29124 (N_29124,N_27137,N_28275);
xor U29125 (N_29125,N_27737,N_27395);
xor U29126 (N_29126,N_27546,N_27785);
or U29127 (N_29127,N_28414,N_28206);
and U29128 (N_29128,N_28227,N_28248);
or U29129 (N_29129,N_27717,N_27980);
and U29130 (N_29130,N_28154,N_27816);
nor U29131 (N_29131,N_28372,N_27456);
and U29132 (N_29132,N_28076,N_27645);
or U29133 (N_29133,N_28238,N_27552);
nand U29134 (N_29134,N_27026,N_27538);
nor U29135 (N_29135,N_27317,N_27486);
or U29136 (N_29136,N_27806,N_28243);
nand U29137 (N_29137,N_28193,N_27237);
xor U29138 (N_29138,N_27637,N_27425);
and U29139 (N_29139,N_27574,N_27913);
nor U29140 (N_29140,N_27571,N_27084);
nor U29141 (N_29141,N_28418,N_27628);
nor U29142 (N_29142,N_28486,N_27464);
nand U29143 (N_29143,N_27072,N_27754);
or U29144 (N_29144,N_27525,N_28469);
nand U29145 (N_29145,N_27111,N_28325);
and U29146 (N_29146,N_27981,N_27670);
or U29147 (N_29147,N_27708,N_28046);
xnor U29148 (N_29148,N_27920,N_28241);
and U29149 (N_29149,N_27006,N_27366);
and U29150 (N_29150,N_28345,N_27093);
or U29151 (N_29151,N_27028,N_27603);
xor U29152 (N_29152,N_27560,N_28013);
nand U29153 (N_29153,N_28178,N_28210);
nand U29154 (N_29154,N_27502,N_28061);
and U29155 (N_29155,N_27903,N_27409);
nand U29156 (N_29156,N_28062,N_27911);
nand U29157 (N_29157,N_28087,N_27450);
xnor U29158 (N_29158,N_28083,N_27154);
or U29159 (N_29159,N_28018,N_27987);
or U29160 (N_29160,N_28005,N_27867);
and U29161 (N_29161,N_27709,N_27068);
or U29162 (N_29162,N_27424,N_27654);
and U29163 (N_29163,N_27942,N_27229);
nor U29164 (N_29164,N_27813,N_28464);
or U29165 (N_29165,N_27454,N_28378);
or U29166 (N_29166,N_27368,N_28394);
nor U29167 (N_29167,N_28339,N_28399);
nand U29168 (N_29168,N_27262,N_27740);
xnor U29169 (N_29169,N_27739,N_27767);
nor U29170 (N_29170,N_27209,N_27444);
xnor U29171 (N_29171,N_27126,N_28402);
xor U29172 (N_29172,N_27573,N_28151);
or U29173 (N_29173,N_28084,N_27682);
or U29174 (N_29174,N_28460,N_27745);
nand U29175 (N_29175,N_27520,N_27757);
nor U29176 (N_29176,N_27240,N_27416);
and U29177 (N_29177,N_28468,N_28461);
xor U29178 (N_29178,N_28353,N_27877);
nand U29179 (N_29179,N_28213,N_27578);
nor U29180 (N_29180,N_27349,N_27830);
xor U29181 (N_29181,N_28163,N_27272);
or U29182 (N_29182,N_27861,N_28155);
and U29183 (N_29183,N_27182,N_28120);
and U29184 (N_29184,N_28122,N_27706);
nor U29185 (N_29185,N_28014,N_27803);
or U29186 (N_29186,N_27559,N_27470);
or U29187 (N_29187,N_27224,N_27326);
xor U29188 (N_29188,N_27243,N_27048);
xnor U29189 (N_29189,N_28308,N_27606);
nor U29190 (N_29190,N_27067,N_27009);
nand U29191 (N_29191,N_28167,N_27461);
xnor U29192 (N_29192,N_28212,N_27919);
nand U29193 (N_29193,N_27947,N_27758);
or U29194 (N_29194,N_27449,N_27081);
nor U29195 (N_29195,N_28482,N_28300);
nor U29196 (N_29196,N_27577,N_27927);
nor U29197 (N_29197,N_28218,N_28103);
nand U29198 (N_29198,N_27704,N_28009);
and U29199 (N_29199,N_27439,N_27664);
nor U29200 (N_29200,N_27624,N_27388);
nand U29201 (N_29201,N_27199,N_27519);
or U29202 (N_29202,N_27011,N_27548);
and U29203 (N_29203,N_27935,N_28030);
nand U29204 (N_29204,N_28235,N_28108);
and U29205 (N_29205,N_28096,N_27514);
xnor U29206 (N_29206,N_27347,N_27720);
nor U29207 (N_29207,N_28348,N_28267);
nand U29208 (N_29208,N_27328,N_28115);
nand U29209 (N_29209,N_28191,N_27695);
xor U29210 (N_29210,N_27685,N_28246);
xnor U29211 (N_29211,N_27396,N_27795);
or U29212 (N_29212,N_27211,N_27715);
or U29213 (N_29213,N_27940,N_27890);
nand U29214 (N_29214,N_27512,N_27868);
nand U29215 (N_29215,N_27002,N_27413);
or U29216 (N_29216,N_28162,N_28470);
and U29217 (N_29217,N_28196,N_28117);
nand U29218 (N_29218,N_27600,N_27690);
or U29219 (N_29219,N_28116,N_28175);
xnor U29220 (N_29220,N_27398,N_28326);
and U29221 (N_29221,N_27566,N_27140);
or U29222 (N_29222,N_27032,N_28127);
nor U29223 (N_29223,N_28313,N_28055);
nand U29224 (N_29224,N_27034,N_27921);
nor U29225 (N_29225,N_27671,N_28228);
or U29226 (N_29226,N_27147,N_27808);
nand U29227 (N_29227,N_28144,N_27222);
and U29228 (N_29228,N_28031,N_28465);
nand U29229 (N_29229,N_27281,N_27099);
xnor U29230 (N_29230,N_27062,N_27151);
and U29231 (N_29231,N_27363,N_27102);
xor U29232 (N_29232,N_28145,N_27996);
or U29233 (N_29233,N_28400,N_28407);
or U29234 (N_29234,N_28182,N_28346);
or U29235 (N_29235,N_27334,N_27866);
or U29236 (N_29236,N_28166,N_28458);
nand U29237 (N_29237,N_28022,N_28285);
and U29238 (N_29238,N_27407,N_27815);
nand U29239 (N_29239,N_27344,N_27805);
xor U29240 (N_29240,N_27627,N_27513);
nand U29241 (N_29241,N_27480,N_27961);
xor U29242 (N_29242,N_28221,N_28205);
nand U29243 (N_29243,N_27496,N_27001);
xor U29244 (N_29244,N_27063,N_27896);
nor U29245 (N_29245,N_27984,N_27822);
xor U29246 (N_29246,N_27286,N_27024);
or U29247 (N_29247,N_27847,N_27917);
nand U29248 (N_29248,N_27916,N_27842);
and U29249 (N_29249,N_27944,N_27656);
and U29250 (N_29250,N_28263,N_27619);
or U29251 (N_29251,N_28419,N_27786);
nor U29252 (N_29252,N_28252,N_28492);
nand U29253 (N_29253,N_27598,N_28370);
or U29254 (N_29254,N_27464,N_28165);
or U29255 (N_29255,N_27502,N_28131);
xnor U29256 (N_29256,N_27717,N_27554);
nand U29257 (N_29257,N_28187,N_28053);
or U29258 (N_29258,N_27196,N_27679);
xor U29259 (N_29259,N_27204,N_27851);
xor U29260 (N_29260,N_27887,N_27412);
or U29261 (N_29261,N_27540,N_28157);
nor U29262 (N_29262,N_27287,N_27325);
nor U29263 (N_29263,N_28062,N_28211);
and U29264 (N_29264,N_27968,N_28416);
and U29265 (N_29265,N_28372,N_27190);
nor U29266 (N_29266,N_28390,N_27249);
xnor U29267 (N_29267,N_27392,N_28483);
and U29268 (N_29268,N_28127,N_27484);
or U29269 (N_29269,N_27637,N_27330);
or U29270 (N_29270,N_27727,N_28099);
and U29271 (N_29271,N_27488,N_28200);
or U29272 (N_29272,N_27096,N_27152);
nor U29273 (N_29273,N_27372,N_27878);
nor U29274 (N_29274,N_27139,N_27060);
nand U29275 (N_29275,N_28403,N_27381);
and U29276 (N_29276,N_28136,N_27960);
or U29277 (N_29277,N_27771,N_27131);
and U29278 (N_29278,N_27094,N_27609);
xor U29279 (N_29279,N_28329,N_28462);
xnor U29280 (N_29280,N_27251,N_28300);
xor U29281 (N_29281,N_28433,N_27834);
or U29282 (N_29282,N_27716,N_27121);
and U29283 (N_29283,N_27859,N_27939);
or U29284 (N_29284,N_27986,N_27666);
xor U29285 (N_29285,N_27706,N_27600);
or U29286 (N_29286,N_27210,N_27939);
xor U29287 (N_29287,N_28282,N_27487);
and U29288 (N_29288,N_27179,N_27836);
and U29289 (N_29289,N_28388,N_28448);
or U29290 (N_29290,N_27111,N_28049);
nor U29291 (N_29291,N_28051,N_27160);
or U29292 (N_29292,N_28452,N_27070);
or U29293 (N_29293,N_27594,N_27928);
and U29294 (N_29294,N_28267,N_28113);
xor U29295 (N_29295,N_28039,N_27704);
xor U29296 (N_29296,N_27072,N_27506);
xor U29297 (N_29297,N_27131,N_27696);
and U29298 (N_29298,N_27616,N_27344);
and U29299 (N_29299,N_27343,N_27997);
and U29300 (N_29300,N_27987,N_27623);
and U29301 (N_29301,N_27845,N_27992);
xor U29302 (N_29302,N_28396,N_27592);
or U29303 (N_29303,N_27761,N_27477);
and U29304 (N_29304,N_27697,N_27799);
nor U29305 (N_29305,N_28231,N_28079);
nor U29306 (N_29306,N_27340,N_27271);
nor U29307 (N_29307,N_28339,N_27683);
or U29308 (N_29308,N_27196,N_27786);
or U29309 (N_29309,N_28485,N_27660);
nor U29310 (N_29310,N_27191,N_27561);
or U29311 (N_29311,N_28319,N_28091);
xnor U29312 (N_29312,N_27252,N_27983);
and U29313 (N_29313,N_27205,N_27775);
or U29314 (N_29314,N_28262,N_27835);
nand U29315 (N_29315,N_27267,N_28319);
or U29316 (N_29316,N_27187,N_27757);
nor U29317 (N_29317,N_27001,N_28410);
nand U29318 (N_29318,N_27845,N_27936);
or U29319 (N_29319,N_27089,N_27480);
or U29320 (N_29320,N_28163,N_27844);
or U29321 (N_29321,N_27857,N_28028);
or U29322 (N_29322,N_27187,N_27490);
or U29323 (N_29323,N_28478,N_27859);
xnor U29324 (N_29324,N_28152,N_27747);
nand U29325 (N_29325,N_27138,N_28107);
or U29326 (N_29326,N_28499,N_27321);
and U29327 (N_29327,N_27734,N_27462);
nor U29328 (N_29328,N_27268,N_27837);
nor U29329 (N_29329,N_28143,N_27679);
or U29330 (N_29330,N_27884,N_27857);
and U29331 (N_29331,N_28467,N_28019);
nand U29332 (N_29332,N_27218,N_28036);
nand U29333 (N_29333,N_28173,N_27325);
and U29334 (N_29334,N_27849,N_27659);
nor U29335 (N_29335,N_28483,N_27371);
or U29336 (N_29336,N_27326,N_28253);
nor U29337 (N_29337,N_27332,N_27886);
nand U29338 (N_29338,N_28263,N_28137);
nor U29339 (N_29339,N_28133,N_27796);
and U29340 (N_29340,N_27198,N_28487);
nor U29341 (N_29341,N_27766,N_28089);
xor U29342 (N_29342,N_28407,N_27118);
nor U29343 (N_29343,N_28394,N_27231);
or U29344 (N_29344,N_27850,N_27026);
nand U29345 (N_29345,N_27171,N_28085);
nor U29346 (N_29346,N_27618,N_28047);
xor U29347 (N_29347,N_28276,N_27193);
nand U29348 (N_29348,N_28193,N_28179);
and U29349 (N_29349,N_27288,N_27878);
xor U29350 (N_29350,N_27580,N_27385);
nand U29351 (N_29351,N_27908,N_27029);
and U29352 (N_29352,N_27841,N_27447);
nand U29353 (N_29353,N_27276,N_28399);
nand U29354 (N_29354,N_28472,N_28073);
xor U29355 (N_29355,N_28268,N_28228);
or U29356 (N_29356,N_28182,N_27037);
or U29357 (N_29357,N_27311,N_27088);
and U29358 (N_29358,N_27109,N_27917);
nor U29359 (N_29359,N_28151,N_28379);
nor U29360 (N_29360,N_28462,N_27928);
and U29361 (N_29361,N_28060,N_28232);
and U29362 (N_29362,N_27281,N_28263);
or U29363 (N_29363,N_28329,N_27259);
nand U29364 (N_29364,N_27552,N_27292);
nand U29365 (N_29365,N_27665,N_27460);
and U29366 (N_29366,N_28372,N_28311);
nor U29367 (N_29367,N_27681,N_28068);
xor U29368 (N_29368,N_28077,N_28115);
and U29369 (N_29369,N_27410,N_28160);
nor U29370 (N_29370,N_28380,N_27209);
xnor U29371 (N_29371,N_27611,N_27182);
or U29372 (N_29372,N_27578,N_28366);
nor U29373 (N_29373,N_27957,N_27298);
nor U29374 (N_29374,N_27774,N_28073);
nor U29375 (N_29375,N_27648,N_27035);
xor U29376 (N_29376,N_27115,N_27641);
nand U29377 (N_29377,N_27956,N_27997);
xor U29378 (N_29378,N_27371,N_27557);
and U29379 (N_29379,N_27867,N_28359);
nand U29380 (N_29380,N_27803,N_28237);
xnor U29381 (N_29381,N_27010,N_27067);
nor U29382 (N_29382,N_27513,N_27723);
or U29383 (N_29383,N_27949,N_27816);
nand U29384 (N_29384,N_27902,N_28338);
and U29385 (N_29385,N_28453,N_27387);
nand U29386 (N_29386,N_27953,N_27399);
xnor U29387 (N_29387,N_27420,N_27332);
xor U29388 (N_29388,N_27881,N_27221);
xor U29389 (N_29389,N_27937,N_27659);
or U29390 (N_29390,N_27023,N_27556);
and U29391 (N_29391,N_27806,N_27548);
nand U29392 (N_29392,N_27791,N_27595);
nand U29393 (N_29393,N_27744,N_28054);
xnor U29394 (N_29394,N_27802,N_28456);
and U29395 (N_29395,N_27116,N_27840);
and U29396 (N_29396,N_27841,N_27244);
nand U29397 (N_29397,N_28338,N_27310);
and U29398 (N_29398,N_27979,N_28404);
nand U29399 (N_29399,N_28442,N_27934);
and U29400 (N_29400,N_27185,N_27961);
nor U29401 (N_29401,N_27138,N_27464);
or U29402 (N_29402,N_27693,N_27894);
or U29403 (N_29403,N_27176,N_28022);
and U29404 (N_29404,N_27627,N_27794);
or U29405 (N_29405,N_28399,N_27938);
and U29406 (N_29406,N_27834,N_27712);
and U29407 (N_29407,N_28484,N_28238);
and U29408 (N_29408,N_28248,N_27610);
or U29409 (N_29409,N_28201,N_28236);
nand U29410 (N_29410,N_27653,N_28365);
nor U29411 (N_29411,N_28085,N_27253);
or U29412 (N_29412,N_27201,N_28177);
nor U29413 (N_29413,N_27196,N_28103);
nor U29414 (N_29414,N_27613,N_27493);
xnor U29415 (N_29415,N_27474,N_28464);
nand U29416 (N_29416,N_28071,N_28272);
xnor U29417 (N_29417,N_27436,N_28170);
xor U29418 (N_29418,N_27670,N_27321);
and U29419 (N_29419,N_28128,N_28271);
and U29420 (N_29420,N_27300,N_28360);
xnor U29421 (N_29421,N_28495,N_27684);
and U29422 (N_29422,N_27298,N_28496);
nand U29423 (N_29423,N_28126,N_27706);
or U29424 (N_29424,N_27178,N_28002);
or U29425 (N_29425,N_28357,N_28331);
nor U29426 (N_29426,N_27748,N_27843);
or U29427 (N_29427,N_28258,N_27813);
xnor U29428 (N_29428,N_28258,N_27143);
xor U29429 (N_29429,N_28462,N_28292);
or U29430 (N_29430,N_27930,N_27251);
nand U29431 (N_29431,N_27613,N_28161);
xor U29432 (N_29432,N_27020,N_27680);
xnor U29433 (N_29433,N_27907,N_28217);
or U29434 (N_29434,N_27718,N_27102);
and U29435 (N_29435,N_27901,N_27110);
xor U29436 (N_29436,N_28290,N_28309);
and U29437 (N_29437,N_27139,N_28478);
or U29438 (N_29438,N_27013,N_27221);
or U29439 (N_29439,N_27842,N_27179);
nand U29440 (N_29440,N_27905,N_27167);
or U29441 (N_29441,N_28008,N_27143);
or U29442 (N_29442,N_27914,N_27468);
xnor U29443 (N_29443,N_28310,N_27108);
or U29444 (N_29444,N_27225,N_27160);
and U29445 (N_29445,N_28239,N_27137);
xor U29446 (N_29446,N_27177,N_27314);
nor U29447 (N_29447,N_28162,N_27325);
nand U29448 (N_29448,N_27122,N_27508);
or U29449 (N_29449,N_27181,N_28221);
or U29450 (N_29450,N_27582,N_28283);
nor U29451 (N_29451,N_28248,N_28362);
nand U29452 (N_29452,N_27697,N_27854);
or U29453 (N_29453,N_27788,N_28135);
and U29454 (N_29454,N_27788,N_27711);
or U29455 (N_29455,N_27739,N_28286);
nor U29456 (N_29456,N_27081,N_27699);
and U29457 (N_29457,N_27763,N_27584);
xor U29458 (N_29458,N_27443,N_28201);
xor U29459 (N_29459,N_27538,N_27750);
and U29460 (N_29460,N_27895,N_28258);
nand U29461 (N_29461,N_28465,N_28372);
nor U29462 (N_29462,N_28430,N_27137);
xnor U29463 (N_29463,N_27959,N_27495);
xnor U29464 (N_29464,N_27579,N_27834);
nand U29465 (N_29465,N_28420,N_27853);
and U29466 (N_29466,N_27147,N_28225);
nand U29467 (N_29467,N_27149,N_27019);
or U29468 (N_29468,N_27340,N_27574);
xor U29469 (N_29469,N_27216,N_27504);
and U29470 (N_29470,N_27931,N_27027);
or U29471 (N_29471,N_28077,N_27600);
nand U29472 (N_29472,N_27060,N_27296);
xor U29473 (N_29473,N_27279,N_27255);
and U29474 (N_29474,N_27488,N_27506);
and U29475 (N_29475,N_27690,N_27628);
nand U29476 (N_29476,N_28487,N_27968);
and U29477 (N_29477,N_27696,N_27695);
and U29478 (N_29478,N_27461,N_27959);
xnor U29479 (N_29479,N_27344,N_27641);
nand U29480 (N_29480,N_27761,N_27858);
nor U29481 (N_29481,N_27405,N_27968);
nor U29482 (N_29482,N_28343,N_27322);
and U29483 (N_29483,N_27976,N_27532);
nor U29484 (N_29484,N_28287,N_27456);
nand U29485 (N_29485,N_28426,N_28361);
nor U29486 (N_29486,N_28241,N_28177);
nor U29487 (N_29487,N_28480,N_28028);
nor U29488 (N_29488,N_28466,N_27411);
xor U29489 (N_29489,N_28454,N_28010);
or U29490 (N_29490,N_27547,N_27981);
and U29491 (N_29491,N_27384,N_27143);
or U29492 (N_29492,N_28326,N_27334);
xnor U29493 (N_29493,N_27591,N_27400);
nor U29494 (N_29494,N_27366,N_27219);
xnor U29495 (N_29495,N_27285,N_28164);
nand U29496 (N_29496,N_28322,N_27627);
and U29497 (N_29497,N_28147,N_27074);
nand U29498 (N_29498,N_27389,N_27780);
nand U29499 (N_29499,N_28035,N_28369);
xnor U29500 (N_29500,N_27734,N_27036);
nor U29501 (N_29501,N_27963,N_28369);
nor U29502 (N_29502,N_28165,N_27027);
and U29503 (N_29503,N_27439,N_28009);
xor U29504 (N_29504,N_27703,N_28382);
nor U29505 (N_29505,N_27304,N_28432);
nand U29506 (N_29506,N_28405,N_27751);
nand U29507 (N_29507,N_27445,N_27388);
xnor U29508 (N_29508,N_27105,N_28240);
nor U29509 (N_29509,N_27609,N_27836);
xor U29510 (N_29510,N_27956,N_28392);
xnor U29511 (N_29511,N_28247,N_27268);
nand U29512 (N_29512,N_27669,N_28432);
nor U29513 (N_29513,N_28399,N_27829);
nor U29514 (N_29514,N_28417,N_28054);
xnor U29515 (N_29515,N_27633,N_27285);
nand U29516 (N_29516,N_28294,N_27857);
or U29517 (N_29517,N_27254,N_27441);
nand U29518 (N_29518,N_28476,N_28375);
and U29519 (N_29519,N_27487,N_27634);
xor U29520 (N_29520,N_27889,N_27670);
xor U29521 (N_29521,N_27255,N_27759);
nor U29522 (N_29522,N_27622,N_27276);
nor U29523 (N_29523,N_28046,N_27631);
or U29524 (N_29524,N_27812,N_27409);
and U29525 (N_29525,N_28404,N_27373);
nand U29526 (N_29526,N_28467,N_27321);
or U29527 (N_29527,N_27316,N_27954);
nand U29528 (N_29528,N_27918,N_27514);
or U29529 (N_29529,N_27864,N_27662);
and U29530 (N_29530,N_28289,N_27650);
nor U29531 (N_29531,N_27871,N_27111);
and U29532 (N_29532,N_28417,N_27510);
xnor U29533 (N_29533,N_27409,N_27231);
nor U29534 (N_29534,N_28272,N_27724);
xor U29535 (N_29535,N_27714,N_28153);
or U29536 (N_29536,N_27657,N_27350);
or U29537 (N_29537,N_27608,N_27936);
nand U29538 (N_29538,N_28354,N_27851);
xnor U29539 (N_29539,N_27267,N_27173);
and U29540 (N_29540,N_27906,N_27747);
nor U29541 (N_29541,N_27694,N_27887);
xnor U29542 (N_29542,N_27029,N_27399);
xnor U29543 (N_29543,N_28461,N_28495);
nor U29544 (N_29544,N_27239,N_27105);
nor U29545 (N_29545,N_28306,N_28235);
nor U29546 (N_29546,N_27773,N_27698);
nor U29547 (N_29547,N_28081,N_28181);
xnor U29548 (N_29548,N_27032,N_27729);
and U29549 (N_29549,N_27097,N_27608);
or U29550 (N_29550,N_28164,N_27441);
nor U29551 (N_29551,N_27946,N_27755);
nand U29552 (N_29552,N_28486,N_27423);
nor U29553 (N_29553,N_28424,N_28188);
nor U29554 (N_29554,N_27892,N_27412);
xor U29555 (N_29555,N_27905,N_28187);
nand U29556 (N_29556,N_27879,N_27430);
nor U29557 (N_29557,N_27074,N_28376);
nand U29558 (N_29558,N_27087,N_27854);
and U29559 (N_29559,N_28388,N_28017);
xnor U29560 (N_29560,N_27730,N_28326);
and U29561 (N_29561,N_28150,N_27149);
or U29562 (N_29562,N_27868,N_27867);
nor U29563 (N_29563,N_28274,N_27806);
nand U29564 (N_29564,N_27425,N_27176);
xnor U29565 (N_29565,N_27292,N_28402);
and U29566 (N_29566,N_27972,N_27595);
and U29567 (N_29567,N_27132,N_27792);
or U29568 (N_29568,N_27581,N_27106);
nand U29569 (N_29569,N_27385,N_27852);
nand U29570 (N_29570,N_28494,N_27137);
nand U29571 (N_29571,N_27518,N_27649);
nand U29572 (N_29572,N_28280,N_27435);
nor U29573 (N_29573,N_27456,N_28330);
xnor U29574 (N_29574,N_28015,N_28176);
nor U29575 (N_29575,N_27115,N_27302);
and U29576 (N_29576,N_27889,N_27212);
nor U29577 (N_29577,N_27981,N_28434);
and U29578 (N_29578,N_27013,N_27797);
or U29579 (N_29579,N_27127,N_27710);
xnor U29580 (N_29580,N_27980,N_28332);
and U29581 (N_29581,N_28062,N_28269);
xnor U29582 (N_29582,N_28288,N_27605);
xor U29583 (N_29583,N_28348,N_27729);
nand U29584 (N_29584,N_28435,N_27397);
or U29585 (N_29585,N_27205,N_27085);
or U29586 (N_29586,N_28014,N_27673);
xor U29587 (N_29587,N_27995,N_27728);
and U29588 (N_29588,N_27573,N_27374);
and U29589 (N_29589,N_27328,N_28010);
nand U29590 (N_29590,N_28202,N_28482);
or U29591 (N_29591,N_27009,N_27376);
xor U29592 (N_29592,N_28283,N_27838);
and U29593 (N_29593,N_28383,N_27805);
and U29594 (N_29594,N_28233,N_27924);
nor U29595 (N_29595,N_27163,N_27687);
nand U29596 (N_29596,N_28278,N_27455);
or U29597 (N_29597,N_28063,N_28371);
nor U29598 (N_29598,N_28083,N_27346);
nor U29599 (N_29599,N_28095,N_27334);
and U29600 (N_29600,N_27753,N_27132);
nand U29601 (N_29601,N_27532,N_27144);
nand U29602 (N_29602,N_27148,N_28076);
nor U29603 (N_29603,N_27842,N_27154);
nand U29604 (N_29604,N_27002,N_27379);
nor U29605 (N_29605,N_27644,N_28351);
nand U29606 (N_29606,N_27621,N_27953);
and U29607 (N_29607,N_28345,N_28210);
and U29608 (N_29608,N_27875,N_28117);
nor U29609 (N_29609,N_27027,N_27452);
nor U29610 (N_29610,N_28488,N_28013);
or U29611 (N_29611,N_27944,N_27481);
nand U29612 (N_29612,N_27082,N_27404);
and U29613 (N_29613,N_28068,N_27453);
and U29614 (N_29614,N_28492,N_28081);
or U29615 (N_29615,N_27751,N_27206);
or U29616 (N_29616,N_27148,N_27853);
nor U29617 (N_29617,N_27311,N_28359);
xnor U29618 (N_29618,N_28188,N_27113);
nor U29619 (N_29619,N_27403,N_28116);
xnor U29620 (N_29620,N_28476,N_28445);
and U29621 (N_29621,N_28142,N_27061);
xor U29622 (N_29622,N_27040,N_28055);
nand U29623 (N_29623,N_27918,N_28379);
nand U29624 (N_29624,N_27130,N_27175);
or U29625 (N_29625,N_27728,N_27010);
and U29626 (N_29626,N_28361,N_27730);
or U29627 (N_29627,N_27926,N_28402);
and U29628 (N_29628,N_28297,N_27389);
or U29629 (N_29629,N_28331,N_28479);
xor U29630 (N_29630,N_28135,N_28278);
and U29631 (N_29631,N_27930,N_27690);
and U29632 (N_29632,N_28261,N_27678);
nor U29633 (N_29633,N_27645,N_27689);
nor U29634 (N_29634,N_27295,N_27735);
nand U29635 (N_29635,N_27641,N_28002);
and U29636 (N_29636,N_27758,N_27567);
nor U29637 (N_29637,N_27380,N_28427);
xor U29638 (N_29638,N_27785,N_28403);
nand U29639 (N_29639,N_28318,N_27452);
nor U29640 (N_29640,N_27462,N_27132);
and U29641 (N_29641,N_28051,N_27000);
nand U29642 (N_29642,N_27669,N_28293);
xnor U29643 (N_29643,N_28320,N_28407);
and U29644 (N_29644,N_28086,N_27325);
or U29645 (N_29645,N_28419,N_27010);
nand U29646 (N_29646,N_28494,N_27044);
xnor U29647 (N_29647,N_28047,N_27981);
or U29648 (N_29648,N_27312,N_27666);
and U29649 (N_29649,N_28353,N_27526);
or U29650 (N_29650,N_27002,N_27934);
nor U29651 (N_29651,N_28139,N_27957);
and U29652 (N_29652,N_27514,N_27428);
and U29653 (N_29653,N_27561,N_28234);
and U29654 (N_29654,N_27185,N_27231);
or U29655 (N_29655,N_27749,N_27649);
nand U29656 (N_29656,N_28397,N_28095);
and U29657 (N_29657,N_28144,N_27011);
and U29658 (N_29658,N_27434,N_28289);
and U29659 (N_29659,N_27384,N_27372);
nor U29660 (N_29660,N_27162,N_28261);
or U29661 (N_29661,N_27139,N_27202);
or U29662 (N_29662,N_27362,N_27711);
nor U29663 (N_29663,N_27321,N_27037);
and U29664 (N_29664,N_27822,N_27817);
and U29665 (N_29665,N_28343,N_28287);
nand U29666 (N_29666,N_27034,N_27897);
or U29667 (N_29667,N_28478,N_28139);
xnor U29668 (N_29668,N_28263,N_27695);
and U29669 (N_29669,N_27552,N_27290);
xor U29670 (N_29670,N_27187,N_27564);
or U29671 (N_29671,N_28490,N_27521);
or U29672 (N_29672,N_28366,N_27622);
nand U29673 (N_29673,N_27192,N_28019);
nor U29674 (N_29674,N_27262,N_27130);
nor U29675 (N_29675,N_27052,N_27147);
and U29676 (N_29676,N_27594,N_27469);
xor U29677 (N_29677,N_28154,N_27470);
or U29678 (N_29678,N_28219,N_27489);
nand U29679 (N_29679,N_27867,N_27090);
and U29680 (N_29680,N_27676,N_27832);
and U29681 (N_29681,N_27627,N_28453);
nor U29682 (N_29682,N_27113,N_27961);
and U29683 (N_29683,N_28071,N_27031);
xnor U29684 (N_29684,N_28070,N_27380);
and U29685 (N_29685,N_27776,N_27763);
xor U29686 (N_29686,N_28209,N_27361);
and U29687 (N_29687,N_28361,N_27572);
and U29688 (N_29688,N_27880,N_27928);
or U29689 (N_29689,N_28363,N_27135);
and U29690 (N_29690,N_27700,N_27790);
or U29691 (N_29691,N_28484,N_27176);
xnor U29692 (N_29692,N_28230,N_27414);
nor U29693 (N_29693,N_28285,N_27465);
or U29694 (N_29694,N_28389,N_27999);
nand U29695 (N_29695,N_27735,N_28022);
or U29696 (N_29696,N_28261,N_28302);
xor U29697 (N_29697,N_28350,N_27519);
xor U29698 (N_29698,N_27032,N_28253);
nor U29699 (N_29699,N_27285,N_27010);
or U29700 (N_29700,N_27156,N_28011);
and U29701 (N_29701,N_27036,N_27091);
xnor U29702 (N_29702,N_28190,N_27492);
and U29703 (N_29703,N_27846,N_27303);
xnor U29704 (N_29704,N_28074,N_27475);
xnor U29705 (N_29705,N_28172,N_27398);
nand U29706 (N_29706,N_28450,N_27949);
xnor U29707 (N_29707,N_27814,N_27086);
xnor U29708 (N_29708,N_27900,N_27827);
xor U29709 (N_29709,N_28454,N_27812);
nand U29710 (N_29710,N_28364,N_27360);
nand U29711 (N_29711,N_28424,N_28257);
nand U29712 (N_29712,N_27665,N_27146);
nor U29713 (N_29713,N_27295,N_27604);
xnor U29714 (N_29714,N_27239,N_28196);
nor U29715 (N_29715,N_27861,N_27606);
nand U29716 (N_29716,N_27243,N_28177);
and U29717 (N_29717,N_28428,N_27864);
nand U29718 (N_29718,N_27274,N_28196);
and U29719 (N_29719,N_28085,N_28086);
nand U29720 (N_29720,N_27695,N_27424);
nand U29721 (N_29721,N_28134,N_28203);
nand U29722 (N_29722,N_27612,N_28041);
and U29723 (N_29723,N_27979,N_27689);
nor U29724 (N_29724,N_28008,N_27025);
xnor U29725 (N_29725,N_28495,N_27695);
and U29726 (N_29726,N_27574,N_27782);
or U29727 (N_29727,N_27460,N_27638);
or U29728 (N_29728,N_28419,N_27022);
nand U29729 (N_29729,N_27053,N_27976);
and U29730 (N_29730,N_27142,N_27695);
and U29731 (N_29731,N_27400,N_28365);
and U29732 (N_29732,N_28064,N_28102);
nor U29733 (N_29733,N_27790,N_27075);
and U29734 (N_29734,N_28131,N_28310);
or U29735 (N_29735,N_28141,N_27409);
nor U29736 (N_29736,N_28113,N_28347);
xor U29737 (N_29737,N_27468,N_27503);
and U29738 (N_29738,N_27079,N_27122);
xor U29739 (N_29739,N_27800,N_27818);
nor U29740 (N_29740,N_27227,N_28441);
xor U29741 (N_29741,N_28160,N_27746);
nand U29742 (N_29742,N_28300,N_28401);
nand U29743 (N_29743,N_27279,N_28180);
and U29744 (N_29744,N_27666,N_27199);
nor U29745 (N_29745,N_27474,N_27780);
nor U29746 (N_29746,N_27270,N_27189);
and U29747 (N_29747,N_27612,N_27111);
or U29748 (N_29748,N_27248,N_27267);
xor U29749 (N_29749,N_28340,N_27814);
xor U29750 (N_29750,N_27308,N_28182);
or U29751 (N_29751,N_28457,N_27804);
nand U29752 (N_29752,N_27840,N_27638);
nand U29753 (N_29753,N_27912,N_28005);
and U29754 (N_29754,N_27989,N_27070);
nor U29755 (N_29755,N_27550,N_28333);
nand U29756 (N_29756,N_28250,N_27561);
and U29757 (N_29757,N_28112,N_27610);
and U29758 (N_29758,N_27525,N_28389);
nand U29759 (N_29759,N_27827,N_27865);
and U29760 (N_29760,N_27896,N_28324);
xnor U29761 (N_29761,N_27158,N_27129);
nand U29762 (N_29762,N_28237,N_27430);
or U29763 (N_29763,N_27100,N_27020);
nor U29764 (N_29764,N_27266,N_28009);
or U29765 (N_29765,N_27877,N_28146);
nor U29766 (N_29766,N_28049,N_27132);
or U29767 (N_29767,N_27167,N_27964);
or U29768 (N_29768,N_27675,N_27762);
xnor U29769 (N_29769,N_27932,N_28211);
nor U29770 (N_29770,N_28167,N_28124);
or U29771 (N_29771,N_28361,N_28369);
nor U29772 (N_29772,N_27214,N_27753);
nand U29773 (N_29773,N_27433,N_27339);
or U29774 (N_29774,N_28080,N_27655);
and U29775 (N_29775,N_28340,N_28428);
nand U29776 (N_29776,N_28411,N_27815);
or U29777 (N_29777,N_27953,N_28071);
xor U29778 (N_29778,N_27735,N_27122);
or U29779 (N_29779,N_27622,N_27441);
nand U29780 (N_29780,N_27968,N_28479);
or U29781 (N_29781,N_28070,N_27880);
nor U29782 (N_29782,N_27610,N_28129);
or U29783 (N_29783,N_28245,N_27247);
xor U29784 (N_29784,N_28102,N_28447);
xor U29785 (N_29785,N_27496,N_27058);
nor U29786 (N_29786,N_27784,N_28153);
and U29787 (N_29787,N_27021,N_28119);
and U29788 (N_29788,N_27878,N_27244);
xnor U29789 (N_29789,N_28376,N_27230);
nor U29790 (N_29790,N_28440,N_27415);
nand U29791 (N_29791,N_27721,N_28462);
or U29792 (N_29792,N_27863,N_27203);
nor U29793 (N_29793,N_28118,N_27414);
nand U29794 (N_29794,N_28251,N_28250);
and U29795 (N_29795,N_27211,N_27248);
xor U29796 (N_29796,N_28219,N_27910);
and U29797 (N_29797,N_28405,N_27125);
nand U29798 (N_29798,N_27345,N_27557);
nand U29799 (N_29799,N_28454,N_28431);
nand U29800 (N_29800,N_28375,N_27226);
xnor U29801 (N_29801,N_28170,N_27971);
nor U29802 (N_29802,N_27554,N_28270);
and U29803 (N_29803,N_28106,N_27568);
nand U29804 (N_29804,N_27816,N_27373);
nand U29805 (N_29805,N_27476,N_27737);
nor U29806 (N_29806,N_28303,N_27135);
and U29807 (N_29807,N_27938,N_27157);
and U29808 (N_29808,N_28334,N_27661);
xor U29809 (N_29809,N_27668,N_28120);
xnor U29810 (N_29810,N_28150,N_27151);
nor U29811 (N_29811,N_27878,N_27715);
or U29812 (N_29812,N_27095,N_27270);
nor U29813 (N_29813,N_27645,N_28479);
nand U29814 (N_29814,N_27136,N_27656);
xnor U29815 (N_29815,N_27563,N_27036);
or U29816 (N_29816,N_27656,N_27119);
nor U29817 (N_29817,N_27553,N_28146);
and U29818 (N_29818,N_27149,N_28317);
or U29819 (N_29819,N_27407,N_27854);
nand U29820 (N_29820,N_27643,N_27243);
nor U29821 (N_29821,N_27304,N_28377);
and U29822 (N_29822,N_28122,N_27155);
nor U29823 (N_29823,N_28332,N_27529);
or U29824 (N_29824,N_27077,N_27357);
or U29825 (N_29825,N_27776,N_27879);
or U29826 (N_29826,N_27050,N_28022);
and U29827 (N_29827,N_27958,N_27739);
and U29828 (N_29828,N_28134,N_27037);
or U29829 (N_29829,N_27366,N_27887);
xor U29830 (N_29830,N_27431,N_27686);
nor U29831 (N_29831,N_27672,N_28397);
xnor U29832 (N_29832,N_27570,N_27437);
nand U29833 (N_29833,N_28339,N_27116);
and U29834 (N_29834,N_28439,N_27435);
nor U29835 (N_29835,N_28292,N_28458);
or U29836 (N_29836,N_27478,N_28326);
nand U29837 (N_29837,N_27454,N_27957);
nand U29838 (N_29838,N_27165,N_27242);
xnor U29839 (N_29839,N_28291,N_27076);
xor U29840 (N_29840,N_28282,N_28027);
or U29841 (N_29841,N_28303,N_27547);
and U29842 (N_29842,N_27337,N_27612);
nor U29843 (N_29843,N_28429,N_27551);
nand U29844 (N_29844,N_27678,N_27741);
nand U29845 (N_29845,N_28141,N_27629);
nor U29846 (N_29846,N_27591,N_27487);
and U29847 (N_29847,N_27009,N_28398);
and U29848 (N_29848,N_27079,N_27306);
nor U29849 (N_29849,N_27360,N_27055);
or U29850 (N_29850,N_27172,N_27001);
or U29851 (N_29851,N_27917,N_27660);
xor U29852 (N_29852,N_27788,N_28310);
nand U29853 (N_29853,N_27665,N_27053);
nand U29854 (N_29854,N_27745,N_28047);
nor U29855 (N_29855,N_28168,N_27205);
nor U29856 (N_29856,N_27953,N_28214);
nand U29857 (N_29857,N_27844,N_27858);
and U29858 (N_29858,N_28419,N_27750);
nand U29859 (N_29859,N_28068,N_27025);
or U29860 (N_29860,N_27547,N_27362);
nor U29861 (N_29861,N_27362,N_28485);
or U29862 (N_29862,N_27676,N_27112);
or U29863 (N_29863,N_28489,N_27082);
nor U29864 (N_29864,N_28122,N_27029);
or U29865 (N_29865,N_27335,N_28360);
or U29866 (N_29866,N_27308,N_27316);
nor U29867 (N_29867,N_27743,N_28073);
and U29868 (N_29868,N_28306,N_27874);
and U29869 (N_29869,N_27802,N_28342);
nand U29870 (N_29870,N_27818,N_28200);
nor U29871 (N_29871,N_27555,N_28161);
xor U29872 (N_29872,N_27705,N_28307);
or U29873 (N_29873,N_28220,N_28007);
and U29874 (N_29874,N_27094,N_27793);
nor U29875 (N_29875,N_27030,N_27854);
nand U29876 (N_29876,N_27323,N_28212);
and U29877 (N_29877,N_28249,N_27578);
xor U29878 (N_29878,N_28480,N_27922);
and U29879 (N_29879,N_28253,N_28054);
xor U29880 (N_29880,N_27870,N_27420);
xnor U29881 (N_29881,N_28023,N_27142);
nand U29882 (N_29882,N_27345,N_28409);
or U29883 (N_29883,N_28369,N_27908);
nor U29884 (N_29884,N_27773,N_27606);
and U29885 (N_29885,N_28003,N_27344);
nor U29886 (N_29886,N_27914,N_28145);
nor U29887 (N_29887,N_28356,N_27723);
xor U29888 (N_29888,N_28389,N_28393);
xnor U29889 (N_29889,N_27526,N_28292);
and U29890 (N_29890,N_28496,N_27907);
nand U29891 (N_29891,N_28126,N_28399);
and U29892 (N_29892,N_27273,N_28353);
and U29893 (N_29893,N_27366,N_27915);
nor U29894 (N_29894,N_28358,N_27646);
or U29895 (N_29895,N_28113,N_27189);
xnor U29896 (N_29896,N_27792,N_27747);
nor U29897 (N_29897,N_27351,N_27288);
xor U29898 (N_29898,N_27909,N_28125);
nand U29899 (N_29899,N_28438,N_27644);
nand U29900 (N_29900,N_27294,N_27020);
or U29901 (N_29901,N_28032,N_28288);
and U29902 (N_29902,N_27659,N_27197);
or U29903 (N_29903,N_27011,N_28377);
nor U29904 (N_29904,N_28411,N_27693);
nor U29905 (N_29905,N_27152,N_28269);
and U29906 (N_29906,N_28148,N_27246);
or U29907 (N_29907,N_27655,N_28352);
nand U29908 (N_29908,N_28307,N_27856);
and U29909 (N_29909,N_27068,N_27752);
nor U29910 (N_29910,N_27126,N_28093);
nor U29911 (N_29911,N_28491,N_27626);
and U29912 (N_29912,N_28345,N_27646);
nor U29913 (N_29913,N_27661,N_28266);
nand U29914 (N_29914,N_27040,N_27641);
nand U29915 (N_29915,N_27606,N_27578);
nor U29916 (N_29916,N_27948,N_27179);
or U29917 (N_29917,N_27583,N_27800);
xor U29918 (N_29918,N_28273,N_27524);
nand U29919 (N_29919,N_28196,N_28105);
or U29920 (N_29920,N_27427,N_27355);
or U29921 (N_29921,N_27376,N_27591);
and U29922 (N_29922,N_27303,N_27121);
nand U29923 (N_29923,N_27477,N_28437);
and U29924 (N_29924,N_27686,N_27858);
or U29925 (N_29925,N_28409,N_27221);
xnor U29926 (N_29926,N_28381,N_27417);
xnor U29927 (N_29927,N_27247,N_27273);
and U29928 (N_29928,N_27716,N_27587);
or U29929 (N_29929,N_27541,N_28222);
or U29930 (N_29930,N_28262,N_27927);
and U29931 (N_29931,N_27270,N_28005);
xnor U29932 (N_29932,N_27680,N_28389);
nand U29933 (N_29933,N_27665,N_27737);
nor U29934 (N_29934,N_28399,N_27649);
nand U29935 (N_29935,N_27320,N_27558);
nand U29936 (N_29936,N_28314,N_27356);
nand U29937 (N_29937,N_27136,N_28413);
or U29938 (N_29938,N_27794,N_27831);
nor U29939 (N_29939,N_28243,N_27076);
nor U29940 (N_29940,N_27246,N_27504);
and U29941 (N_29941,N_28009,N_28330);
or U29942 (N_29942,N_27275,N_27321);
or U29943 (N_29943,N_28177,N_27237);
and U29944 (N_29944,N_28310,N_27466);
xor U29945 (N_29945,N_28246,N_27223);
nor U29946 (N_29946,N_28194,N_27963);
xor U29947 (N_29947,N_27612,N_28334);
nand U29948 (N_29948,N_27429,N_28116);
and U29949 (N_29949,N_27905,N_27343);
nor U29950 (N_29950,N_28229,N_28098);
or U29951 (N_29951,N_28160,N_27446);
xnor U29952 (N_29952,N_27435,N_27607);
or U29953 (N_29953,N_28209,N_27677);
or U29954 (N_29954,N_27422,N_27830);
or U29955 (N_29955,N_28234,N_28071);
xor U29956 (N_29956,N_27581,N_27467);
or U29957 (N_29957,N_28356,N_27893);
and U29958 (N_29958,N_27814,N_28479);
or U29959 (N_29959,N_27769,N_27668);
or U29960 (N_29960,N_28426,N_27092);
and U29961 (N_29961,N_28400,N_27760);
xor U29962 (N_29962,N_28178,N_28417);
and U29963 (N_29963,N_27593,N_28181);
or U29964 (N_29964,N_27140,N_27755);
or U29965 (N_29965,N_27198,N_27333);
nand U29966 (N_29966,N_28431,N_27146);
nor U29967 (N_29967,N_28440,N_27947);
nor U29968 (N_29968,N_28011,N_27947);
nand U29969 (N_29969,N_27373,N_27326);
nand U29970 (N_29970,N_27828,N_28305);
nor U29971 (N_29971,N_27607,N_27634);
xor U29972 (N_29972,N_27826,N_27499);
and U29973 (N_29973,N_28271,N_27098);
xnor U29974 (N_29974,N_27843,N_28198);
nand U29975 (N_29975,N_27614,N_28464);
and U29976 (N_29976,N_28176,N_28234);
or U29977 (N_29977,N_27835,N_27513);
xnor U29978 (N_29978,N_27750,N_28195);
nand U29979 (N_29979,N_28363,N_28359);
nand U29980 (N_29980,N_27551,N_28407);
or U29981 (N_29981,N_27823,N_28136);
or U29982 (N_29982,N_28432,N_27473);
or U29983 (N_29983,N_28220,N_27734);
nand U29984 (N_29984,N_28442,N_28355);
nand U29985 (N_29985,N_28276,N_28443);
nor U29986 (N_29986,N_27452,N_27781);
or U29987 (N_29987,N_27999,N_28239);
and U29988 (N_29988,N_27243,N_28379);
nor U29989 (N_29989,N_28094,N_27448);
and U29990 (N_29990,N_27018,N_27186);
xnor U29991 (N_29991,N_27146,N_28055);
nand U29992 (N_29992,N_28384,N_28269);
or U29993 (N_29993,N_27221,N_28190);
and U29994 (N_29994,N_27570,N_27701);
and U29995 (N_29995,N_27276,N_27781);
or U29996 (N_29996,N_27246,N_27708);
and U29997 (N_29997,N_27900,N_28006);
xnor U29998 (N_29998,N_27832,N_28219);
or U29999 (N_29999,N_27011,N_28138);
nand UO_0 (O_0,N_29753,N_28734);
nor UO_1 (O_1,N_29050,N_28582);
or UO_2 (O_2,N_29589,N_29970);
nor UO_3 (O_3,N_28685,N_28592);
xor UO_4 (O_4,N_29631,N_29131);
and UO_5 (O_5,N_29088,N_28828);
nor UO_6 (O_6,N_28961,N_28895);
xnor UO_7 (O_7,N_29504,N_28645);
and UO_8 (O_8,N_29007,N_29355);
or UO_9 (O_9,N_28767,N_29892);
xor UO_10 (O_10,N_29690,N_29220);
nor UO_11 (O_11,N_29662,N_29773);
and UO_12 (O_12,N_29678,N_29240);
nand UO_13 (O_13,N_28712,N_29483);
nor UO_14 (O_14,N_29744,N_29223);
nor UO_15 (O_15,N_28525,N_28687);
or UO_16 (O_16,N_28669,N_29335);
nor UO_17 (O_17,N_29058,N_28880);
xnor UO_18 (O_18,N_28771,N_28719);
and UO_19 (O_19,N_28954,N_29983);
or UO_20 (O_20,N_28979,N_29768);
or UO_21 (O_21,N_29352,N_29913);
nor UO_22 (O_22,N_29497,N_28883);
and UO_23 (O_23,N_28824,N_28947);
nand UO_24 (O_24,N_29023,N_29495);
nor UO_25 (O_25,N_29942,N_28623);
nor UO_26 (O_26,N_29717,N_28703);
and UO_27 (O_27,N_29969,N_28556);
or UO_28 (O_28,N_28717,N_29436);
xor UO_29 (O_29,N_28584,N_28742);
xor UO_30 (O_30,N_28833,N_29967);
xnor UO_31 (O_31,N_29470,N_28773);
and UO_32 (O_32,N_28672,N_28951);
and UO_33 (O_33,N_29109,N_29803);
or UO_34 (O_34,N_29151,N_29257);
and UO_35 (O_35,N_29968,N_29784);
or UO_36 (O_36,N_28626,N_28689);
and UO_37 (O_37,N_28643,N_29127);
and UO_38 (O_38,N_29858,N_29905);
nor UO_39 (O_39,N_28813,N_29111);
nand UO_40 (O_40,N_29906,N_28573);
or UO_41 (O_41,N_28809,N_29519);
nand UO_42 (O_42,N_29345,N_29565);
or UO_43 (O_43,N_29965,N_29617);
and UO_44 (O_44,N_29539,N_29532);
nor UO_45 (O_45,N_29751,N_28612);
and UO_46 (O_46,N_28735,N_28905);
or UO_47 (O_47,N_29912,N_29908);
nand UO_48 (O_48,N_29601,N_29988);
xor UO_49 (O_49,N_28991,N_29999);
or UO_50 (O_50,N_28786,N_28968);
or UO_51 (O_51,N_29471,N_28577);
nor UO_52 (O_52,N_28743,N_29747);
or UO_53 (O_53,N_28962,N_29191);
nand UO_54 (O_54,N_29450,N_28714);
and UO_55 (O_55,N_29206,N_28635);
and UO_56 (O_56,N_29701,N_28907);
or UO_57 (O_57,N_29693,N_29719);
xnor UO_58 (O_58,N_29552,N_28845);
or UO_59 (O_59,N_28692,N_28914);
and UO_60 (O_60,N_29344,N_28513);
nand UO_61 (O_61,N_28535,N_28680);
or UO_62 (O_62,N_29775,N_29266);
and UO_63 (O_63,N_29762,N_28705);
xnor UO_64 (O_64,N_29243,N_29273);
nor UO_65 (O_65,N_28957,N_28909);
or UO_66 (O_66,N_29125,N_28620);
and UO_67 (O_67,N_29432,N_29829);
or UO_68 (O_68,N_29417,N_29840);
nor UO_69 (O_69,N_29544,N_29196);
or UO_70 (O_70,N_28554,N_29161);
and UO_71 (O_71,N_29216,N_29666);
nor UO_72 (O_72,N_29576,N_29478);
nand UO_73 (O_73,N_29425,N_29353);
nor UO_74 (O_74,N_29779,N_29697);
nor UO_75 (O_75,N_29136,N_29440);
and UO_76 (O_76,N_29072,N_29336);
or UO_77 (O_77,N_29713,N_29537);
or UO_78 (O_78,N_28980,N_28775);
xor UO_79 (O_79,N_29807,N_29868);
nor UO_80 (O_80,N_29742,N_29357);
and UO_81 (O_81,N_28528,N_28625);
and UO_82 (O_82,N_28811,N_29252);
nand UO_83 (O_83,N_29839,N_29083);
or UO_84 (O_84,N_28572,N_29499);
and UO_85 (O_85,N_29330,N_29994);
xor UO_86 (O_86,N_29210,N_29361);
nor UO_87 (O_87,N_29479,N_29397);
or UO_88 (O_88,N_28978,N_29493);
nand UO_89 (O_89,N_28722,N_29384);
xnor UO_90 (O_90,N_29961,N_28842);
and UO_91 (O_91,N_28658,N_28996);
or UO_92 (O_92,N_29780,N_29932);
and UO_93 (O_93,N_29267,N_28605);
or UO_94 (O_94,N_29838,N_29806);
xor UO_95 (O_95,N_28870,N_28855);
and UO_96 (O_96,N_28606,N_28506);
xnor UO_97 (O_97,N_29523,N_29649);
or UO_98 (O_98,N_28732,N_29958);
and UO_99 (O_99,N_29230,N_29006);
nand UO_100 (O_100,N_28729,N_28519);
and UO_101 (O_101,N_29319,N_28631);
or UO_102 (O_102,N_28945,N_29706);
nor UO_103 (O_103,N_28936,N_29106);
and UO_104 (O_104,N_29886,N_29563);
nor UO_105 (O_105,N_29094,N_29178);
or UO_106 (O_106,N_28790,N_29653);
nor UO_107 (O_107,N_29192,N_28723);
nor UO_108 (O_108,N_29110,N_28608);
or UO_109 (O_109,N_28686,N_29016);
nand UO_110 (O_110,N_29062,N_29317);
and UO_111 (O_111,N_29102,N_29786);
and UO_112 (O_112,N_29882,N_28699);
nor UO_113 (O_113,N_28896,N_29696);
or UO_114 (O_114,N_28718,N_29323);
xnor UO_115 (O_115,N_29571,N_29239);
nor UO_116 (O_116,N_29399,N_28733);
nor UO_117 (O_117,N_29503,N_28863);
nor UO_118 (O_118,N_29846,N_28949);
nand UO_119 (O_119,N_28921,N_28799);
nand UO_120 (O_120,N_28507,N_29769);
nor UO_121 (O_121,N_29652,N_28546);
nand UO_122 (O_122,N_28776,N_29457);
nand UO_123 (O_123,N_29376,N_28761);
nand UO_124 (O_124,N_29669,N_29554);
xor UO_125 (O_125,N_29512,N_28558);
nor UO_126 (O_126,N_29730,N_29893);
or UO_127 (O_127,N_28762,N_29297);
nor UO_128 (O_128,N_29797,N_29040);
or UO_129 (O_129,N_28831,N_28797);
nand UO_130 (O_130,N_29671,N_28868);
xnor UO_131 (O_131,N_28964,N_28690);
xnor UO_132 (O_132,N_28515,N_29001);
or UO_133 (O_133,N_29670,N_29386);
nand UO_134 (O_134,N_29320,N_29644);
xor UO_135 (O_135,N_29261,N_29657);
or UO_136 (O_136,N_29279,N_29326);
nand UO_137 (O_137,N_29205,N_29595);
and UO_138 (O_138,N_29656,N_29809);
or UO_139 (O_139,N_29877,N_28518);
or UO_140 (O_140,N_28826,N_29931);
xor UO_141 (O_141,N_28886,N_29569);
nor UO_142 (O_142,N_28911,N_29603);
nor UO_143 (O_143,N_29574,N_29314);
and UO_144 (O_144,N_28580,N_28505);
nor UO_145 (O_145,N_29650,N_29978);
xor UO_146 (O_146,N_29280,N_28562);
or UO_147 (O_147,N_29150,N_29464);
and UO_148 (O_148,N_29985,N_29406);
xor UO_149 (O_149,N_29518,N_29513);
or UO_150 (O_150,N_28578,N_29638);
nor UO_151 (O_151,N_28759,N_29259);
xor UO_152 (O_152,N_29146,N_29919);
nor UO_153 (O_153,N_29682,N_29374);
nor UO_154 (O_154,N_29822,N_28881);
nor UO_155 (O_155,N_29881,N_28902);
and UO_156 (O_156,N_29204,N_29447);
nand UO_157 (O_157,N_28610,N_28878);
or UO_158 (O_158,N_29920,N_29458);
nand UO_159 (O_159,N_28866,N_28641);
xor UO_160 (O_160,N_28851,N_28698);
nand UO_161 (O_161,N_29392,N_29300);
or UO_162 (O_162,N_29089,N_29416);
nor UO_163 (O_163,N_29026,N_29745);
and UO_164 (O_164,N_29788,N_28696);
and UO_165 (O_165,N_29590,N_29667);
xnor UO_166 (O_166,N_29575,N_29098);
nand UO_167 (O_167,N_29844,N_29443);
xor UO_168 (O_168,N_28653,N_29366);
or UO_169 (O_169,N_28874,N_29270);
nand UO_170 (O_170,N_29129,N_29229);
xnor UO_171 (O_171,N_29872,N_28854);
or UO_172 (O_172,N_28816,N_29910);
or UO_173 (O_173,N_29039,N_29343);
nor UO_174 (O_174,N_28670,N_29845);
or UO_175 (O_175,N_29453,N_29289);
xnor UO_176 (O_176,N_28983,N_29375);
nor UO_177 (O_177,N_29095,N_29939);
nor UO_178 (O_178,N_29276,N_29249);
xor UO_179 (O_179,N_28511,N_29372);
or UO_180 (O_180,N_29287,N_29430);
xor UO_181 (O_181,N_28912,N_28649);
and UO_182 (O_182,N_28810,N_29414);
nand UO_183 (O_183,N_28887,N_29577);
or UO_184 (O_184,N_28925,N_28557);
xnor UO_185 (O_185,N_29799,N_29284);
nand UO_186 (O_186,N_29277,N_28959);
nor UO_187 (O_187,N_28544,N_29472);
nand UO_188 (O_188,N_29302,N_29348);
nor UO_189 (O_189,N_29263,N_28716);
or UO_190 (O_190,N_28527,N_29468);
and UO_191 (O_191,N_28531,N_29195);
and UO_192 (O_192,N_29560,N_28995);
or UO_193 (O_193,N_28969,N_29048);
nand UO_194 (O_194,N_29708,N_28640);
xor UO_195 (O_195,N_29077,N_29727);
nand UO_196 (O_196,N_29226,N_28622);
or UO_197 (O_197,N_29438,N_29043);
xor UO_198 (O_198,N_28656,N_29180);
and UO_199 (O_199,N_28588,N_29736);
xnor UO_200 (O_200,N_28609,N_29188);
nor UO_201 (O_201,N_28987,N_29976);
nor UO_202 (O_202,N_29757,N_29303);
xor UO_203 (O_203,N_28568,N_29804);
nand UO_204 (O_204,N_29524,N_29897);
or UO_205 (O_205,N_29288,N_29632);
and UO_206 (O_206,N_28857,N_29911);
nor UO_207 (O_207,N_29278,N_28632);
xnor UO_208 (O_208,N_29238,N_29930);
or UO_209 (O_209,N_29256,N_29028);
xor UO_210 (O_210,N_29242,N_28940);
xnor UO_211 (O_211,N_29347,N_28836);
nand UO_212 (O_212,N_29707,N_29814);
and UO_213 (O_213,N_29036,N_28832);
xnor UO_214 (O_214,N_29936,N_29076);
or UO_215 (O_215,N_29553,N_29860);
nor UO_216 (O_216,N_28749,N_28893);
xor UO_217 (O_217,N_29274,N_29579);
nand UO_218 (O_218,N_29451,N_29620);
and UO_219 (O_219,N_29469,N_29581);
and UO_220 (O_220,N_28785,N_28700);
or UO_221 (O_221,N_29199,N_28872);
and UO_222 (O_222,N_29455,N_29415);
nand UO_223 (O_223,N_28958,N_29624);
or UO_224 (O_224,N_28756,N_29668);
or UO_225 (O_225,N_29090,N_29369);
nor UO_226 (O_226,N_29140,N_28710);
nand UO_227 (O_227,N_28667,N_29012);
or UO_228 (O_228,N_29827,N_29435);
nor UO_229 (O_229,N_29639,N_29431);
nand UO_230 (O_230,N_29311,N_28955);
xor UO_231 (O_231,N_29408,N_28989);
or UO_232 (O_232,N_28726,N_29365);
or UO_233 (O_233,N_29253,N_29625);
and UO_234 (O_234,N_29496,N_29895);
xor UO_235 (O_235,N_29128,N_28611);
nand UO_236 (O_236,N_29709,N_29733);
or UO_237 (O_237,N_28618,N_29449);
nand UO_238 (O_238,N_29534,N_28988);
nor UO_239 (O_239,N_29789,N_28655);
nor UO_240 (O_240,N_29360,N_28861);
and UO_241 (O_241,N_29658,N_28839);
or UO_242 (O_242,N_28850,N_29025);
and UO_243 (O_243,N_28569,N_29413);
xnor UO_244 (O_244,N_29771,N_29465);
nand UO_245 (O_245,N_28574,N_29694);
and UO_246 (O_246,N_29852,N_29531);
xor UO_247 (O_247,N_29866,N_29142);
or UO_248 (O_248,N_28899,N_29429);
or UO_249 (O_249,N_28589,N_29074);
nand UO_250 (O_250,N_28637,N_28848);
xnor UO_251 (O_251,N_29339,N_29830);
or UO_252 (O_252,N_29993,N_29189);
and UO_253 (O_253,N_28924,N_29086);
nor UO_254 (O_254,N_29227,N_29373);
nor UO_255 (O_255,N_28966,N_29057);
or UO_256 (O_256,N_29865,N_29591);
and UO_257 (O_257,N_29281,N_28688);
and UO_258 (O_258,N_29686,N_28748);
nand UO_259 (O_259,N_29139,N_29712);
and UO_260 (O_260,N_29855,N_29763);
xor UO_261 (O_261,N_29953,N_28744);
and UO_262 (O_262,N_28789,N_29502);
xnor UO_263 (O_263,N_29957,N_28898);
and UO_264 (O_264,N_29309,N_29525);
and UO_265 (O_265,N_29538,N_29507);
or UO_266 (O_266,N_29175,N_29857);
nor UO_267 (O_267,N_29896,N_29987);
xor UO_268 (O_268,N_29182,N_28805);
or UO_269 (O_269,N_29460,N_28849);
xnor UO_270 (O_270,N_29186,N_29116);
nand UO_271 (O_271,N_29456,N_29641);
and UO_272 (O_272,N_29726,N_29214);
nor UO_273 (O_273,N_29124,N_29029);
and UO_274 (O_274,N_29955,N_29015);
nor UO_275 (O_275,N_29848,N_29391);
nand UO_276 (O_276,N_29740,N_29437);
xor UO_277 (O_277,N_29433,N_29246);
and UO_278 (O_278,N_28906,N_28662);
or UO_279 (O_279,N_29032,N_29647);
nand UO_280 (O_280,N_29236,N_29648);
xor UO_281 (O_281,N_28939,N_28757);
nor UO_282 (O_282,N_29067,N_29557);
xnor UO_283 (O_283,N_29020,N_28946);
or UO_284 (O_284,N_29593,N_29698);
or UO_285 (O_285,N_28539,N_28815);
nor UO_286 (O_286,N_28512,N_29586);
nand UO_287 (O_287,N_29514,N_29021);
and UO_288 (O_288,N_29138,N_29980);
xor UO_289 (O_289,N_29444,N_29732);
xnor UO_290 (O_290,N_28534,N_29903);
nand UO_291 (O_291,N_29202,N_29511);
or UO_292 (O_292,N_29526,N_29411);
nor UO_293 (O_293,N_29439,N_28600);
or UO_294 (O_294,N_29388,N_29222);
and UO_295 (O_295,N_29307,N_29568);
nand UO_296 (O_296,N_29673,N_29285);
and UO_297 (O_297,N_29609,N_29211);
nand UO_298 (O_298,N_29901,N_28990);
or UO_299 (O_299,N_29722,N_29940);
nor UO_300 (O_300,N_29646,N_28950);
or UO_301 (O_301,N_29914,N_29061);
xor UO_302 (O_302,N_28616,N_28801);
xnor UO_303 (O_303,N_29824,N_28882);
and UO_304 (O_304,N_29370,N_28774);
and UO_305 (O_305,N_29003,N_29615);
or UO_306 (O_306,N_29849,N_29545);
or UO_307 (O_307,N_29183,N_29718);
nor UO_308 (O_308,N_29876,N_29572);
nand UO_309 (O_309,N_28794,N_28751);
and UO_310 (O_310,N_28587,N_28739);
nand UO_311 (O_311,N_28942,N_28792);
nand UO_312 (O_312,N_29772,N_29703);
xor UO_313 (O_313,N_29442,N_28728);
xnor UO_314 (O_314,N_28536,N_29541);
nand UO_315 (O_315,N_29924,N_29152);
or UO_316 (O_316,N_29390,N_29597);
nand UO_317 (O_317,N_29543,N_29165);
xnor UO_318 (O_318,N_29305,N_28843);
and UO_319 (O_319,N_29643,N_28594);
xor UO_320 (O_320,N_29782,N_29163);
or UO_321 (O_321,N_29010,N_29917);
and UO_322 (O_322,N_29559,N_29611);
nor UO_323 (O_323,N_28904,N_29680);
xnor UO_324 (O_324,N_29520,N_29066);
and UO_325 (O_325,N_29405,N_29331);
nor UO_326 (O_326,N_29996,N_28681);
nand UO_327 (O_327,N_28526,N_28927);
xnor UO_328 (O_328,N_29833,N_28884);
nor UO_329 (O_329,N_28533,N_29508);
or UO_330 (O_330,N_29337,N_28754);
nor UO_331 (O_331,N_28553,N_28509);
and UO_332 (O_332,N_28550,N_29594);
or UO_333 (O_333,N_29764,N_29765);
and UO_334 (O_334,N_29810,N_28846);
xor UO_335 (O_335,N_28971,N_29255);
nor UO_336 (O_336,N_29380,N_29823);
xnor UO_337 (O_337,N_28768,N_29837);
or UO_338 (O_338,N_28998,N_29234);
xor UO_339 (O_339,N_28956,N_29721);
and UO_340 (O_340,N_28825,N_28559);
xor UO_341 (O_341,N_29925,N_29723);
and UO_342 (O_342,N_29927,N_29306);
xor UO_343 (O_343,N_29946,N_29466);
and UO_344 (O_344,N_28701,N_29327);
xnor UO_345 (O_345,N_29082,N_28860);
xnor UO_346 (O_346,N_28778,N_28668);
and UO_347 (O_347,N_29777,N_29422);
nor UO_348 (O_348,N_28595,N_29423);
nor UO_349 (O_349,N_29748,N_29861);
and UO_350 (O_350,N_28781,N_29509);
and UO_351 (O_351,N_28674,N_29561);
nor UO_352 (O_352,N_28697,N_29699);
or UO_353 (O_353,N_29123,N_28943);
and UO_354 (O_354,N_29756,N_29659);
or UO_355 (O_355,N_29835,N_29087);
xnor UO_356 (O_356,N_29042,N_29517);
nor UO_357 (O_357,N_28806,N_29785);
nor UO_358 (O_358,N_29071,N_29847);
or UO_359 (O_359,N_29915,N_29655);
or UO_360 (O_360,N_28565,N_28741);
and UO_361 (O_361,N_29622,N_29299);
or UO_362 (O_362,N_29052,N_29613);
and UO_363 (O_363,N_28840,N_29084);
or UO_364 (O_364,N_29971,N_29219);
xor UO_365 (O_365,N_28915,N_28865);
and UO_366 (O_366,N_28615,N_28607);
nand UO_367 (O_367,N_29692,N_28639);
nor UO_368 (O_368,N_29724,N_29900);
xor UO_369 (O_369,N_28522,N_29530);
and UO_370 (O_370,N_29332,N_29168);
xor UO_371 (O_371,N_29929,N_29008);
nor UO_372 (O_372,N_29793,N_28597);
or UO_373 (O_373,N_28901,N_29301);
nand UO_374 (O_374,N_28708,N_29918);
and UO_375 (O_375,N_29290,N_29621);
and UO_376 (O_376,N_29759,N_29612);
xnor UO_377 (O_377,N_28910,N_29367);
nand UO_378 (O_378,N_28928,N_29731);
nand UO_379 (O_379,N_29966,N_29169);
or UO_380 (O_380,N_28837,N_29739);
or UO_381 (O_381,N_28581,N_29051);
and UO_382 (O_382,N_28523,N_29318);
xor UO_383 (O_383,N_28633,N_29688);
nor UO_384 (O_384,N_29185,N_29328);
nor UO_385 (O_385,N_29542,N_29956);
and UO_386 (O_386,N_29033,N_29022);
and UO_387 (O_387,N_29776,N_28934);
nor UO_388 (O_388,N_29122,N_28817);
nor UO_389 (O_389,N_29019,N_29049);
or UO_390 (O_390,N_29529,N_28583);
nand UO_391 (O_391,N_28709,N_29292);
xor UO_392 (O_392,N_29935,N_29774);
nor UO_393 (O_393,N_29158,N_29283);
and UO_394 (O_394,N_28847,N_29676);
and UO_395 (O_395,N_29338,N_29660);
nor UO_396 (O_396,N_29093,N_28879);
and UO_397 (O_397,N_29426,N_29761);
nor UO_398 (O_398,N_28974,N_29684);
and UO_399 (O_399,N_29009,N_29153);
and UO_400 (O_400,N_29884,N_28788);
nand UO_401 (O_401,N_28900,N_29677);
or UO_402 (O_402,N_28579,N_29841);
or UO_403 (O_403,N_29754,N_29528);
and UO_404 (O_404,N_28521,N_29060);
xor UO_405 (O_405,N_29645,N_28844);
or UO_406 (O_406,N_29843,N_28981);
and UO_407 (O_407,N_29928,N_29115);
nand UO_408 (O_408,N_29490,N_29818);
nor UO_409 (O_409,N_29385,N_29176);
nand UO_410 (O_410,N_29623,N_29218);
and UO_411 (O_411,N_29304,N_28693);
and UO_412 (O_412,N_28654,N_28772);
nand UO_413 (O_413,N_29825,N_29610);
and UO_414 (O_414,N_28760,N_28769);
or UO_415 (O_415,N_29923,N_29663);
nor UO_416 (O_416,N_29500,N_28624);
nor UO_417 (O_417,N_29393,N_29959);
and UO_418 (O_418,N_29729,N_29381);
nand UO_419 (O_419,N_28517,N_29636);
nor UO_420 (O_420,N_28869,N_28941);
xnor UO_421 (O_421,N_28691,N_28972);
or UO_422 (O_422,N_28830,N_29056);
nand UO_423 (O_423,N_29629,N_29398);
nor UO_424 (O_424,N_29272,N_29190);
and UO_425 (O_425,N_29446,N_29467);
nand UO_426 (O_426,N_29986,N_28746);
and UO_427 (O_427,N_29329,N_29027);
xor UO_428 (O_428,N_29584,N_28876);
nand UO_429 (O_429,N_29533,N_28571);
nor UO_430 (O_430,N_28711,N_29879);
or UO_431 (O_431,N_29489,N_28619);
nand UO_432 (O_432,N_28814,N_29149);
nand UO_433 (O_433,N_29081,N_29364);
xor UO_434 (O_434,N_29427,N_29002);
and UO_435 (O_435,N_28682,N_28798);
nor UO_436 (O_436,N_29474,N_28764);
and UO_437 (O_437,N_29394,N_29888);
or UO_438 (O_438,N_29949,N_29237);
nand UO_439 (O_439,N_29527,N_29952);
nand UO_440 (O_440,N_29781,N_29035);
or UO_441 (O_441,N_29325,N_29975);
xor UO_442 (O_442,N_29291,N_28986);
nor UO_443 (O_443,N_29606,N_29853);
and UO_444 (O_444,N_28730,N_28783);
nand UO_445 (O_445,N_28665,N_28638);
nor UO_446 (O_446,N_29148,N_29113);
nand UO_447 (O_447,N_28864,N_29296);
nor UO_448 (O_448,N_28777,N_28694);
nor UO_449 (O_449,N_29618,N_28908);
and UO_450 (O_450,N_29247,N_28675);
xnor UO_451 (O_451,N_29434,N_28802);
and UO_452 (O_452,N_29783,N_28540);
nor UO_453 (O_453,N_29535,N_28821);
or UO_454 (O_454,N_29420,N_29598);
nand UO_455 (O_455,N_29550,N_28695);
nor UO_456 (O_456,N_28938,N_29194);
xor UO_457 (O_457,N_29547,N_29979);
nand UO_458 (O_458,N_29995,N_28782);
nor UO_459 (O_459,N_29147,N_29485);
or UO_460 (O_460,N_28551,N_28875);
nand UO_461 (O_461,N_28599,N_28724);
xor UO_462 (O_462,N_28916,N_29602);
xor UO_463 (O_463,N_29548,N_28935);
or UO_464 (O_464,N_29831,N_29120);
xor UO_465 (O_465,N_29691,N_29982);
and UO_466 (O_466,N_28931,N_28500);
xor UO_467 (O_467,N_29501,N_28858);
and UO_468 (O_468,N_28629,N_28560);
nor UO_469 (O_469,N_29600,N_28793);
and UO_470 (O_470,N_29024,N_29642);
or UO_471 (O_471,N_29859,N_29546);
xor UO_472 (O_472,N_29412,N_29794);
nor UO_473 (O_473,N_29564,N_29567);
nor UO_474 (O_474,N_29461,N_29184);
nor UO_475 (O_475,N_29171,N_28603);
nor UO_476 (O_476,N_29637,N_29791);
nand UO_477 (O_477,N_28780,N_28627);
nor UO_478 (O_478,N_28702,N_29515);
xor UO_479 (O_479,N_29133,N_29197);
xnor UO_480 (O_480,N_28917,N_29716);
and UO_481 (O_481,N_29310,N_28953);
or UO_482 (O_482,N_29419,N_28923);
and UO_483 (O_483,N_29203,N_28903);
and UO_484 (O_484,N_28976,N_29981);
and UO_485 (O_485,N_29044,N_29254);
nor UO_486 (O_486,N_29588,N_29145);
and UO_487 (O_487,N_29977,N_28576);
xnor UO_488 (O_488,N_28720,N_29135);
and UO_489 (O_489,N_29972,N_29941);
and UO_490 (O_490,N_29570,N_29080);
and UO_491 (O_491,N_29038,N_29635);
nand UO_492 (O_492,N_29119,N_29396);
nor UO_493 (O_493,N_29863,N_29587);
or UO_494 (O_494,N_29938,N_28888);
xor UO_495 (O_495,N_29902,N_29651);
nand UO_496 (O_496,N_28684,N_28725);
nor UO_497 (O_497,N_28504,N_28807);
xnor UO_498 (O_498,N_29681,N_29954);
xnor UO_499 (O_499,N_29004,N_29944);
nor UO_500 (O_500,N_29251,N_29556);
xnor UO_501 (O_501,N_29358,N_28779);
or UO_502 (O_502,N_29126,N_28604);
nand UO_503 (O_503,N_29614,N_29482);
and UO_504 (O_504,N_29231,N_28548);
and UO_505 (O_505,N_29143,N_29487);
or UO_506 (O_506,N_29402,N_29400);
and UO_507 (O_507,N_29078,N_29134);
or UO_508 (O_508,N_29069,N_29316);
nand UO_509 (O_509,N_28920,N_29767);
nor UO_510 (O_510,N_29282,N_29187);
nor UO_511 (O_511,N_28676,N_28918);
nor UO_512 (O_512,N_28963,N_29313);
and UO_513 (O_513,N_29407,N_28894);
and UO_514 (O_514,N_29179,N_29492);
xnor UO_515 (O_515,N_29815,N_29989);
nand UO_516 (O_516,N_29633,N_28890);
nor UO_517 (O_517,N_29735,N_29990);
and UO_518 (O_518,N_28970,N_28508);
nor UO_519 (O_519,N_29137,N_29268);
and UO_520 (O_520,N_29018,N_28997);
and UO_521 (O_521,N_29221,N_28795);
xor UO_522 (O_522,N_28852,N_29679);
or UO_523 (O_523,N_29728,N_29177);
and UO_524 (O_524,N_28530,N_29964);
and UO_525 (O_525,N_28661,N_28929);
or UO_526 (O_526,N_29898,N_28891);
or UO_527 (O_527,N_28784,N_29752);
or UO_528 (O_528,N_29921,N_28570);
nor UO_529 (O_529,N_29308,N_29063);
nor UO_530 (O_530,N_29974,N_29616);
nor UO_531 (O_531,N_29037,N_29607);
nor UO_532 (O_532,N_29262,N_29382);
nand UO_533 (O_533,N_29948,N_29459);
or UO_534 (O_534,N_29909,N_29805);
and UO_535 (O_535,N_29264,N_29826);
xor UO_536 (O_536,N_28706,N_28892);
or UO_537 (O_537,N_29473,N_29766);
nand UO_538 (O_538,N_29675,N_28873);
or UO_539 (O_539,N_29795,N_29715);
and UO_540 (O_540,N_29295,N_28736);
or UO_541 (O_541,N_29000,N_28856);
and UO_542 (O_542,N_28967,N_28516);
nor UO_543 (O_543,N_28563,N_28930);
nand UO_544 (O_544,N_29992,N_29141);
and UO_545 (O_545,N_29934,N_29269);
or UO_546 (O_546,N_29091,N_28952);
and UO_547 (O_547,N_29480,N_28673);
nor UO_548 (O_548,N_28913,N_29802);
xor UO_549 (O_549,N_29286,N_28834);
and UO_550 (O_550,N_28984,N_29462);
or UO_551 (O_551,N_29476,N_29630);
nand UO_552 (O_552,N_29808,N_29064);
xor UO_553 (O_553,N_29207,N_28671);
nand UO_554 (O_554,N_28753,N_29628);
or UO_555 (O_555,N_29105,N_29013);
and UO_556 (O_556,N_28713,N_29555);
nor UO_557 (O_557,N_29549,N_28885);
nand UO_558 (O_558,N_28591,N_29816);
xnor UO_559 (O_559,N_29755,N_29208);
nor UO_560 (O_560,N_29608,N_28948);
or UO_561 (O_561,N_29383,N_29798);
or UO_562 (O_562,N_28965,N_29583);
nand UO_563 (O_563,N_29836,N_29951);
nand UO_564 (O_564,N_29359,N_28707);
and UO_565 (O_565,N_28985,N_29079);
nor UO_566 (O_566,N_28659,N_29484);
nor UO_567 (O_567,N_28666,N_28598);
nand UO_568 (O_568,N_29265,N_28982);
and UO_569 (O_569,N_29410,N_29562);
or UO_570 (O_570,N_29585,N_28663);
and UO_571 (O_571,N_28752,N_29362);
nor UO_572 (O_572,N_29813,N_29167);
and UO_573 (O_573,N_29689,N_29070);
or UO_574 (O_574,N_29734,N_28650);
xnor UO_575 (O_575,N_28590,N_29101);
xor UO_576 (O_576,N_29403,N_29045);
nor UO_577 (O_577,N_29626,N_29228);
nor UO_578 (O_578,N_29540,N_29215);
and UO_579 (O_579,N_29672,N_29275);
or UO_580 (O_580,N_28715,N_28819);
nand UO_581 (O_581,N_29922,N_28822);
or UO_582 (O_582,N_28514,N_29293);
and UO_583 (O_583,N_28549,N_28827);
nor UO_584 (O_584,N_28642,N_29842);
nor UO_585 (O_585,N_29770,N_29047);
xor UO_586 (O_586,N_29998,N_28601);
nand UO_587 (O_587,N_28862,N_29121);
xor UO_588 (O_588,N_28575,N_29350);
nand UO_589 (O_589,N_29962,N_29108);
and UO_590 (O_590,N_28960,N_29573);
nand UO_591 (O_591,N_28602,N_28763);
or UO_592 (O_592,N_29741,N_29201);
or UO_593 (O_593,N_28867,N_29245);
or UO_594 (O_594,N_28804,N_29801);
or UO_595 (O_595,N_29099,N_29937);
xnor UO_596 (O_596,N_29448,N_29832);
and UO_597 (O_597,N_29878,N_28977);
xor UO_598 (O_598,N_29916,N_29880);
nand UO_599 (O_599,N_28731,N_28648);
and UO_600 (O_600,N_29907,N_29424);
nand UO_601 (O_601,N_29404,N_28630);
nor UO_602 (O_602,N_29475,N_28537);
nor UO_603 (O_603,N_28677,N_28561);
nand UO_604 (O_604,N_29217,N_29200);
or UO_605 (O_605,N_28721,N_29005);
and UO_606 (O_606,N_29170,N_29619);
or UO_607 (O_607,N_29506,N_28841);
xnor UO_608 (O_608,N_29271,N_29714);
nand UO_609 (O_609,N_29592,N_29241);
xnor UO_610 (O_610,N_29695,N_29349);
xor UO_611 (O_611,N_29864,N_28973);
and UO_612 (O_612,N_29322,N_29418);
nand UO_613 (O_613,N_29851,N_28992);
and UO_614 (O_614,N_28614,N_29743);
xnor UO_615 (O_615,N_29702,N_29212);
xor UO_616 (O_616,N_29758,N_29341);
or UO_617 (O_617,N_29796,N_29820);
nand UO_618 (O_618,N_29685,N_29354);
and UO_619 (O_619,N_29871,N_29821);
nand UO_620 (O_620,N_29711,N_28758);
and UO_621 (O_621,N_28796,N_29378);
nor UO_622 (O_622,N_29874,N_29209);
xor UO_623 (O_623,N_29092,N_29068);
or UO_624 (O_624,N_28766,N_29224);
and UO_625 (O_625,N_28555,N_28897);
nor UO_626 (O_626,N_29867,N_29578);
or UO_627 (O_627,N_29132,N_28727);
nand UO_628 (O_628,N_29627,N_28502);
and UO_629 (O_629,N_29580,N_28529);
and UO_630 (O_630,N_29582,N_28541);
nand UO_631 (O_631,N_28937,N_29075);
or UO_632 (O_632,N_28628,N_29750);
xnor UO_633 (O_633,N_28791,N_29011);
xnor UO_634 (O_634,N_28634,N_29883);
nand UO_635 (O_635,N_29790,N_28738);
nor UO_636 (O_636,N_29258,N_28820);
xnor UO_637 (O_637,N_28678,N_28566);
nor UO_638 (O_638,N_29819,N_29891);
and UO_639 (O_639,N_29596,N_29387);
or UO_640 (O_640,N_29664,N_29854);
nor UO_641 (O_641,N_29661,N_28593);
xor UO_642 (O_642,N_29486,N_28919);
nand UO_643 (O_643,N_28999,N_28765);
nand UO_644 (O_644,N_29097,N_28652);
nor UO_645 (O_645,N_29333,N_29850);
or UO_646 (O_646,N_29065,N_28646);
nand UO_647 (O_647,N_29046,N_29683);
and UO_648 (O_648,N_29409,N_29085);
or UO_649 (O_649,N_29324,N_29233);
xnor UO_650 (O_650,N_29260,N_29862);
xnor UO_651 (O_651,N_29894,N_29198);
nor UO_652 (O_652,N_29834,N_28944);
or UO_653 (O_653,N_29991,N_29704);
nor UO_654 (O_654,N_28838,N_29159);
xnor UO_655 (O_655,N_28679,N_29312);
and UO_656 (O_656,N_29445,N_29904);
nor UO_657 (O_657,N_28532,N_28543);
nand UO_658 (O_658,N_28755,N_29890);
nand UO_659 (O_659,N_29760,N_28818);
xor UO_660 (O_660,N_29950,N_28740);
nand UO_661 (O_661,N_29984,N_29160);
nor UO_662 (O_662,N_29053,N_29193);
nand UO_663 (O_663,N_29792,N_29389);
or UO_664 (O_664,N_28542,N_29017);
nor UO_665 (O_665,N_29340,N_29250);
and UO_666 (O_666,N_28613,N_29454);
nor UO_667 (O_667,N_29114,N_29130);
nand UO_668 (O_668,N_28510,N_29599);
and UO_669 (O_669,N_28501,N_29298);
nor UO_670 (O_670,N_28636,N_29705);
xnor UO_671 (O_671,N_29488,N_28993);
and UO_672 (O_672,N_28545,N_29510);
and UO_673 (O_673,N_28617,N_29498);
nor UO_674 (O_674,N_29899,N_29738);
and UO_675 (O_675,N_28889,N_29933);
and UO_676 (O_676,N_29379,N_29100);
nand UO_677 (O_677,N_28877,N_29041);
nand UO_678 (O_678,N_29604,N_29963);
and UO_679 (O_679,N_29720,N_29516);
xnor UO_680 (O_680,N_29875,N_29395);
nor UO_681 (O_681,N_29887,N_29112);
nand UO_682 (O_682,N_29059,N_29173);
nand UO_683 (O_683,N_28994,N_29232);
xor UO_684 (O_684,N_29749,N_28787);
or UO_685 (O_685,N_29371,N_29166);
or UO_686 (O_686,N_29162,N_29947);
or UO_687 (O_687,N_28975,N_29441);
and UO_688 (O_688,N_28808,N_29155);
xor UO_689 (O_689,N_29181,N_28835);
nor UO_690 (O_690,N_28524,N_29674);
and UO_691 (O_691,N_29031,N_28750);
nor UO_692 (O_692,N_29665,N_29014);
xnor UO_693 (O_693,N_29926,N_29356);
xnor UO_694 (O_694,N_29558,N_29885);
and UO_695 (O_695,N_29244,N_28547);
nor UO_696 (O_696,N_28812,N_29522);
or UO_697 (O_697,N_29873,N_29725);
and UO_698 (O_698,N_28503,N_29491);
xnor UO_699 (O_699,N_28644,N_29421);
nor UO_700 (O_700,N_28621,N_29107);
or UO_701 (O_701,N_29164,N_29960);
or UO_702 (O_702,N_28803,N_28770);
or UO_703 (O_703,N_28596,N_28853);
and UO_704 (O_704,N_28586,N_29828);
xnor UO_705 (O_705,N_29943,N_29869);
nand UO_706 (O_706,N_29737,N_28829);
xor UO_707 (O_707,N_29945,N_29640);
nor UO_708 (O_708,N_28660,N_29144);
nand UO_709 (O_709,N_29235,N_28585);
and UO_710 (O_710,N_29368,N_28823);
xor UO_711 (O_711,N_29156,N_29342);
nand UO_712 (O_712,N_29213,N_29997);
nor UO_713 (O_713,N_29157,N_29452);
or UO_714 (O_714,N_29055,N_29030);
and UO_715 (O_715,N_29154,N_29321);
and UO_716 (O_716,N_28564,N_29073);
nor UO_717 (O_717,N_29377,N_28704);
and UO_718 (O_718,N_29654,N_29856);
or UO_719 (O_719,N_29778,N_29812);
xnor UO_720 (O_720,N_28520,N_29463);
and UO_721 (O_721,N_29811,N_29334);
or UO_722 (O_722,N_29566,N_29521);
nor UO_723 (O_723,N_28647,N_28538);
nand UO_724 (O_724,N_29889,N_28800);
nor UO_725 (O_725,N_28859,N_29536);
and UO_726 (O_726,N_28664,N_28871);
or UO_727 (O_727,N_28932,N_29117);
nor UO_728 (O_728,N_29817,N_29605);
xnor UO_729 (O_729,N_29428,N_28651);
nor UO_730 (O_730,N_29481,N_29687);
nor UO_731 (O_731,N_28922,N_29505);
or UO_732 (O_732,N_29787,N_29118);
or UO_733 (O_733,N_28926,N_29346);
and UO_734 (O_734,N_29294,N_29494);
or UO_735 (O_735,N_29034,N_28745);
xor UO_736 (O_736,N_29225,N_29800);
xnor UO_737 (O_737,N_28657,N_29477);
nor UO_738 (O_738,N_29363,N_29401);
xor UO_739 (O_739,N_28552,N_28737);
nand UO_740 (O_740,N_29054,N_29551);
nand UO_741 (O_741,N_28683,N_29634);
or UO_742 (O_742,N_29174,N_29248);
and UO_743 (O_743,N_29172,N_29103);
nand UO_744 (O_744,N_29096,N_29973);
nand UO_745 (O_745,N_29710,N_28933);
nand UO_746 (O_746,N_28567,N_29351);
nor UO_747 (O_747,N_29746,N_29104);
or UO_748 (O_748,N_29315,N_29870);
and UO_749 (O_749,N_28747,N_29700);
xnor UO_750 (O_750,N_28504,N_29405);
nand UO_751 (O_751,N_29911,N_29832);
nor UO_752 (O_752,N_28988,N_28875);
or UO_753 (O_753,N_29092,N_29549);
nor UO_754 (O_754,N_28586,N_28937);
and UO_755 (O_755,N_29144,N_29026);
xnor UO_756 (O_756,N_29256,N_29190);
nand UO_757 (O_757,N_29355,N_29069);
nor UO_758 (O_758,N_29461,N_29433);
nand UO_759 (O_759,N_28845,N_28902);
nand UO_760 (O_760,N_29142,N_29978);
and UO_761 (O_761,N_29644,N_29666);
nor UO_762 (O_762,N_29690,N_28922);
and UO_763 (O_763,N_29812,N_29833);
and UO_764 (O_764,N_29165,N_29796);
nand UO_765 (O_765,N_28796,N_29660);
or UO_766 (O_766,N_29395,N_28926);
or UO_767 (O_767,N_29319,N_29438);
xnor UO_768 (O_768,N_29450,N_28891);
nand UO_769 (O_769,N_28820,N_28589);
xor UO_770 (O_770,N_29927,N_29650);
nor UO_771 (O_771,N_29169,N_29699);
nand UO_772 (O_772,N_28638,N_29062);
or UO_773 (O_773,N_29315,N_29474);
xor UO_774 (O_774,N_29992,N_29646);
nand UO_775 (O_775,N_29478,N_29474);
or UO_776 (O_776,N_29165,N_29239);
or UO_777 (O_777,N_29073,N_29833);
or UO_778 (O_778,N_29397,N_28749);
or UO_779 (O_779,N_28824,N_29493);
xnor UO_780 (O_780,N_28610,N_29425);
nand UO_781 (O_781,N_29087,N_29360);
or UO_782 (O_782,N_29420,N_28665);
and UO_783 (O_783,N_28981,N_29428);
or UO_784 (O_784,N_28927,N_28588);
nor UO_785 (O_785,N_29113,N_28982);
nand UO_786 (O_786,N_28985,N_29104);
nand UO_787 (O_787,N_29916,N_28931);
or UO_788 (O_788,N_29377,N_28535);
and UO_789 (O_789,N_29740,N_28973);
or UO_790 (O_790,N_28948,N_29044);
xnor UO_791 (O_791,N_29596,N_29547);
and UO_792 (O_792,N_28678,N_29552);
or UO_793 (O_793,N_29752,N_29470);
nand UO_794 (O_794,N_29560,N_28765);
and UO_795 (O_795,N_29242,N_29956);
xor UO_796 (O_796,N_29402,N_29210);
nor UO_797 (O_797,N_29299,N_29597);
and UO_798 (O_798,N_29266,N_29317);
or UO_799 (O_799,N_28817,N_29029);
nand UO_800 (O_800,N_29161,N_29725);
nand UO_801 (O_801,N_29990,N_29425);
and UO_802 (O_802,N_28727,N_29191);
or UO_803 (O_803,N_28893,N_29425);
and UO_804 (O_804,N_28681,N_28587);
nand UO_805 (O_805,N_28541,N_29125);
and UO_806 (O_806,N_28669,N_28723);
and UO_807 (O_807,N_28933,N_29269);
and UO_808 (O_808,N_29699,N_29230);
nand UO_809 (O_809,N_29130,N_29426);
or UO_810 (O_810,N_29956,N_28706);
and UO_811 (O_811,N_29088,N_29542);
and UO_812 (O_812,N_29299,N_29023);
nor UO_813 (O_813,N_28501,N_29177);
nor UO_814 (O_814,N_29303,N_28708);
nand UO_815 (O_815,N_28768,N_28943);
nor UO_816 (O_816,N_29410,N_28533);
nand UO_817 (O_817,N_28891,N_29522);
or UO_818 (O_818,N_29614,N_29527);
nand UO_819 (O_819,N_28810,N_29135);
xor UO_820 (O_820,N_28856,N_29246);
xnor UO_821 (O_821,N_28737,N_29280);
xnor UO_822 (O_822,N_29598,N_29190);
nand UO_823 (O_823,N_29128,N_29712);
and UO_824 (O_824,N_28651,N_29974);
or UO_825 (O_825,N_29187,N_29821);
and UO_826 (O_826,N_28560,N_29705);
xor UO_827 (O_827,N_28607,N_28510);
and UO_828 (O_828,N_29744,N_29836);
nor UO_829 (O_829,N_29768,N_28875);
and UO_830 (O_830,N_29479,N_28684);
xor UO_831 (O_831,N_29969,N_29604);
xnor UO_832 (O_832,N_29241,N_28833);
xnor UO_833 (O_833,N_29437,N_29259);
nand UO_834 (O_834,N_28665,N_29080);
nor UO_835 (O_835,N_29560,N_28809);
xor UO_836 (O_836,N_29019,N_29398);
or UO_837 (O_837,N_28613,N_29147);
nor UO_838 (O_838,N_29594,N_29057);
and UO_839 (O_839,N_29019,N_28653);
nand UO_840 (O_840,N_28706,N_28758);
nand UO_841 (O_841,N_29020,N_28892);
xor UO_842 (O_842,N_29385,N_28793);
xnor UO_843 (O_843,N_28537,N_29605);
nand UO_844 (O_844,N_29375,N_29941);
and UO_845 (O_845,N_29661,N_29853);
nor UO_846 (O_846,N_29019,N_29926);
and UO_847 (O_847,N_28779,N_29746);
and UO_848 (O_848,N_28884,N_28628);
nor UO_849 (O_849,N_28993,N_28672);
or UO_850 (O_850,N_28861,N_29687);
nand UO_851 (O_851,N_28817,N_29824);
xor UO_852 (O_852,N_29786,N_28871);
xnor UO_853 (O_853,N_29272,N_29500);
and UO_854 (O_854,N_29051,N_29580);
and UO_855 (O_855,N_28970,N_29574);
nand UO_856 (O_856,N_29995,N_28686);
nand UO_857 (O_857,N_28818,N_29356);
nor UO_858 (O_858,N_28813,N_29067);
nor UO_859 (O_859,N_29987,N_29439);
nor UO_860 (O_860,N_29830,N_29479);
nand UO_861 (O_861,N_29155,N_29640);
xor UO_862 (O_862,N_29829,N_29315);
and UO_863 (O_863,N_29820,N_28777);
and UO_864 (O_864,N_28840,N_28900);
xor UO_865 (O_865,N_29873,N_29229);
nor UO_866 (O_866,N_28907,N_28569);
nor UO_867 (O_867,N_29991,N_28770);
and UO_868 (O_868,N_29508,N_28655);
xnor UO_869 (O_869,N_29713,N_28813);
nor UO_870 (O_870,N_29631,N_29800);
nor UO_871 (O_871,N_29445,N_29475);
nor UO_872 (O_872,N_29589,N_29368);
nand UO_873 (O_873,N_29092,N_28747);
xor UO_874 (O_874,N_29004,N_29561);
or UO_875 (O_875,N_29238,N_29218);
or UO_876 (O_876,N_29526,N_29870);
nor UO_877 (O_877,N_29710,N_28891);
and UO_878 (O_878,N_28502,N_29043);
or UO_879 (O_879,N_29945,N_29594);
nor UO_880 (O_880,N_29774,N_29379);
xor UO_881 (O_881,N_29409,N_29125);
and UO_882 (O_882,N_28801,N_29552);
or UO_883 (O_883,N_28559,N_29759);
xor UO_884 (O_884,N_28740,N_29848);
or UO_885 (O_885,N_29045,N_29431);
or UO_886 (O_886,N_28688,N_28673);
xnor UO_887 (O_887,N_29546,N_28977);
or UO_888 (O_888,N_29571,N_28668);
nand UO_889 (O_889,N_29032,N_28605);
nor UO_890 (O_890,N_29069,N_28771);
nor UO_891 (O_891,N_29081,N_28532);
and UO_892 (O_892,N_29380,N_28612);
or UO_893 (O_893,N_29947,N_29568);
or UO_894 (O_894,N_28663,N_29487);
or UO_895 (O_895,N_29299,N_29793);
xor UO_896 (O_896,N_29155,N_28666);
nor UO_897 (O_897,N_29674,N_29901);
and UO_898 (O_898,N_29828,N_28634);
and UO_899 (O_899,N_29440,N_29345);
nand UO_900 (O_900,N_29083,N_29406);
or UO_901 (O_901,N_29990,N_29192);
nor UO_902 (O_902,N_29901,N_28570);
xor UO_903 (O_903,N_29565,N_28716);
or UO_904 (O_904,N_29027,N_29296);
xnor UO_905 (O_905,N_29707,N_28712);
xor UO_906 (O_906,N_29515,N_28670);
nor UO_907 (O_907,N_29011,N_29741);
nor UO_908 (O_908,N_29447,N_29435);
nor UO_909 (O_909,N_28934,N_28507);
and UO_910 (O_910,N_29199,N_29972);
and UO_911 (O_911,N_28846,N_29455);
xnor UO_912 (O_912,N_29528,N_28822);
or UO_913 (O_913,N_29913,N_29247);
or UO_914 (O_914,N_29362,N_29217);
nor UO_915 (O_915,N_28838,N_29486);
or UO_916 (O_916,N_29951,N_28672);
and UO_917 (O_917,N_28744,N_29384);
or UO_918 (O_918,N_29465,N_29082);
xor UO_919 (O_919,N_29754,N_29554);
or UO_920 (O_920,N_29331,N_29819);
nand UO_921 (O_921,N_29868,N_29336);
or UO_922 (O_922,N_29677,N_29573);
nand UO_923 (O_923,N_29115,N_29488);
or UO_924 (O_924,N_28970,N_29603);
nand UO_925 (O_925,N_28748,N_29940);
or UO_926 (O_926,N_29580,N_29702);
nor UO_927 (O_927,N_28961,N_29191);
or UO_928 (O_928,N_28610,N_29221);
xor UO_929 (O_929,N_29210,N_28614);
or UO_930 (O_930,N_28606,N_28544);
nor UO_931 (O_931,N_29080,N_28973);
nor UO_932 (O_932,N_28693,N_28550);
xnor UO_933 (O_933,N_28840,N_29031);
nand UO_934 (O_934,N_28676,N_29937);
or UO_935 (O_935,N_28712,N_29206);
nor UO_936 (O_936,N_28987,N_29494);
nand UO_937 (O_937,N_28766,N_28735);
or UO_938 (O_938,N_29874,N_29865);
or UO_939 (O_939,N_29954,N_29503);
nand UO_940 (O_940,N_29967,N_29080);
and UO_941 (O_941,N_28821,N_28674);
or UO_942 (O_942,N_28687,N_29249);
and UO_943 (O_943,N_29859,N_29405);
nand UO_944 (O_944,N_29562,N_29792);
nand UO_945 (O_945,N_29519,N_29997);
xor UO_946 (O_946,N_28598,N_29326);
or UO_947 (O_947,N_29890,N_29859);
nand UO_948 (O_948,N_29305,N_28507);
nand UO_949 (O_949,N_29145,N_29676);
or UO_950 (O_950,N_29034,N_28696);
and UO_951 (O_951,N_29531,N_29203);
or UO_952 (O_952,N_29027,N_28618);
or UO_953 (O_953,N_29400,N_29859);
nand UO_954 (O_954,N_28984,N_29883);
or UO_955 (O_955,N_28521,N_28959);
xor UO_956 (O_956,N_29693,N_28830);
nor UO_957 (O_957,N_28905,N_29168);
or UO_958 (O_958,N_29908,N_28759);
and UO_959 (O_959,N_28695,N_28786);
xnor UO_960 (O_960,N_28547,N_29034);
xor UO_961 (O_961,N_29013,N_29858);
xnor UO_962 (O_962,N_28573,N_28941);
and UO_963 (O_963,N_28767,N_28714);
and UO_964 (O_964,N_29399,N_29061);
xor UO_965 (O_965,N_29050,N_29421);
and UO_966 (O_966,N_28815,N_29409);
nand UO_967 (O_967,N_29683,N_29808);
and UO_968 (O_968,N_29208,N_29142);
nand UO_969 (O_969,N_29056,N_28929);
nor UO_970 (O_970,N_29494,N_29477);
nor UO_971 (O_971,N_28681,N_29434);
and UO_972 (O_972,N_29378,N_29001);
or UO_973 (O_973,N_29530,N_29034);
nand UO_974 (O_974,N_28611,N_28716);
nand UO_975 (O_975,N_29005,N_29404);
xnor UO_976 (O_976,N_29711,N_29670);
nand UO_977 (O_977,N_29066,N_29490);
nand UO_978 (O_978,N_28765,N_29329);
nand UO_979 (O_979,N_28903,N_29393);
xnor UO_980 (O_980,N_29742,N_28963);
or UO_981 (O_981,N_29920,N_29249);
nand UO_982 (O_982,N_29520,N_28634);
or UO_983 (O_983,N_28716,N_29377);
xnor UO_984 (O_984,N_29016,N_28759);
nand UO_985 (O_985,N_28714,N_29587);
nand UO_986 (O_986,N_29287,N_29264);
nor UO_987 (O_987,N_29051,N_28507);
and UO_988 (O_988,N_29227,N_29381);
and UO_989 (O_989,N_28647,N_29056);
or UO_990 (O_990,N_28535,N_28989);
and UO_991 (O_991,N_29243,N_29563);
and UO_992 (O_992,N_29956,N_28968);
nor UO_993 (O_993,N_29400,N_28574);
or UO_994 (O_994,N_29280,N_29652);
nor UO_995 (O_995,N_28650,N_29244);
or UO_996 (O_996,N_29462,N_28680);
or UO_997 (O_997,N_28950,N_28788);
nor UO_998 (O_998,N_29202,N_28521);
and UO_999 (O_999,N_29017,N_29289);
nor UO_1000 (O_1000,N_28539,N_29338);
nor UO_1001 (O_1001,N_28865,N_28859);
and UO_1002 (O_1002,N_29721,N_29901);
nand UO_1003 (O_1003,N_29076,N_28523);
and UO_1004 (O_1004,N_29085,N_28702);
nor UO_1005 (O_1005,N_29524,N_28972);
nand UO_1006 (O_1006,N_29801,N_29136);
and UO_1007 (O_1007,N_29010,N_29321);
nand UO_1008 (O_1008,N_28650,N_29008);
nor UO_1009 (O_1009,N_28590,N_29366);
and UO_1010 (O_1010,N_29850,N_29887);
nand UO_1011 (O_1011,N_29780,N_28608);
nor UO_1012 (O_1012,N_28717,N_29012);
or UO_1013 (O_1013,N_29987,N_28941);
nand UO_1014 (O_1014,N_28633,N_29677);
or UO_1015 (O_1015,N_29377,N_29531);
nand UO_1016 (O_1016,N_28753,N_29116);
or UO_1017 (O_1017,N_29386,N_28656);
nand UO_1018 (O_1018,N_28809,N_29687);
nand UO_1019 (O_1019,N_29883,N_29863);
or UO_1020 (O_1020,N_29819,N_29525);
nand UO_1021 (O_1021,N_28856,N_29829);
xor UO_1022 (O_1022,N_29091,N_28878);
nor UO_1023 (O_1023,N_28934,N_28769);
nor UO_1024 (O_1024,N_29712,N_29652);
or UO_1025 (O_1025,N_29264,N_29101);
xor UO_1026 (O_1026,N_29146,N_29058);
xor UO_1027 (O_1027,N_29771,N_29132);
xor UO_1028 (O_1028,N_28597,N_29737);
or UO_1029 (O_1029,N_28953,N_29932);
xor UO_1030 (O_1030,N_29975,N_29259);
nor UO_1031 (O_1031,N_28729,N_28579);
nand UO_1032 (O_1032,N_29751,N_29450);
nand UO_1033 (O_1033,N_29502,N_29240);
or UO_1034 (O_1034,N_29583,N_29352);
nand UO_1035 (O_1035,N_29824,N_28899);
xnor UO_1036 (O_1036,N_29564,N_29229);
xnor UO_1037 (O_1037,N_29768,N_28982);
xor UO_1038 (O_1038,N_28891,N_29403);
nor UO_1039 (O_1039,N_29966,N_29055);
or UO_1040 (O_1040,N_29674,N_29797);
nand UO_1041 (O_1041,N_28880,N_29208);
xor UO_1042 (O_1042,N_29238,N_29082);
or UO_1043 (O_1043,N_29129,N_28566);
or UO_1044 (O_1044,N_29047,N_28872);
nor UO_1045 (O_1045,N_28549,N_29670);
and UO_1046 (O_1046,N_28864,N_29656);
nor UO_1047 (O_1047,N_29214,N_29734);
or UO_1048 (O_1048,N_29872,N_29084);
and UO_1049 (O_1049,N_29059,N_29956);
and UO_1050 (O_1050,N_29612,N_29524);
or UO_1051 (O_1051,N_29347,N_29670);
nor UO_1052 (O_1052,N_28579,N_28524);
xor UO_1053 (O_1053,N_29895,N_28671);
nor UO_1054 (O_1054,N_29361,N_29619);
xnor UO_1055 (O_1055,N_29764,N_29780);
or UO_1056 (O_1056,N_29431,N_29133);
and UO_1057 (O_1057,N_28936,N_29994);
xor UO_1058 (O_1058,N_29000,N_28952);
nor UO_1059 (O_1059,N_29797,N_28848);
or UO_1060 (O_1060,N_29070,N_28761);
nor UO_1061 (O_1061,N_28733,N_28698);
or UO_1062 (O_1062,N_29713,N_29456);
nand UO_1063 (O_1063,N_29901,N_29557);
nand UO_1064 (O_1064,N_28660,N_28865);
or UO_1065 (O_1065,N_29409,N_29009);
and UO_1066 (O_1066,N_29539,N_28563);
xnor UO_1067 (O_1067,N_29543,N_29702);
and UO_1068 (O_1068,N_29939,N_29561);
xor UO_1069 (O_1069,N_28992,N_29983);
nor UO_1070 (O_1070,N_29953,N_29932);
and UO_1071 (O_1071,N_29461,N_29458);
or UO_1072 (O_1072,N_29299,N_28708);
nand UO_1073 (O_1073,N_29489,N_28873);
and UO_1074 (O_1074,N_28752,N_28920);
nand UO_1075 (O_1075,N_29892,N_28829);
or UO_1076 (O_1076,N_29778,N_29541);
xnor UO_1077 (O_1077,N_29918,N_29882);
and UO_1078 (O_1078,N_29018,N_28909);
nand UO_1079 (O_1079,N_28636,N_28739);
nand UO_1080 (O_1080,N_29127,N_29512);
nor UO_1081 (O_1081,N_28872,N_29168);
xor UO_1082 (O_1082,N_29809,N_29061);
nor UO_1083 (O_1083,N_28650,N_29259);
and UO_1084 (O_1084,N_29532,N_29901);
nor UO_1085 (O_1085,N_28701,N_29459);
nor UO_1086 (O_1086,N_29178,N_29620);
nor UO_1087 (O_1087,N_29350,N_29558);
and UO_1088 (O_1088,N_28997,N_28784);
or UO_1089 (O_1089,N_29558,N_28741);
nand UO_1090 (O_1090,N_28832,N_28724);
xor UO_1091 (O_1091,N_28992,N_28730);
nor UO_1092 (O_1092,N_29552,N_29932);
nand UO_1093 (O_1093,N_29272,N_29242);
nor UO_1094 (O_1094,N_29297,N_28554);
xnor UO_1095 (O_1095,N_29555,N_29442);
and UO_1096 (O_1096,N_29627,N_29450);
nor UO_1097 (O_1097,N_28537,N_29521);
xor UO_1098 (O_1098,N_29799,N_29912);
or UO_1099 (O_1099,N_28981,N_29534);
and UO_1100 (O_1100,N_28683,N_29134);
xor UO_1101 (O_1101,N_29932,N_29145);
nand UO_1102 (O_1102,N_29993,N_29064);
nand UO_1103 (O_1103,N_29043,N_29566);
nor UO_1104 (O_1104,N_28585,N_28704);
and UO_1105 (O_1105,N_29850,N_28678);
or UO_1106 (O_1106,N_28655,N_29474);
nand UO_1107 (O_1107,N_29373,N_29509);
or UO_1108 (O_1108,N_29121,N_29337);
nor UO_1109 (O_1109,N_28511,N_28911);
and UO_1110 (O_1110,N_29159,N_29861);
nor UO_1111 (O_1111,N_29326,N_29827);
xnor UO_1112 (O_1112,N_29698,N_28663);
nand UO_1113 (O_1113,N_29832,N_29302);
and UO_1114 (O_1114,N_28944,N_28864);
xor UO_1115 (O_1115,N_28589,N_29302);
and UO_1116 (O_1116,N_29620,N_29593);
or UO_1117 (O_1117,N_29161,N_29999);
and UO_1118 (O_1118,N_28683,N_29793);
nand UO_1119 (O_1119,N_29795,N_29145);
or UO_1120 (O_1120,N_29954,N_28971);
xnor UO_1121 (O_1121,N_29345,N_29575);
and UO_1122 (O_1122,N_28659,N_29446);
xor UO_1123 (O_1123,N_29412,N_28750);
and UO_1124 (O_1124,N_29810,N_29453);
nor UO_1125 (O_1125,N_29103,N_29625);
or UO_1126 (O_1126,N_29222,N_29560);
and UO_1127 (O_1127,N_28574,N_28726);
and UO_1128 (O_1128,N_29193,N_28845);
nand UO_1129 (O_1129,N_28590,N_29476);
or UO_1130 (O_1130,N_29894,N_29319);
or UO_1131 (O_1131,N_29019,N_28765);
and UO_1132 (O_1132,N_29937,N_29891);
or UO_1133 (O_1133,N_29451,N_28942);
or UO_1134 (O_1134,N_29447,N_28533);
nand UO_1135 (O_1135,N_28700,N_29812);
nor UO_1136 (O_1136,N_29909,N_29858);
or UO_1137 (O_1137,N_28759,N_29632);
and UO_1138 (O_1138,N_29103,N_29487);
or UO_1139 (O_1139,N_29182,N_28874);
xor UO_1140 (O_1140,N_28954,N_29262);
nor UO_1141 (O_1141,N_29879,N_29633);
or UO_1142 (O_1142,N_29089,N_29305);
and UO_1143 (O_1143,N_28942,N_28532);
xnor UO_1144 (O_1144,N_28588,N_29396);
or UO_1145 (O_1145,N_29142,N_28737);
or UO_1146 (O_1146,N_29028,N_29824);
and UO_1147 (O_1147,N_29182,N_29102);
or UO_1148 (O_1148,N_29433,N_29408);
xnor UO_1149 (O_1149,N_29621,N_29347);
nor UO_1150 (O_1150,N_29478,N_28847);
and UO_1151 (O_1151,N_28773,N_29701);
xor UO_1152 (O_1152,N_29921,N_29314);
xnor UO_1153 (O_1153,N_28574,N_29827);
nand UO_1154 (O_1154,N_29234,N_28631);
nand UO_1155 (O_1155,N_28900,N_28752);
xor UO_1156 (O_1156,N_29613,N_28888);
and UO_1157 (O_1157,N_28646,N_29238);
nor UO_1158 (O_1158,N_29813,N_28902);
xor UO_1159 (O_1159,N_28890,N_29281);
and UO_1160 (O_1160,N_29855,N_28703);
xnor UO_1161 (O_1161,N_28644,N_29054);
nor UO_1162 (O_1162,N_29272,N_28996);
or UO_1163 (O_1163,N_29456,N_28995);
nor UO_1164 (O_1164,N_29864,N_28936);
and UO_1165 (O_1165,N_28970,N_29006);
nor UO_1166 (O_1166,N_29958,N_28921);
xor UO_1167 (O_1167,N_29044,N_29120);
nor UO_1168 (O_1168,N_29039,N_28890);
xor UO_1169 (O_1169,N_29833,N_29786);
and UO_1170 (O_1170,N_29144,N_28813);
nor UO_1171 (O_1171,N_29121,N_29178);
or UO_1172 (O_1172,N_29847,N_29141);
nand UO_1173 (O_1173,N_29552,N_28725);
nor UO_1174 (O_1174,N_29899,N_29924);
or UO_1175 (O_1175,N_28773,N_29950);
and UO_1176 (O_1176,N_29413,N_29980);
or UO_1177 (O_1177,N_29079,N_29180);
nor UO_1178 (O_1178,N_28549,N_29461);
xnor UO_1179 (O_1179,N_28753,N_29597);
and UO_1180 (O_1180,N_28617,N_29868);
nor UO_1181 (O_1181,N_29581,N_28850);
nand UO_1182 (O_1182,N_29171,N_29107);
and UO_1183 (O_1183,N_29315,N_29780);
and UO_1184 (O_1184,N_28677,N_28939);
or UO_1185 (O_1185,N_29061,N_29438);
or UO_1186 (O_1186,N_29169,N_28856);
or UO_1187 (O_1187,N_28529,N_29371);
nor UO_1188 (O_1188,N_28743,N_28541);
or UO_1189 (O_1189,N_29763,N_29290);
and UO_1190 (O_1190,N_29570,N_29963);
or UO_1191 (O_1191,N_29917,N_29653);
nor UO_1192 (O_1192,N_29975,N_29888);
nor UO_1193 (O_1193,N_29336,N_29405);
and UO_1194 (O_1194,N_29389,N_29974);
xnor UO_1195 (O_1195,N_29664,N_29634);
or UO_1196 (O_1196,N_29616,N_29844);
nor UO_1197 (O_1197,N_29363,N_29410);
nand UO_1198 (O_1198,N_29778,N_28588);
and UO_1199 (O_1199,N_28810,N_28510);
or UO_1200 (O_1200,N_28777,N_29178);
nand UO_1201 (O_1201,N_28936,N_29510);
xor UO_1202 (O_1202,N_28982,N_29344);
xnor UO_1203 (O_1203,N_29755,N_29780);
xor UO_1204 (O_1204,N_28712,N_29202);
xnor UO_1205 (O_1205,N_29927,N_29372);
nand UO_1206 (O_1206,N_29871,N_29926);
nor UO_1207 (O_1207,N_29057,N_29486);
or UO_1208 (O_1208,N_29344,N_29040);
or UO_1209 (O_1209,N_29631,N_28524);
xnor UO_1210 (O_1210,N_28706,N_29929);
and UO_1211 (O_1211,N_29286,N_29145);
or UO_1212 (O_1212,N_28708,N_29931);
xor UO_1213 (O_1213,N_29534,N_29447);
nand UO_1214 (O_1214,N_29846,N_28655);
and UO_1215 (O_1215,N_29980,N_29729);
nor UO_1216 (O_1216,N_29874,N_29342);
and UO_1217 (O_1217,N_29588,N_28969);
and UO_1218 (O_1218,N_29522,N_29861);
and UO_1219 (O_1219,N_29251,N_29340);
xor UO_1220 (O_1220,N_29034,N_29950);
or UO_1221 (O_1221,N_29000,N_29564);
and UO_1222 (O_1222,N_28550,N_28628);
nor UO_1223 (O_1223,N_29020,N_28536);
and UO_1224 (O_1224,N_28824,N_28724);
or UO_1225 (O_1225,N_28710,N_29253);
xor UO_1226 (O_1226,N_29754,N_29750);
xnor UO_1227 (O_1227,N_29769,N_28920);
nor UO_1228 (O_1228,N_29148,N_28827);
and UO_1229 (O_1229,N_29852,N_28556);
or UO_1230 (O_1230,N_29085,N_29469);
or UO_1231 (O_1231,N_29906,N_28650);
xnor UO_1232 (O_1232,N_29579,N_29071);
or UO_1233 (O_1233,N_29459,N_29083);
xor UO_1234 (O_1234,N_29997,N_28666);
xnor UO_1235 (O_1235,N_28526,N_28948);
or UO_1236 (O_1236,N_29207,N_28563);
xor UO_1237 (O_1237,N_28827,N_29500);
or UO_1238 (O_1238,N_29950,N_29231);
and UO_1239 (O_1239,N_29108,N_29436);
or UO_1240 (O_1240,N_29000,N_29072);
nor UO_1241 (O_1241,N_28747,N_29684);
or UO_1242 (O_1242,N_29010,N_29803);
nand UO_1243 (O_1243,N_28559,N_29687);
nand UO_1244 (O_1244,N_29931,N_28767);
and UO_1245 (O_1245,N_29554,N_29111);
nand UO_1246 (O_1246,N_29984,N_29535);
nand UO_1247 (O_1247,N_28849,N_29369);
xor UO_1248 (O_1248,N_28640,N_28946);
nor UO_1249 (O_1249,N_29089,N_29447);
or UO_1250 (O_1250,N_28711,N_28575);
or UO_1251 (O_1251,N_29800,N_29146);
nor UO_1252 (O_1252,N_29078,N_28554);
nand UO_1253 (O_1253,N_28962,N_29013);
xnor UO_1254 (O_1254,N_28646,N_28838);
xnor UO_1255 (O_1255,N_28521,N_29167);
nand UO_1256 (O_1256,N_29743,N_29579);
or UO_1257 (O_1257,N_28536,N_28641);
or UO_1258 (O_1258,N_28561,N_29667);
and UO_1259 (O_1259,N_29704,N_29979);
xor UO_1260 (O_1260,N_29762,N_29265);
and UO_1261 (O_1261,N_29006,N_28963);
or UO_1262 (O_1262,N_29516,N_29180);
nand UO_1263 (O_1263,N_28918,N_29997);
or UO_1264 (O_1264,N_29412,N_28607);
and UO_1265 (O_1265,N_28975,N_28802);
and UO_1266 (O_1266,N_29091,N_29848);
or UO_1267 (O_1267,N_29786,N_28868);
xor UO_1268 (O_1268,N_28916,N_28732);
or UO_1269 (O_1269,N_29347,N_29019);
nor UO_1270 (O_1270,N_28829,N_29362);
nor UO_1271 (O_1271,N_29716,N_29486);
and UO_1272 (O_1272,N_28887,N_29888);
or UO_1273 (O_1273,N_29941,N_28974);
or UO_1274 (O_1274,N_29897,N_29816);
nor UO_1275 (O_1275,N_29388,N_29019);
or UO_1276 (O_1276,N_28689,N_29655);
and UO_1277 (O_1277,N_29618,N_28857);
xor UO_1278 (O_1278,N_29259,N_29721);
and UO_1279 (O_1279,N_28811,N_29166);
nor UO_1280 (O_1280,N_29650,N_28540);
nor UO_1281 (O_1281,N_28715,N_29122);
nand UO_1282 (O_1282,N_29953,N_28508);
xnor UO_1283 (O_1283,N_29828,N_28546);
and UO_1284 (O_1284,N_29679,N_29364);
nor UO_1285 (O_1285,N_29892,N_29793);
or UO_1286 (O_1286,N_29239,N_29823);
xor UO_1287 (O_1287,N_29216,N_29076);
or UO_1288 (O_1288,N_28764,N_28969);
nand UO_1289 (O_1289,N_29399,N_29067);
nand UO_1290 (O_1290,N_29030,N_29124);
nand UO_1291 (O_1291,N_29868,N_28543);
or UO_1292 (O_1292,N_29433,N_28921);
and UO_1293 (O_1293,N_29029,N_29773);
xnor UO_1294 (O_1294,N_29442,N_29956);
nand UO_1295 (O_1295,N_29136,N_29595);
or UO_1296 (O_1296,N_29586,N_28722);
nand UO_1297 (O_1297,N_28944,N_28933);
xor UO_1298 (O_1298,N_29924,N_29916);
and UO_1299 (O_1299,N_28833,N_29199);
and UO_1300 (O_1300,N_29176,N_29997);
xnor UO_1301 (O_1301,N_29378,N_28688);
nand UO_1302 (O_1302,N_29898,N_28852);
xnor UO_1303 (O_1303,N_28811,N_29516);
nand UO_1304 (O_1304,N_29740,N_28729);
and UO_1305 (O_1305,N_28640,N_28863);
nand UO_1306 (O_1306,N_28678,N_28712);
nand UO_1307 (O_1307,N_28870,N_29686);
xor UO_1308 (O_1308,N_29004,N_28775);
xnor UO_1309 (O_1309,N_29194,N_29886);
xor UO_1310 (O_1310,N_29577,N_28937);
nand UO_1311 (O_1311,N_29700,N_29368);
and UO_1312 (O_1312,N_29600,N_29006);
or UO_1313 (O_1313,N_29468,N_29816);
and UO_1314 (O_1314,N_29374,N_29093);
nor UO_1315 (O_1315,N_28629,N_29967);
and UO_1316 (O_1316,N_29636,N_29112);
xor UO_1317 (O_1317,N_29859,N_28945);
nand UO_1318 (O_1318,N_29680,N_28814);
nor UO_1319 (O_1319,N_29881,N_29386);
nand UO_1320 (O_1320,N_29314,N_29949);
and UO_1321 (O_1321,N_29009,N_29853);
or UO_1322 (O_1322,N_29144,N_29931);
or UO_1323 (O_1323,N_29652,N_29440);
or UO_1324 (O_1324,N_28849,N_29742);
nand UO_1325 (O_1325,N_28893,N_29564);
nand UO_1326 (O_1326,N_29838,N_29019);
or UO_1327 (O_1327,N_29170,N_29142);
nor UO_1328 (O_1328,N_28511,N_29692);
or UO_1329 (O_1329,N_29342,N_28791);
and UO_1330 (O_1330,N_29599,N_28957);
nand UO_1331 (O_1331,N_29410,N_29791);
and UO_1332 (O_1332,N_29810,N_28796);
xnor UO_1333 (O_1333,N_29294,N_29011);
xor UO_1334 (O_1334,N_28771,N_29859);
xnor UO_1335 (O_1335,N_28753,N_29683);
and UO_1336 (O_1336,N_28500,N_29402);
nor UO_1337 (O_1337,N_28578,N_29794);
nor UO_1338 (O_1338,N_28687,N_29407);
xnor UO_1339 (O_1339,N_28526,N_29869);
xor UO_1340 (O_1340,N_29050,N_29514);
xnor UO_1341 (O_1341,N_29310,N_29575);
xor UO_1342 (O_1342,N_28984,N_29759);
or UO_1343 (O_1343,N_29497,N_29687);
or UO_1344 (O_1344,N_29246,N_29642);
xnor UO_1345 (O_1345,N_29008,N_29535);
and UO_1346 (O_1346,N_28657,N_29708);
nor UO_1347 (O_1347,N_29433,N_29960);
nand UO_1348 (O_1348,N_29162,N_29570);
nand UO_1349 (O_1349,N_28973,N_29381);
xnor UO_1350 (O_1350,N_28871,N_29128);
nand UO_1351 (O_1351,N_29517,N_28836);
and UO_1352 (O_1352,N_29627,N_29171);
and UO_1353 (O_1353,N_29701,N_29022);
xnor UO_1354 (O_1354,N_29927,N_28950);
xnor UO_1355 (O_1355,N_28757,N_29122);
or UO_1356 (O_1356,N_29572,N_29654);
nor UO_1357 (O_1357,N_29979,N_29206);
or UO_1358 (O_1358,N_29781,N_28664);
nor UO_1359 (O_1359,N_29138,N_29702);
or UO_1360 (O_1360,N_28725,N_29365);
and UO_1361 (O_1361,N_29215,N_29619);
nor UO_1362 (O_1362,N_28670,N_29928);
xnor UO_1363 (O_1363,N_29320,N_29564);
nand UO_1364 (O_1364,N_28944,N_28953);
and UO_1365 (O_1365,N_28622,N_29829);
xor UO_1366 (O_1366,N_29300,N_29568);
and UO_1367 (O_1367,N_29826,N_28846);
xnor UO_1368 (O_1368,N_28758,N_29760);
nand UO_1369 (O_1369,N_29466,N_28630);
and UO_1370 (O_1370,N_29152,N_29786);
nor UO_1371 (O_1371,N_28698,N_28813);
xor UO_1372 (O_1372,N_29030,N_29058);
nand UO_1373 (O_1373,N_29588,N_28516);
nor UO_1374 (O_1374,N_29571,N_29475);
xnor UO_1375 (O_1375,N_28937,N_28636);
and UO_1376 (O_1376,N_29245,N_29035);
nor UO_1377 (O_1377,N_28699,N_29573);
nor UO_1378 (O_1378,N_29445,N_28848);
and UO_1379 (O_1379,N_29937,N_28905);
xor UO_1380 (O_1380,N_29254,N_29084);
xor UO_1381 (O_1381,N_29392,N_29528);
nand UO_1382 (O_1382,N_29104,N_29793);
nand UO_1383 (O_1383,N_28922,N_29642);
nand UO_1384 (O_1384,N_28755,N_29129);
and UO_1385 (O_1385,N_29594,N_28698);
nand UO_1386 (O_1386,N_29283,N_29372);
or UO_1387 (O_1387,N_29713,N_28513);
nand UO_1388 (O_1388,N_28924,N_29239);
xor UO_1389 (O_1389,N_29451,N_29944);
nand UO_1390 (O_1390,N_28982,N_29398);
or UO_1391 (O_1391,N_29072,N_28959);
nand UO_1392 (O_1392,N_29138,N_29713);
xnor UO_1393 (O_1393,N_28975,N_28749);
nand UO_1394 (O_1394,N_28831,N_29466);
and UO_1395 (O_1395,N_29980,N_28680);
nor UO_1396 (O_1396,N_29203,N_28810);
or UO_1397 (O_1397,N_29609,N_29526);
and UO_1398 (O_1398,N_29596,N_29314);
nand UO_1399 (O_1399,N_29054,N_29492);
or UO_1400 (O_1400,N_28900,N_28556);
and UO_1401 (O_1401,N_29150,N_29448);
nand UO_1402 (O_1402,N_28963,N_29931);
and UO_1403 (O_1403,N_29254,N_29395);
or UO_1404 (O_1404,N_29805,N_29889);
nor UO_1405 (O_1405,N_29250,N_28959);
or UO_1406 (O_1406,N_28977,N_28871);
nor UO_1407 (O_1407,N_28567,N_28756);
and UO_1408 (O_1408,N_28665,N_28664);
nand UO_1409 (O_1409,N_29169,N_28855);
or UO_1410 (O_1410,N_28749,N_28729);
xor UO_1411 (O_1411,N_28911,N_28836);
nand UO_1412 (O_1412,N_28690,N_29530);
or UO_1413 (O_1413,N_29472,N_28983);
and UO_1414 (O_1414,N_29757,N_29061);
nand UO_1415 (O_1415,N_29022,N_29058);
and UO_1416 (O_1416,N_28961,N_29511);
xor UO_1417 (O_1417,N_28943,N_28505);
nand UO_1418 (O_1418,N_29635,N_29384);
or UO_1419 (O_1419,N_28821,N_28732);
and UO_1420 (O_1420,N_29240,N_28820);
xor UO_1421 (O_1421,N_29305,N_29469);
nor UO_1422 (O_1422,N_29365,N_29636);
and UO_1423 (O_1423,N_29808,N_29229);
nand UO_1424 (O_1424,N_29888,N_29056);
nand UO_1425 (O_1425,N_29574,N_29215);
and UO_1426 (O_1426,N_29550,N_29418);
nor UO_1427 (O_1427,N_29685,N_29204);
nand UO_1428 (O_1428,N_29957,N_29906);
and UO_1429 (O_1429,N_29565,N_28623);
xor UO_1430 (O_1430,N_28531,N_29216);
xnor UO_1431 (O_1431,N_28860,N_28891);
and UO_1432 (O_1432,N_29220,N_29689);
and UO_1433 (O_1433,N_28790,N_28974);
and UO_1434 (O_1434,N_28588,N_28650);
or UO_1435 (O_1435,N_29926,N_29277);
nor UO_1436 (O_1436,N_28722,N_29163);
xor UO_1437 (O_1437,N_29995,N_29670);
or UO_1438 (O_1438,N_28790,N_29731);
and UO_1439 (O_1439,N_28652,N_28704);
nand UO_1440 (O_1440,N_29234,N_28911);
xor UO_1441 (O_1441,N_29988,N_29915);
or UO_1442 (O_1442,N_29807,N_29555);
or UO_1443 (O_1443,N_29478,N_28894);
xor UO_1444 (O_1444,N_29390,N_29473);
nand UO_1445 (O_1445,N_28636,N_29244);
or UO_1446 (O_1446,N_29044,N_29590);
or UO_1447 (O_1447,N_29964,N_28866);
nor UO_1448 (O_1448,N_29632,N_29975);
or UO_1449 (O_1449,N_29232,N_29198);
nor UO_1450 (O_1450,N_28992,N_29324);
nand UO_1451 (O_1451,N_29135,N_29025);
xnor UO_1452 (O_1452,N_29567,N_29187);
xor UO_1453 (O_1453,N_28742,N_29558);
nand UO_1454 (O_1454,N_28539,N_29638);
nand UO_1455 (O_1455,N_29181,N_29206);
or UO_1456 (O_1456,N_29161,N_28758);
xor UO_1457 (O_1457,N_29621,N_29821);
xnor UO_1458 (O_1458,N_28637,N_28794);
nand UO_1459 (O_1459,N_29095,N_28592);
and UO_1460 (O_1460,N_29598,N_29738);
nor UO_1461 (O_1461,N_28629,N_29499);
nor UO_1462 (O_1462,N_29493,N_29711);
and UO_1463 (O_1463,N_29108,N_28651);
or UO_1464 (O_1464,N_29547,N_29129);
nand UO_1465 (O_1465,N_28995,N_28684);
xnor UO_1466 (O_1466,N_29732,N_28780);
nand UO_1467 (O_1467,N_29231,N_29809);
nor UO_1468 (O_1468,N_28636,N_29609);
nor UO_1469 (O_1469,N_29672,N_29226);
and UO_1470 (O_1470,N_29078,N_29089);
nand UO_1471 (O_1471,N_29481,N_29108);
xnor UO_1472 (O_1472,N_29427,N_29677);
xor UO_1473 (O_1473,N_29497,N_28895);
xnor UO_1474 (O_1474,N_29812,N_28890);
and UO_1475 (O_1475,N_29468,N_29071);
or UO_1476 (O_1476,N_28621,N_28833);
xnor UO_1477 (O_1477,N_29989,N_29713);
and UO_1478 (O_1478,N_28824,N_28876);
and UO_1479 (O_1479,N_28910,N_29502);
or UO_1480 (O_1480,N_28724,N_29328);
nor UO_1481 (O_1481,N_28842,N_28682);
xor UO_1482 (O_1482,N_28949,N_29848);
nor UO_1483 (O_1483,N_29910,N_29361);
xor UO_1484 (O_1484,N_28916,N_29698);
xnor UO_1485 (O_1485,N_28537,N_28524);
nor UO_1486 (O_1486,N_28803,N_28950);
xnor UO_1487 (O_1487,N_28980,N_29477);
or UO_1488 (O_1488,N_29159,N_28748);
nand UO_1489 (O_1489,N_29877,N_29118);
nor UO_1490 (O_1490,N_28943,N_28767);
nand UO_1491 (O_1491,N_28861,N_29107);
and UO_1492 (O_1492,N_29797,N_28587);
and UO_1493 (O_1493,N_28841,N_29210);
nand UO_1494 (O_1494,N_29202,N_28519);
and UO_1495 (O_1495,N_28681,N_29533);
xnor UO_1496 (O_1496,N_29928,N_28761);
nor UO_1497 (O_1497,N_29483,N_29187);
and UO_1498 (O_1498,N_29444,N_28856);
nand UO_1499 (O_1499,N_29711,N_29758);
or UO_1500 (O_1500,N_29446,N_28955);
xor UO_1501 (O_1501,N_29303,N_29651);
nand UO_1502 (O_1502,N_29338,N_29012);
nor UO_1503 (O_1503,N_29734,N_29081);
and UO_1504 (O_1504,N_29648,N_29658);
xnor UO_1505 (O_1505,N_29589,N_29792);
xor UO_1506 (O_1506,N_28638,N_29171);
nor UO_1507 (O_1507,N_28774,N_29287);
nor UO_1508 (O_1508,N_28907,N_29406);
and UO_1509 (O_1509,N_29221,N_28990);
and UO_1510 (O_1510,N_28512,N_29271);
or UO_1511 (O_1511,N_29120,N_29709);
nor UO_1512 (O_1512,N_28991,N_28909);
or UO_1513 (O_1513,N_29622,N_29442);
nor UO_1514 (O_1514,N_29269,N_28700);
nand UO_1515 (O_1515,N_28605,N_28901);
xnor UO_1516 (O_1516,N_29901,N_28973);
nand UO_1517 (O_1517,N_29527,N_29217);
or UO_1518 (O_1518,N_28993,N_28645);
xnor UO_1519 (O_1519,N_29954,N_29847);
nor UO_1520 (O_1520,N_29572,N_29665);
nand UO_1521 (O_1521,N_28582,N_28798);
and UO_1522 (O_1522,N_28692,N_28548);
nand UO_1523 (O_1523,N_29738,N_29712);
and UO_1524 (O_1524,N_29243,N_28994);
nand UO_1525 (O_1525,N_28962,N_29118);
nand UO_1526 (O_1526,N_29457,N_29380);
nand UO_1527 (O_1527,N_29635,N_29126);
or UO_1528 (O_1528,N_28864,N_29317);
nand UO_1529 (O_1529,N_29655,N_29342);
and UO_1530 (O_1530,N_28524,N_28831);
nand UO_1531 (O_1531,N_29208,N_28715);
and UO_1532 (O_1532,N_29625,N_28578);
and UO_1533 (O_1533,N_28643,N_29079);
nand UO_1534 (O_1534,N_29790,N_29883);
xor UO_1535 (O_1535,N_29387,N_29188);
or UO_1536 (O_1536,N_29974,N_29952);
xor UO_1537 (O_1537,N_29256,N_29933);
xor UO_1538 (O_1538,N_28812,N_28992);
xnor UO_1539 (O_1539,N_29991,N_29234);
or UO_1540 (O_1540,N_29426,N_29436);
xor UO_1541 (O_1541,N_28509,N_28582);
or UO_1542 (O_1542,N_29605,N_29099);
and UO_1543 (O_1543,N_29732,N_29662);
nor UO_1544 (O_1544,N_28840,N_29304);
and UO_1545 (O_1545,N_29510,N_29264);
and UO_1546 (O_1546,N_29223,N_29960);
xor UO_1547 (O_1547,N_28936,N_29533);
nor UO_1548 (O_1548,N_28942,N_28727);
nor UO_1549 (O_1549,N_29795,N_29680);
xnor UO_1550 (O_1550,N_29028,N_29628);
or UO_1551 (O_1551,N_29467,N_28735);
and UO_1552 (O_1552,N_29637,N_28802);
and UO_1553 (O_1553,N_29707,N_29123);
nand UO_1554 (O_1554,N_29772,N_29576);
nand UO_1555 (O_1555,N_29449,N_29995);
nor UO_1556 (O_1556,N_29502,N_28859);
and UO_1557 (O_1557,N_28919,N_29388);
and UO_1558 (O_1558,N_29017,N_28611);
nand UO_1559 (O_1559,N_28708,N_29136);
nand UO_1560 (O_1560,N_29828,N_29536);
and UO_1561 (O_1561,N_28984,N_29623);
xnor UO_1562 (O_1562,N_28581,N_28626);
or UO_1563 (O_1563,N_29296,N_29167);
nand UO_1564 (O_1564,N_29873,N_28878);
nor UO_1565 (O_1565,N_29979,N_29346);
and UO_1566 (O_1566,N_28996,N_28929);
nand UO_1567 (O_1567,N_29552,N_28850);
and UO_1568 (O_1568,N_28574,N_28667);
and UO_1569 (O_1569,N_28683,N_29382);
nor UO_1570 (O_1570,N_29332,N_29446);
or UO_1571 (O_1571,N_29472,N_29951);
nand UO_1572 (O_1572,N_29516,N_28664);
xor UO_1573 (O_1573,N_29202,N_29975);
or UO_1574 (O_1574,N_29337,N_29384);
xor UO_1575 (O_1575,N_29714,N_29364);
nand UO_1576 (O_1576,N_29239,N_28654);
and UO_1577 (O_1577,N_29445,N_28679);
nor UO_1578 (O_1578,N_28691,N_28699);
nor UO_1579 (O_1579,N_28978,N_28708);
or UO_1580 (O_1580,N_29891,N_29244);
and UO_1581 (O_1581,N_29599,N_29000);
nand UO_1582 (O_1582,N_28901,N_28877);
xnor UO_1583 (O_1583,N_29432,N_28805);
or UO_1584 (O_1584,N_28928,N_29068);
nor UO_1585 (O_1585,N_29842,N_29599);
nor UO_1586 (O_1586,N_28720,N_29963);
nor UO_1587 (O_1587,N_29628,N_28554);
nand UO_1588 (O_1588,N_28887,N_29925);
and UO_1589 (O_1589,N_28808,N_29447);
and UO_1590 (O_1590,N_29957,N_29266);
nand UO_1591 (O_1591,N_28798,N_29639);
nor UO_1592 (O_1592,N_29972,N_29214);
nor UO_1593 (O_1593,N_28815,N_29268);
and UO_1594 (O_1594,N_28601,N_29342);
and UO_1595 (O_1595,N_28744,N_28663);
nor UO_1596 (O_1596,N_29284,N_28850);
and UO_1597 (O_1597,N_28624,N_29925);
nand UO_1598 (O_1598,N_29140,N_29317);
xnor UO_1599 (O_1599,N_29535,N_29706);
xnor UO_1600 (O_1600,N_29084,N_29465);
nor UO_1601 (O_1601,N_29733,N_29902);
or UO_1602 (O_1602,N_29618,N_29138);
and UO_1603 (O_1603,N_29594,N_28610);
nand UO_1604 (O_1604,N_29655,N_29137);
or UO_1605 (O_1605,N_29952,N_28902);
nor UO_1606 (O_1606,N_29008,N_29344);
or UO_1607 (O_1607,N_28656,N_29049);
nand UO_1608 (O_1608,N_29152,N_29541);
and UO_1609 (O_1609,N_29903,N_29389);
nor UO_1610 (O_1610,N_29788,N_29613);
nor UO_1611 (O_1611,N_29489,N_29477);
nor UO_1612 (O_1612,N_28790,N_29550);
or UO_1613 (O_1613,N_29262,N_29430);
nand UO_1614 (O_1614,N_29288,N_28849);
xor UO_1615 (O_1615,N_29709,N_29126);
nand UO_1616 (O_1616,N_29932,N_28864);
nand UO_1617 (O_1617,N_29871,N_29297);
xor UO_1618 (O_1618,N_29442,N_28779);
nor UO_1619 (O_1619,N_29507,N_28994);
xnor UO_1620 (O_1620,N_29563,N_28595);
and UO_1621 (O_1621,N_29887,N_29085);
xnor UO_1622 (O_1622,N_28838,N_28563);
xnor UO_1623 (O_1623,N_28816,N_28791);
xor UO_1624 (O_1624,N_28823,N_29123);
nand UO_1625 (O_1625,N_28549,N_29677);
and UO_1626 (O_1626,N_28559,N_29971);
nand UO_1627 (O_1627,N_29164,N_29195);
xnor UO_1628 (O_1628,N_29576,N_29377);
xor UO_1629 (O_1629,N_29202,N_29914);
or UO_1630 (O_1630,N_29201,N_29596);
xor UO_1631 (O_1631,N_29276,N_29713);
and UO_1632 (O_1632,N_28782,N_29794);
or UO_1633 (O_1633,N_29939,N_29500);
or UO_1634 (O_1634,N_28606,N_29395);
or UO_1635 (O_1635,N_28890,N_28698);
nor UO_1636 (O_1636,N_29122,N_29591);
and UO_1637 (O_1637,N_29565,N_28641);
or UO_1638 (O_1638,N_28821,N_29431);
and UO_1639 (O_1639,N_29094,N_29698);
or UO_1640 (O_1640,N_28877,N_29721);
or UO_1641 (O_1641,N_29670,N_29379);
or UO_1642 (O_1642,N_29968,N_28960);
nor UO_1643 (O_1643,N_28930,N_28935);
nand UO_1644 (O_1644,N_29023,N_29736);
nand UO_1645 (O_1645,N_28577,N_29391);
or UO_1646 (O_1646,N_29297,N_29973);
and UO_1647 (O_1647,N_29069,N_29757);
nor UO_1648 (O_1648,N_29902,N_29337);
nand UO_1649 (O_1649,N_28929,N_29902);
or UO_1650 (O_1650,N_29056,N_29533);
and UO_1651 (O_1651,N_29013,N_29286);
or UO_1652 (O_1652,N_28922,N_29969);
and UO_1653 (O_1653,N_29916,N_28691);
nand UO_1654 (O_1654,N_29610,N_29625);
or UO_1655 (O_1655,N_29456,N_29721);
nor UO_1656 (O_1656,N_29530,N_29766);
or UO_1657 (O_1657,N_28829,N_29324);
xnor UO_1658 (O_1658,N_29677,N_29132);
nor UO_1659 (O_1659,N_28548,N_28843);
xnor UO_1660 (O_1660,N_28515,N_29821);
or UO_1661 (O_1661,N_28548,N_28902);
nor UO_1662 (O_1662,N_29258,N_28829);
nor UO_1663 (O_1663,N_29683,N_28676);
nor UO_1664 (O_1664,N_29215,N_29936);
nor UO_1665 (O_1665,N_29690,N_29829);
or UO_1666 (O_1666,N_29539,N_29759);
xor UO_1667 (O_1667,N_29032,N_28955);
xor UO_1668 (O_1668,N_29802,N_29297);
or UO_1669 (O_1669,N_29095,N_28994);
xnor UO_1670 (O_1670,N_29911,N_28970);
or UO_1671 (O_1671,N_29938,N_28793);
nor UO_1672 (O_1672,N_28562,N_29392);
xnor UO_1673 (O_1673,N_28664,N_29907);
and UO_1674 (O_1674,N_29485,N_29076);
nor UO_1675 (O_1675,N_29333,N_29443);
nor UO_1676 (O_1676,N_29021,N_28770);
nor UO_1677 (O_1677,N_29280,N_29597);
or UO_1678 (O_1678,N_28648,N_29450);
nand UO_1679 (O_1679,N_29783,N_29411);
nand UO_1680 (O_1680,N_29193,N_28981);
xnor UO_1681 (O_1681,N_28897,N_29860);
xor UO_1682 (O_1682,N_29482,N_29101);
or UO_1683 (O_1683,N_29416,N_29719);
xnor UO_1684 (O_1684,N_29290,N_29462);
nor UO_1685 (O_1685,N_29784,N_29395);
nand UO_1686 (O_1686,N_29216,N_29517);
nor UO_1687 (O_1687,N_29109,N_28736);
and UO_1688 (O_1688,N_29874,N_29379);
nor UO_1689 (O_1689,N_29765,N_28705);
xnor UO_1690 (O_1690,N_29449,N_29922);
and UO_1691 (O_1691,N_29414,N_28590);
nor UO_1692 (O_1692,N_28594,N_29902);
and UO_1693 (O_1693,N_29923,N_29566);
nand UO_1694 (O_1694,N_28822,N_29442);
xor UO_1695 (O_1695,N_28793,N_29354);
xor UO_1696 (O_1696,N_29616,N_28770);
nand UO_1697 (O_1697,N_28867,N_29947);
and UO_1698 (O_1698,N_28636,N_29728);
or UO_1699 (O_1699,N_29729,N_29311);
nand UO_1700 (O_1700,N_28888,N_29095);
or UO_1701 (O_1701,N_29020,N_29901);
and UO_1702 (O_1702,N_28746,N_29726);
nor UO_1703 (O_1703,N_28966,N_28586);
nand UO_1704 (O_1704,N_28791,N_29808);
xor UO_1705 (O_1705,N_29595,N_28975);
and UO_1706 (O_1706,N_29824,N_28943);
nor UO_1707 (O_1707,N_29471,N_29691);
xnor UO_1708 (O_1708,N_28857,N_29432);
or UO_1709 (O_1709,N_28709,N_29874);
xor UO_1710 (O_1710,N_28515,N_28826);
nand UO_1711 (O_1711,N_29306,N_28867);
nand UO_1712 (O_1712,N_29347,N_29084);
nor UO_1713 (O_1713,N_29397,N_28985);
nor UO_1714 (O_1714,N_28939,N_29963);
or UO_1715 (O_1715,N_29464,N_29555);
or UO_1716 (O_1716,N_29965,N_28686);
and UO_1717 (O_1717,N_29136,N_28685);
or UO_1718 (O_1718,N_29386,N_29299);
and UO_1719 (O_1719,N_28950,N_29872);
nand UO_1720 (O_1720,N_29186,N_28775);
and UO_1721 (O_1721,N_28923,N_29205);
nor UO_1722 (O_1722,N_29360,N_29555);
nor UO_1723 (O_1723,N_29132,N_29293);
nor UO_1724 (O_1724,N_29990,N_28820);
nor UO_1725 (O_1725,N_28812,N_29784);
nand UO_1726 (O_1726,N_28721,N_28814);
xnor UO_1727 (O_1727,N_29914,N_29949);
nand UO_1728 (O_1728,N_29426,N_29594);
xnor UO_1729 (O_1729,N_29203,N_28896);
nand UO_1730 (O_1730,N_29755,N_28995);
and UO_1731 (O_1731,N_29655,N_29886);
or UO_1732 (O_1732,N_29510,N_28891);
and UO_1733 (O_1733,N_29102,N_28647);
and UO_1734 (O_1734,N_29393,N_29290);
and UO_1735 (O_1735,N_29133,N_29641);
xnor UO_1736 (O_1736,N_29900,N_28546);
or UO_1737 (O_1737,N_29610,N_28992);
nand UO_1738 (O_1738,N_29348,N_29964);
xnor UO_1739 (O_1739,N_29929,N_28549);
xnor UO_1740 (O_1740,N_29546,N_29101);
nor UO_1741 (O_1741,N_29133,N_29501);
nor UO_1742 (O_1742,N_28700,N_28594);
or UO_1743 (O_1743,N_28743,N_29955);
xnor UO_1744 (O_1744,N_29906,N_29336);
and UO_1745 (O_1745,N_28918,N_28602);
xnor UO_1746 (O_1746,N_28542,N_28673);
and UO_1747 (O_1747,N_29733,N_28577);
nand UO_1748 (O_1748,N_29349,N_28531);
or UO_1749 (O_1749,N_28676,N_29204);
or UO_1750 (O_1750,N_28833,N_28946);
or UO_1751 (O_1751,N_28551,N_28570);
and UO_1752 (O_1752,N_28968,N_29323);
nor UO_1753 (O_1753,N_28810,N_28998);
and UO_1754 (O_1754,N_29331,N_29085);
nand UO_1755 (O_1755,N_29181,N_29835);
nand UO_1756 (O_1756,N_28826,N_29536);
nor UO_1757 (O_1757,N_29032,N_29017);
or UO_1758 (O_1758,N_29938,N_29220);
and UO_1759 (O_1759,N_29417,N_29047);
nand UO_1760 (O_1760,N_29505,N_29661);
xnor UO_1761 (O_1761,N_29838,N_29950);
and UO_1762 (O_1762,N_29974,N_29170);
or UO_1763 (O_1763,N_29378,N_29070);
xnor UO_1764 (O_1764,N_29266,N_29337);
or UO_1765 (O_1765,N_29190,N_29138);
xnor UO_1766 (O_1766,N_28584,N_29055);
nand UO_1767 (O_1767,N_29712,N_28602);
or UO_1768 (O_1768,N_29137,N_29247);
and UO_1769 (O_1769,N_29538,N_28530);
nand UO_1770 (O_1770,N_29244,N_28918);
xor UO_1771 (O_1771,N_29519,N_28701);
nor UO_1772 (O_1772,N_28967,N_28932);
or UO_1773 (O_1773,N_29742,N_29901);
nor UO_1774 (O_1774,N_28955,N_29642);
and UO_1775 (O_1775,N_29129,N_28651);
xor UO_1776 (O_1776,N_28869,N_28704);
nor UO_1777 (O_1777,N_29032,N_29849);
or UO_1778 (O_1778,N_28618,N_29362);
and UO_1779 (O_1779,N_29411,N_28744);
and UO_1780 (O_1780,N_28600,N_29393);
xnor UO_1781 (O_1781,N_29440,N_29937);
nor UO_1782 (O_1782,N_29357,N_29541);
or UO_1783 (O_1783,N_29879,N_29671);
nor UO_1784 (O_1784,N_28634,N_28910);
and UO_1785 (O_1785,N_29867,N_28952);
or UO_1786 (O_1786,N_29928,N_29896);
and UO_1787 (O_1787,N_29915,N_29116);
or UO_1788 (O_1788,N_29883,N_28903);
xnor UO_1789 (O_1789,N_29513,N_28746);
and UO_1790 (O_1790,N_29958,N_28583);
and UO_1791 (O_1791,N_29592,N_29801);
or UO_1792 (O_1792,N_28529,N_29514);
and UO_1793 (O_1793,N_28720,N_29014);
and UO_1794 (O_1794,N_29364,N_29580);
nor UO_1795 (O_1795,N_29658,N_29952);
nand UO_1796 (O_1796,N_28564,N_28812);
or UO_1797 (O_1797,N_29980,N_29548);
nand UO_1798 (O_1798,N_28677,N_29808);
or UO_1799 (O_1799,N_29960,N_29853);
and UO_1800 (O_1800,N_28555,N_29823);
or UO_1801 (O_1801,N_28993,N_29842);
nand UO_1802 (O_1802,N_29351,N_28772);
and UO_1803 (O_1803,N_29075,N_29407);
and UO_1804 (O_1804,N_29968,N_29106);
or UO_1805 (O_1805,N_28824,N_29834);
xnor UO_1806 (O_1806,N_29913,N_29506);
xor UO_1807 (O_1807,N_29639,N_29864);
xnor UO_1808 (O_1808,N_28620,N_29106);
xnor UO_1809 (O_1809,N_29004,N_29017);
nand UO_1810 (O_1810,N_29925,N_29765);
xnor UO_1811 (O_1811,N_29565,N_29854);
or UO_1812 (O_1812,N_28584,N_28895);
xor UO_1813 (O_1813,N_29462,N_29955);
xor UO_1814 (O_1814,N_29376,N_29890);
or UO_1815 (O_1815,N_29143,N_29183);
nand UO_1816 (O_1816,N_29888,N_29373);
nor UO_1817 (O_1817,N_29685,N_29849);
and UO_1818 (O_1818,N_29080,N_29485);
xor UO_1819 (O_1819,N_29233,N_29134);
or UO_1820 (O_1820,N_29308,N_29746);
and UO_1821 (O_1821,N_29468,N_28551);
and UO_1822 (O_1822,N_29985,N_29612);
or UO_1823 (O_1823,N_28792,N_29203);
or UO_1824 (O_1824,N_29102,N_29643);
nand UO_1825 (O_1825,N_28972,N_28889);
nand UO_1826 (O_1826,N_28897,N_29045);
nand UO_1827 (O_1827,N_29755,N_29201);
or UO_1828 (O_1828,N_28953,N_29563);
xnor UO_1829 (O_1829,N_28563,N_29634);
nor UO_1830 (O_1830,N_29950,N_29573);
nand UO_1831 (O_1831,N_29910,N_29305);
and UO_1832 (O_1832,N_29714,N_29522);
or UO_1833 (O_1833,N_29118,N_29984);
xnor UO_1834 (O_1834,N_29647,N_29272);
nor UO_1835 (O_1835,N_28511,N_28845);
and UO_1836 (O_1836,N_28676,N_28535);
xor UO_1837 (O_1837,N_29383,N_28549);
nand UO_1838 (O_1838,N_29774,N_29677);
nor UO_1839 (O_1839,N_28638,N_29699);
or UO_1840 (O_1840,N_28773,N_29683);
nand UO_1841 (O_1841,N_29631,N_29683);
nor UO_1842 (O_1842,N_28795,N_29259);
and UO_1843 (O_1843,N_29810,N_29544);
and UO_1844 (O_1844,N_29441,N_29267);
nor UO_1845 (O_1845,N_29164,N_29792);
xor UO_1846 (O_1846,N_29919,N_29351);
xor UO_1847 (O_1847,N_28607,N_29202);
or UO_1848 (O_1848,N_29932,N_29523);
nand UO_1849 (O_1849,N_29265,N_29774);
nor UO_1850 (O_1850,N_28897,N_29008);
or UO_1851 (O_1851,N_29497,N_29510);
or UO_1852 (O_1852,N_28599,N_29751);
and UO_1853 (O_1853,N_28850,N_29336);
and UO_1854 (O_1854,N_29149,N_29283);
xnor UO_1855 (O_1855,N_28751,N_29491);
nor UO_1856 (O_1856,N_29308,N_29809);
or UO_1857 (O_1857,N_28769,N_29017);
and UO_1858 (O_1858,N_28666,N_29375);
nand UO_1859 (O_1859,N_28922,N_29487);
nor UO_1860 (O_1860,N_29079,N_29976);
or UO_1861 (O_1861,N_29651,N_28614);
nand UO_1862 (O_1862,N_29434,N_29303);
nand UO_1863 (O_1863,N_29389,N_29437);
xnor UO_1864 (O_1864,N_29131,N_29013);
nor UO_1865 (O_1865,N_28621,N_29420);
xor UO_1866 (O_1866,N_29536,N_28915);
and UO_1867 (O_1867,N_29274,N_28617);
xor UO_1868 (O_1868,N_29678,N_28576);
nor UO_1869 (O_1869,N_29341,N_28663);
and UO_1870 (O_1870,N_29259,N_29959);
or UO_1871 (O_1871,N_29236,N_28558);
and UO_1872 (O_1872,N_29907,N_29313);
or UO_1873 (O_1873,N_28572,N_28769);
and UO_1874 (O_1874,N_29482,N_29471);
nand UO_1875 (O_1875,N_28977,N_29914);
nand UO_1876 (O_1876,N_28622,N_29171);
nor UO_1877 (O_1877,N_28608,N_29387);
nand UO_1878 (O_1878,N_29366,N_29491);
xnor UO_1879 (O_1879,N_29722,N_29872);
xor UO_1880 (O_1880,N_29695,N_29263);
nand UO_1881 (O_1881,N_28931,N_29345);
xor UO_1882 (O_1882,N_29538,N_29074);
and UO_1883 (O_1883,N_28594,N_28751);
xor UO_1884 (O_1884,N_29658,N_29705);
or UO_1885 (O_1885,N_28661,N_29231);
and UO_1886 (O_1886,N_29986,N_29724);
and UO_1887 (O_1887,N_29917,N_29450);
nor UO_1888 (O_1888,N_28533,N_28851);
and UO_1889 (O_1889,N_28595,N_29527);
nor UO_1890 (O_1890,N_29488,N_29195);
xnor UO_1891 (O_1891,N_29237,N_29735);
nor UO_1892 (O_1892,N_29082,N_28939);
and UO_1893 (O_1893,N_29691,N_28810);
nor UO_1894 (O_1894,N_28956,N_29190);
nor UO_1895 (O_1895,N_28917,N_28612);
xnor UO_1896 (O_1896,N_29532,N_29192);
xnor UO_1897 (O_1897,N_29969,N_29874);
nand UO_1898 (O_1898,N_29930,N_29170);
nand UO_1899 (O_1899,N_28992,N_29801);
nor UO_1900 (O_1900,N_29399,N_28640);
or UO_1901 (O_1901,N_29420,N_29919);
or UO_1902 (O_1902,N_28873,N_28553);
and UO_1903 (O_1903,N_28738,N_29095);
xor UO_1904 (O_1904,N_29560,N_28794);
xor UO_1905 (O_1905,N_29432,N_28664);
nor UO_1906 (O_1906,N_29496,N_29745);
and UO_1907 (O_1907,N_29864,N_29279);
nand UO_1908 (O_1908,N_29546,N_29096);
nand UO_1909 (O_1909,N_29409,N_29649);
and UO_1910 (O_1910,N_29471,N_28504);
nor UO_1911 (O_1911,N_28843,N_29165);
and UO_1912 (O_1912,N_28820,N_28730);
or UO_1913 (O_1913,N_29433,N_29754);
and UO_1914 (O_1914,N_29292,N_29803);
or UO_1915 (O_1915,N_29496,N_29343);
or UO_1916 (O_1916,N_29722,N_29030);
or UO_1917 (O_1917,N_29484,N_29668);
nor UO_1918 (O_1918,N_29697,N_29309);
nand UO_1919 (O_1919,N_28637,N_29483);
nand UO_1920 (O_1920,N_29958,N_29767);
xnor UO_1921 (O_1921,N_29389,N_28805);
and UO_1922 (O_1922,N_28503,N_28729);
nor UO_1923 (O_1923,N_28636,N_29347);
and UO_1924 (O_1924,N_29264,N_28621);
nor UO_1925 (O_1925,N_29432,N_28677);
xnor UO_1926 (O_1926,N_29645,N_29551);
nand UO_1927 (O_1927,N_28954,N_28743);
nor UO_1928 (O_1928,N_29353,N_28747);
xor UO_1929 (O_1929,N_29499,N_28773);
and UO_1930 (O_1930,N_29389,N_29964);
xor UO_1931 (O_1931,N_29892,N_29632);
nand UO_1932 (O_1932,N_28808,N_28602);
nor UO_1933 (O_1933,N_28973,N_28878);
nor UO_1934 (O_1934,N_28933,N_28545);
nand UO_1935 (O_1935,N_28725,N_29860);
or UO_1936 (O_1936,N_29237,N_29289);
and UO_1937 (O_1937,N_28878,N_29922);
xnor UO_1938 (O_1938,N_29675,N_29790);
or UO_1939 (O_1939,N_29199,N_28638);
and UO_1940 (O_1940,N_28935,N_28634);
nor UO_1941 (O_1941,N_29509,N_28800);
nand UO_1942 (O_1942,N_29428,N_29072);
and UO_1943 (O_1943,N_29947,N_29041);
xnor UO_1944 (O_1944,N_28936,N_28878);
nand UO_1945 (O_1945,N_29408,N_29397);
or UO_1946 (O_1946,N_29667,N_29062);
and UO_1947 (O_1947,N_28642,N_29417);
or UO_1948 (O_1948,N_29523,N_29056);
and UO_1949 (O_1949,N_29206,N_29267);
nand UO_1950 (O_1950,N_28791,N_29935);
nand UO_1951 (O_1951,N_29438,N_29279);
nor UO_1952 (O_1952,N_28946,N_29224);
nand UO_1953 (O_1953,N_28710,N_29292);
xnor UO_1954 (O_1954,N_29917,N_28782);
nor UO_1955 (O_1955,N_29756,N_29163);
xnor UO_1956 (O_1956,N_29538,N_29715);
and UO_1957 (O_1957,N_28769,N_29514);
nor UO_1958 (O_1958,N_28583,N_29922);
nand UO_1959 (O_1959,N_29696,N_28524);
and UO_1960 (O_1960,N_29046,N_28705);
xor UO_1961 (O_1961,N_29196,N_29661);
or UO_1962 (O_1962,N_28874,N_29927);
nor UO_1963 (O_1963,N_28501,N_28585);
nand UO_1964 (O_1964,N_29312,N_29757);
xor UO_1965 (O_1965,N_29607,N_28745);
and UO_1966 (O_1966,N_29319,N_29574);
or UO_1967 (O_1967,N_29104,N_29541);
nand UO_1968 (O_1968,N_28648,N_29702);
and UO_1969 (O_1969,N_28577,N_28870);
and UO_1970 (O_1970,N_29838,N_29249);
nand UO_1971 (O_1971,N_28852,N_29933);
and UO_1972 (O_1972,N_29442,N_29523);
or UO_1973 (O_1973,N_29790,N_28818);
and UO_1974 (O_1974,N_29638,N_29507);
or UO_1975 (O_1975,N_29752,N_28786);
or UO_1976 (O_1976,N_29434,N_29922);
nand UO_1977 (O_1977,N_29900,N_28611);
nand UO_1978 (O_1978,N_29830,N_29222);
nor UO_1979 (O_1979,N_29069,N_28613);
and UO_1980 (O_1980,N_29245,N_28758);
nor UO_1981 (O_1981,N_28708,N_29340);
and UO_1982 (O_1982,N_29676,N_29231);
xnor UO_1983 (O_1983,N_29679,N_29758);
and UO_1984 (O_1984,N_29168,N_29674);
nand UO_1985 (O_1985,N_29618,N_29773);
nor UO_1986 (O_1986,N_29614,N_28547);
and UO_1987 (O_1987,N_29329,N_28641);
and UO_1988 (O_1988,N_29613,N_29870);
nand UO_1989 (O_1989,N_29070,N_28863);
or UO_1990 (O_1990,N_29565,N_29138);
nand UO_1991 (O_1991,N_29292,N_28678);
nor UO_1992 (O_1992,N_28512,N_29194);
nor UO_1993 (O_1993,N_28929,N_29886);
or UO_1994 (O_1994,N_29021,N_28872);
xnor UO_1995 (O_1995,N_29382,N_29851);
nand UO_1996 (O_1996,N_29806,N_28543);
and UO_1997 (O_1997,N_28881,N_29400);
or UO_1998 (O_1998,N_29126,N_28536);
xor UO_1999 (O_1999,N_29391,N_28860);
nor UO_2000 (O_2000,N_29364,N_29826);
and UO_2001 (O_2001,N_29649,N_29994);
and UO_2002 (O_2002,N_29924,N_28827);
or UO_2003 (O_2003,N_29631,N_29196);
nor UO_2004 (O_2004,N_29972,N_28663);
and UO_2005 (O_2005,N_29356,N_29116);
nor UO_2006 (O_2006,N_28512,N_28563);
and UO_2007 (O_2007,N_28822,N_29155);
xnor UO_2008 (O_2008,N_29517,N_28741);
nand UO_2009 (O_2009,N_29373,N_28715);
or UO_2010 (O_2010,N_29154,N_29584);
or UO_2011 (O_2011,N_28929,N_29887);
nand UO_2012 (O_2012,N_29829,N_29055);
nand UO_2013 (O_2013,N_29845,N_28534);
or UO_2014 (O_2014,N_28797,N_29594);
xnor UO_2015 (O_2015,N_28761,N_28746);
nor UO_2016 (O_2016,N_28644,N_29934);
and UO_2017 (O_2017,N_28543,N_28849);
xnor UO_2018 (O_2018,N_29956,N_28787);
xor UO_2019 (O_2019,N_29585,N_29521);
and UO_2020 (O_2020,N_28782,N_28617);
and UO_2021 (O_2021,N_29529,N_28869);
nand UO_2022 (O_2022,N_28661,N_29505);
xnor UO_2023 (O_2023,N_29270,N_28608);
nor UO_2024 (O_2024,N_29144,N_28693);
nor UO_2025 (O_2025,N_29909,N_29124);
or UO_2026 (O_2026,N_28949,N_28957);
xnor UO_2027 (O_2027,N_28575,N_28972);
or UO_2028 (O_2028,N_29606,N_28915);
and UO_2029 (O_2029,N_29180,N_28695);
nor UO_2030 (O_2030,N_29351,N_29253);
nand UO_2031 (O_2031,N_28762,N_29339);
nand UO_2032 (O_2032,N_29750,N_28623);
or UO_2033 (O_2033,N_28957,N_29244);
or UO_2034 (O_2034,N_28813,N_28952);
nor UO_2035 (O_2035,N_29865,N_28671);
xor UO_2036 (O_2036,N_29221,N_29977);
xor UO_2037 (O_2037,N_28786,N_28890);
xor UO_2038 (O_2038,N_28973,N_29791);
and UO_2039 (O_2039,N_29238,N_29474);
or UO_2040 (O_2040,N_29347,N_29428);
xor UO_2041 (O_2041,N_29839,N_29656);
nand UO_2042 (O_2042,N_29458,N_29522);
and UO_2043 (O_2043,N_29234,N_29000);
or UO_2044 (O_2044,N_29355,N_29120);
and UO_2045 (O_2045,N_29516,N_29372);
or UO_2046 (O_2046,N_29664,N_28673);
and UO_2047 (O_2047,N_29762,N_29927);
or UO_2048 (O_2048,N_28507,N_29048);
and UO_2049 (O_2049,N_29687,N_29763);
nor UO_2050 (O_2050,N_29542,N_28746);
nor UO_2051 (O_2051,N_29818,N_29657);
nor UO_2052 (O_2052,N_29899,N_29354);
nand UO_2053 (O_2053,N_29057,N_29352);
xnor UO_2054 (O_2054,N_28791,N_29894);
nor UO_2055 (O_2055,N_28805,N_28903);
and UO_2056 (O_2056,N_29985,N_28552);
xnor UO_2057 (O_2057,N_29702,N_29248);
nor UO_2058 (O_2058,N_29786,N_29348);
and UO_2059 (O_2059,N_29725,N_28742);
nand UO_2060 (O_2060,N_29438,N_29110);
xor UO_2061 (O_2061,N_28511,N_29363);
and UO_2062 (O_2062,N_29823,N_29082);
nand UO_2063 (O_2063,N_28535,N_28903);
nor UO_2064 (O_2064,N_29100,N_29075);
and UO_2065 (O_2065,N_29711,N_28823);
nor UO_2066 (O_2066,N_29480,N_29669);
nand UO_2067 (O_2067,N_28712,N_29659);
and UO_2068 (O_2068,N_29978,N_29191);
nand UO_2069 (O_2069,N_28726,N_29333);
nand UO_2070 (O_2070,N_28508,N_29184);
or UO_2071 (O_2071,N_28971,N_28999);
or UO_2072 (O_2072,N_28535,N_29722);
or UO_2073 (O_2073,N_28674,N_28570);
xnor UO_2074 (O_2074,N_29061,N_29729);
and UO_2075 (O_2075,N_29045,N_29437);
nor UO_2076 (O_2076,N_29451,N_28725);
xor UO_2077 (O_2077,N_29153,N_28962);
nor UO_2078 (O_2078,N_29771,N_29161);
nand UO_2079 (O_2079,N_28649,N_28745);
or UO_2080 (O_2080,N_28837,N_28846);
or UO_2081 (O_2081,N_29615,N_28681);
and UO_2082 (O_2082,N_29973,N_29272);
or UO_2083 (O_2083,N_28570,N_29828);
or UO_2084 (O_2084,N_29778,N_29858);
nor UO_2085 (O_2085,N_29491,N_29658);
or UO_2086 (O_2086,N_29195,N_29823);
nand UO_2087 (O_2087,N_28811,N_28524);
xnor UO_2088 (O_2088,N_29912,N_28619);
or UO_2089 (O_2089,N_29829,N_28661);
or UO_2090 (O_2090,N_29431,N_29727);
nor UO_2091 (O_2091,N_28597,N_29448);
or UO_2092 (O_2092,N_29349,N_29586);
nand UO_2093 (O_2093,N_29709,N_29029);
or UO_2094 (O_2094,N_28580,N_29457);
xor UO_2095 (O_2095,N_29438,N_29193);
nor UO_2096 (O_2096,N_29805,N_29432);
or UO_2097 (O_2097,N_29625,N_28654);
and UO_2098 (O_2098,N_28506,N_29992);
nand UO_2099 (O_2099,N_28965,N_28939);
nor UO_2100 (O_2100,N_28793,N_29910);
nor UO_2101 (O_2101,N_29302,N_29357);
nor UO_2102 (O_2102,N_29760,N_29667);
nor UO_2103 (O_2103,N_29913,N_29183);
nand UO_2104 (O_2104,N_29745,N_29683);
or UO_2105 (O_2105,N_28830,N_29402);
or UO_2106 (O_2106,N_29317,N_29702);
or UO_2107 (O_2107,N_28611,N_29569);
nor UO_2108 (O_2108,N_28673,N_28751);
nand UO_2109 (O_2109,N_29192,N_29230);
or UO_2110 (O_2110,N_28900,N_28989);
or UO_2111 (O_2111,N_29013,N_29519);
nand UO_2112 (O_2112,N_29245,N_29875);
and UO_2113 (O_2113,N_29673,N_29714);
or UO_2114 (O_2114,N_29686,N_29914);
xnor UO_2115 (O_2115,N_29723,N_29569);
nand UO_2116 (O_2116,N_29107,N_29798);
nand UO_2117 (O_2117,N_29175,N_29865);
nand UO_2118 (O_2118,N_28679,N_29395);
or UO_2119 (O_2119,N_29359,N_28852);
xor UO_2120 (O_2120,N_29814,N_28932);
nand UO_2121 (O_2121,N_29063,N_29770);
nor UO_2122 (O_2122,N_29646,N_28785);
nor UO_2123 (O_2123,N_29800,N_28628);
xor UO_2124 (O_2124,N_28611,N_29911);
or UO_2125 (O_2125,N_28717,N_29838);
nor UO_2126 (O_2126,N_28954,N_28769);
and UO_2127 (O_2127,N_29665,N_28965);
nand UO_2128 (O_2128,N_28706,N_29403);
xnor UO_2129 (O_2129,N_29169,N_28560);
nor UO_2130 (O_2130,N_29960,N_28894);
xnor UO_2131 (O_2131,N_29914,N_28657);
xnor UO_2132 (O_2132,N_29302,N_29470);
nor UO_2133 (O_2133,N_29646,N_29149);
nor UO_2134 (O_2134,N_28540,N_28883);
nand UO_2135 (O_2135,N_28665,N_29229);
nor UO_2136 (O_2136,N_29925,N_29184);
nor UO_2137 (O_2137,N_29041,N_29612);
nand UO_2138 (O_2138,N_29836,N_29295);
or UO_2139 (O_2139,N_29232,N_28988);
xor UO_2140 (O_2140,N_29635,N_29849);
and UO_2141 (O_2141,N_28933,N_29477);
xor UO_2142 (O_2142,N_29742,N_28537);
and UO_2143 (O_2143,N_29243,N_29827);
or UO_2144 (O_2144,N_29917,N_29368);
or UO_2145 (O_2145,N_29518,N_29220);
or UO_2146 (O_2146,N_28544,N_28996);
nand UO_2147 (O_2147,N_29803,N_28799);
xnor UO_2148 (O_2148,N_29053,N_29470);
nand UO_2149 (O_2149,N_29687,N_29403);
and UO_2150 (O_2150,N_28871,N_28809);
nor UO_2151 (O_2151,N_29401,N_28793);
or UO_2152 (O_2152,N_28649,N_28547);
or UO_2153 (O_2153,N_29492,N_29752);
or UO_2154 (O_2154,N_29587,N_28761);
nor UO_2155 (O_2155,N_29371,N_28840);
and UO_2156 (O_2156,N_28609,N_28585);
or UO_2157 (O_2157,N_29909,N_28501);
nor UO_2158 (O_2158,N_28810,N_28592);
and UO_2159 (O_2159,N_28932,N_29818);
xor UO_2160 (O_2160,N_29177,N_29788);
and UO_2161 (O_2161,N_28642,N_29348);
nand UO_2162 (O_2162,N_29373,N_29088);
and UO_2163 (O_2163,N_29924,N_29346);
and UO_2164 (O_2164,N_28768,N_29433);
nor UO_2165 (O_2165,N_28828,N_29578);
or UO_2166 (O_2166,N_28808,N_29825);
nor UO_2167 (O_2167,N_28810,N_28746);
xor UO_2168 (O_2168,N_29804,N_28983);
nand UO_2169 (O_2169,N_29781,N_28990);
and UO_2170 (O_2170,N_29541,N_29030);
nand UO_2171 (O_2171,N_29468,N_29825);
nand UO_2172 (O_2172,N_28882,N_29717);
or UO_2173 (O_2173,N_29871,N_28946);
xnor UO_2174 (O_2174,N_28711,N_29588);
and UO_2175 (O_2175,N_29972,N_28778);
nand UO_2176 (O_2176,N_29545,N_28964);
xor UO_2177 (O_2177,N_29970,N_29309);
xnor UO_2178 (O_2178,N_29389,N_29271);
xor UO_2179 (O_2179,N_29116,N_29327);
or UO_2180 (O_2180,N_28633,N_29529);
nand UO_2181 (O_2181,N_28510,N_29611);
or UO_2182 (O_2182,N_28975,N_29308);
or UO_2183 (O_2183,N_28967,N_29739);
and UO_2184 (O_2184,N_28799,N_28766);
or UO_2185 (O_2185,N_29307,N_28855);
or UO_2186 (O_2186,N_29709,N_29396);
and UO_2187 (O_2187,N_29916,N_29807);
nor UO_2188 (O_2188,N_29322,N_28553);
or UO_2189 (O_2189,N_28645,N_28547);
nor UO_2190 (O_2190,N_29778,N_29696);
nor UO_2191 (O_2191,N_29829,N_29853);
and UO_2192 (O_2192,N_28965,N_29392);
or UO_2193 (O_2193,N_29219,N_29732);
xor UO_2194 (O_2194,N_29928,N_29358);
or UO_2195 (O_2195,N_29729,N_29629);
xor UO_2196 (O_2196,N_29226,N_29820);
nand UO_2197 (O_2197,N_28786,N_29340);
and UO_2198 (O_2198,N_28761,N_29654);
nor UO_2199 (O_2199,N_29564,N_29877);
and UO_2200 (O_2200,N_29216,N_29632);
xnor UO_2201 (O_2201,N_28510,N_29727);
nand UO_2202 (O_2202,N_29297,N_28639);
or UO_2203 (O_2203,N_29818,N_29549);
nor UO_2204 (O_2204,N_29870,N_29886);
xor UO_2205 (O_2205,N_29196,N_29790);
nand UO_2206 (O_2206,N_29641,N_28743);
nand UO_2207 (O_2207,N_29445,N_29214);
or UO_2208 (O_2208,N_29197,N_29489);
or UO_2209 (O_2209,N_28637,N_29348);
and UO_2210 (O_2210,N_29650,N_29364);
and UO_2211 (O_2211,N_29177,N_28709);
xor UO_2212 (O_2212,N_28502,N_29423);
xor UO_2213 (O_2213,N_29520,N_29872);
nand UO_2214 (O_2214,N_29114,N_29710);
xnor UO_2215 (O_2215,N_29287,N_28903);
or UO_2216 (O_2216,N_29646,N_28840);
nor UO_2217 (O_2217,N_29795,N_28553);
nor UO_2218 (O_2218,N_29850,N_28990);
xnor UO_2219 (O_2219,N_29046,N_29045);
nor UO_2220 (O_2220,N_29789,N_29205);
or UO_2221 (O_2221,N_28675,N_29449);
and UO_2222 (O_2222,N_28886,N_28730);
and UO_2223 (O_2223,N_29197,N_28660);
or UO_2224 (O_2224,N_29030,N_29205);
nor UO_2225 (O_2225,N_29479,N_28771);
nand UO_2226 (O_2226,N_29976,N_29316);
or UO_2227 (O_2227,N_29241,N_29420);
xnor UO_2228 (O_2228,N_29744,N_29770);
or UO_2229 (O_2229,N_28938,N_29496);
and UO_2230 (O_2230,N_28944,N_28783);
nand UO_2231 (O_2231,N_29240,N_28769);
and UO_2232 (O_2232,N_28838,N_29642);
xor UO_2233 (O_2233,N_29338,N_28953);
and UO_2234 (O_2234,N_29404,N_28733);
nor UO_2235 (O_2235,N_29077,N_29744);
and UO_2236 (O_2236,N_29807,N_29326);
or UO_2237 (O_2237,N_29287,N_28531);
nand UO_2238 (O_2238,N_29419,N_29974);
or UO_2239 (O_2239,N_29744,N_29522);
xnor UO_2240 (O_2240,N_29249,N_29061);
or UO_2241 (O_2241,N_28948,N_29594);
nor UO_2242 (O_2242,N_28790,N_29819);
or UO_2243 (O_2243,N_29256,N_29390);
or UO_2244 (O_2244,N_28695,N_29091);
nor UO_2245 (O_2245,N_29843,N_28883);
nor UO_2246 (O_2246,N_29243,N_29138);
or UO_2247 (O_2247,N_29488,N_28980);
xnor UO_2248 (O_2248,N_29985,N_29099);
or UO_2249 (O_2249,N_29833,N_29952);
xor UO_2250 (O_2250,N_29761,N_29081);
nand UO_2251 (O_2251,N_28886,N_29285);
and UO_2252 (O_2252,N_29082,N_29718);
xnor UO_2253 (O_2253,N_29033,N_29425);
and UO_2254 (O_2254,N_29227,N_29916);
or UO_2255 (O_2255,N_29758,N_29403);
xnor UO_2256 (O_2256,N_28646,N_28919);
or UO_2257 (O_2257,N_28647,N_29427);
or UO_2258 (O_2258,N_29308,N_29447);
or UO_2259 (O_2259,N_29170,N_28862);
or UO_2260 (O_2260,N_29490,N_29168);
and UO_2261 (O_2261,N_29868,N_29482);
or UO_2262 (O_2262,N_29976,N_29633);
and UO_2263 (O_2263,N_28993,N_29315);
and UO_2264 (O_2264,N_29917,N_29338);
nand UO_2265 (O_2265,N_28763,N_29149);
and UO_2266 (O_2266,N_28703,N_29080);
nor UO_2267 (O_2267,N_29929,N_29136);
nand UO_2268 (O_2268,N_29213,N_29438);
or UO_2269 (O_2269,N_29481,N_29797);
and UO_2270 (O_2270,N_29575,N_28573);
and UO_2271 (O_2271,N_28699,N_29622);
nor UO_2272 (O_2272,N_29090,N_29835);
nor UO_2273 (O_2273,N_28673,N_29048);
nor UO_2274 (O_2274,N_28534,N_29482);
or UO_2275 (O_2275,N_29817,N_29781);
xnor UO_2276 (O_2276,N_28914,N_29480);
nor UO_2277 (O_2277,N_29529,N_28621);
nand UO_2278 (O_2278,N_28990,N_29211);
nor UO_2279 (O_2279,N_29914,N_29324);
nand UO_2280 (O_2280,N_28873,N_29933);
xnor UO_2281 (O_2281,N_29875,N_29347);
nor UO_2282 (O_2282,N_29908,N_29694);
nor UO_2283 (O_2283,N_29063,N_29792);
and UO_2284 (O_2284,N_28882,N_29414);
nand UO_2285 (O_2285,N_29418,N_28804);
and UO_2286 (O_2286,N_28915,N_28864);
or UO_2287 (O_2287,N_28625,N_29542);
nor UO_2288 (O_2288,N_29350,N_29813);
nor UO_2289 (O_2289,N_29605,N_29868);
and UO_2290 (O_2290,N_29502,N_29857);
or UO_2291 (O_2291,N_29559,N_29373);
nand UO_2292 (O_2292,N_29857,N_28571);
or UO_2293 (O_2293,N_29621,N_29799);
and UO_2294 (O_2294,N_29140,N_28971);
and UO_2295 (O_2295,N_29870,N_29124);
and UO_2296 (O_2296,N_29498,N_29084);
and UO_2297 (O_2297,N_29696,N_29333);
nor UO_2298 (O_2298,N_29763,N_28989);
and UO_2299 (O_2299,N_29252,N_28649);
xnor UO_2300 (O_2300,N_28861,N_28675);
or UO_2301 (O_2301,N_28810,N_28628);
xor UO_2302 (O_2302,N_29442,N_28637);
nor UO_2303 (O_2303,N_28682,N_29431);
xor UO_2304 (O_2304,N_28642,N_28863);
xnor UO_2305 (O_2305,N_29228,N_29413);
nand UO_2306 (O_2306,N_29878,N_29409);
nand UO_2307 (O_2307,N_29867,N_29167);
xor UO_2308 (O_2308,N_29717,N_28616);
nor UO_2309 (O_2309,N_29048,N_29880);
and UO_2310 (O_2310,N_29372,N_28885);
nor UO_2311 (O_2311,N_29637,N_28539);
and UO_2312 (O_2312,N_29856,N_29984);
nand UO_2313 (O_2313,N_29562,N_28841);
nor UO_2314 (O_2314,N_29837,N_28823);
nand UO_2315 (O_2315,N_29317,N_29453);
xor UO_2316 (O_2316,N_29396,N_28501);
or UO_2317 (O_2317,N_29770,N_28629);
nand UO_2318 (O_2318,N_28804,N_29947);
and UO_2319 (O_2319,N_29156,N_29737);
nand UO_2320 (O_2320,N_29166,N_29615);
nand UO_2321 (O_2321,N_29456,N_28850);
and UO_2322 (O_2322,N_29140,N_29636);
and UO_2323 (O_2323,N_29763,N_28906);
nand UO_2324 (O_2324,N_29866,N_28971);
nand UO_2325 (O_2325,N_29282,N_29656);
xnor UO_2326 (O_2326,N_29824,N_29692);
nor UO_2327 (O_2327,N_29491,N_29247);
nor UO_2328 (O_2328,N_29388,N_29921);
nor UO_2329 (O_2329,N_28666,N_29067);
nor UO_2330 (O_2330,N_29383,N_29391);
nor UO_2331 (O_2331,N_29280,N_28508);
and UO_2332 (O_2332,N_29649,N_29063);
or UO_2333 (O_2333,N_29663,N_28608);
nor UO_2334 (O_2334,N_29239,N_29726);
or UO_2335 (O_2335,N_28877,N_29364);
xor UO_2336 (O_2336,N_29243,N_28836);
or UO_2337 (O_2337,N_29890,N_29735);
nand UO_2338 (O_2338,N_29498,N_29610);
and UO_2339 (O_2339,N_29764,N_28979);
nand UO_2340 (O_2340,N_29789,N_29052);
nor UO_2341 (O_2341,N_28682,N_29323);
and UO_2342 (O_2342,N_29487,N_29155);
xnor UO_2343 (O_2343,N_29425,N_28781);
and UO_2344 (O_2344,N_29336,N_29691);
nor UO_2345 (O_2345,N_29942,N_29394);
and UO_2346 (O_2346,N_29831,N_29784);
and UO_2347 (O_2347,N_28525,N_29144);
and UO_2348 (O_2348,N_29747,N_28937);
xor UO_2349 (O_2349,N_28669,N_29004);
and UO_2350 (O_2350,N_29902,N_29546);
xnor UO_2351 (O_2351,N_29057,N_29192);
nand UO_2352 (O_2352,N_29872,N_29551);
nand UO_2353 (O_2353,N_29223,N_28519);
nor UO_2354 (O_2354,N_29886,N_29204);
nor UO_2355 (O_2355,N_29567,N_29044);
and UO_2356 (O_2356,N_28643,N_29590);
or UO_2357 (O_2357,N_28505,N_29293);
and UO_2358 (O_2358,N_29395,N_29768);
xnor UO_2359 (O_2359,N_29573,N_29968);
nand UO_2360 (O_2360,N_29445,N_28830);
nor UO_2361 (O_2361,N_29106,N_28746);
nand UO_2362 (O_2362,N_29282,N_28692);
nand UO_2363 (O_2363,N_28978,N_29194);
nand UO_2364 (O_2364,N_29705,N_29499);
nor UO_2365 (O_2365,N_28565,N_29698);
nor UO_2366 (O_2366,N_29117,N_28791);
or UO_2367 (O_2367,N_28623,N_29057);
or UO_2368 (O_2368,N_28913,N_28914);
xnor UO_2369 (O_2369,N_29041,N_28807);
xnor UO_2370 (O_2370,N_29843,N_29237);
and UO_2371 (O_2371,N_29037,N_29387);
nor UO_2372 (O_2372,N_29128,N_29589);
or UO_2373 (O_2373,N_28682,N_29293);
nand UO_2374 (O_2374,N_29497,N_29839);
nand UO_2375 (O_2375,N_28595,N_29994);
or UO_2376 (O_2376,N_29886,N_28797);
or UO_2377 (O_2377,N_29764,N_29124);
and UO_2378 (O_2378,N_29534,N_29140);
nand UO_2379 (O_2379,N_29954,N_28902);
and UO_2380 (O_2380,N_28927,N_29367);
or UO_2381 (O_2381,N_29693,N_29691);
nor UO_2382 (O_2382,N_29210,N_29970);
or UO_2383 (O_2383,N_29219,N_29719);
and UO_2384 (O_2384,N_28646,N_29521);
and UO_2385 (O_2385,N_29213,N_29902);
nand UO_2386 (O_2386,N_29574,N_29967);
nand UO_2387 (O_2387,N_29674,N_29228);
nand UO_2388 (O_2388,N_29209,N_29746);
nor UO_2389 (O_2389,N_28549,N_29780);
and UO_2390 (O_2390,N_29208,N_29045);
nor UO_2391 (O_2391,N_28886,N_29739);
or UO_2392 (O_2392,N_29322,N_28615);
nor UO_2393 (O_2393,N_29296,N_28926);
nor UO_2394 (O_2394,N_29345,N_28704);
nor UO_2395 (O_2395,N_29366,N_29176);
or UO_2396 (O_2396,N_29787,N_29542);
xor UO_2397 (O_2397,N_29654,N_28770);
nand UO_2398 (O_2398,N_28619,N_28668);
or UO_2399 (O_2399,N_29834,N_29929);
nor UO_2400 (O_2400,N_28821,N_29252);
xnor UO_2401 (O_2401,N_29578,N_29032);
xor UO_2402 (O_2402,N_29618,N_29870);
or UO_2403 (O_2403,N_29484,N_28839);
and UO_2404 (O_2404,N_29201,N_29268);
and UO_2405 (O_2405,N_29688,N_29980);
and UO_2406 (O_2406,N_29371,N_28959);
or UO_2407 (O_2407,N_29927,N_29824);
or UO_2408 (O_2408,N_29276,N_29497);
nor UO_2409 (O_2409,N_29349,N_28613);
and UO_2410 (O_2410,N_28667,N_29612);
xor UO_2411 (O_2411,N_29734,N_29899);
nand UO_2412 (O_2412,N_28917,N_28539);
xor UO_2413 (O_2413,N_28730,N_29674);
nand UO_2414 (O_2414,N_29759,N_29357);
xnor UO_2415 (O_2415,N_28763,N_29611);
or UO_2416 (O_2416,N_29167,N_29038);
xnor UO_2417 (O_2417,N_29296,N_28806);
xor UO_2418 (O_2418,N_29355,N_29596);
xor UO_2419 (O_2419,N_29442,N_29656);
xnor UO_2420 (O_2420,N_29389,N_28758);
nand UO_2421 (O_2421,N_28811,N_29659);
nand UO_2422 (O_2422,N_28960,N_29457);
and UO_2423 (O_2423,N_29275,N_29250);
nor UO_2424 (O_2424,N_29358,N_28646);
and UO_2425 (O_2425,N_29365,N_29621);
nor UO_2426 (O_2426,N_29273,N_28833);
xor UO_2427 (O_2427,N_29222,N_28613);
nand UO_2428 (O_2428,N_28580,N_29785);
or UO_2429 (O_2429,N_28535,N_28551);
or UO_2430 (O_2430,N_29720,N_29657);
xor UO_2431 (O_2431,N_28543,N_29246);
and UO_2432 (O_2432,N_29353,N_29475);
nor UO_2433 (O_2433,N_29267,N_29144);
nor UO_2434 (O_2434,N_28836,N_29190);
nand UO_2435 (O_2435,N_28560,N_28955);
and UO_2436 (O_2436,N_28838,N_29282);
nand UO_2437 (O_2437,N_28952,N_28807);
xor UO_2438 (O_2438,N_29255,N_29258);
or UO_2439 (O_2439,N_29665,N_28511);
nor UO_2440 (O_2440,N_29214,N_29612);
nand UO_2441 (O_2441,N_29944,N_29930);
nor UO_2442 (O_2442,N_28696,N_28775);
nor UO_2443 (O_2443,N_28614,N_29618);
and UO_2444 (O_2444,N_28947,N_29966);
and UO_2445 (O_2445,N_28970,N_29815);
or UO_2446 (O_2446,N_29246,N_29764);
nand UO_2447 (O_2447,N_29558,N_29457);
nor UO_2448 (O_2448,N_29648,N_28738);
xor UO_2449 (O_2449,N_29986,N_28904);
xor UO_2450 (O_2450,N_29294,N_28813);
or UO_2451 (O_2451,N_28817,N_29097);
nand UO_2452 (O_2452,N_29623,N_29616);
xnor UO_2453 (O_2453,N_29499,N_29748);
or UO_2454 (O_2454,N_29246,N_29358);
nor UO_2455 (O_2455,N_29596,N_28796);
and UO_2456 (O_2456,N_28696,N_29095);
nand UO_2457 (O_2457,N_29573,N_28735);
xor UO_2458 (O_2458,N_29974,N_28955);
and UO_2459 (O_2459,N_29907,N_28902);
nor UO_2460 (O_2460,N_28720,N_29450);
or UO_2461 (O_2461,N_29151,N_29147);
nand UO_2462 (O_2462,N_28647,N_28532);
nand UO_2463 (O_2463,N_29131,N_28944);
and UO_2464 (O_2464,N_29175,N_29271);
or UO_2465 (O_2465,N_28689,N_29186);
and UO_2466 (O_2466,N_29844,N_29332);
xor UO_2467 (O_2467,N_29332,N_29642);
nor UO_2468 (O_2468,N_29178,N_29388);
nor UO_2469 (O_2469,N_28767,N_28940);
nand UO_2470 (O_2470,N_29250,N_28521);
nor UO_2471 (O_2471,N_29001,N_29333);
xnor UO_2472 (O_2472,N_29881,N_29963);
nor UO_2473 (O_2473,N_28723,N_29386);
nand UO_2474 (O_2474,N_28949,N_28816);
nand UO_2475 (O_2475,N_29920,N_29157);
nand UO_2476 (O_2476,N_28954,N_29303);
nor UO_2477 (O_2477,N_29189,N_29555);
or UO_2478 (O_2478,N_28715,N_29216);
nor UO_2479 (O_2479,N_29496,N_29530);
and UO_2480 (O_2480,N_28528,N_28995);
nor UO_2481 (O_2481,N_28965,N_29987);
nand UO_2482 (O_2482,N_28829,N_28767);
or UO_2483 (O_2483,N_28955,N_29285);
xor UO_2484 (O_2484,N_28887,N_28587);
nor UO_2485 (O_2485,N_28615,N_29737);
xor UO_2486 (O_2486,N_29391,N_29647);
xor UO_2487 (O_2487,N_29947,N_29708);
xor UO_2488 (O_2488,N_28874,N_29943);
nor UO_2489 (O_2489,N_29885,N_29306);
nand UO_2490 (O_2490,N_28570,N_29577);
nor UO_2491 (O_2491,N_29733,N_29578);
and UO_2492 (O_2492,N_29120,N_29947);
and UO_2493 (O_2493,N_29221,N_28952);
nor UO_2494 (O_2494,N_29140,N_29715);
xor UO_2495 (O_2495,N_29659,N_28585);
nor UO_2496 (O_2496,N_28559,N_29055);
or UO_2497 (O_2497,N_29397,N_29402);
nor UO_2498 (O_2498,N_29574,N_29742);
xor UO_2499 (O_2499,N_28851,N_28514);
or UO_2500 (O_2500,N_28842,N_28537);
xor UO_2501 (O_2501,N_28729,N_28620);
or UO_2502 (O_2502,N_29868,N_28699);
and UO_2503 (O_2503,N_29837,N_29631);
and UO_2504 (O_2504,N_28825,N_29567);
or UO_2505 (O_2505,N_29265,N_29590);
and UO_2506 (O_2506,N_29017,N_29638);
and UO_2507 (O_2507,N_29786,N_28696);
nand UO_2508 (O_2508,N_28684,N_28908);
nand UO_2509 (O_2509,N_29713,N_29271);
and UO_2510 (O_2510,N_29682,N_28914);
nor UO_2511 (O_2511,N_29044,N_29232);
nand UO_2512 (O_2512,N_29215,N_29631);
nand UO_2513 (O_2513,N_29630,N_29536);
nor UO_2514 (O_2514,N_28942,N_29056);
nand UO_2515 (O_2515,N_29959,N_29462);
nor UO_2516 (O_2516,N_28951,N_29156);
or UO_2517 (O_2517,N_29278,N_29937);
xor UO_2518 (O_2518,N_28816,N_29474);
nand UO_2519 (O_2519,N_29705,N_28542);
or UO_2520 (O_2520,N_29075,N_29785);
nor UO_2521 (O_2521,N_28814,N_29429);
nand UO_2522 (O_2522,N_29060,N_29048);
or UO_2523 (O_2523,N_29874,N_29725);
nor UO_2524 (O_2524,N_29646,N_28856);
or UO_2525 (O_2525,N_29167,N_29236);
nor UO_2526 (O_2526,N_29908,N_28690);
xor UO_2527 (O_2527,N_28755,N_29642);
nor UO_2528 (O_2528,N_29927,N_28858);
nor UO_2529 (O_2529,N_28686,N_28957);
or UO_2530 (O_2530,N_29793,N_28834);
or UO_2531 (O_2531,N_29286,N_28594);
nor UO_2532 (O_2532,N_29238,N_29197);
and UO_2533 (O_2533,N_29881,N_29068);
and UO_2534 (O_2534,N_28760,N_29628);
and UO_2535 (O_2535,N_29502,N_29532);
or UO_2536 (O_2536,N_28898,N_28619);
and UO_2537 (O_2537,N_28557,N_29726);
or UO_2538 (O_2538,N_28673,N_28691);
and UO_2539 (O_2539,N_29793,N_29585);
xnor UO_2540 (O_2540,N_29525,N_28855);
nand UO_2541 (O_2541,N_28524,N_29100);
xnor UO_2542 (O_2542,N_28872,N_29666);
nand UO_2543 (O_2543,N_28678,N_29281);
or UO_2544 (O_2544,N_29233,N_29539);
nand UO_2545 (O_2545,N_29464,N_29043);
nand UO_2546 (O_2546,N_29180,N_28980);
nor UO_2547 (O_2547,N_29403,N_28888);
or UO_2548 (O_2548,N_29933,N_28978);
and UO_2549 (O_2549,N_29132,N_29712);
nor UO_2550 (O_2550,N_29218,N_29922);
or UO_2551 (O_2551,N_29841,N_28633);
xor UO_2552 (O_2552,N_28597,N_28791);
and UO_2553 (O_2553,N_29232,N_29594);
xnor UO_2554 (O_2554,N_28513,N_29536);
and UO_2555 (O_2555,N_29837,N_29093);
xnor UO_2556 (O_2556,N_29600,N_29617);
xnor UO_2557 (O_2557,N_29307,N_28614);
and UO_2558 (O_2558,N_28919,N_28707);
xnor UO_2559 (O_2559,N_29787,N_29299);
or UO_2560 (O_2560,N_28607,N_28771);
or UO_2561 (O_2561,N_28621,N_28650);
xnor UO_2562 (O_2562,N_29569,N_29369);
nand UO_2563 (O_2563,N_29361,N_28587);
xnor UO_2564 (O_2564,N_29992,N_29616);
and UO_2565 (O_2565,N_29830,N_29493);
and UO_2566 (O_2566,N_28677,N_29998);
xor UO_2567 (O_2567,N_29386,N_28988);
or UO_2568 (O_2568,N_29770,N_28653);
or UO_2569 (O_2569,N_29371,N_29551);
and UO_2570 (O_2570,N_29730,N_29695);
nor UO_2571 (O_2571,N_29695,N_29093);
nor UO_2572 (O_2572,N_29880,N_29248);
nor UO_2573 (O_2573,N_29663,N_29334);
and UO_2574 (O_2574,N_29087,N_29735);
nor UO_2575 (O_2575,N_29313,N_29703);
and UO_2576 (O_2576,N_29163,N_29904);
and UO_2577 (O_2577,N_29984,N_28979);
and UO_2578 (O_2578,N_28654,N_29171);
or UO_2579 (O_2579,N_28868,N_28717);
or UO_2580 (O_2580,N_28906,N_29066);
nor UO_2581 (O_2581,N_29286,N_28802);
nor UO_2582 (O_2582,N_28909,N_28519);
nor UO_2583 (O_2583,N_29517,N_29554);
nor UO_2584 (O_2584,N_29617,N_29411);
and UO_2585 (O_2585,N_29936,N_29733);
xor UO_2586 (O_2586,N_29009,N_29257);
nand UO_2587 (O_2587,N_28519,N_29512);
nand UO_2588 (O_2588,N_29010,N_28806);
and UO_2589 (O_2589,N_28933,N_28563);
nor UO_2590 (O_2590,N_29851,N_29668);
and UO_2591 (O_2591,N_29917,N_29419);
nor UO_2592 (O_2592,N_28859,N_29004);
nor UO_2593 (O_2593,N_29720,N_29894);
xnor UO_2594 (O_2594,N_29854,N_28731);
and UO_2595 (O_2595,N_28805,N_28642);
xor UO_2596 (O_2596,N_29303,N_29051);
nor UO_2597 (O_2597,N_28955,N_29009);
or UO_2598 (O_2598,N_28792,N_28751);
nand UO_2599 (O_2599,N_28851,N_29148);
or UO_2600 (O_2600,N_29762,N_29689);
nor UO_2601 (O_2601,N_29039,N_28873);
and UO_2602 (O_2602,N_29631,N_28618);
nor UO_2603 (O_2603,N_29454,N_28529);
or UO_2604 (O_2604,N_29129,N_29437);
nor UO_2605 (O_2605,N_28806,N_29343);
or UO_2606 (O_2606,N_28739,N_29210);
nor UO_2607 (O_2607,N_29287,N_28959);
and UO_2608 (O_2608,N_29872,N_28690);
or UO_2609 (O_2609,N_29413,N_29280);
xnor UO_2610 (O_2610,N_29979,N_28817);
nor UO_2611 (O_2611,N_28577,N_29285);
and UO_2612 (O_2612,N_28526,N_29599);
xnor UO_2613 (O_2613,N_29632,N_29645);
nor UO_2614 (O_2614,N_28856,N_29601);
xnor UO_2615 (O_2615,N_28662,N_28705);
xnor UO_2616 (O_2616,N_29089,N_28863);
and UO_2617 (O_2617,N_29898,N_29243);
nor UO_2618 (O_2618,N_29511,N_29887);
xor UO_2619 (O_2619,N_29211,N_28609);
or UO_2620 (O_2620,N_29920,N_28700);
xor UO_2621 (O_2621,N_29939,N_29327);
and UO_2622 (O_2622,N_29247,N_29686);
nand UO_2623 (O_2623,N_28687,N_29538);
nand UO_2624 (O_2624,N_29242,N_29277);
nand UO_2625 (O_2625,N_29364,N_29406);
xnor UO_2626 (O_2626,N_29863,N_29785);
nand UO_2627 (O_2627,N_29502,N_29287);
xor UO_2628 (O_2628,N_29815,N_28766);
nor UO_2629 (O_2629,N_29919,N_29022);
nor UO_2630 (O_2630,N_29741,N_28701);
nand UO_2631 (O_2631,N_29368,N_28935);
or UO_2632 (O_2632,N_29845,N_29905);
and UO_2633 (O_2633,N_29978,N_29501);
nor UO_2634 (O_2634,N_28748,N_29267);
nand UO_2635 (O_2635,N_29035,N_29996);
nor UO_2636 (O_2636,N_29279,N_29032);
nand UO_2637 (O_2637,N_29806,N_28720);
nand UO_2638 (O_2638,N_29187,N_29348);
xnor UO_2639 (O_2639,N_29952,N_29808);
nor UO_2640 (O_2640,N_28930,N_29355);
xor UO_2641 (O_2641,N_29011,N_29016);
or UO_2642 (O_2642,N_29900,N_29365);
and UO_2643 (O_2643,N_28712,N_29911);
or UO_2644 (O_2644,N_29070,N_28898);
xnor UO_2645 (O_2645,N_29507,N_29411);
and UO_2646 (O_2646,N_29741,N_28592);
and UO_2647 (O_2647,N_29409,N_29835);
and UO_2648 (O_2648,N_29109,N_29121);
or UO_2649 (O_2649,N_28966,N_29796);
nand UO_2650 (O_2650,N_29715,N_29654);
or UO_2651 (O_2651,N_28593,N_28903);
xnor UO_2652 (O_2652,N_28555,N_28777);
xor UO_2653 (O_2653,N_29531,N_29293);
nor UO_2654 (O_2654,N_29651,N_29907);
or UO_2655 (O_2655,N_29381,N_29901);
and UO_2656 (O_2656,N_29646,N_28952);
nand UO_2657 (O_2657,N_28883,N_29481);
xor UO_2658 (O_2658,N_29909,N_28869);
nand UO_2659 (O_2659,N_28713,N_29705);
nand UO_2660 (O_2660,N_28700,N_28722);
or UO_2661 (O_2661,N_29603,N_29347);
nor UO_2662 (O_2662,N_28746,N_29155);
nor UO_2663 (O_2663,N_29261,N_29037);
xnor UO_2664 (O_2664,N_29541,N_29753);
or UO_2665 (O_2665,N_29133,N_29414);
nand UO_2666 (O_2666,N_28866,N_29526);
nor UO_2667 (O_2667,N_29072,N_29387);
nand UO_2668 (O_2668,N_29551,N_28746);
and UO_2669 (O_2669,N_28624,N_29061);
nor UO_2670 (O_2670,N_28936,N_29599);
or UO_2671 (O_2671,N_29323,N_29413);
xor UO_2672 (O_2672,N_28662,N_28688);
xnor UO_2673 (O_2673,N_29785,N_28940);
nand UO_2674 (O_2674,N_29805,N_29509);
nand UO_2675 (O_2675,N_29108,N_28642);
nand UO_2676 (O_2676,N_28936,N_29465);
and UO_2677 (O_2677,N_28580,N_29589);
or UO_2678 (O_2678,N_28893,N_29207);
nand UO_2679 (O_2679,N_28551,N_28622);
xnor UO_2680 (O_2680,N_29916,N_28986);
xor UO_2681 (O_2681,N_29204,N_28631);
xor UO_2682 (O_2682,N_29280,N_28639);
nand UO_2683 (O_2683,N_29720,N_29084);
nand UO_2684 (O_2684,N_28821,N_29466);
nand UO_2685 (O_2685,N_28747,N_28760);
nor UO_2686 (O_2686,N_29107,N_29242);
nand UO_2687 (O_2687,N_28941,N_29438);
xnor UO_2688 (O_2688,N_28552,N_29970);
nand UO_2689 (O_2689,N_28774,N_29413);
or UO_2690 (O_2690,N_28552,N_29582);
nand UO_2691 (O_2691,N_29565,N_29692);
nor UO_2692 (O_2692,N_29890,N_28965);
or UO_2693 (O_2693,N_28770,N_29031);
nor UO_2694 (O_2694,N_28631,N_29975);
xnor UO_2695 (O_2695,N_28709,N_28780);
and UO_2696 (O_2696,N_29943,N_28726);
nand UO_2697 (O_2697,N_28819,N_28531);
or UO_2698 (O_2698,N_28644,N_29840);
nor UO_2699 (O_2699,N_29883,N_29006);
nand UO_2700 (O_2700,N_29424,N_29551);
and UO_2701 (O_2701,N_29974,N_29194);
nand UO_2702 (O_2702,N_29598,N_28654);
nand UO_2703 (O_2703,N_29602,N_28569);
xor UO_2704 (O_2704,N_29334,N_29723);
nor UO_2705 (O_2705,N_28744,N_29454);
nand UO_2706 (O_2706,N_28992,N_28735);
or UO_2707 (O_2707,N_28786,N_28640);
nand UO_2708 (O_2708,N_28909,N_28736);
and UO_2709 (O_2709,N_29929,N_28622);
nor UO_2710 (O_2710,N_28564,N_29228);
and UO_2711 (O_2711,N_28771,N_29036);
xnor UO_2712 (O_2712,N_29525,N_28658);
nor UO_2713 (O_2713,N_29017,N_29371);
nand UO_2714 (O_2714,N_28585,N_29243);
or UO_2715 (O_2715,N_29999,N_29816);
and UO_2716 (O_2716,N_28743,N_29895);
and UO_2717 (O_2717,N_29744,N_29620);
xnor UO_2718 (O_2718,N_28858,N_29334);
and UO_2719 (O_2719,N_29073,N_29889);
and UO_2720 (O_2720,N_29562,N_28889);
nand UO_2721 (O_2721,N_28789,N_28761);
or UO_2722 (O_2722,N_29097,N_29453);
and UO_2723 (O_2723,N_29238,N_28638);
xnor UO_2724 (O_2724,N_29563,N_28515);
or UO_2725 (O_2725,N_28954,N_28608);
nor UO_2726 (O_2726,N_29341,N_28947);
xor UO_2727 (O_2727,N_29916,N_29504);
and UO_2728 (O_2728,N_28712,N_29708);
nand UO_2729 (O_2729,N_29114,N_28507);
xor UO_2730 (O_2730,N_29629,N_28518);
and UO_2731 (O_2731,N_28929,N_28503);
nand UO_2732 (O_2732,N_28800,N_28826);
xor UO_2733 (O_2733,N_29417,N_29054);
xor UO_2734 (O_2734,N_29940,N_29570);
xnor UO_2735 (O_2735,N_28558,N_29348);
and UO_2736 (O_2736,N_28695,N_28893);
and UO_2737 (O_2737,N_28846,N_29361);
nand UO_2738 (O_2738,N_29659,N_28680);
nand UO_2739 (O_2739,N_28545,N_29371);
xnor UO_2740 (O_2740,N_29332,N_29831);
and UO_2741 (O_2741,N_29799,N_28770);
nor UO_2742 (O_2742,N_29427,N_28760);
nand UO_2743 (O_2743,N_28622,N_29987);
and UO_2744 (O_2744,N_29248,N_29160);
xnor UO_2745 (O_2745,N_28767,N_29808);
or UO_2746 (O_2746,N_29292,N_28825);
nor UO_2747 (O_2747,N_29737,N_28600);
and UO_2748 (O_2748,N_29039,N_29582);
xor UO_2749 (O_2749,N_28528,N_29597);
and UO_2750 (O_2750,N_29761,N_29985);
nor UO_2751 (O_2751,N_29115,N_29229);
nor UO_2752 (O_2752,N_29168,N_29605);
and UO_2753 (O_2753,N_28545,N_28526);
nand UO_2754 (O_2754,N_28671,N_29544);
or UO_2755 (O_2755,N_29966,N_29930);
or UO_2756 (O_2756,N_28905,N_29056);
nand UO_2757 (O_2757,N_28758,N_29494);
or UO_2758 (O_2758,N_29617,N_29695);
nor UO_2759 (O_2759,N_28900,N_28636);
nor UO_2760 (O_2760,N_29600,N_29587);
nor UO_2761 (O_2761,N_28600,N_28640);
or UO_2762 (O_2762,N_28611,N_28895);
or UO_2763 (O_2763,N_29373,N_28717);
or UO_2764 (O_2764,N_29121,N_28972);
and UO_2765 (O_2765,N_29084,N_29257);
and UO_2766 (O_2766,N_28872,N_29762);
nor UO_2767 (O_2767,N_29139,N_29199);
and UO_2768 (O_2768,N_28821,N_29392);
nand UO_2769 (O_2769,N_29283,N_29918);
or UO_2770 (O_2770,N_29912,N_29532);
and UO_2771 (O_2771,N_28907,N_28832);
or UO_2772 (O_2772,N_29097,N_28543);
or UO_2773 (O_2773,N_29000,N_29219);
and UO_2774 (O_2774,N_28558,N_29324);
nor UO_2775 (O_2775,N_29449,N_28615);
nand UO_2776 (O_2776,N_29984,N_29654);
or UO_2777 (O_2777,N_29245,N_29628);
and UO_2778 (O_2778,N_29202,N_29000);
or UO_2779 (O_2779,N_29622,N_28978);
xnor UO_2780 (O_2780,N_29428,N_28989);
or UO_2781 (O_2781,N_29929,N_29982);
xor UO_2782 (O_2782,N_29158,N_29519);
nor UO_2783 (O_2783,N_28952,N_29117);
nand UO_2784 (O_2784,N_29765,N_29401);
xnor UO_2785 (O_2785,N_29884,N_28558);
nand UO_2786 (O_2786,N_29392,N_28557);
and UO_2787 (O_2787,N_29931,N_29426);
or UO_2788 (O_2788,N_29921,N_29583);
nand UO_2789 (O_2789,N_29310,N_29863);
nor UO_2790 (O_2790,N_29736,N_28544);
and UO_2791 (O_2791,N_29778,N_28775);
and UO_2792 (O_2792,N_29670,N_29811);
xnor UO_2793 (O_2793,N_29060,N_29783);
and UO_2794 (O_2794,N_28634,N_28777);
or UO_2795 (O_2795,N_29656,N_29176);
xor UO_2796 (O_2796,N_28850,N_28825);
nand UO_2797 (O_2797,N_29443,N_29760);
xnor UO_2798 (O_2798,N_28702,N_29934);
or UO_2799 (O_2799,N_29949,N_28836);
nand UO_2800 (O_2800,N_28746,N_29302);
nor UO_2801 (O_2801,N_29201,N_29563);
xor UO_2802 (O_2802,N_29676,N_28646);
nand UO_2803 (O_2803,N_29370,N_29760);
or UO_2804 (O_2804,N_28543,N_28977);
nand UO_2805 (O_2805,N_28940,N_28507);
nor UO_2806 (O_2806,N_29927,N_28690);
nor UO_2807 (O_2807,N_28980,N_29701);
nand UO_2808 (O_2808,N_28935,N_29092);
nand UO_2809 (O_2809,N_29388,N_29072);
nor UO_2810 (O_2810,N_29643,N_29599);
xnor UO_2811 (O_2811,N_28927,N_29630);
or UO_2812 (O_2812,N_29563,N_29124);
and UO_2813 (O_2813,N_29283,N_29666);
or UO_2814 (O_2814,N_29880,N_28613);
and UO_2815 (O_2815,N_28834,N_28867);
nor UO_2816 (O_2816,N_29495,N_29255);
nand UO_2817 (O_2817,N_29982,N_28738);
nand UO_2818 (O_2818,N_28875,N_28545);
and UO_2819 (O_2819,N_29272,N_29837);
and UO_2820 (O_2820,N_29651,N_28948);
nor UO_2821 (O_2821,N_29608,N_28614);
and UO_2822 (O_2822,N_28941,N_29802);
or UO_2823 (O_2823,N_29665,N_28553);
xnor UO_2824 (O_2824,N_28791,N_29528);
or UO_2825 (O_2825,N_28834,N_29473);
or UO_2826 (O_2826,N_29637,N_29011);
nand UO_2827 (O_2827,N_28733,N_29680);
nor UO_2828 (O_2828,N_29883,N_28948);
nor UO_2829 (O_2829,N_29037,N_29382);
xnor UO_2830 (O_2830,N_29103,N_28585);
xnor UO_2831 (O_2831,N_29883,N_29637);
or UO_2832 (O_2832,N_29639,N_28779);
nor UO_2833 (O_2833,N_29819,N_28540);
or UO_2834 (O_2834,N_28635,N_29620);
nor UO_2835 (O_2835,N_29980,N_28979);
xnor UO_2836 (O_2836,N_29140,N_29956);
and UO_2837 (O_2837,N_28577,N_29843);
nand UO_2838 (O_2838,N_29979,N_28840);
nor UO_2839 (O_2839,N_28607,N_28924);
xnor UO_2840 (O_2840,N_28846,N_28502);
or UO_2841 (O_2841,N_28668,N_29699);
or UO_2842 (O_2842,N_29729,N_28999);
xnor UO_2843 (O_2843,N_29788,N_29792);
or UO_2844 (O_2844,N_28691,N_29018);
or UO_2845 (O_2845,N_28971,N_28515);
xor UO_2846 (O_2846,N_28623,N_29777);
nor UO_2847 (O_2847,N_29425,N_29967);
nand UO_2848 (O_2848,N_29018,N_29971);
and UO_2849 (O_2849,N_28706,N_28613);
xnor UO_2850 (O_2850,N_29700,N_28552);
or UO_2851 (O_2851,N_29802,N_29504);
nand UO_2852 (O_2852,N_29261,N_29460);
nand UO_2853 (O_2853,N_29188,N_29651);
and UO_2854 (O_2854,N_29965,N_29808);
nand UO_2855 (O_2855,N_28761,N_29355);
nor UO_2856 (O_2856,N_29788,N_29290);
and UO_2857 (O_2857,N_29072,N_29094);
and UO_2858 (O_2858,N_29525,N_28672);
nor UO_2859 (O_2859,N_29104,N_28982);
and UO_2860 (O_2860,N_29018,N_29448);
xnor UO_2861 (O_2861,N_29658,N_29493);
or UO_2862 (O_2862,N_29616,N_28961);
and UO_2863 (O_2863,N_29525,N_29824);
nor UO_2864 (O_2864,N_28555,N_29008);
nand UO_2865 (O_2865,N_28997,N_28673);
or UO_2866 (O_2866,N_29129,N_28892);
xnor UO_2867 (O_2867,N_28611,N_29445);
nor UO_2868 (O_2868,N_29053,N_29832);
or UO_2869 (O_2869,N_29646,N_28850);
nand UO_2870 (O_2870,N_29546,N_29514);
and UO_2871 (O_2871,N_29637,N_29227);
nor UO_2872 (O_2872,N_29996,N_29167);
xor UO_2873 (O_2873,N_29883,N_29636);
or UO_2874 (O_2874,N_28669,N_29526);
and UO_2875 (O_2875,N_29379,N_29273);
nand UO_2876 (O_2876,N_28807,N_29261);
nand UO_2877 (O_2877,N_29200,N_28948);
nor UO_2878 (O_2878,N_28997,N_29390);
and UO_2879 (O_2879,N_29914,N_28634);
and UO_2880 (O_2880,N_29911,N_29716);
or UO_2881 (O_2881,N_29673,N_28662);
nand UO_2882 (O_2882,N_29703,N_29592);
nand UO_2883 (O_2883,N_29073,N_29459);
and UO_2884 (O_2884,N_29482,N_29605);
xnor UO_2885 (O_2885,N_29486,N_29799);
xnor UO_2886 (O_2886,N_28982,N_29941);
and UO_2887 (O_2887,N_29254,N_29480);
nand UO_2888 (O_2888,N_29195,N_29454);
and UO_2889 (O_2889,N_28905,N_29021);
nor UO_2890 (O_2890,N_29183,N_29946);
nand UO_2891 (O_2891,N_28735,N_29822);
nor UO_2892 (O_2892,N_29922,N_29524);
or UO_2893 (O_2893,N_29350,N_29401);
nor UO_2894 (O_2894,N_29177,N_29942);
and UO_2895 (O_2895,N_29057,N_29120);
or UO_2896 (O_2896,N_29987,N_28589);
and UO_2897 (O_2897,N_29808,N_29555);
or UO_2898 (O_2898,N_29737,N_28958);
xor UO_2899 (O_2899,N_29740,N_29516);
nor UO_2900 (O_2900,N_29542,N_29867);
and UO_2901 (O_2901,N_29136,N_29612);
xnor UO_2902 (O_2902,N_29987,N_29582);
nand UO_2903 (O_2903,N_28773,N_28513);
or UO_2904 (O_2904,N_28982,N_29289);
and UO_2905 (O_2905,N_28626,N_29706);
or UO_2906 (O_2906,N_28577,N_28680);
or UO_2907 (O_2907,N_29986,N_29612);
and UO_2908 (O_2908,N_28527,N_29442);
nor UO_2909 (O_2909,N_29815,N_29411);
or UO_2910 (O_2910,N_28839,N_29392);
or UO_2911 (O_2911,N_29400,N_28755);
nor UO_2912 (O_2912,N_28824,N_28733);
xor UO_2913 (O_2913,N_29867,N_29702);
and UO_2914 (O_2914,N_28594,N_29024);
xnor UO_2915 (O_2915,N_29583,N_28739);
nand UO_2916 (O_2916,N_29530,N_28942);
nor UO_2917 (O_2917,N_29579,N_29422);
nor UO_2918 (O_2918,N_29391,N_28571);
and UO_2919 (O_2919,N_29730,N_29950);
nor UO_2920 (O_2920,N_28729,N_28759);
or UO_2921 (O_2921,N_29717,N_28636);
or UO_2922 (O_2922,N_29354,N_29941);
or UO_2923 (O_2923,N_29396,N_29365);
and UO_2924 (O_2924,N_28577,N_29090);
or UO_2925 (O_2925,N_29595,N_29477);
xor UO_2926 (O_2926,N_28762,N_28796);
nand UO_2927 (O_2927,N_28540,N_28594);
nor UO_2928 (O_2928,N_28871,N_29807);
xnor UO_2929 (O_2929,N_28759,N_29975);
and UO_2930 (O_2930,N_29993,N_29186);
xor UO_2931 (O_2931,N_28659,N_28985);
nand UO_2932 (O_2932,N_29603,N_29693);
and UO_2933 (O_2933,N_29956,N_29610);
nand UO_2934 (O_2934,N_28572,N_29202);
nand UO_2935 (O_2935,N_28602,N_29072);
or UO_2936 (O_2936,N_29744,N_29419);
or UO_2937 (O_2937,N_29094,N_29646);
nand UO_2938 (O_2938,N_29519,N_29662);
or UO_2939 (O_2939,N_28944,N_29184);
or UO_2940 (O_2940,N_28707,N_29383);
nor UO_2941 (O_2941,N_29893,N_29837);
nand UO_2942 (O_2942,N_29265,N_29327);
and UO_2943 (O_2943,N_29541,N_29135);
and UO_2944 (O_2944,N_29771,N_28811);
nand UO_2945 (O_2945,N_28810,N_29589);
nand UO_2946 (O_2946,N_28728,N_28735);
or UO_2947 (O_2947,N_29117,N_29123);
or UO_2948 (O_2948,N_28685,N_29056);
nand UO_2949 (O_2949,N_28672,N_28849);
nand UO_2950 (O_2950,N_29732,N_29622);
xnor UO_2951 (O_2951,N_29481,N_28964);
and UO_2952 (O_2952,N_28974,N_29496);
or UO_2953 (O_2953,N_29232,N_28765);
and UO_2954 (O_2954,N_29894,N_28894);
or UO_2955 (O_2955,N_28804,N_29309);
and UO_2956 (O_2956,N_29406,N_29699);
nor UO_2957 (O_2957,N_29946,N_29780);
nor UO_2958 (O_2958,N_29757,N_29579);
and UO_2959 (O_2959,N_29654,N_29193);
nand UO_2960 (O_2960,N_28937,N_29083);
and UO_2961 (O_2961,N_29174,N_29496);
xor UO_2962 (O_2962,N_29431,N_28901);
or UO_2963 (O_2963,N_29962,N_28896);
nand UO_2964 (O_2964,N_29608,N_29980);
xnor UO_2965 (O_2965,N_29572,N_29964);
nand UO_2966 (O_2966,N_29361,N_29383);
and UO_2967 (O_2967,N_28522,N_28721);
xnor UO_2968 (O_2968,N_29672,N_29294);
and UO_2969 (O_2969,N_28799,N_29805);
and UO_2970 (O_2970,N_29479,N_29846);
and UO_2971 (O_2971,N_29260,N_29079);
xnor UO_2972 (O_2972,N_28818,N_28867);
or UO_2973 (O_2973,N_28822,N_29571);
or UO_2974 (O_2974,N_29582,N_29119);
or UO_2975 (O_2975,N_29961,N_29695);
nand UO_2976 (O_2976,N_29255,N_29605);
and UO_2977 (O_2977,N_29742,N_29923);
nor UO_2978 (O_2978,N_29832,N_28734);
or UO_2979 (O_2979,N_28933,N_29065);
nor UO_2980 (O_2980,N_28825,N_29431);
or UO_2981 (O_2981,N_29775,N_28789);
nand UO_2982 (O_2982,N_28971,N_28565);
nor UO_2983 (O_2983,N_29890,N_29764);
or UO_2984 (O_2984,N_29206,N_29826);
or UO_2985 (O_2985,N_28934,N_29754);
and UO_2986 (O_2986,N_29412,N_29071);
or UO_2987 (O_2987,N_29573,N_29651);
and UO_2988 (O_2988,N_29264,N_29759);
xor UO_2989 (O_2989,N_28838,N_28507);
nand UO_2990 (O_2990,N_29830,N_29174);
nor UO_2991 (O_2991,N_29072,N_29589);
nor UO_2992 (O_2992,N_28678,N_29953);
nand UO_2993 (O_2993,N_29526,N_29089);
and UO_2994 (O_2994,N_29938,N_28675);
and UO_2995 (O_2995,N_28721,N_29154);
or UO_2996 (O_2996,N_29424,N_29654);
xor UO_2997 (O_2997,N_28732,N_29093);
nor UO_2998 (O_2998,N_29045,N_29705);
nor UO_2999 (O_2999,N_28787,N_29246);
and UO_3000 (O_3000,N_29879,N_28869);
xor UO_3001 (O_3001,N_29609,N_28722);
nor UO_3002 (O_3002,N_29755,N_28571);
nand UO_3003 (O_3003,N_29775,N_28576);
xnor UO_3004 (O_3004,N_28618,N_29727);
nor UO_3005 (O_3005,N_28694,N_28601);
nand UO_3006 (O_3006,N_29742,N_28535);
xnor UO_3007 (O_3007,N_28995,N_29263);
or UO_3008 (O_3008,N_29484,N_28583);
and UO_3009 (O_3009,N_29587,N_29233);
nand UO_3010 (O_3010,N_28716,N_29226);
and UO_3011 (O_3011,N_28670,N_29848);
xnor UO_3012 (O_3012,N_28930,N_29819);
and UO_3013 (O_3013,N_28907,N_28915);
xnor UO_3014 (O_3014,N_28866,N_28695);
xor UO_3015 (O_3015,N_28862,N_29299);
xor UO_3016 (O_3016,N_29893,N_29639);
xnor UO_3017 (O_3017,N_28694,N_29502);
nand UO_3018 (O_3018,N_29989,N_29366);
nand UO_3019 (O_3019,N_28870,N_29714);
nand UO_3020 (O_3020,N_29821,N_29484);
nor UO_3021 (O_3021,N_28622,N_29421);
nor UO_3022 (O_3022,N_28591,N_29977);
and UO_3023 (O_3023,N_29275,N_29042);
or UO_3024 (O_3024,N_28691,N_29805);
nor UO_3025 (O_3025,N_29985,N_29253);
and UO_3026 (O_3026,N_29733,N_29189);
nand UO_3027 (O_3027,N_29001,N_29922);
nor UO_3028 (O_3028,N_28934,N_28903);
xnor UO_3029 (O_3029,N_29277,N_29979);
or UO_3030 (O_3030,N_29391,N_28634);
or UO_3031 (O_3031,N_29885,N_29541);
and UO_3032 (O_3032,N_28613,N_28936);
xor UO_3033 (O_3033,N_29149,N_28533);
nor UO_3034 (O_3034,N_29743,N_29431);
xnor UO_3035 (O_3035,N_29771,N_29287);
and UO_3036 (O_3036,N_29047,N_28786);
nor UO_3037 (O_3037,N_29625,N_28872);
nand UO_3038 (O_3038,N_29662,N_29771);
nor UO_3039 (O_3039,N_29731,N_28517);
or UO_3040 (O_3040,N_29207,N_29496);
and UO_3041 (O_3041,N_28877,N_28783);
or UO_3042 (O_3042,N_29810,N_29258);
xnor UO_3043 (O_3043,N_28846,N_28797);
or UO_3044 (O_3044,N_28666,N_29795);
xor UO_3045 (O_3045,N_29774,N_29505);
or UO_3046 (O_3046,N_28968,N_29557);
or UO_3047 (O_3047,N_28553,N_29195);
or UO_3048 (O_3048,N_29467,N_29742);
or UO_3049 (O_3049,N_29609,N_28988);
xor UO_3050 (O_3050,N_28933,N_28887);
nand UO_3051 (O_3051,N_29622,N_29750);
nand UO_3052 (O_3052,N_29495,N_29593);
nor UO_3053 (O_3053,N_29022,N_28647);
nand UO_3054 (O_3054,N_28788,N_28735);
xnor UO_3055 (O_3055,N_29344,N_29872);
xnor UO_3056 (O_3056,N_29737,N_29982);
and UO_3057 (O_3057,N_29459,N_29256);
nor UO_3058 (O_3058,N_29432,N_29570);
xnor UO_3059 (O_3059,N_29089,N_28916);
and UO_3060 (O_3060,N_29632,N_29500);
nor UO_3061 (O_3061,N_29939,N_28802);
or UO_3062 (O_3062,N_29049,N_28611);
and UO_3063 (O_3063,N_29555,N_29683);
or UO_3064 (O_3064,N_29390,N_29800);
or UO_3065 (O_3065,N_29666,N_28642);
xor UO_3066 (O_3066,N_29017,N_29949);
nor UO_3067 (O_3067,N_29602,N_28932);
nand UO_3068 (O_3068,N_29318,N_28858);
and UO_3069 (O_3069,N_29412,N_29030);
xor UO_3070 (O_3070,N_29802,N_29649);
nor UO_3071 (O_3071,N_29730,N_28883);
xnor UO_3072 (O_3072,N_29140,N_29642);
nor UO_3073 (O_3073,N_28503,N_29243);
and UO_3074 (O_3074,N_28838,N_29849);
or UO_3075 (O_3075,N_29302,N_28562);
xnor UO_3076 (O_3076,N_29793,N_29730);
or UO_3077 (O_3077,N_29357,N_29054);
nand UO_3078 (O_3078,N_28977,N_29060);
or UO_3079 (O_3079,N_29394,N_29478);
nor UO_3080 (O_3080,N_29834,N_29616);
or UO_3081 (O_3081,N_29929,N_29022);
or UO_3082 (O_3082,N_29896,N_29461);
and UO_3083 (O_3083,N_29412,N_28697);
xor UO_3084 (O_3084,N_29704,N_29018);
xor UO_3085 (O_3085,N_28844,N_29059);
and UO_3086 (O_3086,N_29847,N_28699);
nor UO_3087 (O_3087,N_29061,N_29465);
xor UO_3088 (O_3088,N_29511,N_29085);
nor UO_3089 (O_3089,N_29395,N_29110);
and UO_3090 (O_3090,N_29445,N_28505);
xor UO_3091 (O_3091,N_29032,N_29689);
xnor UO_3092 (O_3092,N_28507,N_28670);
and UO_3093 (O_3093,N_28631,N_29862);
xnor UO_3094 (O_3094,N_29439,N_29374);
and UO_3095 (O_3095,N_28862,N_29946);
and UO_3096 (O_3096,N_28758,N_28669);
nor UO_3097 (O_3097,N_29698,N_28715);
nor UO_3098 (O_3098,N_28882,N_29608);
and UO_3099 (O_3099,N_29741,N_28839);
xnor UO_3100 (O_3100,N_28859,N_29191);
and UO_3101 (O_3101,N_29119,N_29010);
xnor UO_3102 (O_3102,N_29143,N_29402);
nand UO_3103 (O_3103,N_28751,N_28900);
nand UO_3104 (O_3104,N_29317,N_28911);
or UO_3105 (O_3105,N_29067,N_29665);
nor UO_3106 (O_3106,N_29070,N_29963);
or UO_3107 (O_3107,N_28946,N_29583);
or UO_3108 (O_3108,N_29574,N_29404);
nor UO_3109 (O_3109,N_29236,N_29072);
or UO_3110 (O_3110,N_28556,N_28891);
xnor UO_3111 (O_3111,N_29831,N_29099);
xor UO_3112 (O_3112,N_29219,N_28500);
or UO_3113 (O_3113,N_29307,N_29270);
xnor UO_3114 (O_3114,N_29617,N_29276);
nand UO_3115 (O_3115,N_29097,N_28519);
or UO_3116 (O_3116,N_29526,N_29180);
and UO_3117 (O_3117,N_28638,N_29885);
and UO_3118 (O_3118,N_29394,N_29549);
and UO_3119 (O_3119,N_28521,N_29494);
xor UO_3120 (O_3120,N_29931,N_29448);
xor UO_3121 (O_3121,N_29751,N_28739);
or UO_3122 (O_3122,N_29865,N_28842);
nand UO_3123 (O_3123,N_29694,N_28853);
or UO_3124 (O_3124,N_29788,N_29578);
nand UO_3125 (O_3125,N_29723,N_29491);
or UO_3126 (O_3126,N_28873,N_29580);
or UO_3127 (O_3127,N_29754,N_28993);
or UO_3128 (O_3128,N_29093,N_29993);
and UO_3129 (O_3129,N_29165,N_29235);
and UO_3130 (O_3130,N_29752,N_28575);
nor UO_3131 (O_3131,N_28552,N_29899);
and UO_3132 (O_3132,N_29221,N_28685);
nand UO_3133 (O_3133,N_29165,N_29162);
or UO_3134 (O_3134,N_29091,N_29788);
xor UO_3135 (O_3135,N_28964,N_29870);
and UO_3136 (O_3136,N_29501,N_28677);
and UO_3137 (O_3137,N_29044,N_29277);
nor UO_3138 (O_3138,N_28791,N_29088);
or UO_3139 (O_3139,N_28887,N_29270);
nor UO_3140 (O_3140,N_29254,N_29924);
nor UO_3141 (O_3141,N_29438,N_28585);
and UO_3142 (O_3142,N_29650,N_29551);
nand UO_3143 (O_3143,N_29581,N_29350);
nand UO_3144 (O_3144,N_29779,N_29625);
xor UO_3145 (O_3145,N_29217,N_29091);
nor UO_3146 (O_3146,N_29824,N_29158);
and UO_3147 (O_3147,N_28974,N_29582);
and UO_3148 (O_3148,N_29914,N_29991);
and UO_3149 (O_3149,N_29351,N_28625);
nor UO_3150 (O_3150,N_29725,N_28545);
or UO_3151 (O_3151,N_29460,N_28663);
nor UO_3152 (O_3152,N_29773,N_29835);
xnor UO_3153 (O_3153,N_28585,N_28871);
or UO_3154 (O_3154,N_29401,N_29599);
and UO_3155 (O_3155,N_28834,N_29726);
nand UO_3156 (O_3156,N_29798,N_29413);
or UO_3157 (O_3157,N_29453,N_29157);
nor UO_3158 (O_3158,N_29117,N_29829);
or UO_3159 (O_3159,N_28530,N_29617);
or UO_3160 (O_3160,N_29720,N_29881);
or UO_3161 (O_3161,N_28571,N_29599);
or UO_3162 (O_3162,N_29429,N_29187);
and UO_3163 (O_3163,N_29298,N_29598);
xor UO_3164 (O_3164,N_28782,N_29660);
and UO_3165 (O_3165,N_28697,N_29963);
and UO_3166 (O_3166,N_29626,N_29774);
nor UO_3167 (O_3167,N_29885,N_29660);
nor UO_3168 (O_3168,N_29995,N_29604);
nor UO_3169 (O_3169,N_29588,N_29737);
or UO_3170 (O_3170,N_29749,N_29930);
nand UO_3171 (O_3171,N_29569,N_29994);
nand UO_3172 (O_3172,N_29391,N_29975);
and UO_3173 (O_3173,N_28972,N_28739);
or UO_3174 (O_3174,N_29239,N_28847);
and UO_3175 (O_3175,N_28965,N_29414);
nand UO_3176 (O_3176,N_28572,N_29813);
xor UO_3177 (O_3177,N_29447,N_28589);
nor UO_3178 (O_3178,N_29903,N_29828);
xor UO_3179 (O_3179,N_28806,N_28881);
xnor UO_3180 (O_3180,N_28668,N_29119);
nand UO_3181 (O_3181,N_28717,N_28530);
nor UO_3182 (O_3182,N_28918,N_29231);
xor UO_3183 (O_3183,N_29975,N_28854);
or UO_3184 (O_3184,N_28914,N_29537);
nand UO_3185 (O_3185,N_29505,N_29003);
xnor UO_3186 (O_3186,N_29504,N_29673);
nand UO_3187 (O_3187,N_28879,N_29831);
nor UO_3188 (O_3188,N_28907,N_29290);
nand UO_3189 (O_3189,N_29527,N_29699);
or UO_3190 (O_3190,N_29892,N_28538);
xnor UO_3191 (O_3191,N_29640,N_28751);
nor UO_3192 (O_3192,N_28971,N_29339);
nor UO_3193 (O_3193,N_28763,N_29222);
nand UO_3194 (O_3194,N_28914,N_29769);
xor UO_3195 (O_3195,N_28557,N_28963);
or UO_3196 (O_3196,N_29267,N_28670);
xnor UO_3197 (O_3197,N_28907,N_29675);
or UO_3198 (O_3198,N_28752,N_29667);
nand UO_3199 (O_3199,N_28866,N_29578);
nand UO_3200 (O_3200,N_29565,N_29500);
or UO_3201 (O_3201,N_29941,N_29044);
and UO_3202 (O_3202,N_29970,N_29772);
nand UO_3203 (O_3203,N_29910,N_29081);
nand UO_3204 (O_3204,N_28873,N_29422);
xnor UO_3205 (O_3205,N_29434,N_28676);
and UO_3206 (O_3206,N_29980,N_28751);
nand UO_3207 (O_3207,N_29124,N_28696);
nor UO_3208 (O_3208,N_28979,N_29804);
nand UO_3209 (O_3209,N_29959,N_29338);
nand UO_3210 (O_3210,N_29504,N_29404);
or UO_3211 (O_3211,N_28794,N_29829);
nand UO_3212 (O_3212,N_29519,N_28869);
and UO_3213 (O_3213,N_28609,N_29511);
or UO_3214 (O_3214,N_28675,N_29144);
nor UO_3215 (O_3215,N_29498,N_29256);
and UO_3216 (O_3216,N_29723,N_28727);
or UO_3217 (O_3217,N_29230,N_29540);
and UO_3218 (O_3218,N_29036,N_29624);
nand UO_3219 (O_3219,N_29122,N_29564);
xnor UO_3220 (O_3220,N_28771,N_29788);
and UO_3221 (O_3221,N_29812,N_29932);
or UO_3222 (O_3222,N_29695,N_29246);
or UO_3223 (O_3223,N_29627,N_29546);
or UO_3224 (O_3224,N_28514,N_29525);
and UO_3225 (O_3225,N_29859,N_28759);
or UO_3226 (O_3226,N_29489,N_29683);
xnor UO_3227 (O_3227,N_29749,N_29563);
nor UO_3228 (O_3228,N_29686,N_29911);
or UO_3229 (O_3229,N_28717,N_28936);
or UO_3230 (O_3230,N_28577,N_29263);
nor UO_3231 (O_3231,N_29278,N_28710);
or UO_3232 (O_3232,N_28705,N_29179);
nor UO_3233 (O_3233,N_29062,N_29346);
xnor UO_3234 (O_3234,N_28695,N_28696);
and UO_3235 (O_3235,N_29734,N_28814);
or UO_3236 (O_3236,N_29996,N_28661);
or UO_3237 (O_3237,N_29063,N_28651);
xnor UO_3238 (O_3238,N_29157,N_28500);
and UO_3239 (O_3239,N_29903,N_29593);
or UO_3240 (O_3240,N_28502,N_28974);
nor UO_3241 (O_3241,N_29309,N_28869);
nor UO_3242 (O_3242,N_29513,N_28920);
or UO_3243 (O_3243,N_28812,N_29353);
nand UO_3244 (O_3244,N_29303,N_28655);
or UO_3245 (O_3245,N_29087,N_29925);
nor UO_3246 (O_3246,N_29754,N_28530);
xnor UO_3247 (O_3247,N_29564,N_29804);
and UO_3248 (O_3248,N_28918,N_29931);
or UO_3249 (O_3249,N_28688,N_29675);
xnor UO_3250 (O_3250,N_29844,N_29297);
nor UO_3251 (O_3251,N_29564,N_28910);
and UO_3252 (O_3252,N_29070,N_28994);
xor UO_3253 (O_3253,N_28560,N_28613);
nor UO_3254 (O_3254,N_28854,N_29449);
xor UO_3255 (O_3255,N_29039,N_29263);
and UO_3256 (O_3256,N_28762,N_29812);
xor UO_3257 (O_3257,N_28762,N_28511);
or UO_3258 (O_3258,N_29695,N_28565);
nor UO_3259 (O_3259,N_28896,N_28918);
and UO_3260 (O_3260,N_29520,N_29751);
nor UO_3261 (O_3261,N_29756,N_28533);
or UO_3262 (O_3262,N_29097,N_29762);
xor UO_3263 (O_3263,N_29438,N_29799);
or UO_3264 (O_3264,N_29682,N_28733);
xor UO_3265 (O_3265,N_28634,N_29568);
or UO_3266 (O_3266,N_29622,N_29252);
nor UO_3267 (O_3267,N_29373,N_28937);
nand UO_3268 (O_3268,N_29868,N_29010);
nor UO_3269 (O_3269,N_29644,N_28585);
xnor UO_3270 (O_3270,N_29434,N_28769);
nand UO_3271 (O_3271,N_29995,N_29512);
xor UO_3272 (O_3272,N_28892,N_28896);
nor UO_3273 (O_3273,N_28977,N_29849);
nand UO_3274 (O_3274,N_29748,N_29683);
nand UO_3275 (O_3275,N_29527,N_29482);
nor UO_3276 (O_3276,N_28812,N_29345);
xor UO_3277 (O_3277,N_28791,N_28678);
nand UO_3278 (O_3278,N_28909,N_29920);
xnor UO_3279 (O_3279,N_29805,N_28651);
nand UO_3280 (O_3280,N_29674,N_29964);
or UO_3281 (O_3281,N_29519,N_28561);
nand UO_3282 (O_3282,N_29812,N_28759);
nor UO_3283 (O_3283,N_28562,N_29177);
and UO_3284 (O_3284,N_29802,N_29998);
or UO_3285 (O_3285,N_29412,N_29041);
nor UO_3286 (O_3286,N_29566,N_29193);
or UO_3287 (O_3287,N_28687,N_29682);
or UO_3288 (O_3288,N_29334,N_29716);
or UO_3289 (O_3289,N_29450,N_28586);
nand UO_3290 (O_3290,N_28593,N_29658);
nor UO_3291 (O_3291,N_28981,N_28788);
and UO_3292 (O_3292,N_28805,N_29139);
and UO_3293 (O_3293,N_28846,N_29977);
xor UO_3294 (O_3294,N_29252,N_29436);
nand UO_3295 (O_3295,N_29502,N_28897);
nand UO_3296 (O_3296,N_29182,N_29794);
nand UO_3297 (O_3297,N_28876,N_29558);
nor UO_3298 (O_3298,N_29310,N_29843);
nor UO_3299 (O_3299,N_28584,N_28608);
and UO_3300 (O_3300,N_28954,N_29214);
or UO_3301 (O_3301,N_29940,N_29672);
nor UO_3302 (O_3302,N_28730,N_29757);
and UO_3303 (O_3303,N_28763,N_29427);
and UO_3304 (O_3304,N_29116,N_29293);
xnor UO_3305 (O_3305,N_29669,N_28874);
xor UO_3306 (O_3306,N_29620,N_29378);
xnor UO_3307 (O_3307,N_29442,N_29274);
and UO_3308 (O_3308,N_29261,N_29329);
and UO_3309 (O_3309,N_29678,N_29709);
nand UO_3310 (O_3310,N_29741,N_29898);
and UO_3311 (O_3311,N_29026,N_29545);
nand UO_3312 (O_3312,N_29891,N_28954);
nand UO_3313 (O_3313,N_29194,N_29706);
nor UO_3314 (O_3314,N_28812,N_28804);
or UO_3315 (O_3315,N_28792,N_29390);
or UO_3316 (O_3316,N_28945,N_29403);
nand UO_3317 (O_3317,N_29669,N_29904);
xnor UO_3318 (O_3318,N_29404,N_28858);
nand UO_3319 (O_3319,N_28839,N_29949);
or UO_3320 (O_3320,N_29618,N_29585);
nor UO_3321 (O_3321,N_29143,N_29462);
nor UO_3322 (O_3322,N_28888,N_29902);
nand UO_3323 (O_3323,N_29810,N_29355);
xnor UO_3324 (O_3324,N_29141,N_29500);
and UO_3325 (O_3325,N_29636,N_29437);
or UO_3326 (O_3326,N_29939,N_29126);
nor UO_3327 (O_3327,N_29093,N_28530);
nand UO_3328 (O_3328,N_29098,N_29569);
nand UO_3329 (O_3329,N_29965,N_29210);
xor UO_3330 (O_3330,N_29332,N_29902);
xnor UO_3331 (O_3331,N_29628,N_28533);
nor UO_3332 (O_3332,N_29895,N_29341);
and UO_3333 (O_3333,N_29239,N_28805);
xnor UO_3334 (O_3334,N_29450,N_29060);
and UO_3335 (O_3335,N_28850,N_28879);
nand UO_3336 (O_3336,N_29318,N_28555);
and UO_3337 (O_3337,N_28545,N_29658);
or UO_3338 (O_3338,N_29044,N_28536);
xor UO_3339 (O_3339,N_29801,N_29349);
nor UO_3340 (O_3340,N_29084,N_29008);
and UO_3341 (O_3341,N_29744,N_28509);
or UO_3342 (O_3342,N_28649,N_28830);
and UO_3343 (O_3343,N_28682,N_29000);
and UO_3344 (O_3344,N_28683,N_29094);
xnor UO_3345 (O_3345,N_28575,N_29530);
or UO_3346 (O_3346,N_29139,N_28643);
or UO_3347 (O_3347,N_29227,N_28676);
nor UO_3348 (O_3348,N_29052,N_29903);
xnor UO_3349 (O_3349,N_29491,N_29517);
and UO_3350 (O_3350,N_28713,N_28683);
and UO_3351 (O_3351,N_29412,N_29197);
xor UO_3352 (O_3352,N_28528,N_28801);
nor UO_3353 (O_3353,N_29007,N_28909);
xor UO_3354 (O_3354,N_29296,N_29999);
xor UO_3355 (O_3355,N_29616,N_29395);
nor UO_3356 (O_3356,N_29649,N_28866);
nand UO_3357 (O_3357,N_29172,N_29482);
or UO_3358 (O_3358,N_28871,N_29646);
nand UO_3359 (O_3359,N_29375,N_28525);
xnor UO_3360 (O_3360,N_29461,N_28798);
nor UO_3361 (O_3361,N_28608,N_28667);
xor UO_3362 (O_3362,N_29593,N_29867);
and UO_3363 (O_3363,N_29738,N_28860);
and UO_3364 (O_3364,N_28930,N_29934);
nand UO_3365 (O_3365,N_29444,N_29871);
nor UO_3366 (O_3366,N_28979,N_29456);
xnor UO_3367 (O_3367,N_28864,N_29316);
xor UO_3368 (O_3368,N_29657,N_29645);
nand UO_3369 (O_3369,N_28813,N_29228);
or UO_3370 (O_3370,N_28980,N_29106);
and UO_3371 (O_3371,N_28861,N_29262);
xor UO_3372 (O_3372,N_29788,N_28844);
xor UO_3373 (O_3373,N_29436,N_29439);
nor UO_3374 (O_3374,N_29333,N_29314);
and UO_3375 (O_3375,N_29842,N_29048);
nand UO_3376 (O_3376,N_28535,N_29727);
and UO_3377 (O_3377,N_29549,N_29449);
xnor UO_3378 (O_3378,N_29836,N_28699);
nor UO_3379 (O_3379,N_29950,N_28528);
or UO_3380 (O_3380,N_29766,N_28894);
nand UO_3381 (O_3381,N_29018,N_29466);
and UO_3382 (O_3382,N_28735,N_29007);
xor UO_3383 (O_3383,N_28725,N_28547);
and UO_3384 (O_3384,N_28898,N_28880);
nor UO_3385 (O_3385,N_28926,N_29277);
nand UO_3386 (O_3386,N_29572,N_28802);
nand UO_3387 (O_3387,N_28573,N_29086);
or UO_3388 (O_3388,N_29760,N_29546);
xor UO_3389 (O_3389,N_29809,N_29691);
nand UO_3390 (O_3390,N_28797,N_29622);
or UO_3391 (O_3391,N_29068,N_29565);
or UO_3392 (O_3392,N_29640,N_29541);
nand UO_3393 (O_3393,N_29206,N_29070);
nand UO_3394 (O_3394,N_29260,N_29504);
xor UO_3395 (O_3395,N_29605,N_28854);
xnor UO_3396 (O_3396,N_28579,N_29052);
xnor UO_3397 (O_3397,N_29264,N_28634);
nor UO_3398 (O_3398,N_28521,N_29234);
and UO_3399 (O_3399,N_29289,N_28971);
and UO_3400 (O_3400,N_28820,N_28595);
xnor UO_3401 (O_3401,N_29985,N_28791);
nor UO_3402 (O_3402,N_29827,N_29652);
and UO_3403 (O_3403,N_29211,N_28591);
nor UO_3404 (O_3404,N_28753,N_29693);
nor UO_3405 (O_3405,N_29370,N_29177);
nand UO_3406 (O_3406,N_28911,N_29826);
or UO_3407 (O_3407,N_29090,N_28770);
xor UO_3408 (O_3408,N_29178,N_29645);
nor UO_3409 (O_3409,N_28528,N_29673);
nor UO_3410 (O_3410,N_28532,N_29217);
xor UO_3411 (O_3411,N_29221,N_28733);
or UO_3412 (O_3412,N_29771,N_29517);
or UO_3413 (O_3413,N_29372,N_28723);
or UO_3414 (O_3414,N_28635,N_29319);
and UO_3415 (O_3415,N_28626,N_29385);
or UO_3416 (O_3416,N_29983,N_29607);
xnor UO_3417 (O_3417,N_29928,N_28879);
nor UO_3418 (O_3418,N_28786,N_29319);
xor UO_3419 (O_3419,N_29765,N_28714);
nor UO_3420 (O_3420,N_28800,N_28581);
nand UO_3421 (O_3421,N_29834,N_29364);
nand UO_3422 (O_3422,N_29554,N_29398);
or UO_3423 (O_3423,N_29021,N_29634);
and UO_3424 (O_3424,N_29302,N_28748);
xnor UO_3425 (O_3425,N_29118,N_29922);
and UO_3426 (O_3426,N_29972,N_28531);
and UO_3427 (O_3427,N_29961,N_29354);
or UO_3428 (O_3428,N_28822,N_29018);
or UO_3429 (O_3429,N_29244,N_28956);
nor UO_3430 (O_3430,N_28622,N_29877);
or UO_3431 (O_3431,N_28567,N_28713);
and UO_3432 (O_3432,N_29883,N_29493);
or UO_3433 (O_3433,N_29810,N_28721);
xor UO_3434 (O_3434,N_29266,N_29534);
and UO_3435 (O_3435,N_28704,N_29386);
xor UO_3436 (O_3436,N_28588,N_29165);
nand UO_3437 (O_3437,N_29782,N_28808);
or UO_3438 (O_3438,N_29863,N_29476);
nor UO_3439 (O_3439,N_28878,N_29865);
nor UO_3440 (O_3440,N_29331,N_29946);
and UO_3441 (O_3441,N_28732,N_28972);
or UO_3442 (O_3442,N_29142,N_29574);
and UO_3443 (O_3443,N_29436,N_28990);
nand UO_3444 (O_3444,N_29430,N_29691);
nand UO_3445 (O_3445,N_29689,N_29784);
nand UO_3446 (O_3446,N_29394,N_29383);
nor UO_3447 (O_3447,N_29188,N_29623);
or UO_3448 (O_3448,N_28629,N_29529);
xor UO_3449 (O_3449,N_28707,N_29833);
xnor UO_3450 (O_3450,N_29376,N_29054);
and UO_3451 (O_3451,N_29431,N_29848);
xor UO_3452 (O_3452,N_28898,N_28577);
nor UO_3453 (O_3453,N_28822,N_28617);
xor UO_3454 (O_3454,N_28969,N_29457);
nand UO_3455 (O_3455,N_29406,N_29846);
nor UO_3456 (O_3456,N_29765,N_29366);
and UO_3457 (O_3457,N_29724,N_29396);
nand UO_3458 (O_3458,N_28567,N_29912);
and UO_3459 (O_3459,N_28684,N_29046);
and UO_3460 (O_3460,N_28919,N_28700);
nand UO_3461 (O_3461,N_29248,N_28952);
nand UO_3462 (O_3462,N_29138,N_29609);
or UO_3463 (O_3463,N_28897,N_28660);
and UO_3464 (O_3464,N_28868,N_28912);
xnor UO_3465 (O_3465,N_28643,N_29070);
nand UO_3466 (O_3466,N_29216,N_29993);
nand UO_3467 (O_3467,N_28950,N_29493);
and UO_3468 (O_3468,N_29479,N_29249);
xnor UO_3469 (O_3469,N_29326,N_28666);
nand UO_3470 (O_3470,N_29258,N_29151);
or UO_3471 (O_3471,N_29803,N_28716);
nand UO_3472 (O_3472,N_29150,N_29946);
nand UO_3473 (O_3473,N_29238,N_29544);
xnor UO_3474 (O_3474,N_29426,N_29653);
and UO_3475 (O_3475,N_29595,N_29312);
or UO_3476 (O_3476,N_29271,N_29273);
xor UO_3477 (O_3477,N_29841,N_29846);
nand UO_3478 (O_3478,N_29916,N_29885);
xor UO_3479 (O_3479,N_29868,N_28579);
and UO_3480 (O_3480,N_28756,N_29199);
xnor UO_3481 (O_3481,N_29587,N_29347);
or UO_3482 (O_3482,N_29916,N_29498);
xnor UO_3483 (O_3483,N_29439,N_29445);
xnor UO_3484 (O_3484,N_28515,N_28807);
nor UO_3485 (O_3485,N_29688,N_29300);
and UO_3486 (O_3486,N_28792,N_29899);
xor UO_3487 (O_3487,N_29747,N_29678);
and UO_3488 (O_3488,N_29228,N_29283);
nand UO_3489 (O_3489,N_29733,N_28805);
or UO_3490 (O_3490,N_28755,N_29592);
nand UO_3491 (O_3491,N_29401,N_28576);
or UO_3492 (O_3492,N_29525,N_29885);
xor UO_3493 (O_3493,N_29631,N_29648);
or UO_3494 (O_3494,N_28751,N_29982);
nand UO_3495 (O_3495,N_28918,N_29074);
nor UO_3496 (O_3496,N_28815,N_29139);
xnor UO_3497 (O_3497,N_28788,N_29516);
xor UO_3498 (O_3498,N_29627,N_29265);
nor UO_3499 (O_3499,N_29735,N_29484);
endmodule