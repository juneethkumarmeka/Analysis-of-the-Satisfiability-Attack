module basic_3000_30000_3500_25_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
and U0 (N_0,In_1012,In_2596);
nor U1 (N_1,In_2470,In_1126);
nor U2 (N_2,In_425,In_1317);
or U3 (N_3,In_433,In_1952);
nand U4 (N_4,In_2809,In_202);
or U5 (N_5,In_60,In_364);
xnor U6 (N_6,In_343,In_2553);
nor U7 (N_7,In_20,In_1459);
nand U8 (N_8,In_2451,In_1139);
xor U9 (N_9,In_824,In_1706);
and U10 (N_10,In_352,In_1632);
and U11 (N_11,In_1556,In_536);
and U12 (N_12,In_2731,In_1691);
xnor U13 (N_13,In_505,In_2964);
and U14 (N_14,In_1409,In_707);
and U15 (N_15,In_1599,In_2317);
or U16 (N_16,In_2562,In_658);
nor U17 (N_17,In_2131,In_2225);
or U18 (N_18,In_1526,In_1291);
xnor U19 (N_19,In_78,In_2036);
nor U20 (N_20,In_388,In_926);
nor U21 (N_21,In_937,In_1513);
xor U22 (N_22,In_2408,In_1813);
nand U23 (N_23,In_2091,In_1949);
xor U24 (N_24,In_142,In_633);
or U25 (N_25,In_448,In_1715);
nor U26 (N_26,In_1087,In_538);
and U27 (N_27,In_1730,In_2968);
nand U28 (N_28,In_28,In_1580);
xnor U29 (N_29,In_1907,In_1314);
nor U30 (N_30,In_1649,In_999);
nor U31 (N_31,In_1812,In_2815);
nor U32 (N_32,In_506,In_831);
xor U33 (N_33,In_544,In_2838);
nand U34 (N_34,In_2659,In_1720);
nand U35 (N_35,In_71,In_1829);
or U36 (N_36,In_2276,In_2593);
xnor U37 (N_37,In_1563,In_2250);
xor U38 (N_38,In_1711,In_981);
or U39 (N_39,In_1175,In_1413);
or U40 (N_40,In_1230,In_1477);
or U41 (N_41,In_1024,In_1849);
xnor U42 (N_42,In_1955,In_1495);
nor U43 (N_43,In_1609,In_2613);
or U44 (N_44,In_603,In_2241);
nand U45 (N_45,In_684,In_2874);
or U46 (N_46,In_1861,In_468);
nand U47 (N_47,In_2146,In_2827);
or U48 (N_48,In_2464,In_1075);
or U49 (N_49,In_222,In_488);
or U50 (N_50,In_106,In_1132);
nand U51 (N_51,In_2935,In_1886);
nor U52 (N_52,In_2009,In_2712);
and U53 (N_53,In_313,In_457);
and U54 (N_54,In_769,In_311);
and U55 (N_55,In_1005,In_455);
and U56 (N_56,In_1496,In_1173);
or U57 (N_57,In_2875,In_2352);
xnor U58 (N_58,In_366,In_2298);
nand U59 (N_59,In_1925,In_2488);
xnor U60 (N_60,In_569,In_263);
xnor U61 (N_61,In_1480,In_2567);
nor U62 (N_62,In_2856,In_80);
nor U63 (N_63,In_2386,In_2524);
xor U64 (N_64,In_1362,In_733);
nand U65 (N_65,In_1148,In_445);
and U66 (N_66,In_1670,In_694);
or U67 (N_67,In_1214,In_2042);
and U68 (N_68,In_1555,In_189);
and U69 (N_69,In_1160,In_1636);
nand U70 (N_70,In_2020,In_51);
or U71 (N_71,In_1524,In_2228);
nand U72 (N_72,In_1252,In_721);
and U73 (N_73,In_2871,In_2019);
nand U74 (N_74,In_2118,In_330);
and U75 (N_75,In_1419,In_1961);
or U76 (N_76,In_3,In_1177);
nor U77 (N_77,In_2061,In_868);
and U78 (N_78,In_107,In_1327);
nand U79 (N_79,In_643,In_1666);
or U80 (N_80,In_262,In_1509);
nand U81 (N_81,In_551,In_1656);
and U82 (N_82,In_2765,In_486);
and U83 (N_83,In_2672,In_2989);
xnor U84 (N_84,In_323,In_989);
xor U85 (N_85,In_2975,In_577);
and U86 (N_86,In_1262,In_594);
nor U87 (N_87,In_1390,In_2919);
nand U88 (N_88,In_1144,In_2259);
xnor U89 (N_89,In_2961,In_37);
and U90 (N_90,In_2040,In_676);
nand U91 (N_91,In_2338,In_776);
nor U92 (N_92,In_392,In_2550);
or U93 (N_93,In_2291,In_251);
and U94 (N_94,In_2954,In_1470);
or U95 (N_95,In_639,In_1533);
or U96 (N_96,In_1653,In_714);
nor U97 (N_97,In_2478,In_545);
nand U98 (N_98,In_988,In_2175);
or U99 (N_99,In_645,In_1371);
and U100 (N_100,In_1518,In_480);
or U101 (N_101,In_914,In_1573);
and U102 (N_102,In_2165,In_2667);
xnor U103 (N_103,In_2437,In_229);
nand U104 (N_104,In_1796,In_2327);
xor U105 (N_105,In_124,In_960);
nand U106 (N_106,In_1931,In_2139);
and U107 (N_107,In_2158,In_1425);
nor U108 (N_108,In_2491,In_1777);
nand U109 (N_109,In_165,In_2654);
nand U110 (N_110,In_956,In_1800);
and U111 (N_111,In_2407,In_2400);
or U112 (N_112,In_2404,In_2329);
nand U113 (N_113,In_1932,In_1919);
nand U114 (N_114,In_1402,In_784);
xor U115 (N_115,In_1866,In_2472);
and U116 (N_116,In_895,In_159);
nor U117 (N_117,In_504,In_2958);
nor U118 (N_118,In_365,In_2280);
nand U119 (N_119,In_1911,In_2173);
or U120 (N_120,In_257,In_68);
nor U121 (N_121,In_2963,In_2744);
nand U122 (N_122,In_1780,In_1523);
or U123 (N_123,In_2354,In_2418);
xnor U124 (N_124,In_295,In_377);
nand U125 (N_125,In_958,In_834);
xnor U126 (N_126,In_12,In_414);
nand U127 (N_127,In_192,In_2434);
and U128 (N_128,In_79,In_2249);
nor U129 (N_129,In_2232,In_1123);
xor U130 (N_130,In_617,In_2342);
xor U131 (N_131,In_781,In_111);
xnor U132 (N_132,In_1452,In_1428);
nor U133 (N_133,In_2145,In_1850);
nor U134 (N_134,In_1584,In_94);
xnor U135 (N_135,In_1156,In_2784);
or U136 (N_136,In_510,In_614);
xor U137 (N_137,In_1909,In_2599);
and U138 (N_138,In_2920,In_1270);
or U139 (N_139,In_2068,In_2864);
nor U140 (N_140,In_410,In_1388);
and U141 (N_141,In_1628,In_2912);
or U142 (N_142,In_2001,In_1340);
nand U143 (N_143,In_289,In_2150);
or U144 (N_144,In_1544,In_2906);
and U145 (N_145,In_867,In_1629);
xor U146 (N_146,In_2051,In_1195);
or U147 (N_147,In_660,In_2515);
and U148 (N_148,In_400,In_1115);
nand U149 (N_149,In_2527,In_2032);
and U150 (N_150,In_794,In_44);
xnor U151 (N_151,In_268,In_2718);
and U152 (N_152,In_344,In_25);
nor U153 (N_153,In_767,In_1970);
xor U154 (N_154,In_1639,In_2284);
nor U155 (N_155,In_2835,In_135);
or U156 (N_156,In_1983,In_1664);
nor U157 (N_157,In_663,In_523);
and U158 (N_158,In_2081,In_2587);
nand U159 (N_159,In_147,In_2083);
nor U160 (N_160,In_1254,In_487);
xnor U161 (N_161,In_1121,In_2626);
and U162 (N_162,In_6,In_2096);
xnor U163 (N_163,In_2569,In_2710);
or U164 (N_164,In_2701,In_860);
or U165 (N_165,In_1166,In_496);
xor U166 (N_166,In_217,In_2349);
and U167 (N_167,In_2192,In_1529);
or U168 (N_168,In_314,In_819);
xor U169 (N_169,In_2714,In_1681);
xnor U170 (N_170,In_2277,In_1086);
or U171 (N_171,In_2104,In_2444);
nand U172 (N_172,In_1065,In_945);
and U173 (N_173,In_1978,In_1015);
nand U174 (N_174,In_2006,In_149);
or U175 (N_175,In_665,In_898);
nand U176 (N_176,In_1038,In_167);
nand U177 (N_177,In_1228,In_59);
nand U178 (N_178,In_34,In_1076);
nor U179 (N_179,In_1511,In_1378);
and U180 (N_180,In_2431,In_2373);
nor U181 (N_181,In_650,In_1267);
xnor U182 (N_182,In_611,In_2521);
nand U183 (N_183,In_140,In_1635);
and U184 (N_184,In_1348,In_1458);
nand U185 (N_185,In_1683,In_292);
xor U186 (N_186,In_264,In_1747);
nand U187 (N_187,In_1082,In_2293);
nor U188 (N_188,In_1958,In_965);
and U189 (N_189,In_2558,In_2829);
nand U190 (N_190,In_1892,In_2732);
nor U191 (N_191,In_690,In_2043);
and U192 (N_192,In_948,In_765);
or U193 (N_193,In_472,In_2119);
nor U194 (N_194,In_2087,In_2579);
nand U195 (N_195,In_105,In_494);
or U196 (N_196,In_1610,In_1534);
and U197 (N_197,In_2870,In_308);
and U198 (N_198,In_52,In_1028);
or U199 (N_199,In_2676,In_342);
nor U200 (N_200,In_2059,In_2965);
nor U201 (N_201,In_1724,In_2614);
and U202 (N_202,In_1827,In_1366);
nor U203 (N_203,In_1149,In_351);
xor U204 (N_204,In_1631,In_1094);
xnor U205 (N_205,In_288,In_282);
nand U206 (N_206,In_119,In_1306);
nor U207 (N_207,In_728,In_1017);
xor U208 (N_208,In_230,In_1997);
and U209 (N_209,In_1570,In_2541);
and U210 (N_210,In_276,In_334);
or U211 (N_211,In_2566,In_1799);
nor U212 (N_212,In_1441,In_373);
xor U213 (N_213,In_1238,In_2411);
or U214 (N_214,In_1862,In_2722);
or U215 (N_215,In_2024,In_384);
nand U216 (N_216,In_2790,In_2759);
and U217 (N_217,In_1844,In_1297);
xnor U218 (N_218,In_1290,In_408);
and U219 (N_219,In_2755,In_1307);
nor U220 (N_220,In_2600,In_2687);
nor U221 (N_221,In_387,In_980);
or U222 (N_222,In_2883,In_1321);
nand U223 (N_223,In_1543,In_2719);
xor U224 (N_224,In_1232,In_533);
xnor U225 (N_225,In_1237,In_502);
xor U226 (N_226,In_451,In_1727);
or U227 (N_227,In_8,In_2302);
nand U228 (N_228,In_1426,In_2267);
nand U229 (N_229,In_889,In_768);
or U230 (N_230,In_371,In_2092);
xnor U231 (N_231,In_2559,In_874);
xnor U232 (N_232,In_2988,In_1257);
or U233 (N_233,In_1700,In_574);
xor U234 (N_234,In_1220,In_2505);
nor U235 (N_235,In_137,In_2756);
xor U236 (N_236,In_2084,In_876);
xor U237 (N_237,In_69,In_1045);
or U238 (N_238,In_994,In_2742);
or U239 (N_239,In_1400,In_162);
xor U240 (N_240,In_998,In_7);
or U241 (N_241,In_2943,In_1179);
nor U242 (N_242,In_522,In_2760);
nor U243 (N_243,In_205,In_2052);
and U244 (N_244,In_2178,In_2598);
nor U245 (N_245,In_207,In_1743);
or U246 (N_246,In_1295,In_1790);
or U247 (N_247,In_1036,In_1326);
nand U248 (N_248,In_169,In_1097);
xor U249 (N_249,In_2448,In_1926);
and U250 (N_250,In_1155,In_1697);
or U251 (N_251,In_1644,In_2575);
nor U252 (N_252,In_1616,In_1938);
or U253 (N_253,In_1746,In_420);
and U254 (N_254,In_1410,In_1190);
nand U255 (N_255,In_789,In_1093);
or U256 (N_256,In_2154,In_2849);
or U257 (N_257,In_2612,In_2057);
nor U258 (N_258,In_286,In_422);
nand U259 (N_259,In_2269,In_578);
xnor U260 (N_260,In_1916,In_1084);
xor U261 (N_261,In_2427,In_1211);
nor U262 (N_262,In_771,In_2738);
nand U263 (N_263,In_67,In_2876);
nor U264 (N_264,In_2463,In_2322);
xor U265 (N_265,In_791,In_1007);
xnor U266 (N_266,In_2435,In_442);
or U267 (N_267,In_426,In_716);
and U268 (N_268,In_1025,In_1948);
xor U269 (N_269,In_235,In_1192);
and U270 (N_270,In_877,In_2877);
xnor U271 (N_271,In_2243,In_2275);
and U272 (N_272,In_2247,In_1551);
or U273 (N_273,In_1180,In_2980);
and U274 (N_274,In_2683,In_2905);
nor U275 (N_275,In_2405,In_531);
nor U276 (N_276,In_1993,In_1201);
nand U277 (N_277,In_2823,In_1826);
nor U278 (N_278,In_918,In_1310);
or U279 (N_279,In_2737,In_1112);
nor U280 (N_280,In_2328,In_829);
nor U281 (N_281,In_627,In_326);
or U282 (N_282,In_2027,In_1448);
or U283 (N_283,In_1022,In_2697);
and U284 (N_284,In_711,In_842);
or U285 (N_285,In_1251,In_1331);
or U286 (N_286,In_1437,In_823);
or U287 (N_287,In_2851,In_528);
xor U288 (N_288,In_1501,In_1601);
xor U289 (N_289,In_1839,In_109);
or U290 (N_290,In_409,In_1595);
nor U291 (N_291,In_1131,In_2998);
nor U292 (N_292,In_598,In_2359);
xor U293 (N_293,In_150,In_2806);
nor U294 (N_294,In_2333,In_2378);
and U295 (N_295,In_2462,In_1225);
or U296 (N_296,In_2113,In_766);
or U297 (N_297,In_2079,In_2611);
and U298 (N_298,In_2071,In_2987);
nand U299 (N_299,In_979,In_1871);
nand U300 (N_300,In_1651,In_1941);
nor U301 (N_301,In_1991,In_1966);
xnor U302 (N_302,In_1316,In_2666);
xor U303 (N_303,In_353,In_1538);
nand U304 (N_304,In_117,In_462);
xnor U305 (N_305,In_1749,In_2054);
nor U306 (N_306,In_53,In_1301);
and U307 (N_307,In_2376,In_1185);
nor U308 (N_308,In_717,In_1944);
nand U309 (N_309,In_924,In_640);
and U310 (N_310,In_1673,In_2021);
xnor U311 (N_311,In_724,In_2257);
xnor U312 (N_312,In_2771,In_2326);
xnor U313 (N_313,In_1578,In_570);
or U314 (N_314,In_2179,In_2481);
or U315 (N_315,In_13,In_2775);
and U316 (N_316,In_1264,In_491);
nand U317 (N_317,In_513,In_1935);
nand U318 (N_318,In_1519,In_411);
nand U319 (N_319,In_1210,In_1078);
nor U320 (N_320,In_2907,In_729);
xor U321 (N_321,In_1176,In_2459);
nor U322 (N_322,In_2752,In_1728);
nand U323 (N_323,In_2708,In_2690);
xor U324 (N_324,In_1939,In_73);
xnor U325 (N_325,In_940,In_1748);
nand U326 (N_326,In_1379,In_1924);
and U327 (N_327,In_2533,In_530);
nor U328 (N_328,In_2741,In_1263);
and U329 (N_329,In_861,In_2453);
and U330 (N_330,In_2060,In_2450);
and U331 (N_331,In_2604,In_1053);
nand U332 (N_332,In_1494,In_2502);
or U333 (N_333,In_1250,In_332);
nor U334 (N_334,In_1994,In_1215);
and U335 (N_335,In_753,In_291);
nor U336 (N_336,In_1980,In_703);
and U337 (N_337,In_243,In_112);
xnor U338 (N_338,In_622,In_559);
xor U339 (N_339,In_2078,In_403);
nand U340 (N_340,In_1268,In_2547);
nor U341 (N_341,In_1350,In_904);
and U342 (N_342,In_2381,In_281);
nand U343 (N_343,In_1421,In_1286);
nor U344 (N_344,In_2107,In_816);
and U345 (N_345,In_585,In_1424);
nor U346 (N_346,In_1479,In_83);
nand U347 (N_347,In_1877,In_969);
and U348 (N_348,In_2970,In_2215);
and U349 (N_349,In_674,In_1404);
or U350 (N_350,In_2540,In_290);
or U351 (N_351,In_2424,In_2205);
or U352 (N_352,In_2216,In_554);
xnor U353 (N_353,In_1873,In_278);
and U354 (N_354,In_63,In_1565);
nor U355 (N_355,In_1446,In_413);
xnor U356 (N_356,In_2955,In_2772);
nand U357 (N_357,In_1200,In_1946);
xnor U358 (N_358,In_2630,In_550);
nor U359 (N_359,In_2642,In_2563);
nor U360 (N_360,In_1129,In_2446);
nand U361 (N_361,In_484,In_120);
nand U362 (N_362,In_595,In_685);
nand U363 (N_363,In_540,In_1856);
nor U364 (N_364,In_1193,In_2461);
and U365 (N_365,In_1240,In_2747);
nor U366 (N_366,In_11,In_563);
xnor U367 (N_367,In_240,In_1751);
xnor U368 (N_368,In_1592,In_1823);
or U369 (N_369,In_1559,In_1761);
or U370 (N_370,In_1408,In_896);
xor U371 (N_371,In_1898,In_252);
nor U372 (N_372,In_1789,In_1619);
nor U373 (N_373,In_2285,In_1450);
and U374 (N_374,In_453,In_1779);
and U375 (N_375,In_199,In_1169);
and U376 (N_376,In_1389,In_1550);
nand U377 (N_377,In_1642,In_815);
nor U378 (N_378,In_133,In_709);
and U379 (N_379,In_2582,In_2425);
xor U380 (N_380,In_1589,In_1540);
and U381 (N_381,In_2555,In_2231);
nor U382 (N_382,In_744,In_1539);
nand U383 (N_383,In_1521,In_2572);
xnor U384 (N_384,In_1217,In_1344);
or U385 (N_385,In_2049,In_656);
and U386 (N_386,In_1324,In_499);
or U387 (N_387,In_1954,In_1285);
or U388 (N_388,In_2236,In_1641);
xor U389 (N_389,In_2251,In_2615);
nor U390 (N_390,In_628,In_2886);
nand U391 (N_391,In_2884,In_638);
nand U392 (N_392,In_1895,In_1760);
and U393 (N_393,In_2286,In_1708);
xor U394 (N_394,In_1449,In_2270);
nor U395 (N_395,In_1066,In_936);
nand U396 (N_396,In_2689,In_1034);
nand U397 (N_397,In_2220,In_2416);
nand U398 (N_398,In_2069,In_1178);
or U399 (N_399,In_2273,In_725);
nand U400 (N_400,In_1026,In_62);
xor U401 (N_401,In_2012,In_212);
xor U402 (N_402,In_474,In_1655);
or U403 (N_403,In_2176,In_427);
or U404 (N_404,In_1890,In_2723);
xor U405 (N_405,In_2029,In_280);
xnor U406 (N_406,In_385,In_1973);
and U407 (N_407,In_1633,In_2106);
nor U408 (N_408,In_1884,In_1041);
xor U409 (N_409,In_1814,In_1834);
nand U410 (N_410,In_2500,In_183);
and U411 (N_411,In_2341,In_534);
or U412 (N_412,In_1933,In_2413);
and U413 (N_413,In_2254,In_2063);
and U414 (N_414,In_503,In_1957);
nor U415 (N_415,In_798,In_700);
xnor U416 (N_416,In_302,In_2217);
nand U417 (N_417,In_943,In_1863);
xnor U418 (N_418,In_1434,In_1279);
nor U419 (N_419,In_2831,In_2584);
or U420 (N_420,In_587,In_1569);
nor U421 (N_421,In_2925,In_2332);
nand U422 (N_422,In_2788,In_697);
nand U423 (N_423,In_1382,In_284);
nor U424 (N_424,In_1657,In_2423);
nand U425 (N_425,In_1491,In_779);
or U426 (N_426,In_2163,In_1908);
or U427 (N_427,In_1598,In_2388);
nor U428 (N_428,In_87,In_1956);
and U429 (N_429,In_1549,In_1902);
and U430 (N_430,In_2229,In_2312);
nand U431 (N_431,In_2945,In_2570);
and U432 (N_432,In_754,In_1774);
nand U433 (N_433,In_1186,In_2415);
xnor U434 (N_434,In_1373,In_2014);
xnor U435 (N_435,In_1968,In_1794);
nor U436 (N_436,In_748,In_1455);
and U437 (N_437,In_607,In_95);
nand U438 (N_438,In_2658,In_2819);
xnor U439 (N_439,In_2585,In_2896);
or U440 (N_440,In_2634,In_1090);
nand U441 (N_441,In_1158,In_2565);
or U442 (N_442,In_2868,In_1581);
xor U443 (N_443,In_613,In_362);
nor U444 (N_444,In_1484,In_2393);
xnor U445 (N_445,In_2255,In_2962);
or U446 (N_446,In_838,In_2223);
nor U447 (N_447,In_2169,In_2366);
nor U448 (N_448,In_2136,In_2580);
nand U449 (N_449,In_1342,In_2350);
or U450 (N_450,In_1386,In_256);
and U451 (N_451,In_430,In_2080);
nor U452 (N_452,In_1880,In_2123);
nor U453 (N_453,In_953,In_1611);
xor U454 (N_454,In_26,In_210);
and U455 (N_455,In_1021,In_884);
nor U456 (N_456,In_1744,In_1457);
and U457 (N_457,In_2132,In_2159);
nand U458 (N_458,In_325,In_2624);
nor U459 (N_459,In_1236,In_865);
or U460 (N_460,In_75,In_1397);
xnor U461 (N_461,In_565,In_952);
and U462 (N_462,In_2960,In_2351);
and U463 (N_463,In_85,In_880);
nand U464 (N_464,In_220,In_655);
or U465 (N_465,In_1051,In_987);
and U466 (N_466,In_1292,In_116);
nand U467 (N_467,In_2053,In_1689);
nor U468 (N_468,In_1204,In_1652);
or U469 (N_469,In_1050,In_1912);
nor U470 (N_470,In_546,In_1772);
or U471 (N_471,In_1614,In_2991);
or U472 (N_472,In_661,In_1124);
nand U473 (N_473,In_938,In_2959);
nor U474 (N_474,In_1802,In_1695);
and U475 (N_475,In_2631,In_340);
nor U476 (N_476,In_172,In_481);
nor U477 (N_477,In_158,In_2357);
or U478 (N_478,In_187,In_1412);
and U479 (N_479,In_871,In_1564);
nor U480 (N_480,In_2937,In_156);
and U481 (N_481,In_1665,In_2863);
xor U482 (N_482,In_2300,In_1183);
nor U483 (N_483,In_1859,In_592);
nand U484 (N_484,In_2361,In_375);
xor U485 (N_485,In_1558,In_2212);
and U486 (N_486,In_1816,In_2953);
or U487 (N_487,In_1338,In_141);
nor U488 (N_488,In_1767,In_33);
xnor U489 (N_489,In_378,In_2);
nand U490 (N_490,In_803,In_2544);
nand U491 (N_491,In_2705,In_2665);
or U492 (N_492,In_84,In_1977);
nand U493 (N_493,In_1756,In_2619);
nor U494 (N_494,In_687,In_2385);
nand U495 (N_495,In_456,In_2733);
xnor U496 (N_496,In_2686,In_1913);
nand U497 (N_497,In_2841,In_1466);
nor U498 (N_498,In_2675,In_2836);
nand U499 (N_499,In_588,In_2454);
nand U500 (N_500,In_933,In_21);
and U501 (N_501,In_1209,In_347);
xnor U502 (N_502,In_317,In_1133);
and U503 (N_503,In_294,In_1253);
or U504 (N_504,In_778,In_2694);
nand U505 (N_505,In_2153,In_299);
nand U506 (N_506,In_2813,In_283);
and U507 (N_507,In_495,In_1394);
nor U508 (N_508,In_699,In_1414);
nor U509 (N_509,In_320,In_215);
nand U510 (N_510,In_2143,In_2939);
nand U511 (N_511,In_2785,In_2184);
xor U512 (N_512,In_1337,In_2782);
or U513 (N_513,In_1303,In_782);
and U514 (N_514,In_1246,In_2993);
or U515 (N_515,In_2487,In_103);
or U516 (N_516,In_2893,In_848);
nor U517 (N_517,In_27,In_2356);
and U518 (N_518,In_1537,In_736);
and U519 (N_519,In_678,In_1415);
and U520 (N_520,In_1300,In_2278);
nand U521 (N_521,In_1891,In_482);
or U522 (N_522,In_1737,In_2601);
nand U523 (N_523,In_1258,In_2325);
or U524 (N_524,In_600,In_2039);
nor U525 (N_525,In_1505,In_657);
or U526 (N_526,In_1759,In_2010);
nor U527 (N_527,In_507,In_449);
or U528 (N_528,In_1853,In_99);
or U529 (N_529,In_2637,In_2130);
nand U530 (N_530,In_1369,In_2469);
and U531 (N_531,In_1016,In_529);
xor U532 (N_532,In_2607,In_1679);
nor U533 (N_533,In_321,In_128);
and U534 (N_534,In_1702,In_393);
and U535 (N_535,In_424,In_389);
and U536 (N_536,In_127,In_1284);
nor U537 (N_537,In_376,In_727);
and U538 (N_538,In_248,In_1515);
nand U539 (N_539,In_2114,In_1318);
xor U540 (N_540,In_2258,In_2412);
nand U541 (N_541,In_901,In_2290);
or U542 (N_542,In_2064,In_2193);
nor U543 (N_543,In_1161,In_1398);
xor U544 (N_544,In_1194,In_993);
and U545 (N_545,In_1343,In_2272);
or U546 (N_546,In_270,In_2616);
xor U547 (N_547,In_1566,In_1810);
xor U548 (N_548,In_2292,In_810);
nor U549 (N_549,In_1889,In_2888);
and U550 (N_550,In_2516,In_897);
xor U551 (N_551,In_1623,In_1848);
nor U552 (N_552,In_1803,In_2717);
nand U553 (N_553,In_1287,In_2307);
and U554 (N_554,In_108,In_992);
or U555 (N_555,In_2147,In_2869);
xor U556 (N_556,In_1381,In_1153);
nor U557 (N_557,In_1499,In_1781);
or U558 (N_558,In_2832,In_2045);
xnor U559 (N_559,In_1127,In_1921);
and U560 (N_560,In_1981,In_370);
and U561 (N_561,In_1739,In_372);
or U562 (N_562,In_1778,In_2828);
xnor U563 (N_563,In_226,In_2735);
xnor U564 (N_564,In_1039,In_1710);
or U565 (N_565,In_864,In_1847);
and U566 (N_566,In_2026,In_331);
nand U567 (N_567,In_882,In_1478);
nand U568 (N_568,In_1103,In_2798);
nor U569 (N_569,In_2000,In_760);
nand U570 (N_570,In_1120,In_548);
nor U571 (N_571,In_517,In_1219);
nand U572 (N_572,In_206,In_1137);
or U573 (N_573,In_1741,In_245);
and U574 (N_574,In_177,In_1585);
nand U575 (N_575,In_2213,In_333);
and U576 (N_576,In_1135,In_648);
or U577 (N_577,In_968,In_2695);
nor U578 (N_578,In_1048,In_2882);
nor U579 (N_579,In_1661,In_742);
xnor U580 (N_580,In_2996,In_1191);
or U581 (N_581,In_1420,In_675);
and U582 (N_582,In_1792,In_2237);
or U583 (N_583,In_886,In_1299);
or U584 (N_584,In_909,In_2878);
nand U585 (N_585,In_1881,In_2432);
nand U586 (N_586,In_1032,In_1722);
nand U587 (N_587,In_2923,In_912);
nand U588 (N_588,In_2934,In_143);
nand U589 (N_589,In_827,In_2323);
nand U590 (N_590,In_2265,In_1463);
and U591 (N_591,In_1199,In_2129);
nand U592 (N_592,In_817,In_2844);
nor U593 (N_593,In_2852,In_698);
xnor U594 (N_594,In_2618,In_2640);
nand U595 (N_595,In_878,In_2363);
nand U596 (N_596,In_1031,In_888);
nor U597 (N_597,In_2535,In_2439);
and U598 (N_598,In_1358,In_2921);
nor U599 (N_599,In_2668,In_1352);
and U600 (N_600,In_790,In_310);
or U601 (N_601,In_1712,In_1060);
xnor U602 (N_602,In_1858,In_208);
xor U603 (N_603,In_1485,In_2873);
xnor U604 (N_604,In_242,In_361);
nand U605 (N_605,In_1527,In_2507);
xor U606 (N_606,In_632,In_218);
or U607 (N_607,In_795,In_2620);
or U608 (N_608,In_2670,In_807);
nor U609 (N_609,In_931,In_2916);
xnor U610 (N_610,In_303,In_305);
and U611 (N_611,In_2810,In_2940);
or U612 (N_612,In_1332,In_2680);
xnor U613 (N_613,In_14,In_2409);
xor U614 (N_614,In_1542,In_88);
nand U615 (N_615,In_136,In_1234);
nor U616 (N_616,In_1920,In_1869);
nand U617 (N_617,In_836,In_421);
nor U618 (N_618,In_2930,In_804);
nor U619 (N_619,In_1502,In_1080);
and U620 (N_620,In_2606,In_862);
xor U621 (N_621,In_1857,In_1018);
nand U622 (N_622,In_511,In_144);
or U623 (N_623,In_843,In_1092);
or U624 (N_624,In_1675,In_1713);
xor U625 (N_625,In_1998,In_1701);
nand U626 (N_626,In_2070,In_1714);
xnor U627 (N_627,In_1828,In_2804);
xnor U628 (N_628,In_1198,In_2944);
nor U629 (N_629,In_346,In_1807);
nor U630 (N_630,In_2443,In_1647);
xnor U631 (N_631,In_2037,In_1359);
and U632 (N_632,In_1298,In_2304);
xnor U633 (N_633,In_234,In_2008);
or U634 (N_634,In_35,In_173);
nor U635 (N_635,In_1383,In_852);
nand U636 (N_636,In_2282,In_471);
nor U637 (N_637,In_2651,In_191);
and U638 (N_638,In_597,In_2344);
or U639 (N_639,In_715,In_2075);
nand U640 (N_640,In_2414,In_2142);
nand U641 (N_641,In_605,In_2834);
nand U642 (N_642,In_1182,In_2936);
nor U643 (N_643,In_2713,In_443);
nor U644 (N_644,In_2149,In_1662);
xnor U645 (N_645,In_1927,In_2379);
and U646 (N_646,In_1406,In_1081);
nand U647 (N_647,In_812,In_2949);
and U648 (N_648,In_2514,In_1213);
and U649 (N_649,In_825,In_254);
or U650 (N_650,In_386,In_1498);
and U651 (N_651,In_561,In_950);
xnor U652 (N_652,In_2401,In_826);
nand U653 (N_653,In_2981,In_2209);
and U654 (N_654,In_1669,In_1787);
nand U655 (N_655,In_2047,In_2183);
and U656 (N_656,In_1953,In_2525);
and U657 (N_657,In_2560,In_271);
and U658 (N_658,In_2471,In_1615);
nand U659 (N_659,In_2479,In_1357);
or U660 (N_660,In_1841,In_2763);
xor U661 (N_661,In_70,In_2495);
xor U662 (N_662,In_923,In_647);
or U663 (N_663,In_2120,In_2296);
and U664 (N_664,In_66,In_2156);
nand U665 (N_665,In_747,In_1878);
nand U666 (N_666,In_1736,In_1308);
nand U667 (N_667,In_602,In_2779);
xor U668 (N_668,In_1377,In_830);
and U669 (N_669,In_2458,In_2984);
xnor U670 (N_670,In_2198,In_1830);
nor U671 (N_671,In_2610,In_2133);
or U672 (N_672,In_2764,In_957);
nor U673 (N_673,In_297,In_2554);
xnor U674 (N_674,In_2486,In_2861);
xnor U675 (N_675,In_2546,In_350);
and U676 (N_676,In_2090,In_1506);
or U677 (N_677,In_1842,In_1208);
xor U678 (N_678,In_97,In_2028);
and U679 (N_679,In_2808,In_1003);
and U680 (N_680,In_2551,In_2498);
or U681 (N_681,In_1947,In_1872);
or U682 (N_682,In_1259,In_1845);
or U683 (N_683,In_2857,In_1899);
nor U684 (N_684,In_2167,In_19);
xnor U685 (N_685,In_844,In_906);
xor U686 (N_686,In_2002,In_2324);
or U687 (N_687,In_2484,In_535);
nand U688 (N_688,In_318,In_1427);
xnor U689 (N_689,In_1432,In_821);
or U690 (N_690,In_2181,In_2824);
or U691 (N_691,In_2306,In_1995);
or U692 (N_692,In_1687,In_179);
xor U693 (N_693,In_1030,In_802);
and U694 (N_694,In_478,In_2177);
or U695 (N_695,In_31,In_907);
xnor U696 (N_696,In_1010,In_2557);
or U697 (N_697,In_2754,In_2098);
and U698 (N_698,In_114,In_153);
or U699 (N_699,In_2913,In_1627);
and U700 (N_700,In_1659,In_198);
or U701 (N_701,In_2433,In_1151);
and U702 (N_702,In_783,In_2780);
and U703 (N_703,In_1618,In_1013);
nand U704 (N_704,In_1281,In_2235);
xor U705 (N_705,In_1271,In_1469);
nand U706 (N_706,In_718,In_1429);
and U707 (N_707,In_2283,In_1951);
nand U708 (N_708,In_549,In_1068);
and U709 (N_709,In_1154,In_1770);
or U710 (N_710,In_2086,In_1396);
and U711 (N_711,In_2441,In_1876);
or U712 (N_712,In_2517,In_1860);
and U713 (N_713,In_1212,In_406);
or U714 (N_714,In_696,In_1668);
nor U715 (N_715,In_2428,In_2826);
nor U716 (N_716,In_668,In_2793);
or U717 (N_717,In_2529,In_2736);
and U718 (N_718,In_2345,In_2067);
xnor U719 (N_719,In_2140,In_2872);
or U720 (N_720,In_356,In_160);
nand U721 (N_721,In_1255,In_1593);
or U722 (N_722,In_2066,In_1833);
xor U723 (N_723,In_1355,In_2436);
xor U724 (N_724,In_327,In_15);
and U725 (N_725,In_2885,In_516);
nand U726 (N_726,In_1172,In_1482);
nand U727 (N_727,In_2904,In_394);
nand U728 (N_728,In_1440,In_2703);
xor U729 (N_729,In_2062,In_477);
nor U730 (N_730,In_851,In_1811);
xor U731 (N_731,In_555,In_2704);
xor U732 (N_732,In_1118,In_572);
or U733 (N_733,In_145,In_2702);
xnor U734 (N_734,In_1798,In_151);
or U735 (N_735,In_237,In_1989);
nor U736 (N_736,In_244,In_2240);
xnor U737 (N_737,In_1805,In_1269);
xor U738 (N_738,In_922,In_1522);
and U739 (N_739,In_2590,In_2187);
and U740 (N_740,In_473,In_2663);
nor U741 (N_741,In_2889,In_1107);
nor U742 (N_742,In_176,In_2303);
nor U743 (N_743,In_2992,In_38);
nor U744 (N_744,In_423,In_1468);
or U745 (N_745,In_2268,In_1831);
nand U746 (N_746,In_1822,In_383);
nor U747 (N_747,In_2777,In_18);
nand U748 (N_748,In_125,In_223);
nor U749 (N_749,In_1407,In_2410);
xnor U750 (N_750,In_1335,In_955);
and U751 (N_751,In_1607,In_2266);
nand U752 (N_752,In_2238,In_2467);
nor U753 (N_753,In_2942,In_1893);
and U754 (N_754,In_900,In_90);
xnor U755 (N_755,In_2046,In_946);
xor U756 (N_756,In_1922,In_593);
nor U757 (N_757,In_139,In_1645);
or U758 (N_758,In_265,In_971);
xor U759 (N_759,In_1033,In_2501);
or U760 (N_760,In_2188,In_197);
nor U761 (N_761,In_203,In_2319);
xnor U762 (N_762,In_2692,In_1603);
nand U763 (N_763,In_1606,In_437);
xnor U764 (N_764,In_713,In_2245);
or U765 (N_765,In_2148,In_1548);
nand U766 (N_766,In_809,In_800);
and U767 (N_767,In_92,In_2758);
nor U768 (N_768,In_1319,In_1367);
nor U769 (N_769,In_1245,In_2537);
nand U770 (N_770,In_2025,In_1073);
xnor U771 (N_771,In_2396,In_2116);
xnor U772 (N_772,In_2649,In_1276);
xnor U773 (N_773,In_2837,In_1572);
or U774 (N_774,In_1353,In_1923);
nor U775 (N_775,In_2315,In_1650);
and U776 (N_776,In_2508,In_441);
or U777 (N_777,In_0,In_1049);
nor U778 (N_778,In_2483,In_76);
xor U779 (N_779,In_730,In_562);
or U780 (N_780,In_1100,In_1818);
or U781 (N_781,In_1597,In_2833);
and U782 (N_782,In_726,In_2222);
or U783 (N_783,In_1604,In_1840);
or U784 (N_784,In_1821,In_2227);
or U785 (N_785,In_606,In_1442);
and U786 (N_786,In_2652,In_582);
xor U787 (N_787,In_2155,In_1242);
nand U788 (N_788,In_2073,In_996);
nand U789 (N_789,In_2406,In_273);
and U790 (N_790,In_1698,In_1113);
nor U791 (N_791,In_2395,In_885);
xnor U792 (N_792,In_1738,In_532);
nor U793 (N_793,In_64,In_2202);
and U794 (N_794,In_2748,In_2706);
nand U795 (N_795,In_1638,In_1771);
xnor U796 (N_796,In_623,In_2108);
nand U797 (N_797,In_1162,In_2561);
nand U798 (N_798,In_194,In_695);
and U799 (N_799,In_1901,In_1786);
or U800 (N_800,In_1114,In_2340);
nand U801 (N_801,In_514,In_1574);
and U802 (N_802,In_2743,In_2468);
and U803 (N_803,In_369,In_2197);
and U804 (N_804,In_1405,In_2493);
nor U805 (N_805,In_2966,In_2948);
or U806 (N_806,In_2035,In_1465);
xnor U807 (N_807,In_1562,In_2757);
nor U808 (N_808,In_1788,In_722);
nor U809 (N_809,In_2506,In_2931);
or U810 (N_810,In_723,In_2594);
and U811 (N_811,In_161,In_1079);
and U812 (N_812,In_764,In_2568);
nand U813 (N_813,In_1110,In_1532);
and U814 (N_814,In_2099,In_1782);
and U815 (N_815,In_309,In_417);
or U816 (N_816,In_2825,In_1202);
or U817 (N_817,In_576,In_2330);
and U818 (N_818,In_2803,In_1699);
xnor U819 (N_819,In_431,In_1203);
or U820 (N_820,In_104,In_1059);
nor U821 (N_821,In_2812,In_2693);
xnor U822 (N_822,In_2420,In_591);
or U823 (N_823,In_1145,In_196);
nand U824 (N_824,In_796,In_1500);
xnor U825 (N_825,In_543,In_2750);
and U826 (N_826,In_2321,In_2952);
xor U827 (N_827,In_121,In_2480);
nand U828 (N_828,In_2538,In_1963);
and U829 (N_829,In_1273,In_2520);
nor U830 (N_830,In_2093,In_2842);
or U831 (N_831,In_2440,In_232);
and U832 (N_832,In_1704,In_2058);
and U833 (N_833,In_2674,In_2682);
or U834 (N_834,In_667,In_601);
nand U835 (N_835,In_1773,In_115);
nor U836 (N_836,In_2011,In_1489);
nand U837 (N_837,In_1027,In_1102);
or U838 (N_838,In_2219,In_512);
or U839 (N_839,In_959,In_875);
nand U840 (N_840,In_2972,In_1507);
and U841 (N_841,In_932,In_1376);
nor U842 (N_842,In_163,In_942);
and U843 (N_843,In_973,In_2309);
nand U844 (N_844,In_1205,In_811);
or U845 (N_845,In_312,In_2914);
and U846 (N_846,In_1972,In_1265);
nand U847 (N_847,In_2800,In_964);
xor U848 (N_848,In_2512,In_2577);
and U849 (N_849,In_1764,In_1227);
and U850 (N_850,In_872,In_893);
and U851 (N_851,In_560,In_2716);
xnor U852 (N_852,In_2211,In_1399);
xor U853 (N_853,In_1608,In_1733);
nor U854 (N_854,In_2374,In_329);
nand U855 (N_855,In_1043,In_1009);
nor U856 (N_856,In_2822,In_2003);
nor U857 (N_857,In_168,In_2632);
xnor U858 (N_858,In_2795,In_2391);
or U859 (N_859,In_2766,In_1368);
nand U860 (N_860,In_2473,In_479);
xnor U861 (N_861,In_2794,In_1734);
or U862 (N_862,In_349,In_743);
nor U863 (N_863,In_1052,In_985);
nor U864 (N_864,In_450,In_1375);
and U865 (N_865,In_2364,In_1339);
nand U866 (N_866,In_828,In_98);
nor U867 (N_867,In_2681,In_2890);
and U868 (N_868,In_274,In_1928);
nor U869 (N_869,In_467,In_40);
nor U870 (N_870,In_483,In_2455);
nand U871 (N_871,In_2168,In_1766);
xor U872 (N_872,In_476,In_338);
or U873 (N_873,In_2574,In_253);
nand U874 (N_874,In_2727,In_2050);
or U875 (N_875,In_2623,In_1600);
nor U876 (N_876,In_2170,In_2597);
xor U877 (N_877,In_2739,In_224);
nand U878 (N_878,In_786,In_2128);
xor U879 (N_879,In_1815,In_1740);
nor U880 (N_880,In_1241,In_2331);
or U881 (N_881,In_972,In_2127);
xor U882 (N_882,In_583,In_39);
xnor U883 (N_883,In_184,In_732);
or U884 (N_884,In_246,In_2203);
nand U885 (N_885,In_788,In_390);
nor U886 (N_886,In_2734,In_2578);
nand U887 (N_887,In_2720,In_845);
nand U888 (N_888,In_170,In_1577);
xor U889 (N_889,In_322,In_2635);
nor U890 (N_890,In_1809,In_2974);
nand U891 (N_891,In_2218,In_671);
xnor U892 (N_892,In_1940,In_738);
and U893 (N_893,In_1422,In_2421);
or U894 (N_894,In_2892,In_2880);
xnor U895 (N_895,In_941,In_2271);
and U896 (N_896,In_1481,In_2839);
xnor U897 (N_897,In_374,In_266);
xor U898 (N_898,In_905,In_2171);
or U899 (N_899,In_1416,In_432);
and U900 (N_900,In_1763,In_2125);
nand U901 (N_901,In_1900,In_395);
or U902 (N_902,In_681,In_2301);
xnor U903 (N_903,In_2253,In_1630);
xnor U904 (N_904,In_929,In_2336);
nand U905 (N_905,In_618,In_2072);
or U906 (N_906,In_662,In_1910);
or U907 (N_907,In_637,In_2023);
nand U908 (N_908,In_1851,In_2768);
nor U909 (N_909,In_1937,In_935);
and U910 (N_910,In_2190,In_201);
nand U911 (N_911,In_2530,In_1221);
nor U912 (N_912,In_2699,In_745);
or U913 (N_913,In_780,In_939);
nand U914 (N_914,In_757,In_2583);
or U915 (N_915,In_416,In_2430);
nor U916 (N_916,In_32,In_566);
nor U917 (N_917,In_2767,In_2088);
nor U918 (N_918,In_2191,In_391);
nand U919 (N_919,In_2489,In_1894);
and U920 (N_920,In_2274,In_2602);
nand U921 (N_921,In_651,In_849);
nand U922 (N_922,In_2986,In_2281);
nand U923 (N_923,In_1754,In_2371);
and U924 (N_924,In_853,In_1677);
nand U925 (N_925,In_1456,In_401);
nand U926 (N_926,In_1654,In_1006);
nor U927 (N_927,In_1443,In_1384);
or U928 (N_928,In_2684,In_586);
and U929 (N_929,In_1044,In_358);
and U930 (N_930,In_2698,In_2536);
nor U931 (N_931,In_927,In_470);
xnor U932 (N_932,In_1004,In_1197);
xnor U933 (N_933,In_1089,In_213);
nor U934 (N_934,In_1174,In_556);
xnor U935 (N_935,In_2671,In_2185);
and U936 (N_936,In_2504,In_1159);
xnor U937 (N_937,In_1520,In_200);
and U938 (N_938,In_1329,In_2814);
and U939 (N_939,In_1487,In_1431);
xor U940 (N_940,In_1231,In_188);
xnor U941 (N_941,In_746,In_2761);
xnor U942 (N_942,In_2457,In_1438);
or U943 (N_943,In_2909,In_620);
and U944 (N_944,In_636,In_348);
and U945 (N_945,In_1723,In_775);
nor U946 (N_946,In_2816,In_154);
xor U947 (N_947,In_130,In_2030);
or U948 (N_948,In_813,In_1660);
and U949 (N_949,In_461,In_2466);
and U950 (N_950,In_755,In_526);
nor U951 (N_951,In_1461,In_1959);
or U952 (N_952,In_2346,In_801);
nand U953 (N_953,In_1224,In_2879);
and U954 (N_954,In_1266,In_1020);
or U955 (N_955,In_1312,In_749);
and U956 (N_956,In_2077,In_2977);
or U957 (N_957,In_30,In_1985);
nand U958 (N_958,In_2497,In_1793);
or U959 (N_959,In_428,In_1721);
nor U960 (N_960,In_997,In_2807);
nand U961 (N_961,In_2152,In_1690);
nand U962 (N_962,In_315,In_1735);
nand U963 (N_963,In_524,In_241);
nor U964 (N_964,In_1347,In_2648);
nand U965 (N_965,In_691,In_2233);
nand U966 (N_966,In_991,In_806);
or U967 (N_967,In_881,In_363);
xor U968 (N_968,In_2859,In_2669);
or U969 (N_969,In_1099,In_1703);
nor U970 (N_970,In_2976,In_181);
nand U971 (N_971,In_710,In_2985);
nand U972 (N_972,In_1784,In_962);
or U973 (N_973,In_1280,In_81);
xnor U974 (N_974,In_5,In_2164);
nand U975 (N_975,In_1260,In_2375);
and U976 (N_976,In_216,In_1986);
nor U977 (N_977,In_2452,In_892);
nand U978 (N_978,In_1436,In_1879);
or U979 (N_979,In_129,In_2646);
nor U980 (N_980,In_2194,In_1492);
nor U981 (N_981,In_930,In_1077);
or U982 (N_982,In_1546,In_1333);
nand U983 (N_983,In_2866,In_1672);
and U984 (N_984,In_2117,In_1168);
and U985 (N_985,In_854,In_773);
and U986 (N_986,In_934,In_1626);
nor U987 (N_987,In_236,In_1411);
nand U988 (N_988,In_2382,In_1106);
nor U989 (N_989,In_277,In_1023);
and U990 (N_990,In_976,In_1417);
or U991 (N_991,In_1541,In_1745);
or U992 (N_992,In_761,In_2627);
xor U993 (N_993,In_1768,In_1311);
nand U994 (N_994,In_2082,In_1817);
nor U995 (N_995,In_693,In_1887);
and U996 (N_996,In_1594,In_404);
nand U997 (N_997,In_2339,In_1883);
or U998 (N_998,In_916,In_857);
or U999 (N_999,In_45,In_1288);
xor U1000 (N_1000,In_1248,In_2564);
and U1001 (N_1001,In_975,In_1);
nand U1002 (N_1002,In_2843,In_1216);
nor U1003 (N_1003,In_1447,In_459);
xor U1004 (N_1004,In_2172,In_2475);
xnor U1005 (N_1005,In_43,In_1620);
or U1006 (N_1006,In_2449,In_2485);
xnor U1007 (N_1007,In_2978,In_1531);
or U1008 (N_1008,In_1783,In_818);
xor U1009 (N_1009,In_475,In_339);
xnor U1010 (N_1010,In_2811,In_2242);
or U1011 (N_1011,In_452,In_134);
xnor U1012 (N_1012,In_54,In_1930);
and U1013 (N_1013,In_1622,In_1648);
nor U1014 (N_1014,In_1753,In_239);
nor U1015 (N_1015,In_2922,In_1218);
nor U1016 (N_1016,In_2509,In_1063);
and U1017 (N_1017,In_131,In_2367);
nor U1018 (N_1018,In_1206,In_677);
and U1019 (N_1019,In_1716,In_2311);
or U1020 (N_1020,In_2111,In_2791);
nor U1021 (N_1021,In_1474,In_2621);
nand U1022 (N_1022,In_2244,In_772);
nand U1023 (N_1023,In_1945,In_2089);
nand U1024 (N_1024,In_307,In_2821);
nor U1025 (N_1025,In_1062,In_493);
and U1026 (N_1026,In_1101,In_1011);
or U1027 (N_1027,In_190,In_2162);
or U1028 (N_1028,In_1692,In_579);
nand U1029 (N_1029,In_2369,In_2999);
or U1030 (N_1030,In_1865,In_2353);
or U1031 (N_1031,In_770,In_436);
nor U1032 (N_1032,In_2397,In_2881);
or U1033 (N_1033,In_1108,In_2264);
nand U1034 (N_1034,In_759,In_412);
xor U1035 (N_1035,In_2786,In_1686);
nand U1036 (N_1036,In_1854,In_557);
and U1037 (N_1037,In_1451,In_2845);
and U1038 (N_1038,In_1875,In_609);
xnor U1039 (N_1039,In_547,In_604);
and U1040 (N_1040,In_539,In_1984);
and U1041 (N_1041,In_1726,In_683);
or U1042 (N_1042,In_2260,In_525);
nor U1043 (N_1043,In_1445,In_1244);
xnor U1044 (N_1044,In_537,In_1646);
nor U1045 (N_1045,In_963,In_2477);
nand U1046 (N_1046,In_610,In_2137);
and U1047 (N_1047,In_209,In_2318);
nand U1048 (N_1048,In_164,In_1962);
and U1049 (N_1049,In_1361,In_2645);
nand U1050 (N_1050,In_2662,In_2161);
nor U1051 (N_1051,In_1897,In_1561);
nand U1052 (N_1052,In_2112,In_2134);
nor U1053 (N_1053,In_293,In_2494);
xor U1054 (N_1054,In_1694,In_2532);
nand U1055 (N_1055,In_797,In_1187);
nor U1056 (N_1056,In_847,In_267);
nand U1057 (N_1057,In_1590,In_1806);
nand U1058 (N_1058,In_429,In_1971);
and U1059 (N_1059,In_2895,In_1170);
nor U1060 (N_1060,In_2915,In_2979);
or U1061 (N_1061,In_1943,In_463);
or U1062 (N_1062,In_464,In_1140);
xor U1063 (N_1063,In_808,In_659);
and U1064 (N_1064,In_435,In_846);
or U1065 (N_1065,In_634,In_1934);
nand U1066 (N_1066,In_1688,In_204);
nor U1067 (N_1067,In_2609,In_285);
or U1068 (N_1068,In_96,In_2368);
nand U1069 (N_1069,In_152,In_65);
and U1070 (N_1070,In_1464,In_324);
and U1071 (N_1071,In_2817,In_56);
and U1072 (N_1072,In_490,In_1001);
or U1073 (N_1073,In_2121,In_1732);
nor U1074 (N_1074,In_2474,In_1801);
or U1075 (N_1075,In_832,In_306);
or U1076 (N_1076,In_185,In_1838);
nand U1077 (N_1077,In_221,In_440);
xnor U1078 (N_1078,In_1530,In_255);
xnor U1079 (N_1079,In_1987,In_1836);
or U1080 (N_1080,In_2038,In_1235);
or U1081 (N_1081,In_2850,In_1575);
nor U1082 (N_1082,In_2214,In_1804);
nor U1083 (N_1083,In_74,In_1917);
nor U1084 (N_1084,In_1617,In_2034);
nor U1085 (N_1085,In_1557,In_1996);
xnor U1086 (N_1086,In_407,In_2522);
or U1087 (N_1087,In_2355,In_1825);
xor U1088 (N_1088,In_899,In_2995);
nand U1089 (N_1089,In_2402,In_2017);
and U1090 (N_1090,In_89,In_2372);
xor U1091 (N_1091,In_2097,In_863);
nand U1092 (N_1092,In_72,In_1545);
nand U1093 (N_1093,In_261,In_2387);
or U1094 (N_1094,In_567,In_2655);
nand U1095 (N_1095,In_2201,In_1742);
and U1096 (N_1096,In_589,In_688);
nor U1097 (N_1097,In_258,In_1758);
or U1098 (N_1098,In_805,In_629);
or U1099 (N_1099,In_642,In_2548);
or U1100 (N_1100,In_2588,In_2951);
xnor U1101 (N_1101,In_2707,In_995);
or U1102 (N_1102,In_1868,In_1274);
and U1103 (N_1103,In_741,In_2650);
nor U1104 (N_1104,In_1560,In_180);
nand U1105 (N_1105,In_902,In_93);
and U1106 (N_1106,In_1184,In_785);
and U1107 (N_1107,In_1037,In_1967);
xnor U1108 (N_1108,In_46,In_1567);
nand U1109 (N_1109,In_731,In_1096);
nor U1110 (N_1110,In_1444,In_2513);
and U1111 (N_1111,In_2639,In_799);
nand U1112 (N_1112,In_951,In_2730);
xor U1113 (N_1113,In_2745,In_664);
nor U1114 (N_1114,In_1936,In_1508);
xnor U1115 (N_1115,In_1718,In_2773);
nor U1116 (N_1116,In_2065,In_2528);
nor U1117 (N_1117,In_2005,In_110);
nor U1118 (N_1118,In_1320,In_2004);
nand U1119 (N_1119,In_1085,In_840);
nor U1120 (N_1120,In_2234,In_2126);
nor U1121 (N_1121,In_915,In_1035);
or U1122 (N_1122,In_2860,In_2740);
xnor U1123 (N_1123,In_1471,In_49);
xnor U1124 (N_1124,In_792,In_1488);
nor U1125 (N_1125,In_1497,In_2033);
and U1126 (N_1126,In_2711,In_269);
nor U1127 (N_1127,In_465,In_2022);
or U1128 (N_1128,In_1122,In_2776);
nand U1129 (N_1129,In_615,In_616);
xnor U1130 (N_1130,In_29,In_735);
or U1131 (N_1131,In_1387,In_1731);
nand U1132 (N_1132,In_82,In_101);
and U1133 (N_1133,In_1167,In_214);
or U1134 (N_1134,In_644,In_335);
and U1135 (N_1135,In_2677,In_1914);
nand U1136 (N_1136,In_612,In_2314);
or U1137 (N_1137,In_1512,In_669);
xnor U1138 (N_1138,In_2900,In_1385);
and U1139 (N_1139,In_2783,In_1119);
or U1140 (N_1140,In_1765,In_1134);
or U1141 (N_1141,In_1056,In_2586);
and U1142 (N_1142,In_122,In_2552);
or U1143 (N_1143,In_2617,In_2313);
nor U1144 (N_1144,In_653,In_1852);
nand U1145 (N_1145,In_1315,In_77);
nand U1146 (N_1146,In_1988,In_2924);
or U1147 (N_1147,In_316,In_175);
nor U1148 (N_1148,In_2055,In_2377);
or U1149 (N_1149,In_2334,In_1334);
nand U1150 (N_1150,In_2426,In_1819);
nor U1151 (N_1151,In_814,In_2753);
nand U1152 (N_1152,In_1671,In_1364);
xor U1153 (N_1153,In_2358,In_1222);
and U1154 (N_1154,In_763,In_686);
or U1155 (N_1155,In_1824,In_856);
or U1156 (N_1156,In_1019,In_1008);
xnor U1157 (N_1157,In_336,In_466);
or U1158 (N_1158,In_2206,In_36);
or U1159 (N_1159,In_2715,In_2746);
and U1160 (N_1160,In_1249,In_1658);
nand U1161 (N_1161,In_1882,In_1503);
nor U1162 (N_1162,In_2348,In_558);
nor U1163 (N_1163,In_123,In_2902);
nand U1164 (N_1164,In_1322,In_1678);
and U1165 (N_1165,In_2031,In_61);
and U1166 (N_1166,In_460,In_2343);
xnor U1167 (N_1167,In_2335,In_2279);
nor U1168 (N_1168,In_859,In_2770);
nand U1169 (N_1169,In_1374,In_552);
and U1170 (N_1170,In_9,In_298);
nand U1171 (N_1171,In_171,In_1643);
nor U1172 (N_1172,In_1640,In_2189);
xor U1173 (N_1173,In_498,In_359);
nor U1174 (N_1174,In_1239,In_405);
or U1175 (N_1175,In_1165,In_1360);
nor U1176 (N_1176,In_1002,In_42);
xor U1177 (N_1177,In_913,In_444);
nor U1178 (N_1178,In_1067,In_2543);
nand U1179 (N_1179,In_2370,In_2638);
nand U1180 (N_1180,In_367,In_2496);
and U1181 (N_1181,In_1305,In_890);
and U1182 (N_1182,In_2262,In_970);
or U1183 (N_1183,In_2956,In_2287);
and U1184 (N_1184,In_1855,In_527);
and U1185 (N_1185,In_758,In_944);
or U1186 (N_1186,In_438,In_1493);
or U1187 (N_1187,In_328,In_2608);
or U1188 (N_1188,In_379,In_1181);
and U1189 (N_1189,In_2941,In_2207);
nor U1190 (N_1190,In_2911,In_1990);
and U1191 (N_1191,In_2679,In_2762);
nor U1192 (N_1192,In_966,In_57);
and U1193 (N_1193,In_756,In_2818);
nor U1194 (N_1194,In_2460,In_1719);
nand U1195 (N_1195,In_961,In_1277);
nand U1196 (N_1196,In_908,In_682);
xor U1197 (N_1197,In_1663,In_2186);
and U1198 (N_1198,In_2969,In_1864);
or U1199 (N_1199,In_1554,In_1976);
nor U1200 (N_1200,N_1170,N_679);
nand U1201 (N_1201,In_928,N_751);
and U1202 (N_1202,N_1050,N_118);
or U1203 (N_1203,N_537,In_1460);
or U1204 (N_1204,N_710,N_802);
nor U1205 (N_1205,In_2957,N_867);
or U1206 (N_1206,In_1074,N_809);
and U1207 (N_1207,N_22,In_2523);
nor U1208 (N_1208,N_574,In_2769);
nor U1209 (N_1209,N_995,In_2865);
and U1210 (N_1210,In_1752,N_371);
or U1211 (N_1211,In_1380,In_50);
nor U1212 (N_1212,N_116,In_1042);
and U1213 (N_1213,N_74,N_81);
nor U1214 (N_1214,N_536,N_0);
xor U1215 (N_1215,In_1423,In_2556);
nor U1216 (N_1216,N_17,N_1047);
or U1217 (N_1217,N_1080,N_305);
nand U1218 (N_1218,N_1163,N_839);
nand U1219 (N_1219,In_520,N_317);
nand U1220 (N_1220,N_390,In_737);
xor U1221 (N_1221,In_2103,N_420);
and U1222 (N_1222,N_324,N_38);
and U1223 (N_1223,N_300,N_443);
nor U1224 (N_1224,N_267,N_766);
xor U1225 (N_1225,In_584,N_911);
xor U1226 (N_1226,In_2438,N_963);
nand U1227 (N_1227,In_1061,In_2950);
and U1228 (N_1228,N_812,N_554);
xor U1229 (N_1229,In_1278,N_470);
xnor U1230 (N_1230,In_399,N_858);
nand U1231 (N_1231,N_1040,N_992);
and U1232 (N_1232,N_769,N_152);
and U1233 (N_1233,N_1157,In_2721);
and U1234 (N_1234,N_861,N_343);
and U1235 (N_1235,N_738,N_688);
or U1236 (N_1236,In_2305,N_345);
or U1237 (N_1237,In_1000,In_974);
or U1238 (N_1238,In_1229,N_850);
nor U1239 (N_1239,N_314,N_180);
nor U1240 (N_1240,N_1165,In_917);
nor U1241 (N_1241,In_1392,In_2224);
nor U1242 (N_1242,In_2230,In_2657);
and U1243 (N_1243,N_277,In_568);
or U1244 (N_1244,N_755,N_583);
and U1245 (N_1245,N_296,N_23);
or U1246 (N_1246,N_313,N_76);
or U1247 (N_1247,N_650,N_1090);
nand U1248 (N_1248,N_818,N_1147);
xor U1249 (N_1249,N_582,N_524);
nand U1250 (N_1250,N_288,In_1475);
xnor U1251 (N_1251,In_720,N_978);
or U1252 (N_1252,In_841,N_547);
or U1253 (N_1253,In_219,In_2422);
nand U1254 (N_1254,In_949,In_2910);
nand U1255 (N_1255,N_286,In_1621);
nand U1256 (N_1256,N_223,In_2289);
or U1257 (N_1257,N_873,N_311);
nand U1258 (N_1258,N_432,N_1005);
nor U1259 (N_1259,N_778,In_2248);
nor U1260 (N_1260,N_681,In_2862);
xor U1261 (N_1261,N_323,N_170);
nor U1262 (N_1262,N_438,In_2797);
or U1263 (N_1263,In_977,N_25);
nor U1264 (N_1264,N_393,In_2545);
xor U1265 (N_1265,N_217,In_1064);
or U1266 (N_1266,N_959,In_751);
or U1267 (N_1267,N_897,N_764);
and U1268 (N_1268,N_527,N_977);
nor U1269 (N_1269,In_1047,N_927);
nor U1270 (N_1270,In_2846,In_1552);
nor U1271 (N_1271,In_345,N_303);
xnor U1272 (N_1272,In_1289,In_1553);
nand U1273 (N_1273,N_1117,N_1175);
nor U1274 (N_1274,N_558,N_991);
nand U1275 (N_1275,N_147,N_204);
or U1276 (N_1276,N_875,N_1176);
xor U1277 (N_1277,N_670,In_1354);
xor U1278 (N_1278,N_1191,N_306);
xnor U1279 (N_1279,N_689,In_1163);
and U1280 (N_1280,N_246,N_120);
nor U1281 (N_1281,N_731,N_381);
and U1282 (N_1282,N_785,N_95);
nand U1283 (N_1283,N_335,N_326);
and U1284 (N_1284,N_194,In_1171);
and U1285 (N_1285,N_1186,In_2709);
nor U1286 (N_1286,N_829,In_879);
or U1287 (N_1287,N_621,N_932);
nor U1288 (N_1288,N_505,In_249);
and U1289 (N_1289,N_484,In_382);
nand U1290 (N_1290,In_787,N_700);
nor U1291 (N_1291,N_1143,N_1011);
xor U1292 (N_1292,N_803,In_1750);
nor U1293 (N_1293,N_433,In_2200);
xnor U1294 (N_1294,N_685,In_599);
or U1295 (N_1295,N_151,In_666);
xor U1296 (N_1296,In_2854,In_2643);
and U1297 (N_1297,N_713,In_1929);
nor U1298 (N_1298,In_1975,N_287);
and U1299 (N_1299,N_653,N_881);
or U1300 (N_1300,N_1142,N_570);
and U1301 (N_1301,N_395,N_447);
xor U1302 (N_1302,N_934,In_1605);
nor U1303 (N_1303,In_1504,In_1486);
and U1304 (N_1304,N_1067,N_889);
nand U1305 (N_1305,N_942,N_592);
nor U1306 (N_1306,N_66,N_12);
or U1307 (N_1307,In_497,In_2208);
xor U1308 (N_1308,In_2166,In_1029);
xor U1309 (N_1309,In_446,N_55);
or U1310 (N_1310,N_131,N_290);
xnor U1311 (N_1311,N_789,N_801);
nand U1312 (N_1312,N_657,In_2967);
and U1313 (N_1313,N_195,In_469);
or U1314 (N_1314,In_1586,N_871);
and U1315 (N_1315,N_140,N_816);
nand U1316 (N_1316,In_1111,N_855);
and U1317 (N_1317,In_2983,In_1791);
nand U1318 (N_1318,In_1904,N_815);
or U1319 (N_1319,In_2997,N_580);
nor U1320 (N_1320,N_1035,In_1582);
or U1321 (N_1321,In_233,N_316);
nor U1322 (N_1322,N_788,N_509);
nor U1323 (N_1323,N_322,In_1674);
nand U1324 (N_1324,In_573,N_754);
and U1325 (N_1325,N_783,N_627);
nor U1326 (N_1326,N_595,N_649);
nor U1327 (N_1327,N_844,In_2383);
and U1328 (N_1328,N_464,In_2151);
xor U1329 (N_1329,N_89,In_2542);
nor U1330 (N_1330,N_284,N_1032);
nor U1331 (N_1331,N_355,In_2636);
nand U1332 (N_1332,N_28,N_215);
xnor U1333 (N_1333,N_918,N_282);
or U1334 (N_1334,N_1189,N_704);
and U1335 (N_1335,N_1138,N_511);
or U1336 (N_1336,N_373,N_1199);
or U1337 (N_1337,In_2394,N_672);
or U1338 (N_1338,In_1684,N_758);
or U1339 (N_1339,N_996,N_687);
nor U1340 (N_1340,N_849,N_763);
or U1341 (N_1341,N_13,In_2664);
or U1342 (N_1342,N_436,N_930);
xnor U1343 (N_1343,In_2389,N_218);
and U1344 (N_1344,N_986,In_1969);
or U1345 (N_1345,N_709,N_281);
or U1346 (N_1346,N_94,N_1064);
nor U1347 (N_1347,N_1108,N_1187);
or U1348 (N_1348,In_1104,In_1164);
xnor U1349 (N_1349,N_1000,N_361);
xnor U1350 (N_1350,N_1159,N_923);
xnor U1351 (N_1351,N_34,N_877);
nand U1352 (N_1352,In_1083,N_1169);
and U1353 (N_1353,N_571,N_837);
and U1354 (N_1354,N_890,N_581);
nor U1355 (N_1355,In_701,N_42);
xor U1356 (N_1356,N_833,In_2661);
and U1357 (N_1357,N_888,N_1131);
and U1358 (N_1358,N_944,In_2246);
and U1359 (N_1359,In_705,N_1043);
xnor U1360 (N_1360,N_1155,N_775);
xor U1361 (N_1361,N_185,N_784);
and U1362 (N_1362,N_500,In_2076);
or U1363 (N_1363,N_1190,N_382);
nand U1364 (N_1364,N_933,In_2802);
nor U1365 (N_1365,In_2347,In_2696);
xor U1366 (N_1366,In_1325,N_544);
nand U1367 (N_1367,In_1974,N_123);
nand U1368 (N_1368,N_1072,In_22);
and U1369 (N_1369,N_734,In_1146);
and U1370 (N_1370,In_2122,In_186);
nand U1371 (N_1371,In_1370,N_901);
and U1372 (N_1372,In_2015,N_1110);
or U1373 (N_1373,N_533,N_675);
or U1374 (N_1374,N_411,N_1078);
nor U1375 (N_1375,N_646,N_82);
nor U1376 (N_1376,N_1181,N_517);
or U1377 (N_1377,N_1174,N_232);
or U1378 (N_1378,N_872,In_2447);
nand U1379 (N_1379,N_456,In_1345);
nand U1380 (N_1380,In_1757,N_1087);
xor U1381 (N_1381,N_946,N_78);
nor U1382 (N_1382,N_656,N_273);
nor U1383 (N_1383,N_454,N_61);
or U1384 (N_1384,In_1693,N_668);
or U1385 (N_1385,N_422,N_1178);
or U1386 (N_1386,N_1122,In_211);
and U1387 (N_1387,In_2728,In_2647);
nand U1388 (N_1388,N_762,In_2101);
nand U1389 (N_1389,N_884,In_1808);
or U1390 (N_1390,N_1034,N_1133);
or U1391 (N_1391,In_704,N_136);
or U1392 (N_1392,N_201,N_701);
or U1393 (N_1393,N_1009,N_935);
nor U1394 (N_1394,N_642,N_980);
nor U1395 (N_1395,N_851,N_974);
and U1396 (N_1396,N_431,N_1082);
nor U1397 (N_1397,N_260,N_9);
xor U1398 (N_1398,N_637,N_444);
and U1399 (N_1399,In_2417,N_599);
or U1400 (N_1400,N_631,N_961);
or U1401 (N_1401,In_1517,N_33);
xor U1402 (N_1402,N_1070,In_1058);
or U1403 (N_1403,N_718,In_2095);
or U1404 (N_1404,N_47,In_1188);
nor U1405 (N_1405,N_612,N_245);
and U1406 (N_1406,N_402,N_1008);
and U1407 (N_1407,In_24,N_674);
nor U1408 (N_1408,N_920,In_1328);
nand U1409 (N_1409,N_58,N_418);
nor U1410 (N_1410,In_626,N_838);
nor U1411 (N_1411,N_467,N_548);
nand U1412 (N_1412,N_272,N_1049);
xnor U1413 (N_1413,N_430,N_1135);
nand U1414 (N_1414,N_825,N_985);
or U1415 (N_1415,N_87,In_869);
or U1416 (N_1416,N_1168,N_318);
xor U1417 (N_1417,N_1028,N_663);
nor U1418 (N_1418,In_279,In_2603);
nand U1419 (N_1419,In_2226,N_57);
nor U1420 (N_1420,N_477,In_55);
nor U1421 (N_1421,N_109,In_2990);
or U1422 (N_1422,In_2007,N_952);
xnor U1423 (N_1423,N_513,N_1145);
or U1424 (N_1424,N_31,In_259);
nand U1425 (N_1425,N_1152,N_146);
and U1426 (N_1426,N_144,N_578);
nor U1427 (N_1427,In_91,In_2499);
nor U1428 (N_1428,In_2932,N_231);
nor U1429 (N_1429,In_1837,N_613);
nor U1430 (N_1430,N_1154,N_37);
xor U1431 (N_1431,N_230,N_63);
xnor U1432 (N_1432,In_1283,N_234);
nor U1433 (N_1433,In_2725,N_1111);
or U1434 (N_1434,In_2908,N_153);
or U1435 (N_1435,In_1525,In_1014);
and U1436 (N_1436,N_45,N_161);
and U1437 (N_1437,N_224,N_1184);
or U1438 (N_1438,N_501,N_575);
xor U1439 (N_1439,N_384,N_665);
and U1440 (N_1440,N_865,In_2316);
xnor U1441 (N_1441,N_647,N_293);
nand U1442 (N_1442,N_966,In_2320);
xor U1443 (N_1443,In_518,N_666);
or U1444 (N_1444,N_807,N_53);
xnor U1445 (N_1445,N_417,N_327);
and U1446 (N_1446,N_869,In_1196);
and U1447 (N_1447,In_911,N_1093);
nor U1448 (N_1448,In_1992,N_310);
nor U1449 (N_1449,N_552,N_494);
nor U1450 (N_1450,N_1031,N_834);
or U1451 (N_1451,N_496,N_354);
and U1452 (N_1452,In_1304,N_1015);
nand U1453 (N_1453,In_719,In_2518);
xor U1454 (N_1454,In_1874,N_1068);
or U1455 (N_1455,N_1021,N_465);
or U1456 (N_1456,N_100,N_486);
nand U1457 (N_1457,N_392,N_192);
nand U1458 (N_1458,N_266,In_1105);
nand U1459 (N_1459,In_2539,N_958);
nand U1460 (N_1460,In_2917,N_307);
xnor U1461 (N_1461,N_439,In_1341);
nor U1462 (N_1462,N_60,N_683);
nor U1463 (N_1463,N_360,N_619);
nor U1464 (N_1464,N_940,N_828);
and U1465 (N_1465,N_423,N_673);
nor U1466 (N_1466,N_761,In_740);
nor U1467 (N_1467,N_474,In_1795);
nand U1468 (N_1468,In_947,In_835);
nand U1469 (N_1469,N_261,N_1010);
nor U1470 (N_1470,N_862,In_2918);
nand U1471 (N_1471,N_1029,In_1142);
xnor U1472 (N_1472,In_275,N_387);
or U1473 (N_1473,In_2629,N_122);
and U1474 (N_1474,N_169,N_705);
and U1475 (N_1475,N_1048,N_1179);
nand U1476 (N_1476,N_154,N_1006);
and U1477 (N_1477,N_1148,N_1037);
and U1478 (N_1478,N_32,N_950);
and U1479 (N_1479,In_1587,N_883);
xnor U1480 (N_1480,N_1183,N_1177);
xor U1481 (N_1481,N_577,In_673);
nand U1482 (N_1482,N_1128,In_2531);
and U1483 (N_1483,In_2789,In_1302);
nor U1484 (N_1484,N_655,In_1117);
nand U1485 (N_1485,N_479,N_448);
or U1486 (N_1486,N_229,N_150);
or U1487 (N_1487,N_110,In_287);
or U1488 (N_1488,In_1391,N_951);
or U1489 (N_1489,N_208,N_75);
nor U1490 (N_1490,In_1676,In_454);
or U1491 (N_1491,In_157,N_1158);
nand U1492 (N_1492,N_863,N_589);
nor U1493 (N_1493,N_400,N_104);
xnor U1494 (N_1494,In_2199,N_896);
and U1495 (N_1495,N_1098,N_606);
xnor U1496 (N_1496,In_1785,N_732);
and U1497 (N_1497,N_878,In_670);
xnor U1498 (N_1498,N_347,N_566);
or U1499 (N_1499,N_244,In_689);
and U1500 (N_1500,N_1081,In_509);
and U1501 (N_1501,N_915,N_835);
nor U1502 (N_1502,In_850,N_199);
nor U1503 (N_1503,N_598,In_2044);
nand U1504 (N_1504,N_600,In_447);
nand U1505 (N_1505,N_771,N_1060);
and U1506 (N_1506,In_1602,N_279);
and U1507 (N_1507,N_913,N_69);
or U1508 (N_1508,In_231,N_782);
nor U1509 (N_1509,N_591,N_259);
nand U1510 (N_1510,N_939,N_960);
nor U1511 (N_1511,In_1776,N_325);
xor U1512 (N_1512,In_894,N_954);
and U1513 (N_1513,In_2465,N_895);
or U1514 (N_1514,N_587,In_1707);
or U1515 (N_1515,N_730,N_328);
nor U1516 (N_1516,In_887,In_739);
nor U1517 (N_1517,N_483,N_810);
nand U1518 (N_1518,N_765,N_520);
nand U1519 (N_1519,In_132,N_105);
and U1520 (N_1520,N_178,N_112);
or U1521 (N_1521,N_1124,In_2926);
or U1522 (N_1522,N_96,In_1906);
nor U1523 (N_1523,In_300,N_1182);
nor U1524 (N_1524,N_874,N_1153);
nand U1525 (N_1525,In_146,In_2174);
and U1526 (N_1526,N_337,N_319);
nor U1527 (N_1527,N_396,N_356);
nor U1528 (N_1528,In_250,N_125);
or U1529 (N_1529,In_396,N_793);
nor U1530 (N_1530,N_880,N_1160);
xnor U1531 (N_1531,N_1099,N_622);
nand U1532 (N_1532,N_706,N_248);
or U1533 (N_1533,In_2288,N_969);
xnor U1534 (N_1534,In_515,In_1336);
nand U1535 (N_1535,In_1762,In_397);
nand U1536 (N_1536,N_220,N_879);
nor U1537 (N_1537,N_492,N_126);
and U1538 (N_1538,In_1439,N_737);
and U1539 (N_1539,N_508,In_2041);
or U1540 (N_1540,N_545,N_295);
xor U1541 (N_1541,N_528,N_906);
or U1542 (N_1542,N_725,N_590);
xor U1543 (N_1543,In_2899,N_1046);
or U1544 (N_1544,N_117,N_389);
nor U1545 (N_1545,In_2100,N_553);
nand U1546 (N_1546,N_945,In_1069);
or U1547 (N_1547,N_183,N_712);
xnor U1548 (N_1548,In_138,N_143);
nor U1549 (N_1549,N_635,In_1624);
nand U1550 (N_1550,N_956,In_1797);
nor U1551 (N_1551,N_611,N_241);
or U1552 (N_1552,N_957,In_402);
xor U1553 (N_1553,N_19,In_2160);
or U1554 (N_1554,In_2685,In_2482);
xnor U1555 (N_1555,In_489,N_502);
or U1556 (N_1556,N_1024,N_106);
nor U1557 (N_1557,In_635,In_1591);
or U1558 (N_1558,In_1372,N_555);
xor U1559 (N_1559,N_214,N_588);
and U1560 (N_1560,In_1454,In_625);
nor U1561 (N_1561,In_1330,In_1040);
xor U1562 (N_1562,N_1065,In_1950);
or U1563 (N_1563,N_1071,N_79);
nor U1564 (N_1564,In_692,N_461);
xnor U1565 (N_1565,In_1282,In_1261);
xor U1566 (N_1566,N_249,In_434);
and U1567 (N_1567,In_2628,N_20);
and U1568 (N_1568,N_336,N_206);
nor U1569 (N_1569,N_735,In_1625);
nor U1570 (N_1570,In_2898,N_690);
nand U1571 (N_1571,N_349,In_1125);
nor U1572 (N_1572,N_405,N_363);
nor U1573 (N_1573,In_1568,N_830);
xor U1574 (N_1574,N_333,In_360);
or U1575 (N_1575,N_716,In_2691);
nand U1576 (N_1576,N_891,N_164);
and U1577 (N_1577,In_2796,N_276);
nor U1578 (N_1578,N_852,N_275);
nand U1579 (N_1579,N_383,N_1198);
and U1580 (N_1580,N_813,In_1467);
nor U1581 (N_1581,N_222,In_954);
and U1582 (N_1582,N_1053,N_845);
nor U1583 (N_1583,In_2653,In_301);
xnor U1584 (N_1584,N_15,N_997);
xor U1585 (N_1585,N_943,N_184);
or U1586 (N_1586,N_854,N_601);
and U1587 (N_1587,In_354,N_593);
or U1588 (N_1588,N_727,In_2048);
nand U1589 (N_1589,N_175,N_301);
nand U1590 (N_1590,In_621,In_1905);
nand U1591 (N_1591,N_1086,N_573);
and U1592 (N_1592,N_667,N_1141);
or U1593 (N_1593,In_1088,N_1134);
nand U1594 (N_1594,In_4,N_289);
or U1595 (N_1595,N_129,In_2490);
xor U1596 (N_1596,N_119,N_999);
xnor U1597 (N_1597,N_1149,N_1089);
xnor U1598 (N_1598,N_767,N_614);
and U1599 (N_1599,N_269,In_439);
xnor U1600 (N_1600,N_584,N_556);
xnor U1601 (N_1601,In_870,In_2678);
nand U1602 (N_1602,N_252,N_348);
or U1603 (N_1603,N_937,N_346);
xnor U1604 (N_1604,In_1296,N_714);
nor U1605 (N_1605,N_226,In_1888);
nor U1606 (N_1606,N_842,N_831);
or U1607 (N_1607,In_1365,N_907);
and U1608 (N_1608,N_86,N_207);
nor U1609 (N_1609,N_676,N_46);
xor U1610 (N_1610,In_1637,In_1942);
or U1611 (N_1611,In_2141,In_2903);
nor U1612 (N_1612,N_72,In_1070);
nor U1613 (N_1613,N_334,N_680);
or U1614 (N_1614,N_1042,N_497);
or U1615 (N_1615,N_107,In_762);
or U1616 (N_1616,N_83,N_750);
and U1617 (N_1617,In_193,N_662);
and U1618 (N_1618,N_882,N_1118);
nor U1619 (N_1619,N_299,N_724);
xnor U1620 (N_1620,N_359,In_1918);
nor U1621 (N_1621,N_250,N_525);
and U1622 (N_1622,N_610,In_17);
xor U1623 (N_1623,N_742,N_264);
and U1624 (N_1624,N_753,N_40);
nand U1625 (N_1625,In_1667,N_693);
nor U1626 (N_1626,N_466,In_2157);
xor U1627 (N_1627,In_590,In_2390);
or U1628 (N_1628,N_777,In_624);
xor U1629 (N_1629,In_1547,In_1430);
nor U1630 (N_1630,N_186,N_684);
nand U1631 (N_1631,N_428,N_427);
or U1632 (N_1632,In_596,In_2891);
nand U1633 (N_1633,N_510,In_2994);
or U1634 (N_1634,In_16,N_399);
or U1635 (N_1635,In_2929,In_2360);
or U1636 (N_1636,N_1018,N_671);
nor U1637 (N_1637,N_805,N_10);
or U1638 (N_1638,In_1583,N_190);
nor U1639 (N_1639,N_1023,In_646);
xor U1640 (N_1640,N_274,N_521);
nand U1641 (N_1641,N_962,N_1094);
or U1642 (N_1642,N_166,In_2510);
xnor U1643 (N_1643,N_696,N_233);
nand U1644 (N_1644,N_885,N_437);
xor U1645 (N_1645,N_221,N_955);
and U1646 (N_1646,N_795,N_235);
nand U1647 (N_1647,N_168,N_44);
or U1648 (N_1648,N_538,N_1014);
nor U1649 (N_1649,N_350,N_173);
nand U1650 (N_1650,N_859,N_564);
xnor U1651 (N_1651,N_351,In_1820);
nand U1652 (N_1652,In_712,In_1516);
nand U1653 (N_1653,N_529,In_1514);
and U1654 (N_1654,N_139,N_64);
nand U1655 (N_1655,N_506,N_242);
and U1656 (N_1656,In_1528,N_973);
nand U1657 (N_1657,In_654,N_216);
xnor U1658 (N_1658,In_1612,N_133);
nand U1659 (N_1659,N_1054,N_375);
and U1660 (N_1660,N_924,N_237);
nand U1661 (N_1661,N_617,N_1129);
and U1662 (N_1662,N_263,N_62);
and U1663 (N_1663,N_177,In_2549);
nor U1664 (N_1664,N_625,In_319);
xnor U1665 (N_1665,In_1835,In_2138);
or U1666 (N_1666,N_604,In_2182);
xnor U1667 (N_1667,N_472,N_603);
and U1668 (N_1668,In_1903,N_787);
nand U1669 (N_1669,N_569,In_415);
and U1670 (N_1670,N_342,N_378);
and U1671 (N_1671,In_2105,N_182);
nand U1672 (N_1672,In_1685,In_982);
and U1673 (N_1673,N_41,N_929);
xor U1674 (N_1674,In_2641,N_534);
nand U1675 (N_1675,N_377,N_847);
nor U1676 (N_1676,N_1033,In_1571);
nand U1677 (N_1677,N_644,N_315);
nand U1678 (N_1678,N_137,In_2625);
and U1679 (N_1679,N_132,N_141);
nor U1680 (N_1680,N_2,N_608);
xnor U1681 (N_1681,N_557,N_928);
or U1682 (N_1682,N_899,N_715);
xnor U1683 (N_1683,N_1001,In_1072);
nand U1684 (N_1684,In_2144,N_243);
nor U1685 (N_1685,N_451,N_1016);
xor U1686 (N_1686,N_794,N_507);
nand U1687 (N_1687,In_1207,N_56);
and U1688 (N_1688,N_128,In_2456);
nor U1689 (N_1689,N_826,N_925);
or U1690 (N_1690,N_172,N_605);
xor U1691 (N_1691,N_1162,In_2947);
nor U1692 (N_1692,N_408,N_35);
xor U1693 (N_1693,In_2673,N_101);
nand U1694 (N_1694,N_814,N_870);
nand U1695 (N_1695,N_54,N_8);
or U1696 (N_1696,N_824,N_904);
xor U1697 (N_1697,In_2195,In_148);
xor U1698 (N_1698,N_388,N_134);
and U1699 (N_1699,In_575,N_340);
nor U1700 (N_1700,N_1103,N_191);
nand U1701 (N_1701,N_1059,N_984);
nor U1702 (N_1702,N_941,N_341);
nand U1703 (N_1703,In_564,N_618);
nor U1704 (N_1704,In_2855,N_6);
and U1705 (N_1705,N_493,In_820);
nor U1706 (N_1706,N_745,N_546);
or U1707 (N_1707,N_623,N_434);
and U1708 (N_1708,N_531,N_1195);
and U1709 (N_1709,In_2398,N_298);
and U1710 (N_1710,In_1717,In_708);
and U1711 (N_1711,N_320,In_793);
xor U1712 (N_1712,N_752,In_1755);
xor U1713 (N_1713,In_1349,N_516);
nand U1714 (N_1714,In_919,In_984);
nand U1715 (N_1715,In_2971,In_1275);
nand U1716 (N_1716,N_1137,N_791);
and U1717 (N_1717,In_883,In_672);
nor U1718 (N_1718,N_1116,N_512);
or U1719 (N_1719,N_271,N_450);
xor U1720 (N_1720,N_926,N_1004);
and U1721 (N_1721,N_70,N_265);
nand U1722 (N_1722,In_1138,N_1020);
and U1723 (N_1723,N_1109,N_616);
xor U1724 (N_1724,N_1125,N_1156);
nor U1725 (N_1725,N_1105,In_2056);
xor U1726 (N_1726,In_1682,In_1098);
or U1727 (N_1727,N_998,N_692);
or U1728 (N_1728,N_975,N_1120);
and U1729 (N_1729,In_381,N_567);
nor U1730 (N_1730,N_1030,N_864);
nand U1731 (N_1731,N_856,In_1510);
xor U1732 (N_1732,N_722,N_482);
xor U1733 (N_1733,N_452,N_948);
nor U1734 (N_1734,In_2589,N_968);
nor U1735 (N_1735,N_979,N_398);
or U1736 (N_1736,N_202,In_2403);
or U1737 (N_1737,In_1433,In_1596);
nand U1738 (N_1738,N_179,N_189);
or U1739 (N_1739,In_2337,N_990);
nor U1740 (N_1740,In_2399,N_659);
nor U1741 (N_1741,N_425,N_744);
nor U1742 (N_1742,N_550,N_846);
nor U1743 (N_1743,N_702,In_1055);
nand U1744 (N_1744,N_1104,In_337);
xnor U1745 (N_1745,In_2928,N_549);
nand U1746 (N_1746,N_628,N_1188);
xnor U1747 (N_1747,N_1,N_386);
xor U1748 (N_1748,In_2591,In_501);
xnor U1749 (N_1749,In_839,N_1185);
nand U1750 (N_1750,In_2503,N_48);
xnor U1751 (N_1751,N_1013,N_11);
nand U1752 (N_1752,In_641,In_986);
nor U1753 (N_1753,In_608,N_772);
or U1754 (N_1754,N_379,N_660);
and U1755 (N_1755,N_357,N_385);
xnor U1756 (N_1756,In_2840,N_736);
and U1757 (N_1757,In_752,In_2887);
nor U1758 (N_1758,N_495,N_3);
xor U1759 (N_1759,N_409,N_394);
nor U1760 (N_1760,In_1393,N_1039);
nand U1761 (N_1761,In_2644,N_304);
xor U1762 (N_1762,N_1083,In_10);
xnor U1763 (N_1763,N_596,N_1114);
or U1764 (N_1764,N_406,In_418);
xor U1765 (N_1765,N_756,N_124);
xnor U1766 (N_1766,N_1100,In_1472);
nand U1767 (N_1767,N_1161,N_779);
and U1768 (N_1768,N_1172,N_993);
or U1769 (N_1769,N_648,N_808);
xor U1770 (N_1770,N_1063,In_1832);
nor U1771 (N_1771,N_238,N_1119);
xor U1772 (N_1772,N_415,In_2365);
or U1773 (N_1773,N_982,N_97);
nor U1774 (N_1774,N_1113,N_163);
and U1775 (N_1775,N_770,N_1058);
or U1776 (N_1776,N_121,N_167);
nor U1777 (N_1777,N_914,N_424);
or U1778 (N_1778,In_649,N_1077);
and U1779 (N_1779,N_1003,N_843);
and U1780 (N_1780,In_1157,N_330);
nor U1781 (N_1781,N_130,In_1243);
and U1782 (N_1782,N_585,N_98);
xnor U1783 (N_1783,N_99,In_1870);
and U1784 (N_1784,N_607,In_1401);
nand U1785 (N_1785,In_2392,N_445);
and U1786 (N_1786,N_840,N_142);
xor U1787 (N_1787,N_212,N_1096);
or U1788 (N_1788,N_916,N_632);
and U1789 (N_1789,In_174,In_2180);
xnor U1790 (N_1790,N_799,N_630);
xnor U1791 (N_1791,N_1144,In_2308);
and U1792 (N_1792,In_1490,N_1126);
and U1793 (N_1793,In_1729,In_2476);
nand U1794 (N_1794,N_1192,N_638);
and U1795 (N_1795,In_1054,N_412);
or U1796 (N_1796,In_921,In_521);
nand U1797 (N_1797,N_760,N_698);
xnor U1798 (N_1798,N_894,N_703);
and U1799 (N_1799,N_720,In_2573);
nor U1800 (N_1800,In_398,In_368);
xor U1801 (N_1801,N_746,In_2805);
nand U1802 (N_1802,N_380,N_919);
or U1803 (N_1803,N_900,N_353);
nor U1804 (N_1804,N_292,N_1196);
nand U1805 (N_1805,N_435,N_898);
or U1806 (N_1806,In_419,N_970);
xnor U1807 (N_1807,N_741,In_1346);
and U1808 (N_1808,N_518,N_719);
or U1809 (N_1809,N_490,In_2362);
nand U1810 (N_1810,N_1002,N_219);
and U1811 (N_1811,N_115,In_652);
xor U1812 (N_1812,N_661,N_504);
xnor U1813 (N_1813,In_630,N_374);
xor U1814 (N_1814,N_774,N_26);
or U1815 (N_1815,N_446,N_790);
xnor U1816 (N_1816,In_1476,In_1843);
xnor U1817 (N_1817,N_489,In_458);
and U1818 (N_1818,N_102,In_247);
xor U1819 (N_1819,N_27,In_967);
xor U1820 (N_1820,In_925,In_2204);
nor U1821 (N_1821,N_171,N_478);
nand U1822 (N_1822,In_619,N_678);
or U1823 (N_1823,N_416,N_67);
nand U1824 (N_1824,N_485,N_197);
xnor U1825 (N_1825,In_1483,In_1964);
and U1826 (N_1826,N_14,N_338);
nor U1827 (N_1827,N_1041,N_227);
and U1828 (N_1828,In_858,N_832);
and U1829 (N_1829,In_1147,In_1846);
nor U1830 (N_1830,N_468,In_2820);
and U1831 (N_1831,N_114,In_1233);
and U1832 (N_1832,N_254,N_1166);
and U1833 (N_1833,N_519,N_1027);
or U1834 (N_1834,N_1130,In_2897);
or U1835 (N_1835,In_1309,N_1193);
xnor U1836 (N_1836,N_697,In_2380);
nor U1837 (N_1837,N_181,In_2858);
or U1838 (N_1838,N_270,N_165);
or U1839 (N_1839,N_640,N_449);
or U1840 (N_1840,N_453,In_541);
or U1841 (N_1841,N_535,In_58);
and U1842 (N_1842,In_1095,In_23);
and U1843 (N_1843,N_1097,N_362);
nand U1844 (N_1844,N_358,In_774);
nor U1845 (N_1845,N_366,N_247);
nand U1846 (N_1846,N_976,N_156);
and U1847 (N_1847,N_475,In_2787);
xnor U1848 (N_1848,In_822,N_85);
nor U1849 (N_1849,In_2013,N_108);
and U1850 (N_1850,N_403,N_594);
nor U1851 (N_1851,N_258,N_329);
or U1852 (N_1852,In_1223,N_971);
nor U1853 (N_1853,N_694,N_344);
nor U1854 (N_1854,N_1136,N_677);
nand U1855 (N_1855,In_380,N_823);
or U1856 (N_1856,N_551,N_902);
and U1857 (N_1857,N_768,In_2901);
xnor U1858 (N_1858,In_113,N_645);
xnor U1859 (N_1859,N_52,N_294);
xor U1860 (N_1860,N_29,In_2799);
nor U1861 (N_1861,N_636,N_481);
nand U1862 (N_1862,In_2511,In_2135);
nand U1863 (N_1863,In_1867,N_972);
or U1864 (N_1864,N_391,In_1272);
and U1865 (N_1865,N_624,N_938);
and U1866 (N_1866,N_1115,In_837);
xnor U1867 (N_1867,N_1045,N_1057);
xnor U1868 (N_1868,N_857,N_68);
nor U1869 (N_1869,N_749,N_1052);
nor U1870 (N_1870,N_16,In_580);
or U1871 (N_1871,In_2294,N_160);
nand U1872 (N_1872,N_18,In_2688);
xor U1873 (N_1873,N_200,N_278);
or U1874 (N_1874,N_860,N_989);
or U1875 (N_1875,In_1046,In_1965);
nand U1876 (N_1876,N_283,In_155);
nand U1877 (N_1877,In_2299,N_987);
nor U1878 (N_1878,N_917,In_1143);
or U1879 (N_1879,N_733,N_407);
nor U1880 (N_1880,In_1152,N_255);
nand U1881 (N_1881,In_571,In_2894);
or U1882 (N_1882,In_341,N_1051);
xor U1883 (N_1883,N_542,N_1074);
nor U1884 (N_1884,N_1164,N_135);
xnor U1885 (N_1885,In_1709,N_1026);
and U1886 (N_1886,N_1069,In_1999);
nand U1887 (N_1887,N_138,In_2595);
nand U1888 (N_1888,In_891,N_30);
xnor U1889 (N_1889,N_695,N_251);
nand U1890 (N_1890,In_2210,N_776);
nor U1891 (N_1891,In_1403,In_631);
xnor U1892 (N_1892,N_1107,N_321);
or U1893 (N_1893,N_711,N_1171);
nand U1894 (N_1894,In_228,N_747);
nand U1895 (N_1895,N_205,N_176);
or U1896 (N_1896,N_498,N_365);
nor U1897 (N_1897,N_480,In_1150);
or U1898 (N_1898,In_2801,In_1293);
or U1899 (N_1899,N_1044,In_304);
nand U1900 (N_1900,In_2751,N_213);
nand U1901 (N_1901,N_297,N_965);
nand U1902 (N_1902,N_1123,N_225);
nor U1903 (N_1903,N_983,N_1167);
nand U1904 (N_1904,N_1085,N_658);
and U1905 (N_1905,N_532,N_936);
nand U1906 (N_1906,In_355,N_626);
or U1907 (N_1907,In_1705,In_1453);
or U1908 (N_1908,N_1075,N_51);
and U1909 (N_1909,N_786,In_706);
nor U1910 (N_1910,In_357,In_1473);
nor U1911 (N_1911,N_949,N_876);
and U1912 (N_1912,N_209,N_49);
nor U1913 (N_1913,N_1079,N_780);
or U1914 (N_1914,N_90,In_485);
xnor U1915 (N_1915,In_102,In_1960);
and U1916 (N_1916,In_1588,In_1247);
and U1917 (N_1917,N_539,N_5);
nand U1918 (N_1918,N_488,N_796);
or U1919 (N_1919,N_1038,N_691);
and U1920 (N_1920,In_1395,N_699);
xnor U1921 (N_1921,In_2109,In_2094);
and U1922 (N_1922,N_634,In_1323);
and U1923 (N_1923,In_2239,In_519);
nor U1924 (N_1924,N_332,N_1073);
xnor U1925 (N_1925,In_296,N_65);
nor U1926 (N_1926,In_1418,N_530);
and U1927 (N_1927,N_1062,N_804);
xor U1928 (N_1928,N_563,N_368);
nand U1929 (N_1929,N_460,In_1896);
or U1930 (N_1930,In_581,N_312);
nor U1931 (N_1931,In_166,N_739);
or U1932 (N_1932,In_272,In_903);
and U1933 (N_1933,N_757,N_469);
or U1934 (N_1934,N_291,N_651);
nor U1935 (N_1935,N_523,N_113);
or U1936 (N_1936,In_702,In_2729);
nand U1937 (N_1937,N_50,N_198);
xor U1938 (N_1938,N_561,N_819);
or U1939 (N_1939,N_285,N_841);
or U1940 (N_1940,In_1116,N_1101);
nor U1941 (N_1941,N_413,N_473);
nand U1942 (N_1942,N_1102,In_1725);
nand U1943 (N_1943,N_4,In_1613);
and U1944 (N_1944,N_88,N_455);
xor U1945 (N_1945,N_1012,N_908);
or U1946 (N_1946,N_463,N_905);
xor U1947 (N_1947,In_2295,In_2297);
nand U1948 (N_1948,In_2445,N_155);
or U1949 (N_1949,In_2196,N_127);
and U1950 (N_1950,N_21,In_2263);
and U1951 (N_1951,N_148,N_903);
xor U1952 (N_1952,N_262,In_2526);
nand U1953 (N_1953,N_397,N_71);
or U1954 (N_1954,N_43,In_2018);
or U1955 (N_1955,N_239,In_2016);
or U1956 (N_1956,N_723,In_750);
nor U1957 (N_1957,In_1982,N_158);
xor U1958 (N_1958,N_352,In_2519);
or U1959 (N_1959,In_2933,N_1132);
or U1960 (N_1960,N_421,In_126);
nor U1961 (N_1961,N_80,N_629);
xnor U1962 (N_1962,N_1017,In_1979);
or U1963 (N_1963,N_560,N_1055);
nor U1964 (N_1964,N_1139,N_821);
xor U1965 (N_1965,N_602,N_240);
nand U1966 (N_1966,N_7,N_1194);
nor U1967 (N_1967,In_1535,In_2700);
xor U1968 (N_1968,N_1197,N_910);
xor U1969 (N_1969,N_620,N_597);
nor U1970 (N_1970,N_1151,In_983);
or U1971 (N_1971,In_2592,In_1256);
or U1972 (N_1972,In_238,In_2781);
xor U1973 (N_1973,In_86,In_1634);
xor U1974 (N_1974,In_777,N_404);
nor U1975 (N_1975,N_1180,N_91);
xnor U1976 (N_1976,In_2310,In_1136);
or U1977 (N_1977,N_664,In_2847);
nor U1978 (N_1978,In_48,In_118);
or U1979 (N_1979,N_953,In_1536);
xor U1980 (N_1980,In_2256,N_372);
and U1981 (N_1981,In_1130,In_2384);
nor U1982 (N_1982,In_1435,N_268);
nand U1983 (N_1983,N_339,In_2867);
nor U1984 (N_1984,N_822,In_920);
and U1985 (N_1985,N_893,N_892);
or U1986 (N_1986,N_806,N_931);
xor U1987 (N_1987,In_178,N_419);
nor U1988 (N_1988,In_2853,N_540);
xnor U1989 (N_1989,In_1057,N_1019);
or U1990 (N_1990,In_1363,N_866);
xor U1991 (N_1991,N_1112,N_641);
nor U1992 (N_1992,In_855,N_1095);
nor U1993 (N_1993,N_84,In_1696);
xor U1994 (N_1994,In_260,N_203);
or U1995 (N_1995,N_1140,In_1769);
xnor U1996 (N_1996,N_36,In_2927);
xnor U1997 (N_1997,In_2726,N_1076);
xor U1998 (N_1998,N_159,In_910);
xor U1999 (N_1999,N_526,N_886);
xor U2000 (N_2000,N_639,In_47);
nand U2001 (N_2001,N_426,N_414);
or U2002 (N_2002,N_1084,In_2622);
or U2003 (N_2003,In_1680,N_309);
nand U2004 (N_2004,In_833,In_2085);
nor U2005 (N_2005,N_1106,In_2946);
xnor U2006 (N_2006,N_24,N_820);
xor U2007 (N_2007,In_2442,In_2724);
and U2008 (N_2008,N_708,N_559);
nand U2009 (N_2009,N_836,N_157);
nor U2010 (N_2010,In_2848,N_1056);
and U2011 (N_2011,N_503,N_964);
nand U2012 (N_2012,In_1356,N_1022);
nand U2013 (N_2013,N_981,N_77);
or U2014 (N_2014,N_541,N_188);
and U2015 (N_2015,N_773,N_609);
nand U2016 (N_2016,N_514,N_792);
nor U2017 (N_2017,In_2633,N_643);
xnor U2018 (N_2018,N_476,N_562);
and U2019 (N_2019,In_2973,N_827);
nand U2020 (N_2020,N_1036,N_654);
nor U2021 (N_2021,N_515,N_728);
xor U2022 (N_2022,N_633,N_800);
nand U2023 (N_2023,N_73,N_256);
nand U2024 (N_2024,N_92,N_798);
or U2025 (N_2025,N_210,In_2102);
and U2026 (N_2026,In_1141,N_994);
xor U2027 (N_2027,In_2581,N_280);
and U2028 (N_2028,N_187,N_748);
and U2029 (N_2029,N_543,In_734);
and U2030 (N_2030,N_302,In_2656);
nor U2031 (N_2031,N_522,In_2774);
and U2032 (N_2032,In_873,In_225);
or U2033 (N_2033,N_1127,N_471);
xor U2034 (N_2034,N_721,In_1226);
or U2035 (N_2035,In_1071,N_457);
and U2036 (N_2036,N_707,In_1091);
nor U2037 (N_2037,In_2534,N_410);
nand U2038 (N_2038,N_1146,N_1007);
nor U2039 (N_2039,In_1462,In_542);
nor U2040 (N_2040,In_2419,N_429);
and U2041 (N_2041,N_367,N_576);
xor U2042 (N_2042,N_499,In_2115);
xor U2043 (N_2043,In_2124,N_743);
and U2044 (N_2044,N_1025,In_2110);
nand U2045 (N_2045,In_990,N_257);
nor U2046 (N_2046,N_93,In_2830);
and U2047 (N_2047,In_100,N_579);
nand U2048 (N_2048,N_811,N_401);
nor U2049 (N_2049,N_853,N_111);
nor U2050 (N_2050,N_912,In_680);
and U2051 (N_2051,N_568,N_462);
or U2052 (N_2052,N_370,In_2571);
nor U2053 (N_2053,N_887,N_253);
nand U2054 (N_2054,In_508,In_1579);
or U2055 (N_2055,N_59,N_331);
nor U2056 (N_2056,N_236,N_459);
nand U2057 (N_2057,N_162,In_978);
nand U2058 (N_2058,N_441,In_866);
xnor U2059 (N_2059,N_1121,In_1576);
and U2060 (N_2060,In_553,N_1066);
nor U2061 (N_2061,N_211,In_492);
xnor U2062 (N_2062,N_717,In_2605);
nor U2063 (N_2063,In_2492,In_2074);
xnor U2064 (N_2064,N_988,N_682);
and U2065 (N_2065,N_615,N_149);
xor U2066 (N_2066,N_967,In_2982);
xor U2067 (N_2067,N_491,In_195);
nor U2068 (N_2068,N_740,In_1915);
nor U2069 (N_2069,N_922,In_2792);
nor U2070 (N_2070,N_1088,N_376);
nor U2071 (N_2071,N_1061,In_2261);
and U2072 (N_2072,N_1173,In_41);
xor U2073 (N_2073,N_458,N_487);
xnor U2074 (N_2074,N_686,N_565);
or U2075 (N_2075,N_726,In_1351);
xor U2076 (N_2076,N_1150,In_1109);
nand U2077 (N_2077,N_364,N_652);
nor U2078 (N_2078,In_2429,In_1313);
nand U2079 (N_2079,N_759,N_145);
nor U2080 (N_2080,In_1885,N_1092);
and U2081 (N_2081,In_1128,N_848);
nor U2082 (N_2082,N_797,N_442);
xnor U2083 (N_2083,N_817,In_227);
nor U2084 (N_2084,In_182,In_1294);
nor U2085 (N_2085,In_679,N_868);
or U2086 (N_2086,N_572,N_369);
xor U2087 (N_2087,N_174,N_440);
nor U2088 (N_2088,In_2778,N_39);
or U2089 (N_2089,N_729,In_1775);
and U2090 (N_2090,N_947,N_308);
xor U2091 (N_2091,N_921,In_2221);
or U2092 (N_2092,In_1189,N_781);
nor U2093 (N_2093,In_2938,N_586);
or U2094 (N_2094,In_2749,N_669);
nand U2095 (N_2095,N_1091,In_500);
and U2096 (N_2096,N_909,In_2252);
nand U2097 (N_2097,N_193,N_103);
nand U2098 (N_2098,In_2576,N_228);
nor U2099 (N_2099,N_196,In_2660);
or U2100 (N_2100,In_983,N_376);
or U2101 (N_2101,In_47,N_750);
nor U2102 (N_2102,N_493,In_1904);
nand U2103 (N_2103,N_871,N_787);
nor U2104 (N_2104,In_1392,N_153);
and U2105 (N_2105,N_853,N_887);
xnor U2106 (N_2106,N_521,In_1950);
or U2107 (N_2107,In_1054,In_986);
and U2108 (N_2108,N_809,N_307);
nand U2109 (N_2109,N_608,N_398);
xnor U2110 (N_2110,N_1174,N_880);
or U2111 (N_2111,In_1395,In_419);
xnor U2112 (N_2112,N_496,N_305);
nor U2113 (N_2113,In_2199,N_1090);
and U2114 (N_2114,In_2894,N_681);
or U2115 (N_2115,In_2085,N_1018);
or U2116 (N_2116,In_1014,N_479);
or U2117 (N_2117,N_591,In_2894);
or U2118 (N_2118,In_2519,N_533);
nand U2119 (N_2119,In_2157,N_967);
nor U2120 (N_2120,N_692,N_622);
xor U2121 (N_2121,N_569,In_1867);
or U2122 (N_2122,N_203,N_26);
xnor U2123 (N_2123,N_443,N_196);
nand U2124 (N_2124,N_294,N_600);
or U2125 (N_2125,N_180,N_152);
xnor U2126 (N_2126,N_1021,N_789);
and U2127 (N_2127,N_128,In_148);
nor U2128 (N_2128,N_607,N_951);
nand U2129 (N_2129,N_6,N_617);
xnor U2130 (N_2130,N_640,N_218);
nor U2131 (N_2131,In_1929,In_2261);
xor U2132 (N_2132,N_996,N_440);
xor U2133 (N_2133,In_2726,N_1048);
or U2134 (N_2134,N_248,N_838);
nor U2135 (N_2135,N_329,N_468);
nor U2136 (N_2136,N_65,N_22);
and U2137 (N_2137,N_75,In_1040);
nand U2138 (N_2138,N_832,N_1026);
and U2139 (N_2139,N_124,N_621);
or U2140 (N_2140,In_1083,N_40);
nor U2141 (N_2141,N_432,N_344);
nor U2142 (N_2142,N_424,N_657);
xnor U2143 (N_2143,N_176,N_12);
xnor U2144 (N_2144,N_334,In_2622);
nand U2145 (N_2145,N_18,In_2085);
nand U2146 (N_2146,N_990,In_2589);
and U2147 (N_2147,N_734,N_56);
or U2148 (N_2148,N_304,N_570);
and U2149 (N_2149,N_143,In_2595);
and U2150 (N_2150,In_132,In_625);
or U2151 (N_2151,In_2210,N_343);
and U2152 (N_2152,N_1075,N_833);
nor U2153 (N_2153,N_7,N_275);
nand U2154 (N_2154,N_25,In_1904);
xor U2155 (N_2155,N_738,N_877);
or U2156 (N_2156,In_2248,In_1476);
nand U2157 (N_2157,In_1064,N_254);
nor U2158 (N_2158,In_1363,In_571);
xnor U2159 (N_2159,N_521,In_2854);
or U2160 (N_2160,In_2422,N_892);
xor U2161 (N_2161,N_733,N_1007);
and U2162 (N_2162,N_547,N_924);
nor U2163 (N_2163,N_1148,N_256);
or U2164 (N_2164,N_783,N_132);
or U2165 (N_2165,N_874,In_739);
or U2166 (N_2166,N_143,N_331);
and U2167 (N_2167,N_1091,In_2095);
or U2168 (N_2168,In_2927,In_24);
nand U2169 (N_2169,N_347,N_981);
and U2170 (N_2170,N_674,In_1309);
or U2171 (N_2171,N_684,N_769);
or U2172 (N_2172,N_282,N_0);
nand U2173 (N_2173,N_517,N_587);
nand U2174 (N_2174,N_1173,In_2647);
nand U2175 (N_2175,N_516,In_2797);
and U2176 (N_2176,N_687,N_1145);
xor U2177 (N_2177,In_447,In_2310);
xnor U2178 (N_2178,N_1162,N_166);
and U2179 (N_2179,N_1033,N_405);
and U2180 (N_2180,N_460,In_2297);
nor U2181 (N_2181,N_289,N_902);
or U2182 (N_2182,N_298,N_982);
or U2183 (N_2183,N_747,N_382);
or U2184 (N_2184,N_362,In_2100);
nor U2185 (N_2185,N_931,N_1013);
and U2186 (N_2186,N_436,In_1682);
or U2187 (N_2187,N_468,N_558);
xor U2188 (N_2188,In_458,In_1074);
xor U2189 (N_2189,N_63,In_501);
or U2190 (N_2190,N_910,N_930);
nand U2191 (N_2191,N_348,In_1282);
and U2192 (N_2192,N_1137,In_2573);
xor U2193 (N_2193,N_184,N_544);
nor U2194 (N_2194,In_2685,In_1128);
nor U2195 (N_2195,In_2239,N_824);
or U2196 (N_2196,In_1061,N_187);
xor U2197 (N_2197,In_1613,N_338);
and U2198 (N_2198,N_145,N_780);
or U2199 (N_2199,N_329,N_389);
xnor U2200 (N_2200,N_520,N_1052);
or U2201 (N_2201,N_1138,N_939);
and U2202 (N_2202,N_670,N_556);
and U2203 (N_2203,In_2595,N_554);
nand U2204 (N_2204,N_968,In_489);
and U2205 (N_2205,In_1261,N_1038);
nor U2206 (N_2206,N_127,N_239);
xnor U2207 (N_2207,N_655,N_219);
or U2208 (N_2208,N_517,N_811);
and U2209 (N_2209,N_691,N_763);
xnor U2210 (N_2210,N_369,N_903);
xnor U2211 (N_2211,N_1007,N_115);
or U2212 (N_2212,N_652,N_57);
xnor U2213 (N_2213,N_25,N_1192);
xnor U2214 (N_2214,In_1693,N_604);
and U2215 (N_2215,N_665,N_913);
nand U2216 (N_2216,In_1975,N_975);
xor U2217 (N_2217,N_131,In_1430);
or U2218 (N_2218,N_526,N_190);
nand U2219 (N_2219,N_1034,N_252);
xnor U2220 (N_2220,N_397,N_567);
xor U2221 (N_2221,In_166,N_93);
or U2222 (N_2222,N_1007,In_1256);
xnor U2223 (N_2223,In_2950,N_913);
and U2224 (N_2224,In_870,N_593);
and U2225 (N_2225,N_626,N_652);
xor U2226 (N_2226,N_1140,N_566);
and U2227 (N_2227,N_187,In_508);
or U2228 (N_2228,In_2891,In_446);
xnor U2229 (N_2229,N_475,N_723);
and U2230 (N_2230,N_361,N_630);
xnor U2231 (N_2231,In_774,In_2248);
and U2232 (N_2232,N_465,N_892);
or U2233 (N_2233,In_2751,In_654);
and U2234 (N_2234,N_64,In_1750);
or U2235 (N_2235,In_2519,N_503);
xnor U2236 (N_2236,In_1104,In_2523);
and U2237 (N_2237,N_360,N_104);
xor U2238 (N_2238,N_102,N_139);
nor U2239 (N_2239,N_1063,N_107);
nor U2240 (N_2240,N_887,In_1453);
nand U2241 (N_2241,N_92,N_947);
or U2242 (N_2242,N_961,N_1150);
and U2243 (N_2243,N_13,N_392);
xnor U2244 (N_2244,N_486,N_612);
nor U2245 (N_2245,N_855,In_1294);
or U2246 (N_2246,In_1820,N_591);
or U2247 (N_2247,In_2094,In_2933);
nand U2248 (N_2248,N_758,N_241);
nand U2249 (N_2249,N_199,In_2898);
or U2250 (N_2250,N_337,In_398);
and U2251 (N_2251,N_1085,N_57);
nor U2252 (N_2252,N_1071,N_588);
nand U2253 (N_2253,N_67,In_1136);
nand U2254 (N_2254,N_830,N_597);
nor U2255 (N_2255,In_2239,N_670);
and U2256 (N_2256,N_307,N_934);
and U2257 (N_2257,N_290,N_891);
xnor U2258 (N_2258,In_2721,In_2545);
and U2259 (N_2259,N_650,N_972);
nor U2260 (N_2260,N_999,N_1148);
nand U2261 (N_2261,In_1363,N_378);
nor U2262 (N_2262,In_1054,N_1004);
nand U2263 (N_2263,N_486,N_680);
xor U2264 (N_2264,N_799,N_675);
nor U2265 (N_2265,N_711,In_2862);
xor U2266 (N_2266,In_1582,N_37);
nor U2267 (N_2267,In_247,N_663);
and U2268 (N_2268,N_104,In_485);
xor U2269 (N_2269,N_580,In_2534);
nor U2270 (N_2270,N_983,N_60);
nand U2271 (N_2271,In_631,N_93);
and U2272 (N_2272,In_259,N_162);
xnor U2273 (N_2273,N_875,In_1490);
nand U2274 (N_2274,In_2539,N_72);
nand U2275 (N_2275,N_837,N_715);
or U2276 (N_2276,N_993,N_810);
nand U2277 (N_2277,N_1188,N_56);
nor U2278 (N_2278,N_967,N_257);
and U2279 (N_2279,In_2897,N_812);
nor U2280 (N_2280,N_236,In_2947);
nand U2281 (N_2281,In_679,N_951);
or U2282 (N_2282,N_85,In_1223);
or U2283 (N_2283,N_239,In_1680);
xor U2284 (N_2284,N_138,In_1313);
xnor U2285 (N_2285,N_503,N_603);
nand U2286 (N_2286,N_1012,In_381);
nor U2287 (N_2287,In_1083,N_596);
and U2288 (N_2288,N_77,N_253);
and U2289 (N_2289,N_402,N_521);
nor U2290 (N_2290,N_446,In_1365);
or U2291 (N_2291,In_2115,In_2774);
or U2292 (N_2292,In_2419,In_2928);
and U2293 (N_2293,N_755,In_2653);
and U2294 (N_2294,In_631,N_35);
xor U2295 (N_2295,In_2526,N_414);
and U2296 (N_2296,N_604,In_2967);
xnor U2297 (N_2297,N_868,In_2422);
xnor U2298 (N_2298,In_619,N_280);
xor U2299 (N_2299,N_186,N_376);
xnor U2300 (N_2300,In_2115,N_633);
nand U2301 (N_2301,In_762,N_903);
xor U2302 (N_2302,In_1709,N_1016);
nand U2303 (N_2303,N_96,N_258);
nor U2304 (N_2304,In_2688,N_518);
and U2305 (N_2305,N_979,N_499);
and U2306 (N_2306,In_2195,N_351);
nand U2307 (N_2307,N_67,N_742);
or U2308 (N_2308,N_816,N_245);
nand U2309 (N_2309,N_772,In_1064);
xor U2310 (N_2310,In_2256,In_489);
nor U2311 (N_2311,N_889,N_986);
nor U2312 (N_2312,N_988,N_11);
and U2313 (N_2313,N_300,N_719);
xnor U2314 (N_2314,In_259,In_1164);
or U2315 (N_2315,N_1082,N_674);
and U2316 (N_2316,N_155,N_214);
or U2317 (N_2317,N_1047,N_410);
or U2318 (N_2318,N_1080,In_1684);
nor U2319 (N_2319,N_964,N_212);
nor U2320 (N_2320,N_740,In_793);
xor U2321 (N_2321,N_705,N_77);
or U2322 (N_2322,N_349,N_158);
nor U2323 (N_2323,N_674,N_329);
xnor U2324 (N_2324,N_499,N_1158);
nand U2325 (N_2325,In_1579,N_389);
xor U2326 (N_2326,N_1119,N_1019);
nor U2327 (N_2327,N_423,N_852);
nand U2328 (N_2328,N_556,N_150);
nor U2329 (N_2329,N_1163,N_247);
xnor U2330 (N_2330,N_898,N_830);
or U2331 (N_2331,N_816,N_306);
xnor U2332 (N_2332,N_148,In_2200);
nor U2333 (N_2333,N_248,N_593);
nand U2334 (N_2334,N_749,In_1163);
nor U2335 (N_2335,In_380,In_41);
nor U2336 (N_2336,In_919,N_955);
xor U2337 (N_2337,N_961,In_469);
or U2338 (N_2338,N_126,N_266);
nor U2339 (N_2339,N_136,N_1094);
nand U2340 (N_2340,N_567,N_960);
nor U2341 (N_2341,N_464,N_602);
nor U2342 (N_2342,In_1870,In_2661);
or U2343 (N_2343,N_974,N_108);
xnor U2344 (N_2344,N_958,N_759);
nor U2345 (N_2345,N_83,N_622);
nand U2346 (N_2346,In_1808,N_1164);
xnor U2347 (N_2347,N_984,N_53);
xor U2348 (N_2348,N_797,In_903);
and U2349 (N_2349,N_1062,In_178);
nor U2350 (N_2350,N_781,In_1982);
or U2351 (N_2351,N_344,N_688);
xnor U2352 (N_2352,In_2629,In_1680);
and U2353 (N_2353,N_239,N_316);
xnor U2354 (N_2354,N_217,In_750);
nand U2355 (N_2355,In_1846,In_2160);
nand U2356 (N_2356,In_2603,In_2180);
xor U2357 (N_2357,In_355,In_2603);
xnor U2358 (N_2358,In_2725,N_300);
xor U2359 (N_2359,In_319,N_210);
or U2360 (N_2360,N_688,N_997);
xnor U2361 (N_2361,N_1116,N_522);
nand U2362 (N_2362,N_8,N_35);
or U2363 (N_2363,In_118,N_886);
nor U2364 (N_2364,N_566,In_2534);
nor U2365 (N_2365,N_3,In_978);
xnor U2366 (N_2366,In_300,N_385);
or U2367 (N_2367,N_1150,In_2709);
or U2368 (N_2368,N_615,N_356);
and U2369 (N_2369,In_2226,In_2929);
xor U2370 (N_2370,In_1272,N_34);
xnor U2371 (N_2371,N_500,N_950);
xnor U2372 (N_2372,N_380,N_191);
xnor U2373 (N_2373,N_91,N_19);
xor U2374 (N_2374,N_147,In_820);
nand U2375 (N_2375,N_55,N_306);
nand U2376 (N_2376,N_26,N_1083);
or U2377 (N_2377,In_762,N_54);
nand U2378 (N_2378,In_920,In_1757);
nor U2379 (N_2379,N_648,N_981);
or U2380 (N_2380,In_1903,N_951);
nor U2381 (N_2381,N_344,In_679);
and U2382 (N_2382,In_1514,N_405);
nand U2383 (N_2383,N_1196,N_606);
nor U2384 (N_2384,In_1365,N_418);
and U2385 (N_2385,N_581,N_512);
or U2386 (N_2386,In_2678,N_270);
nor U2387 (N_2387,In_1709,N_486);
or U2388 (N_2388,N_1042,In_2263);
xnor U2389 (N_2389,N_806,N_441);
nand U2390 (N_2390,In_1345,In_1040);
or U2391 (N_2391,N_1196,N_1094);
and U2392 (N_2392,N_190,N_31);
or U2393 (N_2393,N_1145,N_50);
nand U2394 (N_2394,N_525,N_967);
and U2395 (N_2395,In_2847,In_2510);
nand U2396 (N_2396,In_2947,N_121);
xor U2397 (N_2397,N_133,In_1472);
nand U2398 (N_2398,N_931,In_458);
nor U2399 (N_2399,N_1151,N_615);
or U2400 (N_2400,N_2354,N_1944);
nor U2401 (N_2401,N_1267,N_1912);
nor U2402 (N_2402,N_1535,N_1402);
nand U2403 (N_2403,N_2343,N_1653);
nor U2404 (N_2404,N_1579,N_2010);
nand U2405 (N_2405,N_1597,N_2009);
nand U2406 (N_2406,N_1308,N_1565);
xor U2407 (N_2407,N_1886,N_1715);
nand U2408 (N_2408,N_2303,N_1992);
xnor U2409 (N_2409,N_1297,N_1950);
and U2410 (N_2410,N_1998,N_1778);
and U2411 (N_2411,N_2129,N_2309);
nor U2412 (N_2412,N_1916,N_1711);
or U2413 (N_2413,N_2295,N_1758);
nor U2414 (N_2414,N_1929,N_1343);
and U2415 (N_2415,N_1456,N_2375);
nand U2416 (N_2416,N_1980,N_1249);
xnor U2417 (N_2417,N_2321,N_1789);
and U2418 (N_2418,N_1207,N_1482);
and U2419 (N_2419,N_2172,N_2358);
or U2420 (N_2420,N_2016,N_1461);
nor U2421 (N_2421,N_2175,N_1364);
and U2422 (N_2422,N_1898,N_1940);
nor U2423 (N_2423,N_2111,N_1312);
xor U2424 (N_2424,N_1558,N_1733);
or U2425 (N_2425,N_1770,N_2152);
xnor U2426 (N_2426,N_2042,N_1477);
or U2427 (N_2427,N_1515,N_1702);
nand U2428 (N_2428,N_1592,N_1787);
or U2429 (N_2429,N_2248,N_1977);
xnor U2430 (N_2430,N_1253,N_2018);
xor U2431 (N_2431,N_2277,N_1652);
and U2432 (N_2432,N_2045,N_1547);
xnor U2433 (N_2433,N_1348,N_2299);
nor U2434 (N_2434,N_2083,N_1559);
nand U2435 (N_2435,N_1372,N_2069);
nor U2436 (N_2436,N_2314,N_1225);
or U2437 (N_2437,N_1208,N_1818);
or U2438 (N_2438,N_1603,N_2229);
or U2439 (N_2439,N_1452,N_2361);
nor U2440 (N_2440,N_1423,N_1393);
or U2441 (N_2441,N_2384,N_1400);
xor U2442 (N_2442,N_1618,N_1917);
or U2443 (N_2443,N_1230,N_1427);
or U2444 (N_2444,N_2266,N_1630);
nor U2445 (N_2445,N_2251,N_1536);
xor U2446 (N_2446,N_1488,N_1808);
xnor U2447 (N_2447,N_2388,N_2119);
nand U2448 (N_2448,N_2164,N_1797);
and U2449 (N_2449,N_1712,N_2139);
xor U2450 (N_2450,N_1451,N_1600);
and U2451 (N_2451,N_2125,N_1700);
nor U2452 (N_2452,N_2256,N_1891);
nand U2453 (N_2453,N_1810,N_1632);
or U2454 (N_2454,N_1594,N_2238);
and U2455 (N_2455,N_1543,N_2262);
or U2456 (N_2456,N_1970,N_1206);
or U2457 (N_2457,N_1305,N_1245);
xor U2458 (N_2458,N_1792,N_2312);
or U2459 (N_2459,N_1324,N_1766);
nand U2460 (N_2460,N_2211,N_2234);
or U2461 (N_2461,N_1760,N_1595);
nand U2462 (N_2462,N_1222,N_1218);
and U2463 (N_2463,N_1649,N_1410);
or U2464 (N_2464,N_1708,N_1280);
or U2465 (N_2465,N_1775,N_2133);
and U2466 (N_2466,N_1752,N_2316);
and U2467 (N_2467,N_2094,N_2052);
nand U2468 (N_2468,N_1448,N_1949);
nand U2469 (N_2469,N_1344,N_2027);
nor U2470 (N_2470,N_1593,N_1602);
xnor U2471 (N_2471,N_1415,N_1954);
nand U2472 (N_2472,N_2216,N_2392);
or U2473 (N_2473,N_1391,N_2143);
xor U2474 (N_2474,N_1417,N_1303);
nand U2475 (N_2475,N_2379,N_1441);
nor U2476 (N_2476,N_1633,N_2031);
and U2477 (N_2477,N_2174,N_1825);
nor U2478 (N_2478,N_2285,N_2260);
xor U2479 (N_2479,N_2193,N_1588);
or U2480 (N_2480,N_1832,N_2291);
or U2481 (N_2481,N_1629,N_1378);
nand U2482 (N_2482,N_2037,N_1573);
and U2483 (N_2483,N_1903,N_1861);
nor U2484 (N_2484,N_2134,N_2236);
nand U2485 (N_2485,N_1566,N_2355);
nor U2486 (N_2486,N_2104,N_1691);
and U2487 (N_2487,N_2160,N_1822);
and U2488 (N_2488,N_1676,N_2223);
nor U2489 (N_2489,N_1354,N_2386);
nor U2490 (N_2490,N_1377,N_2186);
or U2491 (N_2491,N_2398,N_1533);
and U2492 (N_2492,N_1576,N_2023);
nand U2493 (N_2493,N_1902,N_1921);
and U2494 (N_2494,N_1498,N_1826);
and U2495 (N_2495,N_1495,N_2092);
or U2496 (N_2496,N_1295,N_1741);
nand U2497 (N_2497,N_1472,N_2212);
nor U2498 (N_2498,N_2363,N_2300);
or U2499 (N_2499,N_2353,N_1754);
and U2500 (N_2500,N_1358,N_2207);
xor U2501 (N_2501,N_1981,N_1635);
or U2502 (N_2502,N_1731,N_1663);
nand U2503 (N_2503,N_2304,N_1835);
or U2504 (N_2504,N_1529,N_2327);
nand U2505 (N_2505,N_2219,N_1571);
nand U2506 (N_2506,N_1336,N_1221);
and U2507 (N_2507,N_1493,N_1746);
nand U2508 (N_2508,N_1900,N_1394);
or U2509 (N_2509,N_1985,N_1881);
xor U2510 (N_2510,N_1743,N_2153);
nor U2511 (N_2511,N_1580,N_2073);
xor U2512 (N_2512,N_1445,N_1233);
nand U2513 (N_2513,N_1931,N_1475);
nor U2514 (N_2514,N_1436,N_1729);
nor U2515 (N_2515,N_1260,N_1425);
xnor U2516 (N_2516,N_2096,N_1335);
and U2517 (N_2517,N_1721,N_1266);
and U2518 (N_2518,N_2043,N_1480);
and U2519 (N_2519,N_1310,N_2306);
and U2520 (N_2520,N_2012,N_1933);
and U2521 (N_2521,N_1341,N_1447);
nand U2522 (N_2522,N_1357,N_1627);
or U2523 (N_2523,N_1411,N_1901);
and U2524 (N_2524,N_1544,N_1730);
nor U2525 (N_2525,N_2350,N_1673);
nand U2526 (N_2526,N_2039,N_1925);
xor U2527 (N_2527,N_1512,N_2025);
nand U2528 (N_2528,N_2318,N_1859);
nand U2529 (N_2529,N_1942,N_1965);
or U2530 (N_2530,N_1522,N_1621);
or U2531 (N_2531,N_2197,N_2278);
or U2532 (N_2532,N_1928,N_1203);
xor U2533 (N_2533,N_1761,N_1874);
or U2534 (N_2534,N_2249,N_1323);
and U2535 (N_2535,N_2372,N_2368);
xnor U2536 (N_2536,N_2336,N_1385);
nor U2537 (N_2537,N_1459,N_1416);
xor U2538 (N_2538,N_1922,N_1541);
nand U2539 (N_2539,N_1785,N_2138);
or U2540 (N_2540,N_2100,N_1418);
and U2541 (N_2541,N_1413,N_1687);
and U2542 (N_2542,N_1604,N_1392);
nand U2543 (N_2543,N_1705,N_2187);
or U2544 (N_2544,N_1484,N_1888);
and U2545 (N_2545,N_1894,N_1987);
or U2546 (N_2546,N_1867,N_2275);
or U2547 (N_2547,N_1626,N_1375);
xor U2548 (N_2548,N_1241,N_1381);
or U2549 (N_2549,N_1382,N_1285);
xor U2550 (N_2550,N_1742,N_2032);
or U2551 (N_2551,N_1899,N_2188);
and U2552 (N_2552,N_2021,N_1283);
nor U2553 (N_2553,N_2163,N_1645);
xor U2554 (N_2554,N_1855,N_1470);
nand U2555 (N_2555,N_2381,N_1848);
nor U2556 (N_2556,N_2024,N_2245);
nand U2557 (N_2557,N_1856,N_2036);
or U2558 (N_2558,N_1857,N_2099);
nand U2559 (N_2559,N_1707,N_2078);
and U2560 (N_2560,N_1257,N_1596);
or U2561 (N_2561,N_1246,N_1306);
or U2562 (N_2562,N_2206,N_2136);
and U2563 (N_2563,N_1293,N_2101);
or U2564 (N_2564,N_1804,N_1386);
nor U2565 (N_2565,N_1564,N_1973);
nand U2566 (N_2566,N_1226,N_1767);
or U2567 (N_2567,N_1947,N_1232);
xor U2568 (N_2568,N_1757,N_2151);
nor U2569 (N_2569,N_1732,N_2272);
or U2570 (N_2570,N_1248,N_2185);
and U2571 (N_2571,N_1548,N_1585);
xor U2572 (N_2572,N_1996,N_2259);
xnor U2573 (N_2573,N_1780,N_1842);
and U2574 (N_2574,N_1771,N_1840);
nor U2575 (N_2575,N_2017,N_2086);
and U2576 (N_2576,N_2098,N_1224);
or U2577 (N_2577,N_1332,N_1525);
xor U2578 (N_2578,N_1943,N_1955);
nand U2579 (N_2579,N_1816,N_2268);
or U2580 (N_2580,N_1471,N_2195);
nor U2581 (N_2581,N_1279,N_2257);
nor U2582 (N_2582,N_2061,N_1667);
and U2583 (N_2583,N_2367,N_1419);
xor U2584 (N_2584,N_1318,N_2054);
nand U2585 (N_2585,N_1750,N_1795);
and U2586 (N_2586,N_1836,N_2399);
nor U2587 (N_2587,N_2385,N_2250);
and U2588 (N_2588,N_1906,N_2141);
or U2589 (N_2589,N_2351,N_1969);
nand U2590 (N_2590,N_1510,N_1328);
xnor U2591 (N_2591,N_2233,N_1496);
xnor U2592 (N_2592,N_1674,N_1647);
nand U2593 (N_2593,N_2040,N_1317);
xor U2594 (N_2594,N_1744,N_2357);
or U2595 (N_2595,N_1424,N_1869);
nor U2596 (N_2596,N_1607,N_1932);
or U2597 (N_2597,N_1827,N_2371);
nand U2598 (N_2598,N_1934,N_2204);
nand U2599 (N_2599,N_2217,N_1429);
or U2600 (N_2600,N_1964,N_1453);
xnor U2601 (N_2601,N_2289,N_1408);
nand U2602 (N_2602,N_1952,N_1262);
nor U2603 (N_2603,N_1569,N_2364);
and U2604 (N_2604,N_1514,N_2106);
and U2605 (N_2605,N_1399,N_2062);
or U2606 (N_2606,N_1777,N_2166);
nand U2607 (N_2607,N_1374,N_1698);
nor U2608 (N_2608,N_1763,N_1736);
or U2609 (N_2609,N_2382,N_1956);
nor U2610 (N_2610,N_1269,N_2270);
and U2611 (N_2611,N_1586,N_1352);
xnor U2612 (N_2612,N_2057,N_1613);
xor U2613 (N_2613,N_1554,N_1885);
or U2614 (N_2614,N_2090,N_1682);
and U2615 (N_2615,N_2243,N_2342);
nor U2616 (N_2616,N_1422,N_1745);
xor U2617 (N_2617,N_1738,N_2019);
or U2618 (N_2618,N_1572,N_1255);
and U2619 (N_2619,N_1551,N_1656);
or U2620 (N_2620,N_1521,N_1365);
xor U2621 (N_2621,N_1534,N_1718);
xor U2622 (N_2622,N_1575,N_1923);
xnor U2623 (N_2623,N_1710,N_1237);
or U2624 (N_2624,N_1974,N_2228);
or U2625 (N_2625,N_1713,N_2003);
xor U2626 (N_2626,N_2394,N_1622);
nand U2627 (N_2627,N_2297,N_1466);
nor U2628 (N_2628,N_2205,N_1908);
nor U2629 (N_2629,N_2066,N_1839);
nand U2630 (N_2630,N_2264,N_2232);
and U2631 (N_2631,N_1948,N_2047);
or U2632 (N_2632,N_1847,N_1798);
and U2633 (N_2633,N_1236,N_1568);
xnor U2634 (N_2634,N_2352,N_1567);
and U2635 (N_2635,N_1314,N_2029);
nand U2636 (N_2636,N_2183,N_1578);
nand U2637 (N_2637,N_1937,N_1537);
nand U2638 (N_2638,N_1990,N_1824);
or U2639 (N_2639,N_1539,N_1485);
and U2640 (N_2640,N_1759,N_1722);
nand U2641 (N_2641,N_1409,N_1945);
xor U2642 (N_2642,N_1963,N_2209);
nor U2643 (N_2643,N_1388,N_1489);
and U2644 (N_2644,N_2286,N_1258);
nand U2645 (N_2645,N_1774,N_1939);
or U2646 (N_2646,N_1250,N_2079);
and U2647 (N_2647,N_1333,N_1214);
xnor U2648 (N_2648,N_2390,N_1251);
and U2649 (N_2649,N_2004,N_1756);
and U2650 (N_2650,N_1773,N_2137);
nand U2651 (N_2651,N_2144,N_1697);
and U2652 (N_2652,N_1984,N_2146);
xor U2653 (N_2653,N_2269,N_1628);
xnor U2654 (N_2654,N_2159,N_1648);
and U2655 (N_2655,N_2180,N_1930);
xnor U2656 (N_2656,N_2051,N_1611);
xor U2657 (N_2657,N_1864,N_2347);
nand U2658 (N_2658,N_1844,N_2189);
xnor U2659 (N_2659,N_1669,N_1666);
or U2660 (N_2660,N_1693,N_1644);
and U2661 (N_2661,N_2080,N_2389);
or U2662 (N_2662,N_1538,N_1696);
nor U2663 (N_2663,N_1846,N_1342);
nor U2664 (N_2664,N_1871,N_1454);
and U2665 (N_2665,N_1972,N_1728);
and U2666 (N_2666,N_1828,N_1499);
nand U2667 (N_2667,N_1264,N_1820);
nand U2668 (N_2668,N_2377,N_2328);
and U2669 (N_2669,N_1866,N_2182);
or U2670 (N_2670,N_1369,N_1806);
nor U2671 (N_2671,N_1662,N_2369);
xor U2672 (N_2672,N_1803,N_2201);
nand U2673 (N_2673,N_1527,N_1234);
nor U2674 (N_2674,N_1706,N_1443);
xor U2675 (N_2675,N_1877,N_1805);
nor U2676 (N_2676,N_1389,N_1716);
nor U2677 (N_2677,N_1300,N_1455);
nor U2678 (N_2678,N_2356,N_2091);
xnor U2679 (N_2679,N_2127,N_1503);
or U2680 (N_2680,N_1468,N_1583);
or U2681 (N_2681,N_2199,N_2178);
nand U2682 (N_2682,N_1502,N_1213);
nand U2683 (N_2683,N_1688,N_1247);
and U2684 (N_2684,N_1720,N_1494);
and U2685 (N_2685,N_1617,N_2114);
or U2686 (N_2686,N_1670,N_2282);
nand U2687 (N_2687,N_1403,N_2341);
or U2688 (N_2688,N_2165,N_1740);
or U2689 (N_2689,N_2319,N_1360);
and U2690 (N_2690,N_2022,N_1244);
nand U2691 (N_2691,N_2097,N_1426);
nor U2692 (N_2692,N_1265,N_1909);
nor U2693 (N_2693,N_1227,N_1353);
nand U2694 (N_2694,N_1788,N_1776);
nor U2695 (N_2695,N_2184,N_1723);
and U2696 (N_2696,N_1813,N_2373);
xor U2697 (N_2697,N_2161,N_1914);
xnor U2698 (N_2698,N_1517,N_1887);
or U2699 (N_2699,N_1675,N_1557);
xor U2700 (N_2700,N_2095,N_1833);
nor U2701 (N_2701,N_1790,N_1555);
nand U2702 (N_2702,N_1272,N_1434);
nand U2703 (N_2703,N_2064,N_1211);
or U2704 (N_2704,N_2391,N_1988);
and U2705 (N_2705,N_1467,N_1817);
xnor U2706 (N_2706,N_1487,N_2005);
nand U2707 (N_2707,N_1997,N_1420);
nand U2708 (N_2708,N_2240,N_1202);
and U2709 (N_2709,N_1508,N_1714);
nand U2710 (N_2710,N_1524,N_1542);
xor U2711 (N_2711,N_2340,N_1892);
nor U2712 (N_2712,N_1681,N_1589);
nand U2713 (N_2713,N_1646,N_1680);
nand U2714 (N_2714,N_2322,N_1811);
and U2715 (N_2715,N_1958,N_1553);
xor U2716 (N_2716,N_1546,N_2044);
or U2717 (N_2717,N_1500,N_2276);
xnor U2718 (N_2718,N_1384,N_1768);
nor U2719 (N_2719,N_2292,N_1501);
xor U2720 (N_2720,N_1747,N_1699);
and U2721 (N_2721,N_1296,N_1860);
and U2722 (N_2722,N_1347,N_1562);
nand U2723 (N_2723,N_1240,N_1291);
or U2724 (N_2724,N_1404,N_2181);
nand U2725 (N_2725,N_1516,N_2013);
nand U2726 (N_2726,N_2162,N_1220);
nor U2727 (N_2727,N_1946,N_1582);
nand U2728 (N_2728,N_2337,N_2107);
nand U2729 (N_2729,N_1229,N_2030);
nor U2730 (N_2730,N_1528,N_1913);
nor U2731 (N_2731,N_1651,N_1753);
or U2732 (N_2732,N_1837,N_2071);
nor U2733 (N_2733,N_1491,N_1563);
and U2734 (N_2734,N_2123,N_1560);
xnor U2735 (N_2735,N_1363,N_1590);
nand U2736 (N_2736,N_1412,N_1276);
and U2737 (N_2737,N_2171,N_2124);
xor U2738 (N_2738,N_2192,N_1793);
or U2739 (N_2739,N_1725,N_2068);
and U2740 (N_2740,N_1504,N_1879);
or U2741 (N_2741,N_1889,N_1277);
and U2742 (N_2742,N_1823,N_1918);
nor U2743 (N_2743,N_1966,N_1853);
nand U2744 (N_2744,N_1460,N_1625);
xnor U2745 (N_2745,N_1786,N_2049);
xor U2746 (N_2746,N_2370,N_2215);
xor U2747 (N_2747,N_1330,N_1406);
nor U2748 (N_2748,N_2033,N_2102);
or U2749 (N_2749,N_2169,N_2158);
nand U2750 (N_2750,N_2378,N_2315);
or U2751 (N_2751,N_1339,N_1978);
nor U2752 (N_2752,N_2105,N_2235);
xor U2753 (N_2753,N_1637,N_2084);
or U2754 (N_2754,N_2149,N_1371);
xnor U2755 (N_2755,N_1897,N_2220);
and U2756 (N_2756,N_2231,N_1672);
xor U2757 (N_2757,N_2271,N_1668);
nor U2758 (N_2758,N_1684,N_1801);
nor U2759 (N_2759,N_2121,N_1623);
xnor U2760 (N_2760,N_1709,N_1338);
or U2761 (N_2761,N_2082,N_2011);
xnor U2762 (N_2762,N_1995,N_2020);
xor U2763 (N_2763,N_1830,N_1307);
and U2764 (N_2764,N_1319,N_1976);
nand U2765 (N_2765,N_2148,N_1320);
nor U2766 (N_2766,N_1254,N_1507);
nor U2767 (N_2767,N_2311,N_1421);
nand U2768 (N_2768,N_1215,N_1858);
and U2769 (N_2769,N_1380,N_2001);
nor U2770 (N_2770,N_1938,N_1390);
xor U2771 (N_2771,N_2065,N_1911);
nand U2772 (N_2772,N_2307,N_2281);
or U2773 (N_2773,N_1959,N_1287);
and U2774 (N_2774,N_1896,N_2155);
nor U2775 (N_2775,N_1231,N_1549);
and U2776 (N_2776,N_1610,N_2150);
nand U2777 (N_2777,N_1642,N_2335);
and U2778 (N_2778,N_1446,N_1634);
nor U2779 (N_2779,N_2075,N_2214);
nand U2780 (N_2780,N_2239,N_1289);
xor U2781 (N_2781,N_2060,N_1552);
nor U2782 (N_2782,N_1657,N_1373);
or U2783 (N_2783,N_1505,N_1658);
nor U2784 (N_2784,N_2313,N_1337);
xor U2785 (N_2785,N_1935,N_2128);
and U2786 (N_2786,N_2059,N_1368);
nor U2787 (N_2787,N_1994,N_1523);
or U2788 (N_2788,N_2048,N_1927);
or U2789 (N_2789,N_1288,N_2323);
and U2790 (N_2790,N_1719,N_1986);
xor U2791 (N_2791,N_1735,N_2374);
nor U2792 (N_2792,N_2331,N_1953);
and U2793 (N_2793,N_1762,N_1217);
nor U2794 (N_2794,N_2122,N_2326);
nand U2795 (N_2795,N_1216,N_1812);
and U2796 (N_2796,N_2140,N_1821);
or U2797 (N_2797,N_1481,N_1252);
or U2798 (N_2798,N_1957,N_1960);
and U2799 (N_2799,N_2387,N_1870);
nor U2800 (N_2800,N_1263,N_1270);
and U2801 (N_2801,N_1298,N_1407);
and U2802 (N_2802,N_2274,N_2147);
or U2803 (N_2803,N_1614,N_1570);
nor U2804 (N_2804,N_2261,N_2000);
xnor U2805 (N_2805,N_1223,N_2273);
nand U2806 (N_2806,N_1431,N_1556);
and U2807 (N_2807,N_1587,N_1704);
nor U2808 (N_2808,N_1598,N_1619);
nor U2809 (N_2809,N_1641,N_2076);
nor U2810 (N_2810,N_1796,N_2063);
nand U2811 (N_2811,N_2190,N_1606);
and U2812 (N_2812,N_2208,N_2310);
and U2813 (N_2813,N_2108,N_2093);
or U2814 (N_2814,N_1506,N_2298);
nor U2815 (N_2815,N_2154,N_1545);
nand U2816 (N_2816,N_1784,N_1450);
nor U2817 (N_2817,N_2288,N_1346);
nand U2818 (N_2818,N_1281,N_2324);
nor U2819 (N_2819,N_1640,N_2296);
and U2820 (N_2820,N_1999,N_1904);
nor U2821 (N_2821,N_1726,N_1694);
nor U2822 (N_2822,N_2002,N_2202);
nand U2823 (N_2823,N_1791,N_2284);
nand U2824 (N_2824,N_1638,N_1851);
nor U2825 (N_2825,N_2007,N_1852);
nor U2826 (N_2826,N_2074,N_1239);
nand U2827 (N_2827,N_1893,N_2346);
nand U2828 (N_2828,N_1609,N_1843);
xnor U2829 (N_2829,N_2087,N_1993);
and U2830 (N_2830,N_1275,N_2191);
xor U2831 (N_2831,N_1863,N_1478);
nand U2832 (N_2832,N_1794,N_1463);
nand U2833 (N_2833,N_1951,N_1620);
xnor U2834 (N_2834,N_1340,N_2302);
and U2835 (N_2835,N_1316,N_2041);
nand U2836 (N_2836,N_2058,N_1301);
xnor U2837 (N_2837,N_1398,N_2227);
and U2838 (N_2838,N_1473,N_2305);
or U2839 (N_2839,N_1321,N_2308);
and U2840 (N_2840,N_2397,N_2120);
and U2841 (N_2841,N_1854,N_2067);
or U2842 (N_2842,N_2330,N_2258);
or U2843 (N_2843,N_1469,N_1361);
xnor U2844 (N_2844,N_1474,N_2246);
nand U2845 (N_2845,N_1261,N_1437);
or U2846 (N_2846,N_1772,N_1540);
nor U2847 (N_2847,N_1873,N_2225);
xor U2848 (N_2848,N_2349,N_1397);
nor U2849 (N_2849,N_1350,N_1751);
nor U2850 (N_2850,N_2131,N_1615);
and U2851 (N_2851,N_1574,N_2116);
xor U2852 (N_2852,N_2365,N_1961);
or U2853 (N_2853,N_1329,N_1290);
nand U2854 (N_2854,N_2038,N_1677);
nor U2855 (N_2855,N_1243,N_1802);
nor U2856 (N_2856,N_2213,N_1238);
nand U2857 (N_2857,N_1479,N_1414);
and U2858 (N_2858,N_1880,N_1210);
and U2859 (N_2859,N_1345,N_2115);
nor U2860 (N_2860,N_2173,N_1692);
nor U2861 (N_2861,N_1660,N_2015);
and U2862 (N_2862,N_1204,N_1513);
and U2863 (N_2863,N_2203,N_1490);
nor U2864 (N_2864,N_2109,N_1807);
and U2865 (N_2865,N_1483,N_2253);
xor U2866 (N_2866,N_1862,N_2218);
xnor U2867 (N_2867,N_2334,N_1616);
and U2868 (N_2868,N_2376,N_1727);
or U2869 (N_2869,N_1608,N_1520);
xor U2870 (N_2870,N_2026,N_2055);
and U2871 (N_2871,N_2194,N_2383);
xnor U2872 (N_2872,N_2301,N_2126);
and U2873 (N_2873,N_1286,N_1430);
nand U2874 (N_2874,N_1282,N_1591);
nor U2875 (N_2875,N_2293,N_1829);
nand U2876 (N_2876,N_1865,N_1313);
nand U2877 (N_2877,N_1351,N_2221);
nand U2878 (N_2878,N_1268,N_1878);
or U2879 (N_2879,N_1831,N_1359);
nand U2880 (N_2880,N_1650,N_1433);
nand U2881 (N_2881,N_2283,N_2226);
nor U2882 (N_2882,N_1782,N_2333);
nand U2883 (N_2883,N_2196,N_1737);
and U2884 (N_2884,N_2339,N_2089);
nor U2885 (N_2885,N_2252,N_1331);
xor U2886 (N_2886,N_1671,N_1205);
xnor U2887 (N_2887,N_1876,N_1294);
nor U2888 (N_2888,N_1967,N_2396);
xnor U2889 (N_2889,N_2360,N_2263);
and U2890 (N_2890,N_2070,N_1284);
nor U2891 (N_2891,N_1631,N_1497);
nand U2892 (N_2892,N_1882,N_2035);
or U2893 (N_2893,N_2279,N_1449);
xnor U2894 (N_2894,N_2198,N_1532);
or U2895 (N_2895,N_2244,N_1356);
or U2896 (N_2896,N_1884,N_1868);
nand U2897 (N_2897,N_1936,N_2380);
and U2898 (N_2898,N_1654,N_2362);
xor U2899 (N_2899,N_1685,N_1201);
nand U2900 (N_2900,N_2014,N_1428);
or U2901 (N_2901,N_1850,N_1924);
nor U2902 (N_2902,N_2088,N_1905);
nor U2903 (N_2903,N_1519,N_1926);
nor U2904 (N_2904,N_1326,N_1432);
nand U2905 (N_2905,N_1561,N_1971);
or U2906 (N_2906,N_1370,N_2338);
and U2907 (N_2907,N_2179,N_1975);
or U2908 (N_2908,N_1815,N_2028);
and U2909 (N_2909,N_2177,N_2085);
or U2910 (N_2910,N_1781,N_1989);
and U2911 (N_2911,N_1678,N_2320);
xor U2912 (N_2912,N_2113,N_1783);
or U2913 (N_2913,N_1531,N_1883);
or U2914 (N_2914,N_1376,N_1509);
and U2915 (N_2915,N_2034,N_1695);
nor U2916 (N_2916,N_1349,N_2008);
xor U2917 (N_2917,N_1438,N_2393);
or U2918 (N_2918,N_2265,N_1442);
or U2919 (N_2919,N_1259,N_1299);
nor U2920 (N_2920,N_2344,N_2135);
nor U2921 (N_2921,N_1486,N_1439);
or U2922 (N_2922,N_1809,N_1362);
nand U2923 (N_2923,N_1612,N_1749);
or U2924 (N_2924,N_1209,N_1465);
or U2925 (N_2925,N_2345,N_1895);
and U2926 (N_2926,N_1395,N_1550);
or U2927 (N_2927,N_1962,N_2294);
xor U2928 (N_2928,N_2222,N_1584);
xnor U2929 (N_2929,N_1366,N_2130);
or U2930 (N_2930,N_2046,N_2329);
nor U2931 (N_2931,N_1982,N_2053);
nand U2932 (N_2932,N_1689,N_2237);
xnor U2933 (N_2933,N_1511,N_1387);
nor U2934 (N_2934,N_1779,N_2224);
nor U2935 (N_2935,N_1703,N_2081);
and U2936 (N_2936,N_1665,N_1383);
nand U2937 (N_2937,N_1683,N_2132);
nand U2938 (N_2938,N_1405,N_1636);
or U2939 (N_2939,N_1581,N_1769);
or U2940 (N_2940,N_1526,N_1872);
xnor U2941 (N_2941,N_1764,N_2117);
xnor U2942 (N_2942,N_1800,N_1601);
nand U2943 (N_2943,N_1910,N_1661);
nor U2944 (N_2944,N_2254,N_1664);
xnor U2945 (N_2945,N_2242,N_1492);
nand U2946 (N_2946,N_2267,N_2395);
and U2947 (N_2947,N_2112,N_1274);
nand U2948 (N_2948,N_2056,N_2167);
nand U2949 (N_2949,N_1396,N_1941);
xnor U2950 (N_2950,N_1799,N_1212);
and U2951 (N_2951,N_2247,N_1278);
and U2952 (N_2952,N_1577,N_2118);
and U2953 (N_2953,N_1219,N_1235);
nand U2954 (N_2954,N_1679,N_1435);
or U2955 (N_2955,N_1273,N_2359);
and U2956 (N_2956,N_1302,N_1462);
nor U2957 (N_2957,N_1849,N_2168);
and U2958 (N_2958,N_2287,N_1327);
or U2959 (N_2959,N_1686,N_1890);
or U2960 (N_2960,N_1228,N_2317);
xor U2961 (N_2961,N_1271,N_1367);
nand U2962 (N_2962,N_1518,N_1325);
or U2963 (N_2963,N_2200,N_1690);
or U2964 (N_2964,N_1915,N_1643);
xnor U2965 (N_2965,N_1464,N_2077);
and U2966 (N_2966,N_1717,N_2145);
nand U2967 (N_2967,N_2050,N_2156);
nand U2968 (N_2968,N_1379,N_2142);
and U2969 (N_2969,N_2110,N_1919);
or U2970 (N_2970,N_2348,N_2157);
or U2971 (N_2971,N_1907,N_1920);
nor U2972 (N_2972,N_1624,N_2280);
and U2973 (N_2973,N_2170,N_2325);
or U2974 (N_2974,N_1355,N_1599);
nand U2975 (N_2975,N_2241,N_1765);
nand U2976 (N_2976,N_1444,N_1322);
or U2977 (N_2977,N_1979,N_1814);
and U2978 (N_2978,N_1983,N_1991);
or U2979 (N_2979,N_1819,N_2230);
or U2980 (N_2980,N_1701,N_1311);
or U2981 (N_2981,N_1841,N_2176);
nand U2982 (N_2982,N_1875,N_1605);
xnor U2983 (N_2983,N_1834,N_1457);
xnor U2984 (N_2984,N_1292,N_2366);
and U2985 (N_2985,N_2103,N_1401);
xor U2986 (N_2986,N_1458,N_2332);
and U2987 (N_2987,N_2255,N_1659);
or U2988 (N_2988,N_1748,N_1315);
nor U2989 (N_2989,N_1845,N_1755);
or U2990 (N_2990,N_1968,N_2210);
nor U2991 (N_2991,N_2006,N_1639);
and U2992 (N_2992,N_1476,N_1739);
xnor U2993 (N_2993,N_1309,N_1304);
or U2994 (N_2994,N_1440,N_1242);
nor U2995 (N_2995,N_1655,N_2072);
or U2996 (N_2996,N_1530,N_2290);
xor U2997 (N_2997,N_1256,N_1724);
and U2998 (N_2998,N_1734,N_1838);
and U2999 (N_2999,N_1334,N_1200);
or U3000 (N_3000,N_2206,N_1862);
nor U3001 (N_3001,N_1774,N_1836);
nor U3002 (N_3002,N_1462,N_1671);
nand U3003 (N_3003,N_1498,N_1468);
nand U3004 (N_3004,N_1322,N_1503);
and U3005 (N_3005,N_2036,N_2396);
or U3006 (N_3006,N_1247,N_1463);
xnor U3007 (N_3007,N_1989,N_1209);
or U3008 (N_3008,N_1495,N_2363);
or U3009 (N_3009,N_1343,N_1778);
or U3010 (N_3010,N_2009,N_1499);
nor U3011 (N_3011,N_2245,N_1500);
xnor U3012 (N_3012,N_1583,N_1602);
and U3013 (N_3013,N_1756,N_1738);
xnor U3014 (N_3014,N_2075,N_2140);
or U3015 (N_3015,N_1371,N_1782);
and U3016 (N_3016,N_1419,N_1989);
or U3017 (N_3017,N_1871,N_2079);
nor U3018 (N_3018,N_2359,N_1541);
xor U3019 (N_3019,N_1973,N_1823);
or U3020 (N_3020,N_2154,N_2331);
nand U3021 (N_3021,N_2204,N_2077);
nand U3022 (N_3022,N_2342,N_1290);
nand U3023 (N_3023,N_1234,N_2041);
and U3024 (N_3024,N_1297,N_1938);
or U3025 (N_3025,N_2024,N_2107);
or U3026 (N_3026,N_2022,N_1824);
xnor U3027 (N_3027,N_1958,N_1418);
and U3028 (N_3028,N_1352,N_1406);
nand U3029 (N_3029,N_1923,N_1924);
nor U3030 (N_3030,N_2294,N_1593);
and U3031 (N_3031,N_2205,N_2240);
xnor U3032 (N_3032,N_1859,N_1362);
nand U3033 (N_3033,N_1952,N_2105);
nor U3034 (N_3034,N_1661,N_1938);
nor U3035 (N_3035,N_1256,N_2372);
nand U3036 (N_3036,N_1954,N_1484);
and U3037 (N_3037,N_2375,N_2176);
and U3038 (N_3038,N_2152,N_2248);
xnor U3039 (N_3039,N_2239,N_2163);
xnor U3040 (N_3040,N_1820,N_2312);
nor U3041 (N_3041,N_1283,N_1899);
or U3042 (N_3042,N_1394,N_2394);
nand U3043 (N_3043,N_1243,N_1285);
and U3044 (N_3044,N_1973,N_1744);
nor U3045 (N_3045,N_1850,N_1441);
nand U3046 (N_3046,N_2163,N_1612);
and U3047 (N_3047,N_1605,N_1650);
or U3048 (N_3048,N_1489,N_1690);
nand U3049 (N_3049,N_2011,N_1713);
or U3050 (N_3050,N_2186,N_2075);
and U3051 (N_3051,N_1485,N_1829);
or U3052 (N_3052,N_1736,N_1600);
and U3053 (N_3053,N_1676,N_2304);
nand U3054 (N_3054,N_1431,N_1250);
or U3055 (N_3055,N_1791,N_1745);
xnor U3056 (N_3056,N_1822,N_2015);
nand U3057 (N_3057,N_2108,N_1882);
xor U3058 (N_3058,N_1225,N_2025);
or U3059 (N_3059,N_2181,N_1491);
nand U3060 (N_3060,N_2301,N_1369);
and U3061 (N_3061,N_1680,N_1665);
xor U3062 (N_3062,N_2098,N_2052);
nand U3063 (N_3063,N_1465,N_1676);
nand U3064 (N_3064,N_1655,N_1258);
nor U3065 (N_3065,N_2284,N_2111);
or U3066 (N_3066,N_2338,N_2387);
nor U3067 (N_3067,N_1905,N_1973);
nor U3068 (N_3068,N_2371,N_1320);
or U3069 (N_3069,N_1588,N_1348);
nor U3070 (N_3070,N_2157,N_1912);
nor U3071 (N_3071,N_1369,N_1459);
and U3072 (N_3072,N_1945,N_1778);
nand U3073 (N_3073,N_1304,N_1421);
nand U3074 (N_3074,N_1944,N_2386);
xnor U3075 (N_3075,N_1614,N_2270);
nor U3076 (N_3076,N_1922,N_1870);
xnor U3077 (N_3077,N_1704,N_1287);
xor U3078 (N_3078,N_1730,N_1828);
nand U3079 (N_3079,N_1463,N_2084);
nand U3080 (N_3080,N_2241,N_1977);
nor U3081 (N_3081,N_2255,N_2336);
xor U3082 (N_3082,N_1418,N_1489);
nor U3083 (N_3083,N_1716,N_2200);
nor U3084 (N_3084,N_1628,N_1928);
xor U3085 (N_3085,N_2079,N_1586);
xnor U3086 (N_3086,N_1390,N_1853);
and U3087 (N_3087,N_1632,N_1300);
and U3088 (N_3088,N_1294,N_1675);
nand U3089 (N_3089,N_2055,N_1434);
and U3090 (N_3090,N_2058,N_1275);
xnor U3091 (N_3091,N_1528,N_2079);
nand U3092 (N_3092,N_1444,N_1357);
and U3093 (N_3093,N_2088,N_1440);
nor U3094 (N_3094,N_1806,N_1282);
and U3095 (N_3095,N_1266,N_1906);
or U3096 (N_3096,N_2359,N_1338);
nand U3097 (N_3097,N_1357,N_2386);
and U3098 (N_3098,N_1607,N_1985);
or U3099 (N_3099,N_2330,N_1894);
nand U3100 (N_3100,N_2073,N_1783);
and U3101 (N_3101,N_2141,N_1323);
or U3102 (N_3102,N_2347,N_1358);
xor U3103 (N_3103,N_1936,N_1549);
xor U3104 (N_3104,N_1645,N_1400);
xnor U3105 (N_3105,N_2247,N_2009);
nand U3106 (N_3106,N_1365,N_2010);
nand U3107 (N_3107,N_1730,N_1643);
or U3108 (N_3108,N_1792,N_2271);
or U3109 (N_3109,N_1517,N_2164);
nor U3110 (N_3110,N_2077,N_1512);
xor U3111 (N_3111,N_1715,N_2225);
or U3112 (N_3112,N_1931,N_2089);
xnor U3113 (N_3113,N_1883,N_2013);
xnor U3114 (N_3114,N_1311,N_2363);
and U3115 (N_3115,N_2326,N_1452);
and U3116 (N_3116,N_1901,N_2253);
nand U3117 (N_3117,N_1448,N_2123);
xor U3118 (N_3118,N_1833,N_1523);
or U3119 (N_3119,N_1787,N_1951);
and U3120 (N_3120,N_1270,N_1830);
xnor U3121 (N_3121,N_1934,N_1638);
and U3122 (N_3122,N_2116,N_2333);
and U3123 (N_3123,N_1739,N_2385);
xnor U3124 (N_3124,N_1458,N_1698);
nand U3125 (N_3125,N_1884,N_1369);
and U3126 (N_3126,N_1716,N_1423);
or U3127 (N_3127,N_2184,N_1621);
xor U3128 (N_3128,N_2052,N_1449);
or U3129 (N_3129,N_1516,N_1693);
and U3130 (N_3130,N_1369,N_1231);
nor U3131 (N_3131,N_1934,N_2035);
xnor U3132 (N_3132,N_1867,N_2391);
and U3133 (N_3133,N_1372,N_2175);
or U3134 (N_3134,N_2072,N_1478);
xnor U3135 (N_3135,N_1586,N_1845);
or U3136 (N_3136,N_1235,N_2005);
or U3137 (N_3137,N_2124,N_1284);
nor U3138 (N_3138,N_1435,N_2213);
xnor U3139 (N_3139,N_1812,N_1549);
nor U3140 (N_3140,N_2128,N_2335);
xor U3141 (N_3141,N_1213,N_2002);
or U3142 (N_3142,N_1459,N_1862);
nand U3143 (N_3143,N_1644,N_1268);
nand U3144 (N_3144,N_1293,N_2163);
and U3145 (N_3145,N_1725,N_2224);
xnor U3146 (N_3146,N_2195,N_1719);
nand U3147 (N_3147,N_2301,N_2025);
nor U3148 (N_3148,N_2252,N_1997);
or U3149 (N_3149,N_1534,N_1671);
and U3150 (N_3150,N_1879,N_1588);
nor U3151 (N_3151,N_1292,N_1905);
and U3152 (N_3152,N_1720,N_1570);
nor U3153 (N_3153,N_1544,N_1689);
xor U3154 (N_3154,N_1955,N_1271);
nor U3155 (N_3155,N_1852,N_1433);
nor U3156 (N_3156,N_2105,N_1810);
nor U3157 (N_3157,N_1351,N_1307);
nand U3158 (N_3158,N_2256,N_1218);
nand U3159 (N_3159,N_1891,N_1526);
nand U3160 (N_3160,N_2133,N_1684);
xor U3161 (N_3161,N_1836,N_1438);
xor U3162 (N_3162,N_2065,N_1653);
xnor U3163 (N_3163,N_1418,N_1579);
nor U3164 (N_3164,N_2253,N_1978);
xnor U3165 (N_3165,N_2094,N_1742);
or U3166 (N_3166,N_1896,N_1217);
nor U3167 (N_3167,N_1203,N_1647);
or U3168 (N_3168,N_2110,N_1250);
xor U3169 (N_3169,N_1236,N_1999);
or U3170 (N_3170,N_2049,N_1864);
and U3171 (N_3171,N_1665,N_2074);
and U3172 (N_3172,N_1404,N_2175);
or U3173 (N_3173,N_2198,N_2190);
xnor U3174 (N_3174,N_1503,N_1876);
or U3175 (N_3175,N_1405,N_2292);
nand U3176 (N_3176,N_2284,N_1663);
nand U3177 (N_3177,N_1793,N_1837);
xor U3178 (N_3178,N_1877,N_1938);
or U3179 (N_3179,N_2037,N_1495);
xor U3180 (N_3180,N_2392,N_2246);
xnor U3181 (N_3181,N_1662,N_2385);
nor U3182 (N_3182,N_1332,N_2105);
or U3183 (N_3183,N_1458,N_2342);
or U3184 (N_3184,N_1426,N_1291);
nand U3185 (N_3185,N_1832,N_1706);
and U3186 (N_3186,N_1553,N_2076);
xor U3187 (N_3187,N_1399,N_2238);
and U3188 (N_3188,N_2135,N_1620);
nor U3189 (N_3189,N_2276,N_2328);
or U3190 (N_3190,N_1920,N_1707);
and U3191 (N_3191,N_2158,N_1949);
nand U3192 (N_3192,N_1288,N_2256);
or U3193 (N_3193,N_2216,N_1739);
nand U3194 (N_3194,N_1670,N_1734);
or U3195 (N_3195,N_2165,N_1968);
nand U3196 (N_3196,N_1823,N_1889);
and U3197 (N_3197,N_1717,N_1770);
nand U3198 (N_3198,N_1855,N_2178);
xnor U3199 (N_3199,N_2314,N_1879);
xnor U3200 (N_3200,N_1889,N_1303);
or U3201 (N_3201,N_1216,N_1494);
and U3202 (N_3202,N_1378,N_1530);
or U3203 (N_3203,N_2037,N_2116);
or U3204 (N_3204,N_1255,N_1247);
and U3205 (N_3205,N_1872,N_1815);
xnor U3206 (N_3206,N_1471,N_1523);
xor U3207 (N_3207,N_1272,N_1956);
xnor U3208 (N_3208,N_1775,N_2091);
xor U3209 (N_3209,N_1800,N_1710);
nor U3210 (N_3210,N_1856,N_2137);
and U3211 (N_3211,N_2302,N_2328);
nand U3212 (N_3212,N_2125,N_2173);
xnor U3213 (N_3213,N_1636,N_1876);
and U3214 (N_3214,N_1576,N_1561);
nand U3215 (N_3215,N_1491,N_2295);
nor U3216 (N_3216,N_1749,N_2167);
nor U3217 (N_3217,N_1425,N_1623);
or U3218 (N_3218,N_1737,N_2065);
and U3219 (N_3219,N_1787,N_1794);
xnor U3220 (N_3220,N_2207,N_1422);
or U3221 (N_3221,N_1466,N_2301);
xnor U3222 (N_3222,N_2386,N_2377);
and U3223 (N_3223,N_1795,N_2237);
nand U3224 (N_3224,N_1406,N_1231);
nand U3225 (N_3225,N_2019,N_1407);
xnor U3226 (N_3226,N_1596,N_2256);
or U3227 (N_3227,N_1665,N_1581);
nor U3228 (N_3228,N_2290,N_2189);
nor U3229 (N_3229,N_1813,N_1321);
xnor U3230 (N_3230,N_1531,N_1310);
nor U3231 (N_3231,N_2000,N_2301);
nand U3232 (N_3232,N_1568,N_1763);
xor U3233 (N_3233,N_1788,N_1674);
nand U3234 (N_3234,N_2284,N_2366);
and U3235 (N_3235,N_1867,N_1563);
or U3236 (N_3236,N_2273,N_1220);
or U3237 (N_3237,N_1634,N_1298);
xor U3238 (N_3238,N_1839,N_1812);
or U3239 (N_3239,N_1761,N_2290);
nand U3240 (N_3240,N_2253,N_2058);
nand U3241 (N_3241,N_2050,N_1478);
and U3242 (N_3242,N_1964,N_1714);
nand U3243 (N_3243,N_1665,N_2375);
or U3244 (N_3244,N_2006,N_1389);
and U3245 (N_3245,N_2002,N_1202);
and U3246 (N_3246,N_1376,N_2216);
nor U3247 (N_3247,N_1928,N_1361);
or U3248 (N_3248,N_1554,N_2378);
nand U3249 (N_3249,N_1876,N_2009);
and U3250 (N_3250,N_1295,N_1633);
and U3251 (N_3251,N_2224,N_1326);
xor U3252 (N_3252,N_2005,N_2357);
xnor U3253 (N_3253,N_1275,N_1823);
nand U3254 (N_3254,N_1743,N_1394);
or U3255 (N_3255,N_1866,N_1405);
or U3256 (N_3256,N_1492,N_1814);
xnor U3257 (N_3257,N_1263,N_1840);
nor U3258 (N_3258,N_1703,N_2399);
xor U3259 (N_3259,N_1326,N_1615);
nor U3260 (N_3260,N_1517,N_1466);
nor U3261 (N_3261,N_2216,N_1325);
nand U3262 (N_3262,N_1346,N_1467);
or U3263 (N_3263,N_2176,N_1351);
xor U3264 (N_3264,N_1532,N_1774);
and U3265 (N_3265,N_1289,N_1582);
and U3266 (N_3266,N_1512,N_2184);
or U3267 (N_3267,N_1956,N_1571);
or U3268 (N_3268,N_1860,N_1409);
and U3269 (N_3269,N_1945,N_1515);
and U3270 (N_3270,N_2320,N_1277);
nand U3271 (N_3271,N_1553,N_2101);
xor U3272 (N_3272,N_2017,N_1526);
nand U3273 (N_3273,N_2232,N_2091);
or U3274 (N_3274,N_1494,N_1725);
xnor U3275 (N_3275,N_2344,N_1479);
or U3276 (N_3276,N_2082,N_2183);
and U3277 (N_3277,N_1414,N_1280);
or U3278 (N_3278,N_1372,N_1639);
xor U3279 (N_3279,N_1342,N_1874);
nor U3280 (N_3280,N_2221,N_2234);
nor U3281 (N_3281,N_2157,N_1349);
xnor U3282 (N_3282,N_2331,N_1266);
nor U3283 (N_3283,N_2088,N_2272);
nand U3284 (N_3284,N_2115,N_2313);
nand U3285 (N_3285,N_1692,N_1753);
xnor U3286 (N_3286,N_1228,N_1972);
and U3287 (N_3287,N_1671,N_1552);
xor U3288 (N_3288,N_1273,N_1422);
or U3289 (N_3289,N_1633,N_2207);
nor U3290 (N_3290,N_2111,N_1967);
xnor U3291 (N_3291,N_2271,N_2003);
nand U3292 (N_3292,N_2052,N_1667);
or U3293 (N_3293,N_1673,N_1636);
nand U3294 (N_3294,N_2196,N_2002);
nand U3295 (N_3295,N_2373,N_2015);
nand U3296 (N_3296,N_1921,N_1660);
nand U3297 (N_3297,N_1796,N_1570);
nor U3298 (N_3298,N_2284,N_1657);
or U3299 (N_3299,N_1828,N_2292);
and U3300 (N_3300,N_1458,N_2037);
xnor U3301 (N_3301,N_2392,N_1811);
nand U3302 (N_3302,N_1968,N_1905);
nand U3303 (N_3303,N_1506,N_1386);
nand U3304 (N_3304,N_2386,N_1286);
nor U3305 (N_3305,N_1986,N_1438);
nand U3306 (N_3306,N_1289,N_2166);
xor U3307 (N_3307,N_1519,N_1678);
xor U3308 (N_3308,N_1421,N_1986);
and U3309 (N_3309,N_1502,N_1348);
nand U3310 (N_3310,N_2219,N_1685);
xnor U3311 (N_3311,N_1463,N_1966);
and U3312 (N_3312,N_1841,N_2371);
nand U3313 (N_3313,N_2214,N_2177);
and U3314 (N_3314,N_1704,N_1806);
or U3315 (N_3315,N_1489,N_1217);
or U3316 (N_3316,N_1607,N_1406);
xnor U3317 (N_3317,N_1679,N_1969);
xor U3318 (N_3318,N_2286,N_1715);
and U3319 (N_3319,N_1419,N_1460);
and U3320 (N_3320,N_1359,N_1207);
and U3321 (N_3321,N_1694,N_2378);
nor U3322 (N_3322,N_2346,N_1427);
and U3323 (N_3323,N_1919,N_2244);
xor U3324 (N_3324,N_2202,N_2213);
and U3325 (N_3325,N_1860,N_2226);
xnor U3326 (N_3326,N_1663,N_1654);
and U3327 (N_3327,N_2336,N_2182);
or U3328 (N_3328,N_1705,N_1609);
xnor U3329 (N_3329,N_1558,N_1623);
or U3330 (N_3330,N_2157,N_1628);
and U3331 (N_3331,N_1989,N_2195);
or U3332 (N_3332,N_2183,N_1958);
or U3333 (N_3333,N_1524,N_2141);
nand U3334 (N_3334,N_1256,N_2298);
xnor U3335 (N_3335,N_2316,N_2314);
or U3336 (N_3336,N_2002,N_2121);
nor U3337 (N_3337,N_1467,N_1516);
or U3338 (N_3338,N_1648,N_1412);
nor U3339 (N_3339,N_1623,N_1957);
and U3340 (N_3340,N_1981,N_1913);
nor U3341 (N_3341,N_1474,N_2396);
and U3342 (N_3342,N_1802,N_1291);
nor U3343 (N_3343,N_1278,N_1477);
or U3344 (N_3344,N_2095,N_2399);
and U3345 (N_3345,N_1602,N_1475);
nand U3346 (N_3346,N_2056,N_2273);
and U3347 (N_3347,N_1843,N_2321);
nand U3348 (N_3348,N_1631,N_1451);
or U3349 (N_3349,N_1927,N_1891);
nand U3350 (N_3350,N_2232,N_2394);
xnor U3351 (N_3351,N_2334,N_2356);
nand U3352 (N_3352,N_1983,N_1939);
or U3353 (N_3353,N_1509,N_2146);
nand U3354 (N_3354,N_2255,N_2081);
and U3355 (N_3355,N_1679,N_2285);
and U3356 (N_3356,N_1358,N_1313);
xor U3357 (N_3357,N_1850,N_2284);
or U3358 (N_3358,N_2062,N_1825);
nor U3359 (N_3359,N_1549,N_2172);
nand U3360 (N_3360,N_2277,N_1788);
and U3361 (N_3361,N_1330,N_1650);
and U3362 (N_3362,N_1335,N_1325);
or U3363 (N_3363,N_1581,N_1235);
and U3364 (N_3364,N_1527,N_1680);
nand U3365 (N_3365,N_2009,N_2106);
nand U3366 (N_3366,N_1441,N_2040);
nand U3367 (N_3367,N_1615,N_1750);
or U3368 (N_3368,N_1438,N_1253);
or U3369 (N_3369,N_1310,N_2126);
or U3370 (N_3370,N_2000,N_1805);
xnor U3371 (N_3371,N_2381,N_1512);
xor U3372 (N_3372,N_2038,N_1732);
and U3373 (N_3373,N_1910,N_1291);
or U3374 (N_3374,N_1277,N_2092);
and U3375 (N_3375,N_1352,N_2053);
or U3376 (N_3376,N_1612,N_1229);
nand U3377 (N_3377,N_1905,N_2287);
and U3378 (N_3378,N_1428,N_1496);
nand U3379 (N_3379,N_2319,N_1585);
or U3380 (N_3380,N_1247,N_2371);
xor U3381 (N_3381,N_2015,N_1369);
and U3382 (N_3382,N_1306,N_1858);
and U3383 (N_3383,N_1943,N_1284);
and U3384 (N_3384,N_1210,N_2020);
nand U3385 (N_3385,N_1559,N_1871);
nor U3386 (N_3386,N_1760,N_1880);
or U3387 (N_3387,N_2318,N_2310);
xnor U3388 (N_3388,N_2295,N_1762);
nor U3389 (N_3389,N_1344,N_1410);
nand U3390 (N_3390,N_1555,N_1396);
and U3391 (N_3391,N_2162,N_1706);
nand U3392 (N_3392,N_2069,N_2145);
nor U3393 (N_3393,N_2072,N_1488);
xnor U3394 (N_3394,N_1273,N_2069);
xor U3395 (N_3395,N_1213,N_1482);
and U3396 (N_3396,N_2292,N_1820);
or U3397 (N_3397,N_1417,N_1368);
nand U3398 (N_3398,N_2159,N_1300);
xnor U3399 (N_3399,N_1843,N_1664);
xnor U3400 (N_3400,N_2287,N_1911);
nand U3401 (N_3401,N_1269,N_1831);
xor U3402 (N_3402,N_1817,N_1941);
and U3403 (N_3403,N_1475,N_1587);
and U3404 (N_3404,N_1791,N_1940);
or U3405 (N_3405,N_1796,N_1660);
xor U3406 (N_3406,N_1206,N_1929);
nor U3407 (N_3407,N_1344,N_2087);
nor U3408 (N_3408,N_1382,N_1554);
and U3409 (N_3409,N_1298,N_1506);
xnor U3410 (N_3410,N_1557,N_1594);
nor U3411 (N_3411,N_1414,N_2266);
or U3412 (N_3412,N_2174,N_2371);
xor U3413 (N_3413,N_1768,N_2369);
nor U3414 (N_3414,N_1959,N_1970);
nand U3415 (N_3415,N_1459,N_2262);
xor U3416 (N_3416,N_1314,N_1561);
or U3417 (N_3417,N_1762,N_1944);
nand U3418 (N_3418,N_2133,N_1925);
and U3419 (N_3419,N_1713,N_2120);
nor U3420 (N_3420,N_2040,N_2172);
xor U3421 (N_3421,N_2027,N_2039);
and U3422 (N_3422,N_1788,N_1243);
and U3423 (N_3423,N_1808,N_1434);
and U3424 (N_3424,N_1699,N_1924);
and U3425 (N_3425,N_1733,N_2320);
and U3426 (N_3426,N_1448,N_2258);
nor U3427 (N_3427,N_1873,N_1594);
and U3428 (N_3428,N_1633,N_2085);
nand U3429 (N_3429,N_1889,N_2139);
and U3430 (N_3430,N_2026,N_1327);
or U3431 (N_3431,N_1693,N_1629);
nand U3432 (N_3432,N_1870,N_2238);
or U3433 (N_3433,N_1875,N_1726);
or U3434 (N_3434,N_2362,N_1255);
xor U3435 (N_3435,N_2124,N_1326);
or U3436 (N_3436,N_2132,N_1920);
xor U3437 (N_3437,N_2380,N_2173);
xnor U3438 (N_3438,N_1360,N_2262);
xnor U3439 (N_3439,N_1326,N_1743);
xnor U3440 (N_3440,N_1347,N_1995);
xnor U3441 (N_3441,N_1947,N_2217);
and U3442 (N_3442,N_2094,N_2228);
xnor U3443 (N_3443,N_1228,N_1248);
nand U3444 (N_3444,N_2058,N_1962);
and U3445 (N_3445,N_1362,N_2355);
nand U3446 (N_3446,N_1594,N_1294);
nor U3447 (N_3447,N_1409,N_1459);
nand U3448 (N_3448,N_1562,N_2345);
nand U3449 (N_3449,N_1442,N_2226);
nand U3450 (N_3450,N_2074,N_1368);
nand U3451 (N_3451,N_1723,N_2316);
and U3452 (N_3452,N_2153,N_1972);
xnor U3453 (N_3453,N_2268,N_2043);
nor U3454 (N_3454,N_2206,N_1271);
xor U3455 (N_3455,N_1715,N_1636);
or U3456 (N_3456,N_1864,N_1979);
or U3457 (N_3457,N_1760,N_2059);
and U3458 (N_3458,N_1426,N_1809);
nand U3459 (N_3459,N_2355,N_1657);
xor U3460 (N_3460,N_1853,N_1396);
xnor U3461 (N_3461,N_1265,N_1343);
xor U3462 (N_3462,N_2298,N_1516);
and U3463 (N_3463,N_2030,N_2178);
nor U3464 (N_3464,N_2074,N_1688);
nor U3465 (N_3465,N_2125,N_2269);
and U3466 (N_3466,N_1201,N_1241);
xnor U3467 (N_3467,N_1257,N_2213);
and U3468 (N_3468,N_2087,N_1531);
nor U3469 (N_3469,N_1295,N_1911);
nand U3470 (N_3470,N_1410,N_1770);
and U3471 (N_3471,N_1821,N_1418);
or U3472 (N_3472,N_1685,N_1396);
and U3473 (N_3473,N_1485,N_1809);
and U3474 (N_3474,N_1280,N_1737);
xor U3475 (N_3475,N_1803,N_1620);
xnor U3476 (N_3476,N_1928,N_2340);
nor U3477 (N_3477,N_2043,N_2172);
xor U3478 (N_3478,N_1858,N_2221);
or U3479 (N_3479,N_2011,N_2076);
or U3480 (N_3480,N_1966,N_1976);
and U3481 (N_3481,N_1684,N_1361);
and U3482 (N_3482,N_1201,N_2345);
nand U3483 (N_3483,N_1655,N_1646);
nor U3484 (N_3484,N_1250,N_1756);
nand U3485 (N_3485,N_1871,N_1228);
nand U3486 (N_3486,N_1783,N_1510);
and U3487 (N_3487,N_1620,N_2089);
nand U3488 (N_3488,N_1485,N_1939);
nor U3489 (N_3489,N_1753,N_2213);
or U3490 (N_3490,N_2359,N_1256);
nor U3491 (N_3491,N_2273,N_2331);
nor U3492 (N_3492,N_1220,N_1240);
nand U3493 (N_3493,N_2337,N_1633);
nor U3494 (N_3494,N_1218,N_2361);
nand U3495 (N_3495,N_2221,N_2171);
xnor U3496 (N_3496,N_2003,N_1796);
and U3497 (N_3497,N_1803,N_1887);
and U3498 (N_3498,N_1254,N_1249);
or U3499 (N_3499,N_2068,N_2273);
xnor U3500 (N_3500,N_1946,N_2039);
xor U3501 (N_3501,N_1834,N_1889);
xor U3502 (N_3502,N_2238,N_2240);
nand U3503 (N_3503,N_1811,N_1973);
xor U3504 (N_3504,N_1399,N_2370);
nand U3505 (N_3505,N_1472,N_1299);
nand U3506 (N_3506,N_2068,N_2093);
xor U3507 (N_3507,N_1241,N_1408);
nor U3508 (N_3508,N_1662,N_2211);
and U3509 (N_3509,N_1352,N_2061);
nand U3510 (N_3510,N_2189,N_1823);
or U3511 (N_3511,N_1404,N_2026);
or U3512 (N_3512,N_2192,N_1978);
nand U3513 (N_3513,N_1953,N_1974);
xnor U3514 (N_3514,N_1624,N_1465);
and U3515 (N_3515,N_2145,N_1255);
and U3516 (N_3516,N_1413,N_2086);
xor U3517 (N_3517,N_1531,N_1598);
xor U3518 (N_3518,N_1792,N_2348);
and U3519 (N_3519,N_1303,N_1798);
nor U3520 (N_3520,N_1700,N_2005);
nand U3521 (N_3521,N_1586,N_1411);
or U3522 (N_3522,N_2039,N_1951);
nor U3523 (N_3523,N_1355,N_1931);
nor U3524 (N_3524,N_1838,N_1910);
xnor U3525 (N_3525,N_1329,N_1996);
nor U3526 (N_3526,N_2107,N_1522);
nand U3527 (N_3527,N_2093,N_2064);
nor U3528 (N_3528,N_1224,N_1799);
and U3529 (N_3529,N_2276,N_1744);
and U3530 (N_3530,N_1597,N_1203);
xor U3531 (N_3531,N_1985,N_1599);
nor U3532 (N_3532,N_2022,N_2177);
and U3533 (N_3533,N_1620,N_2228);
or U3534 (N_3534,N_1703,N_1580);
nand U3535 (N_3535,N_2262,N_1535);
nor U3536 (N_3536,N_2002,N_2108);
and U3537 (N_3537,N_1609,N_1672);
or U3538 (N_3538,N_1638,N_1572);
xnor U3539 (N_3539,N_1918,N_1737);
xnor U3540 (N_3540,N_1907,N_2113);
and U3541 (N_3541,N_1998,N_2004);
nor U3542 (N_3542,N_1641,N_2293);
xnor U3543 (N_3543,N_1601,N_2121);
nor U3544 (N_3544,N_1293,N_1549);
or U3545 (N_3545,N_1937,N_1217);
and U3546 (N_3546,N_2108,N_1333);
nand U3547 (N_3547,N_1432,N_1579);
or U3548 (N_3548,N_1673,N_1736);
or U3549 (N_3549,N_1358,N_1461);
and U3550 (N_3550,N_1378,N_1279);
and U3551 (N_3551,N_1431,N_2341);
nand U3552 (N_3552,N_1910,N_1766);
or U3553 (N_3553,N_1252,N_1429);
nor U3554 (N_3554,N_2198,N_1266);
or U3555 (N_3555,N_1320,N_1344);
and U3556 (N_3556,N_2130,N_1994);
or U3557 (N_3557,N_1416,N_2035);
xor U3558 (N_3558,N_2271,N_2010);
or U3559 (N_3559,N_2085,N_1660);
or U3560 (N_3560,N_1400,N_2094);
or U3561 (N_3561,N_1467,N_2208);
and U3562 (N_3562,N_1413,N_2095);
xnor U3563 (N_3563,N_1675,N_2313);
nand U3564 (N_3564,N_1924,N_1572);
nand U3565 (N_3565,N_1872,N_2211);
nor U3566 (N_3566,N_1882,N_1884);
nand U3567 (N_3567,N_1688,N_2128);
or U3568 (N_3568,N_1798,N_1525);
nand U3569 (N_3569,N_2212,N_1743);
nor U3570 (N_3570,N_1357,N_1943);
xnor U3571 (N_3571,N_1832,N_2377);
xor U3572 (N_3572,N_2080,N_1924);
and U3573 (N_3573,N_1849,N_2215);
nor U3574 (N_3574,N_2116,N_2370);
nand U3575 (N_3575,N_1665,N_1984);
nand U3576 (N_3576,N_1843,N_2078);
nand U3577 (N_3577,N_1269,N_1828);
nor U3578 (N_3578,N_2380,N_1599);
and U3579 (N_3579,N_1468,N_1959);
or U3580 (N_3580,N_1850,N_1358);
nor U3581 (N_3581,N_2266,N_2159);
xnor U3582 (N_3582,N_2077,N_2133);
xnor U3583 (N_3583,N_1435,N_1785);
xnor U3584 (N_3584,N_1491,N_1770);
and U3585 (N_3585,N_1832,N_1513);
nor U3586 (N_3586,N_2196,N_1757);
xnor U3587 (N_3587,N_1692,N_1747);
xor U3588 (N_3588,N_1868,N_1756);
xor U3589 (N_3589,N_1475,N_1346);
and U3590 (N_3590,N_1865,N_1569);
nand U3591 (N_3591,N_1592,N_2285);
nor U3592 (N_3592,N_2005,N_1853);
nor U3593 (N_3593,N_1509,N_1446);
or U3594 (N_3594,N_1303,N_1988);
nand U3595 (N_3595,N_1280,N_1764);
or U3596 (N_3596,N_1692,N_1592);
nor U3597 (N_3597,N_1390,N_1384);
nand U3598 (N_3598,N_1879,N_2184);
and U3599 (N_3599,N_1258,N_2017);
or U3600 (N_3600,N_2527,N_3230);
and U3601 (N_3601,N_3388,N_3091);
nand U3602 (N_3602,N_3469,N_3081);
xor U3603 (N_3603,N_2532,N_3251);
nand U3604 (N_3604,N_2590,N_3221);
nand U3605 (N_3605,N_3396,N_3033);
nand U3606 (N_3606,N_2434,N_3143);
xnor U3607 (N_3607,N_3341,N_2539);
and U3608 (N_3608,N_2880,N_2691);
nand U3609 (N_3609,N_2760,N_3038);
xnor U3610 (N_3610,N_2877,N_2730);
nor U3611 (N_3611,N_3229,N_3591);
xor U3612 (N_3612,N_2946,N_3334);
or U3613 (N_3613,N_3022,N_2411);
nor U3614 (N_3614,N_2862,N_3294);
nand U3615 (N_3615,N_3574,N_3529);
xor U3616 (N_3616,N_3531,N_3084);
or U3617 (N_3617,N_3534,N_2910);
nand U3618 (N_3618,N_2766,N_3519);
xnor U3619 (N_3619,N_3487,N_3235);
nand U3620 (N_3620,N_2895,N_2911);
or U3621 (N_3621,N_2899,N_2721);
nor U3622 (N_3622,N_2927,N_3359);
or U3623 (N_3623,N_2738,N_3323);
nand U3624 (N_3624,N_2933,N_2792);
nand U3625 (N_3625,N_2664,N_3111);
nor U3626 (N_3626,N_3215,N_2837);
and U3627 (N_3627,N_3029,N_3062);
or U3628 (N_3628,N_3048,N_3035);
xnor U3629 (N_3629,N_2656,N_3288);
xor U3630 (N_3630,N_3289,N_3416);
or U3631 (N_3631,N_3045,N_2676);
xnor U3632 (N_3632,N_2867,N_2740);
or U3633 (N_3633,N_2875,N_3583);
nand U3634 (N_3634,N_2629,N_3197);
or U3635 (N_3635,N_3172,N_2553);
and U3636 (N_3636,N_2719,N_3060);
and U3637 (N_3637,N_2701,N_3043);
and U3638 (N_3638,N_2936,N_2608);
nor U3639 (N_3639,N_2761,N_2972);
and U3640 (N_3640,N_3198,N_2441);
and U3641 (N_3641,N_2923,N_2796);
nor U3642 (N_3642,N_3053,N_2826);
nor U3643 (N_3643,N_2457,N_3509);
and U3644 (N_3644,N_2703,N_2660);
and U3645 (N_3645,N_2401,N_2913);
nand U3646 (N_3646,N_3112,N_3241);
nor U3647 (N_3647,N_3319,N_3152);
xor U3648 (N_3648,N_3086,N_3131);
nor U3649 (N_3649,N_3597,N_2589);
or U3650 (N_3650,N_2777,N_2617);
nor U3651 (N_3651,N_3077,N_2484);
xor U3652 (N_3652,N_3391,N_3103);
nand U3653 (N_3653,N_2483,N_3495);
or U3654 (N_3654,N_2635,N_2773);
nand U3655 (N_3655,N_2602,N_2770);
and U3656 (N_3656,N_3484,N_2555);
or U3657 (N_3657,N_2799,N_2898);
or U3658 (N_3658,N_3122,N_2502);
xor U3659 (N_3659,N_2426,N_2612);
nor U3660 (N_3660,N_2958,N_2450);
and U3661 (N_3661,N_3355,N_2797);
and U3662 (N_3662,N_3194,N_2978);
or U3663 (N_3663,N_3080,N_2726);
nand U3664 (N_3664,N_2813,N_3119);
xor U3665 (N_3665,N_2588,N_3299);
and U3666 (N_3666,N_3558,N_3508);
nand U3667 (N_3667,N_3559,N_2666);
nand U3668 (N_3668,N_3343,N_3339);
xnor U3669 (N_3669,N_2914,N_2506);
nand U3670 (N_3670,N_3503,N_3256);
xor U3671 (N_3671,N_3335,N_3114);
xor U3672 (N_3672,N_2607,N_3375);
nor U3673 (N_3673,N_3521,N_3490);
xor U3674 (N_3674,N_3063,N_3496);
or U3675 (N_3675,N_2793,N_3201);
xor U3676 (N_3676,N_2685,N_3144);
or U3677 (N_3677,N_3020,N_2771);
nand U3678 (N_3678,N_2474,N_2892);
xor U3679 (N_3679,N_3464,N_2592);
nor U3680 (N_3680,N_3378,N_2560);
or U3681 (N_3681,N_3065,N_3403);
xor U3682 (N_3682,N_2470,N_3439);
xnor U3683 (N_3683,N_2584,N_2780);
nor U3684 (N_3684,N_2807,N_3097);
nand U3685 (N_3685,N_3382,N_3115);
and U3686 (N_3686,N_3417,N_3088);
nor U3687 (N_3687,N_3457,N_2767);
nor U3688 (N_3688,N_2732,N_3407);
and U3689 (N_3689,N_3567,N_2653);
and U3690 (N_3690,N_2815,N_2670);
nand U3691 (N_3691,N_2987,N_2804);
xor U3692 (N_3692,N_2577,N_2782);
nor U3693 (N_3693,N_2501,N_3171);
and U3694 (N_3694,N_2728,N_3433);
nor U3695 (N_3695,N_2665,N_2999);
and U3696 (N_3696,N_3147,N_2843);
or U3697 (N_3697,N_3575,N_2684);
nor U3698 (N_3698,N_3493,N_3419);
xor U3699 (N_3699,N_3264,N_2624);
xor U3700 (N_3700,N_3428,N_2802);
or U3701 (N_3701,N_2884,N_2791);
nand U3702 (N_3702,N_3465,N_2749);
nand U3703 (N_3703,N_3116,N_3523);
or U3704 (N_3704,N_3373,N_3432);
or U3705 (N_3705,N_3308,N_2601);
nand U3706 (N_3706,N_2836,N_2647);
or U3707 (N_3707,N_2998,N_2768);
or U3708 (N_3708,N_2979,N_2654);
xor U3709 (N_3709,N_2774,N_2904);
xor U3710 (N_3710,N_3213,N_3217);
xnor U3711 (N_3711,N_2544,N_3340);
nand U3712 (N_3712,N_2471,N_2615);
nor U3713 (N_3713,N_3546,N_2631);
xor U3714 (N_3714,N_3214,N_3446);
nor U3715 (N_3715,N_2893,N_2430);
nand U3716 (N_3716,N_2948,N_3431);
nor U3717 (N_3717,N_2757,N_3581);
nand U3718 (N_3718,N_3379,N_3386);
xor U3719 (N_3719,N_3442,N_3422);
and U3720 (N_3720,N_3021,N_2717);
and U3721 (N_3721,N_2762,N_3268);
nor U3722 (N_3722,N_2954,N_2578);
xor U3723 (N_3723,N_2551,N_3309);
or U3724 (N_3724,N_2498,N_3402);
nor U3725 (N_3725,N_2462,N_3146);
xor U3726 (N_3726,N_3526,N_2934);
or U3727 (N_3727,N_2447,N_3459);
nand U3728 (N_3728,N_3209,N_2897);
nand U3729 (N_3729,N_3205,N_3480);
nor U3730 (N_3730,N_2481,N_3538);
nand U3731 (N_3731,N_2627,N_3248);
and U3732 (N_3732,N_2412,N_3301);
or U3733 (N_3733,N_3117,N_2810);
xor U3734 (N_3734,N_3224,N_2517);
and U3735 (N_3735,N_2930,N_3506);
xnor U3736 (N_3736,N_3188,N_2870);
nor U3737 (N_3737,N_2865,N_2745);
xor U3738 (N_3738,N_2781,N_3515);
or U3739 (N_3739,N_3360,N_3192);
or U3740 (N_3740,N_3032,N_3260);
xnor U3741 (N_3741,N_3313,N_2931);
and U3742 (N_3742,N_3349,N_3336);
nor U3743 (N_3743,N_2682,N_2747);
nand U3744 (N_3744,N_3276,N_2929);
and U3745 (N_3745,N_2821,N_2764);
nor U3746 (N_3746,N_3039,N_3399);
and U3747 (N_3747,N_3453,N_3505);
nor U3748 (N_3748,N_2418,N_3489);
and U3749 (N_3749,N_2603,N_2846);
or U3750 (N_3750,N_3377,N_3383);
or U3751 (N_3751,N_2473,N_3070);
nand U3752 (N_3752,N_2431,N_2966);
nand U3753 (N_3753,N_2983,N_2794);
nand U3754 (N_3754,N_2622,N_3105);
or U3755 (N_3755,N_2822,N_2960);
and U3756 (N_3756,N_2504,N_3000);
nor U3757 (N_3757,N_2640,N_2596);
xor U3758 (N_3758,N_2487,N_3332);
or U3759 (N_3759,N_3311,N_3278);
and U3760 (N_3760,N_3579,N_3361);
nand U3761 (N_3761,N_2633,N_2790);
nor U3762 (N_3762,N_2550,N_3404);
xor U3763 (N_3763,N_2806,N_3145);
and U3764 (N_3764,N_3456,N_2452);
nand U3765 (N_3765,N_3445,N_3321);
nand U3766 (N_3766,N_2708,N_2533);
or U3767 (N_3767,N_3389,N_2569);
nor U3768 (N_3768,N_2787,N_3189);
or U3769 (N_3769,N_3483,N_2723);
nand U3770 (N_3770,N_3364,N_2872);
nand U3771 (N_3771,N_2585,N_2926);
nand U3772 (N_3772,N_2632,N_3303);
nand U3773 (N_3773,N_2696,N_2641);
or U3774 (N_3774,N_3199,N_3369);
nor U3775 (N_3775,N_2439,N_3544);
or U3776 (N_3776,N_2969,N_2456);
nand U3777 (N_3777,N_3387,N_2976);
nor U3778 (N_3778,N_3418,N_2964);
xor U3779 (N_3779,N_2658,N_2642);
nor U3780 (N_3780,N_2557,N_2683);
nand U3781 (N_3781,N_2851,N_3061);
xor U3782 (N_3782,N_3517,N_2536);
xnor U3783 (N_3783,N_3239,N_3392);
xor U3784 (N_3784,N_3525,N_3316);
or U3785 (N_3785,N_3073,N_3025);
or U3786 (N_3786,N_3331,N_2834);
xor U3787 (N_3787,N_3592,N_3076);
nand U3788 (N_3788,N_2838,N_3223);
nand U3789 (N_3789,N_2988,N_3176);
nand U3790 (N_3790,N_3167,N_2814);
xor U3791 (N_3791,N_2494,N_2572);
xor U3792 (N_3792,N_3085,N_3121);
nand U3793 (N_3793,N_3002,N_2547);
nor U3794 (N_3794,N_3072,N_3202);
nand U3795 (N_3795,N_3552,N_2419);
nand U3796 (N_3796,N_3139,N_3220);
or U3797 (N_3797,N_2522,N_2621);
and U3798 (N_3798,N_2800,N_2742);
or U3799 (N_3799,N_3587,N_2945);
or U3800 (N_3800,N_2811,N_2543);
nor U3801 (N_3801,N_3380,N_2619);
and U3802 (N_3802,N_2702,N_2485);
xor U3803 (N_3803,N_3598,N_3012);
and U3804 (N_3804,N_3550,N_2965);
and U3805 (N_3805,N_2967,N_3155);
nand U3806 (N_3806,N_3140,N_3173);
nor U3807 (N_3807,N_3051,N_3082);
nand U3808 (N_3808,N_2659,N_2463);
or U3809 (N_3809,N_3129,N_2570);
nor U3810 (N_3810,N_3158,N_3018);
and U3811 (N_3811,N_3008,N_2499);
or U3812 (N_3812,N_3153,N_3227);
nand U3813 (N_3813,N_2906,N_2446);
xnor U3814 (N_3814,N_2783,N_3047);
nand U3815 (N_3815,N_2962,N_3367);
xnor U3816 (N_3816,N_2680,N_2593);
nor U3817 (N_3817,N_2679,N_2460);
xnor U3818 (N_3818,N_2743,N_3074);
and U3819 (N_3819,N_2751,N_2818);
nor U3820 (N_3820,N_3485,N_2488);
xnor U3821 (N_3821,N_3482,N_3259);
nor U3822 (N_3822,N_3046,N_2510);
nand U3823 (N_3823,N_3599,N_3249);
or U3824 (N_3824,N_3518,N_3222);
and U3825 (N_3825,N_3477,N_2516);
nand U3826 (N_3826,N_2402,N_3580);
nand U3827 (N_3827,N_2748,N_3430);
nor U3828 (N_3828,N_2545,N_3555);
xor U3829 (N_3829,N_3578,N_2912);
or U3830 (N_3830,N_2706,N_2848);
nor U3831 (N_3831,N_3543,N_3098);
nand U3832 (N_3832,N_2478,N_3150);
nand U3833 (N_3833,N_3514,N_3400);
nand U3834 (N_3834,N_2531,N_3540);
or U3835 (N_3835,N_2772,N_3314);
nand U3836 (N_3836,N_3193,N_3004);
nand U3837 (N_3837,N_3411,N_2951);
and U3838 (N_3838,N_2508,N_2663);
nand U3839 (N_3839,N_2973,N_2563);
nor U3840 (N_3840,N_2961,N_2825);
nand U3841 (N_3841,N_2404,N_2514);
or U3842 (N_3842,N_2681,N_2876);
nor U3843 (N_3843,N_3187,N_3243);
or U3844 (N_3844,N_3190,N_2630);
and U3845 (N_3845,N_3306,N_3041);
nand U3846 (N_3846,N_2405,N_3504);
nor U3847 (N_3847,N_2610,N_2817);
or U3848 (N_3848,N_3545,N_3551);
nor U3849 (N_3849,N_3476,N_2469);
nand U3850 (N_3850,N_2963,N_2921);
and U3851 (N_3851,N_3405,N_3120);
or U3852 (N_3852,N_2465,N_2943);
xor U3853 (N_3853,N_3136,N_2886);
and U3854 (N_3854,N_3437,N_2480);
and U3855 (N_3855,N_2556,N_2493);
nor U3856 (N_3856,N_3015,N_3354);
xor U3857 (N_3857,N_2538,N_2495);
nand U3858 (N_3858,N_2707,N_3110);
or U3859 (N_3859,N_2582,N_3159);
nor U3860 (N_3860,N_3013,N_3244);
nand U3861 (N_3861,N_3317,N_3582);
or U3862 (N_3862,N_3196,N_3478);
nand U3863 (N_3863,N_2724,N_2779);
xor U3864 (N_3864,N_2686,N_3246);
xor U3865 (N_3865,N_2968,N_3133);
or U3866 (N_3866,N_3195,N_3141);
and U3867 (N_3867,N_2731,N_3440);
xor U3868 (N_3868,N_2918,N_3058);
or U3869 (N_3869,N_3312,N_3100);
and U3870 (N_3870,N_2992,N_3398);
nor U3871 (N_3871,N_2537,N_2651);
nand U3872 (N_3872,N_3044,N_3204);
nand U3873 (N_3873,N_3408,N_2406);
xnor U3874 (N_3874,N_3185,N_3421);
and U3875 (N_3875,N_2753,N_2736);
or U3876 (N_3876,N_3151,N_2775);
xnor U3877 (N_3877,N_3412,N_3471);
nor U3878 (N_3878,N_3184,N_2981);
or U3879 (N_3879,N_2595,N_3560);
and U3880 (N_3880,N_3003,N_2733);
or U3881 (N_3881,N_3434,N_3287);
or U3882 (N_3882,N_3595,N_2917);
or U3883 (N_3883,N_3585,N_2700);
or U3884 (N_3884,N_3238,N_3106);
nor U3885 (N_3885,N_2885,N_2888);
nand U3886 (N_3886,N_3182,N_3553);
or U3887 (N_3887,N_3468,N_2648);
nor U3888 (N_3888,N_2626,N_3094);
nand U3889 (N_3889,N_2580,N_3109);
and U3890 (N_3890,N_3071,N_3448);
and U3891 (N_3891,N_3590,N_2662);
nor U3892 (N_3892,N_3451,N_2518);
nor U3893 (N_3893,N_3160,N_3068);
nand U3894 (N_3894,N_2859,N_3011);
xor U3895 (N_3895,N_2809,N_3102);
nor U3896 (N_3896,N_3372,N_2491);
and U3897 (N_3897,N_2715,N_2819);
or U3898 (N_3898,N_2451,N_3267);
nor U3899 (N_3899,N_2689,N_3031);
nor U3900 (N_3900,N_3090,N_2565);
or U3901 (N_3901,N_3092,N_2455);
or U3902 (N_3902,N_3232,N_3539);
or U3903 (N_3903,N_3397,N_3449);
or U3904 (N_3904,N_3385,N_3203);
and U3905 (N_3905,N_3059,N_2863);
or U3906 (N_3906,N_2986,N_3271);
nor U3907 (N_3907,N_3165,N_3528);
nand U3908 (N_3908,N_2438,N_2829);
nor U3909 (N_3909,N_2938,N_3118);
xnor U3910 (N_3910,N_3363,N_2750);
or U3911 (N_3911,N_3353,N_2554);
or U3912 (N_3912,N_3516,N_2526);
nor U3913 (N_3913,N_3272,N_2704);
and U3914 (N_3914,N_3257,N_3512);
or U3915 (N_3915,N_2823,N_3036);
nor U3916 (N_3916,N_2901,N_3329);
xor U3917 (N_3917,N_3183,N_2652);
xnor U3918 (N_3918,N_3325,N_2878);
xor U3919 (N_3919,N_3023,N_2552);
xor U3920 (N_3920,N_3123,N_2711);
nand U3921 (N_3921,N_2959,N_2645);
nor U3922 (N_3922,N_2669,N_3357);
or U3923 (N_3923,N_2869,N_3577);
and U3924 (N_3924,N_2925,N_3305);
and U3925 (N_3925,N_2932,N_3338);
nand U3926 (N_3926,N_3450,N_2840);
and U3927 (N_3927,N_2600,N_3502);
nor U3928 (N_3928,N_3064,N_2883);
xor U3929 (N_3929,N_2908,N_2515);
or U3930 (N_3930,N_3030,N_3414);
or U3931 (N_3931,N_2841,N_3371);
and U3932 (N_3932,N_3568,N_2692);
xnor U3933 (N_3933,N_2882,N_2941);
nand U3934 (N_3934,N_3328,N_2407);
and U3935 (N_3935,N_3454,N_3576);
xnor U3936 (N_3936,N_2739,N_2606);
xnor U3937 (N_3937,N_2524,N_3573);
xor U3938 (N_3938,N_3275,N_3542);
and U3939 (N_3939,N_2849,N_3548);
xnor U3940 (N_3940,N_3298,N_2693);
nor U3941 (N_3941,N_3310,N_3208);
xnor U3942 (N_3942,N_3207,N_3569);
nor U3943 (N_3943,N_3138,N_2828);
or U3944 (N_3944,N_2984,N_2905);
xnor U3945 (N_3945,N_3154,N_3127);
or U3946 (N_3946,N_3099,N_2970);
or U3947 (N_3947,N_3438,N_2646);
or U3948 (N_3948,N_2586,N_2765);
nor U3949 (N_3949,N_3566,N_2718);
and U3950 (N_3950,N_3280,N_3420);
nor U3951 (N_3951,N_3034,N_3443);
or U3952 (N_3952,N_3324,N_2778);
and U3953 (N_3953,N_2467,N_2448);
nor U3954 (N_3954,N_3107,N_3500);
and U3955 (N_3955,N_2808,N_2940);
nand U3956 (N_3956,N_3593,N_3206);
nor U3957 (N_3957,N_3010,N_3441);
and U3958 (N_3958,N_2678,N_3472);
xnor U3959 (N_3959,N_2637,N_3017);
nand U3960 (N_3960,N_2939,N_3237);
or U3961 (N_3961,N_2466,N_2920);
or U3962 (N_3962,N_3535,N_2655);
xnor U3963 (N_3963,N_2812,N_3491);
nand U3964 (N_3964,N_2564,N_2861);
and U3965 (N_3965,N_2534,N_2511);
xor U3966 (N_3966,N_3087,N_2425);
xor U3967 (N_3967,N_3586,N_2628);
or U3968 (N_3968,N_3296,N_3458);
and U3969 (N_3969,N_3473,N_3293);
and U3970 (N_3970,N_2786,N_3093);
or U3971 (N_3971,N_3390,N_3219);
xor U3972 (N_3972,N_2479,N_3350);
xnor U3973 (N_3973,N_3262,N_3588);
nand U3974 (N_3974,N_2847,N_3024);
xnor U3975 (N_3975,N_2614,N_3149);
nand U3976 (N_3976,N_3269,N_3498);
xnor U3977 (N_3977,N_3384,N_2649);
and U3978 (N_3978,N_3265,N_3424);
nor U3979 (N_3979,N_2873,N_2667);
or U3980 (N_3980,N_3242,N_2436);
or U3981 (N_3981,N_2996,N_2675);
xnor U3982 (N_3982,N_2587,N_3300);
or U3983 (N_3983,N_3320,N_2519);
and U3984 (N_3984,N_2618,N_3066);
or U3985 (N_3985,N_3089,N_2997);
xor U3986 (N_3986,N_3401,N_3596);
xnor U3987 (N_3987,N_2424,N_2744);
and U3988 (N_3988,N_2896,N_3026);
or U3989 (N_3989,N_2435,N_3137);
xnor U3990 (N_3990,N_2725,N_3212);
or U3991 (N_3991,N_3284,N_3014);
nand U3992 (N_3992,N_3104,N_3344);
nand U3993 (N_3993,N_2443,N_2900);
xor U3994 (N_3994,N_3270,N_3322);
or U3995 (N_3995,N_2427,N_2705);
nor U3996 (N_3996,N_3096,N_3253);
xor U3997 (N_3997,N_2529,N_3494);
nor U3998 (N_3998,N_3368,N_3462);
and U3999 (N_3999,N_3006,N_3436);
xor U4000 (N_4000,N_2830,N_2548);
and U4001 (N_4001,N_3163,N_2604);
and U4002 (N_4002,N_2453,N_2839);
nand U4003 (N_4003,N_3460,N_2575);
nand U4004 (N_4004,N_3162,N_3083);
or U4005 (N_4005,N_2638,N_3056);
nand U4006 (N_4006,N_2650,N_2489);
nor U4007 (N_4007,N_2852,N_2400);
xor U4008 (N_4008,N_2408,N_2525);
nor U4009 (N_4009,N_3486,N_3124);
nand U4010 (N_4010,N_2503,N_3040);
and U4011 (N_4011,N_2980,N_2422);
xor U4012 (N_4012,N_3180,N_3547);
nand U4013 (N_4013,N_3095,N_3532);
nand U4014 (N_4014,N_3170,N_2890);
or U4015 (N_4015,N_2975,N_2581);
nor U4016 (N_4016,N_2576,N_2541);
nor U4017 (N_4017,N_3524,N_3522);
and U4018 (N_4018,N_3225,N_3481);
nor U4019 (N_4019,N_3236,N_2801);
xor U4020 (N_4020,N_2428,N_3148);
and U4021 (N_4021,N_2845,N_3467);
nor U4022 (N_4022,N_2530,N_3016);
and U4023 (N_4023,N_3282,N_2421);
xnor U4024 (N_4024,N_2720,N_3435);
xor U4025 (N_4025,N_2674,N_2523);
and U4026 (N_4026,N_2623,N_2468);
and U4027 (N_4027,N_2985,N_2416);
xor U4028 (N_4028,N_2879,N_2758);
nor U4029 (N_4029,N_3274,N_3218);
or U4030 (N_4030,N_2716,N_3005);
and U4031 (N_4031,N_3429,N_3455);
and U4032 (N_4032,N_3290,N_2887);
nor U4033 (N_4033,N_3285,N_2505);
xor U4034 (N_4034,N_2928,N_2990);
or U4035 (N_4035,N_3307,N_2475);
xnor U4036 (N_4036,N_3277,N_3563);
or U4037 (N_4037,N_2472,N_2889);
and U4038 (N_4038,N_3067,N_2982);
nor U4039 (N_4039,N_2597,N_3266);
and U4040 (N_4040,N_3169,N_3174);
xnor U4041 (N_4041,N_3142,N_2866);
and U4042 (N_4042,N_3200,N_3594);
nor U4043 (N_4043,N_2727,N_2609);
and U4044 (N_4044,N_3536,N_2995);
nor U4045 (N_4045,N_2500,N_2858);
nand U4046 (N_4046,N_2476,N_3113);
nor U4047 (N_4047,N_3479,N_2417);
xor U4048 (N_4048,N_3234,N_2625);
xnor U4049 (N_4049,N_2558,N_3295);
or U4050 (N_4050,N_3181,N_2714);
nand U4051 (N_4051,N_2611,N_2513);
nand U4052 (N_4052,N_2432,N_2562);
nand U4053 (N_4053,N_2423,N_3501);
and U4054 (N_4054,N_3283,N_3463);
or U4055 (N_4055,N_3028,N_3423);
xnor U4056 (N_4056,N_3302,N_2445);
and U4057 (N_4057,N_2613,N_2713);
nor U4058 (N_4058,N_3132,N_3584);
xor U4059 (N_4059,N_3572,N_3342);
or U4060 (N_4060,N_3279,N_3250);
or U4061 (N_4061,N_2492,N_2694);
or U4062 (N_4062,N_3019,N_2850);
xor U4063 (N_4063,N_3315,N_3079);
xor U4064 (N_4064,N_3211,N_2734);
and U4065 (N_4065,N_3130,N_2835);
nor U4066 (N_4066,N_2712,N_3252);
nand U4067 (N_4067,N_2521,N_3520);
or U4068 (N_4068,N_3168,N_2752);
and U4069 (N_4069,N_3541,N_2831);
nor U4070 (N_4070,N_3530,N_2433);
nand U4071 (N_4071,N_2490,N_2737);
and U4072 (N_4072,N_2403,N_2784);
or U4073 (N_4073,N_2891,N_3395);
or U4074 (N_4074,N_3556,N_3304);
nor U4075 (N_4075,N_3027,N_3497);
xor U4076 (N_4076,N_3179,N_2729);
nor U4077 (N_4077,N_2415,N_3492);
or U4078 (N_4078,N_2853,N_3425);
xor U4079 (N_4079,N_3210,N_2871);
and U4080 (N_4080,N_2697,N_2549);
and U4081 (N_4081,N_2854,N_2566);
or U4082 (N_4082,N_2953,N_2464);
and U4083 (N_4083,N_3134,N_3337);
and U4084 (N_4084,N_3409,N_2444);
or U4085 (N_4085,N_2755,N_2709);
and U4086 (N_4086,N_2661,N_2785);
nor U4087 (N_4087,N_3037,N_2909);
nand U4088 (N_4088,N_2842,N_2789);
and U4089 (N_4089,N_2699,N_2579);
xnor U4090 (N_4090,N_2594,N_2429);
nor U4091 (N_4091,N_3488,N_2950);
nand U4092 (N_4092,N_3326,N_3426);
nor U4093 (N_4093,N_2956,N_2599);
nand U4094 (N_4094,N_3365,N_2952);
nand U4095 (N_4095,N_2437,N_2677);
or U4096 (N_4096,N_3470,N_3240);
or U4097 (N_4097,N_3161,N_3356);
nand U4098 (N_4098,N_3042,N_2741);
or U4099 (N_4099,N_2915,N_2542);
and U4100 (N_4100,N_3410,N_3049);
nand U4101 (N_4101,N_2949,N_3054);
xnor U4102 (N_4102,N_3177,N_2788);
xnor U4103 (N_4103,N_2832,N_3466);
nor U4104 (N_4104,N_3549,N_2413);
nand U4105 (N_4105,N_2820,N_2833);
and U4106 (N_4106,N_3231,N_3318);
nand U4107 (N_4107,N_2710,N_2568);
or U4108 (N_4108,N_2722,N_3475);
xnor U4109 (N_4109,N_3191,N_2440);
xnor U4110 (N_4110,N_2688,N_2894);
and U4111 (N_4111,N_2535,N_3247);
or U4112 (N_4112,N_2924,N_3376);
xor U4113 (N_4113,N_3507,N_3554);
xnor U4114 (N_4114,N_3351,N_3128);
nand U4115 (N_4115,N_2583,N_2643);
or U4116 (N_4116,N_3108,N_2458);
or U4117 (N_4117,N_3135,N_2512);
nor U4118 (N_4118,N_2573,N_3156);
and U4119 (N_4119,N_2509,N_3444);
xor U4120 (N_4120,N_3452,N_2414);
nor U4121 (N_4121,N_3333,N_2574);
and U4122 (N_4122,N_3533,N_2971);
and U4123 (N_4123,N_2571,N_2844);
nor U4124 (N_4124,N_2634,N_2827);
nand U4125 (N_4125,N_3415,N_3254);
nand U4126 (N_4126,N_2546,N_2922);
xnor U4127 (N_4127,N_2420,N_3537);
xnor U4128 (N_4128,N_2916,N_3226);
nor U4129 (N_4129,N_2759,N_2977);
nand U4130 (N_4130,N_3510,N_2857);
nor U4131 (N_4131,N_3078,N_3001);
and U4132 (N_4132,N_2805,N_2903);
and U4133 (N_4133,N_2454,N_2528);
xor U4134 (N_4134,N_3589,N_3370);
nor U4135 (N_4135,N_3157,N_2461);
xnor U4136 (N_4136,N_2695,N_3164);
or U4137 (N_4137,N_2559,N_2735);
nor U4138 (N_4138,N_3178,N_2591);
or U4139 (N_4139,N_2947,N_2449);
nand U4140 (N_4140,N_3406,N_2482);
xor U4141 (N_4141,N_3447,N_2860);
nand U4142 (N_4142,N_3216,N_2868);
xnor U4143 (N_4143,N_2935,N_2561);
and U4144 (N_4144,N_2957,N_2795);
nor U4145 (N_4145,N_2881,N_3348);
nand U4146 (N_4146,N_2856,N_3394);
nor U4147 (N_4147,N_2687,N_3125);
xor U4148 (N_4148,N_2520,N_3075);
or U4149 (N_4149,N_3557,N_3461);
nor U4150 (N_4150,N_3186,N_2942);
nor U4151 (N_4151,N_2902,N_3297);
and U4152 (N_4152,N_2668,N_2955);
nand U4153 (N_4153,N_2698,N_2639);
nor U4154 (N_4154,N_3362,N_2540);
and U4155 (N_4155,N_3233,N_3413);
nand U4156 (N_4156,N_3286,N_2410);
nand U4157 (N_4157,N_2769,N_3327);
nor U4158 (N_4158,N_3255,N_3513);
nor U4159 (N_4159,N_3345,N_3273);
nand U4160 (N_4160,N_3263,N_3258);
and U4161 (N_4161,N_2636,N_3571);
or U4162 (N_4162,N_3055,N_2673);
nor U4163 (N_4163,N_3291,N_2991);
xor U4164 (N_4164,N_2974,N_3562);
and U4165 (N_4165,N_2756,N_3570);
xor U4166 (N_4166,N_2497,N_2507);
or U4167 (N_4167,N_2763,N_2496);
xor U4168 (N_4168,N_2567,N_3366);
or U4169 (N_4169,N_3352,N_3393);
and U4170 (N_4170,N_3499,N_3228);
xnor U4171 (N_4171,N_3565,N_3281);
xor U4172 (N_4172,N_2993,N_3292);
xnor U4173 (N_4173,N_3050,N_2776);
xnor U4174 (N_4174,N_3561,N_2409);
or U4175 (N_4175,N_2644,N_2620);
nor U4176 (N_4176,N_2855,N_2746);
xnor U4177 (N_4177,N_2798,N_3009);
or U4178 (N_4178,N_2442,N_2937);
and U4179 (N_4179,N_3245,N_3374);
nor U4180 (N_4180,N_2824,N_3057);
nor U4181 (N_4181,N_2944,N_2598);
nand U4182 (N_4182,N_2690,N_3346);
and U4183 (N_4183,N_3358,N_2907);
nor U4184 (N_4184,N_2657,N_3427);
nand U4185 (N_4185,N_3069,N_3527);
and U4186 (N_4186,N_2864,N_3007);
xor U4187 (N_4187,N_3511,N_2919);
and U4188 (N_4188,N_2671,N_3052);
and U4189 (N_4189,N_2754,N_3126);
xor U4190 (N_4190,N_2672,N_2477);
and U4191 (N_4191,N_2459,N_2989);
nand U4192 (N_4192,N_3175,N_2605);
nand U4193 (N_4193,N_3330,N_3474);
nand U4194 (N_4194,N_3381,N_3261);
nand U4195 (N_4195,N_3166,N_2994);
nor U4196 (N_4196,N_2486,N_2803);
nand U4197 (N_4197,N_3564,N_3347);
nor U4198 (N_4198,N_2616,N_2816);
and U4199 (N_4199,N_3101,N_2874);
nor U4200 (N_4200,N_3237,N_2632);
xnor U4201 (N_4201,N_3139,N_3350);
and U4202 (N_4202,N_2908,N_3049);
nand U4203 (N_4203,N_2725,N_2424);
xor U4204 (N_4204,N_2713,N_3213);
nor U4205 (N_4205,N_2810,N_2678);
xor U4206 (N_4206,N_2711,N_3478);
nor U4207 (N_4207,N_2464,N_3021);
and U4208 (N_4208,N_3086,N_3361);
and U4209 (N_4209,N_2424,N_3148);
and U4210 (N_4210,N_3019,N_3045);
or U4211 (N_4211,N_3537,N_3131);
nand U4212 (N_4212,N_3187,N_3479);
nor U4213 (N_4213,N_3145,N_3048);
xnor U4214 (N_4214,N_3127,N_3464);
nor U4215 (N_4215,N_2827,N_3169);
or U4216 (N_4216,N_2814,N_3088);
nor U4217 (N_4217,N_2698,N_3468);
or U4218 (N_4218,N_2879,N_2930);
or U4219 (N_4219,N_2701,N_2746);
xnor U4220 (N_4220,N_3187,N_2812);
xnor U4221 (N_4221,N_2429,N_3565);
and U4222 (N_4222,N_2760,N_2736);
xor U4223 (N_4223,N_3523,N_2511);
nor U4224 (N_4224,N_3177,N_2895);
or U4225 (N_4225,N_2788,N_3430);
and U4226 (N_4226,N_3440,N_2527);
nor U4227 (N_4227,N_2903,N_2409);
nand U4228 (N_4228,N_3101,N_3115);
nor U4229 (N_4229,N_3543,N_3348);
nand U4230 (N_4230,N_2438,N_2695);
xnor U4231 (N_4231,N_3452,N_2818);
and U4232 (N_4232,N_2962,N_3292);
xor U4233 (N_4233,N_3160,N_3153);
nand U4234 (N_4234,N_2991,N_3544);
and U4235 (N_4235,N_2755,N_3018);
nand U4236 (N_4236,N_2421,N_2819);
or U4237 (N_4237,N_2638,N_3393);
or U4238 (N_4238,N_3524,N_3025);
nor U4239 (N_4239,N_3308,N_3225);
and U4240 (N_4240,N_2990,N_2676);
and U4241 (N_4241,N_3313,N_3584);
or U4242 (N_4242,N_3494,N_3480);
nor U4243 (N_4243,N_2514,N_2444);
nand U4244 (N_4244,N_2717,N_3584);
and U4245 (N_4245,N_2612,N_3291);
or U4246 (N_4246,N_2753,N_3501);
nand U4247 (N_4247,N_2724,N_3314);
nand U4248 (N_4248,N_3420,N_3343);
nor U4249 (N_4249,N_3220,N_2615);
xor U4250 (N_4250,N_2985,N_2728);
and U4251 (N_4251,N_3538,N_2584);
nor U4252 (N_4252,N_2978,N_3299);
xor U4253 (N_4253,N_3314,N_3326);
xor U4254 (N_4254,N_3302,N_2710);
and U4255 (N_4255,N_2625,N_3375);
xor U4256 (N_4256,N_3566,N_2853);
and U4257 (N_4257,N_2575,N_3158);
nor U4258 (N_4258,N_2498,N_3068);
nand U4259 (N_4259,N_3105,N_3066);
xor U4260 (N_4260,N_3416,N_2858);
nand U4261 (N_4261,N_3347,N_2689);
or U4262 (N_4262,N_3499,N_2484);
nor U4263 (N_4263,N_2788,N_2752);
nand U4264 (N_4264,N_2668,N_3597);
nor U4265 (N_4265,N_2402,N_3554);
xnor U4266 (N_4266,N_3187,N_3378);
nor U4267 (N_4267,N_2452,N_2576);
or U4268 (N_4268,N_3013,N_3167);
nor U4269 (N_4269,N_2579,N_3380);
nor U4270 (N_4270,N_2992,N_3262);
and U4271 (N_4271,N_2485,N_3113);
and U4272 (N_4272,N_3178,N_3025);
xor U4273 (N_4273,N_2459,N_2573);
nand U4274 (N_4274,N_3298,N_3209);
xnor U4275 (N_4275,N_2815,N_3227);
and U4276 (N_4276,N_3148,N_2572);
nor U4277 (N_4277,N_2867,N_3170);
or U4278 (N_4278,N_2898,N_2481);
nor U4279 (N_4279,N_2819,N_3303);
or U4280 (N_4280,N_3212,N_3428);
or U4281 (N_4281,N_2640,N_2413);
or U4282 (N_4282,N_2547,N_3475);
or U4283 (N_4283,N_3198,N_2595);
nor U4284 (N_4284,N_2751,N_3526);
nand U4285 (N_4285,N_2994,N_3137);
and U4286 (N_4286,N_3034,N_3246);
and U4287 (N_4287,N_2704,N_2895);
xnor U4288 (N_4288,N_2520,N_2428);
nand U4289 (N_4289,N_2592,N_2892);
xnor U4290 (N_4290,N_2634,N_3410);
and U4291 (N_4291,N_3378,N_3505);
and U4292 (N_4292,N_2800,N_3495);
or U4293 (N_4293,N_3284,N_2424);
nand U4294 (N_4294,N_2622,N_3151);
xnor U4295 (N_4295,N_3171,N_3165);
nor U4296 (N_4296,N_2608,N_2700);
nand U4297 (N_4297,N_3398,N_3107);
xnor U4298 (N_4298,N_3548,N_3115);
xnor U4299 (N_4299,N_2868,N_2432);
and U4300 (N_4300,N_2565,N_3198);
or U4301 (N_4301,N_3312,N_3023);
nor U4302 (N_4302,N_3397,N_2842);
or U4303 (N_4303,N_3516,N_2703);
and U4304 (N_4304,N_2827,N_2862);
nor U4305 (N_4305,N_2969,N_2724);
or U4306 (N_4306,N_2881,N_3293);
and U4307 (N_4307,N_2761,N_3595);
or U4308 (N_4308,N_2817,N_3447);
and U4309 (N_4309,N_2454,N_2792);
xnor U4310 (N_4310,N_3262,N_2728);
and U4311 (N_4311,N_2633,N_3595);
or U4312 (N_4312,N_3590,N_3416);
nand U4313 (N_4313,N_3211,N_3544);
and U4314 (N_4314,N_3172,N_2868);
and U4315 (N_4315,N_2902,N_3427);
and U4316 (N_4316,N_2725,N_2564);
xnor U4317 (N_4317,N_3138,N_2638);
and U4318 (N_4318,N_2586,N_2605);
nand U4319 (N_4319,N_2859,N_3056);
or U4320 (N_4320,N_2824,N_2998);
nand U4321 (N_4321,N_3222,N_3225);
and U4322 (N_4322,N_2751,N_3291);
nor U4323 (N_4323,N_2783,N_2893);
nand U4324 (N_4324,N_3407,N_2669);
nand U4325 (N_4325,N_3389,N_3152);
xnor U4326 (N_4326,N_3081,N_2871);
xnor U4327 (N_4327,N_3219,N_3217);
and U4328 (N_4328,N_2887,N_3409);
nand U4329 (N_4329,N_3345,N_3464);
or U4330 (N_4330,N_2813,N_2440);
nor U4331 (N_4331,N_3527,N_2719);
nor U4332 (N_4332,N_2672,N_3398);
xor U4333 (N_4333,N_3152,N_3201);
and U4334 (N_4334,N_3027,N_3396);
xor U4335 (N_4335,N_3264,N_3048);
and U4336 (N_4336,N_2956,N_2586);
nand U4337 (N_4337,N_3036,N_3249);
and U4338 (N_4338,N_2656,N_3382);
xor U4339 (N_4339,N_3591,N_3142);
nand U4340 (N_4340,N_3094,N_3233);
or U4341 (N_4341,N_2901,N_2934);
xnor U4342 (N_4342,N_2990,N_3127);
nand U4343 (N_4343,N_3374,N_3027);
nor U4344 (N_4344,N_3149,N_2458);
nand U4345 (N_4345,N_3578,N_2486);
xor U4346 (N_4346,N_3377,N_2573);
xor U4347 (N_4347,N_2986,N_2489);
nor U4348 (N_4348,N_2411,N_3313);
xnor U4349 (N_4349,N_3371,N_3409);
or U4350 (N_4350,N_3581,N_2489);
xnor U4351 (N_4351,N_3029,N_2404);
nand U4352 (N_4352,N_3235,N_2478);
or U4353 (N_4353,N_2953,N_2525);
or U4354 (N_4354,N_3023,N_3497);
or U4355 (N_4355,N_3103,N_3298);
and U4356 (N_4356,N_3344,N_3340);
or U4357 (N_4357,N_3048,N_2859);
nor U4358 (N_4358,N_2763,N_3488);
or U4359 (N_4359,N_3001,N_3400);
nand U4360 (N_4360,N_3367,N_2982);
nand U4361 (N_4361,N_3038,N_3107);
and U4362 (N_4362,N_2957,N_2489);
xnor U4363 (N_4363,N_2918,N_3411);
nor U4364 (N_4364,N_2757,N_3364);
nand U4365 (N_4365,N_3169,N_2579);
or U4366 (N_4366,N_3404,N_3281);
nor U4367 (N_4367,N_2695,N_3112);
or U4368 (N_4368,N_3581,N_3409);
xnor U4369 (N_4369,N_2811,N_2714);
xor U4370 (N_4370,N_3587,N_2661);
xor U4371 (N_4371,N_3404,N_2554);
nor U4372 (N_4372,N_3416,N_2870);
nor U4373 (N_4373,N_2989,N_2944);
xor U4374 (N_4374,N_2809,N_3031);
nand U4375 (N_4375,N_3420,N_3406);
and U4376 (N_4376,N_3244,N_3398);
and U4377 (N_4377,N_3374,N_3304);
and U4378 (N_4378,N_2829,N_2770);
or U4379 (N_4379,N_2624,N_2535);
xnor U4380 (N_4380,N_2730,N_3582);
xor U4381 (N_4381,N_3509,N_2446);
nor U4382 (N_4382,N_2983,N_2462);
nor U4383 (N_4383,N_2413,N_3533);
and U4384 (N_4384,N_3330,N_3031);
nand U4385 (N_4385,N_2513,N_2484);
nand U4386 (N_4386,N_3257,N_2705);
nor U4387 (N_4387,N_2949,N_2627);
or U4388 (N_4388,N_3164,N_3262);
nor U4389 (N_4389,N_3022,N_3511);
xor U4390 (N_4390,N_3403,N_2445);
or U4391 (N_4391,N_2667,N_2692);
nand U4392 (N_4392,N_2551,N_3030);
nand U4393 (N_4393,N_3468,N_3472);
and U4394 (N_4394,N_3534,N_2935);
or U4395 (N_4395,N_3190,N_3063);
xor U4396 (N_4396,N_3515,N_3125);
nand U4397 (N_4397,N_3070,N_3139);
xnor U4398 (N_4398,N_2418,N_3178);
and U4399 (N_4399,N_3168,N_3083);
or U4400 (N_4400,N_2492,N_3472);
nor U4401 (N_4401,N_2757,N_2539);
xor U4402 (N_4402,N_3325,N_3423);
nand U4403 (N_4403,N_2968,N_3124);
nor U4404 (N_4404,N_3406,N_2871);
and U4405 (N_4405,N_3287,N_2969);
nor U4406 (N_4406,N_3050,N_2622);
and U4407 (N_4407,N_2720,N_3318);
nor U4408 (N_4408,N_3432,N_3353);
nand U4409 (N_4409,N_3569,N_2756);
xnor U4410 (N_4410,N_3540,N_3154);
nand U4411 (N_4411,N_2837,N_2681);
or U4412 (N_4412,N_3431,N_2671);
and U4413 (N_4413,N_3256,N_2569);
or U4414 (N_4414,N_3301,N_3351);
nand U4415 (N_4415,N_3242,N_2920);
and U4416 (N_4416,N_2853,N_2774);
or U4417 (N_4417,N_2779,N_3120);
or U4418 (N_4418,N_2463,N_2915);
nor U4419 (N_4419,N_3411,N_2795);
and U4420 (N_4420,N_3330,N_2652);
or U4421 (N_4421,N_2671,N_2549);
nand U4422 (N_4422,N_3599,N_3331);
or U4423 (N_4423,N_2677,N_2538);
and U4424 (N_4424,N_3319,N_3475);
and U4425 (N_4425,N_3069,N_2781);
and U4426 (N_4426,N_3162,N_2591);
or U4427 (N_4427,N_3100,N_2807);
and U4428 (N_4428,N_3598,N_3022);
xnor U4429 (N_4429,N_2888,N_3585);
nand U4430 (N_4430,N_3004,N_2655);
and U4431 (N_4431,N_3273,N_2452);
or U4432 (N_4432,N_2416,N_3336);
and U4433 (N_4433,N_2560,N_2617);
nor U4434 (N_4434,N_3018,N_3555);
or U4435 (N_4435,N_2988,N_3112);
xor U4436 (N_4436,N_3101,N_2663);
and U4437 (N_4437,N_2517,N_3424);
and U4438 (N_4438,N_3030,N_2403);
nand U4439 (N_4439,N_3539,N_2430);
or U4440 (N_4440,N_3078,N_2579);
nor U4441 (N_4441,N_2575,N_2922);
nor U4442 (N_4442,N_2474,N_2430);
nor U4443 (N_4443,N_2501,N_3555);
nand U4444 (N_4444,N_3192,N_3282);
xnor U4445 (N_4445,N_2496,N_2418);
xnor U4446 (N_4446,N_3203,N_3491);
nor U4447 (N_4447,N_3160,N_3454);
xor U4448 (N_4448,N_2609,N_2672);
xor U4449 (N_4449,N_3503,N_3444);
nand U4450 (N_4450,N_2481,N_3218);
or U4451 (N_4451,N_3273,N_3227);
and U4452 (N_4452,N_2519,N_2614);
nor U4453 (N_4453,N_2756,N_3231);
and U4454 (N_4454,N_3545,N_2890);
xnor U4455 (N_4455,N_2920,N_2903);
xnor U4456 (N_4456,N_3322,N_2469);
or U4457 (N_4457,N_3530,N_2949);
and U4458 (N_4458,N_3234,N_3033);
and U4459 (N_4459,N_3327,N_2512);
xnor U4460 (N_4460,N_2607,N_2675);
nor U4461 (N_4461,N_2698,N_2653);
nor U4462 (N_4462,N_3171,N_3599);
nand U4463 (N_4463,N_3494,N_2736);
or U4464 (N_4464,N_3512,N_2909);
and U4465 (N_4465,N_2637,N_3465);
nor U4466 (N_4466,N_2916,N_2457);
nand U4467 (N_4467,N_2481,N_3447);
xor U4468 (N_4468,N_3235,N_3123);
and U4469 (N_4469,N_2483,N_3480);
or U4470 (N_4470,N_2635,N_2956);
nand U4471 (N_4471,N_2876,N_2967);
nor U4472 (N_4472,N_2811,N_3500);
nand U4473 (N_4473,N_2522,N_2720);
and U4474 (N_4474,N_3230,N_3187);
and U4475 (N_4475,N_2421,N_2815);
nand U4476 (N_4476,N_2951,N_3468);
nand U4477 (N_4477,N_3560,N_2926);
nor U4478 (N_4478,N_3089,N_3283);
nor U4479 (N_4479,N_2843,N_3579);
nor U4480 (N_4480,N_3521,N_2532);
and U4481 (N_4481,N_2928,N_2443);
nand U4482 (N_4482,N_3333,N_2439);
or U4483 (N_4483,N_3593,N_2700);
xor U4484 (N_4484,N_3220,N_3102);
nor U4485 (N_4485,N_2566,N_2428);
nand U4486 (N_4486,N_2688,N_3431);
and U4487 (N_4487,N_2411,N_2814);
nor U4488 (N_4488,N_2923,N_3133);
nand U4489 (N_4489,N_3191,N_2675);
or U4490 (N_4490,N_3507,N_2743);
nor U4491 (N_4491,N_3137,N_2527);
nor U4492 (N_4492,N_3418,N_2767);
xnor U4493 (N_4493,N_3346,N_3120);
xnor U4494 (N_4494,N_2611,N_2849);
nor U4495 (N_4495,N_3220,N_2983);
nor U4496 (N_4496,N_3252,N_3118);
or U4497 (N_4497,N_3441,N_2582);
or U4498 (N_4498,N_3071,N_3073);
nand U4499 (N_4499,N_3321,N_3581);
xor U4500 (N_4500,N_2656,N_3542);
and U4501 (N_4501,N_3182,N_3316);
and U4502 (N_4502,N_3355,N_2946);
xnor U4503 (N_4503,N_3449,N_2922);
nand U4504 (N_4504,N_2410,N_3113);
and U4505 (N_4505,N_3190,N_2511);
and U4506 (N_4506,N_2586,N_2596);
nand U4507 (N_4507,N_3298,N_3285);
nand U4508 (N_4508,N_2692,N_3026);
nor U4509 (N_4509,N_2803,N_2602);
nor U4510 (N_4510,N_2720,N_2987);
xnor U4511 (N_4511,N_2682,N_2867);
nor U4512 (N_4512,N_2792,N_3583);
nor U4513 (N_4513,N_2690,N_2937);
or U4514 (N_4514,N_2950,N_3009);
or U4515 (N_4515,N_2502,N_2678);
xnor U4516 (N_4516,N_2818,N_2471);
and U4517 (N_4517,N_2690,N_3360);
and U4518 (N_4518,N_2462,N_3104);
nor U4519 (N_4519,N_2742,N_3135);
xor U4520 (N_4520,N_2845,N_3352);
nand U4521 (N_4521,N_2924,N_3188);
and U4522 (N_4522,N_2915,N_2976);
nand U4523 (N_4523,N_3420,N_3325);
nand U4524 (N_4524,N_3478,N_3075);
or U4525 (N_4525,N_3228,N_2444);
and U4526 (N_4526,N_3492,N_2866);
nand U4527 (N_4527,N_3299,N_3521);
and U4528 (N_4528,N_2524,N_3489);
and U4529 (N_4529,N_2760,N_2885);
and U4530 (N_4530,N_3547,N_3053);
nand U4531 (N_4531,N_2859,N_2430);
xnor U4532 (N_4532,N_3210,N_2553);
or U4533 (N_4533,N_3222,N_3299);
and U4534 (N_4534,N_2423,N_2902);
xor U4535 (N_4535,N_3456,N_2705);
xnor U4536 (N_4536,N_2508,N_2857);
xor U4537 (N_4537,N_3009,N_3049);
nor U4538 (N_4538,N_3534,N_2899);
xnor U4539 (N_4539,N_2778,N_2496);
or U4540 (N_4540,N_2661,N_3334);
nand U4541 (N_4541,N_2779,N_2616);
or U4542 (N_4542,N_3359,N_2784);
nand U4543 (N_4543,N_2518,N_3497);
nand U4544 (N_4544,N_3220,N_2952);
nand U4545 (N_4545,N_3399,N_3004);
nor U4546 (N_4546,N_2413,N_2650);
nand U4547 (N_4547,N_3062,N_2857);
xor U4548 (N_4548,N_3025,N_2822);
xor U4549 (N_4549,N_2628,N_3552);
xor U4550 (N_4550,N_3577,N_2915);
nand U4551 (N_4551,N_2495,N_2615);
or U4552 (N_4552,N_2537,N_3463);
nand U4553 (N_4553,N_3265,N_3371);
and U4554 (N_4554,N_2619,N_3122);
nand U4555 (N_4555,N_3285,N_2907);
xnor U4556 (N_4556,N_2777,N_2792);
xnor U4557 (N_4557,N_2645,N_3225);
nor U4558 (N_4558,N_2499,N_2734);
and U4559 (N_4559,N_3192,N_3349);
and U4560 (N_4560,N_2476,N_2743);
xor U4561 (N_4561,N_2933,N_2868);
or U4562 (N_4562,N_2511,N_2660);
or U4563 (N_4563,N_3421,N_2651);
and U4564 (N_4564,N_3509,N_2407);
nor U4565 (N_4565,N_2861,N_2883);
xor U4566 (N_4566,N_3420,N_2740);
nand U4567 (N_4567,N_3073,N_3205);
xnor U4568 (N_4568,N_2761,N_3122);
xnor U4569 (N_4569,N_3582,N_2511);
and U4570 (N_4570,N_2467,N_2553);
xnor U4571 (N_4571,N_3028,N_3086);
nand U4572 (N_4572,N_3373,N_2688);
nor U4573 (N_4573,N_3265,N_2710);
nand U4574 (N_4574,N_3224,N_2440);
or U4575 (N_4575,N_3102,N_3226);
and U4576 (N_4576,N_3474,N_2835);
or U4577 (N_4577,N_3407,N_3317);
xnor U4578 (N_4578,N_2964,N_3519);
xnor U4579 (N_4579,N_2828,N_3578);
and U4580 (N_4580,N_2612,N_2787);
or U4581 (N_4581,N_3443,N_2951);
nor U4582 (N_4582,N_2737,N_2625);
xor U4583 (N_4583,N_2715,N_3586);
nor U4584 (N_4584,N_3321,N_3549);
and U4585 (N_4585,N_2618,N_3582);
or U4586 (N_4586,N_3148,N_2728);
or U4587 (N_4587,N_3419,N_3563);
or U4588 (N_4588,N_3558,N_2809);
or U4589 (N_4589,N_3557,N_2797);
nand U4590 (N_4590,N_2520,N_3070);
nand U4591 (N_4591,N_3346,N_3272);
or U4592 (N_4592,N_3541,N_2777);
or U4593 (N_4593,N_2911,N_3214);
xor U4594 (N_4594,N_2611,N_2754);
nor U4595 (N_4595,N_3485,N_2438);
xnor U4596 (N_4596,N_3028,N_3537);
or U4597 (N_4597,N_2507,N_3253);
nor U4598 (N_4598,N_2511,N_3435);
nor U4599 (N_4599,N_3246,N_2591);
and U4600 (N_4600,N_3098,N_3313);
nand U4601 (N_4601,N_2644,N_2701);
and U4602 (N_4602,N_2653,N_3370);
nand U4603 (N_4603,N_2918,N_2815);
or U4604 (N_4604,N_3360,N_2479);
nand U4605 (N_4605,N_3104,N_3205);
nor U4606 (N_4606,N_3591,N_2540);
and U4607 (N_4607,N_3125,N_3211);
nand U4608 (N_4608,N_2648,N_2981);
nor U4609 (N_4609,N_3526,N_3309);
nor U4610 (N_4610,N_3085,N_2679);
nand U4611 (N_4611,N_3001,N_2926);
nor U4612 (N_4612,N_2763,N_3407);
or U4613 (N_4613,N_3469,N_3531);
or U4614 (N_4614,N_2854,N_3448);
and U4615 (N_4615,N_3000,N_2564);
nand U4616 (N_4616,N_2758,N_2615);
or U4617 (N_4617,N_3044,N_2965);
nor U4618 (N_4618,N_3474,N_3079);
nor U4619 (N_4619,N_2480,N_3103);
or U4620 (N_4620,N_3172,N_2623);
and U4621 (N_4621,N_2548,N_3247);
and U4622 (N_4622,N_3148,N_2771);
nor U4623 (N_4623,N_2986,N_2755);
nor U4624 (N_4624,N_3509,N_2907);
and U4625 (N_4625,N_3001,N_3027);
xor U4626 (N_4626,N_2475,N_3547);
and U4627 (N_4627,N_2838,N_3213);
nor U4628 (N_4628,N_3427,N_3014);
and U4629 (N_4629,N_2980,N_2929);
nor U4630 (N_4630,N_3241,N_3046);
and U4631 (N_4631,N_2579,N_2661);
nand U4632 (N_4632,N_2808,N_3382);
or U4633 (N_4633,N_3568,N_3561);
nand U4634 (N_4634,N_2524,N_3547);
xor U4635 (N_4635,N_2749,N_3018);
nor U4636 (N_4636,N_2998,N_3568);
nand U4637 (N_4637,N_3266,N_3146);
nor U4638 (N_4638,N_3389,N_3438);
or U4639 (N_4639,N_2818,N_2908);
or U4640 (N_4640,N_2802,N_2944);
nor U4641 (N_4641,N_3079,N_3019);
nand U4642 (N_4642,N_2786,N_3265);
nand U4643 (N_4643,N_3028,N_2665);
nand U4644 (N_4644,N_3494,N_3495);
or U4645 (N_4645,N_3403,N_2684);
nand U4646 (N_4646,N_3167,N_3402);
or U4647 (N_4647,N_2890,N_3008);
and U4648 (N_4648,N_3218,N_3032);
xor U4649 (N_4649,N_3491,N_3369);
or U4650 (N_4650,N_3568,N_3090);
and U4651 (N_4651,N_2426,N_2770);
or U4652 (N_4652,N_2824,N_2930);
or U4653 (N_4653,N_3064,N_3571);
xnor U4654 (N_4654,N_3595,N_2440);
and U4655 (N_4655,N_2449,N_3225);
nand U4656 (N_4656,N_3353,N_2548);
and U4657 (N_4657,N_3594,N_3390);
nor U4658 (N_4658,N_2927,N_3329);
nor U4659 (N_4659,N_2834,N_3513);
nand U4660 (N_4660,N_3028,N_2788);
or U4661 (N_4661,N_2940,N_2502);
nand U4662 (N_4662,N_3118,N_2893);
and U4663 (N_4663,N_3169,N_2923);
and U4664 (N_4664,N_2740,N_2718);
xnor U4665 (N_4665,N_3001,N_2529);
and U4666 (N_4666,N_2963,N_3446);
nor U4667 (N_4667,N_2807,N_3214);
and U4668 (N_4668,N_3257,N_2585);
nor U4669 (N_4669,N_3382,N_3235);
xor U4670 (N_4670,N_3236,N_2412);
or U4671 (N_4671,N_2810,N_3507);
nand U4672 (N_4672,N_2706,N_3103);
xor U4673 (N_4673,N_3300,N_3247);
xnor U4674 (N_4674,N_2423,N_2716);
or U4675 (N_4675,N_3491,N_2669);
or U4676 (N_4676,N_2506,N_2853);
nand U4677 (N_4677,N_3306,N_3129);
and U4678 (N_4678,N_2604,N_2925);
or U4679 (N_4679,N_3292,N_3587);
nand U4680 (N_4680,N_3141,N_2453);
xnor U4681 (N_4681,N_2608,N_2964);
xnor U4682 (N_4682,N_3015,N_3254);
nand U4683 (N_4683,N_3595,N_2400);
and U4684 (N_4684,N_3529,N_2987);
nand U4685 (N_4685,N_3190,N_2750);
xnor U4686 (N_4686,N_3232,N_3237);
or U4687 (N_4687,N_2539,N_2864);
and U4688 (N_4688,N_2736,N_2568);
or U4689 (N_4689,N_2922,N_3009);
or U4690 (N_4690,N_2543,N_3345);
or U4691 (N_4691,N_3417,N_3396);
nand U4692 (N_4692,N_3006,N_3159);
nand U4693 (N_4693,N_2958,N_2638);
nor U4694 (N_4694,N_3300,N_2690);
nor U4695 (N_4695,N_2552,N_3259);
or U4696 (N_4696,N_3267,N_2706);
nor U4697 (N_4697,N_3331,N_3334);
nand U4698 (N_4698,N_2976,N_3536);
nand U4699 (N_4699,N_2517,N_2506);
nor U4700 (N_4700,N_2853,N_3100);
or U4701 (N_4701,N_2989,N_2518);
nor U4702 (N_4702,N_3090,N_2992);
nand U4703 (N_4703,N_2638,N_2810);
xor U4704 (N_4704,N_2858,N_3578);
nor U4705 (N_4705,N_3208,N_2598);
or U4706 (N_4706,N_2872,N_3481);
or U4707 (N_4707,N_3339,N_3069);
or U4708 (N_4708,N_2511,N_2607);
xor U4709 (N_4709,N_3184,N_2537);
nor U4710 (N_4710,N_2448,N_3202);
xor U4711 (N_4711,N_3045,N_3306);
and U4712 (N_4712,N_3351,N_3002);
and U4713 (N_4713,N_3140,N_3186);
nor U4714 (N_4714,N_3544,N_2686);
nand U4715 (N_4715,N_3189,N_3127);
or U4716 (N_4716,N_2654,N_2766);
or U4717 (N_4717,N_2901,N_2522);
or U4718 (N_4718,N_2943,N_3217);
and U4719 (N_4719,N_2904,N_2464);
nand U4720 (N_4720,N_2435,N_3442);
nor U4721 (N_4721,N_2461,N_3477);
nand U4722 (N_4722,N_3562,N_3523);
nor U4723 (N_4723,N_3102,N_3190);
nor U4724 (N_4724,N_2635,N_2530);
nor U4725 (N_4725,N_3595,N_2809);
nor U4726 (N_4726,N_2678,N_2456);
or U4727 (N_4727,N_3490,N_2824);
and U4728 (N_4728,N_2583,N_2964);
nor U4729 (N_4729,N_2595,N_2568);
nand U4730 (N_4730,N_2584,N_2859);
nand U4731 (N_4731,N_2844,N_2728);
nor U4732 (N_4732,N_2514,N_3285);
or U4733 (N_4733,N_2929,N_2500);
nand U4734 (N_4734,N_3272,N_2675);
or U4735 (N_4735,N_2708,N_3504);
nor U4736 (N_4736,N_2535,N_3092);
xnor U4737 (N_4737,N_2526,N_2865);
or U4738 (N_4738,N_2836,N_2985);
nand U4739 (N_4739,N_2778,N_2692);
and U4740 (N_4740,N_2459,N_2557);
xor U4741 (N_4741,N_3294,N_2774);
nand U4742 (N_4742,N_2522,N_3146);
nor U4743 (N_4743,N_3075,N_2468);
nor U4744 (N_4744,N_2411,N_3271);
or U4745 (N_4745,N_2931,N_3392);
or U4746 (N_4746,N_3183,N_3158);
and U4747 (N_4747,N_2667,N_2409);
and U4748 (N_4748,N_2552,N_3460);
nand U4749 (N_4749,N_2738,N_2586);
nand U4750 (N_4750,N_3265,N_3033);
xnor U4751 (N_4751,N_3491,N_3388);
nor U4752 (N_4752,N_3335,N_3080);
xnor U4753 (N_4753,N_3164,N_3136);
xor U4754 (N_4754,N_3423,N_3095);
nand U4755 (N_4755,N_3296,N_3407);
nor U4756 (N_4756,N_2426,N_3092);
xnor U4757 (N_4757,N_3509,N_2995);
or U4758 (N_4758,N_2550,N_3117);
nor U4759 (N_4759,N_3479,N_3165);
nor U4760 (N_4760,N_3553,N_2920);
xnor U4761 (N_4761,N_3171,N_2753);
nand U4762 (N_4762,N_3548,N_3164);
nor U4763 (N_4763,N_2705,N_2621);
nor U4764 (N_4764,N_3418,N_2443);
xor U4765 (N_4765,N_3002,N_3017);
nor U4766 (N_4766,N_3454,N_2656);
or U4767 (N_4767,N_2642,N_3564);
nand U4768 (N_4768,N_2727,N_2756);
xnor U4769 (N_4769,N_2982,N_3470);
or U4770 (N_4770,N_2820,N_2607);
and U4771 (N_4771,N_2835,N_2832);
nor U4772 (N_4772,N_3544,N_2744);
and U4773 (N_4773,N_2759,N_3350);
xor U4774 (N_4774,N_2437,N_3259);
and U4775 (N_4775,N_2743,N_3451);
xnor U4776 (N_4776,N_2652,N_2616);
nor U4777 (N_4777,N_2584,N_3113);
or U4778 (N_4778,N_2471,N_2435);
nor U4779 (N_4779,N_2580,N_3297);
or U4780 (N_4780,N_2982,N_3484);
nand U4781 (N_4781,N_2833,N_3405);
and U4782 (N_4782,N_2744,N_2601);
nand U4783 (N_4783,N_3575,N_3521);
or U4784 (N_4784,N_3398,N_3405);
nor U4785 (N_4785,N_2523,N_3119);
xor U4786 (N_4786,N_2724,N_2505);
or U4787 (N_4787,N_2883,N_3590);
xnor U4788 (N_4788,N_2881,N_3458);
xor U4789 (N_4789,N_2430,N_2870);
nand U4790 (N_4790,N_2720,N_3180);
xnor U4791 (N_4791,N_3262,N_3347);
or U4792 (N_4792,N_2517,N_2991);
nor U4793 (N_4793,N_3112,N_3345);
and U4794 (N_4794,N_2946,N_3031);
nor U4795 (N_4795,N_3333,N_2584);
and U4796 (N_4796,N_2833,N_3347);
xor U4797 (N_4797,N_3310,N_3089);
nand U4798 (N_4798,N_3383,N_3380);
xnor U4799 (N_4799,N_2568,N_2669);
nand U4800 (N_4800,N_3947,N_3723);
or U4801 (N_4801,N_4731,N_3914);
nor U4802 (N_4802,N_3776,N_4673);
nand U4803 (N_4803,N_3644,N_4751);
and U4804 (N_4804,N_3890,N_4363);
xor U4805 (N_4805,N_4374,N_4015);
nand U4806 (N_4806,N_4065,N_4432);
xnor U4807 (N_4807,N_3635,N_4658);
nor U4808 (N_4808,N_3604,N_4072);
xor U4809 (N_4809,N_4637,N_4055);
nor U4810 (N_4810,N_4563,N_4570);
nand U4811 (N_4811,N_4586,N_3922);
or U4812 (N_4812,N_3896,N_3891);
nand U4813 (N_4813,N_4705,N_4499);
or U4814 (N_4814,N_4041,N_3892);
nor U4815 (N_4815,N_4361,N_4407);
or U4816 (N_4816,N_4051,N_3984);
nor U4817 (N_4817,N_4423,N_3902);
and U4818 (N_4818,N_4193,N_4201);
nand U4819 (N_4819,N_3870,N_3679);
xnor U4820 (N_4820,N_4300,N_3652);
xnor U4821 (N_4821,N_4073,N_4607);
xor U4822 (N_4822,N_4305,N_3658);
and U4823 (N_4823,N_4153,N_4270);
or U4824 (N_4824,N_3881,N_4544);
nor U4825 (N_4825,N_4319,N_4483);
xor U4826 (N_4826,N_3729,N_4753);
xnor U4827 (N_4827,N_3805,N_4220);
nand U4828 (N_4828,N_4615,N_4525);
and U4829 (N_4829,N_4265,N_4160);
or U4830 (N_4830,N_4442,N_4140);
nor U4831 (N_4831,N_4333,N_4258);
xor U4832 (N_4832,N_3637,N_4727);
or U4833 (N_4833,N_4368,N_4448);
xnor U4834 (N_4834,N_4500,N_3919);
nor U4835 (N_4835,N_4094,N_4137);
and U4836 (N_4836,N_4564,N_4697);
and U4837 (N_4837,N_4578,N_3921);
nor U4838 (N_4838,N_4548,N_4255);
or U4839 (N_4839,N_4659,N_4004);
and U4840 (N_4840,N_3838,N_3960);
or U4841 (N_4841,N_4491,N_4469);
nor U4842 (N_4842,N_3704,N_4622);
xor U4843 (N_4843,N_4005,N_4164);
or U4844 (N_4844,N_4696,N_4032);
nor U4845 (N_4845,N_4117,N_3707);
nor U4846 (N_4846,N_4463,N_4262);
and U4847 (N_4847,N_4416,N_3811);
and U4848 (N_4848,N_4735,N_4334);
xor U4849 (N_4849,N_4694,N_4415);
nand U4850 (N_4850,N_4272,N_4573);
nor U4851 (N_4851,N_3972,N_4326);
xnor U4852 (N_4852,N_4531,N_4708);
or U4853 (N_4853,N_4211,N_3760);
nand U4854 (N_4854,N_3939,N_4171);
or U4855 (N_4855,N_4046,N_3906);
or U4856 (N_4856,N_3730,N_4189);
nand U4857 (N_4857,N_4760,N_4489);
nand U4858 (N_4858,N_4386,N_4454);
and U4859 (N_4859,N_4278,N_4769);
or U4860 (N_4860,N_4438,N_3618);
nor U4861 (N_4861,N_3852,N_4188);
or U4862 (N_4862,N_4605,N_3950);
and U4863 (N_4863,N_4453,N_4667);
nand U4864 (N_4864,N_4232,N_4569);
and U4865 (N_4865,N_3755,N_4774);
or U4866 (N_4866,N_4641,N_4468);
or U4867 (N_4867,N_3695,N_3630);
nand U4868 (N_4868,N_3908,N_4179);
or U4869 (N_4869,N_4308,N_4204);
and U4870 (N_4870,N_3886,N_3989);
or U4871 (N_4871,N_3762,N_4379);
xor U4872 (N_4872,N_4657,N_4192);
xor U4873 (N_4873,N_4364,N_4090);
nor U4874 (N_4874,N_4693,N_4481);
nand U4875 (N_4875,N_4547,N_4150);
xnor U4876 (N_4876,N_3705,N_3844);
and U4877 (N_4877,N_4465,N_4620);
nor U4878 (N_4878,N_4163,N_4585);
or U4879 (N_4879,N_3834,N_4449);
xnor U4880 (N_4880,N_3994,N_4538);
nand U4881 (N_4881,N_4422,N_3779);
nand U4882 (N_4882,N_4409,N_3615);
and U4883 (N_4883,N_4315,N_3692);
or U4884 (N_4884,N_4619,N_4329);
xor U4885 (N_4885,N_4011,N_4384);
xor U4886 (N_4886,N_4207,N_4277);
nor U4887 (N_4887,N_4116,N_4035);
xnor U4888 (N_4888,N_3636,N_4097);
and U4889 (N_4889,N_4478,N_4391);
and U4890 (N_4890,N_3613,N_4248);
nand U4891 (N_4891,N_4310,N_4624);
xor U4892 (N_4892,N_4691,N_4718);
and U4893 (N_4893,N_4758,N_4653);
and U4894 (N_4894,N_3653,N_4555);
nor U4895 (N_4895,N_4515,N_4664);
and U4896 (N_4896,N_3968,N_3926);
nand U4897 (N_4897,N_3718,N_4053);
nand U4898 (N_4898,N_4723,N_4195);
nand U4899 (N_4899,N_4459,N_3976);
nand U4900 (N_4900,N_4318,N_3975);
or U4901 (N_4901,N_4047,N_4429);
or U4902 (N_4902,N_4689,N_3693);
xor U4903 (N_4903,N_4155,N_4773);
xor U4904 (N_4904,N_3710,N_3807);
xor U4905 (N_4905,N_4796,N_4467);
nand U4906 (N_4906,N_3985,N_4063);
nor U4907 (N_4907,N_3845,N_4198);
and U4908 (N_4908,N_4001,N_3849);
or U4909 (N_4909,N_3702,N_4381);
xnor U4910 (N_4910,N_3943,N_3715);
and U4911 (N_4911,N_4768,N_3874);
or U4912 (N_4912,N_3664,N_4746);
xnor U4913 (N_4913,N_3603,N_4599);
or U4914 (N_4914,N_4743,N_3753);
nand U4915 (N_4915,N_4686,N_4572);
or U4916 (N_4916,N_4021,N_3750);
or U4917 (N_4917,N_4427,N_3732);
and U4918 (N_4918,N_3769,N_4656);
nand U4919 (N_4919,N_4726,N_4335);
nor U4920 (N_4920,N_3856,N_4301);
and U4921 (N_4921,N_3969,N_4474);
xor U4922 (N_4922,N_3713,N_3859);
and U4923 (N_4923,N_4722,N_3864);
xor U4924 (N_4924,N_3949,N_4725);
and U4925 (N_4925,N_3833,N_4492);
nand U4926 (N_4926,N_4102,N_4156);
nand U4927 (N_4927,N_4304,N_3792);
and U4928 (N_4928,N_3764,N_4575);
xor U4929 (N_4929,N_3946,N_4792);
nor U4930 (N_4930,N_3818,N_4762);
nor U4931 (N_4931,N_4124,N_4370);
xor U4932 (N_4932,N_4212,N_3809);
or U4933 (N_4933,N_4707,N_4321);
xnor U4934 (N_4934,N_3773,N_4601);
xnor U4935 (N_4935,N_4222,N_3829);
nor U4936 (N_4936,N_3823,N_4505);
nor U4937 (N_4937,N_4238,N_4397);
xor U4938 (N_4938,N_3673,N_3749);
nor U4939 (N_4939,N_4190,N_3677);
and U4940 (N_4940,N_3726,N_4518);
nor U4941 (N_4941,N_3662,N_3665);
or U4942 (N_4942,N_3815,N_4299);
and U4943 (N_4943,N_4181,N_3940);
xnor U4944 (N_4944,N_4733,N_4458);
nor U4945 (N_4945,N_3991,N_4236);
and U4946 (N_4946,N_4464,N_3952);
nor U4947 (N_4947,N_4439,N_4230);
or U4948 (N_4948,N_3992,N_4100);
and U4949 (N_4949,N_4085,N_4522);
or U4950 (N_4950,N_4710,N_3721);
nand U4951 (N_4951,N_4413,N_4777);
or U4952 (N_4952,N_3682,N_3909);
nand U4953 (N_4953,N_4023,N_3619);
nor U4954 (N_4954,N_4594,N_4057);
xnor U4955 (N_4955,N_4676,N_4237);
or U4956 (N_4956,N_3782,N_4376);
and U4957 (N_4957,N_3904,N_4618);
xor U4958 (N_4958,N_4147,N_3649);
or U4959 (N_4959,N_3915,N_4457);
and U4960 (N_4960,N_4681,N_4152);
nor U4961 (N_4961,N_3967,N_3885);
nand U4962 (N_4962,N_3611,N_4730);
or U4963 (N_4963,N_3614,N_3607);
nor U4964 (N_4964,N_4685,N_4486);
xnor U4965 (N_4965,N_4480,N_4034);
nand U4966 (N_4966,N_4672,N_3822);
or U4967 (N_4967,N_3962,N_3990);
xnor U4968 (N_4968,N_3785,N_4744);
nor U4969 (N_4969,N_4075,N_3798);
and U4970 (N_4970,N_3888,N_4396);
or U4971 (N_4971,N_4446,N_4614);
or U4972 (N_4972,N_4695,N_4497);
or U4973 (N_4973,N_4706,N_4789);
xor U4974 (N_4974,N_4540,N_4663);
xor U4975 (N_4975,N_3629,N_3736);
or U4976 (N_4976,N_3802,N_3795);
and U4977 (N_4977,N_3741,N_3646);
xor U4978 (N_4978,N_4530,N_4332);
and U4979 (N_4979,N_4025,N_3907);
nor U4980 (N_4980,N_4249,N_3767);
nor U4981 (N_4981,N_4290,N_4349);
nand U4982 (N_4982,N_4093,N_4020);
nand U4983 (N_4983,N_3851,N_4761);
or U4984 (N_4984,N_4780,N_4286);
nor U4985 (N_4985,N_4040,N_4354);
xnor U4986 (N_4986,N_4408,N_4141);
xnor U4987 (N_4987,N_3625,N_3731);
and U4988 (N_4988,N_4729,N_3772);
or U4989 (N_4989,N_4136,N_4414);
nor U4990 (N_4990,N_4214,N_4008);
xnor U4991 (N_4991,N_4394,N_4307);
xor U4992 (N_4992,N_4024,N_3979);
and U4993 (N_4993,N_4581,N_4510);
or U4994 (N_4994,N_4552,N_4677);
or U4995 (N_4995,N_3935,N_3880);
xor U4996 (N_4996,N_4610,N_3757);
and U4997 (N_4997,N_4461,N_4567);
nor U4998 (N_4998,N_4081,N_4353);
nor U4999 (N_4999,N_4395,N_4595);
or U5000 (N_5000,N_4640,N_4279);
or U5001 (N_5001,N_4589,N_3812);
or U5002 (N_5002,N_3956,N_3694);
and U5003 (N_5003,N_4553,N_4247);
and U5004 (N_5004,N_4297,N_3642);
nand U5005 (N_5005,N_3810,N_3806);
or U5006 (N_5006,N_4635,N_4782);
or U5007 (N_5007,N_4360,N_4042);
and U5008 (N_5008,N_4330,N_3790);
nor U5009 (N_5009,N_3712,N_3944);
nor U5010 (N_5010,N_4148,N_3987);
nor U5011 (N_5011,N_4403,N_3836);
xor U5012 (N_5012,N_4609,N_4390);
xor U5013 (N_5013,N_3711,N_3608);
and U5014 (N_5014,N_4501,N_4314);
or U5015 (N_5015,N_4690,N_3925);
xnor U5016 (N_5016,N_3884,N_3899);
nor U5017 (N_5017,N_4625,N_4221);
or U5018 (N_5018,N_4675,N_4433);
and U5019 (N_5019,N_4752,N_3918);
xnor U5020 (N_5020,N_4235,N_4537);
nor U5021 (N_5021,N_4512,N_3727);
or U5022 (N_5022,N_4017,N_3617);
nor U5023 (N_5023,N_4006,N_4289);
or U5024 (N_5024,N_3774,N_4130);
or U5025 (N_5025,N_4582,N_4131);
nand U5026 (N_5026,N_4161,N_3848);
nand U5027 (N_5027,N_3696,N_3936);
nand U5028 (N_5028,N_3980,N_4291);
xor U5029 (N_5029,N_4060,N_4602);
nor U5030 (N_5030,N_3828,N_4346);
and U5031 (N_5031,N_4739,N_4378);
nor U5032 (N_5032,N_3878,N_4312);
xor U5033 (N_5033,N_3748,N_4591);
nand U5034 (N_5034,N_4080,N_4187);
or U5035 (N_5035,N_3628,N_4404);
and U5036 (N_5036,N_3835,N_4728);
nor U5037 (N_5037,N_3839,N_3824);
xor U5038 (N_5038,N_4703,N_3759);
or U5039 (N_5039,N_4166,N_4071);
or U5040 (N_5040,N_4078,N_4388);
nand U5041 (N_5041,N_4514,N_4475);
and U5042 (N_5042,N_4382,N_3672);
and U5043 (N_5043,N_4292,N_4083);
or U5044 (N_5044,N_3725,N_4028);
and U5045 (N_5045,N_4186,N_4369);
nand U5046 (N_5046,N_3675,N_3786);
or U5047 (N_5047,N_3854,N_4447);
nand U5048 (N_5048,N_4546,N_4227);
or U5049 (N_5049,N_4048,N_3971);
xor U5050 (N_5050,N_3966,N_3620);
or U5051 (N_5051,N_4061,N_4668);
nand U5052 (N_5052,N_3965,N_4120);
and U5053 (N_5053,N_4473,N_4260);
nor U5054 (N_5054,N_4632,N_4642);
and U5055 (N_5055,N_4082,N_4139);
or U5056 (N_5056,N_3895,N_4778);
or U5057 (N_5057,N_4764,N_4029);
nor U5058 (N_5058,N_4639,N_4417);
and U5059 (N_5059,N_4527,N_4755);
nor U5060 (N_5060,N_3763,N_4484);
nor U5061 (N_5061,N_4385,N_4246);
nor U5062 (N_5062,N_4245,N_4180);
or U5063 (N_5063,N_4434,N_4151);
xnor U5064 (N_5064,N_4033,N_4003);
nand U5065 (N_5065,N_4571,N_3813);
xnor U5066 (N_5066,N_4347,N_4142);
xnor U5067 (N_5067,N_4256,N_3645);
nor U5068 (N_5068,N_4062,N_4742);
nor U5069 (N_5069,N_3651,N_4772);
xnor U5070 (N_5070,N_3709,N_4740);
and U5071 (N_5071,N_3938,N_4425);
nand U5072 (N_5072,N_4219,N_4557);
and U5073 (N_5073,N_4266,N_3837);
xor U5074 (N_5074,N_4074,N_4146);
xnor U5075 (N_5075,N_4365,N_4284);
and U5076 (N_5076,N_4646,N_3616);
nor U5077 (N_5077,N_4182,N_3735);
nand U5078 (N_5078,N_4562,N_3791);
nor U5079 (N_5079,N_4580,N_3793);
or U5080 (N_5080,N_3905,N_4328);
or U5081 (N_5081,N_3610,N_3643);
xor U5082 (N_5082,N_3742,N_4317);
nor U5083 (N_5083,N_4183,N_4217);
nor U5084 (N_5084,N_4086,N_3631);
and U5085 (N_5085,N_4437,N_4406);
nand U5086 (N_5086,N_4282,N_4617);
and U5087 (N_5087,N_4627,N_4600);
and U5088 (N_5088,N_4785,N_3998);
nor U5089 (N_5089,N_4398,N_4628);
and U5090 (N_5090,N_4239,N_4472);
or U5091 (N_5091,N_4419,N_3780);
or U5092 (N_5092,N_4767,N_4526);
nand U5093 (N_5093,N_4529,N_4377);
and U5094 (N_5094,N_4669,N_4325);
xnor U5095 (N_5095,N_4014,N_3771);
nor U5096 (N_5096,N_4405,N_3758);
xor U5097 (N_5097,N_4295,N_4231);
nor U5098 (N_5098,N_3996,N_3747);
nand U5099 (N_5099,N_3701,N_4634);
xnor U5100 (N_5100,N_3789,N_4296);
or U5101 (N_5101,N_4528,N_4233);
nand U5102 (N_5102,N_4477,N_4223);
nand U5103 (N_5103,N_4159,N_4392);
xnor U5104 (N_5104,N_4508,N_4597);
and U5105 (N_5105,N_4110,N_3986);
and U5106 (N_5106,N_4534,N_3941);
nand U5107 (N_5107,N_3819,N_4283);
nand U5108 (N_5108,N_4587,N_4494);
nand U5109 (N_5109,N_4303,N_3784);
and U5110 (N_5110,N_3800,N_3691);
and U5111 (N_5111,N_4340,N_3602);
nand U5112 (N_5112,N_3601,N_4367);
and U5113 (N_5113,N_4674,N_4424);
xnor U5114 (N_5114,N_4079,N_4502);
xnor U5115 (N_5115,N_3910,N_3777);
or U5116 (N_5116,N_3840,N_3957);
nand U5117 (N_5117,N_3681,N_4643);
nor U5118 (N_5118,N_4242,N_4089);
nor U5119 (N_5119,N_4660,N_3841);
nor U5120 (N_5120,N_4178,N_4748);
nand U5121 (N_5121,N_4462,N_3842);
nand U5122 (N_5122,N_4795,N_3847);
and U5123 (N_5123,N_3901,N_3794);
nor U5124 (N_5124,N_4630,N_4022);
or U5125 (N_5125,N_4016,N_4234);
and U5126 (N_5126,N_4049,N_3923);
xor U5127 (N_5127,N_4076,N_4732);
xnor U5128 (N_5128,N_3942,N_4545);
nor U5129 (N_5129,N_4206,N_4698);
xnor U5130 (N_5130,N_4466,N_4067);
nor U5131 (N_5131,N_3916,N_4504);
or U5132 (N_5132,N_4476,N_3817);
nand U5133 (N_5133,N_4185,N_3804);
and U5134 (N_5134,N_4254,N_4616);
nor U5135 (N_5135,N_4679,N_4412);
nor U5136 (N_5136,N_3846,N_4513);
xor U5137 (N_5137,N_4253,N_4197);
or U5138 (N_5138,N_4267,N_3827);
and U5139 (N_5139,N_4633,N_4177);
nand U5140 (N_5140,N_4336,N_3924);
or U5141 (N_5141,N_4561,N_3959);
or U5142 (N_5142,N_4455,N_3927);
and U5143 (N_5143,N_3797,N_4584);
xor U5144 (N_5144,N_4274,N_4426);
xor U5145 (N_5145,N_3871,N_3622);
nand U5146 (N_5146,N_4787,N_3783);
nand U5147 (N_5147,N_3728,N_4747);
or U5148 (N_5148,N_4556,N_3768);
nor U5149 (N_5149,N_4281,N_4650);
nor U5150 (N_5150,N_3716,N_4551);
xor U5151 (N_5151,N_3605,N_4018);
nand U5152 (N_5152,N_4608,N_4054);
or U5153 (N_5153,N_3638,N_3743);
or U5154 (N_5154,N_4104,N_4655);
or U5155 (N_5155,N_3974,N_3714);
nand U5156 (N_5156,N_4688,N_4542);
xor U5157 (N_5157,N_4109,N_4339);
nor U5158 (N_5158,N_4532,N_4680);
nand U5159 (N_5159,N_4158,N_3659);
xor U5160 (N_5160,N_3873,N_3781);
or U5161 (N_5161,N_4338,N_4479);
or U5162 (N_5162,N_3708,N_3937);
nor U5163 (N_5163,N_3897,N_4263);
nand U5164 (N_5164,N_3740,N_4019);
and U5165 (N_5165,N_4383,N_4273);
and U5166 (N_5166,N_4175,N_3893);
xor U5167 (N_5167,N_4699,N_4052);
and U5168 (N_5168,N_3678,N_4692);
xnor U5169 (N_5169,N_3703,N_4129);
nand U5170 (N_5170,N_3639,N_3650);
nor U5171 (N_5171,N_4754,N_3738);
nor U5172 (N_5172,N_4135,N_4757);
nand U5173 (N_5173,N_4096,N_3913);
nor U5174 (N_5174,N_4554,N_4157);
xnor U5175 (N_5175,N_4106,N_4162);
xnor U5176 (N_5176,N_3684,N_3820);
or U5177 (N_5177,N_4145,N_4064);
xnor U5178 (N_5178,N_4058,N_4560);
xnor U5179 (N_5179,N_3719,N_4783);
nand U5180 (N_5180,N_4498,N_4088);
or U5181 (N_5181,N_4490,N_4343);
and U5182 (N_5182,N_4331,N_4240);
or U5183 (N_5183,N_4421,N_4523);
nand U5184 (N_5184,N_4344,N_4621);
xnor U5185 (N_5185,N_4357,N_4786);
or U5186 (N_5186,N_4375,N_4765);
nor U5187 (N_5187,N_4348,N_4350);
and U5188 (N_5188,N_3752,N_4122);
and U5189 (N_5189,N_4320,N_3932);
or U5190 (N_5190,N_4030,N_4000);
nor U5191 (N_5191,N_4173,N_4684);
or U5192 (N_5192,N_4176,N_4598);
or U5193 (N_5193,N_4393,N_3656);
or U5194 (N_5194,N_4506,N_4037);
nand U5195 (N_5195,N_3978,N_4036);
nand U5196 (N_5196,N_4411,N_4521);
or U5197 (N_5197,N_3843,N_4202);
nand U5198 (N_5198,N_4613,N_3997);
nand U5199 (N_5199,N_3995,N_3663);
and U5200 (N_5200,N_3686,N_4662);
nor U5201 (N_5201,N_4652,N_3993);
or U5202 (N_5202,N_4536,N_3654);
nand U5203 (N_5203,N_4487,N_4056);
or U5204 (N_5204,N_4351,N_4683);
and U5205 (N_5205,N_4362,N_4496);
nand U5206 (N_5206,N_4066,N_3830);
xor U5207 (N_5207,N_4734,N_3808);
and U5208 (N_5208,N_4645,N_4128);
nor U5209 (N_5209,N_3977,N_3756);
nor U5210 (N_5210,N_3761,N_4168);
xnor U5211 (N_5211,N_4210,N_4741);
or U5212 (N_5212,N_3626,N_4196);
or U5213 (N_5213,N_4027,N_3688);
nor U5214 (N_5214,N_4517,N_4191);
and U5215 (N_5215,N_3867,N_3861);
or U5216 (N_5216,N_3850,N_4345);
nand U5217 (N_5217,N_4737,N_4002);
nor U5218 (N_5218,N_4644,N_4420);
xor U5219 (N_5219,N_3816,N_3929);
nand U5220 (N_5220,N_3722,N_4134);
nand U5221 (N_5221,N_3999,N_3700);
nand U5222 (N_5222,N_4797,N_3648);
nor U5223 (N_5223,N_4358,N_4293);
nor U5224 (N_5224,N_3745,N_4038);
nor U5225 (N_5225,N_3911,N_3883);
nand U5226 (N_5226,N_4103,N_4402);
nor U5227 (N_5227,N_3685,N_4794);
xor U5228 (N_5228,N_4559,N_4118);
nand U5229 (N_5229,N_4126,N_3954);
nand U5230 (N_5230,N_4269,N_4215);
nor U5231 (N_5231,N_4205,N_3744);
xor U5232 (N_5232,N_3900,N_4714);
or U5233 (N_5233,N_4380,N_4719);
xor U5234 (N_5234,N_4170,N_4533);
or U5235 (N_5235,N_3933,N_4341);
xor U5236 (N_5236,N_3687,N_4264);
and U5237 (N_5237,N_4276,N_4576);
xor U5238 (N_5238,N_4013,N_4558);
nand U5239 (N_5239,N_4252,N_4099);
xor U5240 (N_5240,N_3875,N_4138);
xor U5241 (N_5241,N_4793,N_3746);
and U5242 (N_5242,N_4045,N_3641);
xnor U5243 (N_5243,N_3609,N_4111);
and U5244 (N_5244,N_3866,N_3788);
or U5245 (N_5245,N_4717,N_3857);
nand U5246 (N_5246,N_4199,N_3621);
and U5247 (N_5247,N_4372,N_3787);
or U5248 (N_5248,N_4460,N_4213);
and U5249 (N_5249,N_4647,N_4631);
xor U5250 (N_5250,N_4366,N_4450);
xor U5251 (N_5251,N_4091,N_4009);
xnor U5252 (N_5252,N_4784,N_4194);
nor U5253 (N_5253,N_4208,N_4323);
xnor U5254 (N_5254,N_4456,N_4174);
nor U5255 (N_5255,N_4121,N_4298);
or U5256 (N_5256,N_4108,N_4776);
nand U5257 (N_5257,N_4488,N_4068);
and U5258 (N_5258,N_3931,N_4451);
nand U5259 (N_5259,N_4039,N_3706);
or U5260 (N_5260,N_4799,N_4127);
nor U5261 (N_5261,N_3733,N_3877);
nor U5262 (N_5262,N_3930,N_3917);
nand U5263 (N_5263,N_4649,N_4250);
and U5264 (N_5264,N_3894,N_4724);
or U5265 (N_5265,N_4745,N_4125);
nand U5266 (N_5266,N_3683,N_3889);
nand U5267 (N_5267,N_4050,N_4709);
nand U5268 (N_5268,N_4574,N_3882);
or U5269 (N_5269,N_3814,N_4132);
or U5270 (N_5270,N_3983,N_4026);
nor U5271 (N_5271,N_4400,N_4716);
and U5272 (N_5272,N_4520,N_4687);
or U5273 (N_5273,N_4519,N_3831);
nand U5274 (N_5274,N_4418,N_3868);
xnor U5275 (N_5275,N_4781,N_3948);
nand U5276 (N_5276,N_4638,N_4241);
nor U5277 (N_5277,N_4495,N_4588);
xor U5278 (N_5278,N_4311,N_3803);
xor U5279 (N_5279,N_3689,N_4119);
or U5280 (N_5280,N_4114,N_4541);
nand U5281 (N_5281,N_4577,N_4216);
or U5282 (N_5282,N_4516,N_4203);
nand U5283 (N_5283,N_4549,N_4623);
or U5284 (N_5284,N_4105,N_3627);
nand U5285 (N_5285,N_3657,N_4288);
nand U5286 (N_5286,N_4579,N_4763);
and U5287 (N_5287,N_4543,N_4771);
xnor U5288 (N_5288,N_3640,N_4606);
nor U5289 (N_5289,N_3970,N_4359);
nor U5290 (N_5290,N_4324,N_4313);
or U5291 (N_5291,N_4069,N_3860);
xnor U5292 (N_5292,N_4144,N_4791);
nor U5293 (N_5293,N_4440,N_4604);
nand U5294 (N_5294,N_4107,N_4123);
or U5295 (N_5295,N_4702,N_3796);
and U5296 (N_5296,N_3988,N_4651);
and U5297 (N_5297,N_4268,N_4285);
nand U5298 (N_5298,N_4770,N_4611);
xnor U5299 (N_5299,N_3697,N_4671);
nor U5300 (N_5300,N_4738,N_4670);
or U5301 (N_5301,N_4566,N_4636);
xnor U5302 (N_5302,N_4715,N_4084);
xor U5303 (N_5303,N_4373,N_3826);
and U5304 (N_5304,N_4010,N_4509);
xnor U5305 (N_5305,N_4444,N_4713);
xor U5306 (N_5306,N_3612,N_4322);
or U5307 (N_5307,N_4275,N_3898);
and U5308 (N_5308,N_3801,N_4736);
nand U5309 (N_5309,N_4749,N_3961);
xnor U5310 (N_5310,N_4271,N_4261);
nor U5311 (N_5311,N_4441,N_3766);
nor U5312 (N_5312,N_4470,N_3770);
or U5313 (N_5313,N_4389,N_4209);
xnor U5314 (N_5314,N_3862,N_3953);
nor U5315 (N_5315,N_4115,N_3832);
nor U5316 (N_5316,N_3666,N_4229);
or U5317 (N_5317,N_4154,N_3674);
xor U5318 (N_5318,N_3778,N_3858);
or U5319 (N_5319,N_4720,N_4790);
nand U5320 (N_5320,N_3690,N_3724);
and U5321 (N_5321,N_3955,N_4565);
or U5322 (N_5322,N_4428,N_3928);
and U5323 (N_5323,N_3734,N_4251);
xor U5324 (N_5324,N_3668,N_4309);
and U5325 (N_5325,N_3660,N_4788);
and U5326 (N_5326,N_3903,N_3606);
nor U5327 (N_5327,N_4524,N_3634);
xor U5328 (N_5328,N_3855,N_4485);
and U5329 (N_5329,N_4280,N_4779);
and U5330 (N_5330,N_3655,N_3945);
or U5331 (N_5331,N_4539,N_4678);
and U5332 (N_5332,N_3973,N_3775);
and U5333 (N_5333,N_3661,N_4503);
and U5334 (N_5334,N_4399,N_4493);
and U5335 (N_5335,N_4098,N_3717);
xnor U5336 (N_5336,N_4302,N_3698);
nor U5337 (N_5337,N_4629,N_4228);
and U5338 (N_5338,N_4244,N_3879);
xor U5339 (N_5339,N_4603,N_4243);
or U5340 (N_5340,N_4568,N_4165);
xnor U5341 (N_5341,N_4452,N_4059);
xnor U5342 (N_5342,N_4342,N_4401);
xor U5343 (N_5343,N_3720,N_4661);
and U5344 (N_5344,N_3765,N_4410);
nor U5345 (N_5345,N_4756,N_3964);
xnor U5346 (N_5346,N_4200,N_4766);
nand U5347 (N_5347,N_4593,N_3739);
or U5348 (N_5348,N_4583,N_3600);
nor U5349 (N_5349,N_3887,N_4007);
or U5350 (N_5350,N_4218,N_3825);
xor U5351 (N_5351,N_4224,N_4700);
or U5352 (N_5352,N_4775,N_3951);
or U5353 (N_5353,N_3958,N_4798);
nor U5354 (N_5354,N_3912,N_4337);
nand U5355 (N_5355,N_4226,N_4550);
or U5356 (N_5356,N_4387,N_4167);
or U5357 (N_5357,N_4113,N_4682);
or U5358 (N_5358,N_3669,N_4101);
and U5359 (N_5359,N_4654,N_4184);
or U5360 (N_5360,N_4070,N_4612);
nand U5361 (N_5361,N_4759,N_4712);
nor U5362 (N_5362,N_3699,N_4287);
or U5363 (N_5363,N_3667,N_4666);
nand U5364 (N_5364,N_4306,N_4043);
nor U5365 (N_5365,N_4435,N_3799);
or U5366 (N_5366,N_3872,N_4143);
and U5367 (N_5367,N_4701,N_4356);
and U5368 (N_5368,N_4750,N_4430);
and U5369 (N_5369,N_4648,N_4371);
nand U5370 (N_5370,N_4077,N_4704);
and U5371 (N_5371,N_3865,N_3633);
nand U5372 (N_5372,N_4590,N_4172);
nand U5373 (N_5373,N_4112,N_4087);
xor U5374 (N_5374,N_3623,N_3876);
nor U5375 (N_5375,N_3751,N_3863);
xnor U5376 (N_5376,N_3934,N_3920);
and U5377 (N_5377,N_4471,N_4482);
nand U5378 (N_5378,N_3982,N_4012);
nand U5379 (N_5379,N_4169,N_4225);
and U5380 (N_5380,N_3680,N_4445);
nand U5381 (N_5381,N_4095,N_3737);
xor U5382 (N_5382,N_4535,N_4294);
and U5383 (N_5383,N_3821,N_4431);
xnor U5384 (N_5384,N_4721,N_3624);
nor U5385 (N_5385,N_4257,N_4352);
nor U5386 (N_5386,N_4592,N_3671);
or U5387 (N_5387,N_4149,N_4092);
nand U5388 (N_5388,N_3676,N_4436);
xnor U5389 (N_5389,N_4327,N_4133);
and U5390 (N_5390,N_3869,N_4596);
or U5391 (N_5391,N_4355,N_4626);
xnor U5392 (N_5392,N_3632,N_3647);
nor U5393 (N_5393,N_4711,N_3754);
xnor U5394 (N_5394,N_3670,N_4443);
and U5395 (N_5395,N_3981,N_4665);
nor U5396 (N_5396,N_3853,N_4507);
nor U5397 (N_5397,N_4259,N_4044);
nand U5398 (N_5398,N_4316,N_4031);
and U5399 (N_5399,N_3963,N_4511);
xnor U5400 (N_5400,N_3977,N_3625);
xor U5401 (N_5401,N_4023,N_3775);
xor U5402 (N_5402,N_4578,N_3756);
xor U5403 (N_5403,N_4261,N_3614);
or U5404 (N_5404,N_3623,N_4756);
and U5405 (N_5405,N_3867,N_4648);
or U5406 (N_5406,N_4684,N_4591);
and U5407 (N_5407,N_4399,N_4172);
or U5408 (N_5408,N_3690,N_4026);
xor U5409 (N_5409,N_4372,N_4041);
nor U5410 (N_5410,N_4330,N_4484);
nor U5411 (N_5411,N_4520,N_3658);
or U5412 (N_5412,N_4554,N_4111);
nand U5413 (N_5413,N_4509,N_4343);
nor U5414 (N_5414,N_4491,N_4200);
nor U5415 (N_5415,N_4080,N_3919);
xor U5416 (N_5416,N_4574,N_3900);
or U5417 (N_5417,N_3850,N_4052);
or U5418 (N_5418,N_4794,N_3866);
and U5419 (N_5419,N_3753,N_3695);
and U5420 (N_5420,N_4601,N_4006);
and U5421 (N_5421,N_4411,N_3876);
or U5422 (N_5422,N_4773,N_3671);
or U5423 (N_5423,N_4364,N_4320);
nand U5424 (N_5424,N_4763,N_4317);
nand U5425 (N_5425,N_4231,N_4720);
nand U5426 (N_5426,N_4170,N_3644);
and U5427 (N_5427,N_4060,N_4600);
and U5428 (N_5428,N_3862,N_4739);
xnor U5429 (N_5429,N_4780,N_3752);
nand U5430 (N_5430,N_4715,N_4409);
and U5431 (N_5431,N_3699,N_4700);
nor U5432 (N_5432,N_4210,N_3790);
or U5433 (N_5433,N_4131,N_4721);
nor U5434 (N_5434,N_3974,N_3644);
nor U5435 (N_5435,N_4512,N_4281);
nand U5436 (N_5436,N_4033,N_4069);
xnor U5437 (N_5437,N_3941,N_4638);
xnor U5438 (N_5438,N_4714,N_3801);
nand U5439 (N_5439,N_3865,N_3794);
nand U5440 (N_5440,N_4377,N_3992);
or U5441 (N_5441,N_4388,N_4433);
nand U5442 (N_5442,N_4573,N_4733);
and U5443 (N_5443,N_4611,N_3868);
nand U5444 (N_5444,N_3972,N_3789);
xnor U5445 (N_5445,N_4546,N_4780);
or U5446 (N_5446,N_4190,N_4498);
xnor U5447 (N_5447,N_4585,N_4779);
nor U5448 (N_5448,N_4044,N_4424);
nor U5449 (N_5449,N_4306,N_4480);
xnor U5450 (N_5450,N_3749,N_4530);
nor U5451 (N_5451,N_4525,N_4652);
nand U5452 (N_5452,N_3623,N_4451);
and U5453 (N_5453,N_4026,N_4070);
nand U5454 (N_5454,N_4278,N_4536);
and U5455 (N_5455,N_4325,N_3784);
nand U5456 (N_5456,N_4773,N_3751);
nor U5457 (N_5457,N_4001,N_4631);
nor U5458 (N_5458,N_4102,N_4379);
nor U5459 (N_5459,N_4155,N_4249);
or U5460 (N_5460,N_4736,N_4456);
nor U5461 (N_5461,N_4700,N_3696);
nor U5462 (N_5462,N_3996,N_4614);
and U5463 (N_5463,N_4547,N_4012);
or U5464 (N_5464,N_4384,N_4260);
xor U5465 (N_5465,N_4043,N_3994);
and U5466 (N_5466,N_3877,N_4258);
xor U5467 (N_5467,N_4479,N_3819);
or U5468 (N_5468,N_3896,N_4787);
nor U5469 (N_5469,N_4427,N_3654);
nor U5470 (N_5470,N_4678,N_4477);
xor U5471 (N_5471,N_3962,N_3979);
xnor U5472 (N_5472,N_3710,N_3721);
or U5473 (N_5473,N_3657,N_4436);
xor U5474 (N_5474,N_4719,N_3819);
nand U5475 (N_5475,N_3723,N_4002);
nor U5476 (N_5476,N_3785,N_4371);
nand U5477 (N_5477,N_4278,N_4405);
nor U5478 (N_5478,N_4606,N_3714);
xor U5479 (N_5479,N_4335,N_3750);
or U5480 (N_5480,N_4219,N_3685);
xor U5481 (N_5481,N_3862,N_3670);
xor U5482 (N_5482,N_3796,N_4191);
nor U5483 (N_5483,N_4519,N_4500);
or U5484 (N_5484,N_4252,N_4066);
and U5485 (N_5485,N_4245,N_3834);
nand U5486 (N_5486,N_3777,N_3951);
and U5487 (N_5487,N_4190,N_4625);
nand U5488 (N_5488,N_4672,N_4137);
nor U5489 (N_5489,N_4063,N_4563);
xnor U5490 (N_5490,N_4472,N_4309);
xor U5491 (N_5491,N_3605,N_3600);
nor U5492 (N_5492,N_4204,N_4442);
nand U5493 (N_5493,N_4158,N_4264);
nand U5494 (N_5494,N_4626,N_3737);
or U5495 (N_5495,N_3799,N_3893);
and U5496 (N_5496,N_4540,N_4311);
nor U5497 (N_5497,N_4127,N_3772);
or U5498 (N_5498,N_4008,N_3702);
nand U5499 (N_5499,N_4477,N_4755);
and U5500 (N_5500,N_4405,N_3766);
nor U5501 (N_5501,N_4474,N_4242);
or U5502 (N_5502,N_4621,N_3923);
nand U5503 (N_5503,N_4579,N_4750);
and U5504 (N_5504,N_3602,N_3956);
xnor U5505 (N_5505,N_4781,N_4566);
xnor U5506 (N_5506,N_3702,N_4656);
nand U5507 (N_5507,N_4577,N_4638);
and U5508 (N_5508,N_4387,N_4186);
nand U5509 (N_5509,N_3859,N_3780);
and U5510 (N_5510,N_4356,N_3672);
nor U5511 (N_5511,N_4365,N_4229);
nand U5512 (N_5512,N_4585,N_4055);
nand U5513 (N_5513,N_3778,N_4200);
nand U5514 (N_5514,N_4250,N_4572);
and U5515 (N_5515,N_4315,N_4753);
xnor U5516 (N_5516,N_4306,N_4596);
or U5517 (N_5517,N_4123,N_4016);
or U5518 (N_5518,N_4300,N_3861);
and U5519 (N_5519,N_4582,N_4259);
and U5520 (N_5520,N_4359,N_3853);
or U5521 (N_5521,N_3924,N_4492);
nand U5522 (N_5522,N_4615,N_4200);
or U5523 (N_5523,N_4141,N_4347);
and U5524 (N_5524,N_4422,N_4247);
nand U5525 (N_5525,N_4053,N_4571);
nor U5526 (N_5526,N_3848,N_4098);
xnor U5527 (N_5527,N_3777,N_3998);
xnor U5528 (N_5528,N_4560,N_4625);
nand U5529 (N_5529,N_4261,N_3797);
nand U5530 (N_5530,N_3922,N_4446);
or U5531 (N_5531,N_4272,N_4685);
xnor U5532 (N_5532,N_4194,N_4282);
and U5533 (N_5533,N_4710,N_4294);
nand U5534 (N_5534,N_4125,N_3650);
xnor U5535 (N_5535,N_4658,N_4797);
nand U5536 (N_5536,N_3640,N_3610);
or U5537 (N_5537,N_3977,N_4042);
and U5538 (N_5538,N_4506,N_4770);
or U5539 (N_5539,N_3624,N_4032);
and U5540 (N_5540,N_4062,N_3682);
xor U5541 (N_5541,N_3846,N_4434);
xnor U5542 (N_5542,N_4797,N_4237);
nand U5543 (N_5543,N_4243,N_4445);
and U5544 (N_5544,N_3840,N_4389);
nor U5545 (N_5545,N_4275,N_4796);
nand U5546 (N_5546,N_4174,N_4680);
and U5547 (N_5547,N_4718,N_4108);
or U5548 (N_5548,N_3944,N_4252);
and U5549 (N_5549,N_4180,N_4260);
xnor U5550 (N_5550,N_4372,N_4049);
and U5551 (N_5551,N_4732,N_4559);
or U5552 (N_5552,N_4106,N_3893);
xnor U5553 (N_5553,N_4024,N_4115);
nand U5554 (N_5554,N_4762,N_3786);
nand U5555 (N_5555,N_4208,N_3820);
nor U5556 (N_5556,N_4419,N_4505);
nor U5557 (N_5557,N_4051,N_4595);
and U5558 (N_5558,N_4180,N_3885);
and U5559 (N_5559,N_3969,N_4136);
and U5560 (N_5560,N_3818,N_4576);
nor U5561 (N_5561,N_4612,N_4336);
or U5562 (N_5562,N_4080,N_4777);
nor U5563 (N_5563,N_4505,N_3957);
xnor U5564 (N_5564,N_4493,N_4387);
and U5565 (N_5565,N_4779,N_3970);
xnor U5566 (N_5566,N_4173,N_3681);
or U5567 (N_5567,N_3798,N_4061);
nand U5568 (N_5568,N_3814,N_4514);
nor U5569 (N_5569,N_3703,N_4061);
xor U5570 (N_5570,N_4419,N_4405);
or U5571 (N_5571,N_3974,N_4770);
nor U5572 (N_5572,N_4305,N_3738);
nor U5573 (N_5573,N_3797,N_4248);
or U5574 (N_5574,N_4599,N_4071);
xor U5575 (N_5575,N_3905,N_3720);
xor U5576 (N_5576,N_4077,N_3986);
xnor U5577 (N_5577,N_4291,N_4432);
nor U5578 (N_5578,N_4111,N_4184);
nand U5579 (N_5579,N_4666,N_4702);
or U5580 (N_5580,N_4318,N_3869);
nor U5581 (N_5581,N_4311,N_4533);
nor U5582 (N_5582,N_4604,N_4041);
and U5583 (N_5583,N_4628,N_3878);
nand U5584 (N_5584,N_3784,N_4528);
xor U5585 (N_5585,N_4397,N_3865);
nand U5586 (N_5586,N_4096,N_4569);
nand U5587 (N_5587,N_4433,N_3653);
xnor U5588 (N_5588,N_4446,N_4777);
or U5589 (N_5589,N_4122,N_3807);
nand U5590 (N_5590,N_4516,N_4594);
xor U5591 (N_5591,N_3839,N_4366);
and U5592 (N_5592,N_4205,N_3715);
or U5593 (N_5593,N_3820,N_4762);
and U5594 (N_5594,N_4162,N_3895);
and U5595 (N_5595,N_4673,N_4534);
and U5596 (N_5596,N_3698,N_4746);
nor U5597 (N_5597,N_4624,N_4768);
and U5598 (N_5598,N_3994,N_3758);
nand U5599 (N_5599,N_4146,N_4758);
xor U5600 (N_5600,N_4355,N_4225);
nor U5601 (N_5601,N_4740,N_4471);
or U5602 (N_5602,N_4156,N_4682);
or U5603 (N_5603,N_4612,N_4112);
or U5604 (N_5604,N_4500,N_4175);
nand U5605 (N_5605,N_4781,N_4581);
xnor U5606 (N_5606,N_4799,N_4374);
nand U5607 (N_5607,N_4433,N_4141);
nor U5608 (N_5608,N_3799,N_4779);
or U5609 (N_5609,N_4301,N_4391);
xnor U5610 (N_5610,N_4438,N_4439);
or U5611 (N_5611,N_4651,N_4392);
nor U5612 (N_5612,N_3660,N_4798);
nor U5613 (N_5613,N_3634,N_4282);
xor U5614 (N_5614,N_4546,N_4152);
nor U5615 (N_5615,N_4411,N_4468);
xor U5616 (N_5616,N_3700,N_4040);
xor U5617 (N_5617,N_4302,N_3761);
nand U5618 (N_5618,N_4590,N_4198);
nand U5619 (N_5619,N_3936,N_4456);
xnor U5620 (N_5620,N_3740,N_4234);
nor U5621 (N_5621,N_3740,N_4231);
nand U5622 (N_5622,N_3739,N_4035);
or U5623 (N_5623,N_4476,N_4427);
and U5624 (N_5624,N_4436,N_3601);
xor U5625 (N_5625,N_4496,N_3867);
nor U5626 (N_5626,N_4205,N_4741);
or U5627 (N_5627,N_4758,N_4236);
and U5628 (N_5628,N_4005,N_4064);
or U5629 (N_5629,N_4405,N_3995);
nor U5630 (N_5630,N_4163,N_3723);
and U5631 (N_5631,N_4057,N_3613);
nor U5632 (N_5632,N_4023,N_4420);
and U5633 (N_5633,N_4033,N_4039);
or U5634 (N_5634,N_3822,N_3777);
and U5635 (N_5635,N_4234,N_4668);
nor U5636 (N_5636,N_4761,N_4300);
xnor U5637 (N_5637,N_4470,N_4740);
nor U5638 (N_5638,N_3747,N_4519);
nand U5639 (N_5639,N_3975,N_4506);
or U5640 (N_5640,N_4278,N_4127);
and U5641 (N_5641,N_4276,N_4748);
nor U5642 (N_5642,N_3675,N_4157);
nor U5643 (N_5643,N_4166,N_4167);
xnor U5644 (N_5644,N_4248,N_4447);
or U5645 (N_5645,N_3704,N_4282);
nor U5646 (N_5646,N_3754,N_4547);
xnor U5647 (N_5647,N_3852,N_3984);
and U5648 (N_5648,N_3923,N_4704);
nand U5649 (N_5649,N_3861,N_4234);
or U5650 (N_5650,N_4076,N_4736);
nand U5651 (N_5651,N_4578,N_4090);
nor U5652 (N_5652,N_4323,N_3790);
xor U5653 (N_5653,N_4788,N_3665);
or U5654 (N_5654,N_4007,N_4315);
and U5655 (N_5655,N_4306,N_4589);
or U5656 (N_5656,N_4330,N_3674);
xor U5657 (N_5657,N_4798,N_4643);
xor U5658 (N_5658,N_4301,N_3933);
and U5659 (N_5659,N_3648,N_3807);
nand U5660 (N_5660,N_3756,N_4131);
xnor U5661 (N_5661,N_4056,N_4009);
xor U5662 (N_5662,N_4189,N_4654);
nand U5663 (N_5663,N_4510,N_4260);
nor U5664 (N_5664,N_4114,N_4356);
or U5665 (N_5665,N_3787,N_3972);
or U5666 (N_5666,N_4085,N_3604);
nor U5667 (N_5667,N_4761,N_4137);
xor U5668 (N_5668,N_3855,N_4015);
or U5669 (N_5669,N_3949,N_4533);
or U5670 (N_5670,N_4726,N_3906);
nand U5671 (N_5671,N_4274,N_3634);
nor U5672 (N_5672,N_3650,N_4644);
xnor U5673 (N_5673,N_3880,N_4606);
nand U5674 (N_5674,N_4732,N_4286);
and U5675 (N_5675,N_4196,N_4104);
and U5676 (N_5676,N_3864,N_4303);
and U5677 (N_5677,N_4140,N_4424);
or U5678 (N_5678,N_4239,N_3828);
nand U5679 (N_5679,N_4301,N_4516);
or U5680 (N_5680,N_4642,N_4578);
and U5681 (N_5681,N_4179,N_4356);
or U5682 (N_5682,N_3766,N_4414);
nor U5683 (N_5683,N_3863,N_4395);
or U5684 (N_5684,N_3946,N_3897);
and U5685 (N_5685,N_3961,N_3770);
nor U5686 (N_5686,N_4251,N_4315);
or U5687 (N_5687,N_3798,N_3710);
nand U5688 (N_5688,N_3798,N_3695);
or U5689 (N_5689,N_4111,N_4752);
nor U5690 (N_5690,N_3937,N_4365);
or U5691 (N_5691,N_4231,N_4449);
nor U5692 (N_5692,N_3834,N_3925);
nand U5693 (N_5693,N_3723,N_4024);
nand U5694 (N_5694,N_4149,N_4011);
xor U5695 (N_5695,N_4701,N_4073);
nand U5696 (N_5696,N_3748,N_4552);
or U5697 (N_5697,N_4539,N_4052);
or U5698 (N_5698,N_4101,N_3920);
xor U5699 (N_5699,N_4122,N_4645);
nor U5700 (N_5700,N_3752,N_4510);
nor U5701 (N_5701,N_4428,N_4321);
nand U5702 (N_5702,N_4027,N_4166);
or U5703 (N_5703,N_4661,N_4552);
nor U5704 (N_5704,N_4331,N_3803);
nor U5705 (N_5705,N_4372,N_4127);
xor U5706 (N_5706,N_4144,N_4440);
nor U5707 (N_5707,N_3951,N_4592);
xnor U5708 (N_5708,N_4153,N_4093);
and U5709 (N_5709,N_3804,N_3749);
and U5710 (N_5710,N_4226,N_4148);
nor U5711 (N_5711,N_3808,N_4640);
and U5712 (N_5712,N_3847,N_4199);
or U5713 (N_5713,N_4538,N_4214);
nand U5714 (N_5714,N_4277,N_3765);
and U5715 (N_5715,N_3664,N_4043);
nand U5716 (N_5716,N_3936,N_4716);
or U5717 (N_5717,N_4516,N_4152);
or U5718 (N_5718,N_4444,N_4331);
and U5719 (N_5719,N_3878,N_3830);
or U5720 (N_5720,N_3646,N_4307);
or U5721 (N_5721,N_4079,N_4683);
nand U5722 (N_5722,N_3851,N_3636);
and U5723 (N_5723,N_3865,N_4199);
xnor U5724 (N_5724,N_4634,N_4718);
and U5725 (N_5725,N_4446,N_4718);
nor U5726 (N_5726,N_3864,N_3813);
and U5727 (N_5727,N_4265,N_4314);
nand U5728 (N_5728,N_3905,N_4074);
nand U5729 (N_5729,N_4236,N_4374);
xnor U5730 (N_5730,N_4611,N_3919);
xnor U5731 (N_5731,N_3616,N_4619);
nand U5732 (N_5732,N_4009,N_4565);
and U5733 (N_5733,N_3618,N_4440);
nand U5734 (N_5734,N_3853,N_4065);
or U5735 (N_5735,N_4160,N_3873);
xnor U5736 (N_5736,N_4404,N_3818);
xor U5737 (N_5737,N_4777,N_4203);
xor U5738 (N_5738,N_4755,N_4730);
and U5739 (N_5739,N_3986,N_4490);
and U5740 (N_5740,N_3941,N_4038);
nor U5741 (N_5741,N_3728,N_3921);
nor U5742 (N_5742,N_4102,N_4349);
and U5743 (N_5743,N_4585,N_4393);
nand U5744 (N_5744,N_4137,N_4360);
nor U5745 (N_5745,N_3838,N_4755);
nand U5746 (N_5746,N_3746,N_4525);
xor U5747 (N_5747,N_4745,N_4064);
nor U5748 (N_5748,N_3920,N_3852);
or U5749 (N_5749,N_4138,N_4512);
and U5750 (N_5750,N_4049,N_3943);
nand U5751 (N_5751,N_4450,N_4672);
xor U5752 (N_5752,N_4058,N_4595);
nor U5753 (N_5753,N_3983,N_4080);
nand U5754 (N_5754,N_3737,N_3616);
or U5755 (N_5755,N_4045,N_4708);
or U5756 (N_5756,N_4128,N_4124);
xnor U5757 (N_5757,N_4364,N_4456);
nor U5758 (N_5758,N_4597,N_4624);
xor U5759 (N_5759,N_4417,N_3650);
or U5760 (N_5760,N_3886,N_4406);
xnor U5761 (N_5761,N_4323,N_4008);
and U5762 (N_5762,N_4134,N_4552);
xor U5763 (N_5763,N_3668,N_3946);
and U5764 (N_5764,N_4110,N_4283);
nand U5765 (N_5765,N_3647,N_3694);
and U5766 (N_5766,N_3765,N_4221);
and U5767 (N_5767,N_4350,N_3690);
nor U5768 (N_5768,N_4692,N_3835);
or U5769 (N_5769,N_3709,N_3884);
or U5770 (N_5770,N_4050,N_4481);
nor U5771 (N_5771,N_4040,N_4092);
nor U5772 (N_5772,N_3860,N_4001);
nand U5773 (N_5773,N_3824,N_4763);
nand U5774 (N_5774,N_4064,N_3796);
nor U5775 (N_5775,N_4438,N_4389);
xor U5776 (N_5776,N_3600,N_4337);
or U5777 (N_5777,N_3839,N_4541);
xnor U5778 (N_5778,N_4134,N_4021);
xor U5779 (N_5779,N_3892,N_4703);
xor U5780 (N_5780,N_4135,N_3903);
nor U5781 (N_5781,N_4133,N_3731);
xnor U5782 (N_5782,N_4410,N_4247);
and U5783 (N_5783,N_4413,N_4500);
and U5784 (N_5784,N_4397,N_4503);
nor U5785 (N_5785,N_4344,N_3994);
nand U5786 (N_5786,N_4072,N_4335);
and U5787 (N_5787,N_4205,N_3915);
xnor U5788 (N_5788,N_4494,N_3944);
or U5789 (N_5789,N_3921,N_3744);
or U5790 (N_5790,N_3735,N_4345);
xnor U5791 (N_5791,N_4476,N_4400);
or U5792 (N_5792,N_3847,N_3837);
and U5793 (N_5793,N_4464,N_4501);
and U5794 (N_5794,N_4650,N_3816);
and U5795 (N_5795,N_4770,N_3754);
or U5796 (N_5796,N_3940,N_4299);
and U5797 (N_5797,N_4416,N_3734);
and U5798 (N_5798,N_3671,N_4047);
nor U5799 (N_5799,N_3604,N_3848);
nand U5800 (N_5800,N_3718,N_4550);
nor U5801 (N_5801,N_4577,N_4306);
xor U5802 (N_5802,N_4699,N_3756);
nand U5803 (N_5803,N_4641,N_3603);
and U5804 (N_5804,N_4651,N_4342);
nand U5805 (N_5805,N_4733,N_4107);
or U5806 (N_5806,N_3886,N_4779);
or U5807 (N_5807,N_3834,N_3998);
or U5808 (N_5808,N_3692,N_3660);
nand U5809 (N_5809,N_4419,N_4720);
xor U5810 (N_5810,N_3888,N_4453);
xor U5811 (N_5811,N_4256,N_3876);
and U5812 (N_5812,N_4065,N_4782);
and U5813 (N_5813,N_3935,N_3984);
nor U5814 (N_5814,N_4547,N_3672);
and U5815 (N_5815,N_3904,N_3727);
nor U5816 (N_5816,N_4746,N_3697);
nor U5817 (N_5817,N_3875,N_4109);
xor U5818 (N_5818,N_4651,N_3718);
nand U5819 (N_5819,N_3761,N_3865);
xor U5820 (N_5820,N_4278,N_4351);
and U5821 (N_5821,N_3954,N_4422);
xor U5822 (N_5822,N_4648,N_3833);
or U5823 (N_5823,N_4133,N_3679);
or U5824 (N_5824,N_4033,N_3870);
nor U5825 (N_5825,N_4167,N_4796);
xor U5826 (N_5826,N_4486,N_4194);
xor U5827 (N_5827,N_3894,N_4234);
xor U5828 (N_5828,N_4630,N_3821);
and U5829 (N_5829,N_3783,N_4326);
nand U5830 (N_5830,N_4127,N_4229);
or U5831 (N_5831,N_4355,N_4285);
nor U5832 (N_5832,N_4056,N_3615);
or U5833 (N_5833,N_3921,N_4197);
and U5834 (N_5834,N_3897,N_4223);
nand U5835 (N_5835,N_4117,N_3973);
and U5836 (N_5836,N_4302,N_3924);
or U5837 (N_5837,N_3935,N_3885);
nor U5838 (N_5838,N_4757,N_4067);
nand U5839 (N_5839,N_4285,N_3711);
or U5840 (N_5840,N_4110,N_3708);
or U5841 (N_5841,N_4411,N_4430);
nand U5842 (N_5842,N_3828,N_4578);
and U5843 (N_5843,N_3778,N_4744);
nand U5844 (N_5844,N_4541,N_3966);
nand U5845 (N_5845,N_3732,N_4496);
xor U5846 (N_5846,N_3966,N_4731);
nor U5847 (N_5847,N_4024,N_4070);
and U5848 (N_5848,N_4156,N_4018);
or U5849 (N_5849,N_4331,N_4271);
nand U5850 (N_5850,N_3965,N_4702);
nor U5851 (N_5851,N_4640,N_4452);
nand U5852 (N_5852,N_4156,N_4385);
xnor U5853 (N_5853,N_4509,N_4709);
xnor U5854 (N_5854,N_4153,N_4475);
and U5855 (N_5855,N_4194,N_3997);
or U5856 (N_5856,N_3891,N_3931);
xnor U5857 (N_5857,N_4336,N_4287);
nor U5858 (N_5858,N_3853,N_3647);
or U5859 (N_5859,N_3817,N_4613);
and U5860 (N_5860,N_4422,N_4259);
and U5861 (N_5861,N_4484,N_4526);
or U5862 (N_5862,N_3725,N_3863);
nor U5863 (N_5863,N_4758,N_3814);
nor U5864 (N_5864,N_4009,N_4708);
or U5865 (N_5865,N_3703,N_4348);
nor U5866 (N_5866,N_4367,N_3821);
or U5867 (N_5867,N_4479,N_4376);
xnor U5868 (N_5868,N_4694,N_4074);
or U5869 (N_5869,N_4608,N_4116);
nor U5870 (N_5870,N_4633,N_4652);
nor U5871 (N_5871,N_4412,N_4483);
xnor U5872 (N_5872,N_4307,N_4137);
xor U5873 (N_5873,N_4798,N_4021);
nand U5874 (N_5874,N_4565,N_4287);
nor U5875 (N_5875,N_3860,N_4418);
nor U5876 (N_5876,N_4259,N_4000);
nand U5877 (N_5877,N_4130,N_3671);
and U5878 (N_5878,N_4011,N_4250);
or U5879 (N_5879,N_4406,N_4281);
nand U5880 (N_5880,N_4004,N_4283);
xor U5881 (N_5881,N_4429,N_4730);
nor U5882 (N_5882,N_4574,N_4003);
nand U5883 (N_5883,N_3803,N_4160);
nor U5884 (N_5884,N_4476,N_4224);
nand U5885 (N_5885,N_4279,N_4738);
or U5886 (N_5886,N_3906,N_3970);
and U5887 (N_5887,N_4607,N_4281);
xor U5888 (N_5888,N_4427,N_4765);
nor U5889 (N_5889,N_4770,N_4496);
or U5890 (N_5890,N_3926,N_4322);
and U5891 (N_5891,N_3706,N_4629);
or U5892 (N_5892,N_4130,N_3915);
and U5893 (N_5893,N_3949,N_3946);
or U5894 (N_5894,N_4647,N_3989);
xnor U5895 (N_5895,N_3888,N_4512);
and U5896 (N_5896,N_4072,N_4409);
nand U5897 (N_5897,N_4433,N_4523);
nor U5898 (N_5898,N_4193,N_4541);
nor U5899 (N_5899,N_4770,N_4245);
nor U5900 (N_5900,N_4350,N_3653);
nand U5901 (N_5901,N_3777,N_4707);
and U5902 (N_5902,N_4406,N_3983);
xor U5903 (N_5903,N_4242,N_4328);
and U5904 (N_5904,N_3883,N_4252);
nand U5905 (N_5905,N_3750,N_4003);
and U5906 (N_5906,N_4589,N_4450);
nand U5907 (N_5907,N_3995,N_3637);
or U5908 (N_5908,N_4037,N_3658);
and U5909 (N_5909,N_4635,N_4243);
or U5910 (N_5910,N_4758,N_3795);
nand U5911 (N_5911,N_4426,N_4042);
or U5912 (N_5912,N_4507,N_4125);
nand U5913 (N_5913,N_4229,N_4305);
xnor U5914 (N_5914,N_4611,N_3665);
or U5915 (N_5915,N_4304,N_4106);
xnor U5916 (N_5916,N_4467,N_3712);
and U5917 (N_5917,N_4760,N_4750);
nor U5918 (N_5918,N_3931,N_3682);
xnor U5919 (N_5919,N_4391,N_4492);
nor U5920 (N_5920,N_4021,N_3680);
nand U5921 (N_5921,N_4391,N_3708);
nor U5922 (N_5922,N_4145,N_4362);
and U5923 (N_5923,N_3656,N_4356);
or U5924 (N_5924,N_4766,N_4101);
or U5925 (N_5925,N_4737,N_3806);
and U5926 (N_5926,N_3884,N_4539);
xnor U5927 (N_5927,N_4334,N_4263);
xor U5928 (N_5928,N_3919,N_4779);
nand U5929 (N_5929,N_4344,N_4254);
and U5930 (N_5930,N_4278,N_4682);
nor U5931 (N_5931,N_4107,N_4469);
xnor U5932 (N_5932,N_4310,N_4696);
xnor U5933 (N_5933,N_4524,N_4566);
and U5934 (N_5934,N_3738,N_4640);
and U5935 (N_5935,N_4697,N_3855);
and U5936 (N_5936,N_4192,N_3624);
nor U5937 (N_5937,N_3652,N_4704);
xor U5938 (N_5938,N_3736,N_4753);
nor U5939 (N_5939,N_4529,N_4526);
or U5940 (N_5940,N_3820,N_3987);
nor U5941 (N_5941,N_3778,N_4473);
and U5942 (N_5942,N_4762,N_3733);
or U5943 (N_5943,N_3924,N_4462);
xor U5944 (N_5944,N_4378,N_4530);
or U5945 (N_5945,N_4002,N_3969);
or U5946 (N_5946,N_4157,N_3789);
nor U5947 (N_5947,N_4236,N_3764);
xor U5948 (N_5948,N_4647,N_3733);
xnor U5949 (N_5949,N_4067,N_4225);
or U5950 (N_5950,N_4119,N_4008);
nand U5951 (N_5951,N_4234,N_4306);
nor U5952 (N_5952,N_4622,N_4720);
and U5953 (N_5953,N_3705,N_4647);
and U5954 (N_5954,N_4146,N_4373);
and U5955 (N_5955,N_4088,N_3935);
and U5956 (N_5956,N_4302,N_3689);
and U5957 (N_5957,N_4762,N_4743);
nor U5958 (N_5958,N_4317,N_4270);
nor U5959 (N_5959,N_3673,N_4112);
or U5960 (N_5960,N_4528,N_3951);
nor U5961 (N_5961,N_3771,N_4795);
and U5962 (N_5962,N_3912,N_4641);
or U5963 (N_5963,N_3840,N_3754);
nor U5964 (N_5964,N_3871,N_4655);
or U5965 (N_5965,N_4411,N_4083);
or U5966 (N_5966,N_3748,N_4794);
nand U5967 (N_5967,N_4240,N_3994);
or U5968 (N_5968,N_3784,N_3914);
nor U5969 (N_5969,N_4067,N_3864);
nor U5970 (N_5970,N_4330,N_4544);
xnor U5971 (N_5971,N_4780,N_4387);
or U5972 (N_5972,N_4525,N_3777);
nand U5973 (N_5973,N_4155,N_4561);
nor U5974 (N_5974,N_3744,N_4321);
xnor U5975 (N_5975,N_4567,N_4458);
and U5976 (N_5976,N_4778,N_3724);
nor U5977 (N_5977,N_3785,N_4622);
nand U5978 (N_5978,N_3829,N_4754);
and U5979 (N_5979,N_4007,N_4509);
or U5980 (N_5980,N_3703,N_4501);
and U5981 (N_5981,N_3981,N_4180);
nor U5982 (N_5982,N_4365,N_3853);
nand U5983 (N_5983,N_4252,N_4488);
nor U5984 (N_5984,N_4767,N_4727);
nand U5985 (N_5985,N_3721,N_4020);
xor U5986 (N_5986,N_4515,N_4003);
and U5987 (N_5987,N_4223,N_4052);
xnor U5988 (N_5988,N_4112,N_4674);
xnor U5989 (N_5989,N_4416,N_4249);
nor U5990 (N_5990,N_4242,N_3782);
or U5991 (N_5991,N_3784,N_3710);
and U5992 (N_5992,N_4109,N_3620);
nor U5993 (N_5993,N_4381,N_4509);
and U5994 (N_5994,N_4500,N_3702);
nor U5995 (N_5995,N_4214,N_4579);
xnor U5996 (N_5996,N_3849,N_4412);
and U5997 (N_5997,N_3935,N_4635);
nor U5998 (N_5998,N_4781,N_3706);
nand U5999 (N_5999,N_3717,N_3866);
nand U6000 (N_6000,N_5836,N_5840);
and U6001 (N_6001,N_5403,N_5070);
or U6002 (N_6002,N_5777,N_5930);
xor U6003 (N_6003,N_5878,N_5555);
and U6004 (N_6004,N_5523,N_5668);
or U6005 (N_6005,N_5263,N_5716);
and U6006 (N_6006,N_5311,N_5073);
and U6007 (N_6007,N_5140,N_5478);
and U6008 (N_6008,N_5879,N_5036);
nor U6009 (N_6009,N_5327,N_5788);
and U6010 (N_6010,N_5155,N_5305);
or U6011 (N_6011,N_5394,N_5886);
xor U6012 (N_6012,N_5134,N_4990);
xor U6013 (N_6013,N_5530,N_5314);
xor U6014 (N_6014,N_5876,N_5321);
nand U6015 (N_6015,N_5242,N_5971);
nand U6016 (N_6016,N_5481,N_4862);
and U6017 (N_6017,N_4907,N_5679);
or U6018 (N_6018,N_4893,N_4816);
or U6019 (N_6019,N_5180,N_5376);
and U6020 (N_6020,N_5737,N_5590);
xor U6021 (N_6021,N_5553,N_5884);
and U6022 (N_6022,N_5994,N_5345);
nor U6023 (N_6023,N_5597,N_5487);
nand U6024 (N_6024,N_5191,N_5343);
and U6025 (N_6025,N_4944,N_4942);
and U6026 (N_6026,N_5386,N_5492);
or U6027 (N_6027,N_5916,N_5429);
and U6028 (N_6028,N_5572,N_5575);
or U6029 (N_6029,N_5402,N_5453);
xnor U6030 (N_6030,N_5577,N_5174);
nor U6031 (N_6031,N_5759,N_5200);
and U6032 (N_6032,N_5820,N_5677);
and U6033 (N_6033,N_5861,N_4805);
xor U6034 (N_6034,N_5604,N_5987);
or U6035 (N_6035,N_5338,N_5703);
nor U6036 (N_6036,N_5982,N_5816);
nand U6037 (N_6037,N_5256,N_5248);
nor U6038 (N_6038,N_4917,N_5819);
xnor U6039 (N_6039,N_5849,N_5011);
nand U6040 (N_6040,N_4953,N_5154);
and U6041 (N_6041,N_5661,N_5326);
nand U6042 (N_6042,N_5917,N_5379);
xnor U6043 (N_6043,N_5937,N_5885);
or U6044 (N_6044,N_5293,N_5302);
and U6045 (N_6045,N_4965,N_4859);
nand U6046 (N_6046,N_5100,N_4898);
or U6047 (N_6047,N_5099,N_5475);
nor U6048 (N_6048,N_5975,N_5583);
nor U6049 (N_6049,N_5556,N_5225);
nand U6050 (N_6050,N_5391,N_5729);
nand U6051 (N_6051,N_5918,N_5244);
nor U6052 (N_6052,N_5924,N_5898);
nor U6053 (N_6053,N_5789,N_5570);
and U6054 (N_6054,N_5694,N_5750);
and U6055 (N_6055,N_5638,N_5347);
and U6056 (N_6056,N_5805,N_5204);
or U6057 (N_6057,N_4939,N_5464);
nor U6058 (N_6058,N_5420,N_4950);
and U6059 (N_6059,N_5418,N_5355);
nand U6060 (N_6060,N_5371,N_5584);
nand U6061 (N_6061,N_5044,N_5760);
and U6062 (N_6062,N_5337,N_5253);
or U6063 (N_6063,N_5156,N_4921);
and U6064 (N_6064,N_5522,N_5881);
nor U6065 (N_6065,N_5657,N_4813);
or U6066 (N_6066,N_5936,N_5166);
nor U6067 (N_6067,N_5368,N_5064);
and U6068 (N_6068,N_5163,N_5037);
and U6069 (N_6069,N_5653,N_5127);
nor U6070 (N_6070,N_4923,N_4909);
nor U6071 (N_6071,N_5565,N_4838);
nor U6072 (N_6072,N_4978,N_5817);
nand U6073 (N_6073,N_5245,N_5187);
and U6074 (N_6074,N_5151,N_5153);
nand U6075 (N_6075,N_5354,N_5656);
xnor U6076 (N_6076,N_5152,N_5755);
and U6077 (N_6077,N_5260,N_5954);
nor U6078 (N_6078,N_4910,N_5602);
and U6079 (N_6079,N_5542,N_5043);
xor U6080 (N_6080,N_5297,N_5366);
or U6081 (N_6081,N_5637,N_4889);
nand U6082 (N_6082,N_5624,N_5614);
and U6083 (N_6083,N_5220,N_5961);
or U6084 (N_6084,N_5065,N_5758);
xnor U6085 (N_6085,N_5616,N_4870);
xnor U6086 (N_6086,N_5844,N_4872);
and U6087 (N_6087,N_5240,N_5528);
and U6088 (N_6088,N_5234,N_5809);
and U6089 (N_6089,N_5102,N_4974);
nor U6090 (N_6090,N_5400,N_5280);
nor U6091 (N_6091,N_5251,N_5459);
xor U6092 (N_6092,N_5821,N_5723);
or U6093 (N_6093,N_5610,N_5237);
nand U6094 (N_6094,N_5843,N_5157);
nand U6095 (N_6095,N_5873,N_5678);
and U6096 (N_6096,N_5667,N_5945);
or U6097 (N_6097,N_4854,N_4997);
and U6098 (N_6098,N_4964,N_5482);
and U6099 (N_6099,N_4967,N_5951);
or U6100 (N_6100,N_5202,N_5933);
xnor U6101 (N_6101,N_5895,N_4962);
nor U6102 (N_6102,N_5005,N_5199);
xor U6103 (N_6103,N_4858,N_5985);
nand U6104 (N_6104,N_5880,N_5589);
nand U6105 (N_6105,N_5865,N_5525);
xnor U6106 (N_6106,N_4820,N_5427);
nor U6107 (N_6107,N_4979,N_5019);
nand U6108 (N_6108,N_4973,N_5634);
xnor U6109 (N_6109,N_5010,N_5130);
xnor U6110 (N_6110,N_5591,N_5718);
nor U6111 (N_6111,N_5664,N_4900);
and U6112 (N_6112,N_5607,N_5193);
nand U6113 (N_6113,N_5052,N_5033);
nor U6114 (N_6114,N_5965,N_5243);
xor U6115 (N_6115,N_5742,N_4951);
and U6116 (N_6116,N_4840,N_5219);
nand U6117 (N_6117,N_4876,N_5324);
or U6118 (N_6118,N_5957,N_5807);
nor U6119 (N_6119,N_5279,N_5491);
and U6120 (N_6120,N_4981,N_4952);
nor U6121 (N_6121,N_5651,N_5135);
xor U6122 (N_6122,N_5644,N_5510);
xnor U6123 (N_6123,N_5440,N_5692);
or U6124 (N_6124,N_5514,N_5516);
xnor U6125 (N_6125,N_5986,N_5801);
nand U6126 (N_6126,N_5210,N_4856);
nand U6127 (N_6127,N_4830,N_4970);
nand U6128 (N_6128,N_5230,N_4968);
or U6129 (N_6129,N_5058,N_5007);
xor U6130 (N_6130,N_5313,N_5900);
xnor U6131 (N_6131,N_5833,N_5866);
nand U6132 (N_6132,N_5619,N_5867);
and U6133 (N_6133,N_5286,N_5796);
or U6134 (N_6134,N_4824,N_5113);
xor U6135 (N_6135,N_5336,N_5888);
xnor U6136 (N_6136,N_5707,N_4972);
nor U6137 (N_6137,N_5015,N_5894);
nand U6138 (N_6138,N_5686,N_5369);
or U6139 (N_6139,N_4928,N_4938);
nor U6140 (N_6140,N_4926,N_4986);
xnor U6141 (N_6141,N_5361,N_5800);
xnor U6142 (N_6142,N_5507,N_5799);
or U6143 (N_6143,N_5068,N_4945);
nor U6144 (N_6144,N_5623,N_5942);
and U6145 (N_6145,N_5483,N_5518);
nor U6146 (N_6146,N_5460,N_5471);
nand U6147 (N_6147,N_4869,N_4918);
xnor U6148 (N_6148,N_5261,N_4943);
and U6149 (N_6149,N_5964,N_5207);
xor U6150 (N_6150,N_4821,N_5098);
nand U6151 (N_6151,N_5477,N_5283);
xnor U6152 (N_6152,N_5693,N_5825);
xor U6153 (N_6153,N_4819,N_5650);
or U6154 (N_6154,N_5559,N_4920);
xor U6155 (N_6155,N_5506,N_5480);
and U6156 (N_6156,N_5672,N_4887);
nor U6157 (N_6157,N_5067,N_5296);
and U6158 (N_6158,N_5598,N_5090);
or U6159 (N_6159,N_5162,N_5288);
or U6160 (N_6160,N_5582,N_5545);
nor U6161 (N_6161,N_5743,N_5103);
nand U6162 (N_6162,N_5050,N_5883);
nor U6163 (N_6163,N_5864,N_4983);
nand U6164 (N_6164,N_5952,N_5276);
or U6165 (N_6165,N_5171,N_5105);
nor U6166 (N_6166,N_5748,N_5762);
xor U6167 (N_6167,N_5787,N_5647);
and U6168 (N_6168,N_5419,N_4879);
or U6169 (N_6169,N_5282,N_5967);
and U6170 (N_6170,N_5824,N_5784);
and U6171 (N_6171,N_5578,N_5786);
nand U6172 (N_6172,N_5983,N_5500);
and U6173 (N_6173,N_4860,N_5332);
xor U6174 (N_6174,N_5791,N_4906);
nand U6175 (N_6175,N_5365,N_5841);
and U6176 (N_6176,N_5995,N_5144);
nor U6177 (N_6177,N_5978,N_5358);
nand U6178 (N_6178,N_4998,N_5869);
and U6179 (N_6179,N_5989,N_5968);
or U6180 (N_6180,N_5740,N_5177);
or U6181 (N_6181,N_5027,N_5505);
and U6182 (N_6182,N_5325,N_4847);
nor U6183 (N_6183,N_5095,N_5689);
nand U6184 (N_6184,N_5695,N_5018);
nor U6185 (N_6185,N_5673,N_5615);
xnor U6186 (N_6186,N_5012,N_5744);
and U6187 (N_6187,N_5030,N_5882);
and U6188 (N_6188,N_5446,N_5124);
and U6189 (N_6189,N_5054,N_5513);
and U6190 (N_6190,N_5367,N_5974);
or U6191 (N_6191,N_5465,N_5990);
nand U6192 (N_6192,N_5097,N_5766);
nand U6193 (N_6193,N_5897,N_5906);
and U6194 (N_6194,N_4886,N_5189);
or U6195 (N_6195,N_4884,N_5573);
xnor U6196 (N_6196,N_5594,N_5811);
xor U6197 (N_6197,N_5736,N_5229);
nand U6198 (N_6198,N_5176,N_5142);
nand U6199 (N_6199,N_5357,N_5250);
xor U6200 (N_6200,N_5851,N_5259);
and U6201 (N_6201,N_5804,N_5392);
nor U6202 (N_6202,N_5870,N_5797);
xor U6203 (N_6203,N_5085,N_4929);
nand U6204 (N_6204,N_5699,N_5449);
nand U6205 (N_6205,N_5309,N_5436);
and U6206 (N_6206,N_5641,N_5104);
or U6207 (N_6207,N_5585,N_5246);
xor U6208 (N_6208,N_5101,N_5398);
nor U6209 (N_6209,N_5441,N_4941);
and U6210 (N_6210,N_5295,N_5258);
nand U6211 (N_6211,N_5706,N_5854);
xor U6212 (N_6212,N_5026,N_5387);
or U6213 (N_6213,N_4896,N_5133);
or U6214 (N_6214,N_5375,N_4806);
xor U6215 (N_6215,N_5221,N_5722);
or U6216 (N_6216,N_4888,N_5117);
xor U6217 (N_6217,N_4848,N_5648);
nand U6218 (N_6218,N_5775,N_4996);
nor U6219 (N_6219,N_5312,N_5108);
nor U6220 (N_6220,N_5136,N_5963);
nor U6221 (N_6221,N_5285,N_4922);
and U6222 (N_6222,N_5874,N_5094);
or U6223 (N_6223,N_5080,N_5197);
nor U6224 (N_6224,N_4958,N_5813);
or U6225 (N_6225,N_5914,N_5034);
xnor U6226 (N_6226,N_5546,N_5999);
and U6227 (N_6227,N_5631,N_4851);
nand U6228 (N_6228,N_5741,N_4829);
or U6229 (N_6229,N_5992,N_4849);
nor U6230 (N_6230,N_4985,N_5928);
and U6231 (N_6231,N_5734,N_5123);
or U6232 (N_6232,N_5909,N_5935);
nand U6233 (N_6233,N_5254,N_5808);
nor U6234 (N_6234,N_5955,N_5915);
nand U6235 (N_6235,N_4809,N_5752);
and U6236 (N_6236,N_5397,N_4864);
xnor U6237 (N_6237,N_5850,N_5426);
or U6238 (N_6238,N_5993,N_5066);
nand U6239 (N_6239,N_5934,N_5960);
or U6240 (N_6240,N_5172,N_4994);
xnor U6241 (N_6241,N_5927,N_5063);
nand U6242 (N_6242,N_5378,N_5349);
nor U6243 (N_6243,N_4932,N_5255);
nor U6244 (N_6244,N_5364,N_4823);
and U6245 (N_6245,N_4988,N_5088);
xor U6246 (N_6246,N_5148,N_5201);
xnor U6247 (N_6247,N_5713,N_5691);
nor U6248 (N_6248,N_4811,N_5318);
or U6249 (N_6249,N_5016,N_5306);
and U6250 (N_6250,N_5399,N_5452);
nor U6251 (N_6251,N_4995,N_4960);
and U6252 (N_6252,N_4815,N_5212);
or U6253 (N_6253,N_5534,N_5020);
nand U6254 (N_6254,N_4825,N_5605);
nand U6255 (N_6255,N_5435,N_4812);
xnor U6256 (N_6256,N_4853,N_5227);
xor U6257 (N_6257,N_5905,N_5508);
or U6258 (N_6258,N_5275,N_5138);
xnor U6259 (N_6259,N_4975,N_5214);
nor U6260 (N_6260,N_5595,N_5447);
and U6261 (N_6261,N_5627,N_5238);
or U6262 (N_6262,N_5941,N_5751);
nand U6263 (N_6263,N_5128,N_5724);
nand U6264 (N_6264,N_4925,N_5970);
and U6265 (N_6265,N_4999,N_5676);
xnor U6266 (N_6266,N_5074,N_5538);
xnor U6267 (N_6267,N_5772,N_5984);
nand U6268 (N_6268,N_5735,N_5490);
and U6269 (N_6269,N_4875,N_5558);
or U6270 (N_6270,N_5473,N_5931);
or U6271 (N_6271,N_5947,N_5511);
nand U6272 (N_6272,N_5298,N_5684);
or U6273 (N_6273,N_5901,N_5083);
and U6274 (N_6274,N_4937,N_5574);
or U6275 (N_6275,N_5862,N_5185);
xor U6276 (N_6276,N_4835,N_5903);
or U6277 (N_6277,N_5976,N_5795);
nor U6278 (N_6278,N_5503,N_5056);
or U6279 (N_6279,N_5890,N_5421);
and U6280 (N_6280,N_5270,N_5596);
and U6281 (N_6281,N_5126,N_5389);
nor U6282 (N_6282,N_4842,N_5443);
or U6283 (N_6283,N_5904,N_5456);
and U6284 (N_6284,N_5669,N_5536);
nand U6285 (N_6285,N_4873,N_5072);
nand U6286 (N_6286,N_5537,N_5738);
xnor U6287 (N_6287,N_5586,N_4880);
or U6288 (N_6288,N_5198,N_5437);
and U6289 (N_6289,N_5145,N_5494);
xor U6290 (N_6290,N_5137,N_5600);
nand U6291 (N_6291,N_5749,N_5708);
xnor U6292 (N_6292,N_5409,N_4895);
nand U6293 (N_6293,N_5544,N_4903);
and U6294 (N_6294,N_5618,N_5024);
or U6295 (N_6295,N_5726,N_5252);
nor U6296 (N_6296,N_4865,N_4959);
nand U6297 (N_6297,N_5329,N_5182);
and U6298 (N_6298,N_5416,N_5444);
xnor U6299 (N_6299,N_5532,N_5632);
nor U6300 (N_6300,N_5075,N_5539);
nor U6301 (N_6301,N_5812,N_4924);
nor U6302 (N_6302,N_5504,N_5265);
or U6303 (N_6303,N_5962,N_5352);
nand U6304 (N_6304,N_5919,N_5649);
or U6305 (N_6305,N_5509,N_4954);
xor U6306 (N_6306,N_5633,N_5654);
or U6307 (N_6307,N_4961,N_5401);
nor U6308 (N_6308,N_5696,N_5793);
and U6309 (N_6309,N_5423,N_5164);
nand U6310 (N_6310,N_5889,N_5169);
xnor U6311 (N_6311,N_5868,N_5988);
nor U6312 (N_6312,N_5038,N_5488);
or U6313 (N_6313,N_5118,N_5146);
nor U6314 (N_6314,N_5489,N_5949);
xnor U6315 (N_6315,N_5388,N_5110);
nor U6316 (N_6316,N_5636,N_5060);
and U6317 (N_6317,N_5776,N_5715);
nor U6318 (N_6318,N_5374,N_5771);
nand U6319 (N_6319,N_5495,N_5685);
or U6320 (N_6320,N_5687,N_4818);
nor U6321 (N_6321,N_5980,N_4837);
and U6322 (N_6322,N_5853,N_4949);
nand U6323 (N_6323,N_5588,N_5408);
nand U6324 (N_6324,N_4861,N_5714);
and U6325 (N_6325,N_5739,N_5300);
xnor U6326 (N_6326,N_5003,N_5131);
nand U6327 (N_6327,N_5533,N_5670);
and U6328 (N_6328,N_5055,N_5404);
or U6329 (N_6329,N_5926,N_5022);
nor U6330 (N_6330,N_5448,N_5173);
or U6331 (N_6331,N_4810,N_4934);
nor U6332 (N_6332,N_5838,N_5032);
nor U6333 (N_6333,N_5896,N_5384);
or U6334 (N_6334,N_5241,N_5877);
or U6335 (N_6335,N_5262,N_5773);
or U6336 (N_6336,N_5733,N_5158);
xnor U6337 (N_6337,N_4946,N_5213);
and U6338 (N_6338,N_5093,N_5428);
or U6339 (N_6339,N_5121,N_5554);
or U6340 (N_6340,N_5639,N_5268);
nand U6341 (N_6341,N_5021,N_5373);
nand U6342 (N_6342,N_5946,N_5304);
nor U6343 (N_6343,N_5139,N_5761);
and U6344 (N_6344,N_4868,N_4894);
or U6345 (N_6345,N_5835,N_5048);
or U6346 (N_6346,N_4871,N_5485);
nand U6347 (N_6347,N_5781,N_5948);
and U6348 (N_6348,N_5730,N_5129);
and U6349 (N_6349,N_5360,N_5450);
or U6350 (N_6350,N_5818,N_5106);
xnor U6351 (N_6351,N_5071,N_5217);
nor U6352 (N_6352,N_5847,N_5161);
and U6353 (N_6353,N_5061,N_5828);
and U6354 (N_6354,N_5697,N_5764);
nor U6355 (N_6355,N_5798,N_5192);
nand U6356 (N_6356,N_5690,N_4802);
nand U6357 (N_6357,N_5496,N_5794);
and U6358 (N_6358,N_5362,N_5266);
nand U6359 (N_6359,N_5159,N_4804);
or U6360 (N_6360,N_5540,N_5863);
xnor U6361 (N_6361,N_5902,N_5042);
or U6362 (N_6362,N_5997,N_5377);
or U6363 (N_6363,N_5548,N_5620);
and U6364 (N_6364,N_5823,N_5560);
and U6365 (N_6365,N_5592,N_4940);
nand U6366 (N_6366,N_5810,N_5603);
or U6367 (N_6367,N_5290,N_5712);
nor U6368 (N_6368,N_5710,N_4948);
nand U6369 (N_6369,N_5175,N_5385);
or U6370 (N_6370,N_5417,N_5287);
or U6371 (N_6371,N_5790,N_5203);
and U6372 (N_6372,N_5049,N_5702);
nor U6373 (N_6373,N_5497,N_5186);
nor U6374 (N_6374,N_4914,N_5660);
nor U6375 (N_6375,N_4883,N_5704);
and U6376 (N_6376,N_5208,N_5587);
nor U6377 (N_6377,N_5893,N_5778);
or U6378 (N_6378,N_5628,N_4897);
or U6379 (N_6379,N_5527,N_5330);
nand U6380 (N_6380,N_5120,N_5316);
and U6381 (N_6381,N_5827,N_5013);
and U6382 (N_6382,N_5267,N_5579);
xnor U6383 (N_6383,N_5765,N_5082);
and U6384 (N_6384,N_5822,N_4885);
xor U6385 (N_6385,N_5233,N_5529);
or U6386 (N_6386,N_4916,N_5451);
nor U6387 (N_6387,N_4839,N_5006);
and U6388 (N_6388,N_5396,N_5216);
and U6389 (N_6389,N_5040,N_5467);
xor U6390 (N_6390,N_5346,N_5950);
or U6391 (N_6391,N_5859,N_5531);
nand U6392 (N_6392,N_5271,N_5745);
and U6393 (N_6393,N_5224,N_5046);
nor U6394 (N_6394,N_5940,N_5476);
xnor U6395 (N_6395,N_5091,N_5087);
xor U6396 (N_6396,N_5593,N_5183);
nand U6397 (N_6397,N_5470,N_5719);
xor U6398 (N_6398,N_4822,N_5269);
or U6399 (N_6399,N_5381,N_5682);
xor U6400 (N_6400,N_5031,N_5576);
xnor U6401 (N_6401,N_5831,N_5837);
and U6402 (N_6402,N_4989,N_5303);
xor U6403 (N_6403,N_4892,N_4915);
or U6404 (N_6404,N_5076,N_5413);
xnor U6405 (N_6405,N_5484,N_5939);
nand U6406 (N_6406,N_5659,N_4874);
nor U6407 (N_6407,N_4850,N_4828);
xnor U6408 (N_6408,N_5756,N_5348);
nand U6409 (N_6409,N_4808,N_5768);
and U6410 (N_6410,N_5194,N_5643);
or U6411 (N_6411,N_5004,N_5335);
and U6412 (N_6412,N_5116,N_5390);
nor U6413 (N_6413,N_4817,N_5683);
nand U6414 (N_6414,N_5168,N_5165);
or U6415 (N_6415,N_5041,N_5721);
nand U6416 (N_6416,N_5350,N_4919);
nor U6417 (N_6417,N_4904,N_5114);
nor U6418 (N_6418,N_5053,N_5769);
or U6419 (N_6419,N_5566,N_5705);
xnor U6420 (N_6420,N_5323,N_4878);
and U6421 (N_6421,N_5674,N_5622);
nand U6422 (N_6422,N_5308,N_5580);
nor U6423 (N_6423,N_5414,N_5564);
or U6424 (N_6424,N_5188,N_5519);
nand U6425 (N_6425,N_5551,N_5938);
or U6426 (N_6426,N_5727,N_5222);
nand U6427 (N_6427,N_5855,N_5433);
xnor U6428 (N_6428,N_4957,N_5609);
or U6429 (N_6429,N_5671,N_5543);
and U6430 (N_6430,N_5395,N_4905);
or U6431 (N_6431,N_5466,N_5057);
nand U6432 (N_6432,N_5953,N_5763);
or U6433 (N_6433,N_5658,N_5458);
nor U6434 (N_6434,N_5150,N_5552);
nand U6435 (N_6435,N_4992,N_4863);
nor U6436 (N_6436,N_5430,N_5785);
or U6437 (N_6437,N_5517,N_5956);
and U6438 (N_6438,N_5912,N_5774);
or U6439 (N_6439,N_5017,N_5342);
and U6440 (N_6440,N_5284,N_5701);
and U6441 (N_6441,N_5249,N_5431);
or U6442 (N_6442,N_5425,N_5081);
and U6443 (N_6443,N_5929,N_5001);
and U6444 (N_6444,N_5943,N_5319);
and U6445 (N_6445,N_5415,N_5331);
nor U6446 (N_6446,N_5645,N_5499);
nand U6447 (N_6447,N_5991,N_5806);
nor U6448 (N_6448,N_5845,N_5132);
nor U6449 (N_6449,N_4976,N_5351);
nand U6450 (N_6450,N_5190,N_4899);
nor U6451 (N_6451,N_5932,N_5062);
nor U6452 (N_6452,N_5257,N_5782);
nor U6453 (N_6453,N_5272,N_5322);
and U6454 (N_6454,N_5317,N_5344);
and U6455 (N_6455,N_5009,N_4993);
or U6456 (N_6456,N_5569,N_5626);
nor U6457 (N_6457,N_5029,N_5493);
nor U6458 (N_6458,N_5205,N_4807);
nand U6459 (N_6459,N_5195,N_5871);
nor U6460 (N_6460,N_5051,N_5218);
nand U6461 (N_6461,N_5662,N_5732);
nor U6462 (N_6462,N_5277,N_4834);
xor U6463 (N_6463,N_5725,N_5802);
xnor U6464 (N_6464,N_5547,N_5625);
nand U6465 (N_6465,N_5226,N_5469);
nor U6466 (N_6466,N_5411,N_5393);
nor U6467 (N_6467,N_5289,N_5112);
nand U6468 (N_6468,N_5754,N_5410);
or U6469 (N_6469,N_5830,N_5521);
xnor U6470 (N_6470,N_4933,N_4852);
xnor U6471 (N_6471,N_5911,N_5512);
or U6472 (N_6472,N_5611,N_5747);
nand U6473 (N_6473,N_5892,N_5178);
xor U6474 (N_6474,N_5872,N_5468);
nor U6475 (N_6475,N_4882,N_5359);
nor U6476 (N_6476,N_5278,N_5728);
nand U6477 (N_6477,N_5315,N_5665);
and U6478 (N_6478,N_5700,N_5612);
nand U6479 (N_6479,N_5299,N_5601);
nor U6480 (N_6480,N_5445,N_4980);
nor U6481 (N_6481,N_5731,N_5328);
nor U6482 (N_6482,N_5424,N_5630);
xor U6483 (N_6483,N_4891,N_4908);
and U6484 (N_6484,N_5111,N_4935);
and U6485 (N_6485,N_5274,N_4841);
nor U6486 (N_6486,N_5406,N_5196);
nor U6487 (N_6487,N_5655,N_5563);
or U6488 (N_6488,N_4991,N_4890);
xnor U6489 (N_6489,N_5709,N_5923);
xnor U6490 (N_6490,N_5606,N_5002);
and U6491 (N_6491,N_4987,N_5977);
nand U6492 (N_6492,N_5652,N_5640);
nor U6493 (N_6493,N_5167,N_5432);
and U6494 (N_6494,N_5921,N_5086);
and U6495 (N_6495,N_5310,N_4801);
nor U6496 (N_6496,N_5228,N_5439);
and U6497 (N_6497,N_5307,N_5535);
and U6498 (N_6498,N_5239,N_4832);
nand U6499 (N_6499,N_5235,N_5363);
and U6500 (N_6500,N_5910,N_4947);
and U6501 (N_6501,N_5996,N_4845);
and U6502 (N_6502,N_5842,N_5206);
and U6503 (N_6503,N_5858,N_5035);
and U6504 (N_6504,N_5125,N_5215);
xor U6505 (N_6505,N_4827,N_5720);
or U6506 (N_6506,N_4803,N_5571);
nand U6507 (N_6507,N_5839,N_5028);
nand U6508 (N_6508,N_5236,N_5079);
xor U6509 (N_6509,N_5479,N_5438);
nor U6510 (N_6510,N_5045,N_4982);
xor U6511 (N_6511,N_4866,N_5550);
and U6512 (N_6512,N_5635,N_5008);
nor U6513 (N_6513,N_5209,N_5292);
nor U6514 (N_6514,N_5000,N_4881);
nor U6515 (N_6515,N_5698,N_5524);
nor U6516 (N_6516,N_5966,N_4833);
xnor U6517 (N_6517,N_5059,N_5958);
or U6518 (N_6518,N_5141,N_5856);
and U6519 (N_6519,N_5998,N_5770);
or U6520 (N_6520,N_5908,N_5143);
and U6521 (N_6521,N_5122,N_5688);
xnor U6522 (N_6522,N_5109,N_4927);
and U6523 (N_6523,N_5568,N_5680);
and U6524 (N_6524,N_5281,N_5077);
nor U6525 (N_6525,N_5852,N_5826);
or U6526 (N_6526,N_4966,N_5023);
nand U6527 (N_6527,N_5792,N_5857);
or U6528 (N_6528,N_5407,N_5541);
or U6529 (N_6529,N_5372,N_5642);
xor U6530 (N_6530,N_5981,N_5846);
nand U6531 (N_6531,N_5084,N_5562);
nor U6532 (N_6532,N_5832,N_5092);
xor U6533 (N_6533,N_5887,N_4800);
nor U6534 (N_6534,N_5333,N_5455);
xor U6535 (N_6535,N_4984,N_5078);
nand U6536 (N_6536,N_5264,N_5179);
nor U6537 (N_6537,N_5457,N_4930);
nor U6538 (N_6538,N_5115,N_5973);
xor U6539 (N_6539,N_5666,N_5412);
nor U6540 (N_6540,N_5422,N_5462);
xnor U6541 (N_6541,N_5211,N_5780);
nor U6542 (N_6542,N_4969,N_4844);
or U6543 (N_6543,N_5223,N_5629);
or U6544 (N_6544,N_5779,N_4843);
nand U6545 (N_6545,N_5463,N_5380);
nand U6546 (N_6546,N_4877,N_5273);
or U6547 (N_6547,N_5096,N_5815);
xnor U6548 (N_6548,N_4831,N_5160);
xor U6549 (N_6549,N_5149,N_4836);
and U6550 (N_6550,N_4971,N_5663);
nand U6551 (N_6551,N_4931,N_5119);
xor U6552 (N_6552,N_5920,N_5907);
nor U6553 (N_6553,N_5599,N_5486);
and U6554 (N_6554,N_5294,N_5944);
nor U6555 (N_6555,N_5320,N_5561);
and U6556 (N_6556,N_4826,N_5442);
and U6557 (N_6557,N_4902,N_5014);
or U6558 (N_6558,N_5383,N_5515);
nand U6559 (N_6559,N_5334,N_4857);
and U6560 (N_6560,N_5613,N_5860);
and U6561 (N_6561,N_4956,N_4867);
nand U6562 (N_6562,N_5803,N_5899);
nor U6563 (N_6563,N_4814,N_5353);
nand U6564 (N_6564,N_4855,N_5047);
nand U6565 (N_6565,N_5979,N_5472);
nor U6566 (N_6566,N_4846,N_5875);
nand U6567 (N_6567,N_5147,N_5291);
xnor U6568 (N_6568,N_5434,N_5498);
or U6569 (N_6569,N_5370,N_5757);
xor U6570 (N_6570,N_5502,N_5025);
nand U6571 (N_6571,N_5567,N_5959);
or U6572 (N_6572,N_5969,N_5675);
and U6573 (N_6573,N_5454,N_5181);
or U6574 (N_6574,N_5069,N_5767);
nand U6575 (N_6575,N_4963,N_4913);
nor U6576 (N_6576,N_5621,N_5356);
and U6577 (N_6577,N_5922,N_5340);
nand U6578 (N_6578,N_5746,N_5581);
nand U6579 (N_6579,N_5972,N_5231);
and U6580 (N_6580,N_5681,N_5753);
or U6581 (N_6581,N_5526,N_5339);
nand U6582 (N_6582,N_5405,N_5646);
xnor U6583 (N_6583,N_5717,N_5170);
and U6584 (N_6584,N_5608,N_5549);
and U6585 (N_6585,N_5461,N_5834);
nor U6586 (N_6586,N_5913,N_5107);
or U6587 (N_6587,N_4911,N_5783);
nor U6588 (N_6588,N_5382,N_4912);
nand U6589 (N_6589,N_5829,N_5341);
nor U6590 (N_6590,N_5617,N_4955);
or U6591 (N_6591,N_5184,N_5520);
or U6592 (N_6592,N_4936,N_5474);
nor U6593 (N_6593,N_5501,N_5247);
nor U6594 (N_6594,N_5039,N_4977);
nand U6595 (N_6595,N_5557,N_4901);
xnor U6596 (N_6596,N_5711,N_5814);
and U6597 (N_6597,N_5848,N_5301);
nand U6598 (N_6598,N_5089,N_5925);
or U6599 (N_6599,N_5891,N_5232);
nand U6600 (N_6600,N_5152,N_5714);
xnor U6601 (N_6601,N_5142,N_4904);
xnor U6602 (N_6602,N_5581,N_5330);
nor U6603 (N_6603,N_5380,N_5006);
nand U6604 (N_6604,N_5082,N_5095);
nand U6605 (N_6605,N_5435,N_4989);
nand U6606 (N_6606,N_5238,N_4918);
and U6607 (N_6607,N_5285,N_5214);
or U6608 (N_6608,N_5032,N_5949);
and U6609 (N_6609,N_5814,N_4925);
xor U6610 (N_6610,N_5534,N_5584);
xor U6611 (N_6611,N_5633,N_4833);
and U6612 (N_6612,N_5702,N_5957);
nor U6613 (N_6613,N_4821,N_5746);
nand U6614 (N_6614,N_5665,N_4905);
nor U6615 (N_6615,N_4862,N_5299);
xnor U6616 (N_6616,N_5337,N_4863);
or U6617 (N_6617,N_5389,N_5383);
nand U6618 (N_6618,N_5790,N_4853);
xor U6619 (N_6619,N_5111,N_5823);
xor U6620 (N_6620,N_4933,N_5232);
nor U6621 (N_6621,N_5160,N_4965);
nor U6622 (N_6622,N_5991,N_5795);
xnor U6623 (N_6623,N_5166,N_5159);
nand U6624 (N_6624,N_5870,N_5374);
nor U6625 (N_6625,N_5598,N_4814);
nand U6626 (N_6626,N_5482,N_5540);
xnor U6627 (N_6627,N_4980,N_5698);
nor U6628 (N_6628,N_5347,N_5422);
or U6629 (N_6629,N_5951,N_4960);
or U6630 (N_6630,N_5697,N_5232);
nor U6631 (N_6631,N_5236,N_5645);
and U6632 (N_6632,N_5922,N_4961);
xor U6633 (N_6633,N_5605,N_5073);
nand U6634 (N_6634,N_5470,N_5595);
or U6635 (N_6635,N_5040,N_5838);
xnor U6636 (N_6636,N_5833,N_5450);
and U6637 (N_6637,N_5965,N_5351);
and U6638 (N_6638,N_5831,N_5722);
and U6639 (N_6639,N_5532,N_5442);
or U6640 (N_6640,N_5785,N_4856);
nand U6641 (N_6641,N_4859,N_5414);
xor U6642 (N_6642,N_5116,N_5127);
or U6643 (N_6643,N_5084,N_5791);
nand U6644 (N_6644,N_4897,N_5885);
xor U6645 (N_6645,N_5914,N_4881);
xnor U6646 (N_6646,N_5193,N_5961);
or U6647 (N_6647,N_5814,N_5965);
and U6648 (N_6648,N_5226,N_5185);
and U6649 (N_6649,N_5722,N_4953);
nor U6650 (N_6650,N_4928,N_5496);
or U6651 (N_6651,N_4836,N_5817);
xnor U6652 (N_6652,N_5062,N_5540);
xor U6653 (N_6653,N_5951,N_5693);
or U6654 (N_6654,N_5890,N_5130);
or U6655 (N_6655,N_5577,N_4883);
nor U6656 (N_6656,N_4870,N_5414);
nand U6657 (N_6657,N_5972,N_5699);
xnor U6658 (N_6658,N_5225,N_5318);
nor U6659 (N_6659,N_4869,N_5389);
and U6660 (N_6660,N_5200,N_5629);
xnor U6661 (N_6661,N_5116,N_5167);
nor U6662 (N_6662,N_5578,N_5799);
nand U6663 (N_6663,N_5024,N_5217);
xor U6664 (N_6664,N_5016,N_5141);
xnor U6665 (N_6665,N_5812,N_5211);
xor U6666 (N_6666,N_5096,N_5035);
and U6667 (N_6667,N_5621,N_4893);
or U6668 (N_6668,N_5101,N_5555);
nand U6669 (N_6669,N_4928,N_5551);
xor U6670 (N_6670,N_5964,N_5595);
nor U6671 (N_6671,N_5341,N_5641);
nor U6672 (N_6672,N_5975,N_5042);
and U6673 (N_6673,N_5799,N_5003);
nor U6674 (N_6674,N_5829,N_4801);
xnor U6675 (N_6675,N_5255,N_5616);
nand U6676 (N_6676,N_5406,N_5581);
xnor U6677 (N_6677,N_5249,N_5575);
xnor U6678 (N_6678,N_5367,N_5203);
and U6679 (N_6679,N_4909,N_5759);
or U6680 (N_6680,N_5190,N_5369);
or U6681 (N_6681,N_5456,N_4937);
nor U6682 (N_6682,N_4928,N_5063);
or U6683 (N_6683,N_5424,N_5211);
nor U6684 (N_6684,N_5465,N_5926);
and U6685 (N_6685,N_5307,N_5981);
nor U6686 (N_6686,N_5306,N_5421);
nor U6687 (N_6687,N_5680,N_5724);
nand U6688 (N_6688,N_5076,N_5694);
and U6689 (N_6689,N_5263,N_5308);
nor U6690 (N_6690,N_5403,N_4827);
xnor U6691 (N_6691,N_5723,N_5784);
xnor U6692 (N_6692,N_5216,N_5289);
nor U6693 (N_6693,N_5504,N_4863);
xnor U6694 (N_6694,N_5714,N_5258);
or U6695 (N_6695,N_5449,N_5708);
xor U6696 (N_6696,N_5948,N_5137);
or U6697 (N_6697,N_5369,N_5392);
or U6698 (N_6698,N_5411,N_5277);
nand U6699 (N_6699,N_5208,N_5603);
xor U6700 (N_6700,N_5206,N_5624);
or U6701 (N_6701,N_5844,N_5379);
or U6702 (N_6702,N_4855,N_5931);
nor U6703 (N_6703,N_5636,N_5912);
or U6704 (N_6704,N_5701,N_5162);
nor U6705 (N_6705,N_4878,N_5473);
xnor U6706 (N_6706,N_5343,N_5965);
xor U6707 (N_6707,N_5479,N_4972);
or U6708 (N_6708,N_5845,N_4803);
nand U6709 (N_6709,N_4971,N_5594);
or U6710 (N_6710,N_4814,N_5684);
xor U6711 (N_6711,N_5851,N_4989);
or U6712 (N_6712,N_5587,N_5636);
xor U6713 (N_6713,N_4822,N_4985);
or U6714 (N_6714,N_5789,N_4917);
or U6715 (N_6715,N_5430,N_5110);
or U6716 (N_6716,N_4849,N_5422);
and U6717 (N_6717,N_5130,N_5175);
and U6718 (N_6718,N_5711,N_5334);
nor U6719 (N_6719,N_5038,N_5206);
or U6720 (N_6720,N_5792,N_5473);
nand U6721 (N_6721,N_5440,N_4884);
and U6722 (N_6722,N_5342,N_5593);
nand U6723 (N_6723,N_4914,N_4812);
or U6724 (N_6724,N_5925,N_5833);
and U6725 (N_6725,N_5606,N_5834);
xor U6726 (N_6726,N_5029,N_5974);
nand U6727 (N_6727,N_5843,N_5275);
nand U6728 (N_6728,N_5404,N_5468);
nor U6729 (N_6729,N_5641,N_5688);
or U6730 (N_6730,N_5286,N_5312);
xnor U6731 (N_6731,N_5437,N_5369);
nor U6732 (N_6732,N_5344,N_5335);
nand U6733 (N_6733,N_5211,N_5975);
xnor U6734 (N_6734,N_5633,N_4853);
or U6735 (N_6735,N_4926,N_5681);
nand U6736 (N_6736,N_5238,N_5904);
nor U6737 (N_6737,N_5472,N_5124);
and U6738 (N_6738,N_5862,N_5153);
nor U6739 (N_6739,N_5932,N_4935);
and U6740 (N_6740,N_5900,N_5212);
nand U6741 (N_6741,N_4944,N_5524);
xnor U6742 (N_6742,N_5943,N_5686);
xnor U6743 (N_6743,N_5781,N_5258);
nand U6744 (N_6744,N_5917,N_5162);
nand U6745 (N_6745,N_5713,N_5224);
or U6746 (N_6746,N_5064,N_5028);
xor U6747 (N_6747,N_5757,N_5005);
nor U6748 (N_6748,N_5236,N_5018);
xor U6749 (N_6749,N_5688,N_5761);
or U6750 (N_6750,N_4879,N_5753);
or U6751 (N_6751,N_5268,N_5368);
xnor U6752 (N_6752,N_5990,N_4834);
nand U6753 (N_6753,N_5919,N_4956);
or U6754 (N_6754,N_5052,N_5070);
or U6755 (N_6755,N_5663,N_4872);
nor U6756 (N_6756,N_5308,N_5131);
nor U6757 (N_6757,N_4839,N_5332);
nor U6758 (N_6758,N_5827,N_4925);
nand U6759 (N_6759,N_5090,N_5010);
xnor U6760 (N_6760,N_5280,N_5248);
nand U6761 (N_6761,N_5128,N_4932);
nor U6762 (N_6762,N_5778,N_5372);
nor U6763 (N_6763,N_5732,N_5017);
nor U6764 (N_6764,N_4959,N_4964);
and U6765 (N_6765,N_5313,N_5340);
xor U6766 (N_6766,N_5795,N_5478);
or U6767 (N_6767,N_5086,N_5467);
and U6768 (N_6768,N_5214,N_5175);
nand U6769 (N_6769,N_4803,N_5065);
nand U6770 (N_6770,N_5400,N_5577);
xnor U6771 (N_6771,N_5935,N_5162);
or U6772 (N_6772,N_5623,N_5591);
nor U6773 (N_6773,N_5021,N_5079);
nor U6774 (N_6774,N_5448,N_5536);
nor U6775 (N_6775,N_5703,N_4840);
or U6776 (N_6776,N_4851,N_5290);
xor U6777 (N_6777,N_5381,N_5271);
nand U6778 (N_6778,N_5645,N_4866);
nand U6779 (N_6779,N_4909,N_5292);
or U6780 (N_6780,N_4961,N_5760);
xor U6781 (N_6781,N_5133,N_5089);
or U6782 (N_6782,N_5354,N_5659);
and U6783 (N_6783,N_5403,N_5960);
nand U6784 (N_6784,N_4943,N_5616);
and U6785 (N_6785,N_5569,N_5027);
nand U6786 (N_6786,N_4962,N_5136);
nor U6787 (N_6787,N_5468,N_4859);
or U6788 (N_6788,N_5861,N_5016);
and U6789 (N_6789,N_5142,N_5245);
xor U6790 (N_6790,N_5815,N_5256);
and U6791 (N_6791,N_5927,N_5928);
or U6792 (N_6792,N_5692,N_5254);
and U6793 (N_6793,N_4834,N_5537);
xnor U6794 (N_6794,N_5953,N_5985);
xor U6795 (N_6795,N_5129,N_5759);
nor U6796 (N_6796,N_5140,N_5578);
and U6797 (N_6797,N_5969,N_5568);
or U6798 (N_6798,N_5086,N_5091);
nand U6799 (N_6799,N_4812,N_5048);
or U6800 (N_6800,N_5452,N_5612);
xnor U6801 (N_6801,N_5252,N_5041);
or U6802 (N_6802,N_5020,N_5077);
nand U6803 (N_6803,N_4933,N_5094);
xor U6804 (N_6804,N_5173,N_5536);
and U6805 (N_6805,N_5532,N_5101);
nand U6806 (N_6806,N_5940,N_5098);
xor U6807 (N_6807,N_5792,N_5406);
and U6808 (N_6808,N_5719,N_5205);
and U6809 (N_6809,N_5501,N_4984);
nand U6810 (N_6810,N_5225,N_4960);
nor U6811 (N_6811,N_5977,N_5916);
and U6812 (N_6812,N_4891,N_5821);
and U6813 (N_6813,N_5056,N_5926);
and U6814 (N_6814,N_5706,N_5450);
nor U6815 (N_6815,N_5025,N_4893);
and U6816 (N_6816,N_5753,N_5462);
or U6817 (N_6817,N_5161,N_5595);
xor U6818 (N_6818,N_5442,N_5553);
xor U6819 (N_6819,N_5298,N_5890);
nor U6820 (N_6820,N_5585,N_4900);
nor U6821 (N_6821,N_5185,N_5740);
xor U6822 (N_6822,N_4845,N_4801);
nand U6823 (N_6823,N_5932,N_4877);
and U6824 (N_6824,N_5034,N_5642);
or U6825 (N_6825,N_5760,N_4962);
nand U6826 (N_6826,N_5668,N_5103);
xnor U6827 (N_6827,N_5087,N_5533);
or U6828 (N_6828,N_5744,N_4809);
nand U6829 (N_6829,N_4859,N_5369);
and U6830 (N_6830,N_4849,N_5624);
or U6831 (N_6831,N_5915,N_4801);
and U6832 (N_6832,N_5760,N_5354);
or U6833 (N_6833,N_5723,N_5391);
and U6834 (N_6834,N_4947,N_5652);
xnor U6835 (N_6835,N_5979,N_4894);
xnor U6836 (N_6836,N_4872,N_5229);
nor U6837 (N_6837,N_5784,N_5293);
and U6838 (N_6838,N_4811,N_5996);
nand U6839 (N_6839,N_5164,N_5309);
nor U6840 (N_6840,N_5820,N_5479);
or U6841 (N_6841,N_4946,N_5783);
or U6842 (N_6842,N_5154,N_4987);
nand U6843 (N_6843,N_5869,N_5806);
xor U6844 (N_6844,N_5248,N_5460);
nor U6845 (N_6845,N_5062,N_4868);
or U6846 (N_6846,N_5805,N_4941);
nand U6847 (N_6847,N_5324,N_5049);
or U6848 (N_6848,N_5115,N_5159);
nand U6849 (N_6849,N_4839,N_5420);
and U6850 (N_6850,N_5095,N_5730);
or U6851 (N_6851,N_5352,N_4911);
and U6852 (N_6852,N_5186,N_5630);
and U6853 (N_6853,N_5415,N_5423);
nor U6854 (N_6854,N_5808,N_5055);
or U6855 (N_6855,N_4978,N_5836);
nand U6856 (N_6856,N_5732,N_5636);
or U6857 (N_6857,N_5357,N_5095);
nor U6858 (N_6858,N_5892,N_5911);
or U6859 (N_6859,N_4883,N_4902);
or U6860 (N_6860,N_5087,N_5916);
and U6861 (N_6861,N_5320,N_5550);
or U6862 (N_6862,N_5171,N_4946);
nand U6863 (N_6863,N_4849,N_5377);
or U6864 (N_6864,N_5920,N_5717);
nor U6865 (N_6865,N_5220,N_5194);
or U6866 (N_6866,N_5525,N_5179);
xor U6867 (N_6867,N_5434,N_5165);
and U6868 (N_6868,N_5075,N_4811);
or U6869 (N_6869,N_5332,N_5629);
xnor U6870 (N_6870,N_5116,N_4940);
nand U6871 (N_6871,N_5554,N_5222);
and U6872 (N_6872,N_5610,N_5333);
xnor U6873 (N_6873,N_5217,N_5001);
or U6874 (N_6874,N_5102,N_4973);
and U6875 (N_6875,N_5778,N_4987);
nor U6876 (N_6876,N_5596,N_5101);
nand U6877 (N_6877,N_5921,N_5197);
or U6878 (N_6878,N_5094,N_5709);
nand U6879 (N_6879,N_4915,N_5317);
and U6880 (N_6880,N_5377,N_5335);
nor U6881 (N_6881,N_5161,N_5209);
and U6882 (N_6882,N_4985,N_5813);
or U6883 (N_6883,N_5627,N_5696);
or U6884 (N_6884,N_5724,N_4959);
or U6885 (N_6885,N_5137,N_5850);
and U6886 (N_6886,N_5583,N_5193);
xnor U6887 (N_6887,N_5616,N_5961);
nor U6888 (N_6888,N_4923,N_4811);
nand U6889 (N_6889,N_5667,N_5892);
xnor U6890 (N_6890,N_5354,N_5055);
and U6891 (N_6891,N_5143,N_5869);
nand U6892 (N_6892,N_5325,N_5305);
or U6893 (N_6893,N_5728,N_5977);
nand U6894 (N_6894,N_4890,N_5123);
nand U6895 (N_6895,N_5454,N_4962);
xor U6896 (N_6896,N_5014,N_5592);
or U6897 (N_6897,N_5139,N_5770);
nor U6898 (N_6898,N_5168,N_5764);
xnor U6899 (N_6899,N_5945,N_5910);
and U6900 (N_6900,N_5878,N_5318);
nor U6901 (N_6901,N_5880,N_5360);
nor U6902 (N_6902,N_5266,N_5031);
or U6903 (N_6903,N_5421,N_5066);
or U6904 (N_6904,N_5150,N_5978);
or U6905 (N_6905,N_5315,N_5430);
or U6906 (N_6906,N_5152,N_5790);
nor U6907 (N_6907,N_5672,N_5736);
and U6908 (N_6908,N_5156,N_5971);
or U6909 (N_6909,N_5311,N_5509);
xor U6910 (N_6910,N_5106,N_5075);
nor U6911 (N_6911,N_5797,N_5605);
and U6912 (N_6912,N_4918,N_5081);
nor U6913 (N_6913,N_5036,N_5568);
xor U6914 (N_6914,N_4826,N_4848);
xor U6915 (N_6915,N_4944,N_5585);
xnor U6916 (N_6916,N_5669,N_5280);
and U6917 (N_6917,N_5789,N_5231);
nand U6918 (N_6918,N_5103,N_4978);
or U6919 (N_6919,N_4856,N_5787);
and U6920 (N_6920,N_5178,N_4916);
nand U6921 (N_6921,N_5313,N_5191);
or U6922 (N_6922,N_5139,N_5881);
nor U6923 (N_6923,N_5117,N_5992);
and U6924 (N_6924,N_5422,N_5056);
and U6925 (N_6925,N_5863,N_4803);
and U6926 (N_6926,N_5943,N_5498);
nand U6927 (N_6927,N_5716,N_5635);
xnor U6928 (N_6928,N_5576,N_5573);
and U6929 (N_6929,N_5397,N_5761);
nor U6930 (N_6930,N_5907,N_5544);
or U6931 (N_6931,N_5594,N_5245);
and U6932 (N_6932,N_5411,N_5787);
and U6933 (N_6933,N_5641,N_5276);
xnor U6934 (N_6934,N_5868,N_5385);
and U6935 (N_6935,N_5235,N_5012);
nor U6936 (N_6936,N_5253,N_4975);
or U6937 (N_6937,N_5920,N_4935);
nor U6938 (N_6938,N_5701,N_5571);
xor U6939 (N_6939,N_5581,N_5726);
xnor U6940 (N_6940,N_5959,N_5501);
nand U6941 (N_6941,N_5447,N_4995);
nand U6942 (N_6942,N_4990,N_5529);
or U6943 (N_6943,N_5294,N_4826);
xor U6944 (N_6944,N_5754,N_5259);
xnor U6945 (N_6945,N_5851,N_5519);
and U6946 (N_6946,N_5567,N_5966);
or U6947 (N_6947,N_5649,N_4809);
nor U6948 (N_6948,N_5639,N_5621);
xor U6949 (N_6949,N_4974,N_5875);
and U6950 (N_6950,N_5482,N_5190);
nand U6951 (N_6951,N_5366,N_5685);
and U6952 (N_6952,N_5538,N_5865);
nand U6953 (N_6953,N_5767,N_5507);
or U6954 (N_6954,N_5270,N_5331);
xnor U6955 (N_6955,N_5926,N_5859);
and U6956 (N_6956,N_5137,N_5028);
xor U6957 (N_6957,N_4953,N_5876);
and U6958 (N_6958,N_4885,N_5626);
xnor U6959 (N_6959,N_5127,N_4971);
nor U6960 (N_6960,N_5117,N_5874);
and U6961 (N_6961,N_5250,N_5285);
or U6962 (N_6962,N_5562,N_5641);
nor U6963 (N_6963,N_5286,N_5485);
xor U6964 (N_6964,N_5311,N_5061);
or U6965 (N_6965,N_5085,N_5341);
and U6966 (N_6966,N_5018,N_5975);
nand U6967 (N_6967,N_5926,N_4998);
or U6968 (N_6968,N_5379,N_5019);
xor U6969 (N_6969,N_5582,N_5623);
nand U6970 (N_6970,N_5356,N_5918);
nand U6971 (N_6971,N_5182,N_4980);
nor U6972 (N_6972,N_5386,N_5363);
or U6973 (N_6973,N_4897,N_5509);
and U6974 (N_6974,N_5245,N_5978);
xor U6975 (N_6975,N_5423,N_4906);
nor U6976 (N_6976,N_5524,N_5858);
and U6977 (N_6977,N_5523,N_5636);
nand U6978 (N_6978,N_5841,N_5134);
nand U6979 (N_6979,N_5731,N_5638);
nor U6980 (N_6980,N_5508,N_5834);
nor U6981 (N_6981,N_5429,N_5274);
and U6982 (N_6982,N_5481,N_5414);
nand U6983 (N_6983,N_5141,N_5535);
and U6984 (N_6984,N_5595,N_5021);
and U6985 (N_6985,N_5499,N_5648);
and U6986 (N_6986,N_4959,N_5896);
and U6987 (N_6987,N_5369,N_4860);
xnor U6988 (N_6988,N_5323,N_5273);
nand U6989 (N_6989,N_4957,N_5339);
or U6990 (N_6990,N_5280,N_5956);
xor U6991 (N_6991,N_5490,N_4814);
nor U6992 (N_6992,N_5749,N_4857);
and U6993 (N_6993,N_5966,N_5854);
nand U6994 (N_6994,N_5983,N_5459);
xnor U6995 (N_6995,N_5874,N_5694);
xnor U6996 (N_6996,N_5867,N_5369);
nor U6997 (N_6997,N_5494,N_5630);
or U6998 (N_6998,N_5150,N_4897);
nor U6999 (N_6999,N_5391,N_5261);
xnor U7000 (N_7000,N_4888,N_5436);
nand U7001 (N_7001,N_5235,N_4886);
nor U7002 (N_7002,N_5042,N_5040);
nand U7003 (N_7003,N_4874,N_5156);
or U7004 (N_7004,N_5824,N_5578);
and U7005 (N_7005,N_5908,N_5917);
or U7006 (N_7006,N_4988,N_4869);
or U7007 (N_7007,N_5884,N_5630);
nor U7008 (N_7008,N_5533,N_5579);
and U7009 (N_7009,N_4909,N_5282);
and U7010 (N_7010,N_5093,N_4852);
and U7011 (N_7011,N_5591,N_5933);
nand U7012 (N_7012,N_5367,N_5366);
nand U7013 (N_7013,N_4909,N_5779);
and U7014 (N_7014,N_5382,N_5726);
nand U7015 (N_7015,N_5995,N_4869);
xnor U7016 (N_7016,N_5504,N_5845);
xor U7017 (N_7017,N_4900,N_4877);
or U7018 (N_7018,N_5724,N_5445);
nor U7019 (N_7019,N_5844,N_4985);
xnor U7020 (N_7020,N_5657,N_5783);
or U7021 (N_7021,N_5477,N_5982);
nor U7022 (N_7022,N_5745,N_5491);
and U7023 (N_7023,N_4885,N_5875);
nand U7024 (N_7024,N_5793,N_5267);
nand U7025 (N_7025,N_4992,N_5818);
or U7026 (N_7026,N_4849,N_5655);
nor U7027 (N_7027,N_5177,N_5179);
and U7028 (N_7028,N_5973,N_5525);
nor U7029 (N_7029,N_5342,N_5652);
xnor U7030 (N_7030,N_5975,N_5250);
nand U7031 (N_7031,N_5943,N_5931);
xnor U7032 (N_7032,N_5447,N_5568);
nand U7033 (N_7033,N_5116,N_5819);
nand U7034 (N_7034,N_5093,N_4892);
xnor U7035 (N_7035,N_5439,N_4996);
nor U7036 (N_7036,N_5657,N_4915);
nand U7037 (N_7037,N_4926,N_5238);
xnor U7038 (N_7038,N_4927,N_5359);
nand U7039 (N_7039,N_5264,N_5723);
and U7040 (N_7040,N_5794,N_5847);
nor U7041 (N_7041,N_5300,N_5036);
or U7042 (N_7042,N_5005,N_4966);
and U7043 (N_7043,N_5192,N_5393);
nor U7044 (N_7044,N_5128,N_4916);
or U7045 (N_7045,N_4972,N_4830);
nand U7046 (N_7046,N_5300,N_5737);
xnor U7047 (N_7047,N_5718,N_5296);
and U7048 (N_7048,N_5575,N_5355);
or U7049 (N_7049,N_5053,N_5101);
and U7050 (N_7050,N_5675,N_5102);
nor U7051 (N_7051,N_5612,N_5208);
xnor U7052 (N_7052,N_5697,N_5215);
nand U7053 (N_7053,N_5163,N_5359);
or U7054 (N_7054,N_5367,N_5198);
nor U7055 (N_7055,N_5217,N_4903);
nor U7056 (N_7056,N_5027,N_5518);
xor U7057 (N_7057,N_4849,N_5865);
or U7058 (N_7058,N_5996,N_4875);
nand U7059 (N_7059,N_5846,N_5814);
nor U7060 (N_7060,N_5420,N_5158);
and U7061 (N_7061,N_5485,N_5085);
nand U7062 (N_7062,N_5172,N_5492);
nand U7063 (N_7063,N_5686,N_5998);
and U7064 (N_7064,N_5826,N_5011);
nor U7065 (N_7065,N_5973,N_5510);
and U7066 (N_7066,N_4833,N_5476);
or U7067 (N_7067,N_5098,N_5243);
or U7068 (N_7068,N_5340,N_5016);
and U7069 (N_7069,N_4926,N_5208);
and U7070 (N_7070,N_5791,N_5805);
or U7071 (N_7071,N_5926,N_4997);
and U7072 (N_7072,N_5387,N_5467);
or U7073 (N_7073,N_5705,N_5886);
and U7074 (N_7074,N_5123,N_5433);
nor U7075 (N_7075,N_5274,N_5602);
nand U7076 (N_7076,N_5494,N_4935);
nand U7077 (N_7077,N_5094,N_5911);
or U7078 (N_7078,N_5535,N_5942);
nand U7079 (N_7079,N_4867,N_5405);
nand U7080 (N_7080,N_4900,N_5054);
nor U7081 (N_7081,N_4917,N_5821);
or U7082 (N_7082,N_5221,N_4859);
or U7083 (N_7083,N_4927,N_5777);
nor U7084 (N_7084,N_4846,N_5499);
nor U7085 (N_7085,N_5331,N_5507);
nand U7086 (N_7086,N_4832,N_5029);
nor U7087 (N_7087,N_5639,N_5847);
nor U7088 (N_7088,N_5591,N_5353);
or U7089 (N_7089,N_5156,N_5538);
and U7090 (N_7090,N_5644,N_5185);
xnor U7091 (N_7091,N_4941,N_5710);
nand U7092 (N_7092,N_5034,N_5593);
or U7093 (N_7093,N_5699,N_5702);
and U7094 (N_7094,N_5381,N_5647);
xor U7095 (N_7095,N_5356,N_5084);
nand U7096 (N_7096,N_5412,N_5029);
xor U7097 (N_7097,N_5008,N_5382);
or U7098 (N_7098,N_5764,N_5732);
and U7099 (N_7099,N_5055,N_5683);
nor U7100 (N_7100,N_5035,N_4967);
xor U7101 (N_7101,N_5592,N_5124);
nor U7102 (N_7102,N_5176,N_4972);
or U7103 (N_7103,N_5372,N_5073);
nor U7104 (N_7104,N_5458,N_5701);
and U7105 (N_7105,N_5532,N_5277);
nor U7106 (N_7106,N_4985,N_5754);
and U7107 (N_7107,N_5833,N_5706);
xnor U7108 (N_7108,N_5678,N_4868);
nand U7109 (N_7109,N_5320,N_5846);
and U7110 (N_7110,N_5512,N_4884);
xor U7111 (N_7111,N_5430,N_5245);
nand U7112 (N_7112,N_5537,N_4887);
xnor U7113 (N_7113,N_4837,N_5936);
xor U7114 (N_7114,N_5972,N_5055);
nor U7115 (N_7115,N_5501,N_5032);
and U7116 (N_7116,N_4890,N_5138);
nand U7117 (N_7117,N_5333,N_5402);
and U7118 (N_7118,N_5702,N_5227);
xnor U7119 (N_7119,N_5255,N_5912);
nand U7120 (N_7120,N_5167,N_5556);
or U7121 (N_7121,N_5113,N_5909);
and U7122 (N_7122,N_5245,N_5639);
xor U7123 (N_7123,N_5939,N_5596);
nand U7124 (N_7124,N_5342,N_5997);
and U7125 (N_7125,N_5189,N_5694);
and U7126 (N_7126,N_4982,N_5992);
or U7127 (N_7127,N_4935,N_5213);
and U7128 (N_7128,N_5156,N_5349);
and U7129 (N_7129,N_5331,N_5532);
or U7130 (N_7130,N_5104,N_5606);
or U7131 (N_7131,N_5645,N_5508);
nor U7132 (N_7132,N_5141,N_5135);
xor U7133 (N_7133,N_5467,N_5827);
nand U7134 (N_7134,N_5642,N_5784);
xnor U7135 (N_7135,N_5465,N_4943);
xor U7136 (N_7136,N_4880,N_5375);
or U7137 (N_7137,N_4940,N_5997);
nand U7138 (N_7138,N_4932,N_5785);
nor U7139 (N_7139,N_5914,N_4961);
nand U7140 (N_7140,N_4919,N_5244);
or U7141 (N_7141,N_5190,N_5012);
xor U7142 (N_7142,N_4855,N_5762);
or U7143 (N_7143,N_5259,N_5669);
nor U7144 (N_7144,N_5905,N_5917);
nand U7145 (N_7145,N_5098,N_4834);
xnor U7146 (N_7146,N_5588,N_5880);
nor U7147 (N_7147,N_5294,N_5286);
or U7148 (N_7148,N_5418,N_4960);
or U7149 (N_7149,N_5854,N_5651);
and U7150 (N_7150,N_4866,N_5702);
xor U7151 (N_7151,N_5489,N_5907);
nor U7152 (N_7152,N_5025,N_5366);
nand U7153 (N_7153,N_5120,N_5366);
xor U7154 (N_7154,N_5235,N_5067);
nor U7155 (N_7155,N_5604,N_5442);
or U7156 (N_7156,N_5497,N_5150);
nand U7157 (N_7157,N_4911,N_5821);
and U7158 (N_7158,N_4813,N_5730);
nand U7159 (N_7159,N_5122,N_5117);
and U7160 (N_7160,N_5998,N_5999);
and U7161 (N_7161,N_5426,N_5595);
nor U7162 (N_7162,N_4937,N_5317);
or U7163 (N_7163,N_5524,N_4992);
xor U7164 (N_7164,N_5321,N_5608);
nand U7165 (N_7165,N_5383,N_5579);
nor U7166 (N_7166,N_5417,N_5289);
and U7167 (N_7167,N_5710,N_5941);
and U7168 (N_7168,N_5738,N_5854);
and U7169 (N_7169,N_4957,N_5617);
nor U7170 (N_7170,N_5428,N_5130);
and U7171 (N_7171,N_4933,N_5469);
xor U7172 (N_7172,N_5272,N_5429);
nor U7173 (N_7173,N_5299,N_5619);
nand U7174 (N_7174,N_5118,N_5444);
or U7175 (N_7175,N_5411,N_5868);
or U7176 (N_7176,N_5915,N_5646);
nor U7177 (N_7177,N_5734,N_5522);
or U7178 (N_7178,N_5237,N_5239);
nor U7179 (N_7179,N_5963,N_5898);
and U7180 (N_7180,N_5813,N_4983);
xnor U7181 (N_7181,N_5094,N_5207);
xnor U7182 (N_7182,N_5218,N_5911);
and U7183 (N_7183,N_5599,N_5462);
nor U7184 (N_7184,N_5970,N_5196);
or U7185 (N_7185,N_5081,N_5454);
or U7186 (N_7186,N_5270,N_5290);
and U7187 (N_7187,N_5223,N_4949);
nand U7188 (N_7188,N_4842,N_4820);
xnor U7189 (N_7189,N_5725,N_5887);
nor U7190 (N_7190,N_5879,N_5998);
xor U7191 (N_7191,N_5501,N_5467);
nor U7192 (N_7192,N_5557,N_5108);
nand U7193 (N_7193,N_5503,N_5733);
nor U7194 (N_7194,N_4996,N_5941);
nand U7195 (N_7195,N_5820,N_5688);
or U7196 (N_7196,N_5002,N_5813);
nor U7197 (N_7197,N_5360,N_5190);
and U7198 (N_7198,N_4864,N_5288);
xor U7199 (N_7199,N_5078,N_5653);
xnor U7200 (N_7200,N_6344,N_6085);
or U7201 (N_7201,N_6368,N_6810);
nand U7202 (N_7202,N_6103,N_6229);
xnor U7203 (N_7203,N_6953,N_6091);
xor U7204 (N_7204,N_6592,N_6398);
or U7205 (N_7205,N_6141,N_6119);
nand U7206 (N_7206,N_6595,N_6753);
xor U7207 (N_7207,N_7025,N_6076);
or U7208 (N_7208,N_6628,N_6213);
xnor U7209 (N_7209,N_6359,N_6513);
nand U7210 (N_7210,N_6916,N_6677);
and U7211 (N_7211,N_6264,N_6335);
xnor U7212 (N_7212,N_6018,N_6489);
and U7213 (N_7213,N_7115,N_6715);
and U7214 (N_7214,N_6280,N_6201);
xor U7215 (N_7215,N_6755,N_6759);
or U7216 (N_7216,N_6912,N_6388);
xnor U7217 (N_7217,N_6927,N_6737);
or U7218 (N_7218,N_6247,N_6090);
or U7219 (N_7219,N_6376,N_6886);
or U7220 (N_7220,N_7066,N_6972);
xor U7221 (N_7221,N_6714,N_6899);
nor U7222 (N_7222,N_6989,N_7079);
xnor U7223 (N_7223,N_6787,N_6722);
xor U7224 (N_7224,N_6414,N_6373);
and U7225 (N_7225,N_6517,N_6370);
nand U7226 (N_7226,N_6033,N_6296);
nor U7227 (N_7227,N_6613,N_6488);
nor U7228 (N_7228,N_6162,N_7156);
nor U7229 (N_7229,N_6256,N_6735);
and U7230 (N_7230,N_6214,N_6003);
nand U7231 (N_7231,N_7058,N_6254);
nand U7232 (N_7232,N_6220,N_6395);
or U7233 (N_7233,N_6780,N_6455);
nand U7234 (N_7234,N_6801,N_7170);
and U7235 (N_7235,N_7045,N_7103);
nor U7236 (N_7236,N_6584,N_6078);
and U7237 (N_7237,N_6881,N_6996);
nor U7238 (N_7238,N_6179,N_6960);
or U7239 (N_7239,N_6364,N_6342);
nand U7240 (N_7240,N_6406,N_6980);
nand U7241 (N_7241,N_6849,N_6295);
xor U7242 (N_7242,N_6415,N_7034);
xnor U7243 (N_7243,N_6439,N_6520);
xor U7244 (N_7244,N_6071,N_6712);
nor U7245 (N_7245,N_6203,N_6487);
and U7246 (N_7246,N_6047,N_6786);
nor U7247 (N_7247,N_6082,N_6619);
xnor U7248 (N_7248,N_6889,N_7029);
nor U7249 (N_7249,N_6000,N_6630);
nand U7250 (N_7250,N_6242,N_6668);
xor U7251 (N_7251,N_6506,N_6053);
xor U7252 (N_7252,N_6063,N_6050);
or U7253 (N_7253,N_6182,N_7085);
xor U7254 (N_7254,N_6074,N_7194);
nor U7255 (N_7255,N_6676,N_6708);
xnor U7256 (N_7256,N_6688,N_6746);
and U7257 (N_7257,N_6130,N_7087);
nor U7258 (N_7258,N_6286,N_6958);
and U7259 (N_7259,N_6404,N_6011);
nor U7260 (N_7260,N_6542,N_7027);
or U7261 (N_7261,N_6466,N_7128);
nor U7262 (N_7262,N_6667,N_6223);
nor U7263 (N_7263,N_6802,N_6217);
nand U7264 (N_7264,N_6720,N_6822);
xor U7265 (N_7265,N_6290,N_6450);
nand U7266 (N_7266,N_6829,N_6212);
and U7267 (N_7267,N_6339,N_6532);
nor U7268 (N_7268,N_6265,N_6828);
and U7269 (N_7269,N_6424,N_6156);
and U7270 (N_7270,N_7179,N_6961);
xnor U7271 (N_7271,N_6571,N_6869);
nand U7272 (N_7272,N_6811,N_6273);
nor U7273 (N_7273,N_7098,N_6436);
and U7274 (N_7274,N_7094,N_6711);
and U7275 (N_7275,N_6258,N_6686);
nand U7276 (N_7276,N_6351,N_6251);
or U7277 (N_7277,N_6921,N_6360);
or U7278 (N_7278,N_7112,N_7032);
or U7279 (N_7279,N_6888,N_7041);
or U7280 (N_7280,N_6172,N_6186);
xor U7281 (N_7281,N_6973,N_6848);
nand U7282 (N_7282,N_6901,N_6143);
nor U7283 (N_7283,N_6678,N_6238);
or U7284 (N_7284,N_6337,N_6456);
or U7285 (N_7285,N_6127,N_6747);
and U7286 (N_7286,N_6583,N_7083);
or U7287 (N_7287,N_6624,N_6627);
and U7288 (N_7288,N_6543,N_6419);
and U7289 (N_7289,N_7157,N_6800);
nand U7290 (N_7290,N_7022,N_7035);
xnor U7291 (N_7291,N_6052,N_6379);
and U7292 (N_7292,N_6476,N_7030);
nor U7293 (N_7293,N_6097,N_6654);
nor U7294 (N_7294,N_6135,N_6355);
and U7295 (N_7295,N_6197,N_6576);
nand U7296 (N_7296,N_6154,N_6494);
nor U7297 (N_7297,N_6025,N_6012);
nand U7298 (N_7298,N_6638,N_6030);
xnor U7299 (N_7299,N_6248,N_6299);
xnor U7300 (N_7300,N_7064,N_6016);
nand U7301 (N_7301,N_6940,N_6483);
nor U7302 (N_7302,N_6727,N_7180);
and U7303 (N_7303,N_6147,N_6365);
nand U7304 (N_7304,N_6323,N_6356);
nand U7305 (N_7305,N_6690,N_7114);
nor U7306 (N_7306,N_7131,N_6637);
nand U7307 (N_7307,N_7165,N_6907);
or U7308 (N_7308,N_7054,N_7100);
and U7309 (N_7309,N_6590,N_6860);
or U7310 (N_7310,N_6357,N_6581);
nand U7311 (N_7311,N_6894,N_6028);
and U7312 (N_7312,N_6228,N_6884);
and U7313 (N_7313,N_6679,N_6896);
nand U7314 (N_7314,N_6334,N_7067);
xor U7315 (N_7315,N_6783,N_6399);
nand U7316 (N_7316,N_7109,N_7120);
xnor U7317 (N_7317,N_6291,N_6305);
or U7318 (N_7318,N_6312,N_7135);
or U7319 (N_7319,N_6361,N_6675);
and U7320 (N_7320,N_6064,N_6540);
xor U7321 (N_7321,N_6683,N_6465);
nand U7322 (N_7322,N_6204,N_6403);
and U7323 (N_7323,N_6218,N_7168);
and U7324 (N_7324,N_6855,N_6577);
xnor U7325 (N_7325,N_6527,N_6648);
xnor U7326 (N_7326,N_6149,N_6748);
nand U7327 (N_7327,N_7024,N_7059);
nor U7328 (N_7328,N_6645,N_6057);
and U7329 (N_7329,N_7148,N_6726);
xor U7330 (N_7330,N_6845,N_7096);
xor U7331 (N_7331,N_6872,N_6417);
and U7332 (N_7332,N_6498,N_6326);
xnor U7333 (N_7333,N_7003,N_6526);
xnor U7334 (N_7334,N_6087,N_6636);
xor U7335 (N_7335,N_6385,N_7061);
xor U7336 (N_7336,N_6689,N_6846);
xnor U7337 (N_7337,N_6122,N_6680);
or U7338 (N_7338,N_7019,N_6084);
and U7339 (N_7339,N_6503,N_6080);
nand U7340 (N_7340,N_6695,N_6387);
nor U7341 (N_7341,N_6731,N_7012);
xnor U7342 (N_7342,N_7127,N_6758);
nor U7343 (N_7343,N_6522,N_6508);
nor U7344 (N_7344,N_7056,N_6614);
xor U7345 (N_7345,N_6175,N_6445);
or U7346 (N_7346,N_6037,N_6706);
and U7347 (N_7347,N_6210,N_6730);
nor U7348 (N_7348,N_6804,N_7046);
or U7349 (N_7349,N_7071,N_6079);
and U7350 (N_7350,N_6552,N_6655);
and U7351 (N_7351,N_7033,N_6020);
and U7352 (N_7352,N_6622,N_6556);
or U7353 (N_7353,N_6525,N_6586);
nand U7354 (N_7354,N_6566,N_6496);
nor U7355 (N_7355,N_6448,N_6168);
and U7356 (N_7356,N_6325,N_7149);
and U7357 (N_7357,N_6742,N_7076);
nor U7358 (N_7358,N_6088,N_6140);
or U7359 (N_7359,N_6844,N_6656);
or U7360 (N_7360,N_6836,N_6701);
nand U7361 (N_7361,N_6126,N_6559);
xor U7362 (N_7362,N_6152,N_6192);
or U7363 (N_7363,N_6150,N_7133);
xor U7364 (N_7364,N_6310,N_6002);
or U7365 (N_7365,N_6393,N_6809);
xnor U7366 (N_7366,N_6954,N_6460);
nand U7367 (N_7367,N_7177,N_6650);
nand U7368 (N_7368,N_6762,N_6651);
nor U7369 (N_7369,N_6382,N_7037);
and U7370 (N_7370,N_6440,N_6100);
xor U7371 (N_7371,N_6131,N_6138);
nor U7372 (N_7372,N_6600,N_6838);
xor U7373 (N_7373,N_6470,N_6641);
nand U7374 (N_7374,N_6852,N_6055);
and U7375 (N_7375,N_6502,N_7020);
nor U7376 (N_7376,N_6114,N_6826);
or U7377 (N_7377,N_6673,N_7092);
nor U7378 (N_7378,N_6536,N_6531);
or U7379 (N_7379,N_6659,N_6582);
or U7380 (N_7380,N_6544,N_6999);
or U7381 (N_7381,N_7173,N_7099);
xor U7382 (N_7382,N_6318,N_6763);
nor U7383 (N_7383,N_6573,N_6660);
xor U7384 (N_7384,N_6877,N_6512);
xor U7385 (N_7385,N_6320,N_6224);
or U7386 (N_7386,N_6952,N_6309);
and U7387 (N_7387,N_6710,N_6322);
and U7388 (N_7388,N_6473,N_6941);
nor U7389 (N_7389,N_6601,N_6068);
and U7390 (N_7390,N_7174,N_6794);
xnor U7391 (N_7391,N_7183,N_6835);
nor U7392 (N_7392,N_6813,N_6463);
nor U7393 (N_7393,N_6277,N_6437);
nand U7394 (N_7394,N_6998,N_6240);
and U7395 (N_7395,N_6430,N_6262);
or U7396 (N_7396,N_7051,N_6793);
and U7397 (N_7397,N_6239,N_6596);
and U7398 (N_7398,N_6685,N_6294);
xor U7399 (N_7399,N_6477,N_6865);
xnor U7400 (N_7400,N_6934,N_6196);
or U7401 (N_7401,N_6158,N_6332);
and U7402 (N_7402,N_7057,N_6065);
nor U7403 (N_7403,N_6891,N_6358);
nand U7404 (N_7404,N_6282,N_6013);
nand U7405 (N_7405,N_6631,N_7182);
nor U7406 (N_7406,N_7060,N_6331);
and U7407 (N_7407,N_6381,N_6259);
nor U7408 (N_7408,N_6541,N_6546);
nand U7409 (N_7409,N_6824,N_6014);
and U7410 (N_7410,N_6283,N_6871);
nand U7411 (N_7411,N_6442,N_6602);
nand U7412 (N_7412,N_6672,N_6160);
or U7413 (N_7413,N_6902,N_6340);
or U7414 (N_7414,N_6920,N_6202);
nand U7415 (N_7415,N_6165,N_6059);
and U7416 (N_7416,N_6411,N_6225);
and U7417 (N_7417,N_6107,N_6607);
nor U7418 (N_7418,N_6657,N_6198);
nand U7419 (N_7419,N_6336,N_6724);
nand U7420 (N_7420,N_6303,N_7078);
and U7421 (N_7421,N_6412,N_7086);
and U7422 (N_7422,N_7063,N_7158);
nand U7423 (N_7423,N_6338,N_7090);
nor U7424 (N_7424,N_7105,N_6092);
and U7425 (N_7425,N_6369,N_6410);
nand U7426 (N_7426,N_7018,N_6478);
xnor U7427 (N_7427,N_7073,N_6752);
nand U7428 (N_7428,N_7088,N_6729);
xor U7429 (N_7429,N_6244,N_7132);
nand U7430 (N_7430,N_6146,N_6408);
nand U7431 (N_7431,N_6977,N_6497);
nand U7432 (N_7432,N_6964,N_6132);
nand U7433 (N_7433,N_6549,N_6567);
xor U7434 (N_7434,N_7040,N_6444);
and U7435 (N_7435,N_6563,N_6618);
or U7436 (N_7436,N_6741,N_7069);
or U7437 (N_7437,N_6620,N_6537);
nor U7438 (N_7438,N_6908,N_6775);
xnor U7439 (N_7439,N_6771,N_7050);
or U7440 (N_7440,N_6278,N_6216);
and U7441 (N_7441,N_6554,N_6950);
nand U7442 (N_7442,N_6640,N_6528);
nand U7443 (N_7443,N_6593,N_6979);
nand U7444 (N_7444,N_6211,N_6102);
xnor U7445 (N_7445,N_6188,N_6591);
and U7446 (N_7446,N_7044,N_7139);
or U7447 (N_7447,N_7187,N_7017);
nand U7448 (N_7448,N_6276,N_6261);
and U7449 (N_7449,N_6313,N_6386);
nand U7450 (N_7450,N_6236,N_6518);
nand U7451 (N_7451,N_6300,N_6096);
and U7452 (N_7452,N_6231,N_6015);
nor U7453 (N_7453,N_6568,N_7163);
nor U7454 (N_7454,N_6986,N_6603);
nand U7455 (N_7455,N_6257,N_6461);
xnor U7456 (N_7456,N_7125,N_6093);
and U7457 (N_7457,N_6446,N_7191);
nand U7458 (N_7458,N_6148,N_6694);
xor U7459 (N_7459,N_6633,N_6232);
xnor U7460 (N_7460,N_7185,N_7146);
and U7461 (N_7461,N_6129,N_6482);
xor U7462 (N_7462,N_7038,N_6709);
nand U7463 (N_7463,N_6199,N_6378);
and U7464 (N_7464,N_7002,N_7042);
or U7465 (N_7465,N_6022,N_6545);
nand U7466 (N_7466,N_6565,N_6062);
nor U7467 (N_7467,N_6017,N_7097);
or U7468 (N_7468,N_6981,N_7113);
or U7469 (N_7469,N_6519,N_6652);
xnor U7470 (N_7470,N_6523,N_6451);
xnor U7471 (N_7471,N_6426,N_6995);
nand U7472 (N_7472,N_7172,N_6562);
or U7473 (N_7473,N_6390,N_6904);
xor U7474 (N_7474,N_6992,N_6302);
xor U7475 (N_7475,N_6459,N_7147);
or U7476 (N_7476,N_6761,N_6665);
and U7477 (N_7477,N_6279,N_6974);
xor U7478 (N_7478,N_7021,N_6985);
or U7479 (N_7479,N_7048,N_6782);
or U7480 (N_7480,N_6432,N_6433);
or U7481 (N_7481,N_7186,N_6825);
and U7482 (N_7482,N_7145,N_6895);
xor U7483 (N_7483,N_6144,N_6321);
nand U7484 (N_7484,N_6384,N_7001);
or U7485 (N_7485,N_6330,N_7000);
or U7486 (N_7486,N_6749,N_7026);
or U7487 (N_7487,N_6831,N_7196);
nor U7488 (N_7488,N_6698,N_6948);
and U7489 (N_7489,N_6550,N_6341);
nand U7490 (N_7490,N_6910,N_7062);
or U7491 (N_7491,N_6863,N_6687);
and U7492 (N_7492,N_7028,N_6452);
xor U7493 (N_7493,N_6599,N_6073);
xor U7494 (N_7494,N_6756,N_7192);
or U7495 (N_7495,N_7124,N_7108);
xnor U7496 (N_7496,N_6113,N_6867);
and U7497 (N_7497,N_6288,N_6789);
or U7498 (N_7498,N_7198,N_7195);
nand U7499 (N_7499,N_6642,N_6589);
and U7500 (N_7500,N_6161,N_6915);
and U7501 (N_7501,N_6447,N_6314);
nand U7502 (N_7502,N_6926,N_6371);
nand U7503 (N_7503,N_6925,N_7118);
xor U7504 (N_7504,N_6971,N_6306);
nor U7505 (N_7505,N_6875,N_6049);
or U7506 (N_7506,N_7080,N_6474);
xnor U7507 (N_7507,N_6389,N_7084);
nor U7508 (N_7508,N_6058,N_6486);
or U7509 (N_7509,N_6994,N_6784);
nor U7510 (N_7510,N_6693,N_6221);
xor U7511 (N_7511,N_7193,N_6555);
and U7512 (N_7512,N_6873,N_6969);
xnor U7513 (N_7513,N_6343,N_6151);
nand U7514 (N_7514,N_7167,N_6109);
or U7515 (N_7515,N_6598,N_6887);
nor U7516 (N_7516,N_7091,N_6352);
nand U7517 (N_7517,N_6798,N_6612);
nand U7518 (N_7518,N_6274,N_6287);
xor U7519 (N_7519,N_6548,N_6048);
and U7520 (N_7520,N_6778,N_6345);
xor U7521 (N_7521,N_6350,N_6529);
or U7522 (N_7522,N_6621,N_6180);
nand U7523 (N_7523,N_6250,N_6785);
xnor U7524 (N_7524,N_6883,N_6515);
nor U7525 (N_7525,N_6070,N_6796);
and U7526 (N_7526,N_6851,N_6010);
xor U7527 (N_7527,N_6733,N_6744);
or U7528 (N_7528,N_6234,N_6157);
or U7529 (N_7529,N_6167,N_6123);
nand U7530 (N_7530,N_7136,N_6978);
nor U7531 (N_7531,N_6159,N_7104);
and U7532 (N_7532,N_6435,N_6346);
or U7533 (N_7533,N_6609,N_6383);
or U7534 (N_7534,N_7082,N_6409);
nor U7535 (N_7535,N_7175,N_6434);
xnor U7536 (N_7536,N_6538,N_6500);
or U7537 (N_7537,N_6133,N_6504);
xnor U7538 (N_7538,N_7110,N_6072);
and U7539 (N_7539,N_6990,N_6604);
or U7540 (N_7540,N_6769,N_6768);
xnor U7541 (N_7541,N_6056,N_6653);
nand U7542 (N_7542,N_6880,N_7164);
or U7543 (N_7543,N_6284,N_6237);
xnor U7544 (N_7544,N_6524,N_6243);
and U7545 (N_7545,N_6416,N_7006);
or U7546 (N_7546,N_6843,N_6441);
and U7547 (N_7547,N_6083,N_6469);
nor U7548 (N_7548,N_6616,N_6821);
and U7549 (N_7549,N_6428,N_6900);
nor U7550 (N_7550,N_6658,N_6935);
and U7551 (N_7551,N_6751,N_7169);
xnor U7552 (N_7552,N_6205,N_7152);
nand U7553 (N_7553,N_7111,N_7137);
nand U7554 (N_7554,N_6081,N_6166);
and U7555 (N_7555,N_6479,N_6551);
or U7556 (N_7556,N_6490,N_6089);
and U7557 (N_7557,N_6570,N_6209);
nor U7558 (N_7558,N_6249,N_7039);
nor U7559 (N_7559,N_6632,N_6105);
nand U7560 (N_7560,N_6454,N_6405);
nor U7561 (N_7561,N_6190,N_6847);
and U7562 (N_7562,N_6840,N_6298);
nor U7563 (N_7563,N_7130,N_6193);
and U7564 (N_7564,N_6818,N_6670);
or U7565 (N_7565,N_6795,N_6625);
or U7566 (N_7566,N_6575,N_6557);
nand U7567 (N_7567,N_6868,N_6580);
xnor U7568 (N_7568,N_6375,N_6951);
nand U7569 (N_7569,N_6098,N_6699);
and U7570 (N_7570,N_6219,N_6363);
nor U7571 (N_7571,N_6206,N_6413);
and U7572 (N_7572,N_6307,N_6245);
and U7573 (N_7573,N_6772,N_6928);
nand U7574 (N_7574,N_6970,N_6707);
and U7575 (N_7575,N_6757,N_6293);
nor U7576 (N_7576,N_6955,N_7049);
or U7577 (N_7577,N_6115,N_6850);
xor U7578 (N_7578,N_6647,N_7072);
or U7579 (N_7579,N_6181,N_6959);
and U7580 (N_7580,N_6853,N_6732);
xnor U7581 (N_7581,N_6233,N_6719);
nor U7582 (N_7582,N_6832,N_7117);
or U7583 (N_7583,N_6521,N_6270);
xnor U7584 (N_7584,N_6713,N_6418);
nor U7585 (N_7585,N_7009,N_6882);
nor U7586 (N_7586,N_6539,N_6226);
and U7587 (N_7587,N_6745,N_7055);
nor U7588 (N_7588,N_6136,N_6480);
nor U7589 (N_7589,N_6776,N_6507);
and U7590 (N_7590,N_6574,N_6036);
nand U7591 (N_7591,N_6856,N_6919);
and U7592 (N_7592,N_6572,N_6696);
nand U7593 (N_7593,N_6449,N_7166);
nand U7594 (N_7594,N_6178,N_7023);
nand U7595 (N_7595,N_6317,N_6924);
nand U7596 (N_7596,N_6215,N_6530);
xnor U7597 (N_7597,N_6605,N_6932);
nand U7598 (N_7598,N_6579,N_6560);
or U7599 (N_7599,N_6608,N_6681);
nor U7600 (N_7600,N_7171,N_6892);
or U7601 (N_7601,N_6792,N_6101);
or U7602 (N_7602,N_7123,N_6866);
or U7603 (N_7603,N_6421,N_6791);
and U7604 (N_7604,N_6173,N_6993);
nand U7605 (N_7605,N_6060,N_6615);
nand U7606 (N_7606,N_6464,N_7181);
nor U7607 (N_7607,N_6492,N_6534);
or U7608 (N_7608,N_6760,N_6807);
or U7609 (N_7609,N_6965,N_7119);
or U7610 (N_7610,N_6635,N_6266);
nor U7611 (N_7611,N_6061,N_6754);
nor U7612 (N_7612,N_6661,N_6235);
nand U7613 (N_7613,N_6118,N_6914);
and U7614 (N_7614,N_7074,N_6725);
xnor U7615 (N_7615,N_6626,N_6922);
or U7616 (N_7616,N_6984,N_6134);
xnor U7617 (N_7617,N_6585,N_6040);
nand U7618 (N_7618,N_7015,N_7184);
xor U7619 (N_7619,N_6968,N_6879);
nand U7620 (N_7620,N_6275,N_6644);
nor U7621 (N_7621,N_6606,N_6425);
nor U7622 (N_7622,N_6738,N_6142);
nor U7623 (N_7623,N_6594,N_6086);
nor U7624 (N_7624,N_6671,N_6740);
or U7625 (N_7625,N_6703,N_6035);
and U7626 (N_7626,N_6643,N_6443);
nor U7627 (N_7627,N_6019,N_7155);
or U7628 (N_7628,N_6718,N_6943);
or U7629 (N_7629,N_7016,N_7197);
xnor U7630 (N_7630,N_6112,N_6044);
and U7631 (N_7631,N_7154,N_6353);
xor U7632 (N_7632,N_6377,N_6816);
xor U7633 (N_7633,N_6702,N_6401);
nand U7634 (N_7634,N_6770,N_6367);
and U7635 (N_7635,N_6111,N_7011);
or U7636 (N_7636,N_6032,N_6790);
and U7637 (N_7637,N_6046,N_6864);
and U7638 (N_7638,N_6402,N_7161);
nor U7639 (N_7639,N_6842,N_6553);
nand U7640 (N_7640,N_6669,N_6145);
and U7641 (N_7641,N_6819,N_6285);
xnor U7642 (N_7642,N_7010,N_6422);
and U7643 (N_7643,N_6649,N_7178);
or U7644 (N_7644,N_6155,N_6929);
or U7645 (N_7645,N_6913,N_6820);
and U7646 (N_7646,N_6903,N_6194);
xor U7647 (N_7647,N_6862,N_6110);
xnor U7648 (N_7648,N_7116,N_6024);
nor U7649 (N_7649,N_6253,N_7134);
nor U7650 (N_7650,N_6876,N_6094);
nor U7651 (N_7651,N_6949,N_6806);
xnor U7652 (N_7652,N_6005,N_6930);
or U7653 (N_7653,N_6991,N_7190);
or U7654 (N_7654,N_6429,N_6983);
nand U7655 (N_7655,N_6918,N_6372);
nand U7656 (N_7656,N_6324,N_6420);
nor U7657 (N_7657,N_6045,N_6639);
or U7658 (N_7658,N_6269,N_6348);
xor U7659 (N_7659,N_6475,N_6739);
nor U7660 (N_7660,N_6610,N_6982);
and U7661 (N_7661,N_6963,N_6031);
and U7662 (N_7662,N_6817,N_7142);
or U7663 (N_7663,N_6128,N_7176);
and U7664 (N_7664,N_6859,N_6117);
or U7665 (N_7665,N_6734,N_6308);
and U7666 (N_7666,N_6195,N_6834);
or U7667 (N_7667,N_6116,N_7068);
nand U7668 (N_7668,N_6774,N_6962);
and U7669 (N_7669,N_7121,N_6623);
nand U7670 (N_7670,N_6797,N_6808);
nor U7671 (N_7671,N_6684,N_6297);
or U7672 (N_7672,N_6137,N_6120);
xor U7673 (N_7673,N_6893,N_6588);
xor U7674 (N_7674,N_7093,N_6458);
or U7675 (N_7675,N_6750,N_7159);
xnor U7676 (N_7676,N_6861,N_6124);
nor U7677 (N_7677,N_7122,N_6779);
nor U7678 (N_7678,N_6717,N_6485);
and U7679 (N_7679,N_6857,N_7070);
nand U7680 (N_7680,N_6077,N_6987);
xor U7681 (N_7681,N_6027,N_6301);
xnor U7682 (N_7682,N_6423,N_6457);
xnor U7683 (N_7683,N_6788,N_6937);
nand U7684 (N_7684,N_6890,N_6905);
nor U7685 (N_7685,N_6564,N_6975);
and U7686 (N_7686,N_6042,N_6260);
nor U7687 (N_7687,N_7081,N_6281);
xor U7688 (N_7688,N_6467,N_6394);
nand U7689 (N_7689,N_6292,N_6736);
or U7690 (N_7690,N_6106,N_6617);
and U7691 (N_7691,N_6646,N_6870);
and U7692 (N_7692,N_6333,N_6252);
and U7693 (N_7693,N_6885,N_6374);
and U7694 (N_7694,N_6004,N_6629);
or U7695 (N_7695,N_6509,N_6805);
nor U7696 (N_7696,N_6666,N_6716);
nor U7697 (N_7697,N_6812,N_7107);
and U7698 (N_7698,N_7089,N_6823);
xnor U7699 (N_7699,N_6946,N_6104);
or U7700 (N_7700,N_6007,N_6505);
nand U7701 (N_7701,N_6453,N_6597);
nand U7702 (N_7702,N_6674,N_6174);
or U7703 (N_7703,N_6267,N_6263);
nor U7704 (N_7704,N_6705,N_6664);
nor U7705 (N_7705,N_6501,N_7047);
xor U7706 (N_7706,N_6272,N_6139);
or U7707 (N_7707,N_6697,N_7160);
nand U7708 (N_7708,N_7008,N_6316);
nand U7709 (N_7709,N_6164,N_6945);
and U7710 (N_7710,N_6909,N_6944);
and U7711 (N_7711,N_6397,N_6976);
or U7712 (N_7712,N_7065,N_6815);
nand U7713 (N_7713,N_6327,N_7007);
nor U7714 (N_7714,N_6578,N_7005);
or U7715 (N_7715,N_6936,N_6183);
or U7716 (N_7716,N_7014,N_6029);
xnor U7717 (N_7717,N_6516,N_6773);
xnor U7718 (N_7718,N_7153,N_6906);
nor U7719 (N_7719,N_6827,N_6108);
and U7720 (N_7720,N_6177,N_6966);
nor U7721 (N_7721,N_6427,N_6765);
and U7722 (N_7722,N_6391,N_6184);
nor U7723 (N_7723,N_6163,N_6311);
or U7724 (N_7724,N_7151,N_6878);
nor U7725 (N_7725,N_6481,N_6099);
xnor U7726 (N_7726,N_6329,N_6533);
nand U7727 (N_7727,N_6006,N_6069);
xor U7728 (N_7728,N_6230,N_6511);
xor U7729 (N_7729,N_7144,N_6034);
xnor U7730 (N_7730,N_6728,N_6535);
nand U7731 (N_7731,N_7126,N_7199);
or U7732 (N_7732,N_6957,N_6704);
nor U7733 (N_7733,N_6366,N_6858);
or U7734 (N_7734,N_6051,N_6938);
xor U7735 (N_7735,N_6988,N_7101);
and U7736 (N_7736,N_6066,N_6043);
or U7737 (N_7737,N_6917,N_6207);
nand U7738 (N_7738,N_6169,N_7043);
nor U7739 (N_7739,N_6255,N_7188);
nand U7740 (N_7740,N_6392,N_6021);
or U7741 (N_7741,N_6227,N_6997);
or U7742 (N_7742,N_6095,N_6246);
and U7743 (N_7743,N_6743,N_6200);
nand U7744 (N_7744,N_6799,N_6484);
xor U7745 (N_7745,N_7102,N_6723);
nor U7746 (N_7746,N_6561,N_7150);
xnor U7747 (N_7747,N_7075,N_6764);
nand U7748 (N_7748,N_7189,N_6289);
and U7749 (N_7749,N_6008,N_6191);
nor U7750 (N_7750,N_6939,N_6777);
xor U7751 (N_7751,N_6125,N_6241);
nand U7752 (N_7752,N_6803,N_7138);
xor U7753 (N_7753,N_6185,N_6328);
xor U7754 (N_7754,N_6897,N_6001);
or U7755 (N_7755,N_6781,N_6026);
xor U7756 (N_7756,N_6569,N_6472);
nand U7757 (N_7757,N_6839,N_6067);
and U7758 (N_7758,N_6942,N_6766);
or U7759 (N_7759,N_6023,N_6471);
nand U7760 (N_7760,N_7095,N_6315);
xor U7761 (N_7761,N_7052,N_6956);
and U7762 (N_7762,N_6304,N_6967);
xor U7763 (N_7763,N_6431,N_6407);
nor U7764 (N_7764,N_6841,N_6438);
and U7765 (N_7765,N_6268,N_6222);
nand U7766 (N_7766,N_6558,N_6187);
or U7767 (N_7767,N_6039,N_6176);
nor U7768 (N_7768,N_6491,N_6499);
nand U7769 (N_7769,N_6208,N_6692);
or U7770 (N_7770,N_7013,N_6931);
nand U7771 (N_7771,N_6462,N_6400);
xor U7772 (N_7772,N_6691,N_6611);
nor U7773 (N_7773,N_6319,N_6923);
nand U7774 (N_7774,N_6547,N_7143);
and U7775 (N_7775,N_6354,N_6349);
nor U7776 (N_7776,N_7004,N_7077);
or U7777 (N_7777,N_7141,N_6830);
xnor U7778 (N_7778,N_6767,N_6153);
nand U7779 (N_7779,N_6396,N_7140);
or U7780 (N_7780,N_6271,N_7036);
or U7781 (N_7781,N_6189,N_6468);
nand U7782 (N_7782,N_6510,N_6898);
nor U7783 (N_7783,N_6700,N_6587);
nand U7784 (N_7784,N_6362,N_6837);
or U7785 (N_7785,N_6682,N_6833);
nor U7786 (N_7786,N_6171,N_6347);
nor U7787 (N_7787,N_6911,N_6663);
and U7788 (N_7788,N_6874,N_7162);
or U7789 (N_7789,N_6947,N_6933);
and U7790 (N_7790,N_6170,N_6662);
nand U7791 (N_7791,N_6380,N_7129);
nand U7792 (N_7792,N_6038,N_6041);
or U7793 (N_7793,N_7106,N_7031);
or U7794 (N_7794,N_6075,N_6009);
and U7795 (N_7795,N_6493,N_6054);
or U7796 (N_7796,N_6854,N_6721);
and U7797 (N_7797,N_6121,N_7053);
xor U7798 (N_7798,N_6514,N_6634);
or U7799 (N_7799,N_6814,N_6495);
or U7800 (N_7800,N_6526,N_6573);
and U7801 (N_7801,N_6284,N_7064);
and U7802 (N_7802,N_6889,N_7113);
xnor U7803 (N_7803,N_6155,N_6619);
and U7804 (N_7804,N_6703,N_7183);
or U7805 (N_7805,N_7046,N_6064);
or U7806 (N_7806,N_6305,N_6574);
nand U7807 (N_7807,N_6798,N_6421);
and U7808 (N_7808,N_6340,N_6576);
xnor U7809 (N_7809,N_6264,N_6691);
and U7810 (N_7810,N_6805,N_6912);
nor U7811 (N_7811,N_6961,N_6342);
nor U7812 (N_7812,N_6847,N_6319);
nor U7813 (N_7813,N_6655,N_7102);
xnor U7814 (N_7814,N_6007,N_6449);
and U7815 (N_7815,N_6614,N_6688);
and U7816 (N_7816,N_6884,N_6139);
nand U7817 (N_7817,N_6318,N_6042);
nand U7818 (N_7818,N_7004,N_6513);
and U7819 (N_7819,N_6666,N_6769);
or U7820 (N_7820,N_6885,N_6939);
nor U7821 (N_7821,N_6890,N_6077);
nor U7822 (N_7822,N_6710,N_6836);
and U7823 (N_7823,N_6561,N_6699);
nand U7824 (N_7824,N_6905,N_6446);
xnor U7825 (N_7825,N_6869,N_6080);
nand U7826 (N_7826,N_6000,N_6618);
or U7827 (N_7827,N_6191,N_6901);
nand U7828 (N_7828,N_6337,N_6453);
and U7829 (N_7829,N_6408,N_6018);
or U7830 (N_7830,N_6724,N_6943);
xnor U7831 (N_7831,N_6351,N_6142);
xnor U7832 (N_7832,N_6068,N_6671);
nand U7833 (N_7833,N_7191,N_6503);
nand U7834 (N_7834,N_7087,N_7063);
xnor U7835 (N_7835,N_6862,N_6780);
nor U7836 (N_7836,N_6334,N_7075);
nor U7837 (N_7837,N_6831,N_6661);
nor U7838 (N_7838,N_6143,N_6690);
nand U7839 (N_7839,N_6454,N_6769);
and U7840 (N_7840,N_7095,N_6352);
or U7841 (N_7841,N_6200,N_6692);
nor U7842 (N_7842,N_6121,N_6979);
xor U7843 (N_7843,N_7114,N_6644);
xor U7844 (N_7844,N_6026,N_6545);
nand U7845 (N_7845,N_7043,N_6512);
and U7846 (N_7846,N_6229,N_6500);
or U7847 (N_7847,N_6125,N_6621);
nand U7848 (N_7848,N_6714,N_6413);
or U7849 (N_7849,N_6255,N_6661);
nor U7850 (N_7850,N_6446,N_6027);
nor U7851 (N_7851,N_6478,N_6750);
or U7852 (N_7852,N_6162,N_6318);
xnor U7853 (N_7853,N_7075,N_6460);
and U7854 (N_7854,N_6199,N_6452);
xor U7855 (N_7855,N_6515,N_6049);
xnor U7856 (N_7856,N_6488,N_6920);
nand U7857 (N_7857,N_7095,N_7190);
xor U7858 (N_7858,N_6185,N_6773);
and U7859 (N_7859,N_7098,N_6797);
or U7860 (N_7860,N_6317,N_6438);
and U7861 (N_7861,N_6712,N_6861);
nand U7862 (N_7862,N_6016,N_6051);
nand U7863 (N_7863,N_7076,N_6893);
or U7864 (N_7864,N_6708,N_6246);
nor U7865 (N_7865,N_6364,N_6257);
or U7866 (N_7866,N_6582,N_6507);
and U7867 (N_7867,N_6497,N_6472);
nor U7868 (N_7868,N_6184,N_6204);
or U7869 (N_7869,N_6453,N_6394);
xnor U7870 (N_7870,N_6309,N_6041);
or U7871 (N_7871,N_6925,N_6548);
nand U7872 (N_7872,N_6033,N_6607);
nor U7873 (N_7873,N_6800,N_6598);
nor U7874 (N_7874,N_7046,N_6098);
nor U7875 (N_7875,N_6797,N_6740);
nand U7876 (N_7876,N_6868,N_6842);
and U7877 (N_7877,N_6850,N_6449);
nand U7878 (N_7878,N_6427,N_7122);
and U7879 (N_7879,N_6810,N_6724);
nor U7880 (N_7880,N_6681,N_7020);
or U7881 (N_7881,N_6430,N_6660);
nand U7882 (N_7882,N_6878,N_6014);
nor U7883 (N_7883,N_6517,N_6961);
or U7884 (N_7884,N_6420,N_6679);
or U7885 (N_7885,N_6416,N_6342);
nand U7886 (N_7886,N_6210,N_6762);
and U7887 (N_7887,N_7064,N_6655);
and U7888 (N_7888,N_6363,N_6518);
nor U7889 (N_7889,N_6041,N_6729);
nor U7890 (N_7890,N_6046,N_6368);
xor U7891 (N_7891,N_7096,N_6390);
and U7892 (N_7892,N_6902,N_6226);
nand U7893 (N_7893,N_6843,N_6303);
nand U7894 (N_7894,N_7054,N_6247);
nand U7895 (N_7895,N_6813,N_6055);
nor U7896 (N_7896,N_6768,N_6035);
or U7897 (N_7897,N_6644,N_6959);
xor U7898 (N_7898,N_7175,N_7198);
xor U7899 (N_7899,N_6046,N_6381);
and U7900 (N_7900,N_6653,N_6587);
or U7901 (N_7901,N_6011,N_6670);
or U7902 (N_7902,N_6772,N_6258);
and U7903 (N_7903,N_6221,N_6877);
and U7904 (N_7904,N_7105,N_6724);
xnor U7905 (N_7905,N_6537,N_6178);
nand U7906 (N_7906,N_6189,N_6063);
and U7907 (N_7907,N_6783,N_6628);
or U7908 (N_7908,N_6011,N_6746);
and U7909 (N_7909,N_6598,N_6372);
xnor U7910 (N_7910,N_6536,N_6925);
xor U7911 (N_7911,N_6474,N_6464);
nor U7912 (N_7912,N_7046,N_6646);
nor U7913 (N_7913,N_7173,N_6944);
xnor U7914 (N_7914,N_7139,N_6721);
nand U7915 (N_7915,N_6841,N_6773);
nor U7916 (N_7916,N_6035,N_7068);
nand U7917 (N_7917,N_6647,N_6857);
nor U7918 (N_7918,N_6827,N_6828);
or U7919 (N_7919,N_6248,N_6442);
nand U7920 (N_7920,N_6326,N_6740);
xor U7921 (N_7921,N_6268,N_6855);
xnor U7922 (N_7922,N_6204,N_6089);
xor U7923 (N_7923,N_6171,N_6757);
or U7924 (N_7924,N_6892,N_6455);
nand U7925 (N_7925,N_6118,N_6154);
nor U7926 (N_7926,N_6532,N_6267);
nor U7927 (N_7927,N_6076,N_6145);
xnor U7928 (N_7928,N_6984,N_6454);
or U7929 (N_7929,N_6906,N_6808);
or U7930 (N_7930,N_6337,N_7193);
or U7931 (N_7931,N_6868,N_6089);
xor U7932 (N_7932,N_6521,N_6737);
nor U7933 (N_7933,N_7184,N_7000);
or U7934 (N_7934,N_6409,N_6122);
nand U7935 (N_7935,N_6100,N_7027);
nor U7936 (N_7936,N_6708,N_6963);
nand U7937 (N_7937,N_6895,N_6334);
nand U7938 (N_7938,N_6387,N_6860);
nand U7939 (N_7939,N_7026,N_7123);
or U7940 (N_7940,N_6001,N_6319);
nand U7941 (N_7941,N_6465,N_6474);
nor U7942 (N_7942,N_7109,N_6242);
and U7943 (N_7943,N_6896,N_6529);
nor U7944 (N_7944,N_6427,N_6356);
nand U7945 (N_7945,N_6356,N_6912);
and U7946 (N_7946,N_6490,N_6267);
xnor U7947 (N_7947,N_6218,N_6885);
nor U7948 (N_7948,N_6626,N_7081);
nor U7949 (N_7949,N_6162,N_7084);
and U7950 (N_7950,N_6055,N_7049);
xnor U7951 (N_7951,N_6028,N_6195);
nand U7952 (N_7952,N_6035,N_6887);
nand U7953 (N_7953,N_6128,N_6310);
xnor U7954 (N_7954,N_6153,N_7113);
and U7955 (N_7955,N_6350,N_7054);
nand U7956 (N_7956,N_6397,N_7180);
and U7957 (N_7957,N_6046,N_6163);
and U7958 (N_7958,N_6716,N_6725);
xnor U7959 (N_7959,N_6611,N_6705);
nand U7960 (N_7960,N_6161,N_7100);
xnor U7961 (N_7961,N_6839,N_6838);
and U7962 (N_7962,N_6851,N_7058);
or U7963 (N_7963,N_7087,N_6654);
nand U7964 (N_7964,N_6631,N_6265);
xnor U7965 (N_7965,N_6590,N_6247);
or U7966 (N_7966,N_6225,N_6136);
and U7967 (N_7967,N_7005,N_7045);
or U7968 (N_7968,N_7134,N_6349);
or U7969 (N_7969,N_7031,N_6707);
nor U7970 (N_7970,N_6021,N_7054);
or U7971 (N_7971,N_6411,N_6758);
and U7972 (N_7972,N_6491,N_6438);
and U7973 (N_7973,N_6514,N_6558);
nand U7974 (N_7974,N_6000,N_6265);
and U7975 (N_7975,N_6764,N_6212);
nor U7976 (N_7976,N_6162,N_6777);
or U7977 (N_7977,N_6852,N_6459);
nor U7978 (N_7978,N_6695,N_6915);
nand U7979 (N_7979,N_7115,N_6131);
or U7980 (N_7980,N_6806,N_6577);
or U7981 (N_7981,N_6321,N_7084);
nor U7982 (N_7982,N_6444,N_6172);
nor U7983 (N_7983,N_6954,N_6358);
or U7984 (N_7984,N_6683,N_7043);
or U7985 (N_7985,N_6094,N_6783);
xor U7986 (N_7986,N_7138,N_6459);
nor U7987 (N_7987,N_7072,N_6237);
nand U7988 (N_7988,N_6029,N_6832);
or U7989 (N_7989,N_6928,N_6461);
and U7990 (N_7990,N_6454,N_6977);
or U7991 (N_7991,N_6519,N_7142);
or U7992 (N_7992,N_6551,N_6645);
and U7993 (N_7993,N_6132,N_6163);
nor U7994 (N_7994,N_6179,N_6224);
xor U7995 (N_7995,N_6810,N_6174);
nand U7996 (N_7996,N_7079,N_6117);
nand U7997 (N_7997,N_6245,N_6660);
or U7998 (N_7998,N_6649,N_7125);
and U7999 (N_7999,N_7183,N_6528);
or U8000 (N_8000,N_7131,N_6396);
xor U8001 (N_8001,N_6497,N_6204);
and U8002 (N_8002,N_6907,N_6613);
and U8003 (N_8003,N_6767,N_6663);
nand U8004 (N_8004,N_6413,N_6288);
and U8005 (N_8005,N_6083,N_6704);
and U8006 (N_8006,N_6341,N_6403);
or U8007 (N_8007,N_6958,N_6519);
nand U8008 (N_8008,N_6951,N_6803);
nand U8009 (N_8009,N_6508,N_6334);
or U8010 (N_8010,N_6245,N_6290);
and U8011 (N_8011,N_6948,N_6230);
nor U8012 (N_8012,N_7177,N_6369);
and U8013 (N_8013,N_6562,N_6694);
xnor U8014 (N_8014,N_6631,N_6991);
nor U8015 (N_8015,N_6303,N_6599);
nor U8016 (N_8016,N_6564,N_6385);
nand U8017 (N_8017,N_6375,N_6092);
or U8018 (N_8018,N_6071,N_6462);
and U8019 (N_8019,N_7089,N_7125);
nand U8020 (N_8020,N_7161,N_6600);
or U8021 (N_8021,N_6644,N_6253);
or U8022 (N_8022,N_6756,N_7125);
nor U8023 (N_8023,N_6735,N_7165);
xnor U8024 (N_8024,N_6743,N_6739);
and U8025 (N_8025,N_6627,N_6656);
xor U8026 (N_8026,N_6140,N_6951);
nand U8027 (N_8027,N_6178,N_6852);
nand U8028 (N_8028,N_6703,N_6069);
nand U8029 (N_8029,N_6761,N_6689);
nand U8030 (N_8030,N_6932,N_6718);
xor U8031 (N_8031,N_6488,N_7007);
xor U8032 (N_8032,N_6227,N_6339);
or U8033 (N_8033,N_6693,N_6578);
nor U8034 (N_8034,N_6142,N_6468);
or U8035 (N_8035,N_6758,N_6734);
nor U8036 (N_8036,N_6832,N_6059);
nor U8037 (N_8037,N_6749,N_6833);
nand U8038 (N_8038,N_6245,N_6113);
nor U8039 (N_8039,N_6008,N_6162);
or U8040 (N_8040,N_6801,N_6104);
and U8041 (N_8041,N_6639,N_6251);
and U8042 (N_8042,N_6767,N_7142);
and U8043 (N_8043,N_7019,N_7188);
or U8044 (N_8044,N_6267,N_6325);
nand U8045 (N_8045,N_6137,N_6018);
nor U8046 (N_8046,N_6678,N_6336);
nor U8047 (N_8047,N_6143,N_6619);
nor U8048 (N_8048,N_6057,N_6464);
xnor U8049 (N_8049,N_7155,N_6837);
and U8050 (N_8050,N_6869,N_6844);
nor U8051 (N_8051,N_6263,N_6121);
xnor U8052 (N_8052,N_6090,N_6215);
xor U8053 (N_8053,N_6881,N_6277);
or U8054 (N_8054,N_6076,N_7177);
xnor U8055 (N_8055,N_6271,N_6971);
and U8056 (N_8056,N_6154,N_6837);
xnor U8057 (N_8057,N_6157,N_6711);
and U8058 (N_8058,N_6662,N_6734);
or U8059 (N_8059,N_7134,N_6857);
nor U8060 (N_8060,N_6715,N_7109);
nand U8061 (N_8061,N_6214,N_6744);
xnor U8062 (N_8062,N_7168,N_7026);
xnor U8063 (N_8063,N_6979,N_7150);
nand U8064 (N_8064,N_6343,N_7019);
nor U8065 (N_8065,N_6017,N_6935);
nand U8066 (N_8066,N_7045,N_6799);
xnor U8067 (N_8067,N_6846,N_6440);
nand U8068 (N_8068,N_6235,N_6445);
nor U8069 (N_8069,N_6948,N_7194);
or U8070 (N_8070,N_6229,N_6993);
nand U8071 (N_8071,N_6167,N_6339);
xnor U8072 (N_8072,N_7127,N_6287);
nand U8073 (N_8073,N_6488,N_6030);
nand U8074 (N_8074,N_6405,N_7024);
or U8075 (N_8075,N_7007,N_6541);
nor U8076 (N_8076,N_6064,N_6414);
nor U8077 (N_8077,N_7108,N_6172);
nand U8078 (N_8078,N_6613,N_6312);
and U8079 (N_8079,N_6284,N_6241);
xnor U8080 (N_8080,N_6859,N_6569);
xor U8081 (N_8081,N_6817,N_6476);
xnor U8082 (N_8082,N_6972,N_7172);
nand U8083 (N_8083,N_6943,N_6759);
nand U8084 (N_8084,N_6246,N_6396);
xnor U8085 (N_8085,N_6956,N_6295);
xnor U8086 (N_8086,N_6520,N_6848);
xnor U8087 (N_8087,N_6314,N_6068);
nand U8088 (N_8088,N_6371,N_6921);
and U8089 (N_8089,N_7173,N_6538);
nor U8090 (N_8090,N_6162,N_7129);
and U8091 (N_8091,N_6476,N_6622);
or U8092 (N_8092,N_6217,N_7034);
and U8093 (N_8093,N_6714,N_6363);
nor U8094 (N_8094,N_6665,N_6653);
and U8095 (N_8095,N_6793,N_6521);
nor U8096 (N_8096,N_6847,N_6983);
nand U8097 (N_8097,N_6419,N_6957);
and U8098 (N_8098,N_6118,N_6067);
nand U8099 (N_8099,N_6125,N_6272);
xor U8100 (N_8100,N_6471,N_6284);
nand U8101 (N_8101,N_7061,N_7165);
or U8102 (N_8102,N_7067,N_6915);
xor U8103 (N_8103,N_6477,N_6055);
and U8104 (N_8104,N_6753,N_6457);
or U8105 (N_8105,N_6241,N_6688);
nor U8106 (N_8106,N_7196,N_6728);
and U8107 (N_8107,N_6329,N_6424);
nor U8108 (N_8108,N_6445,N_7043);
nor U8109 (N_8109,N_6886,N_6651);
and U8110 (N_8110,N_6262,N_6568);
nand U8111 (N_8111,N_6207,N_6075);
and U8112 (N_8112,N_6582,N_6384);
nor U8113 (N_8113,N_7105,N_7012);
or U8114 (N_8114,N_6318,N_6504);
nor U8115 (N_8115,N_6838,N_6695);
and U8116 (N_8116,N_6864,N_6211);
xnor U8117 (N_8117,N_6926,N_6159);
nor U8118 (N_8118,N_7013,N_6340);
or U8119 (N_8119,N_6049,N_6622);
xnor U8120 (N_8120,N_6313,N_6621);
or U8121 (N_8121,N_6423,N_6647);
nand U8122 (N_8122,N_6714,N_7067);
nand U8123 (N_8123,N_6473,N_6505);
or U8124 (N_8124,N_6692,N_6611);
nand U8125 (N_8125,N_6298,N_6624);
xnor U8126 (N_8126,N_6417,N_6505);
xnor U8127 (N_8127,N_6633,N_6844);
or U8128 (N_8128,N_6831,N_6893);
and U8129 (N_8129,N_6336,N_7132);
xor U8130 (N_8130,N_6838,N_7155);
nand U8131 (N_8131,N_6322,N_6789);
and U8132 (N_8132,N_6221,N_6265);
xnor U8133 (N_8133,N_7027,N_6610);
nor U8134 (N_8134,N_6720,N_6469);
nand U8135 (N_8135,N_6483,N_6236);
nor U8136 (N_8136,N_6019,N_6279);
nor U8137 (N_8137,N_6634,N_7181);
xor U8138 (N_8138,N_6498,N_6401);
nor U8139 (N_8139,N_6938,N_6955);
xor U8140 (N_8140,N_6650,N_6438);
xor U8141 (N_8141,N_6002,N_6846);
nand U8142 (N_8142,N_6923,N_6931);
xnor U8143 (N_8143,N_6669,N_6367);
or U8144 (N_8144,N_6872,N_6881);
or U8145 (N_8145,N_6250,N_6360);
nand U8146 (N_8146,N_6926,N_6641);
nand U8147 (N_8147,N_6325,N_6193);
or U8148 (N_8148,N_6230,N_6489);
xor U8149 (N_8149,N_6934,N_6210);
and U8150 (N_8150,N_6892,N_7129);
or U8151 (N_8151,N_6951,N_7190);
nor U8152 (N_8152,N_6475,N_6802);
and U8153 (N_8153,N_6641,N_6507);
nand U8154 (N_8154,N_7038,N_6784);
nand U8155 (N_8155,N_7158,N_6907);
xor U8156 (N_8156,N_6527,N_7050);
xor U8157 (N_8157,N_6038,N_6259);
or U8158 (N_8158,N_6672,N_7053);
and U8159 (N_8159,N_6626,N_7033);
nand U8160 (N_8160,N_6587,N_6655);
nand U8161 (N_8161,N_6824,N_7174);
nand U8162 (N_8162,N_6582,N_6530);
and U8163 (N_8163,N_6257,N_6709);
nand U8164 (N_8164,N_6981,N_6633);
nand U8165 (N_8165,N_6391,N_6380);
and U8166 (N_8166,N_6922,N_7159);
xnor U8167 (N_8167,N_7102,N_7156);
nand U8168 (N_8168,N_6888,N_6603);
nor U8169 (N_8169,N_6928,N_6454);
nand U8170 (N_8170,N_7192,N_7109);
nand U8171 (N_8171,N_7187,N_7088);
nand U8172 (N_8172,N_6827,N_6436);
and U8173 (N_8173,N_6818,N_6166);
and U8174 (N_8174,N_6786,N_6209);
xor U8175 (N_8175,N_6901,N_6839);
nor U8176 (N_8176,N_7058,N_6506);
and U8177 (N_8177,N_6911,N_6380);
or U8178 (N_8178,N_6241,N_6315);
nor U8179 (N_8179,N_6947,N_6591);
nor U8180 (N_8180,N_6979,N_6902);
and U8181 (N_8181,N_6076,N_6433);
and U8182 (N_8182,N_6227,N_6483);
and U8183 (N_8183,N_6534,N_6299);
nand U8184 (N_8184,N_6042,N_6655);
nand U8185 (N_8185,N_6518,N_7098);
nor U8186 (N_8186,N_7088,N_6996);
and U8187 (N_8187,N_6587,N_6428);
nor U8188 (N_8188,N_6099,N_6660);
nand U8189 (N_8189,N_7080,N_6295);
and U8190 (N_8190,N_6809,N_6940);
or U8191 (N_8191,N_6553,N_7165);
and U8192 (N_8192,N_6370,N_6093);
or U8193 (N_8193,N_6915,N_7190);
nand U8194 (N_8194,N_7133,N_7037);
xnor U8195 (N_8195,N_6550,N_6907);
and U8196 (N_8196,N_6660,N_7012);
nor U8197 (N_8197,N_6330,N_6450);
nand U8198 (N_8198,N_6231,N_6087);
xor U8199 (N_8199,N_6951,N_6395);
or U8200 (N_8200,N_6273,N_7028);
and U8201 (N_8201,N_6201,N_6054);
or U8202 (N_8202,N_6614,N_6405);
nand U8203 (N_8203,N_6921,N_6772);
and U8204 (N_8204,N_6317,N_6597);
nor U8205 (N_8205,N_6655,N_6500);
nor U8206 (N_8206,N_6388,N_6236);
nor U8207 (N_8207,N_6499,N_6135);
nand U8208 (N_8208,N_6497,N_6145);
nand U8209 (N_8209,N_6313,N_6381);
and U8210 (N_8210,N_6415,N_6753);
xnor U8211 (N_8211,N_7092,N_6389);
nor U8212 (N_8212,N_6797,N_6071);
or U8213 (N_8213,N_6328,N_6972);
and U8214 (N_8214,N_6203,N_6180);
nor U8215 (N_8215,N_6267,N_6398);
nand U8216 (N_8216,N_6923,N_6276);
or U8217 (N_8217,N_6970,N_6825);
and U8218 (N_8218,N_6564,N_6728);
nor U8219 (N_8219,N_7169,N_7016);
and U8220 (N_8220,N_6046,N_6122);
xnor U8221 (N_8221,N_6260,N_7083);
nand U8222 (N_8222,N_6981,N_6546);
and U8223 (N_8223,N_7190,N_6370);
or U8224 (N_8224,N_6312,N_6208);
or U8225 (N_8225,N_6670,N_7075);
nand U8226 (N_8226,N_6623,N_6060);
nor U8227 (N_8227,N_6854,N_6722);
or U8228 (N_8228,N_6027,N_6666);
xor U8229 (N_8229,N_6734,N_6268);
xnor U8230 (N_8230,N_6266,N_7134);
xnor U8231 (N_8231,N_6137,N_7198);
or U8232 (N_8232,N_6034,N_6870);
nor U8233 (N_8233,N_6511,N_6280);
or U8234 (N_8234,N_6401,N_6505);
or U8235 (N_8235,N_7019,N_6921);
or U8236 (N_8236,N_6321,N_7185);
xnor U8237 (N_8237,N_6307,N_6061);
nor U8238 (N_8238,N_7120,N_7186);
or U8239 (N_8239,N_6148,N_6939);
xnor U8240 (N_8240,N_6351,N_6687);
and U8241 (N_8241,N_6136,N_6234);
nor U8242 (N_8242,N_6027,N_6304);
and U8243 (N_8243,N_6087,N_6734);
nor U8244 (N_8244,N_6851,N_6842);
or U8245 (N_8245,N_6424,N_6361);
nand U8246 (N_8246,N_6455,N_7126);
or U8247 (N_8247,N_6378,N_6054);
or U8248 (N_8248,N_6059,N_6753);
nand U8249 (N_8249,N_6601,N_6463);
nor U8250 (N_8250,N_7088,N_6234);
nand U8251 (N_8251,N_7060,N_6487);
nand U8252 (N_8252,N_6588,N_6879);
nor U8253 (N_8253,N_6610,N_6223);
or U8254 (N_8254,N_6000,N_6106);
or U8255 (N_8255,N_6964,N_6588);
xor U8256 (N_8256,N_6725,N_6502);
nor U8257 (N_8257,N_6009,N_6678);
xnor U8258 (N_8258,N_6024,N_7060);
and U8259 (N_8259,N_7156,N_6464);
nand U8260 (N_8260,N_6696,N_6732);
and U8261 (N_8261,N_6973,N_6335);
nor U8262 (N_8262,N_7168,N_6397);
xor U8263 (N_8263,N_6830,N_6519);
nor U8264 (N_8264,N_6757,N_6975);
and U8265 (N_8265,N_6154,N_6129);
or U8266 (N_8266,N_6457,N_6088);
xnor U8267 (N_8267,N_6410,N_6474);
or U8268 (N_8268,N_6441,N_6181);
or U8269 (N_8269,N_6180,N_6710);
and U8270 (N_8270,N_6778,N_6674);
nand U8271 (N_8271,N_6043,N_6663);
nor U8272 (N_8272,N_7161,N_7143);
xnor U8273 (N_8273,N_6976,N_6553);
xnor U8274 (N_8274,N_6685,N_6887);
xnor U8275 (N_8275,N_6731,N_6400);
and U8276 (N_8276,N_6952,N_6981);
nor U8277 (N_8277,N_6967,N_7193);
or U8278 (N_8278,N_6222,N_6324);
and U8279 (N_8279,N_6014,N_6387);
xnor U8280 (N_8280,N_6217,N_6576);
xnor U8281 (N_8281,N_6132,N_6402);
or U8282 (N_8282,N_6663,N_6722);
nor U8283 (N_8283,N_6481,N_7121);
nor U8284 (N_8284,N_6704,N_6399);
nor U8285 (N_8285,N_6549,N_6535);
nor U8286 (N_8286,N_6548,N_6250);
nand U8287 (N_8287,N_6852,N_6589);
xnor U8288 (N_8288,N_7178,N_6353);
and U8289 (N_8289,N_6731,N_7148);
xnor U8290 (N_8290,N_6471,N_6868);
nor U8291 (N_8291,N_6922,N_6770);
nor U8292 (N_8292,N_6761,N_6801);
xor U8293 (N_8293,N_6033,N_7075);
or U8294 (N_8294,N_6674,N_6436);
and U8295 (N_8295,N_6340,N_6219);
nor U8296 (N_8296,N_6049,N_6267);
nand U8297 (N_8297,N_6723,N_6226);
and U8298 (N_8298,N_7093,N_6278);
and U8299 (N_8299,N_6578,N_6674);
and U8300 (N_8300,N_7187,N_6226);
xnor U8301 (N_8301,N_6813,N_6926);
and U8302 (N_8302,N_6613,N_6392);
and U8303 (N_8303,N_6953,N_6788);
nor U8304 (N_8304,N_6406,N_6582);
xnor U8305 (N_8305,N_7042,N_6699);
and U8306 (N_8306,N_6644,N_6243);
or U8307 (N_8307,N_6478,N_6305);
and U8308 (N_8308,N_6110,N_6090);
nor U8309 (N_8309,N_6360,N_6219);
nand U8310 (N_8310,N_6449,N_6116);
nand U8311 (N_8311,N_6969,N_6124);
or U8312 (N_8312,N_6277,N_6655);
xor U8313 (N_8313,N_7063,N_6793);
or U8314 (N_8314,N_6044,N_6498);
or U8315 (N_8315,N_7011,N_6220);
or U8316 (N_8316,N_6066,N_6502);
or U8317 (N_8317,N_6896,N_6990);
nor U8318 (N_8318,N_6415,N_6770);
xnor U8319 (N_8319,N_6397,N_6236);
xnor U8320 (N_8320,N_6730,N_6044);
nand U8321 (N_8321,N_6421,N_6779);
nor U8322 (N_8322,N_6704,N_6262);
nor U8323 (N_8323,N_6017,N_7025);
nor U8324 (N_8324,N_6693,N_6720);
nor U8325 (N_8325,N_6005,N_6490);
and U8326 (N_8326,N_7028,N_6186);
nand U8327 (N_8327,N_6174,N_6811);
or U8328 (N_8328,N_6707,N_7036);
nor U8329 (N_8329,N_6704,N_6988);
or U8330 (N_8330,N_6599,N_6060);
and U8331 (N_8331,N_6944,N_7154);
xor U8332 (N_8332,N_7008,N_6168);
nand U8333 (N_8333,N_6711,N_6020);
nor U8334 (N_8334,N_7061,N_6249);
and U8335 (N_8335,N_6548,N_6011);
xor U8336 (N_8336,N_6250,N_6874);
xor U8337 (N_8337,N_7183,N_6927);
nor U8338 (N_8338,N_6809,N_7136);
xnor U8339 (N_8339,N_6670,N_6145);
xnor U8340 (N_8340,N_6089,N_7026);
nor U8341 (N_8341,N_7027,N_6170);
nor U8342 (N_8342,N_6853,N_6941);
xnor U8343 (N_8343,N_7007,N_6857);
xnor U8344 (N_8344,N_6235,N_6724);
nand U8345 (N_8345,N_6753,N_6224);
nor U8346 (N_8346,N_6001,N_6012);
xor U8347 (N_8347,N_6362,N_6288);
xor U8348 (N_8348,N_6771,N_6505);
nor U8349 (N_8349,N_6313,N_6529);
nand U8350 (N_8350,N_7024,N_6028);
nor U8351 (N_8351,N_7127,N_6708);
nor U8352 (N_8352,N_7199,N_7107);
and U8353 (N_8353,N_6560,N_6344);
and U8354 (N_8354,N_6537,N_6480);
or U8355 (N_8355,N_6516,N_6134);
nor U8356 (N_8356,N_6078,N_6128);
nand U8357 (N_8357,N_7094,N_7117);
nor U8358 (N_8358,N_6761,N_6119);
or U8359 (N_8359,N_6220,N_6998);
xnor U8360 (N_8360,N_6763,N_7067);
nor U8361 (N_8361,N_6782,N_6282);
and U8362 (N_8362,N_6255,N_6718);
nor U8363 (N_8363,N_6944,N_6580);
nor U8364 (N_8364,N_6120,N_6064);
nand U8365 (N_8365,N_6532,N_6638);
xor U8366 (N_8366,N_7132,N_6308);
and U8367 (N_8367,N_6052,N_7187);
nand U8368 (N_8368,N_6057,N_6867);
xnor U8369 (N_8369,N_7184,N_6690);
or U8370 (N_8370,N_6678,N_6292);
and U8371 (N_8371,N_6193,N_6017);
or U8372 (N_8372,N_6230,N_7005);
xor U8373 (N_8373,N_7101,N_6841);
and U8374 (N_8374,N_6183,N_6425);
xor U8375 (N_8375,N_6999,N_6273);
nand U8376 (N_8376,N_6835,N_6334);
or U8377 (N_8377,N_6068,N_7099);
nor U8378 (N_8378,N_6466,N_6626);
and U8379 (N_8379,N_7073,N_6361);
or U8380 (N_8380,N_6801,N_7150);
and U8381 (N_8381,N_7129,N_7161);
nor U8382 (N_8382,N_6592,N_6564);
nand U8383 (N_8383,N_6733,N_6908);
nand U8384 (N_8384,N_6483,N_6602);
or U8385 (N_8385,N_6214,N_6507);
nor U8386 (N_8386,N_6557,N_6965);
or U8387 (N_8387,N_6789,N_7151);
nand U8388 (N_8388,N_6593,N_6642);
or U8389 (N_8389,N_6807,N_7174);
nand U8390 (N_8390,N_7132,N_6449);
and U8391 (N_8391,N_6483,N_6942);
xor U8392 (N_8392,N_6933,N_7128);
nand U8393 (N_8393,N_6190,N_6944);
and U8394 (N_8394,N_6426,N_6684);
or U8395 (N_8395,N_6805,N_6847);
and U8396 (N_8396,N_6092,N_6320);
or U8397 (N_8397,N_6246,N_7165);
nand U8398 (N_8398,N_6301,N_7038);
nand U8399 (N_8399,N_6615,N_6013);
xnor U8400 (N_8400,N_7482,N_7812);
nor U8401 (N_8401,N_7714,N_7343);
nor U8402 (N_8402,N_8075,N_8388);
nand U8403 (N_8403,N_7425,N_8264);
nand U8404 (N_8404,N_7827,N_8300);
and U8405 (N_8405,N_8230,N_7647);
nor U8406 (N_8406,N_7729,N_7360);
and U8407 (N_8407,N_7591,N_7596);
or U8408 (N_8408,N_7270,N_8223);
nor U8409 (N_8409,N_7765,N_7892);
xnor U8410 (N_8410,N_7675,N_7580);
nor U8411 (N_8411,N_7664,N_7655);
or U8412 (N_8412,N_8181,N_7991);
nand U8413 (N_8413,N_8055,N_7217);
xor U8414 (N_8414,N_7865,N_7480);
nand U8415 (N_8415,N_7720,N_7645);
xnor U8416 (N_8416,N_8294,N_8310);
xnor U8417 (N_8417,N_8398,N_8047);
nor U8418 (N_8418,N_7553,N_8043);
or U8419 (N_8419,N_7285,N_8157);
nand U8420 (N_8420,N_8100,N_7995);
or U8421 (N_8421,N_7309,N_8184);
or U8422 (N_8422,N_8135,N_7884);
nand U8423 (N_8423,N_7815,N_7787);
nor U8424 (N_8424,N_8173,N_7736);
nor U8425 (N_8425,N_8117,N_7862);
or U8426 (N_8426,N_7273,N_7871);
xor U8427 (N_8427,N_7531,N_7274);
and U8428 (N_8428,N_8113,N_7564);
xor U8429 (N_8429,N_7872,N_7811);
xor U8430 (N_8430,N_8316,N_7939);
nor U8431 (N_8431,N_8314,N_7418);
nor U8432 (N_8432,N_7843,N_7701);
nand U8433 (N_8433,N_7784,N_8197);
nand U8434 (N_8434,N_7205,N_7735);
xnor U8435 (N_8435,N_8035,N_7746);
and U8436 (N_8436,N_7390,N_7644);
nand U8437 (N_8437,N_7696,N_8174);
and U8438 (N_8438,N_8204,N_8044);
and U8439 (N_8439,N_8021,N_7755);
nand U8440 (N_8440,N_7248,N_7369);
or U8441 (N_8441,N_7505,N_7403);
nor U8442 (N_8442,N_8238,N_7368);
or U8443 (N_8443,N_7548,N_8236);
nor U8444 (N_8444,N_8217,N_8141);
nor U8445 (N_8445,N_7534,N_7817);
or U8446 (N_8446,N_7299,N_7711);
xor U8447 (N_8447,N_8182,N_7767);
xor U8448 (N_8448,N_7640,N_7389);
nand U8449 (N_8449,N_7351,N_7912);
or U8450 (N_8450,N_7747,N_7652);
nor U8451 (N_8451,N_7972,N_7507);
nand U8452 (N_8452,N_8269,N_7778);
or U8453 (N_8453,N_7933,N_8352);
and U8454 (N_8454,N_8125,N_7410);
or U8455 (N_8455,N_8114,N_7669);
and U8456 (N_8456,N_8088,N_7326);
nor U8457 (N_8457,N_7677,N_7467);
xnor U8458 (N_8458,N_7233,N_7208);
or U8459 (N_8459,N_7211,N_8076);
xor U8460 (N_8460,N_8122,N_8304);
nor U8461 (N_8461,N_8280,N_7760);
or U8462 (N_8462,N_7257,N_7216);
or U8463 (N_8463,N_8385,N_8148);
nand U8464 (N_8464,N_8336,N_7526);
xor U8465 (N_8465,N_7894,N_7443);
nor U8466 (N_8466,N_7291,N_8396);
nand U8467 (N_8467,N_7373,N_7663);
or U8468 (N_8468,N_7569,N_7495);
xor U8469 (N_8469,N_7604,N_7335);
xor U8470 (N_8470,N_7397,N_7960);
and U8471 (N_8471,N_7286,N_7296);
xnor U8472 (N_8472,N_7959,N_7726);
and U8473 (N_8473,N_7610,N_7823);
nand U8474 (N_8474,N_7619,N_7444);
nor U8475 (N_8475,N_7454,N_7931);
xnor U8476 (N_8476,N_8134,N_7824);
and U8477 (N_8477,N_8211,N_7943);
nand U8478 (N_8478,N_7911,N_7997);
nor U8479 (N_8479,N_7998,N_7500);
nor U8480 (N_8480,N_7430,N_8357);
xor U8481 (N_8481,N_7453,N_8131);
and U8482 (N_8482,N_8030,N_8067);
or U8483 (N_8483,N_8019,N_7621);
xor U8484 (N_8484,N_7896,N_7387);
or U8485 (N_8485,N_7409,N_8079);
and U8486 (N_8486,N_7885,N_7574);
nand U8487 (N_8487,N_7268,N_7923);
xnor U8488 (N_8488,N_7856,N_8195);
nand U8489 (N_8489,N_7880,N_8218);
and U8490 (N_8490,N_7751,N_8311);
or U8491 (N_8491,N_7284,N_7733);
nand U8492 (N_8492,N_7512,N_7447);
and U8493 (N_8493,N_8288,N_8291);
or U8494 (N_8494,N_7956,N_8303);
nand U8495 (N_8495,N_7304,N_7223);
xnor U8496 (N_8496,N_8097,N_7316);
and U8497 (N_8497,N_7301,N_7928);
or U8498 (N_8498,N_7420,N_7364);
nor U8499 (N_8499,N_7897,N_8221);
or U8500 (N_8500,N_7702,N_7890);
and U8501 (N_8501,N_7637,N_7977);
nor U8502 (N_8502,N_7497,N_7445);
nand U8503 (N_8503,N_7321,N_7925);
xor U8504 (N_8504,N_7670,N_7879);
and U8505 (N_8505,N_7559,N_7340);
or U8506 (N_8506,N_8198,N_7944);
nor U8507 (N_8507,N_7877,N_7819);
nor U8508 (N_8508,N_7292,N_7816);
or U8509 (N_8509,N_7478,N_7348);
and U8510 (N_8510,N_7642,N_7620);
and U8511 (N_8511,N_7496,N_8200);
nor U8512 (N_8512,N_7535,N_7904);
and U8513 (N_8513,N_7902,N_7648);
or U8514 (N_8514,N_7875,N_7634);
nand U8515 (N_8515,N_7522,N_7305);
and U8516 (N_8516,N_7691,N_7541);
or U8517 (N_8517,N_7797,N_8234);
nand U8518 (N_8518,N_7438,N_7832);
nand U8519 (N_8519,N_7983,N_7985);
xor U8520 (N_8520,N_8123,N_8266);
nor U8521 (N_8521,N_8363,N_7465);
or U8522 (N_8522,N_8282,N_8395);
and U8523 (N_8523,N_7826,N_8175);
and U8524 (N_8524,N_7631,N_7785);
nor U8525 (N_8525,N_8187,N_7848);
and U8526 (N_8526,N_8251,N_7973);
nor U8527 (N_8527,N_7888,N_7909);
xor U8528 (N_8528,N_7560,N_7868);
nand U8529 (N_8529,N_7457,N_7716);
nand U8530 (N_8530,N_8241,N_7311);
nor U8531 (N_8531,N_8330,N_7793);
and U8532 (N_8532,N_8024,N_7250);
and U8533 (N_8533,N_7855,N_7754);
xnor U8534 (N_8534,N_7258,N_8057);
and U8535 (N_8535,N_7988,N_8128);
nand U8536 (N_8536,N_7562,N_7688);
and U8537 (N_8537,N_7431,N_8031);
nand U8538 (N_8538,N_7388,N_7382);
or U8539 (N_8539,N_8351,N_7385);
and U8540 (N_8540,N_7915,N_8028);
or U8541 (N_8541,N_8225,N_7231);
or U8542 (N_8542,N_7759,N_7525);
nor U8543 (N_8543,N_8213,N_8159);
and U8544 (N_8544,N_7448,N_8312);
xnor U8545 (N_8545,N_7969,N_8169);
nor U8546 (N_8546,N_7730,N_7324);
nor U8547 (N_8547,N_8058,N_8380);
nor U8548 (N_8548,N_8228,N_7412);
or U8549 (N_8549,N_8263,N_7656);
nand U8550 (N_8550,N_7707,N_7325);
nor U8551 (N_8551,N_8036,N_8095);
nor U8552 (N_8552,N_7671,N_8318);
or U8553 (N_8553,N_8026,N_7607);
nor U8554 (N_8554,N_8003,N_8186);
and U8555 (N_8555,N_8258,N_7623);
nor U8556 (N_8556,N_8354,N_7616);
and U8557 (N_8557,N_7719,N_8307);
xor U8558 (N_8558,N_8362,N_7563);
or U8559 (N_8559,N_7704,N_7357);
xor U8560 (N_8560,N_7243,N_8137);
or U8561 (N_8561,N_7681,N_7905);
nand U8562 (N_8562,N_8208,N_7966);
xnor U8563 (N_8563,N_7611,N_8235);
nor U8564 (N_8564,N_8015,N_7886);
xor U8565 (N_8565,N_8040,N_7481);
or U8566 (N_8566,N_7212,N_7331);
nand U8567 (N_8567,N_7201,N_7240);
and U8568 (N_8568,N_7841,N_7230);
xor U8569 (N_8569,N_7947,N_7723);
xnor U8570 (N_8570,N_7602,N_8286);
and U8571 (N_8571,N_7678,N_7399);
and U8572 (N_8572,N_7581,N_8391);
and U8573 (N_8573,N_7416,N_7408);
nand U8574 (N_8574,N_7693,N_7506);
nand U8575 (N_8575,N_8140,N_7439);
xor U8576 (N_8576,N_7502,N_8384);
xor U8577 (N_8577,N_7256,N_8147);
xnor U8578 (N_8578,N_7650,N_7770);
nand U8579 (N_8579,N_8360,N_8329);
nor U8580 (N_8580,N_8025,N_7822);
and U8581 (N_8581,N_7279,N_8038);
nand U8582 (N_8582,N_8252,N_7213);
xnor U8583 (N_8583,N_7992,N_7845);
nand U8584 (N_8584,N_7463,N_7614);
and U8585 (N_8585,N_8145,N_7520);
nor U8586 (N_8586,N_7662,N_7336);
nor U8587 (N_8587,N_8016,N_7433);
or U8588 (N_8588,N_8156,N_7910);
nor U8589 (N_8589,N_8356,N_7501);
or U8590 (N_8590,N_7471,N_7539);
nand U8591 (N_8591,N_7741,N_7833);
nand U8592 (N_8592,N_7776,N_8227);
and U8593 (N_8593,N_8377,N_7840);
xnor U8594 (N_8594,N_7202,N_7245);
and U8595 (N_8595,N_7918,N_8041);
or U8596 (N_8596,N_8254,N_8194);
nor U8597 (N_8597,N_7547,N_7781);
and U8598 (N_8598,N_8083,N_7994);
or U8599 (N_8599,N_7979,N_8054);
nand U8600 (N_8600,N_7587,N_8255);
xor U8601 (N_8601,N_8189,N_7695);
xnor U8602 (N_8602,N_8301,N_7990);
xnor U8603 (N_8603,N_7930,N_7750);
and U8604 (N_8604,N_7818,N_8283);
nor U8605 (N_8605,N_7993,N_8249);
nand U8606 (N_8606,N_7281,N_8136);
nor U8607 (N_8607,N_8344,N_7628);
or U8608 (N_8608,N_7734,N_7970);
xor U8609 (N_8609,N_7486,N_7226);
nor U8610 (N_8610,N_7363,N_7253);
nor U8611 (N_8611,N_7401,N_8371);
nand U8612 (N_8612,N_7685,N_7949);
and U8613 (N_8613,N_8144,N_8393);
xor U8614 (N_8614,N_7780,N_7901);
and U8615 (N_8615,N_7940,N_8193);
nor U8616 (N_8616,N_8034,N_7801);
nor U8617 (N_8617,N_7709,N_8081);
and U8618 (N_8618,N_8013,N_8382);
nand U8619 (N_8619,N_7287,N_8381);
xnor U8620 (N_8620,N_7362,N_7713);
nand U8621 (N_8621,N_8212,N_7828);
or U8622 (N_8622,N_7690,N_7545);
or U8623 (N_8623,N_8118,N_8115);
nand U8624 (N_8624,N_8029,N_7870);
nor U8625 (N_8625,N_8281,N_7846);
nand U8626 (N_8626,N_8052,N_7732);
or U8627 (N_8627,N_7951,N_7498);
xnor U8628 (N_8628,N_8000,N_7594);
or U8629 (N_8629,N_8306,N_8270);
nand U8630 (N_8630,N_7898,N_7272);
xnor U8631 (N_8631,N_8168,N_7706);
or U8632 (N_8632,N_8158,N_7661);
nor U8633 (N_8633,N_7267,N_7203);
or U8634 (N_8634,N_8162,N_7352);
nand U8635 (N_8635,N_7579,N_7224);
nor U8636 (N_8636,N_8246,N_8317);
or U8637 (N_8637,N_8290,N_8060);
xnor U8638 (N_8638,N_7882,N_7347);
xor U8639 (N_8639,N_8061,N_7330);
xnor U8640 (N_8640,N_8196,N_8348);
or U8641 (N_8641,N_8143,N_8203);
or U8642 (N_8642,N_8121,N_8201);
and U8643 (N_8643,N_7612,N_7752);
or U8644 (N_8644,N_7679,N_7974);
xor U8645 (N_8645,N_8279,N_8365);
xnor U8646 (N_8646,N_8185,N_7237);
nor U8647 (N_8647,N_8315,N_8350);
nand U8648 (N_8648,N_8099,N_8065);
nor U8649 (N_8649,N_7391,N_7585);
or U8650 (N_8650,N_7963,N_7798);
or U8651 (N_8651,N_8272,N_7519);
nor U8652 (N_8652,N_8338,N_8179);
xnor U8653 (N_8653,N_7544,N_7766);
xor U8654 (N_8654,N_8229,N_7314);
nand U8655 (N_8655,N_8216,N_8242);
nand U8656 (N_8656,N_7289,N_7262);
nand U8657 (N_8657,N_7370,N_8092);
and U8658 (N_8658,N_7852,N_8210);
nand U8659 (N_8659,N_7978,N_8205);
nor U8660 (N_8660,N_7383,N_7996);
or U8661 (N_8661,N_8289,N_8256);
nor U8662 (N_8662,N_7555,N_7375);
xor U8663 (N_8663,N_8299,N_7698);
and U8664 (N_8664,N_7473,N_7715);
or U8665 (N_8665,N_8151,N_7295);
nor U8666 (N_8666,N_7227,N_8383);
xor U8667 (N_8667,N_7571,N_7204);
xnor U8668 (N_8668,N_7639,N_8394);
or U8669 (N_8669,N_8325,N_7532);
nand U8670 (N_8670,N_7572,N_7934);
nor U8671 (N_8671,N_8071,N_8109);
xor U8672 (N_8672,N_8042,N_7633);
xnor U8673 (N_8673,N_8326,N_7850);
xor U8674 (N_8674,N_7967,N_7239);
nand U8675 (N_8675,N_8359,N_8374);
nand U8676 (N_8676,N_7400,N_7813);
nand U8677 (N_8677,N_7586,N_8014);
xnor U8678 (N_8678,N_7860,N_7209);
and U8679 (N_8679,N_7965,N_8002);
and U8680 (N_8680,N_7748,N_7788);
nor U8681 (N_8681,N_7867,N_7568);
and U8682 (N_8682,N_7861,N_7883);
xnor U8683 (N_8683,N_7821,N_7700);
xnor U8684 (N_8684,N_7451,N_8341);
xor U8685 (N_8685,N_7926,N_7603);
nor U8686 (N_8686,N_7953,N_7459);
nor U8687 (N_8687,N_7774,N_7406);
or U8688 (N_8688,N_8078,N_7873);
or U8689 (N_8689,N_7789,N_8387);
nand U8690 (N_8690,N_7524,N_7312);
and U8691 (N_8691,N_7415,N_7627);
nor U8692 (N_8692,N_7651,N_8008);
or U8693 (N_8693,N_7269,N_7942);
nand U8694 (N_8694,N_7777,N_8101);
and U8695 (N_8695,N_8285,N_7405);
nand U8696 (N_8696,N_7315,N_7680);
xor U8697 (N_8697,N_8305,N_7427);
nor U8698 (N_8698,N_7206,N_8392);
and U8699 (N_8699,N_7657,N_7533);
nand U8700 (N_8700,N_7643,N_7288);
and U8701 (N_8701,N_7232,N_7407);
nand U8702 (N_8702,N_7440,N_7460);
nand U8703 (N_8703,N_8370,N_8215);
or U8704 (N_8704,N_7329,N_8389);
or U8705 (N_8705,N_7863,N_8199);
nor U8706 (N_8706,N_7508,N_7929);
nor U8707 (N_8707,N_7356,N_8274);
or U8708 (N_8708,N_7374,N_7493);
and U8709 (N_8709,N_7950,N_8074);
and U8710 (N_8710,N_8265,N_8068);
xnor U8711 (N_8711,N_7844,N_7462);
nand U8712 (N_8712,N_8261,N_7744);
xnor U8713 (N_8713,N_8005,N_7659);
nor U8714 (N_8714,N_8232,N_7999);
nor U8715 (N_8715,N_7836,N_7298);
xnor U8716 (N_8716,N_7536,N_8161);
or U8717 (N_8717,N_7276,N_7874);
nor U8718 (N_8718,N_7542,N_7676);
or U8719 (N_8719,N_7479,N_7492);
xor U8720 (N_8720,N_7540,N_8007);
or U8721 (N_8721,N_7938,N_7386);
and U8722 (N_8722,N_7738,N_7455);
and U8723 (N_8723,N_8347,N_7592);
nor U8724 (N_8724,N_7263,N_8226);
nor U8725 (N_8725,N_7957,N_8017);
nor U8726 (N_8726,N_7491,N_7570);
xor U8727 (N_8727,N_7372,N_8009);
nor U8728 (N_8728,N_8048,N_8051);
and U8729 (N_8729,N_7899,N_7799);
nand U8730 (N_8730,N_7674,N_7831);
or U8731 (N_8731,N_7626,N_7772);
nand U8732 (N_8732,N_7724,N_8006);
nand U8733 (N_8733,N_8166,N_7740);
and U8734 (N_8734,N_8018,N_8105);
or U8735 (N_8735,N_8271,N_7499);
and U8736 (N_8736,N_8070,N_7353);
nand U8737 (N_8737,N_7476,N_7477);
and U8738 (N_8738,N_7487,N_7756);
nand U8739 (N_8739,N_8262,N_7251);
and U8740 (N_8740,N_7921,N_8292);
nand U8741 (N_8741,N_8331,N_7668);
or U8742 (N_8742,N_7834,N_8372);
and U8743 (N_8743,N_7300,N_8219);
or U8744 (N_8744,N_8032,N_7814);
and U8745 (N_8745,N_7332,N_7641);
nand U8746 (N_8746,N_7989,N_7710);
xnor U8747 (N_8747,N_7945,N_8124);
xor U8748 (N_8748,N_7878,N_8077);
nor U8749 (N_8749,N_8257,N_7342);
xor U8750 (N_8750,N_7549,N_8176);
xnor U8751 (N_8751,N_7638,N_7266);
or U8752 (N_8752,N_7396,N_7567);
or U8753 (N_8753,N_7866,N_8190);
nor U8754 (N_8754,N_8375,N_7725);
or U8755 (N_8755,N_7809,N_8379);
and U8756 (N_8756,N_7590,N_8328);
nor U8757 (N_8757,N_7936,N_7413);
xor U8758 (N_8758,N_7229,N_8103);
nor U8759 (N_8759,N_7275,N_7829);
or U8760 (N_8760,N_7575,N_7379);
xor U8761 (N_8761,N_7582,N_7820);
or U8762 (N_8762,N_7552,N_7359);
nor U8763 (N_8763,N_7712,N_8090);
and U8764 (N_8764,N_7728,N_7908);
nand U8765 (N_8765,N_7837,N_7442);
nor U8766 (N_8766,N_7987,N_8037);
nor U8767 (N_8767,N_7247,N_7238);
and U8768 (N_8768,N_7392,N_8165);
nand U8769 (N_8769,N_8001,N_8183);
nand U8770 (N_8770,N_8066,N_7469);
nor U8771 (N_8771,N_7470,N_7854);
xor U8772 (N_8772,N_8155,N_7763);
and U8773 (N_8773,N_7380,N_7566);
and U8774 (N_8774,N_8020,N_7265);
or U8775 (N_8775,N_7743,N_8239);
xnor U8776 (N_8776,N_7920,N_7830);
xor U8777 (N_8777,N_7429,N_7538);
or U8778 (N_8778,N_7509,N_7919);
nor U8779 (N_8779,N_7742,N_8321);
nor U8780 (N_8780,N_8399,N_7761);
or U8781 (N_8781,N_7434,N_7242);
nand U8782 (N_8782,N_7806,N_7718);
and U8783 (N_8783,N_8087,N_8327);
or U8784 (N_8784,N_8233,N_8237);
or U8785 (N_8785,N_7791,N_7218);
or U8786 (N_8786,N_8033,N_8177);
and U8787 (N_8787,N_8098,N_7876);
and U8788 (N_8788,N_7595,N_8010);
or U8789 (N_8789,N_7722,N_8146);
xor U8790 (N_8790,N_7807,N_7293);
or U8791 (N_8791,N_7513,N_7334);
nand U8792 (N_8792,N_8376,N_7895);
nor U8793 (N_8793,N_8231,N_8171);
nor U8794 (N_8794,N_8064,N_7606);
and U8795 (N_8795,N_8346,N_8069);
or U8796 (N_8796,N_7749,N_7757);
nor U8797 (N_8797,N_8053,N_8106);
xor U8798 (N_8798,N_8340,N_7906);
nand U8799 (N_8799,N_7252,N_7589);
nand U8800 (N_8800,N_7510,N_7984);
nand U8801 (N_8801,N_7318,N_7423);
or U8802 (N_8802,N_8191,N_7782);
nor U8803 (N_8803,N_7394,N_8277);
nand U8804 (N_8804,N_7219,N_7236);
and U8805 (N_8805,N_8085,N_7446);
xnor U8806 (N_8806,N_7869,N_8308);
or U8807 (N_8807,N_7697,N_8366);
nand U8808 (N_8808,N_7344,N_7689);
and U8809 (N_8809,N_8022,N_8102);
xor U8810 (N_8810,N_7283,N_7328);
and U8811 (N_8811,N_7786,N_7411);
xnor U8812 (N_8812,N_8367,N_7598);
nand U8813 (N_8813,N_8378,N_8170);
or U8814 (N_8814,N_8345,N_7417);
nand U8815 (N_8815,N_7800,N_7851);
nor U8816 (N_8816,N_7600,N_7672);
nand U8817 (N_8817,N_7558,N_7319);
xor U8818 (N_8818,N_7658,N_7366);
or U8819 (N_8819,N_7775,N_8214);
nand U8820 (N_8820,N_8086,N_8104);
and U8821 (N_8821,N_7864,N_7666);
nand U8822 (N_8822,N_7608,N_7805);
xor U8823 (N_8823,N_7618,N_7764);
or U8824 (N_8824,N_7737,N_8084);
xnor U8825 (N_8825,N_7573,N_8260);
xor U8826 (N_8826,N_7249,N_7523);
xor U8827 (N_8827,N_8355,N_8045);
nand U8828 (N_8828,N_8163,N_7835);
xor U8829 (N_8829,N_7521,N_7297);
nor U8830 (N_8830,N_8295,N_8004);
and U8831 (N_8831,N_8220,N_8172);
or U8832 (N_8832,N_7900,N_8164);
or U8833 (N_8833,N_8333,N_7264);
nor U8834 (N_8834,N_8335,N_8116);
nand U8835 (N_8835,N_7584,N_7527);
nor U8836 (N_8836,N_8108,N_7424);
nand U8837 (N_8837,N_7597,N_7753);
nand U8838 (N_8838,N_7654,N_7794);
nand U8839 (N_8839,N_7768,N_8337);
and U8840 (N_8840,N_7982,N_7282);
xnor U8841 (N_8841,N_8142,N_7913);
or U8842 (N_8842,N_8302,N_7528);
xor U8843 (N_8843,N_7808,N_7889);
nor U8844 (N_8844,N_7530,N_7629);
or U8845 (N_8845,N_7511,N_8245);
xnor U8846 (N_8846,N_7739,N_7474);
or U8847 (N_8847,N_7727,N_8082);
and U8848 (N_8848,N_8150,N_7692);
nand U8849 (N_8849,N_7485,N_8153);
nand U8850 (N_8850,N_7302,N_8273);
or U8851 (N_8851,N_8309,N_7546);
xnor U8852 (N_8852,N_7769,N_7458);
and U8853 (N_8853,N_8152,N_8358);
or U8854 (N_8854,N_7980,N_7986);
or U8855 (N_8855,N_7244,N_7683);
and U8856 (N_8856,N_7414,N_8119);
or U8857 (N_8857,N_7916,N_7557);
nand U8858 (N_8858,N_7554,N_8343);
nor U8859 (N_8859,N_7200,N_8132);
nor U8860 (N_8860,N_7941,N_8222);
or U8861 (N_8861,N_8240,N_7207);
nand U8862 (N_8862,N_7853,N_7367);
nor U8863 (N_8863,N_8243,N_7849);
nand U8864 (N_8864,N_7622,N_7441);
and U8865 (N_8865,N_7613,N_7503);
and U8866 (N_8866,N_7461,N_8178);
xor U8867 (N_8867,N_8276,N_7857);
xor U8868 (N_8868,N_8322,N_8253);
xnor U8869 (N_8869,N_7903,N_7721);
nand U8870 (N_8870,N_7422,N_7588);
nor U8871 (N_8871,N_7346,N_7402);
or U8872 (N_8872,N_7483,N_8342);
or U8873 (N_8873,N_7398,N_7636);
xor U8874 (N_8874,N_7703,N_7303);
or U8875 (N_8875,N_7235,N_8209);
nand U8876 (N_8876,N_7665,N_7395);
and U8877 (N_8877,N_7307,N_7593);
nor U8878 (N_8878,N_7432,N_8129);
nand U8879 (N_8879,N_8323,N_8247);
or U8880 (N_8880,N_8386,N_8091);
nor U8881 (N_8881,N_7518,N_7537);
and U8882 (N_8882,N_7341,N_8046);
and U8883 (N_8883,N_7327,N_8039);
nand U8884 (N_8884,N_8050,N_8324);
nor U8885 (N_8885,N_7731,N_8096);
or U8886 (N_8886,N_8160,N_8130);
nand U8887 (N_8887,N_7682,N_7514);
xor U8888 (N_8888,N_7339,N_8207);
nor U8889 (N_8889,N_7371,N_7630);
and U8890 (N_8890,N_7466,N_7234);
nand U8891 (N_8891,N_8334,N_8397);
or U8892 (N_8892,N_7624,N_7260);
or U8893 (N_8893,N_7290,N_7881);
nand U8894 (N_8894,N_8206,N_7646);
or U8895 (N_8895,N_7948,N_8127);
nor U8896 (N_8896,N_7294,N_7556);
nor U8897 (N_8897,N_7333,N_8133);
nand U8898 (N_8898,N_7419,N_7708);
and U8899 (N_8899,N_7225,N_7228);
or U8900 (N_8900,N_8361,N_7436);
nand U8901 (N_8901,N_7421,N_8368);
nor U8902 (N_8902,N_8332,N_7393);
xor U8903 (N_8903,N_7758,N_8012);
nor U8904 (N_8904,N_8056,N_7802);
or U8905 (N_8905,N_7745,N_7215);
and U8906 (N_8906,N_7261,N_7475);
xor U8907 (N_8907,N_7625,N_7529);
xor U8908 (N_8908,N_7271,N_8275);
or U8909 (N_8909,N_7358,N_7345);
nor U8910 (N_8910,N_8250,N_7660);
xor U8911 (N_8911,N_7705,N_7796);
nor U8912 (N_8912,N_7426,N_7278);
nor U8913 (N_8913,N_7935,N_8111);
xnor U8914 (N_8914,N_8011,N_8167);
xnor U8915 (N_8915,N_7504,N_7803);
or U8916 (N_8916,N_7783,N_7576);
or U8917 (N_8917,N_7214,N_7717);
and U8918 (N_8918,N_7927,N_8073);
or U8919 (N_8919,N_7241,N_7858);
and U8920 (N_8920,N_7338,N_8284);
or U8921 (N_8921,N_7381,N_7551);
nand U8922 (N_8922,N_8080,N_8319);
nand U8923 (N_8923,N_8112,N_7838);
and U8924 (N_8924,N_8059,N_8353);
nor U8925 (N_8925,N_7976,N_8364);
nor U8926 (N_8926,N_8313,N_7349);
or U8927 (N_8927,N_7435,N_8107);
nand U8928 (N_8928,N_7859,N_8268);
or U8929 (N_8929,N_8120,N_8297);
nand U8930 (N_8930,N_7914,N_7561);
nand U8931 (N_8931,N_7583,N_7847);
nor U8932 (N_8932,N_8202,N_7635);
and U8933 (N_8933,N_8089,N_7893);
or U8934 (N_8934,N_7667,N_7221);
nand U8935 (N_8935,N_7810,N_7981);
xnor U8936 (N_8936,N_7254,N_8390);
nor U8937 (N_8937,N_7952,N_7355);
nor U8938 (N_8938,N_7404,N_7792);
nand U8939 (N_8939,N_7464,N_8267);
nor U8940 (N_8940,N_8180,N_8062);
xor U8941 (N_8941,N_7350,N_7322);
nor U8942 (N_8942,N_8093,N_7632);
xnor U8943 (N_8943,N_8154,N_7220);
xnor U8944 (N_8944,N_7790,N_8278);
or U8945 (N_8945,N_7699,N_7246);
and U8946 (N_8946,N_7891,N_7578);
and U8947 (N_8947,N_8298,N_7694);
and U8948 (N_8948,N_7222,N_8192);
and U8949 (N_8949,N_8224,N_7384);
nor U8950 (N_8950,N_8320,N_7773);
or U8951 (N_8951,N_7255,N_7932);
xor U8952 (N_8952,N_7320,N_8023);
or U8953 (N_8953,N_7489,N_7308);
nand U8954 (N_8954,N_7494,N_7565);
or U8955 (N_8955,N_7771,N_7490);
or U8956 (N_8956,N_8138,N_7964);
xor U8957 (N_8957,N_7449,N_7515);
and U8958 (N_8958,N_8139,N_7599);
xnor U8959 (N_8959,N_7825,N_7968);
xor U8960 (N_8960,N_7577,N_7310);
and U8961 (N_8961,N_7543,N_8049);
nor U8962 (N_8962,N_7687,N_7361);
xnor U8963 (N_8963,N_7317,N_8188);
or U8964 (N_8964,N_8369,N_7452);
and U8965 (N_8965,N_8126,N_7354);
nand U8966 (N_8966,N_7450,N_7484);
xnor U8967 (N_8967,N_7946,N_7280);
or U8968 (N_8968,N_7516,N_7955);
nand U8969 (N_8969,N_7259,N_7922);
xnor U8970 (N_8970,N_7210,N_8244);
and U8971 (N_8971,N_7488,N_8287);
or U8972 (N_8972,N_7468,N_7306);
or U8973 (N_8973,N_7795,N_7617);
nor U8974 (N_8974,N_8027,N_8094);
nand U8975 (N_8975,N_7365,N_7842);
xor U8976 (N_8976,N_7958,N_7653);
xor U8977 (N_8977,N_7615,N_7609);
nand U8978 (N_8978,N_8072,N_8349);
or U8979 (N_8979,N_7961,N_7937);
nor U8980 (N_8980,N_7971,N_7472);
nor U8981 (N_8981,N_8149,N_7376);
nand U8982 (N_8982,N_7601,N_8110);
and U8983 (N_8983,N_7887,N_8293);
nor U8984 (N_8984,N_7779,N_8339);
nor U8985 (N_8985,N_8259,N_7277);
and U8986 (N_8986,N_7456,N_7517);
or U8987 (N_8987,N_7954,N_7962);
xnor U8988 (N_8988,N_7605,N_7323);
nand U8989 (N_8989,N_8373,N_7762);
xor U8990 (N_8990,N_7686,N_7684);
and U8991 (N_8991,N_7550,N_7437);
nand U8992 (N_8992,N_7377,N_7428);
nand U8993 (N_8993,N_7378,N_8296);
xnor U8994 (N_8994,N_7907,N_7924);
or U8995 (N_8995,N_8248,N_7673);
and U8996 (N_8996,N_7804,N_7649);
or U8997 (N_8997,N_8063,N_7975);
nor U8998 (N_8998,N_7313,N_7839);
xor U8999 (N_8999,N_7337,N_7917);
nor U9000 (N_9000,N_8019,N_8122);
or U9001 (N_9001,N_7610,N_7703);
and U9002 (N_9002,N_7488,N_8394);
nor U9003 (N_9003,N_7733,N_8351);
xnor U9004 (N_9004,N_7629,N_7275);
xnor U9005 (N_9005,N_7320,N_7855);
nand U9006 (N_9006,N_8092,N_7960);
xnor U9007 (N_9007,N_7799,N_7286);
or U9008 (N_9008,N_8155,N_7620);
nor U9009 (N_9009,N_7672,N_8158);
xnor U9010 (N_9010,N_8083,N_8131);
nor U9011 (N_9011,N_7501,N_7948);
and U9012 (N_9012,N_7848,N_8339);
xnor U9013 (N_9013,N_8305,N_7791);
nor U9014 (N_9014,N_8318,N_8383);
nor U9015 (N_9015,N_7559,N_7978);
xor U9016 (N_9016,N_8303,N_7975);
nand U9017 (N_9017,N_8223,N_7719);
and U9018 (N_9018,N_8173,N_7344);
xor U9019 (N_9019,N_8151,N_7406);
nor U9020 (N_9020,N_7409,N_7374);
xor U9021 (N_9021,N_7470,N_7936);
xor U9022 (N_9022,N_8121,N_7854);
xnor U9023 (N_9023,N_7965,N_8229);
and U9024 (N_9024,N_7710,N_8326);
xor U9025 (N_9025,N_8291,N_7881);
nand U9026 (N_9026,N_7275,N_8018);
and U9027 (N_9027,N_7631,N_7692);
nand U9028 (N_9028,N_7291,N_7410);
and U9029 (N_9029,N_7802,N_7990);
xor U9030 (N_9030,N_8172,N_7855);
nor U9031 (N_9031,N_7809,N_7208);
xnor U9032 (N_9032,N_7856,N_7610);
xnor U9033 (N_9033,N_8155,N_7576);
nor U9034 (N_9034,N_7606,N_7941);
and U9035 (N_9035,N_7760,N_8172);
xor U9036 (N_9036,N_8097,N_7738);
nor U9037 (N_9037,N_8019,N_8174);
nand U9038 (N_9038,N_7664,N_7744);
and U9039 (N_9039,N_7727,N_7601);
nand U9040 (N_9040,N_7258,N_7536);
and U9041 (N_9041,N_8262,N_7573);
nand U9042 (N_9042,N_7470,N_7598);
nand U9043 (N_9043,N_7752,N_7285);
or U9044 (N_9044,N_8246,N_7981);
nor U9045 (N_9045,N_8349,N_7748);
or U9046 (N_9046,N_8213,N_8321);
or U9047 (N_9047,N_7882,N_8053);
and U9048 (N_9048,N_7507,N_7496);
and U9049 (N_9049,N_7834,N_8369);
or U9050 (N_9050,N_8348,N_7945);
or U9051 (N_9051,N_7782,N_7515);
nand U9052 (N_9052,N_7544,N_7443);
nor U9053 (N_9053,N_7206,N_7701);
nor U9054 (N_9054,N_7231,N_7961);
xnor U9055 (N_9055,N_7526,N_7883);
nor U9056 (N_9056,N_8314,N_7394);
nand U9057 (N_9057,N_8084,N_7370);
xor U9058 (N_9058,N_8388,N_7598);
nand U9059 (N_9059,N_7372,N_8343);
or U9060 (N_9060,N_7961,N_7254);
nor U9061 (N_9061,N_7851,N_8227);
nand U9062 (N_9062,N_7773,N_7420);
nand U9063 (N_9063,N_8047,N_7696);
and U9064 (N_9064,N_7925,N_7230);
nor U9065 (N_9065,N_8285,N_7592);
xnor U9066 (N_9066,N_7681,N_7838);
and U9067 (N_9067,N_8119,N_7355);
nand U9068 (N_9068,N_8090,N_7297);
and U9069 (N_9069,N_7996,N_8216);
or U9070 (N_9070,N_7528,N_7482);
nand U9071 (N_9071,N_7591,N_8253);
nand U9072 (N_9072,N_7758,N_8030);
xnor U9073 (N_9073,N_7920,N_8132);
and U9074 (N_9074,N_7564,N_7775);
or U9075 (N_9075,N_8084,N_7644);
nor U9076 (N_9076,N_7358,N_7850);
nor U9077 (N_9077,N_7606,N_8243);
xnor U9078 (N_9078,N_8166,N_8071);
nand U9079 (N_9079,N_8101,N_8359);
xnor U9080 (N_9080,N_8157,N_8103);
nor U9081 (N_9081,N_8021,N_8069);
nor U9082 (N_9082,N_8168,N_7984);
xor U9083 (N_9083,N_7624,N_7855);
xnor U9084 (N_9084,N_7825,N_7798);
nor U9085 (N_9085,N_7655,N_8302);
or U9086 (N_9086,N_7246,N_7468);
xor U9087 (N_9087,N_8075,N_7928);
nand U9088 (N_9088,N_7603,N_7915);
xnor U9089 (N_9089,N_8147,N_7416);
nand U9090 (N_9090,N_8257,N_7623);
or U9091 (N_9091,N_7627,N_7560);
nand U9092 (N_9092,N_8040,N_7891);
or U9093 (N_9093,N_7559,N_7804);
nor U9094 (N_9094,N_7824,N_7838);
and U9095 (N_9095,N_8051,N_7435);
or U9096 (N_9096,N_8388,N_7821);
or U9097 (N_9097,N_8066,N_8024);
or U9098 (N_9098,N_7836,N_7205);
nand U9099 (N_9099,N_7720,N_7605);
xnor U9100 (N_9100,N_7389,N_7735);
nor U9101 (N_9101,N_7570,N_7970);
or U9102 (N_9102,N_8060,N_8144);
or U9103 (N_9103,N_8051,N_7248);
or U9104 (N_9104,N_7294,N_8124);
or U9105 (N_9105,N_8369,N_7422);
and U9106 (N_9106,N_7975,N_7697);
nand U9107 (N_9107,N_7626,N_8296);
xnor U9108 (N_9108,N_7320,N_7304);
or U9109 (N_9109,N_7500,N_7926);
or U9110 (N_9110,N_8300,N_7454);
nand U9111 (N_9111,N_8231,N_8394);
nor U9112 (N_9112,N_8048,N_7764);
xnor U9113 (N_9113,N_8274,N_8257);
xor U9114 (N_9114,N_7647,N_7740);
and U9115 (N_9115,N_8285,N_7679);
and U9116 (N_9116,N_8195,N_7578);
nand U9117 (N_9117,N_7890,N_8079);
nor U9118 (N_9118,N_7798,N_8137);
xor U9119 (N_9119,N_7457,N_7983);
xnor U9120 (N_9120,N_7968,N_8040);
xnor U9121 (N_9121,N_7937,N_8237);
nor U9122 (N_9122,N_7959,N_8070);
xnor U9123 (N_9123,N_7869,N_7473);
and U9124 (N_9124,N_7965,N_7476);
or U9125 (N_9125,N_7542,N_8047);
and U9126 (N_9126,N_7567,N_7229);
nor U9127 (N_9127,N_7757,N_7286);
xor U9128 (N_9128,N_7551,N_7568);
nand U9129 (N_9129,N_7762,N_8074);
or U9130 (N_9130,N_8114,N_7333);
and U9131 (N_9131,N_7684,N_7616);
and U9132 (N_9132,N_8099,N_7877);
and U9133 (N_9133,N_8036,N_8123);
nand U9134 (N_9134,N_7466,N_7902);
or U9135 (N_9135,N_8388,N_7589);
or U9136 (N_9136,N_8347,N_8152);
nand U9137 (N_9137,N_7853,N_7904);
and U9138 (N_9138,N_7464,N_7223);
xnor U9139 (N_9139,N_7233,N_7585);
nor U9140 (N_9140,N_8063,N_7969);
and U9141 (N_9141,N_7432,N_7480);
or U9142 (N_9142,N_8161,N_7214);
and U9143 (N_9143,N_7423,N_7525);
and U9144 (N_9144,N_7446,N_7273);
or U9145 (N_9145,N_8102,N_7598);
nand U9146 (N_9146,N_8234,N_7865);
and U9147 (N_9147,N_7633,N_8073);
or U9148 (N_9148,N_8134,N_7859);
and U9149 (N_9149,N_7875,N_8396);
or U9150 (N_9150,N_8327,N_7998);
or U9151 (N_9151,N_7871,N_8377);
or U9152 (N_9152,N_7316,N_8230);
xnor U9153 (N_9153,N_7365,N_7661);
nor U9154 (N_9154,N_7984,N_7863);
xnor U9155 (N_9155,N_7988,N_7218);
nand U9156 (N_9156,N_7727,N_7728);
nor U9157 (N_9157,N_7277,N_7931);
nor U9158 (N_9158,N_7486,N_7294);
xor U9159 (N_9159,N_7502,N_7929);
xor U9160 (N_9160,N_7884,N_7721);
nor U9161 (N_9161,N_7982,N_7708);
xor U9162 (N_9162,N_8126,N_7477);
nor U9163 (N_9163,N_7539,N_8197);
and U9164 (N_9164,N_7222,N_7778);
nand U9165 (N_9165,N_8178,N_8085);
and U9166 (N_9166,N_8379,N_7901);
or U9167 (N_9167,N_8002,N_7613);
and U9168 (N_9168,N_7388,N_8245);
and U9169 (N_9169,N_7899,N_7507);
or U9170 (N_9170,N_7491,N_7781);
nor U9171 (N_9171,N_7281,N_7582);
xnor U9172 (N_9172,N_8194,N_7800);
and U9173 (N_9173,N_7612,N_8341);
xnor U9174 (N_9174,N_7932,N_7310);
nor U9175 (N_9175,N_7332,N_8370);
nand U9176 (N_9176,N_7876,N_7974);
and U9177 (N_9177,N_7413,N_8252);
and U9178 (N_9178,N_7445,N_7771);
nand U9179 (N_9179,N_8035,N_7815);
and U9180 (N_9180,N_7423,N_7659);
nand U9181 (N_9181,N_7606,N_7664);
xnor U9182 (N_9182,N_8001,N_7649);
or U9183 (N_9183,N_7778,N_7797);
nand U9184 (N_9184,N_7438,N_8080);
nand U9185 (N_9185,N_7445,N_8130);
nor U9186 (N_9186,N_7360,N_7595);
nor U9187 (N_9187,N_7514,N_7243);
or U9188 (N_9188,N_7993,N_7890);
nand U9189 (N_9189,N_7880,N_8323);
nor U9190 (N_9190,N_7529,N_8127);
and U9191 (N_9191,N_7353,N_8134);
nor U9192 (N_9192,N_8128,N_7999);
xnor U9193 (N_9193,N_7562,N_7805);
nor U9194 (N_9194,N_7303,N_7906);
and U9195 (N_9195,N_7758,N_7854);
nor U9196 (N_9196,N_7586,N_8139);
nand U9197 (N_9197,N_7958,N_8140);
xnor U9198 (N_9198,N_7852,N_7913);
or U9199 (N_9199,N_7739,N_7768);
nand U9200 (N_9200,N_7443,N_7219);
nor U9201 (N_9201,N_8008,N_7234);
nor U9202 (N_9202,N_8005,N_7525);
xnor U9203 (N_9203,N_7793,N_7685);
nor U9204 (N_9204,N_8357,N_8023);
or U9205 (N_9205,N_7271,N_7428);
nor U9206 (N_9206,N_7721,N_7289);
nand U9207 (N_9207,N_7522,N_7836);
or U9208 (N_9208,N_8174,N_8254);
nor U9209 (N_9209,N_7628,N_7829);
nor U9210 (N_9210,N_7337,N_7681);
and U9211 (N_9211,N_8121,N_7285);
xor U9212 (N_9212,N_7480,N_7792);
nand U9213 (N_9213,N_8060,N_7211);
nor U9214 (N_9214,N_7239,N_7846);
nand U9215 (N_9215,N_7287,N_7497);
xnor U9216 (N_9216,N_7546,N_7454);
nand U9217 (N_9217,N_7898,N_7510);
xnor U9218 (N_9218,N_7471,N_8161);
nor U9219 (N_9219,N_8331,N_7307);
xor U9220 (N_9220,N_7897,N_8006);
nand U9221 (N_9221,N_7258,N_7701);
or U9222 (N_9222,N_8161,N_7405);
xnor U9223 (N_9223,N_7245,N_7574);
xnor U9224 (N_9224,N_8339,N_7850);
nand U9225 (N_9225,N_7794,N_7200);
or U9226 (N_9226,N_8328,N_7672);
nor U9227 (N_9227,N_7512,N_7710);
nand U9228 (N_9228,N_7748,N_8167);
nand U9229 (N_9229,N_7602,N_7455);
xnor U9230 (N_9230,N_8281,N_8393);
xnor U9231 (N_9231,N_7506,N_7648);
and U9232 (N_9232,N_7472,N_8286);
or U9233 (N_9233,N_7201,N_7379);
xnor U9234 (N_9234,N_7878,N_8215);
and U9235 (N_9235,N_8056,N_7353);
or U9236 (N_9236,N_8049,N_7314);
and U9237 (N_9237,N_7331,N_8001);
or U9238 (N_9238,N_8362,N_8386);
and U9239 (N_9239,N_7360,N_7653);
or U9240 (N_9240,N_8189,N_7430);
and U9241 (N_9241,N_8066,N_7691);
and U9242 (N_9242,N_8187,N_8334);
and U9243 (N_9243,N_7359,N_7738);
xnor U9244 (N_9244,N_7597,N_7665);
and U9245 (N_9245,N_7694,N_7611);
nor U9246 (N_9246,N_7837,N_7431);
nand U9247 (N_9247,N_7666,N_8163);
or U9248 (N_9248,N_7896,N_8380);
xnor U9249 (N_9249,N_8234,N_8277);
nand U9250 (N_9250,N_7808,N_8228);
nand U9251 (N_9251,N_7468,N_8067);
xnor U9252 (N_9252,N_8145,N_7943);
xor U9253 (N_9253,N_7641,N_7286);
or U9254 (N_9254,N_7815,N_7871);
or U9255 (N_9255,N_7758,N_8299);
nand U9256 (N_9256,N_7802,N_7686);
nand U9257 (N_9257,N_8196,N_8376);
and U9258 (N_9258,N_7832,N_7286);
nor U9259 (N_9259,N_8279,N_7700);
xor U9260 (N_9260,N_7204,N_7981);
nor U9261 (N_9261,N_8035,N_7289);
and U9262 (N_9262,N_7515,N_7546);
nand U9263 (N_9263,N_7949,N_8355);
nand U9264 (N_9264,N_8198,N_8293);
nor U9265 (N_9265,N_7448,N_7415);
nand U9266 (N_9266,N_7219,N_7866);
nand U9267 (N_9267,N_8280,N_7726);
or U9268 (N_9268,N_7953,N_7396);
xor U9269 (N_9269,N_8040,N_7445);
nor U9270 (N_9270,N_8114,N_8047);
xor U9271 (N_9271,N_7280,N_7861);
nand U9272 (N_9272,N_7500,N_7833);
xor U9273 (N_9273,N_7228,N_7403);
and U9274 (N_9274,N_7689,N_7928);
or U9275 (N_9275,N_7571,N_8199);
nand U9276 (N_9276,N_7575,N_8260);
xnor U9277 (N_9277,N_7840,N_8028);
or U9278 (N_9278,N_7866,N_7476);
and U9279 (N_9279,N_8362,N_7200);
nand U9280 (N_9280,N_7435,N_7951);
or U9281 (N_9281,N_7735,N_8306);
and U9282 (N_9282,N_8384,N_8191);
nor U9283 (N_9283,N_7390,N_8107);
nor U9284 (N_9284,N_8289,N_7691);
and U9285 (N_9285,N_8256,N_8363);
or U9286 (N_9286,N_7445,N_8224);
nor U9287 (N_9287,N_7369,N_8141);
xor U9288 (N_9288,N_8045,N_7228);
and U9289 (N_9289,N_8217,N_7525);
or U9290 (N_9290,N_8010,N_7962);
xnor U9291 (N_9291,N_7858,N_7901);
and U9292 (N_9292,N_8181,N_7608);
xnor U9293 (N_9293,N_8028,N_7248);
or U9294 (N_9294,N_8325,N_7287);
nand U9295 (N_9295,N_7464,N_7984);
xnor U9296 (N_9296,N_8386,N_7203);
or U9297 (N_9297,N_7643,N_7765);
nand U9298 (N_9298,N_7906,N_7334);
nor U9299 (N_9299,N_7585,N_7603);
nand U9300 (N_9300,N_7930,N_8348);
nor U9301 (N_9301,N_7402,N_8062);
nand U9302 (N_9302,N_7938,N_7724);
nand U9303 (N_9303,N_8036,N_7256);
or U9304 (N_9304,N_8250,N_7716);
or U9305 (N_9305,N_7882,N_8338);
nand U9306 (N_9306,N_8324,N_7564);
xor U9307 (N_9307,N_8047,N_7298);
nand U9308 (N_9308,N_8238,N_8349);
or U9309 (N_9309,N_7558,N_8035);
or U9310 (N_9310,N_7438,N_8043);
nand U9311 (N_9311,N_7912,N_8125);
xnor U9312 (N_9312,N_7682,N_7329);
nor U9313 (N_9313,N_7538,N_7410);
xnor U9314 (N_9314,N_7920,N_8312);
nor U9315 (N_9315,N_7349,N_7772);
nor U9316 (N_9316,N_7369,N_7568);
or U9317 (N_9317,N_7284,N_8212);
or U9318 (N_9318,N_7919,N_7511);
and U9319 (N_9319,N_7699,N_7377);
and U9320 (N_9320,N_7521,N_8200);
nor U9321 (N_9321,N_7409,N_7887);
or U9322 (N_9322,N_8230,N_7836);
and U9323 (N_9323,N_7757,N_7887);
or U9324 (N_9324,N_7223,N_8247);
and U9325 (N_9325,N_7480,N_7656);
nand U9326 (N_9326,N_7445,N_8015);
nor U9327 (N_9327,N_7357,N_7989);
and U9328 (N_9328,N_8339,N_7808);
or U9329 (N_9329,N_8334,N_7957);
xnor U9330 (N_9330,N_8162,N_8148);
nor U9331 (N_9331,N_7454,N_7582);
and U9332 (N_9332,N_8170,N_7378);
nor U9333 (N_9333,N_7322,N_7826);
and U9334 (N_9334,N_7663,N_7841);
or U9335 (N_9335,N_8282,N_7438);
and U9336 (N_9336,N_8271,N_7384);
and U9337 (N_9337,N_7598,N_7347);
and U9338 (N_9338,N_7759,N_7290);
nor U9339 (N_9339,N_7827,N_7417);
nand U9340 (N_9340,N_7360,N_8381);
xnor U9341 (N_9341,N_8099,N_7334);
and U9342 (N_9342,N_8397,N_7352);
and U9343 (N_9343,N_8137,N_7540);
or U9344 (N_9344,N_7887,N_8190);
xnor U9345 (N_9345,N_7342,N_8264);
nand U9346 (N_9346,N_7877,N_7225);
xor U9347 (N_9347,N_8276,N_7207);
and U9348 (N_9348,N_7716,N_7770);
and U9349 (N_9349,N_7545,N_7421);
xnor U9350 (N_9350,N_8318,N_7467);
and U9351 (N_9351,N_7830,N_7442);
nor U9352 (N_9352,N_7711,N_7695);
nor U9353 (N_9353,N_7817,N_7388);
xnor U9354 (N_9354,N_8228,N_7536);
nand U9355 (N_9355,N_8361,N_7415);
xnor U9356 (N_9356,N_7281,N_7389);
and U9357 (N_9357,N_7321,N_7331);
xnor U9358 (N_9358,N_8064,N_7840);
xnor U9359 (N_9359,N_7572,N_7273);
or U9360 (N_9360,N_7380,N_7360);
and U9361 (N_9361,N_7386,N_7622);
nor U9362 (N_9362,N_7995,N_7412);
nand U9363 (N_9363,N_7923,N_7214);
or U9364 (N_9364,N_7500,N_7936);
nor U9365 (N_9365,N_8054,N_7471);
nand U9366 (N_9366,N_7240,N_7575);
or U9367 (N_9367,N_7217,N_7990);
nor U9368 (N_9368,N_7282,N_7787);
nor U9369 (N_9369,N_7291,N_8315);
xor U9370 (N_9370,N_7912,N_7413);
or U9371 (N_9371,N_8221,N_8373);
or U9372 (N_9372,N_7874,N_7419);
xnor U9373 (N_9373,N_8020,N_8380);
or U9374 (N_9374,N_8210,N_7267);
or U9375 (N_9375,N_7514,N_8156);
or U9376 (N_9376,N_7766,N_7969);
nand U9377 (N_9377,N_7922,N_7261);
xnor U9378 (N_9378,N_7786,N_8157);
and U9379 (N_9379,N_7776,N_8204);
and U9380 (N_9380,N_8170,N_7502);
xnor U9381 (N_9381,N_7386,N_7304);
and U9382 (N_9382,N_7462,N_7916);
nand U9383 (N_9383,N_7766,N_8001);
or U9384 (N_9384,N_8022,N_7720);
and U9385 (N_9385,N_7823,N_7873);
nand U9386 (N_9386,N_7520,N_8298);
or U9387 (N_9387,N_7728,N_8331);
nor U9388 (N_9388,N_7963,N_8158);
or U9389 (N_9389,N_7365,N_7441);
and U9390 (N_9390,N_7336,N_7738);
or U9391 (N_9391,N_7910,N_7561);
nor U9392 (N_9392,N_7360,N_7383);
xor U9393 (N_9393,N_8342,N_7329);
and U9394 (N_9394,N_7545,N_7406);
nand U9395 (N_9395,N_8294,N_8057);
xnor U9396 (N_9396,N_7522,N_7779);
nor U9397 (N_9397,N_8384,N_7633);
nand U9398 (N_9398,N_8004,N_7702);
nand U9399 (N_9399,N_8023,N_7576);
or U9400 (N_9400,N_7616,N_7613);
nor U9401 (N_9401,N_8340,N_7286);
and U9402 (N_9402,N_7822,N_8287);
or U9403 (N_9403,N_7861,N_8071);
nor U9404 (N_9404,N_7442,N_7635);
and U9405 (N_9405,N_7367,N_7960);
or U9406 (N_9406,N_7634,N_7521);
nand U9407 (N_9407,N_8039,N_8383);
or U9408 (N_9408,N_8102,N_8351);
nor U9409 (N_9409,N_8119,N_7629);
xor U9410 (N_9410,N_7271,N_8172);
nor U9411 (N_9411,N_8038,N_7687);
nor U9412 (N_9412,N_7938,N_8167);
xnor U9413 (N_9413,N_7993,N_7369);
nor U9414 (N_9414,N_7613,N_7332);
nand U9415 (N_9415,N_7302,N_7703);
and U9416 (N_9416,N_8224,N_8285);
or U9417 (N_9417,N_8238,N_7346);
and U9418 (N_9418,N_8164,N_8396);
xor U9419 (N_9419,N_8209,N_7427);
or U9420 (N_9420,N_7225,N_7222);
or U9421 (N_9421,N_7260,N_7944);
and U9422 (N_9422,N_7733,N_7915);
xnor U9423 (N_9423,N_7855,N_7479);
or U9424 (N_9424,N_7272,N_8105);
nand U9425 (N_9425,N_8098,N_7587);
xnor U9426 (N_9426,N_7616,N_7708);
or U9427 (N_9427,N_8312,N_7918);
nor U9428 (N_9428,N_7491,N_7284);
nor U9429 (N_9429,N_7627,N_7471);
xnor U9430 (N_9430,N_7249,N_8025);
nand U9431 (N_9431,N_8167,N_7697);
or U9432 (N_9432,N_8094,N_7589);
xor U9433 (N_9433,N_7396,N_7643);
nor U9434 (N_9434,N_8073,N_8040);
and U9435 (N_9435,N_7802,N_7996);
or U9436 (N_9436,N_7548,N_8216);
and U9437 (N_9437,N_7641,N_7480);
or U9438 (N_9438,N_7692,N_8215);
xnor U9439 (N_9439,N_7473,N_7632);
nand U9440 (N_9440,N_7824,N_7736);
nand U9441 (N_9441,N_8393,N_8064);
or U9442 (N_9442,N_7367,N_7427);
or U9443 (N_9443,N_7509,N_7476);
or U9444 (N_9444,N_8029,N_7876);
nor U9445 (N_9445,N_7789,N_7209);
nor U9446 (N_9446,N_7487,N_8358);
xor U9447 (N_9447,N_7399,N_7490);
nand U9448 (N_9448,N_7686,N_7474);
nor U9449 (N_9449,N_7372,N_8138);
nor U9450 (N_9450,N_7739,N_7200);
xor U9451 (N_9451,N_7681,N_8011);
or U9452 (N_9452,N_8095,N_8021);
xor U9453 (N_9453,N_7672,N_7931);
nor U9454 (N_9454,N_8254,N_8098);
or U9455 (N_9455,N_7709,N_7656);
xor U9456 (N_9456,N_8276,N_8072);
nor U9457 (N_9457,N_7941,N_7427);
nand U9458 (N_9458,N_8283,N_8375);
nand U9459 (N_9459,N_7906,N_8107);
xnor U9460 (N_9460,N_7548,N_8069);
nand U9461 (N_9461,N_7544,N_8285);
nor U9462 (N_9462,N_7593,N_7356);
and U9463 (N_9463,N_8177,N_7590);
nor U9464 (N_9464,N_7645,N_7956);
xnor U9465 (N_9465,N_7531,N_7994);
and U9466 (N_9466,N_7860,N_8177);
or U9467 (N_9467,N_8177,N_7517);
nor U9468 (N_9468,N_7607,N_8301);
nor U9469 (N_9469,N_8236,N_7627);
and U9470 (N_9470,N_7482,N_7728);
or U9471 (N_9471,N_7375,N_8218);
nor U9472 (N_9472,N_7716,N_8235);
and U9473 (N_9473,N_7416,N_8233);
nor U9474 (N_9474,N_7970,N_7424);
or U9475 (N_9475,N_7330,N_8263);
nand U9476 (N_9476,N_8037,N_7388);
nand U9477 (N_9477,N_7575,N_7550);
and U9478 (N_9478,N_7288,N_7543);
xor U9479 (N_9479,N_7718,N_8234);
or U9480 (N_9480,N_8124,N_7498);
xor U9481 (N_9481,N_8334,N_7461);
and U9482 (N_9482,N_8153,N_7501);
nor U9483 (N_9483,N_7490,N_7564);
xnor U9484 (N_9484,N_7646,N_7711);
and U9485 (N_9485,N_7829,N_8116);
nor U9486 (N_9486,N_7301,N_8232);
and U9487 (N_9487,N_8368,N_7608);
and U9488 (N_9488,N_7995,N_7836);
nand U9489 (N_9489,N_8059,N_7912);
nor U9490 (N_9490,N_7487,N_8055);
or U9491 (N_9491,N_7388,N_7737);
or U9492 (N_9492,N_8081,N_8399);
or U9493 (N_9493,N_7579,N_8139);
nor U9494 (N_9494,N_7655,N_8164);
nand U9495 (N_9495,N_7390,N_7545);
and U9496 (N_9496,N_7817,N_7376);
and U9497 (N_9497,N_7799,N_7207);
xor U9498 (N_9498,N_8045,N_7298);
and U9499 (N_9499,N_8329,N_8054);
nand U9500 (N_9500,N_7879,N_8072);
nor U9501 (N_9501,N_7956,N_8273);
xor U9502 (N_9502,N_8173,N_7504);
xnor U9503 (N_9503,N_8171,N_8133);
or U9504 (N_9504,N_7206,N_8364);
nand U9505 (N_9505,N_8358,N_7866);
and U9506 (N_9506,N_7439,N_7517);
xnor U9507 (N_9507,N_7996,N_7890);
nand U9508 (N_9508,N_8299,N_7776);
and U9509 (N_9509,N_7670,N_8320);
nor U9510 (N_9510,N_7236,N_7980);
nand U9511 (N_9511,N_7949,N_7646);
or U9512 (N_9512,N_7786,N_8128);
and U9513 (N_9513,N_8384,N_7578);
or U9514 (N_9514,N_7394,N_7665);
or U9515 (N_9515,N_8011,N_7231);
nor U9516 (N_9516,N_7989,N_8103);
and U9517 (N_9517,N_8129,N_7693);
xnor U9518 (N_9518,N_7699,N_7582);
nand U9519 (N_9519,N_8353,N_7324);
xnor U9520 (N_9520,N_8295,N_7818);
nand U9521 (N_9521,N_8219,N_7969);
nand U9522 (N_9522,N_7559,N_8018);
nand U9523 (N_9523,N_7981,N_8087);
and U9524 (N_9524,N_7910,N_7829);
nand U9525 (N_9525,N_8046,N_8061);
nand U9526 (N_9526,N_7203,N_7728);
xnor U9527 (N_9527,N_7763,N_8315);
or U9528 (N_9528,N_7760,N_7281);
nor U9529 (N_9529,N_7930,N_8068);
nand U9530 (N_9530,N_7577,N_7521);
and U9531 (N_9531,N_8258,N_7413);
and U9532 (N_9532,N_8282,N_8272);
nand U9533 (N_9533,N_7360,N_8042);
nor U9534 (N_9534,N_8314,N_7508);
xnor U9535 (N_9535,N_8098,N_7991);
or U9536 (N_9536,N_7274,N_7717);
or U9537 (N_9537,N_7768,N_7204);
and U9538 (N_9538,N_8092,N_7335);
and U9539 (N_9539,N_7569,N_8250);
and U9540 (N_9540,N_7488,N_7948);
nand U9541 (N_9541,N_7348,N_7657);
nor U9542 (N_9542,N_7823,N_8375);
and U9543 (N_9543,N_8174,N_7446);
or U9544 (N_9544,N_7666,N_8211);
or U9545 (N_9545,N_7479,N_8127);
nand U9546 (N_9546,N_7529,N_7751);
nor U9547 (N_9547,N_7684,N_8280);
nor U9548 (N_9548,N_7565,N_7877);
xnor U9549 (N_9549,N_8012,N_7500);
and U9550 (N_9550,N_8352,N_7597);
xnor U9551 (N_9551,N_8361,N_7316);
and U9552 (N_9552,N_7691,N_8032);
nor U9553 (N_9553,N_8308,N_7735);
and U9554 (N_9554,N_7893,N_8199);
xor U9555 (N_9555,N_7431,N_7439);
and U9556 (N_9556,N_8127,N_8381);
xnor U9557 (N_9557,N_7276,N_7550);
and U9558 (N_9558,N_7447,N_7877);
nand U9559 (N_9559,N_7246,N_7942);
xnor U9560 (N_9560,N_7338,N_7790);
nor U9561 (N_9561,N_7845,N_7711);
and U9562 (N_9562,N_7658,N_7354);
nor U9563 (N_9563,N_8238,N_8272);
nand U9564 (N_9564,N_7424,N_8083);
xnor U9565 (N_9565,N_7222,N_8298);
xor U9566 (N_9566,N_7814,N_7464);
and U9567 (N_9567,N_7405,N_7456);
xor U9568 (N_9568,N_8072,N_7312);
nor U9569 (N_9569,N_8388,N_8004);
nor U9570 (N_9570,N_7384,N_7982);
and U9571 (N_9571,N_7604,N_7781);
nor U9572 (N_9572,N_8312,N_7225);
nor U9573 (N_9573,N_8184,N_7502);
xnor U9574 (N_9574,N_7971,N_7286);
xnor U9575 (N_9575,N_7214,N_7229);
and U9576 (N_9576,N_7239,N_7792);
or U9577 (N_9577,N_7235,N_8108);
nor U9578 (N_9578,N_7760,N_7378);
xor U9579 (N_9579,N_7708,N_7648);
and U9580 (N_9580,N_7675,N_7314);
or U9581 (N_9581,N_8073,N_7664);
nand U9582 (N_9582,N_7665,N_7509);
or U9583 (N_9583,N_7648,N_7304);
and U9584 (N_9584,N_7998,N_7433);
or U9585 (N_9585,N_7373,N_7322);
and U9586 (N_9586,N_7563,N_8315);
and U9587 (N_9587,N_7219,N_7599);
nor U9588 (N_9588,N_7252,N_7420);
nand U9589 (N_9589,N_8094,N_7704);
nor U9590 (N_9590,N_7369,N_8284);
or U9591 (N_9591,N_7986,N_7467);
and U9592 (N_9592,N_7605,N_7215);
or U9593 (N_9593,N_7795,N_8157);
xor U9594 (N_9594,N_8395,N_8320);
xnor U9595 (N_9595,N_8012,N_7994);
and U9596 (N_9596,N_7521,N_7304);
and U9597 (N_9597,N_7353,N_7233);
or U9598 (N_9598,N_7596,N_8204);
and U9599 (N_9599,N_8317,N_7806);
nor U9600 (N_9600,N_8714,N_8858);
and U9601 (N_9601,N_9322,N_8942);
and U9602 (N_9602,N_8849,N_9187);
or U9603 (N_9603,N_9123,N_9443);
xor U9604 (N_9604,N_9454,N_8591);
or U9605 (N_9605,N_9037,N_8632);
nor U9606 (N_9606,N_9512,N_9175);
and U9607 (N_9607,N_9113,N_8847);
nor U9608 (N_9608,N_8906,N_8732);
and U9609 (N_9609,N_9242,N_8494);
or U9610 (N_9610,N_9588,N_8533);
or U9611 (N_9611,N_9425,N_8894);
nor U9612 (N_9612,N_8963,N_8902);
and U9613 (N_9613,N_8544,N_8603);
nor U9614 (N_9614,N_9134,N_8556);
and U9615 (N_9615,N_9292,N_8552);
xnor U9616 (N_9616,N_9361,N_8650);
nand U9617 (N_9617,N_9332,N_9389);
or U9618 (N_9618,N_8834,N_8829);
or U9619 (N_9619,N_8497,N_9480);
and U9620 (N_9620,N_9135,N_8742);
nor U9621 (N_9621,N_9024,N_8521);
and U9622 (N_9622,N_8947,N_8968);
nand U9623 (N_9623,N_9407,N_8884);
nand U9624 (N_9624,N_9397,N_8867);
nor U9625 (N_9625,N_8637,N_8755);
xor U9626 (N_9626,N_8583,N_9566);
nor U9627 (N_9627,N_8487,N_8741);
xor U9628 (N_9628,N_9234,N_8433);
nor U9629 (N_9629,N_9380,N_9519);
nand U9630 (N_9630,N_8510,N_9367);
xnor U9631 (N_9631,N_8631,N_9260);
nor U9632 (N_9632,N_8720,N_8477);
or U9633 (N_9633,N_9273,N_9093);
nor U9634 (N_9634,N_9471,N_9592);
and U9635 (N_9635,N_9483,N_8406);
or U9636 (N_9636,N_9277,N_8962);
xnor U9637 (N_9637,N_8641,N_9424);
xor U9638 (N_9638,N_9334,N_9415);
nor U9639 (N_9639,N_8657,N_9097);
or U9640 (N_9640,N_9593,N_9092);
or U9641 (N_9641,N_9133,N_9439);
and U9642 (N_9642,N_8473,N_8743);
or U9643 (N_9643,N_9453,N_8970);
or U9644 (N_9644,N_9170,N_9079);
and U9645 (N_9645,N_8917,N_9305);
nor U9646 (N_9646,N_9524,N_9475);
or U9647 (N_9647,N_8600,N_8647);
nand U9648 (N_9648,N_8798,N_9262);
or U9649 (N_9649,N_8581,N_9271);
and U9650 (N_9650,N_8469,N_8653);
nor U9651 (N_9651,N_9243,N_8423);
nand U9652 (N_9652,N_8978,N_8934);
xor U9653 (N_9653,N_9052,N_8957);
and U9654 (N_9654,N_8886,N_9550);
xor U9655 (N_9655,N_8440,N_9213);
nand U9656 (N_9656,N_9573,N_8809);
xnor U9657 (N_9657,N_8693,N_8622);
nand U9658 (N_9658,N_9042,N_9217);
nand U9659 (N_9659,N_9046,N_8515);
nand U9660 (N_9660,N_9560,N_8548);
nand U9661 (N_9661,N_9100,N_9153);
nand U9662 (N_9662,N_9562,N_8746);
nand U9663 (N_9663,N_8682,N_8706);
or U9664 (N_9664,N_8425,N_9120);
xor U9665 (N_9665,N_8453,N_8921);
nand U9666 (N_9666,N_8883,N_8441);
nor U9667 (N_9667,N_9462,N_9055);
nand U9668 (N_9668,N_9574,N_8669);
xnor U9669 (N_9669,N_9326,N_9286);
xnor U9670 (N_9670,N_8655,N_9402);
nor U9671 (N_9671,N_8496,N_8671);
nand U9672 (N_9672,N_9340,N_9142);
nand U9673 (N_9673,N_9222,N_8754);
xor U9674 (N_9674,N_8436,N_8920);
nor U9675 (N_9675,N_9220,N_8846);
xnor U9676 (N_9676,N_9571,N_8447);
or U9677 (N_9677,N_8862,N_8526);
nand U9678 (N_9678,N_9227,N_8553);
xnor U9679 (N_9679,N_9418,N_9096);
and U9680 (N_9680,N_9061,N_9364);
or U9681 (N_9681,N_9004,N_8984);
nand U9682 (N_9682,N_9247,N_8981);
or U9683 (N_9683,N_8745,N_9535);
xor U9684 (N_9684,N_8474,N_9224);
nand U9685 (N_9685,N_8750,N_8504);
nand U9686 (N_9686,N_9285,N_8778);
and U9687 (N_9687,N_9147,N_8617);
and U9688 (N_9688,N_8860,N_8513);
xor U9689 (N_9689,N_8822,N_8676);
nand U9690 (N_9690,N_8488,N_9281);
nor U9691 (N_9691,N_8993,N_9484);
or U9692 (N_9692,N_8446,N_9163);
or U9693 (N_9693,N_8932,N_9396);
xnor U9694 (N_9694,N_8634,N_8456);
nand U9695 (N_9695,N_8989,N_8432);
nand U9696 (N_9696,N_9409,N_9428);
and U9697 (N_9697,N_8564,N_9327);
nand U9698 (N_9698,N_9143,N_9410);
nor U9699 (N_9699,N_9552,N_8520);
nand U9700 (N_9700,N_9017,N_9338);
nand U9701 (N_9701,N_8815,N_8565);
nor U9702 (N_9702,N_8997,N_8592);
nor U9703 (N_9703,N_9118,N_9040);
nor U9704 (N_9704,N_8408,N_9073);
nor U9705 (N_9705,N_9461,N_8568);
nor U9706 (N_9706,N_8787,N_8551);
xor U9707 (N_9707,N_8492,N_8975);
or U9708 (N_9708,N_8639,N_9272);
and U9709 (N_9709,N_9476,N_8752);
nand U9710 (N_9710,N_9282,N_9466);
xnor U9711 (N_9711,N_8943,N_8602);
and U9712 (N_9712,N_8889,N_9577);
nand U9713 (N_9713,N_9493,N_8776);
nor U9714 (N_9714,N_8769,N_8522);
nand U9715 (N_9715,N_9442,N_8500);
and U9716 (N_9716,N_9053,N_8580);
xnor U9717 (N_9717,N_9348,N_8796);
nand U9718 (N_9718,N_8944,N_9164);
nor U9719 (N_9719,N_9275,N_8576);
nor U9720 (N_9720,N_9283,N_9555);
or U9721 (N_9721,N_8797,N_9206);
xnor U9722 (N_9722,N_9506,N_8737);
or U9723 (N_9723,N_8724,N_9357);
xnor U9724 (N_9724,N_9330,N_9300);
nor U9725 (N_9725,N_9490,N_9473);
or U9726 (N_9726,N_9148,N_8900);
nor U9727 (N_9727,N_8470,N_9478);
and U9728 (N_9728,N_8927,N_8559);
nand U9729 (N_9729,N_8897,N_8570);
nor U9730 (N_9730,N_9132,N_9088);
nor U9731 (N_9731,N_9551,N_8407);
xor U9732 (N_9732,N_9501,N_9094);
and U9733 (N_9733,N_9567,N_8539);
or U9734 (N_9734,N_9504,N_8982);
nand U9735 (N_9735,N_9515,N_8810);
or U9736 (N_9736,N_9559,N_8698);
nand U9737 (N_9737,N_9267,N_9549);
nand U9738 (N_9738,N_8690,N_9181);
or U9739 (N_9739,N_9057,N_9505);
xnor U9740 (N_9740,N_9235,N_8793);
and U9741 (N_9741,N_9032,N_8730);
xor U9742 (N_9742,N_9440,N_9117);
and U9743 (N_9743,N_9597,N_9544);
nand U9744 (N_9744,N_9302,N_8431);
nand U9745 (N_9745,N_9511,N_9238);
xor U9746 (N_9746,N_8751,N_9201);
and U9747 (N_9747,N_9180,N_9007);
or U9748 (N_9748,N_8478,N_8926);
or U9749 (N_9749,N_8571,N_8998);
or U9750 (N_9750,N_8842,N_9495);
nor U9751 (N_9751,N_9158,N_8455);
and U9752 (N_9752,N_9006,N_9188);
xnor U9753 (N_9753,N_8645,N_9316);
and U9754 (N_9754,N_9295,N_9075);
and U9755 (N_9755,N_9414,N_9104);
nor U9756 (N_9756,N_8885,N_9304);
and U9757 (N_9757,N_9528,N_8700);
or U9758 (N_9758,N_9569,N_8424);
nor U9759 (N_9759,N_8573,N_8485);
or U9760 (N_9760,N_8722,N_9047);
or U9761 (N_9761,N_8479,N_9189);
nor U9762 (N_9762,N_8615,N_8610);
or U9763 (N_9763,N_9012,N_8877);
nor U9764 (N_9764,N_8620,N_8516);
nor U9765 (N_9765,N_8801,N_8624);
xnor U9766 (N_9766,N_8905,N_8593);
xor U9767 (N_9767,N_9139,N_8996);
nand U9768 (N_9768,N_8726,N_8955);
and U9769 (N_9769,N_9399,N_9353);
and U9770 (N_9770,N_9541,N_9510);
nand U9771 (N_9771,N_9491,N_8910);
nand U9772 (N_9772,N_9202,N_8983);
nor U9773 (N_9773,N_9537,N_8694);
xor U9774 (N_9774,N_9306,N_8691);
or U9775 (N_9775,N_8483,N_8715);
nor U9776 (N_9776,N_8794,N_9179);
and U9777 (N_9777,N_9150,N_8531);
and U9778 (N_9778,N_8563,N_9193);
xor U9779 (N_9779,N_9126,N_8511);
nor U9780 (N_9780,N_8529,N_8458);
xor U9781 (N_9781,N_8940,N_9074);
and U9782 (N_9782,N_8519,N_9563);
or U9783 (N_9783,N_9464,N_8584);
or U9784 (N_9784,N_9077,N_9078);
nor U9785 (N_9785,N_8748,N_9082);
nand U9786 (N_9786,N_8557,N_9323);
xor U9787 (N_9787,N_9536,N_8912);
nor U9788 (N_9788,N_9026,N_8590);
xor U9789 (N_9789,N_9543,N_8566);
or U9790 (N_9790,N_9342,N_8954);
and U9791 (N_9791,N_8892,N_8628);
xnor U9792 (N_9792,N_9433,N_9420);
or U9793 (N_9793,N_8911,N_8501);
or U9794 (N_9794,N_8950,N_9575);
and U9795 (N_9795,N_8859,N_8735);
and U9796 (N_9796,N_9377,N_9056);
xor U9797 (N_9797,N_8712,N_9030);
and U9798 (N_9798,N_9351,N_8833);
nand U9799 (N_9799,N_8802,N_9091);
and U9800 (N_9800,N_9090,N_9246);
and U9801 (N_9801,N_8792,N_9467);
nor U9802 (N_9802,N_9125,N_8874);
nor U9803 (N_9803,N_9130,N_9208);
or U9804 (N_9804,N_8995,N_9025);
xor U9805 (N_9805,N_8870,N_9470);
and U9806 (N_9806,N_9263,N_9161);
and U9807 (N_9807,N_8661,N_9225);
nor U9808 (N_9808,N_9131,N_9412);
or U9809 (N_9809,N_9314,N_9468);
xor U9810 (N_9810,N_8903,N_8916);
xnor U9811 (N_9811,N_8701,N_8744);
nand U9812 (N_9812,N_8648,N_8967);
nor U9813 (N_9813,N_9087,N_9324);
nand U9814 (N_9814,N_9523,N_8974);
and U9815 (N_9815,N_8879,N_9400);
xor U9816 (N_9816,N_9098,N_9028);
and U9817 (N_9817,N_8945,N_8696);
nor U9818 (N_9818,N_9352,N_8465);
xor U9819 (N_9819,N_9223,N_9230);
or U9820 (N_9820,N_8466,N_8820);
or U9821 (N_9821,N_8731,N_9081);
and U9822 (N_9822,N_9394,N_8437);
xnor U9823 (N_9823,N_8536,N_8838);
nor U9824 (N_9824,N_9110,N_8505);
or U9825 (N_9825,N_8625,N_8606);
xor U9826 (N_9826,N_8430,N_9458);
xor U9827 (N_9827,N_8717,N_9381);
and U9828 (N_9828,N_8541,N_9497);
nor U9829 (N_9829,N_8909,N_9533);
and U9830 (N_9830,N_8965,N_8880);
and U9831 (N_9831,N_8758,N_9371);
and U9832 (N_9832,N_9200,N_9146);
or U9833 (N_9833,N_9518,N_9488);
or U9834 (N_9834,N_8946,N_9171);
and U9835 (N_9835,N_9190,N_9438);
xnor U9836 (N_9836,N_9121,N_9391);
xnor U9837 (N_9837,N_8992,N_8991);
or U9838 (N_9838,N_8855,N_8644);
xor U9839 (N_9839,N_8629,N_8422);
xnor U9840 (N_9840,N_9109,N_9197);
and U9841 (N_9841,N_8512,N_8836);
or U9842 (N_9842,N_9259,N_9313);
nand U9843 (N_9843,N_8532,N_9445);
or U9844 (N_9844,N_8609,N_8768);
nand U9845 (N_9845,N_8662,N_8845);
nand U9846 (N_9846,N_9023,N_8938);
or U9847 (N_9847,N_9054,N_8843);
or U9848 (N_9848,N_9565,N_9115);
nor U9849 (N_9849,N_9196,N_8688);
or U9850 (N_9850,N_9296,N_9430);
or U9851 (N_9851,N_9444,N_9261);
nor U9852 (N_9852,N_9219,N_9346);
nor U9853 (N_9853,N_9269,N_9049);
and U9854 (N_9854,N_8537,N_8508);
nor U9855 (N_9855,N_9395,N_9525);
xor U9856 (N_9856,N_8988,N_8756);
nand U9857 (N_9857,N_9048,N_9554);
and U9858 (N_9858,N_8964,N_8543);
nand U9859 (N_9859,N_9513,N_8663);
nand U9860 (N_9860,N_9383,N_9341);
nand U9861 (N_9861,N_9401,N_9336);
or U9862 (N_9862,N_8596,N_8630);
or U9863 (N_9863,N_8826,N_8813);
nand U9864 (N_9864,N_9065,N_8555);
nor U9865 (N_9865,N_9257,N_8907);
xor U9866 (N_9866,N_8540,N_9318);
or U9867 (N_9867,N_8805,N_9003);
and U9868 (N_9868,N_8835,N_8499);
and U9869 (N_9869,N_8651,N_8857);
or U9870 (N_9870,N_9101,N_8994);
or U9871 (N_9871,N_8549,N_9404);
xor U9872 (N_9872,N_8888,N_8454);
nand U9873 (N_9873,N_8811,N_9556);
nor U9874 (N_9874,N_8445,N_9168);
and U9875 (N_9875,N_9485,N_8850);
or U9876 (N_9876,N_8729,N_8438);
and U9877 (N_9877,N_9539,N_9469);
xor U9878 (N_9878,N_8704,N_8604);
and U9879 (N_9879,N_9154,N_8814);
xor U9880 (N_9880,N_8901,N_9591);
xor U9881 (N_9881,N_8525,N_9050);
and U9882 (N_9882,N_8684,N_9116);
or U9883 (N_9883,N_9122,N_8733);
nand U9884 (N_9884,N_8495,N_9522);
nor U9885 (N_9885,N_8839,N_8679);
nor U9886 (N_9886,N_8413,N_9320);
or U9887 (N_9887,N_8868,N_8918);
and U9888 (N_9888,N_9293,N_8670);
and U9889 (N_9889,N_9218,N_9452);
xor U9890 (N_9890,N_9372,N_8558);
and U9891 (N_9891,N_9000,N_9029);
xnor U9892 (N_9892,N_8928,N_8468);
nand U9893 (N_9893,N_8775,N_8844);
and U9894 (N_9894,N_9205,N_8471);
and U9895 (N_9895,N_8827,N_8803);
and U9896 (N_9896,N_9578,N_8482);
nand U9897 (N_9897,N_8535,N_8727);
nand U9898 (N_9898,N_9034,N_9455);
xnor U9899 (N_9899,N_8681,N_8493);
and U9900 (N_9900,N_9041,N_8831);
or U9901 (N_9901,N_9195,N_9038);
or U9902 (N_9902,N_8923,N_8443);
and U9903 (N_9903,N_9514,N_9033);
nand U9904 (N_9904,N_8587,N_8575);
or U9905 (N_9905,N_8875,N_9343);
nor U9906 (N_9906,N_9066,N_9199);
nand U9907 (N_9907,N_9465,N_9449);
nor U9908 (N_9908,N_9328,N_8426);
nor U9909 (N_9909,N_8871,N_9508);
xor U9910 (N_9910,N_9172,N_8891);
and U9911 (N_9911,N_9062,N_8760);
and U9912 (N_9912,N_8817,N_8626);
nand U9913 (N_9913,N_8452,N_9043);
xor U9914 (N_9914,N_8586,N_8611);
nor U9915 (N_9915,N_8716,N_8861);
or U9916 (N_9916,N_8766,N_8614);
nor U9917 (N_9917,N_9553,N_8990);
xnor U9918 (N_9918,N_8898,N_8841);
nand U9919 (N_9919,N_9141,N_9589);
or U9920 (N_9920,N_9398,N_8419);
and U9921 (N_9921,N_9287,N_9446);
and U9922 (N_9922,N_9011,N_9228);
and U9923 (N_9923,N_9317,N_9583);
nor U9924 (N_9924,N_8574,N_8976);
and U9925 (N_9925,N_9308,N_8736);
and U9926 (N_9926,N_8585,N_9312);
nand U9927 (N_9927,N_9157,N_9059);
or U9928 (N_9928,N_8919,N_9595);
and U9929 (N_9929,N_8761,N_8782);
nand U9930 (N_9930,N_8780,N_9347);
and U9931 (N_9931,N_8958,N_8415);
or U9932 (N_9932,N_8764,N_8924);
or U9933 (N_9933,N_9507,N_8759);
and U9934 (N_9934,N_9297,N_8400);
xnor U9935 (N_9935,N_8449,N_9587);
and U9936 (N_9936,N_8507,N_9221);
nand U9937 (N_9937,N_9472,N_9534);
or U9938 (N_9938,N_8589,N_9018);
and U9939 (N_9939,N_9459,N_8800);
nor U9940 (N_9940,N_8824,N_9105);
nor U9941 (N_9941,N_9335,N_9264);
nor U9942 (N_9942,N_8808,N_9112);
nand U9943 (N_9943,N_8770,N_8719);
xor U9944 (N_9944,N_8658,N_8969);
and U9945 (N_9945,N_8692,N_8828);
nor U9946 (N_9946,N_9124,N_9358);
nor U9947 (N_9947,N_9252,N_8598);
xor U9948 (N_9948,N_9384,N_9564);
and U9949 (N_9949,N_9329,N_9226);
xor U9950 (N_9950,N_8542,N_8638);
nor U9951 (N_9951,N_8786,N_8687);
and U9952 (N_9952,N_9063,N_9390);
nand U9953 (N_9953,N_9502,N_9558);
nor U9954 (N_9954,N_8623,N_8523);
or U9955 (N_9955,N_9102,N_9474);
and U9956 (N_9956,N_8594,N_9114);
and U9957 (N_9957,N_9127,N_8935);
and U9958 (N_9958,N_9258,N_8956);
nor U9959 (N_9959,N_8773,N_9517);
or U9960 (N_9960,N_8837,N_9557);
and U9961 (N_9961,N_9129,N_8667);
nand U9962 (N_9962,N_8621,N_9450);
nor U9963 (N_9963,N_9014,N_8685);
nor U9964 (N_9964,N_9568,N_8767);
nor U9965 (N_9965,N_8818,N_9481);
and U9966 (N_9966,N_9451,N_9477);
or U9967 (N_9967,N_8734,N_9002);
nand U9968 (N_9968,N_8922,N_9321);
nand U9969 (N_9969,N_8444,N_9254);
xnor U9970 (N_9970,N_9356,N_8675);
or U9971 (N_9971,N_9067,N_9192);
or U9972 (N_9972,N_9426,N_9266);
nand U9973 (N_9973,N_8547,N_9162);
nand U9974 (N_9974,N_8753,N_9447);
and U9975 (N_9975,N_8749,N_9060);
nand U9976 (N_9976,N_8832,N_9151);
or U9977 (N_9977,N_8977,N_9185);
or U9978 (N_9978,N_9457,N_8779);
and U9979 (N_9979,N_9339,N_9265);
or U9980 (N_9980,N_8649,N_9086);
xor U9981 (N_9981,N_9136,N_8409);
or U9982 (N_9982,N_9255,N_8896);
xor U9983 (N_9983,N_8578,N_9128);
nand U9984 (N_9984,N_8428,N_9406);
xnor U9985 (N_9985,N_9530,N_9108);
nor U9986 (N_9986,N_8403,N_9289);
and U9987 (N_9987,N_8567,N_8789);
nand U9988 (N_9988,N_9435,N_8941);
nor U9989 (N_9989,N_9184,N_8481);
or U9990 (N_9990,N_8689,N_8895);
xnor U9991 (N_9991,N_9076,N_9579);
xnor U9992 (N_9992,N_8527,N_8640);
xnor U9993 (N_9993,N_9432,N_8472);
xnor U9994 (N_9994,N_8777,N_9527);
and U9995 (N_9995,N_9106,N_9279);
nand U9996 (N_9996,N_9210,N_9337);
nand U9997 (N_9997,N_9229,N_9362);
or U9998 (N_9998,N_9355,N_8502);
xnor U9999 (N_9999,N_8709,N_9576);
nand U10000 (N_10000,N_8665,N_9350);
nand U10001 (N_10001,N_9204,N_9194);
nor U10002 (N_10002,N_8616,N_8664);
nand U10003 (N_10003,N_8418,N_9280);
and U10004 (N_10004,N_8613,N_9021);
nor U10005 (N_10005,N_9463,N_8790);
or U10006 (N_10006,N_9027,N_8959);
and U10007 (N_10007,N_8697,N_9392);
or U10008 (N_10008,N_9174,N_8864);
or U10009 (N_10009,N_9370,N_8448);
and U10010 (N_10010,N_8979,N_8763);
or U10011 (N_10011,N_9520,N_8728);
xnor U10012 (N_10012,N_9211,N_8467);
and U10013 (N_10013,N_8673,N_9183);
nand U10014 (N_10014,N_9509,N_9248);
nor U10015 (N_10015,N_8869,N_8972);
nand U10016 (N_10016,N_9429,N_9365);
xor U10017 (N_10017,N_8656,N_9408);
xor U10018 (N_10018,N_8678,N_9270);
xor U10019 (N_10019,N_8881,N_9019);
xor U10020 (N_10020,N_9572,N_8960);
xnor U10021 (N_10021,N_8546,N_9178);
xnor U10022 (N_10022,N_9570,N_8873);
nor U10023 (N_10023,N_8740,N_9311);
nor U10024 (N_10024,N_8784,N_9005);
and U10025 (N_10025,N_9251,N_8659);
nand U10026 (N_10026,N_8416,N_9531);
nor U10027 (N_10027,N_9241,N_9385);
nand U10028 (N_10028,N_9363,N_8601);
nand U10029 (N_10029,N_9421,N_8562);
xnor U10030 (N_10030,N_9582,N_9431);
nor U10031 (N_10031,N_9448,N_8434);
and U10032 (N_10032,N_9159,N_9169);
xor U10033 (N_10033,N_9237,N_9590);
nand U10034 (N_10034,N_9008,N_9010);
nand U10035 (N_10035,N_8904,N_8514);
and U10036 (N_10036,N_8577,N_8410);
xnor U10037 (N_10037,N_8484,N_9207);
and U10038 (N_10038,N_9035,N_9182);
nor U10039 (N_10039,N_8703,N_9290);
nor U10040 (N_10040,N_8660,N_9232);
xnor U10041 (N_10041,N_8804,N_8427);
or U10042 (N_10042,N_8854,N_9494);
or U10043 (N_10043,N_9379,N_9521);
nor U10044 (N_10044,N_9596,N_9249);
and U10045 (N_10045,N_9103,N_8951);
nand U10046 (N_10046,N_8929,N_9538);
nand U10047 (N_10047,N_9268,N_9186);
and U10048 (N_10048,N_8771,N_9016);
xor U10049 (N_10049,N_8939,N_8652);
nor U10050 (N_10050,N_8866,N_9173);
nand U10051 (N_10051,N_8666,N_9291);
nor U10052 (N_10052,N_8710,N_9144);
nand U10053 (N_10053,N_8816,N_9331);
nor U10054 (N_10054,N_8893,N_9039);
or U10055 (N_10055,N_9152,N_9548);
nor U10056 (N_10056,N_9214,N_9434);
nor U10057 (N_10057,N_9354,N_9333);
and U10058 (N_10058,N_8608,N_9250);
or U10059 (N_10059,N_8480,N_9496);
nand U10060 (N_10060,N_9546,N_9532);
and U10061 (N_10061,N_9276,N_9001);
xnor U10062 (N_10062,N_8791,N_8435);
xnor U10063 (N_10063,N_8530,N_8599);
or U10064 (N_10064,N_9099,N_8713);
or U10065 (N_10065,N_9083,N_8627);
or U10066 (N_10066,N_9107,N_9393);
and U10067 (N_10067,N_8607,N_8524);
or U10068 (N_10068,N_9020,N_9441);
and U10069 (N_10069,N_9301,N_9209);
nand U10070 (N_10070,N_9498,N_9138);
or U10071 (N_10071,N_8785,N_9594);
nor U10072 (N_10072,N_9298,N_9310);
and U10073 (N_10073,N_9245,N_8421);
xnor U10074 (N_10074,N_8489,N_9487);
and U10075 (N_10075,N_8491,N_9031);
and U10076 (N_10076,N_8461,N_9111);
nor U10077 (N_10077,N_9547,N_9584);
nand U10078 (N_10078,N_9413,N_9244);
or U10079 (N_10079,N_8757,N_9374);
or U10080 (N_10080,N_8442,N_8686);
nand U10081 (N_10081,N_8459,N_8486);
nand U10082 (N_10082,N_8451,N_8973);
and U10083 (N_10083,N_8463,N_9203);
and U10084 (N_10084,N_8788,N_8987);
or U10085 (N_10085,N_9198,N_9315);
nor U10086 (N_10086,N_9486,N_8457);
nor U10087 (N_10087,N_9149,N_9256);
and U10088 (N_10088,N_8961,N_8937);
nand U10089 (N_10089,N_8545,N_9160);
or U10090 (N_10090,N_8971,N_9499);
xor U10091 (N_10091,N_8560,N_8534);
xnor U10092 (N_10092,N_9419,N_8405);
nand U10093 (N_10093,N_8882,N_9278);
nand U10094 (N_10094,N_8498,N_8420);
xor U10095 (N_10095,N_9095,N_8799);
xnor U10096 (N_10096,N_9303,N_8948);
xor U10097 (N_10097,N_8708,N_8561);
nor U10098 (N_10098,N_8931,N_9526);
and U10099 (N_10099,N_9427,N_9288);
and U10100 (N_10100,N_8747,N_8936);
nand U10101 (N_10101,N_8819,N_9492);
nor U10102 (N_10102,N_9349,N_9360);
or U10103 (N_10103,N_9253,N_9382);
and U10104 (N_10104,N_9411,N_8460);
nor U10105 (N_10105,N_8986,N_8595);
xnor U10106 (N_10106,N_8401,N_8876);
and U10107 (N_10107,N_8643,N_9388);
xor U10108 (N_10108,N_8475,N_9369);
nor U10109 (N_10109,N_8762,N_9216);
or U10110 (N_10110,N_8509,N_8612);
and U10111 (N_10111,N_8852,N_8738);
xor U10112 (N_10112,N_8980,N_9599);
xor U10113 (N_10113,N_8865,N_8404);
xor U10114 (N_10114,N_8538,N_9545);
and U10115 (N_10115,N_8807,N_9284);
nor U10116 (N_10116,N_8439,N_9581);
nor U10117 (N_10117,N_8823,N_9489);
and U10118 (N_10118,N_8774,N_9176);
or U10119 (N_10119,N_8412,N_8569);
nand U10120 (N_10120,N_9165,N_8925);
and U10121 (N_10121,N_8848,N_9080);
nand U10122 (N_10122,N_9013,N_8550);
and U10123 (N_10123,N_9378,N_8506);
or U10124 (N_10124,N_9500,N_8597);
and U10125 (N_10125,N_9540,N_9307);
nand U10126 (N_10126,N_9072,N_8619);
or U10127 (N_10127,N_8795,N_9084);
xor U10128 (N_10128,N_9373,N_8677);
nor U10129 (N_10129,N_9058,N_9069);
nor U10130 (N_10130,N_9516,N_8635);
and U10131 (N_10131,N_9167,N_8825);
nor U10132 (N_10132,N_9437,N_9085);
and U10133 (N_10133,N_8450,N_9009);
or U10134 (N_10134,N_9561,N_9070);
xor U10135 (N_10135,N_8683,N_8668);
xnor U10136 (N_10136,N_9215,N_8707);
nor U10137 (N_10137,N_9145,N_9045);
or U10138 (N_10138,N_9503,N_9366);
or U10139 (N_10139,N_8695,N_9299);
xor U10140 (N_10140,N_9212,N_8464);
or U10141 (N_10141,N_8887,N_8863);
xnor U10142 (N_10142,N_9022,N_9460);
nor U10143 (N_10143,N_9064,N_9376);
xor U10144 (N_10144,N_8518,N_8618);
nand U10145 (N_10145,N_8783,N_9586);
and U10146 (N_10146,N_8721,N_9368);
or U10147 (N_10147,N_9119,N_9479);
and U10148 (N_10148,N_9274,N_8985);
or U10149 (N_10149,N_8476,N_8705);
xor U10150 (N_10150,N_8582,N_9233);
or U10151 (N_10151,N_8908,N_9140);
and U10152 (N_10152,N_8633,N_9344);
nor U10153 (N_10153,N_9325,N_9387);
nand U10154 (N_10154,N_8642,N_8821);
or U10155 (N_10155,N_9155,N_8579);
and U10156 (N_10156,N_9137,N_8588);
nor U10157 (N_10157,N_8806,N_9068);
nand U10158 (N_10158,N_8966,N_9456);
xor U10159 (N_10159,N_8812,N_8999);
xor U10160 (N_10160,N_9231,N_9294);
and U10161 (N_10161,N_9240,N_9482);
xnor U10162 (N_10162,N_8739,N_9071);
and U10163 (N_10163,N_9319,N_9417);
nor U10164 (N_10164,N_8718,N_9375);
and U10165 (N_10165,N_9416,N_9089);
and U10166 (N_10166,N_8872,N_8572);
nor U10167 (N_10167,N_8429,N_9423);
and U10168 (N_10168,N_9191,N_9345);
or U10169 (N_10169,N_8490,N_9405);
nand U10170 (N_10170,N_9044,N_8830);
xnor U10171 (N_10171,N_8680,N_8915);
or U10172 (N_10172,N_8462,N_8711);
nand U10173 (N_10173,N_8674,N_8654);
and U10174 (N_10174,N_8765,N_8851);
and U10175 (N_10175,N_9015,N_8856);
nor U10176 (N_10176,N_8878,N_8725);
nor U10177 (N_10177,N_8402,N_8605);
nor U10178 (N_10178,N_8781,N_8914);
xnor U10179 (N_10179,N_8517,N_8930);
and U10180 (N_10180,N_8890,N_8933);
nand U10181 (N_10181,N_8772,N_8853);
or U10182 (N_10182,N_9166,N_9236);
xnor U10183 (N_10183,N_9422,N_9580);
or U10184 (N_10184,N_8414,N_8554);
nand U10185 (N_10185,N_9309,N_8528);
nor U10186 (N_10186,N_8953,N_8646);
nand U10187 (N_10187,N_9386,N_9177);
or U10188 (N_10188,N_8503,N_9529);
and U10189 (N_10189,N_8672,N_9585);
xnor U10190 (N_10190,N_8702,N_9036);
nand U10191 (N_10191,N_9598,N_9239);
and U10192 (N_10192,N_9359,N_9156);
nor U10193 (N_10193,N_9403,N_8952);
xnor U10194 (N_10194,N_8636,N_8699);
and U10195 (N_10195,N_8913,N_9542);
nor U10196 (N_10196,N_8840,N_8723);
or U10197 (N_10197,N_8949,N_9436);
and U10198 (N_10198,N_8417,N_8411);
xor U10199 (N_10199,N_9051,N_8899);
nand U10200 (N_10200,N_9124,N_8619);
nor U10201 (N_10201,N_9338,N_9478);
nor U10202 (N_10202,N_8438,N_9327);
and U10203 (N_10203,N_9552,N_9274);
or U10204 (N_10204,N_9462,N_8467);
nor U10205 (N_10205,N_8685,N_9193);
xnor U10206 (N_10206,N_9503,N_8600);
nand U10207 (N_10207,N_9126,N_8899);
nand U10208 (N_10208,N_9548,N_8766);
or U10209 (N_10209,N_8654,N_8500);
or U10210 (N_10210,N_8657,N_9315);
nand U10211 (N_10211,N_9432,N_9195);
or U10212 (N_10212,N_8589,N_8839);
or U10213 (N_10213,N_8818,N_9164);
nor U10214 (N_10214,N_9582,N_8984);
nor U10215 (N_10215,N_9492,N_9444);
nor U10216 (N_10216,N_8699,N_8650);
nor U10217 (N_10217,N_9209,N_9498);
xor U10218 (N_10218,N_8790,N_8822);
nor U10219 (N_10219,N_8471,N_9166);
and U10220 (N_10220,N_9488,N_8716);
nand U10221 (N_10221,N_9029,N_8540);
nor U10222 (N_10222,N_9136,N_8515);
nand U10223 (N_10223,N_9088,N_9548);
nand U10224 (N_10224,N_8467,N_8714);
or U10225 (N_10225,N_8900,N_9151);
and U10226 (N_10226,N_9085,N_9441);
xnor U10227 (N_10227,N_8594,N_8939);
or U10228 (N_10228,N_9031,N_9275);
xor U10229 (N_10229,N_9201,N_9479);
nor U10230 (N_10230,N_8968,N_8763);
xor U10231 (N_10231,N_8407,N_8651);
nand U10232 (N_10232,N_9376,N_8677);
nand U10233 (N_10233,N_8996,N_8902);
or U10234 (N_10234,N_9335,N_8966);
xnor U10235 (N_10235,N_9475,N_8976);
nand U10236 (N_10236,N_8941,N_9216);
or U10237 (N_10237,N_8809,N_8623);
and U10238 (N_10238,N_8429,N_9390);
nor U10239 (N_10239,N_9381,N_8528);
nand U10240 (N_10240,N_8465,N_9527);
nor U10241 (N_10241,N_8866,N_9097);
nor U10242 (N_10242,N_9388,N_8770);
or U10243 (N_10243,N_9525,N_9598);
and U10244 (N_10244,N_8894,N_8425);
or U10245 (N_10245,N_8869,N_8430);
nand U10246 (N_10246,N_9074,N_9463);
or U10247 (N_10247,N_9366,N_9078);
nand U10248 (N_10248,N_8892,N_9507);
and U10249 (N_10249,N_9119,N_9530);
or U10250 (N_10250,N_8512,N_9345);
and U10251 (N_10251,N_8746,N_8844);
or U10252 (N_10252,N_9490,N_9370);
and U10253 (N_10253,N_9374,N_8992);
xnor U10254 (N_10254,N_8969,N_9074);
xor U10255 (N_10255,N_8777,N_9021);
xor U10256 (N_10256,N_9171,N_8996);
nand U10257 (N_10257,N_9231,N_8508);
and U10258 (N_10258,N_8607,N_9339);
nand U10259 (N_10259,N_9085,N_9596);
and U10260 (N_10260,N_9386,N_8657);
and U10261 (N_10261,N_9554,N_9509);
nand U10262 (N_10262,N_8439,N_8621);
nand U10263 (N_10263,N_9194,N_9457);
nor U10264 (N_10264,N_9129,N_8673);
and U10265 (N_10265,N_8877,N_9291);
nor U10266 (N_10266,N_9383,N_8649);
nor U10267 (N_10267,N_9337,N_8612);
xor U10268 (N_10268,N_8925,N_9402);
nand U10269 (N_10269,N_9230,N_8822);
and U10270 (N_10270,N_9466,N_9176);
xnor U10271 (N_10271,N_9193,N_8944);
and U10272 (N_10272,N_9138,N_9139);
nor U10273 (N_10273,N_9461,N_8435);
xnor U10274 (N_10274,N_8923,N_9086);
and U10275 (N_10275,N_8549,N_9498);
xnor U10276 (N_10276,N_8972,N_9538);
or U10277 (N_10277,N_9213,N_9384);
or U10278 (N_10278,N_9032,N_9534);
or U10279 (N_10279,N_8564,N_8557);
and U10280 (N_10280,N_8728,N_9169);
nand U10281 (N_10281,N_9396,N_8520);
xor U10282 (N_10282,N_9268,N_8885);
xor U10283 (N_10283,N_9220,N_8579);
nor U10284 (N_10284,N_9530,N_9181);
nor U10285 (N_10285,N_9182,N_8667);
nand U10286 (N_10286,N_9442,N_9118);
xnor U10287 (N_10287,N_9576,N_9555);
and U10288 (N_10288,N_8870,N_9231);
and U10289 (N_10289,N_9375,N_9092);
nor U10290 (N_10290,N_8909,N_9519);
xnor U10291 (N_10291,N_9211,N_8877);
xor U10292 (N_10292,N_8997,N_9346);
xnor U10293 (N_10293,N_9304,N_9327);
nand U10294 (N_10294,N_9546,N_9201);
nor U10295 (N_10295,N_9409,N_8938);
xnor U10296 (N_10296,N_9275,N_9103);
nor U10297 (N_10297,N_8935,N_9599);
nor U10298 (N_10298,N_9307,N_9134);
nand U10299 (N_10299,N_8819,N_9497);
xnor U10300 (N_10300,N_9478,N_9083);
nor U10301 (N_10301,N_9493,N_9109);
nor U10302 (N_10302,N_8616,N_8836);
nand U10303 (N_10303,N_9477,N_8757);
xnor U10304 (N_10304,N_8446,N_8772);
xor U10305 (N_10305,N_8983,N_8500);
xnor U10306 (N_10306,N_9264,N_8827);
nor U10307 (N_10307,N_8420,N_8536);
or U10308 (N_10308,N_9032,N_9502);
xnor U10309 (N_10309,N_8980,N_8972);
or U10310 (N_10310,N_9595,N_9166);
xnor U10311 (N_10311,N_8931,N_8467);
and U10312 (N_10312,N_8732,N_8949);
xnor U10313 (N_10313,N_9542,N_8539);
xnor U10314 (N_10314,N_9455,N_9441);
nor U10315 (N_10315,N_9467,N_9498);
nor U10316 (N_10316,N_8440,N_9138);
nor U10317 (N_10317,N_8552,N_8908);
nand U10318 (N_10318,N_9050,N_8449);
xor U10319 (N_10319,N_9155,N_9156);
nand U10320 (N_10320,N_8406,N_8887);
and U10321 (N_10321,N_9028,N_9271);
and U10322 (N_10322,N_8912,N_9472);
and U10323 (N_10323,N_8445,N_9322);
nand U10324 (N_10324,N_8615,N_9489);
nand U10325 (N_10325,N_9126,N_8603);
nor U10326 (N_10326,N_8952,N_9373);
nand U10327 (N_10327,N_9086,N_8413);
nand U10328 (N_10328,N_8534,N_8618);
xor U10329 (N_10329,N_9383,N_8679);
nor U10330 (N_10330,N_9545,N_9047);
nor U10331 (N_10331,N_8530,N_9449);
xor U10332 (N_10332,N_9127,N_8753);
nand U10333 (N_10333,N_8540,N_9535);
xor U10334 (N_10334,N_9509,N_9562);
xor U10335 (N_10335,N_8971,N_8530);
or U10336 (N_10336,N_9193,N_9454);
xnor U10337 (N_10337,N_9468,N_8418);
or U10338 (N_10338,N_8912,N_8668);
nand U10339 (N_10339,N_8715,N_9377);
xnor U10340 (N_10340,N_8943,N_8416);
or U10341 (N_10341,N_8808,N_9550);
and U10342 (N_10342,N_8582,N_9469);
nor U10343 (N_10343,N_8557,N_9546);
or U10344 (N_10344,N_9489,N_9348);
and U10345 (N_10345,N_9406,N_9337);
nor U10346 (N_10346,N_9319,N_8737);
or U10347 (N_10347,N_8864,N_9158);
and U10348 (N_10348,N_9487,N_8467);
and U10349 (N_10349,N_9323,N_8843);
nor U10350 (N_10350,N_9562,N_9461);
and U10351 (N_10351,N_8982,N_8920);
or U10352 (N_10352,N_8550,N_8616);
nor U10353 (N_10353,N_8707,N_8643);
or U10354 (N_10354,N_8551,N_8963);
or U10355 (N_10355,N_9544,N_8695);
nor U10356 (N_10356,N_8498,N_9184);
and U10357 (N_10357,N_9267,N_8575);
nor U10358 (N_10358,N_8595,N_9504);
nor U10359 (N_10359,N_9413,N_8494);
nor U10360 (N_10360,N_9436,N_9299);
nor U10361 (N_10361,N_9563,N_8642);
nor U10362 (N_10362,N_9543,N_9246);
and U10363 (N_10363,N_9574,N_8760);
nand U10364 (N_10364,N_8645,N_8912);
nand U10365 (N_10365,N_9005,N_9200);
and U10366 (N_10366,N_8473,N_9344);
nand U10367 (N_10367,N_9029,N_8762);
xnor U10368 (N_10368,N_8433,N_9367);
xor U10369 (N_10369,N_8866,N_8642);
and U10370 (N_10370,N_9170,N_9023);
nand U10371 (N_10371,N_9015,N_8805);
or U10372 (N_10372,N_9014,N_9065);
xnor U10373 (N_10373,N_8936,N_8496);
nand U10374 (N_10374,N_8631,N_8884);
nand U10375 (N_10375,N_9170,N_9559);
and U10376 (N_10376,N_9028,N_8952);
or U10377 (N_10377,N_9372,N_8876);
and U10378 (N_10378,N_9235,N_9017);
and U10379 (N_10379,N_9585,N_9155);
xnor U10380 (N_10380,N_9086,N_9045);
nor U10381 (N_10381,N_9302,N_8797);
nand U10382 (N_10382,N_9512,N_8844);
nand U10383 (N_10383,N_8663,N_8725);
xor U10384 (N_10384,N_9022,N_9269);
nand U10385 (N_10385,N_8745,N_9336);
nor U10386 (N_10386,N_9134,N_9504);
nand U10387 (N_10387,N_9202,N_9215);
nor U10388 (N_10388,N_8724,N_8879);
and U10389 (N_10389,N_9223,N_8676);
or U10390 (N_10390,N_8537,N_9415);
and U10391 (N_10391,N_9436,N_8917);
nor U10392 (N_10392,N_8812,N_8664);
nor U10393 (N_10393,N_9029,N_8872);
and U10394 (N_10394,N_8545,N_8541);
nor U10395 (N_10395,N_8921,N_8861);
or U10396 (N_10396,N_8553,N_9522);
nand U10397 (N_10397,N_9488,N_8895);
and U10398 (N_10398,N_9209,N_8512);
and U10399 (N_10399,N_9202,N_9482);
nand U10400 (N_10400,N_9510,N_9418);
xor U10401 (N_10401,N_9391,N_8678);
and U10402 (N_10402,N_9012,N_9491);
or U10403 (N_10403,N_9421,N_9527);
or U10404 (N_10404,N_8891,N_9499);
nor U10405 (N_10405,N_8908,N_8446);
or U10406 (N_10406,N_8682,N_8988);
and U10407 (N_10407,N_9071,N_9432);
nor U10408 (N_10408,N_9024,N_8880);
nand U10409 (N_10409,N_8696,N_9527);
nand U10410 (N_10410,N_9169,N_9446);
nand U10411 (N_10411,N_9185,N_9056);
and U10412 (N_10412,N_8745,N_8573);
nor U10413 (N_10413,N_9378,N_8928);
nor U10414 (N_10414,N_9270,N_9364);
xor U10415 (N_10415,N_8589,N_9007);
nor U10416 (N_10416,N_8887,N_8685);
nand U10417 (N_10417,N_9456,N_8963);
or U10418 (N_10418,N_9279,N_8486);
nand U10419 (N_10419,N_8957,N_8418);
nand U10420 (N_10420,N_8511,N_9571);
nand U10421 (N_10421,N_8745,N_8963);
and U10422 (N_10422,N_8952,N_9045);
and U10423 (N_10423,N_9546,N_9188);
xor U10424 (N_10424,N_8881,N_9354);
nand U10425 (N_10425,N_9416,N_9210);
and U10426 (N_10426,N_8705,N_9250);
xor U10427 (N_10427,N_9392,N_8920);
nand U10428 (N_10428,N_9489,N_9287);
nand U10429 (N_10429,N_9575,N_9111);
nand U10430 (N_10430,N_8425,N_8490);
nand U10431 (N_10431,N_8644,N_8640);
nor U10432 (N_10432,N_9576,N_9365);
or U10433 (N_10433,N_8879,N_8514);
nor U10434 (N_10434,N_8597,N_8796);
and U10435 (N_10435,N_9266,N_9540);
nor U10436 (N_10436,N_8641,N_9439);
nand U10437 (N_10437,N_8594,N_8971);
xnor U10438 (N_10438,N_8981,N_8473);
and U10439 (N_10439,N_8960,N_8591);
and U10440 (N_10440,N_9177,N_8992);
nand U10441 (N_10441,N_8414,N_9306);
nor U10442 (N_10442,N_8847,N_9290);
nand U10443 (N_10443,N_9546,N_8402);
nand U10444 (N_10444,N_8702,N_8519);
nor U10445 (N_10445,N_9014,N_9191);
nor U10446 (N_10446,N_9098,N_9204);
or U10447 (N_10447,N_9574,N_9446);
or U10448 (N_10448,N_9335,N_9035);
xor U10449 (N_10449,N_8661,N_9151);
xnor U10450 (N_10450,N_9457,N_8687);
nand U10451 (N_10451,N_9463,N_9157);
xor U10452 (N_10452,N_8812,N_8590);
nand U10453 (N_10453,N_9494,N_9112);
and U10454 (N_10454,N_9295,N_8825);
xnor U10455 (N_10455,N_9358,N_8450);
or U10456 (N_10456,N_8745,N_8511);
nor U10457 (N_10457,N_9568,N_8531);
and U10458 (N_10458,N_9221,N_8973);
nor U10459 (N_10459,N_9026,N_9418);
or U10460 (N_10460,N_9082,N_9516);
nor U10461 (N_10461,N_8933,N_9262);
nand U10462 (N_10462,N_8838,N_9517);
nor U10463 (N_10463,N_9343,N_9080);
nor U10464 (N_10464,N_9447,N_9319);
or U10465 (N_10465,N_8499,N_9070);
xnor U10466 (N_10466,N_8672,N_8571);
and U10467 (N_10467,N_9190,N_8747);
and U10468 (N_10468,N_9112,N_9276);
nor U10469 (N_10469,N_8683,N_8794);
nand U10470 (N_10470,N_9043,N_8976);
nand U10471 (N_10471,N_8427,N_8861);
nor U10472 (N_10472,N_9118,N_9302);
nor U10473 (N_10473,N_9489,N_8918);
xnor U10474 (N_10474,N_8514,N_9130);
nor U10475 (N_10475,N_8749,N_9051);
and U10476 (N_10476,N_9085,N_8814);
nor U10477 (N_10477,N_8491,N_9280);
nand U10478 (N_10478,N_9097,N_8471);
xor U10479 (N_10479,N_8893,N_9216);
or U10480 (N_10480,N_8829,N_8893);
and U10481 (N_10481,N_8490,N_9555);
nand U10482 (N_10482,N_8903,N_9033);
xor U10483 (N_10483,N_8724,N_8499);
nand U10484 (N_10484,N_8769,N_8911);
nand U10485 (N_10485,N_8457,N_8837);
nand U10486 (N_10486,N_9585,N_8597);
or U10487 (N_10487,N_9551,N_8966);
or U10488 (N_10488,N_9374,N_9079);
and U10489 (N_10489,N_8988,N_8592);
nand U10490 (N_10490,N_9120,N_9384);
nand U10491 (N_10491,N_8891,N_8423);
and U10492 (N_10492,N_8494,N_9324);
xnor U10493 (N_10493,N_8952,N_9571);
or U10494 (N_10494,N_8626,N_8657);
or U10495 (N_10495,N_8701,N_9553);
nand U10496 (N_10496,N_9519,N_9500);
nand U10497 (N_10497,N_9193,N_8715);
xor U10498 (N_10498,N_8807,N_9052);
nand U10499 (N_10499,N_9160,N_9318);
nand U10500 (N_10500,N_8879,N_9317);
xnor U10501 (N_10501,N_8461,N_8997);
nor U10502 (N_10502,N_9519,N_8904);
and U10503 (N_10503,N_8601,N_9117);
nand U10504 (N_10504,N_8780,N_9030);
or U10505 (N_10505,N_8995,N_8511);
or U10506 (N_10506,N_8415,N_8564);
xor U10507 (N_10507,N_9179,N_8792);
nand U10508 (N_10508,N_9452,N_8585);
nor U10509 (N_10509,N_9195,N_9402);
xor U10510 (N_10510,N_9097,N_9223);
and U10511 (N_10511,N_8981,N_8877);
nand U10512 (N_10512,N_8972,N_9035);
xor U10513 (N_10513,N_8812,N_9323);
and U10514 (N_10514,N_8499,N_9338);
and U10515 (N_10515,N_9423,N_9402);
nand U10516 (N_10516,N_8524,N_9062);
and U10517 (N_10517,N_9145,N_8610);
and U10518 (N_10518,N_8608,N_9013);
and U10519 (N_10519,N_9265,N_9287);
xnor U10520 (N_10520,N_9160,N_8588);
or U10521 (N_10521,N_8903,N_9543);
or U10522 (N_10522,N_9425,N_8622);
nand U10523 (N_10523,N_8970,N_8517);
and U10524 (N_10524,N_8565,N_9000);
nor U10525 (N_10525,N_8683,N_9416);
xor U10526 (N_10526,N_9305,N_9004);
or U10527 (N_10527,N_9081,N_9447);
nand U10528 (N_10528,N_8414,N_8484);
xor U10529 (N_10529,N_9527,N_9188);
and U10530 (N_10530,N_9366,N_8671);
and U10531 (N_10531,N_8574,N_8745);
and U10532 (N_10532,N_8865,N_9271);
or U10533 (N_10533,N_9466,N_9185);
or U10534 (N_10534,N_9275,N_8564);
nand U10535 (N_10535,N_9514,N_8976);
xor U10536 (N_10536,N_9153,N_9555);
nor U10537 (N_10537,N_9100,N_8552);
xor U10538 (N_10538,N_8900,N_8855);
or U10539 (N_10539,N_9103,N_9358);
xor U10540 (N_10540,N_8961,N_9144);
and U10541 (N_10541,N_9344,N_8452);
and U10542 (N_10542,N_8597,N_9378);
or U10543 (N_10543,N_9171,N_9000);
xor U10544 (N_10544,N_9169,N_9164);
nor U10545 (N_10545,N_8502,N_9488);
or U10546 (N_10546,N_9111,N_9570);
or U10547 (N_10547,N_9436,N_8964);
and U10548 (N_10548,N_8480,N_9359);
or U10549 (N_10549,N_8777,N_8842);
nor U10550 (N_10550,N_9073,N_9528);
or U10551 (N_10551,N_9580,N_9393);
nand U10552 (N_10552,N_8685,N_9514);
nor U10553 (N_10553,N_9165,N_9418);
xnor U10554 (N_10554,N_9414,N_9480);
xnor U10555 (N_10555,N_9104,N_8842);
nor U10556 (N_10556,N_8778,N_9358);
and U10557 (N_10557,N_9222,N_8653);
or U10558 (N_10558,N_8595,N_8612);
xor U10559 (N_10559,N_8680,N_9499);
nor U10560 (N_10560,N_8676,N_9426);
and U10561 (N_10561,N_8794,N_8978);
xnor U10562 (N_10562,N_8882,N_9060);
and U10563 (N_10563,N_8699,N_9543);
or U10564 (N_10564,N_9026,N_9584);
nand U10565 (N_10565,N_9501,N_8703);
xnor U10566 (N_10566,N_9202,N_8942);
xnor U10567 (N_10567,N_9459,N_8916);
nor U10568 (N_10568,N_9483,N_9323);
xnor U10569 (N_10569,N_9487,N_9366);
nor U10570 (N_10570,N_9219,N_8494);
nor U10571 (N_10571,N_9061,N_8865);
nor U10572 (N_10572,N_8484,N_9402);
nand U10573 (N_10573,N_9095,N_8568);
and U10574 (N_10574,N_9511,N_8881);
and U10575 (N_10575,N_9486,N_9567);
nand U10576 (N_10576,N_8601,N_9068);
xor U10577 (N_10577,N_8535,N_9154);
xnor U10578 (N_10578,N_9176,N_8754);
and U10579 (N_10579,N_9511,N_8654);
nor U10580 (N_10580,N_8640,N_9566);
nor U10581 (N_10581,N_9108,N_9040);
or U10582 (N_10582,N_9388,N_9062);
nor U10583 (N_10583,N_8987,N_8472);
nand U10584 (N_10584,N_9408,N_8934);
nand U10585 (N_10585,N_8956,N_9234);
nand U10586 (N_10586,N_8980,N_9123);
or U10587 (N_10587,N_9223,N_9171);
nor U10588 (N_10588,N_9062,N_8438);
or U10589 (N_10589,N_8822,N_9568);
or U10590 (N_10590,N_9455,N_8580);
and U10591 (N_10591,N_8962,N_8899);
or U10592 (N_10592,N_8752,N_9432);
and U10593 (N_10593,N_9120,N_8532);
xnor U10594 (N_10594,N_8658,N_9299);
or U10595 (N_10595,N_8631,N_9437);
or U10596 (N_10596,N_9577,N_8680);
and U10597 (N_10597,N_8942,N_9560);
or U10598 (N_10598,N_9114,N_9155);
or U10599 (N_10599,N_9294,N_8533);
nor U10600 (N_10600,N_8984,N_8809);
nor U10601 (N_10601,N_9285,N_8618);
nand U10602 (N_10602,N_9171,N_8740);
and U10603 (N_10603,N_8516,N_8618);
nor U10604 (N_10604,N_8793,N_8623);
xnor U10605 (N_10605,N_8755,N_9134);
nand U10606 (N_10606,N_8734,N_8861);
or U10607 (N_10607,N_9490,N_9522);
xnor U10608 (N_10608,N_9469,N_8660);
nand U10609 (N_10609,N_8421,N_8571);
nor U10610 (N_10610,N_9217,N_8714);
nor U10611 (N_10611,N_8898,N_9254);
xnor U10612 (N_10612,N_9519,N_9415);
and U10613 (N_10613,N_9467,N_8484);
or U10614 (N_10614,N_9481,N_8977);
nor U10615 (N_10615,N_8660,N_9093);
nand U10616 (N_10616,N_9100,N_8738);
or U10617 (N_10617,N_8963,N_9444);
and U10618 (N_10618,N_9517,N_8872);
or U10619 (N_10619,N_8682,N_8771);
xor U10620 (N_10620,N_9439,N_9242);
or U10621 (N_10621,N_8823,N_9454);
xor U10622 (N_10622,N_8885,N_8782);
or U10623 (N_10623,N_9268,N_8838);
or U10624 (N_10624,N_9545,N_8748);
or U10625 (N_10625,N_8610,N_8468);
and U10626 (N_10626,N_9246,N_9553);
nand U10627 (N_10627,N_9361,N_8641);
nor U10628 (N_10628,N_8570,N_8747);
nor U10629 (N_10629,N_9301,N_9181);
and U10630 (N_10630,N_8513,N_9180);
nor U10631 (N_10631,N_8522,N_8547);
and U10632 (N_10632,N_9198,N_9490);
xnor U10633 (N_10633,N_9061,N_8700);
xnor U10634 (N_10634,N_8959,N_8734);
nand U10635 (N_10635,N_9271,N_8643);
or U10636 (N_10636,N_8901,N_9431);
nor U10637 (N_10637,N_8979,N_9562);
or U10638 (N_10638,N_8448,N_9287);
xor U10639 (N_10639,N_9422,N_9117);
nor U10640 (N_10640,N_9313,N_8846);
nand U10641 (N_10641,N_8944,N_9257);
nor U10642 (N_10642,N_8418,N_8505);
nor U10643 (N_10643,N_9595,N_9590);
xor U10644 (N_10644,N_8886,N_8596);
xor U10645 (N_10645,N_8686,N_8670);
xnor U10646 (N_10646,N_9376,N_8957);
or U10647 (N_10647,N_8939,N_8908);
or U10648 (N_10648,N_8682,N_9120);
or U10649 (N_10649,N_9214,N_9578);
nand U10650 (N_10650,N_9546,N_9537);
or U10651 (N_10651,N_9085,N_8637);
xor U10652 (N_10652,N_9579,N_8880);
and U10653 (N_10653,N_9244,N_9361);
nand U10654 (N_10654,N_8580,N_8442);
xor U10655 (N_10655,N_9020,N_8875);
and U10656 (N_10656,N_9453,N_9193);
xor U10657 (N_10657,N_8826,N_9383);
and U10658 (N_10658,N_9374,N_8579);
or U10659 (N_10659,N_9574,N_9293);
and U10660 (N_10660,N_8984,N_8910);
or U10661 (N_10661,N_9595,N_8577);
nand U10662 (N_10662,N_8836,N_8863);
nand U10663 (N_10663,N_9024,N_9247);
nor U10664 (N_10664,N_8543,N_8982);
nand U10665 (N_10665,N_8742,N_8986);
or U10666 (N_10666,N_8657,N_9093);
and U10667 (N_10667,N_8849,N_9239);
xnor U10668 (N_10668,N_9341,N_9506);
nor U10669 (N_10669,N_9179,N_9158);
nand U10670 (N_10670,N_8824,N_8752);
nand U10671 (N_10671,N_8550,N_9117);
xnor U10672 (N_10672,N_9133,N_9012);
and U10673 (N_10673,N_9555,N_9192);
and U10674 (N_10674,N_8781,N_8968);
and U10675 (N_10675,N_9269,N_8966);
and U10676 (N_10676,N_9325,N_8757);
or U10677 (N_10677,N_8789,N_9242);
xnor U10678 (N_10678,N_8689,N_9479);
nand U10679 (N_10679,N_8917,N_9273);
xor U10680 (N_10680,N_8867,N_8577);
xor U10681 (N_10681,N_8455,N_8872);
or U10682 (N_10682,N_9224,N_8407);
or U10683 (N_10683,N_9305,N_9451);
or U10684 (N_10684,N_8441,N_9015);
xor U10685 (N_10685,N_8954,N_8871);
nor U10686 (N_10686,N_8901,N_9384);
nor U10687 (N_10687,N_8770,N_8792);
nor U10688 (N_10688,N_9119,N_8541);
xor U10689 (N_10689,N_9420,N_9144);
nand U10690 (N_10690,N_9306,N_9328);
and U10691 (N_10691,N_8695,N_8538);
or U10692 (N_10692,N_9578,N_9587);
xnor U10693 (N_10693,N_8659,N_9086);
and U10694 (N_10694,N_9126,N_9339);
or U10695 (N_10695,N_8981,N_8652);
xnor U10696 (N_10696,N_8453,N_8428);
and U10697 (N_10697,N_9199,N_9208);
and U10698 (N_10698,N_9506,N_9518);
nand U10699 (N_10699,N_8618,N_9357);
xnor U10700 (N_10700,N_8401,N_9533);
and U10701 (N_10701,N_8598,N_9147);
nor U10702 (N_10702,N_9451,N_8435);
and U10703 (N_10703,N_8528,N_9249);
nor U10704 (N_10704,N_8548,N_8579);
nor U10705 (N_10705,N_8728,N_9427);
or U10706 (N_10706,N_8932,N_9285);
nand U10707 (N_10707,N_9082,N_9189);
and U10708 (N_10708,N_8537,N_9252);
or U10709 (N_10709,N_9364,N_8717);
or U10710 (N_10710,N_8431,N_8442);
nand U10711 (N_10711,N_9036,N_8540);
nand U10712 (N_10712,N_9437,N_8413);
and U10713 (N_10713,N_8878,N_9436);
nor U10714 (N_10714,N_9558,N_9212);
nand U10715 (N_10715,N_9126,N_9569);
nor U10716 (N_10716,N_9115,N_8565);
nor U10717 (N_10717,N_9424,N_9489);
nor U10718 (N_10718,N_8959,N_8736);
xnor U10719 (N_10719,N_9449,N_8545);
nand U10720 (N_10720,N_9200,N_8945);
xor U10721 (N_10721,N_8464,N_9279);
or U10722 (N_10722,N_8620,N_9100);
and U10723 (N_10723,N_8643,N_8960);
or U10724 (N_10724,N_8442,N_9394);
xnor U10725 (N_10725,N_8443,N_8625);
nand U10726 (N_10726,N_9190,N_9423);
nand U10727 (N_10727,N_8496,N_9080);
and U10728 (N_10728,N_9599,N_9376);
or U10729 (N_10729,N_8880,N_9477);
xor U10730 (N_10730,N_9273,N_9482);
nor U10731 (N_10731,N_9348,N_8419);
xnor U10732 (N_10732,N_9014,N_8655);
nand U10733 (N_10733,N_8611,N_9075);
or U10734 (N_10734,N_9332,N_8553);
and U10735 (N_10735,N_9496,N_9400);
nand U10736 (N_10736,N_8554,N_9398);
xnor U10737 (N_10737,N_8845,N_9515);
and U10738 (N_10738,N_8855,N_8761);
nand U10739 (N_10739,N_8802,N_8736);
nand U10740 (N_10740,N_9357,N_8416);
or U10741 (N_10741,N_8849,N_8419);
nor U10742 (N_10742,N_8938,N_8753);
and U10743 (N_10743,N_8734,N_8507);
or U10744 (N_10744,N_9344,N_8945);
xnor U10745 (N_10745,N_9294,N_9060);
and U10746 (N_10746,N_8990,N_9008);
nand U10747 (N_10747,N_8923,N_9210);
nor U10748 (N_10748,N_9503,N_9059);
nand U10749 (N_10749,N_9065,N_8659);
and U10750 (N_10750,N_8947,N_8621);
or U10751 (N_10751,N_8955,N_8903);
nand U10752 (N_10752,N_9529,N_9344);
nor U10753 (N_10753,N_8730,N_8940);
nand U10754 (N_10754,N_9271,N_8417);
nand U10755 (N_10755,N_9397,N_9207);
and U10756 (N_10756,N_9407,N_9458);
or U10757 (N_10757,N_8433,N_9269);
and U10758 (N_10758,N_9081,N_8989);
nor U10759 (N_10759,N_9132,N_8414);
xor U10760 (N_10760,N_8970,N_9517);
nand U10761 (N_10761,N_8439,N_9491);
or U10762 (N_10762,N_8891,N_9327);
or U10763 (N_10763,N_9324,N_8681);
nand U10764 (N_10764,N_9395,N_9586);
or U10765 (N_10765,N_9505,N_8723);
xor U10766 (N_10766,N_9349,N_8692);
and U10767 (N_10767,N_9587,N_9246);
xor U10768 (N_10768,N_9471,N_8815);
nand U10769 (N_10769,N_9414,N_8540);
nand U10770 (N_10770,N_9017,N_8836);
nand U10771 (N_10771,N_9528,N_9444);
and U10772 (N_10772,N_8543,N_9449);
xnor U10773 (N_10773,N_8630,N_8619);
nand U10774 (N_10774,N_9159,N_9399);
nor U10775 (N_10775,N_9148,N_9126);
nand U10776 (N_10776,N_8609,N_9176);
nand U10777 (N_10777,N_9014,N_8834);
or U10778 (N_10778,N_8450,N_9453);
or U10779 (N_10779,N_9474,N_8821);
xor U10780 (N_10780,N_9446,N_8492);
xnor U10781 (N_10781,N_9592,N_9229);
nor U10782 (N_10782,N_9216,N_9418);
nand U10783 (N_10783,N_9119,N_8493);
or U10784 (N_10784,N_9495,N_8582);
xor U10785 (N_10785,N_9170,N_9124);
nand U10786 (N_10786,N_8771,N_8491);
nand U10787 (N_10787,N_9064,N_9399);
nand U10788 (N_10788,N_9309,N_9123);
nand U10789 (N_10789,N_8989,N_8529);
xor U10790 (N_10790,N_9165,N_8490);
or U10791 (N_10791,N_8865,N_9127);
nand U10792 (N_10792,N_9268,N_8678);
nand U10793 (N_10793,N_9286,N_9499);
xor U10794 (N_10794,N_9524,N_9055);
xnor U10795 (N_10795,N_8984,N_8739);
nor U10796 (N_10796,N_9373,N_9393);
xor U10797 (N_10797,N_8693,N_8408);
and U10798 (N_10798,N_9544,N_8944);
and U10799 (N_10799,N_8995,N_8640);
nor U10800 (N_10800,N_10042,N_10149);
nand U10801 (N_10801,N_10299,N_9903);
nand U10802 (N_10802,N_10267,N_9651);
nand U10803 (N_10803,N_9889,N_10026);
nor U10804 (N_10804,N_9860,N_10719);
nor U10805 (N_10805,N_10402,N_10414);
nor U10806 (N_10806,N_10656,N_10269);
xnor U10807 (N_10807,N_10016,N_10253);
nand U10808 (N_10808,N_10668,N_10505);
nor U10809 (N_10809,N_9715,N_10798);
xnor U10810 (N_10810,N_9692,N_10660);
nand U10811 (N_10811,N_10006,N_10617);
and U10812 (N_10812,N_9719,N_10662);
nor U10813 (N_10813,N_9825,N_9699);
nor U10814 (N_10814,N_10019,N_10454);
nand U10815 (N_10815,N_10429,N_9911);
nor U10816 (N_10816,N_9686,N_10612);
nor U10817 (N_10817,N_9707,N_10430);
or U10818 (N_10818,N_10121,N_10210);
and U10819 (N_10819,N_9724,N_10373);
nand U10820 (N_10820,N_10475,N_10371);
xor U10821 (N_10821,N_10455,N_9872);
or U10822 (N_10822,N_9722,N_10559);
nand U10823 (N_10823,N_9988,N_10565);
nor U10824 (N_10824,N_10644,N_10465);
and U10825 (N_10825,N_10178,N_10534);
nor U10826 (N_10826,N_10227,N_10793);
and U10827 (N_10827,N_10300,N_10199);
and U10828 (N_10828,N_9972,N_10084);
nand U10829 (N_10829,N_10033,N_10519);
xor U10830 (N_10830,N_10650,N_9964);
nor U10831 (N_10831,N_9613,N_9611);
and U10832 (N_10832,N_10419,N_10604);
xnor U10833 (N_10833,N_9892,N_9704);
nor U10834 (N_10834,N_10352,N_9637);
nor U10835 (N_10835,N_9817,N_10120);
nand U10836 (N_10836,N_10567,N_10574);
xnor U10837 (N_10837,N_10376,N_10637);
and U10838 (N_10838,N_9734,N_9682);
nor U10839 (N_10839,N_9891,N_10357);
nand U10840 (N_10840,N_10052,N_9841);
and U10841 (N_10841,N_10331,N_10190);
xor U10842 (N_10842,N_10374,N_10634);
nor U10843 (N_10843,N_10128,N_9826);
and U10844 (N_10844,N_10593,N_9886);
nor U10845 (N_10845,N_9946,N_9738);
and U10846 (N_10846,N_9997,N_9862);
and U10847 (N_10847,N_10628,N_9920);
nand U10848 (N_10848,N_10720,N_9929);
nand U10849 (N_10849,N_10704,N_9635);
or U10850 (N_10850,N_9813,N_10417);
nand U10851 (N_10851,N_9740,N_10181);
and U10852 (N_10852,N_10481,N_9705);
xnor U10853 (N_10853,N_10492,N_10462);
nand U10854 (N_10854,N_10754,N_10759);
and U10855 (N_10855,N_10609,N_9777);
or U10856 (N_10856,N_10447,N_9633);
and U10857 (N_10857,N_9626,N_10692);
nand U10858 (N_10858,N_10770,N_10170);
nand U10859 (N_10859,N_10551,N_9761);
nor U10860 (N_10860,N_10356,N_10147);
xor U10861 (N_10861,N_10472,N_10739);
and U10862 (N_10862,N_9905,N_10520);
nor U10863 (N_10863,N_9880,N_10048);
nand U10864 (N_10864,N_10530,N_10276);
and U10865 (N_10865,N_10151,N_9876);
xor U10866 (N_10866,N_10708,N_10760);
and U10867 (N_10867,N_10485,N_10382);
nor U10868 (N_10868,N_10761,N_10467);
nor U10869 (N_10869,N_10744,N_10339);
and U10870 (N_10870,N_9790,N_9695);
nor U10871 (N_10871,N_9983,N_10513);
and U10872 (N_10872,N_10018,N_10316);
or U10873 (N_10873,N_10499,N_10030);
or U10874 (N_10874,N_10358,N_10561);
or U10875 (N_10875,N_9853,N_10333);
nor U10876 (N_10876,N_10642,N_10444);
nand U10877 (N_10877,N_9610,N_9832);
and U10878 (N_10878,N_10731,N_10257);
xor U10879 (N_10879,N_10723,N_10610);
xnor U10880 (N_10880,N_10307,N_10193);
nand U10881 (N_10881,N_10289,N_10137);
nor U10882 (N_10882,N_10221,N_10091);
and U10883 (N_10883,N_10491,N_9622);
and U10884 (N_10884,N_9652,N_10431);
nor U10885 (N_10885,N_10787,N_9602);
and U10886 (N_10886,N_10581,N_10734);
or U10887 (N_10887,N_10661,N_9775);
xor U10888 (N_10888,N_10409,N_10663);
xnor U10889 (N_10889,N_9787,N_9956);
nand U10890 (N_10890,N_10456,N_9857);
nand U10891 (N_10891,N_10112,N_10272);
nand U10892 (N_10892,N_9665,N_10250);
xnor U10893 (N_10893,N_10284,N_9882);
and U10894 (N_10894,N_10405,N_9835);
or U10895 (N_10895,N_9642,N_10397);
or U10896 (N_10896,N_10126,N_9819);
nor U10897 (N_10897,N_9907,N_10039);
nand U10898 (N_10898,N_10675,N_10435);
xor U10899 (N_10899,N_10746,N_10175);
and U10900 (N_10900,N_10649,N_10566);
xnor U10901 (N_10901,N_9728,N_9918);
nor U10902 (N_10902,N_10387,N_10424);
or U10903 (N_10903,N_9684,N_10599);
and U10904 (N_10904,N_10647,N_10434);
and U10905 (N_10905,N_9921,N_9914);
nor U10906 (N_10906,N_9890,N_10075);
nand U10907 (N_10907,N_10498,N_9609);
or U10908 (N_10908,N_10234,N_10631);
nand U10909 (N_10909,N_10283,N_9879);
nor U10910 (N_10910,N_9896,N_10230);
nor U10911 (N_10911,N_9616,N_10047);
nand U10912 (N_10912,N_9638,N_10068);
xor U10913 (N_10913,N_9716,N_10347);
nor U10914 (N_10914,N_10304,N_9676);
nand U10915 (N_10915,N_10712,N_10263);
xor U10916 (N_10916,N_10674,N_10482);
and U10917 (N_10917,N_10334,N_9621);
nor U10918 (N_10918,N_9690,N_10738);
nor U10919 (N_10919,N_10683,N_10515);
nor U10920 (N_10920,N_10555,N_10682);
nor U10921 (N_10921,N_10654,N_9623);
nand U10922 (N_10922,N_9675,N_10058);
nand U10923 (N_10923,N_9884,N_10401);
nor U10924 (N_10924,N_10032,N_9978);
or U10925 (N_10925,N_10672,N_10423);
and U10926 (N_10926,N_10632,N_9687);
and U10927 (N_10927,N_9847,N_9620);
xor U10928 (N_10928,N_10527,N_9805);
nor U10929 (N_10929,N_10557,N_9974);
xnor U10930 (N_10930,N_10224,N_10594);
or U10931 (N_10931,N_10422,N_9669);
and U10932 (N_10932,N_9680,N_10057);
and U10933 (N_10933,N_9749,N_9811);
and U10934 (N_10934,N_9765,N_10089);
xnor U10935 (N_10935,N_10406,N_9866);
xnor U10936 (N_10936,N_9953,N_10379);
nand U10937 (N_10937,N_9654,N_9967);
or U10938 (N_10938,N_10795,N_10380);
or U10939 (N_10939,N_10110,N_9888);
xnor U10940 (N_10940,N_10208,N_9781);
nand U10941 (N_10941,N_10785,N_9774);
nand U10942 (N_10942,N_10031,N_10517);
and U10943 (N_10943,N_10732,N_10601);
and U10944 (N_10944,N_10626,N_10319);
or U10945 (N_10945,N_10088,N_10773);
nor U10946 (N_10946,N_10327,N_9748);
or U10947 (N_10947,N_10726,N_10614);
nand U10948 (N_10948,N_9830,N_9958);
nor U10949 (N_10949,N_10616,N_10081);
nor U10950 (N_10950,N_9925,N_10157);
nand U10951 (N_10951,N_9908,N_9976);
nand U10952 (N_10952,N_10141,N_10426);
and U10953 (N_10953,N_10349,N_10781);
or U10954 (N_10954,N_10365,N_10664);
xor U10955 (N_10955,N_10528,N_9657);
nor U10956 (N_10956,N_10449,N_9833);
nand U10957 (N_10957,N_10111,N_10027);
nor U10958 (N_10958,N_9863,N_10092);
or U10959 (N_10959,N_10102,N_9904);
or U10960 (N_10960,N_10148,N_9732);
and U10961 (N_10961,N_10706,N_10524);
and U10962 (N_10962,N_10783,N_10329);
nor U10963 (N_10963,N_10372,N_10343);
or U10964 (N_10964,N_10122,N_9668);
and U10965 (N_10965,N_9899,N_10509);
nand U10966 (N_10966,N_10487,N_10633);
nor U10967 (N_10967,N_10321,N_10443);
and U10968 (N_10968,N_10001,N_10526);
nor U10969 (N_10969,N_10392,N_9844);
and U10970 (N_10970,N_10195,N_10130);
nand U10971 (N_10971,N_9993,N_9725);
and U10972 (N_10972,N_10046,N_10150);
nor U10973 (N_10973,N_9702,N_10015);
nor U10974 (N_10974,N_9723,N_10532);
xor U10975 (N_10975,N_9975,N_9798);
xnor U10976 (N_10976,N_10606,N_10452);
or U10977 (N_10977,N_10619,N_10104);
xnor U10978 (N_10978,N_10060,N_10258);
and U10979 (N_10979,N_10029,N_9937);
xor U10980 (N_10980,N_10236,N_10725);
or U10981 (N_10981,N_10542,N_10588);
nand U10982 (N_10982,N_10375,N_10127);
and U10983 (N_10983,N_10538,N_10337);
and U10984 (N_10984,N_10582,N_9640);
nand U10985 (N_10985,N_10273,N_9917);
and U10986 (N_10986,N_10086,N_9771);
or U10987 (N_10987,N_9791,N_10168);
xnor U10988 (N_10988,N_10737,N_10066);
nand U10989 (N_10989,N_9727,N_10652);
xnor U10990 (N_10990,N_10085,N_9848);
nand U10991 (N_10991,N_9875,N_9731);
xor U10992 (N_10992,N_10314,N_10461);
nand U10993 (N_10993,N_10410,N_9788);
and U10994 (N_10994,N_9701,N_10040);
xor U10995 (N_10995,N_10378,N_10533);
nor U10996 (N_10996,N_10585,N_10394);
nor U10997 (N_10997,N_10219,N_10573);
nor U10998 (N_10998,N_10432,N_10556);
nand U10999 (N_10999,N_10659,N_10070);
nor U11000 (N_11000,N_10301,N_10794);
nand U11001 (N_11001,N_10563,N_10268);
nand U11002 (N_11002,N_9743,N_9912);
nor U11003 (N_11003,N_10460,N_10317);
nand U11004 (N_11004,N_10395,N_9924);
xor U11005 (N_11005,N_10693,N_10736);
nand U11006 (N_11006,N_9944,N_10564);
xnor U11007 (N_11007,N_9672,N_10118);
nor U11008 (N_11008,N_10109,N_9796);
nand U11009 (N_11009,N_9855,N_10722);
nor U11010 (N_11010,N_10554,N_9627);
nor U11011 (N_11011,N_10051,N_10341);
nand U11012 (N_11012,N_9878,N_10421);
and U11013 (N_11013,N_9831,N_10469);
nand U11014 (N_11014,N_10160,N_9927);
xnor U11015 (N_11015,N_9928,N_10735);
or U11016 (N_11016,N_10205,N_9845);
nor U11017 (N_11017,N_10625,N_10763);
nand U11018 (N_11018,N_10182,N_10045);
or U11019 (N_11019,N_10766,N_10177);
nand U11020 (N_11020,N_10694,N_10069);
nand U11021 (N_11021,N_9766,N_9837);
nand U11022 (N_11022,N_9820,N_10142);
xnor U11023 (N_11023,N_9600,N_9733);
and U11024 (N_11024,N_9910,N_10171);
and U11025 (N_11025,N_10361,N_9883);
nor U11026 (N_11026,N_10280,N_10245);
nor U11027 (N_11027,N_10383,N_10540);
or U11028 (N_11028,N_10364,N_10627);
and U11029 (N_11029,N_10144,N_10209);
and U11030 (N_11030,N_9979,N_10302);
xnor U11031 (N_11031,N_10486,N_10484);
nand U11032 (N_11032,N_9793,N_10568);
nand U11033 (N_11033,N_10511,N_10525);
or U11034 (N_11034,N_9643,N_9919);
or U11035 (N_11035,N_9834,N_10370);
nand U11036 (N_11036,N_9641,N_10611);
nand U11037 (N_11037,N_9846,N_10545);
xnor U11038 (N_11038,N_9662,N_9947);
or U11039 (N_11039,N_10011,N_10464);
xor U11040 (N_11040,N_9859,N_10153);
nand U11041 (N_11041,N_10399,N_10711);
and U11042 (N_11042,N_10166,N_10077);
or U11043 (N_11043,N_10255,N_9786);
xnor U11044 (N_11044,N_10641,N_10225);
nor U11045 (N_11045,N_10676,N_10681);
or U11046 (N_11046,N_10458,N_10550);
nor U11047 (N_11047,N_10718,N_10459);
nor U11048 (N_11048,N_9735,N_9823);
nor U11049 (N_11049,N_10035,N_10529);
xor U11050 (N_11050,N_10579,N_10183);
nor U11051 (N_11051,N_9601,N_10586);
nand U11052 (N_11052,N_10105,N_10326);
or U11053 (N_11053,N_10497,N_10214);
or U11054 (N_11054,N_9933,N_9614);
xnor U11055 (N_11055,N_10714,N_10169);
or U11056 (N_11056,N_10340,N_10124);
or U11057 (N_11057,N_10203,N_10727);
xnor U11058 (N_11058,N_10425,N_9708);
or U11059 (N_11059,N_9852,N_10466);
xor U11060 (N_11060,N_10408,N_10325);
or U11061 (N_11061,N_10440,N_9780);
nor U11062 (N_11062,N_9902,N_10493);
nand U11063 (N_11063,N_10173,N_10251);
or U11064 (N_11064,N_10618,N_10648);
xnor U11065 (N_11065,N_9843,N_10320);
and U11066 (N_11066,N_10403,N_9923);
nor U11067 (N_11067,N_10385,N_10293);
or U11068 (N_11068,N_10310,N_10583);
nor U11069 (N_11069,N_9754,N_9850);
nand U11070 (N_11070,N_9968,N_9650);
nor U11071 (N_11071,N_10377,N_9634);
xor U11072 (N_11072,N_10054,N_10353);
nor U11073 (N_11073,N_9801,N_9639);
xnor U11074 (N_11074,N_10782,N_10311);
nor U11075 (N_11075,N_10072,N_10696);
xnor U11076 (N_11076,N_9985,N_10044);
or U11077 (N_11077,N_10716,N_10510);
nand U11078 (N_11078,N_10592,N_10296);
nand U11079 (N_11079,N_10303,N_10322);
and U11080 (N_11080,N_10309,N_9689);
nand U11081 (N_11081,N_9959,N_9840);
or U11082 (N_11082,N_10093,N_9861);
and U11083 (N_11083,N_9785,N_9994);
nand U11084 (N_11084,N_9607,N_10522);
or U11085 (N_11085,N_10764,N_10445);
and U11086 (N_11086,N_9741,N_10348);
and U11087 (N_11087,N_9938,N_9721);
nand U11088 (N_11088,N_9856,N_10413);
and U11089 (N_11089,N_9703,N_9945);
xnor U11090 (N_11090,N_10138,N_9799);
nor U11091 (N_11091,N_9776,N_10715);
nand U11092 (N_11092,N_9778,N_9821);
nor U11093 (N_11093,N_9822,N_10521);
nand U11094 (N_11094,N_10024,N_9827);
or U11095 (N_11095,N_10437,N_10751);
nand U11096 (N_11096,N_10775,N_9632);
nand U11097 (N_11097,N_10721,N_10315);
nor U11098 (N_11098,N_10270,N_10246);
nor U11099 (N_11099,N_9954,N_9982);
nand U11100 (N_11100,N_10106,N_10412);
nor U11101 (N_11101,N_10701,N_9870);
and U11102 (N_11102,N_10184,N_10247);
or U11103 (N_11103,N_10689,N_10595);
or U11104 (N_11104,N_10107,N_9736);
and U11105 (N_11105,N_10501,N_10791);
nor U11106 (N_11106,N_10778,N_9624);
and U11107 (N_11107,N_10477,N_9873);
xor U11108 (N_11108,N_10241,N_9759);
xor U11109 (N_11109,N_10212,N_9810);
or U11110 (N_11110,N_10792,N_10544);
and U11111 (N_11111,N_10025,N_10470);
or U11112 (N_11112,N_10265,N_10129);
nor U11113 (N_11113,N_10670,N_10180);
nand U11114 (N_11114,N_10613,N_10261);
or U11115 (N_11115,N_10640,N_9828);
and U11116 (N_11116,N_10790,N_9842);
nor U11117 (N_11117,N_10012,N_10453);
xnor U11118 (N_11118,N_9694,N_10023);
nand U11119 (N_11119,N_10053,N_10767);
nor U11120 (N_11120,N_10669,N_10589);
nand U11121 (N_11121,N_10546,N_10488);
or U11122 (N_11122,N_10328,N_10765);
nand U11123 (N_11123,N_10264,N_10411);
and U11124 (N_11124,N_10249,N_10771);
nand U11125 (N_11125,N_9999,N_10179);
or U11126 (N_11126,N_9700,N_9760);
nor U11127 (N_11127,N_9935,N_10755);
and U11128 (N_11128,N_10673,N_9679);
and U11129 (N_11129,N_9877,N_9683);
nand U11130 (N_11130,N_10788,N_10577);
nor U11131 (N_11131,N_10125,N_10620);
xor U11132 (N_11132,N_9802,N_10728);
xor U11133 (N_11133,N_10427,N_9966);
nand U11134 (N_11134,N_10285,N_10351);
or U11135 (N_11135,N_10646,N_10446);
nor U11136 (N_11136,N_10238,N_10114);
or U11137 (N_11137,N_10041,N_9674);
nand U11138 (N_11138,N_10717,N_10313);
and U11139 (N_11139,N_10281,N_10176);
nor U11140 (N_11140,N_10748,N_10004);
nand U11141 (N_11141,N_10161,N_9667);
xor U11142 (N_11142,N_10553,N_9815);
and U11143 (N_11143,N_10743,N_9671);
or U11144 (N_11144,N_10123,N_10473);
xnor U11145 (N_11145,N_10433,N_9898);
or U11146 (N_11146,N_9901,N_10503);
and U11147 (N_11147,N_10389,N_9926);
nand U11148 (N_11148,N_9818,N_10239);
nand U11149 (N_11149,N_10132,N_10753);
and U11150 (N_11150,N_9960,N_10476);
or U11151 (N_11151,N_9957,N_9986);
and U11152 (N_11152,N_9768,N_10140);
nor U11153 (N_11153,N_9779,N_9677);
xnor U11154 (N_11154,N_9619,N_10215);
nor U11155 (N_11155,N_9744,N_10645);
and U11156 (N_11156,N_9660,N_9868);
nand U11157 (N_11157,N_10158,N_10441);
nor U11158 (N_11158,N_9906,N_10286);
nand U11159 (N_11159,N_10087,N_9948);
or U11160 (N_11160,N_10096,N_9871);
xnor U11161 (N_11161,N_10658,N_9615);
and U11162 (N_11162,N_10282,N_10490);
and U11163 (N_11163,N_9698,N_9773);
and U11164 (N_11164,N_10164,N_9685);
xnor U11165 (N_11165,N_9804,N_10211);
xnor U11166 (N_11166,N_10222,N_10796);
nand U11167 (N_11167,N_10287,N_10608);
nor U11168 (N_11168,N_10260,N_10667);
nand U11169 (N_11169,N_9992,N_9836);
and U11170 (N_11170,N_10038,N_10451);
xnor U11171 (N_11171,N_10189,N_10428);
nand U11172 (N_11172,N_10500,N_10201);
xnor U11173 (N_11173,N_10635,N_10306);
nand U11174 (N_11174,N_10536,N_10274);
and U11175 (N_11175,N_10095,N_10139);
or U11176 (N_11176,N_10598,N_10702);
nand U11177 (N_11177,N_10777,N_10636);
or U11178 (N_11178,N_10099,N_9795);
nand U11179 (N_11179,N_9981,N_10710);
or U11180 (N_11180,N_9980,N_10548);
and U11181 (N_11181,N_10624,N_9729);
nor U11182 (N_11182,N_10762,N_10185);
nor U11183 (N_11183,N_9991,N_10165);
nand U11184 (N_11184,N_10021,N_10494);
nor U11185 (N_11185,N_10218,N_10295);
xor U11186 (N_11186,N_10686,N_10055);
xnor U11187 (N_11187,N_10400,N_10651);
and U11188 (N_11188,N_10468,N_9648);
and U11189 (N_11189,N_9750,N_10229);
nor U11190 (N_11190,N_9934,N_10240);
nand U11191 (N_11191,N_9763,N_9894);
nand U11192 (N_11192,N_10518,N_9726);
and U11193 (N_11193,N_10009,N_10318);
and U11194 (N_11194,N_9887,N_9604);
nand U11195 (N_11195,N_10688,N_10776);
xor U11196 (N_11196,N_9995,N_10312);
xnor U11197 (N_11197,N_10584,N_9895);
nor U11198 (N_11198,N_10729,N_10008);
or U11199 (N_11199,N_10335,N_10277);
nor U11200 (N_11200,N_9867,N_9936);
nor U11201 (N_11201,N_10294,N_9838);
nor U11202 (N_11202,N_10705,N_10071);
xor U11203 (N_11203,N_9950,N_10100);
nand U11204 (N_11204,N_10439,N_10194);
nand U11205 (N_11205,N_10442,N_9655);
xor U11206 (N_11206,N_10690,N_10391);
or U11207 (N_11207,N_10278,N_9636);
xnor U11208 (N_11208,N_9916,N_10067);
nor U11209 (N_11209,N_10541,N_9897);
or U11210 (N_11210,N_10298,N_9949);
nor U11211 (N_11211,N_9816,N_10639);
and U11212 (N_11212,N_9772,N_10134);
nor U11213 (N_11213,N_9739,N_9742);
nor U11214 (N_11214,N_9913,N_9849);
and U11215 (N_11215,N_10547,N_10502);
xnor U11216 (N_11216,N_10362,N_10297);
or U11217 (N_11217,N_9713,N_10687);
nand U11218 (N_11218,N_9783,N_9893);
nor U11219 (N_11219,N_9653,N_10600);
and U11220 (N_11220,N_10232,N_10275);
nor U11221 (N_11221,N_9656,N_10233);
xor U11222 (N_11222,N_10098,N_9764);
and U11223 (N_11223,N_10366,N_9996);
xor U11224 (N_11224,N_9829,N_10621);
and U11225 (N_11225,N_10064,N_10569);
nand U11226 (N_11226,N_10398,N_9941);
nor U11227 (N_11227,N_10506,N_9720);
nand U11228 (N_11228,N_10156,N_9792);
and U11229 (N_11229,N_9824,N_9987);
xor U11230 (N_11230,N_9617,N_10036);
xor U11231 (N_11231,N_10416,N_9605);
xor U11232 (N_11232,N_10709,N_10543);
nor U11233 (N_11233,N_10248,N_10323);
nand U11234 (N_11234,N_9647,N_10779);
and U11235 (N_11235,N_9961,N_10507);
or U11236 (N_11236,N_10345,N_10733);
and U11237 (N_11237,N_10558,N_10097);
and U11238 (N_11238,N_9646,N_10703);
or U11239 (N_11239,N_10037,N_9681);
or U11240 (N_11240,N_10022,N_10074);
or U11241 (N_11241,N_9955,N_9746);
and U11242 (N_11242,N_10630,N_10677);
and U11243 (N_11243,N_10750,N_10780);
nand U11244 (N_11244,N_10523,N_10216);
or U11245 (N_11245,N_9970,N_10695);
xor U11246 (N_11246,N_9809,N_9730);
and U11247 (N_11247,N_10758,N_10657);
nand U11248 (N_11248,N_10549,N_10381);
nor U11249 (N_11249,N_10073,N_9769);
nor U11250 (N_11250,N_9712,N_10256);
and U11251 (N_11251,N_10336,N_10575);
and U11252 (N_11252,N_10571,N_10350);
nor U11253 (N_11253,N_9612,N_9762);
nor U11254 (N_11254,N_9631,N_9649);
nor U11255 (N_11255,N_10254,N_9909);
and U11256 (N_11256,N_10133,N_10369);
and U11257 (N_11257,N_10010,N_10076);
nand U11258 (N_11258,N_9808,N_9984);
and U11259 (N_11259,N_10288,N_10671);
nor U11260 (N_11260,N_10078,N_10697);
xnor U11261 (N_11261,N_10359,N_10407);
nand U11262 (N_11262,N_10145,N_10082);
or U11263 (N_11263,N_10797,N_10271);
and U11264 (N_11264,N_10570,N_10146);
nand U11265 (N_11265,N_10450,N_10404);
xor U11266 (N_11266,N_9942,N_10065);
or U11267 (N_11267,N_10415,N_10135);
xor U11268 (N_11268,N_10200,N_10242);
and U11269 (N_11269,N_10244,N_10162);
xnor U11270 (N_11270,N_9628,N_10457);
nor U11271 (N_11271,N_10786,N_10596);
nor U11272 (N_11272,N_9711,N_9758);
or U11273 (N_11273,N_10155,N_9965);
nand U11274 (N_11274,N_10784,N_9977);
xnor U11275 (N_11275,N_9706,N_9767);
or U11276 (N_11276,N_9940,N_9869);
and U11277 (N_11277,N_10535,N_10143);
nor U11278 (N_11278,N_9998,N_9658);
nor U11279 (N_11279,N_10745,N_9688);
nor U11280 (N_11280,N_9673,N_10202);
or U11281 (N_11281,N_9858,N_10384);
and U11282 (N_11282,N_10252,N_10489);
and U11283 (N_11283,N_10590,N_9812);
xor U11284 (N_11284,N_9752,N_9753);
nand U11285 (N_11285,N_10393,N_9629);
xnor U11286 (N_11286,N_9864,N_9939);
and U11287 (N_11287,N_9745,N_9770);
xor U11288 (N_11288,N_10438,N_10367);
and U11289 (N_11289,N_10471,N_10386);
nand U11290 (N_11290,N_9932,N_9989);
nand U11291 (N_11291,N_10154,N_9645);
nor U11292 (N_11292,N_10514,N_9943);
nand U11293 (N_11293,N_9755,N_10079);
nand U11294 (N_11294,N_10623,N_10363);
nor U11295 (N_11295,N_10338,N_9814);
xnor U11296 (N_11296,N_10220,N_10576);
nor U11297 (N_11297,N_9990,N_10003);
nor U11298 (N_11298,N_9608,N_10653);
and U11299 (N_11299,N_9661,N_10355);
xnor U11300 (N_11300,N_9606,N_10479);
xnor U11301 (N_11301,N_10560,N_10191);
nand U11302 (N_11302,N_10346,N_10388);
and U11303 (N_11303,N_10108,N_10512);
or U11304 (N_11304,N_9666,N_10152);
or U11305 (N_11305,N_10769,N_10159);
and U11306 (N_11306,N_9714,N_10463);
or U11307 (N_11307,N_9782,N_10094);
xor U11308 (N_11308,N_9630,N_10028);
nor U11309 (N_11309,N_10591,N_10198);
or U11310 (N_11310,N_9664,N_9751);
or U11311 (N_11311,N_10480,N_10213);
xnor U11312 (N_11312,N_10622,N_10603);
or U11313 (N_11313,N_10741,N_10117);
and U11314 (N_11314,N_10390,N_10174);
nand U11315 (N_11315,N_9839,N_9854);
nand U11316 (N_11316,N_10516,N_9963);
or U11317 (N_11317,N_10119,N_10324);
and U11318 (N_11318,N_10204,N_9969);
nor U11319 (N_11319,N_10713,N_10332);
and U11320 (N_11320,N_10629,N_10186);
nand U11321 (N_11321,N_10354,N_10172);
and U11322 (N_11322,N_10685,N_10552);
xor U11323 (N_11323,N_10707,N_10691);
nor U11324 (N_11324,N_10539,N_9709);
nand U11325 (N_11325,N_10014,N_10344);
xnor U11326 (N_11326,N_10083,N_10615);
or U11327 (N_11327,N_10136,N_10103);
and U11328 (N_11328,N_10188,N_10116);
xor U11329 (N_11329,N_10192,N_10207);
or U11330 (N_11330,N_9851,N_10090);
xnor U11331 (N_11331,N_10436,N_10789);
xor U11332 (N_11332,N_10562,N_9973);
nand U11333 (N_11333,N_10580,N_10757);
or U11334 (N_11334,N_10418,N_10050);
or U11335 (N_11335,N_10655,N_10665);
nor U11336 (N_11336,N_9625,N_10495);
and U11337 (N_11337,N_10483,N_10243);
nand U11338 (N_11338,N_9697,N_10005);
xnor U11339 (N_11339,N_10774,N_10291);
xor U11340 (N_11340,N_9885,N_9757);
nand U11341 (N_11341,N_10290,N_10056);
xnor U11342 (N_11342,N_10197,N_10684);
and U11343 (N_11343,N_10020,N_9696);
xor U11344 (N_11344,N_9800,N_9951);
or U11345 (N_11345,N_10308,N_10034);
or U11346 (N_11346,N_9737,N_10017);
xor U11347 (N_11347,N_9881,N_9618);
nand U11348 (N_11348,N_9900,N_10115);
nand U11349 (N_11349,N_10605,N_10007);
xor U11350 (N_11350,N_10131,N_10587);
or U11351 (N_11351,N_10049,N_10643);
and U11352 (N_11352,N_10080,N_10059);
nand U11353 (N_11353,N_10063,N_9922);
nand U11354 (N_11354,N_10666,N_10597);
nand U11355 (N_11355,N_10572,N_10448);
nor U11356 (N_11356,N_10368,N_10113);
nor U11357 (N_11357,N_9659,N_9931);
nor U11358 (N_11358,N_10237,N_9663);
nand U11359 (N_11359,N_10163,N_10002);
nand U11360 (N_11360,N_10749,N_10360);
or U11361 (N_11361,N_10531,N_10061);
nand U11362 (N_11362,N_10747,N_10279);
xnor U11363 (N_11363,N_9915,N_10740);
nor U11364 (N_11364,N_10678,N_9794);
and U11365 (N_11365,N_9930,N_10235);
nor U11366 (N_11366,N_9718,N_10638);
xnor U11367 (N_11367,N_10680,N_9797);
nor U11368 (N_11368,N_10768,N_10508);
nand U11369 (N_11369,N_10396,N_10292);
and U11370 (N_11370,N_10607,N_9807);
or U11371 (N_11371,N_10266,N_9691);
xnor U11372 (N_11372,N_10496,N_9603);
xor U11373 (N_11373,N_10752,N_10187);
nor U11374 (N_11374,N_9971,N_10262);
nor U11375 (N_11375,N_10799,N_10730);
xor U11376 (N_11376,N_10602,N_9756);
or U11377 (N_11377,N_10206,N_10342);
xnor U11378 (N_11378,N_10259,N_10000);
nand U11379 (N_11379,N_10504,N_10167);
nand U11380 (N_11380,N_9865,N_9717);
or U11381 (N_11381,N_9803,N_10223);
or U11382 (N_11382,N_10699,N_10013);
nor U11383 (N_11383,N_10231,N_10474);
nand U11384 (N_11384,N_10196,N_9747);
nor U11385 (N_11385,N_10101,N_10330);
or U11386 (N_11386,N_9784,N_10217);
or U11387 (N_11387,N_9693,N_9710);
and U11388 (N_11388,N_10226,N_10420);
nand U11389 (N_11389,N_10724,N_10742);
xnor U11390 (N_11390,N_10043,N_10578);
nand U11391 (N_11391,N_10537,N_9952);
nand U11392 (N_11392,N_10679,N_10698);
nor U11393 (N_11393,N_9789,N_9806);
nand U11394 (N_11394,N_9670,N_10478);
nor U11395 (N_11395,N_9962,N_10062);
or U11396 (N_11396,N_10700,N_10228);
xor U11397 (N_11397,N_9874,N_10756);
nand U11398 (N_11398,N_9678,N_9644);
or U11399 (N_11399,N_10305,N_10772);
nor U11400 (N_11400,N_10245,N_10232);
or U11401 (N_11401,N_10574,N_10660);
and U11402 (N_11402,N_10423,N_10684);
or U11403 (N_11403,N_10461,N_9867);
or U11404 (N_11404,N_10381,N_10640);
or U11405 (N_11405,N_10413,N_9859);
nor U11406 (N_11406,N_10090,N_9949);
or U11407 (N_11407,N_10520,N_10795);
or U11408 (N_11408,N_9760,N_10004);
and U11409 (N_11409,N_10594,N_9748);
nand U11410 (N_11410,N_10309,N_9790);
and U11411 (N_11411,N_10553,N_10301);
or U11412 (N_11412,N_10707,N_10371);
nand U11413 (N_11413,N_10777,N_9927);
xor U11414 (N_11414,N_10627,N_10653);
xnor U11415 (N_11415,N_10784,N_10251);
or U11416 (N_11416,N_9903,N_9983);
and U11417 (N_11417,N_10684,N_10331);
and U11418 (N_11418,N_10280,N_10073);
nand U11419 (N_11419,N_10666,N_9625);
and U11420 (N_11420,N_10451,N_9655);
nor U11421 (N_11421,N_9917,N_10328);
xnor U11422 (N_11422,N_10068,N_9842);
and U11423 (N_11423,N_10764,N_10444);
nand U11424 (N_11424,N_9669,N_10257);
or U11425 (N_11425,N_10120,N_10397);
xnor U11426 (N_11426,N_9725,N_10577);
nand U11427 (N_11427,N_10751,N_9658);
and U11428 (N_11428,N_9974,N_9685);
and U11429 (N_11429,N_9819,N_9647);
or U11430 (N_11430,N_10534,N_10044);
and U11431 (N_11431,N_10770,N_10413);
nor U11432 (N_11432,N_10506,N_10326);
xnor U11433 (N_11433,N_9775,N_10778);
nor U11434 (N_11434,N_10341,N_9601);
xnor U11435 (N_11435,N_10560,N_10626);
nand U11436 (N_11436,N_9937,N_10031);
nor U11437 (N_11437,N_9826,N_10526);
nor U11438 (N_11438,N_10662,N_10789);
xor U11439 (N_11439,N_9793,N_9952);
nand U11440 (N_11440,N_10061,N_9982);
and U11441 (N_11441,N_9950,N_10025);
and U11442 (N_11442,N_10086,N_9689);
xor U11443 (N_11443,N_9961,N_10436);
xnor U11444 (N_11444,N_9901,N_9915);
xnor U11445 (N_11445,N_10422,N_9788);
and U11446 (N_11446,N_10229,N_10175);
xor U11447 (N_11447,N_10517,N_9990);
nand U11448 (N_11448,N_10574,N_10711);
nand U11449 (N_11449,N_10385,N_10730);
nand U11450 (N_11450,N_10335,N_9749);
and U11451 (N_11451,N_9922,N_10476);
nand U11452 (N_11452,N_10097,N_10155);
nand U11453 (N_11453,N_10711,N_10635);
or U11454 (N_11454,N_10404,N_10368);
xor U11455 (N_11455,N_10663,N_10209);
or U11456 (N_11456,N_9722,N_10471);
nor U11457 (N_11457,N_10467,N_9759);
nand U11458 (N_11458,N_10229,N_10273);
nor U11459 (N_11459,N_9742,N_10773);
and U11460 (N_11460,N_9818,N_10559);
xor U11461 (N_11461,N_10726,N_9622);
nor U11462 (N_11462,N_10606,N_10721);
nand U11463 (N_11463,N_10328,N_9772);
nand U11464 (N_11464,N_10412,N_10411);
xnor U11465 (N_11465,N_9772,N_10069);
xor U11466 (N_11466,N_10584,N_10654);
or U11467 (N_11467,N_9986,N_10401);
or U11468 (N_11468,N_9897,N_10245);
nand U11469 (N_11469,N_10598,N_10405);
xnor U11470 (N_11470,N_10435,N_10051);
xnor U11471 (N_11471,N_10594,N_10287);
nor U11472 (N_11472,N_10280,N_9784);
or U11473 (N_11473,N_9647,N_10003);
or U11474 (N_11474,N_9900,N_10225);
and U11475 (N_11475,N_9611,N_9655);
nand U11476 (N_11476,N_9901,N_10636);
xor U11477 (N_11477,N_10083,N_10378);
or U11478 (N_11478,N_10095,N_10550);
xnor U11479 (N_11479,N_10313,N_10347);
and U11480 (N_11480,N_9828,N_10442);
nand U11481 (N_11481,N_10710,N_10500);
and U11482 (N_11482,N_10482,N_9838);
nor U11483 (N_11483,N_10727,N_10670);
nand U11484 (N_11484,N_10338,N_10266);
nor U11485 (N_11485,N_9767,N_9690);
and U11486 (N_11486,N_10013,N_10190);
nand U11487 (N_11487,N_10463,N_10186);
xor U11488 (N_11488,N_10641,N_10254);
xor U11489 (N_11489,N_10436,N_10787);
and U11490 (N_11490,N_10039,N_10011);
nand U11491 (N_11491,N_10435,N_9864);
nor U11492 (N_11492,N_10446,N_9803);
and U11493 (N_11493,N_10037,N_10411);
and U11494 (N_11494,N_9965,N_9879);
or U11495 (N_11495,N_10145,N_10771);
and U11496 (N_11496,N_10409,N_10477);
nand U11497 (N_11497,N_10431,N_9961);
or U11498 (N_11498,N_10698,N_10704);
or U11499 (N_11499,N_9853,N_9867);
or U11500 (N_11500,N_10488,N_9801);
and U11501 (N_11501,N_9990,N_10303);
nand U11502 (N_11502,N_9604,N_10131);
xnor U11503 (N_11503,N_10732,N_9635);
nor U11504 (N_11504,N_10249,N_10785);
nand U11505 (N_11505,N_10789,N_9808);
and U11506 (N_11506,N_10478,N_10181);
or U11507 (N_11507,N_10175,N_10293);
xor U11508 (N_11508,N_10671,N_10238);
or U11509 (N_11509,N_10055,N_10795);
nor U11510 (N_11510,N_10151,N_9874);
and U11511 (N_11511,N_9966,N_9804);
and U11512 (N_11512,N_10246,N_9823);
or U11513 (N_11513,N_10167,N_10433);
xor U11514 (N_11514,N_10261,N_9986);
nand U11515 (N_11515,N_10154,N_9896);
and U11516 (N_11516,N_9892,N_9877);
or U11517 (N_11517,N_9819,N_9820);
nand U11518 (N_11518,N_10269,N_10633);
and U11519 (N_11519,N_9877,N_9747);
xnor U11520 (N_11520,N_10194,N_10442);
or U11521 (N_11521,N_9753,N_10488);
or U11522 (N_11522,N_10378,N_10560);
and U11523 (N_11523,N_9715,N_10288);
nor U11524 (N_11524,N_9884,N_10190);
nand U11525 (N_11525,N_9623,N_10558);
xnor U11526 (N_11526,N_10155,N_10734);
and U11527 (N_11527,N_9781,N_10155);
nor U11528 (N_11528,N_9640,N_10768);
nor U11529 (N_11529,N_9715,N_9610);
and U11530 (N_11530,N_10633,N_9990);
nor U11531 (N_11531,N_10108,N_10416);
or U11532 (N_11532,N_10401,N_9777);
and U11533 (N_11533,N_10550,N_10396);
nor U11534 (N_11534,N_9936,N_10647);
and U11535 (N_11535,N_10749,N_10032);
or U11536 (N_11536,N_10144,N_10601);
xor U11537 (N_11537,N_10534,N_10463);
nor U11538 (N_11538,N_10226,N_10796);
and U11539 (N_11539,N_10116,N_10767);
and U11540 (N_11540,N_10493,N_9710);
nand U11541 (N_11541,N_10600,N_10033);
nor U11542 (N_11542,N_10792,N_9606);
xor U11543 (N_11543,N_10534,N_10336);
or U11544 (N_11544,N_10677,N_9905);
nand U11545 (N_11545,N_10173,N_10697);
nand U11546 (N_11546,N_10105,N_9924);
xor U11547 (N_11547,N_10060,N_10657);
nand U11548 (N_11548,N_9644,N_9663);
or U11549 (N_11549,N_10316,N_9820);
nor U11550 (N_11550,N_10337,N_10531);
nand U11551 (N_11551,N_10171,N_10510);
or U11552 (N_11552,N_9691,N_10434);
nand U11553 (N_11553,N_9810,N_9879);
nand U11554 (N_11554,N_9622,N_10081);
nor U11555 (N_11555,N_9965,N_10764);
or U11556 (N_11556,N_10109,N_10660);
xnor U11557 (N_11557,N_10616,N_9822);
nand U11558 (N_11558,N_10089,N_10200);
nand U11559 (N_11559,N_10548,N_10567);
nor U11560 (N_11560,N_10611,N_10529);
or U11561 (N_11561,N_10774,N_10425);
xor U11562 (N_11562,N_9996,N_10680);
xor U11563 (N_11563,N_10178,N_10713);
nand U11564 (N_11564,N_9850,N_10064);
nand U11565 (N_11565,N_10584,N_10389);
or U11566 (N_11566,N_10080,N_10643);
nor U11567 (N_11567,N_9728,N_10214);
or U11568 (N_11568,N_10166,N_10410);
nor U11569 (N_11569,N_9928,N_10524);
or U11570 (N_11570,N_9992,N_10036);
or U11571 (N_11571,N_10186,N_10167);
or U11572 (N_11572,N_10200,N_10307);
and U11573 (N_11573,N_10544,N_9856);
nor U11574 (N_11574,N_10450,N_10428);
nand U11575 (N_11575,N_9905,N_10077);
and U11576 (N_11576,N_10325,N_10585);
xnor U11577 (N_11577,N_9957,N_10277);
nor U11578 (N_11578,N_9763,N_10540);
or U11579 (N_11579,N_9847,N_10583);
xnor U11580 (N_11580,N_9742,N_10464);
or U11581 (N_11581,N_10586,N_9976);
nor U11582 (N_11582,N_9711,N_9956);
xnor U11583 (N_11583,N_10666,N_10145);
and U11584 (N_11584,N_10769,N_9914);
nor U11585 (N_11585,N_10336,N_10763);
xnor U11586 (N_11586,N_9663,N_9877);
or U11587 (N_11587,N_10283,N_9615);
nand U11588 (N_11588,N_10457,N_10794);
xor U11589 (N_11589,N_10248,N_10690);
nor U11590 (N_11590,N_10616,N_9935);
xor U11591 (N_11591,N_10664,N_10766);
nand U11592 (N_11592,N_10782,N_10738);
or U11593 (N_11593,N_10002,N_10375);
nor U11594 (N_11594,N_9854,N_10491);
nor U11595 (N_11595,N_10176,N_10755);
nor U11596 (N_11596,N_10310,N_10702);
nor U11597 (N_11597,N_9948,N_10157);
or U11598 (N_11598,N_9722,N_9663);
nor U11599 (N_11599,N_9891,N_10365);
nor U11600 (N_11600,N_10447,N_9647);
nor U11601 (N_11601,N_9751,N_9606);
nor U11602 (N_11602,N_9762,N_9931);
or U11603 (N_11603,N_9823,N_9801);
xor U11604 (N_11604,N_10698,N_10759);
nor U11605 (N_11605,N_10433,N_10427);
xnor U11606 (N_11606,N_9890,N_10072);
nand U11607 (N_11607,N_10699,N_9900);
xnor U11608 (N_11608,N_10184,N_10420);
xor U11609 (N_11609,N_10734,N_10670);
xnor U11610 (N_11610,N_10023,N_10205);
nand U11611 (N_11611,N_9810,N_9975);
or U11612 (N_11612,N_10717,N_10111);
nand U11613 (N_11613,N_9940,N_9742);
and U11614 (N_11614,N_9762,N_10473);
xor U11615 (N_11615,N_10553,N_10438);
and U11616 (N_11616,N_9815,N_10070);
nand U11617 (N_11617,N_10583,N_9973);
nor U11618 (N_11618,N_10612,N_9663);
xnor U11619 (N_11619,N_9895,N_10773);
or U11620 (N_11620,N_10220,N_10423);
nor U11621 (N_11621,N_9748,N_10223);
nor U11622 (N_11622,N_10528,N_10030);
nand U11623 (N_11623,N_9853,N_10316);
or U11624 (N_11624,N_9921,N_9956);
and U11625 (N_11625,N_10045,N_10590);
and U11626 (N_11626,N_10680,N_10506);
and U11627 (N_11627,N_10235,N_9781);
xnor U11628 (N_11628,N_9844,N_10576);
or U11629 (N_11629,N_10048,N_9705);
nand U11630 (N_11630,N_9906,N_10104);
or U11631 (N_11631,N_9951,N_10520);
nor U11632 (N_11632,N_10272,N_9775);
and U11633 (N_11633,N_10205,N_10210);
nor U11634 (N_11634,N_9856,N_10194);
or U11635 (N_11635,N_9816,N_10613);
xor U11636 (N_11636,N_10210,N_10408);
nand U11637 (N_11637,N_10484,N_10229);
xnor U11638 (N_11638,N_9896,N_10078);
or U11639 (N_11639,N_10063,N_10729);
nand U11640 (N_11640,N_10280,N_10020);
and U11641 (N_11641,N_10621,N_10042);
and U11642 (N_11642,N_10769,N_10248);
xnor U11643 (N_11643,N_10665,N_10451);
xnor U11644 (N_11644,N_10038,N_9683);
or U11645 (N_11645,N_10127,N_10452);
or U11646 (N_11646,N_9906,N_10692);
nand U11647 (N_11647,N_10438,N_10798);
or U11648 (N_11648,N_10104,N_10293);
and U11649 (N_11649,N_9928,N_10797);
xor U11650 (N_11650,N_9842,N_10730);
nand U11651 (N_11651,N_10501,N_9604);
and U11652 (N_11652,N_10034,N_9696);
xor U11653 (N_11653,N_10132,N_9809);
and U11654 (N_11654,N_9632,N_10150);
nand U11655 (N_11655,N_10758,N_9929);
xor U11656 (N_11656,N_9793,N_10794);
or U11657 (N_11657,N_10411,N_10381);
nand U11658 (N_11658,N_9865,N_10190);
nor U11659 (N_11659,N_9677,N_10697);
and U11660 (N_11660,N_10056,N_10558);
and U11661 (N_11661,N_10481,N_10718);
nand U11662 (N_11662,N_10161,N_10695);
and U11663 (N_11663,N_10290,N_10687);
or U11664 (N_11664,N_10221,N_10420);
xnor U11665 (N_11665,N_10111,N_9884);
xnor U11666 (N_11666,N_10409,N_9770);
xor U11667 (N_11667,N_10294,N_9666);
and U11668 (N_11668,N_10306,N_10136);
nand U11669 (N_11669,N_9914,N_9737);
and U11670 (N_11670,N_9764,N_10000);
xnor U11671 (N_11671,N_10667,N_10735);
nor U11672 (N_11672,N_9997,N_9989);
xnor U11673 (N_11673,N_10276,N_10204);
or U11674 (N_11674,N_9707,N_10577);
and U11675 (N_11675,N_10768,N_9891);
nor U11676 (N_11676,N_9892,N_9779);
and U11677 (N_11677,N_9640,N_9984);
nor U11678 (N_11678,N_9805,N_10502);
and U11679 (N_11679,N_9982,N_10555);
or U11680 (N_11680,N_10164,N_10157);
xor U11681 (N_11681,N_9656,N_10670);
nor U11682 (N_11682,N_10421,N_10488);
and U11683 (N_11683,N_9867,N_10119);
or U11684 (N_11684,N_10127,N_9681);
nand U11685 (N_11685,N_10696,N_10091);
and U11686 (N_11686,N_9818,N_10179);
nor U11687 (N_11687,N_9963,N_10727);
and U11688 (N_11688,N_10358,N_10568);
or U11689 (N_11689,N_10472,N_9842);
xor U11690 (N_11690,N_9623,N_9923);
nand U11691 (N_11691,N_10321,N_9915);
or U11692 (N_11692,N_10238,N_10477);
and U11693 (N_11693,N_10509,N_10298);
nor U11694 (N_11694,N_10615,N_9710);
and U11695 (N_11695,N_10626,N_9847);
and U11696 (N_11696,N_10430,N_10452);
nand U11697 (N_11697,N_9853,N_9848);
and U11698 (N_11698,N_10316,N_10525);
nand U11699 (N_11699,N_9711,N_10210);
and U11700 (N_11700,N_10092,N_9786);
or U11701 (N_11701,N_10379,N_10769);
or U11702 (N_11702,N_10557,N_9947);
nand U11703 (N_11703,N_10537,N_10387);
nor U11704 (N_11704,N_9727,N_10650);
nand U11705 (N_11705,N_10435,N_9823);
nor U11706 (N_11706,N_10108,N_10473);
and U11707 (N_11707,N_9792,N_10458);
and U11708 (N_11708,N_10644,N_10764);
nor U11709 (N_11709,N_10539,N_10550);
nor U11710 (N_11710,N_10523,N_10477);
nand U11711 (N_11711,N_10185,N_10590);
nor U11712 (N_11712,N_9965,N_10698);
nand U11713 (N_11713,N_10403,N_10602);
nor U11714 (N_11714,N_10135,N_10648);
and U11715 (N_11715,N_9728,N_10732);
nand U11716 (N_11716,N_10381,N_9610);
nor U11717 (N_11717,N_10028,N_9754);
or U11718 (N_11718,N_10446,N_9632);
nand U11719 (N_11719,N_10573,N_10098);
or U11720 (N_11720,N_10699,N_10651);
nor U11721 (N_11721,N_9772,N_9807);
xnor U11722 (N_11722,N_10577,N_10441);
nand U11723 (N_11723,N_9844,N_9946);
nand U11724 (N_11724,N_10042,N_10525);
nor U11725 (N_11725,N_10407,N_10507);
or U11726 (N_11726,N_9801,N_10679);
xnor U11727 (N_11727,N_10755,N_10294);
nor U11728 (N_11728,N_10441,N_10504);
nor U11729 (N_11729,N_10169,N_9867);
xor U11730 (N_11730,N_10375,N_9700);
nor U11731 (N_11731,N_10527,N_9849);
nand U11732 (N_11732,N_10319,N_9680);
nor U11733 (N_11733,N_9950,N_10417);
xor U11734 (N_11734,N_10543,N_10343);
nand U11735 (N_11735,N_10376,N_10238);
and U11736 (N_11736,N_9770,N_10504);
and U11737 (N_11737,N_9748,N_9975);
nand U11738 (N_11738,N_9809,N_10316);
nand U11739 (N_11739,N_10193,N_10777);
nor U11740 (N_11740,N_10772,N_10606);
nand U11741 (N_11741,N_10730,N_10134);
nor U11742 (N_11742,N_10346,N_9649);
xnor U11743 (N_11743,N_10570,N_10560);
and U11744 (N_11744,N_10728,N_10482);
and U11745 (N_11745,N_10745,N_9764);
xnor U11746 (N_11746,N_10267,N_9996);
xor U11747 (N_11747,N_10192,N_10664);
xor U11748 (N_11748,N_9742,N_10111);
nand U11749 (N_11749,N_10721,N_10500);
xor U11750 (N_11750,N_9817,N_9776);
nor U11751 (N_11751,N_10628,N_10062);
nor U11752 (N_11752,N_10301,N_10583);
nor U11753 (N_11753,N_9643,N_10419);
and U11754 (N_11754,N_10187,N_10719);
or U11755 (N_11755,N_10382,N_10581);
nand U11756 (N_11756,N_9790,N_10422);
nand U11757 (N_11757,N_10039,N_9975);
xor U11758 (N_11758,N_10073,N_10502);
and U11759 (N_11759,N_10226,N_9912);
nor U11760 (N_11760,N_10236,N_9625);
or U11761 (N_11761,N_10763,N_10748);
nand U11762 (N_11762,N_10227,N_10535);
or U11763 (N_11763,N_10526,N_10068);
nand U11764 (N_11764,N_10640,N_10779);
or U11765 (N_11765,N_10156,N_10190);
xor U11766 (N_11766,N_9646,N_10205);
xor U11767 (N_11767,N_10129,N_10281);
nor U11768 (N_11768,N_9872,N_10561);
or U11769 (N_11769,N_10779,N_10096);
nand U11770 (N_11770,N_10510,N_10194);
or U11771 (N_11771,N_9623,N_10762);
or U11772 (N_11772,N_10378,N_10603);
and U11773 (N_11773,N_10368,N_9903);
xnor U11774 (N_11774,N_10373,N_10025);
or U11775 (N_11775,N_10310,N_10033);
xnor U11776 (N_11776,N_10616,N_9747);
nor U11777 (N_11777,N_10479,N_9739);
nor U11778 (N_11778,N_10333,N_10332);
xnor U11779 (N_11779,N_10363,N_10238);
or U11780 (N_11780,N_9889,N_9877);
or U11781 (N_11781,N_9999,N_10260);
or U11782 (N_11782,N_10552,N_10276);
nand U11783 (N_11783,N_9864,N_9941);
or U11784 (N_11784,N_10627,N_10048);
nand U11785 (N_11785,N_10398,N_10046);
and U11786 (N_11786,N_9732,N_10488);
xnor U11787 (N_11787,N_10593,N_10564);
nor U11788 (N_11788,N_10072,N_10638);
and U11789 (N_11789,N_9767,N_10027);
and U11790 (N_11790,N_10072,N_10080);
nand U11791 (N_11791,N_10734,N_9643);
nor U11792 (N_11792,N_9834,N_9781);
xor U11793 (N_11793,N_10002,N_10574);
nand U11794 (N_11794,N_10199,N_10343);
nor U11795 (N_11795,N_9895,N_10079);
nor U11796 (N_11796,N_9739,N_9933);
nor U11797 (N_11797,N_9660,N_10270);
nor U11798 (N_11798,N_10782,N_10454);
nand U11799 (N_11799,N_9919,N_10412);
xor U11800 (N_11800,N_9615,N_10366);
or U11801 (N_11801,N_10156,N_10504);
xnor U11802 (N_11802,N_9751,N_9779);
or U11803 (N_11803,N_10528,N_10201);
nand U11804 (N_11804,N_10338,N_10016);
and U11805 (N_11805,N_10506,N_10603);
nor U11806 (N_11806,N_10114,N_10749);
nand U11807 (N_11807,N_10370,N_10641);
or U11808 (N_11808,N_10456,N_9847);
nor U11809 (N_11809,N_10730,N_9641);
nand U11810 (N_11810,N_9783,N_10571);
nand U11811 (N_11811,N_10492,N_10219);
xor U11812 (N_11812,N_10045,N_10750);
or U11813 (N_11813,N_10315,N_10661);
nor U11814 (N_11814,N_9764,N_10292);
xor U11815 (N_11815,N_10222,N_9791);
xor U11816 (N_11816,N_10110,N_10671);
or U11817 (N_11817,N_10417,N_10415);
or U11818 (N_11818,N_10712,N_9888);
xor U11819 (N_11819,N_10195,N_9720);
nor U11820 (N_11820,N_10163,N_9772);
nor U11821 (N_11821,N_10391,N_10797);
nor U11822 (N_11822,N_9872,N_10043);
or U11823 (N_11823,N_10689,N_10332);
or U11824 (N_11824,N_10390,N_10689);
nor U11825 (N_11825,N_10555,N_10451);
and U11826 (N_11826,N_10321,N_9821);
xnor U11827 (N_11827,N_10524,N_10045);
or U11828 (N_11828,N_10623,N_10378);
nor U11829 (N_11829,N_10384,N_10010);
nand U11830 (N_11830,N_9813,N_10079);
nand U11831 (N_11831,N_9942,N_10451);
nor U11832 (N_11832,N_9989,N_9660);
nand U11833 (N_11833,N_10555,N_10155);
and U11834 (N_11834,N_9942,N_10718);
and U11835 (N_11835,N_10400,N_9869);
xnor U11836 (N_11836,N_9722,N_10166);
or U11837 (N_11837,N_10653,N_10045);
nand U11838 (N_11838,N_10387,N_10216);
and U11839 (N_11839,N_10253,N_10258);
nor U11840 (N_11840,N_10222,N_9915);
nor U11841 (N_11841,N_9729,N_10491);
nand U11842 (N_11842,N_10073,N_9969);
xor U11843 (N_11843,N_10276,N_10339);
and U11844 (N_11844,N_9852,N_10470);
and U11845 (N_11845,N_10415,N_10611);
and U11846 (N_11846,N_10224,N_10042);
or U11847 (N_11847,N_10795,N_10626);
xor U11848 (N_11848,N_10478,N_10132);
nor U11849 (N_11849,N_9890,N_10093);
or U11850 (N_11850,N_9972,N_10416);
nand U11851 (N_11851,N_10792,N_10020);
xnor U11852 (N_11852,N_10484,N_9624);
or U11853 (N_11853,N_9870,N_10327);
and U11854 (N_11854,N_10181,N_10544);
nor U11855 (N_11855,N_9647,N_9935);
nand U11856 (N_11856,N_9653,N_10745);
or U11857 (N_11857,N_10576,N_9845);
nand U11858 (N_11858,N_9953,N_9713);
xnor U11859 (N_11859,N_10414,N_10250);
nand U11860 (N_11860,N_10171,N_10263);
nand U11861 (N_11861,N_10338,N_10553);
and U11862 (N_11862,N_10693,N_9749);
nor U11863 (N_11863,N_10093,N_10167);
nor U11864 (N_11864,N_9619,N_10579);
and U11865 (N_11865,N_9940,N_10250);
xnor U11866 (N_11866,N_10204,N_10721);
nor U11867 (N_11867,N_9861,N_10244);
nand U11868 (N_11868,N_9830,N_9840);
xnor U11869 (N_11869,N_10446,N_10797);
xnor U11870 (N_11870,N_9631,N_10100);
or U11871 (N_11871,N_9996,N_9987);
nor U11872 (N_11872,N_9635,N_9910);
nand U11873 (N_11873,N_10573,N_9642);
nand U11874 (N_11874,N_9635,N_9678);
and U11875 (N_11875,N_10256,N_10654);
or U11876 (N_11876,N_9853,N_10713);
xnor U11877 (N_11877,N_10715,N_10357);
nor U11878 (N_11878,N_10031,N_10081);
and U11879 (N_11879,N_10413,N_10589);
and U11880 (N_11880,N_10568,N_10347);
or U11881 (N_11881,N_9656,N_10153);
xor U11882 (N_11882,N_9856,N_10408);
xor U11883 (N_11883,N_10005,N_9602);
xor U11884 (N_11884,N_10596,N_10086);
nor U11885 (N_11885,N_10663,N_10299);
xor U11886 (N_11886,N_9923,N_9673);
nand U11887 (N_11887,N_10199,N_10072);
and U11888 (N_11888,N_10156,N_9827);
and U11889 (N_11889,N_10667,N_9789);
and U11890 (N_11890,N_10551,N_10060);
or U11891 (N_11891,N_10652,N_9770);
nor U11892 (N_11892,N_9691,N_10073);
nand U11893 (N_11893,N_9827,N_10148);
nor U11894 (N_11894,N_10286,N_10486);
and U11895 (N_11895,N_10200,N_9702);
xnor U11896 (N_11896,N_10489,N_9983);
nor U11897 (N_11897,N_10131,N_9891);
nand U11898 (N_11898,N_10206,N_10652);
and U11899 (N_11899,N_10171,N_10205);
or U11900 (N_11900,N_10311,N_10148);
and U11901 (N_11901,N_10562,N_10752);
nor U11902 (N_11902,N_10578,N_10673);
or U11903 (N_11903,N_10787,N_10135);
or U11904 (N_11904,N_9629,N_10370);
nand U11905 (N_11905,N_9627,N_9874);
or U11906 (N_11906,N_10456,N_10759);
nand U11907 (N_11907,N_10049,N_10075);
and U11908 (N_11908,N_9833,N_10349);
and U11909 (N_11909,N_9986,N_9683);
nand U11910 (N_11910,N_10017,N_10030);
nor U11911 (N_11911,N_10404,N_10137);
or U11912 (N_11912,N_9688,N_10032);
or U11913 (N_11913,N_10701,N_9605);
nor U11914 (N_11914,N_10223,N_10066);
nand U11915 (N_11915,N_10514,N_10426);
nand U11916 (N_11916,N_9918,N_10468);
nor U11917 (N_11917,N_10267,N_10321);
nand U11918 (N_11918,N_10067,N_10314);
nor U11919 (N_11919,N_10348,N_9649);
or U11920 (N_11920,N_9951,N_10425);
and U11921 (N_11921,N_10257,N_10551);
nand U11922 (N_11922,N_10136,N_10675);
or U11923 (N_11923,N_9671,N_10715);
nor U11924 (N_11924,N_9722,N_9970);
nor U11925 (N_11925,N_10684,N_10347);
and U11926 (N_11926,N_9927,N_10635);
and U11927 (N_11927,N_9703,N_9751);
and U11928 (N_11928,N_10709,N_10105);
nand U11929 (N_11929,N_10579,N_9887);
nand U11930 (N_11930,N_9934,N_10557);
nor U11931 (N_11931,N_10582,N_9627);
or U11932 (N_11932,N_10522,N_10285);
nor U11933 (N_11933,N_10027,N_9893);
nor U11934 (N_11934,N_10239,N_10712);
and U11935 (N_11935,N_10519,N_9998);
or U11936 (N_11936,N_10780,N_10699);
and U11937 (N_11937,N_9920,N_10023);
and U11938 (N_11938,N_9977,N_9624);
xnor U11939 (N_11939,N_10292,N_10358);
nand U11940 (N_11940,N_10077,N_9623);
xor U11941 (N_11941,N_9867,N_10748);
nor U11942 (N_11942,N_10215,N_10652);
and U11943 (N_11943,N_10170,N_10792);
nor U11944 (N_11944,N_10445,N_10253);
or U11945 (N_11945,N_10004,N_10051);
or U11946 (N_11946,N_10335,N_10246);
and U11947 (N_11947,N_9636,N_10437);
and U11948 (N_11948,N_10107,N_9777);
and U11949 (N_11949,N_9858,N_10661);
nand U11950 (N_11950,N_10223,N_10300);
and U11951 (N_11951,N_9614,N_9815);
and U11952 (N_11952,N_9646,N_10480);
nand U11953 (N_11953,N_9771,N_10462);
xor U11954 (N_11954,N_10107,N_10028);
xnor U11955 (N_11955,N_10226,N_9627);
nor U11956 (N_11956,N_10156,N_10192);
xor U11957 (N_11957,N_9603,N_10377);
nand U11958 (N_11958,N_10206,N_9762);
and U11959 (N_11959,N_9816,N_9660);
and U11960 (N_11960,N_10318,N_10553);
xnor U11961 (N_11961,N_9630,N_10463);
nand U11962 (N_11962,N_10112,N_9935);
and U11963 (N_11963,N_10383,N_9644);
nor U11964 (N_11964,N_9814,N_9916);
and U11965 (N_11965,N_10628,N_9607);
and U11966 (N_11966,N_10157,N_9629);
or U11967 (N_11967,N_10194,N_9996);
and U11968 (N_11968,N_10596,N_10582);
nor U11969 (N_11969,N_9699,N_9869);
nor U11970 (N_11970,N_9605,N_9919);
and U11971 (N_11971,N_9897,N_10212);
nor U11972 (N_11972,N_9606,N_10377);
xnor U11973 (N_11973,N_10711,N_9914);
or U11974 (N_11974,N_10250,N_10625);
or U11975 (N_11975,N_9872,N_9977);
or U11976 (N_11976,N_10720,N_10749);
and U11977 (N_11977,N_10007,N_9733);
nand U11978 (N_11978,N_9676,N_9621);
or U11979 (N_11979,N_9601,N_10087);
nor U11980 (N_11980,N_10190,N_9915);
nand U11981 (N_11981,N_9963,N_10595);
nand U11982 (N_11982,N_10456,N_10680);
xor U11983 (N_11983,N_9812,N_10190);
or U11984 (N_11984,N_10763,N_10637);
nand U11985 (N_11985,N_10447,N_10308);
nor U11986 (N_11986,N_9600,N_10647);
nor U11987 (N_11987,N_9870,N_10438);
nor U11988 (N_11988,N_9890,N_10381);
xnor U11989 (N_11989,N_10384,N_10011);
or U11990 (N_11990,N_10206,N_10767);
or U11991 (N_11991,N_10750,N_10485);
or U11992 (N_11992,N_10568,N_10758);
nand U11993 (N_11993,N_10452,N_9989);
nor U11994 (N_11994,N_10726,N_10233);
and U11995 (N_11995,N_10593,N_10084);
xor U11996 (N_11996,N_10653,N_10441);
nor U11997 (N_11997,N_10744,N_10731);
nand U11998 (N_11998,N_10104,N_10169);
xor U11999 (N_11999,N_10103,N_9653);
xor U12000 (N_12000,N_10924,N_11974);
xor U12001 (N_12001,N_11101,N_11788);
nor U12002 (N_12002,N_11634,N_11786);
or U12003 (N_12003,N_11758,N_11376);
nor U12004 (N_12004,N_11315,N_11585);
nand U12005 (N_12005,N_11571,N_10890);
or U12006 (N_12006,N_11207,N_11105);
xnor U12007 (N_12007,N_11240,N_11936);
nor U12008 (N_12008,N_11458,N_11146);
nand U12009 (N_12009,N_11836,N_10854);
nand U12010 (N_12010,N_10858,N_11116);
nand U12011 (N_12011,N_11384,N_11297);
nor U12012 (N_12012,N_10913,N_11679);
nand U12013 (N_12013,N_11493,N_11397);
and U12014 (N_12014,N_11418,N_11885);
or U12015 (N_12015,N_11552,N_11305);
nand U12016 (N_12016,N_11850,N_11076);
xor U12017 (N_12017,N_11486,N_11094);
nand U12018 (N_12018,N_11524,N_11115);
or U12019 (N_12019,N_11515,N_11341);
and U12020 (N_12020,N_10925,N_11595);
xor U12021 (N_12021,N_11330,N_11112);
nor U12022 (N_12022,N_10977,N_11917);
nor U12023 (N_12023,N_11815,N_11431);
nor U12024 (N_12024,N_11616,N_11513);
xnor U12025 (N_12025,N_10865,N_10881);
or U12026 (N_12026,N_11642,N_11811);
and U12027 (N_12027,N_11137,N_11672);
nand U12028 (N_12028,N_11166,N_11401);
and U12029 (N_12029,N_11230,N_11406);
nand U12030 (N_12030,N_11589,N_10888);
xnor U12031 (N_12031,N_11650,N_11242);
xor U12032 (N_12032,N_11074,N_11109);
or U12033 (N_12033,N_11864,N_11900);
or U12034 (N_12034,N_11689,N_11476);
and U12035 (N_12035,N_10963,N_11421);
nand U12036 (N_12036,N_10841,N_10990);
xnor U12037 (N_12037,N_11235,N_11065);
nor U12038 (N_12038,N_11430,N_11728);
xor U12039 (N_12039,N_10976,N_11807);
and U12040 (N_12040,N_11208,N_11898);
xor U12041 (N_12041,N_11055,N_11972);
xnor U12042 (N_12042,N_11363,N_11499);
or U12043 (N_12043,N_11390,N_11381);
nand U12044 (N_12044,N_11921,N_10823);
nor U12045 (N_12045,N_10973,N_10941);
and U12046 (N_12046,N_11444,N_11959);
or U12047 (N_12047,N_11110,N_11203);
nor U12048 (N_12048,N_10812,N_11837);
xor U12049 (N_12049,N_11429,N_11323);
or U12050 (N_12050,N_11644,N_11639);
and U12051 (N_12051,N_10998,N_10831);
and U12052 (N_12052,N_11262,N_11206);
and U12053 (N_12053,N_11828,N_11988);
nand U12054 (N_12054,N_11852,N_11928);
or U12055 (N_12055,N_11425,N_11286);
nor U12056 (N_12056,N_11756,N_11370);
xor U12057 (N_12057,N_11251,N_10920);
xnor U12058 (N_12058,N_11924,N_11308);
nand U12059 (N_12059,N_11502,N_11749);
nor U12060 (N_12060,N_10992,N_11079);
xnor U12061 (N_12061,N_11598,N_11708);
or U12062 (N_12062,N_11260,N_10949);
nand U12063 (N_12063,N_10936,N_10846);
xor U12064 (N_12064,N_11606,N_11283);
xor U12065 (N_12065,N_10938,N_10814);
nand U12066 (N_12066,N_11744,N_10933);
or U12067 (N_12067,N_11803,N_11880);
nand U12068 (N_12068,N_11800,N_11818);
nand U12069 (N_12069,N_11769,N_11371);
nor U12070 (N_12070,N_11647,N_11239);
or U12071 (N_12071,N_10954,N_11466);
nor U12072 (N_12072,N_11141,N_11993);
nand U12073 (N_12073,N_11142,N_11078);
or U12074 (N_12074,N_11625,N_11271);
or U12075 (N_12075,N_11333,N_11465);
and U12076 (N_12076,N_11931,N_11056);
or U12077 (N_12077,N_11857,N_11562);
nor U12078 (N_12078,N_11643,N_11523);
and U12079 (N_12079,N_11839,N_10826);
and U12080 (N_12080,N_11680,N_11165);
nor U12081 (N_12081,N_10910,N_11001);
or U12082 (N_12082,N_11194,N_11942);
or U12083 (N_12083,N_11045,N_11970);
nor U12084 (N_12084,N_11557,N_10906);
or U12085 (N_12085,N_11368,N_11057);
xor U12086 (N_12086,N_11657,N_11973);
and U12087 (N_12087,N_10830,N_10978);
or U12088 (N_12088,N_11681,N_11159);
nor U12089 (N_12089,N_11725,N_11211);
and U12090 (N_12090,N_10970,N_11426);
nand U12091 (N_12091,N_11899,N_11303);
xor U12092 (N_12092,N_11741,N_11064);
nand U12093 (N_12093,N_11982,N_11382);
and U12094 (N_12094,N_10852,N_11549);
and U12095 (N_12095,N_11578,N_11983);
xnor U12096 (N_12096,N_10834,N_11121);
nand U12097 (N_12097,N_11325,N_11066);
and U12098 (N_12098,N_11449,N_11174);
xnor U12099 (N_12099,N_11574,N_11539);
nor U12100 (N_12100,N_11813,N_11577);
and U12101 (N_12101,N_11007,N_11118);
nand U12102 (N_12102,N_11683,N_11468);
nand U12103 (N_12103,N_11386,N_11560);
xor U12104 (N_12104,N_11534,N_11510);
and U12105 (N_12105,N_11164,N_11031);
nand U12106 (N_12106,N_11307,N_11409);
and U12107 (N_12107,N_11348,N_11796);
nand U12108 (N_12108,N_11313,N_11227);
nor U12109 (N_12109,N_11992,N_11359);
and U12110 (N_12110,N_11096,N_11961);
nand U12111 (N_12111,N_11002,N_11946);
or U12112 (N_12112,N_11608,N_11160);
or U12113 (N_12113,N_11209,N_11067);
and U12114 (N_12114,N_10944,N_10898);
nor U12115 (N_12115,N_11491,N_11025);
nor U12116 (N_12116,N_11049,N_11573);
or U12117 (N_12117,N_10908,N_11331);
nand U12118 (N_12118,N_11790,N_11047);
nor U12119 (N_12119,N_11438,N_11347);
and U12120 (N_12120,N_11247,N_11334);
nand U12121 (N_12121,N_11185,N_11123);
xnor U12122 (N_12122,N_11729,N_11263);
or U12123 (N_12123,N_11832,N_11645);
and U12124 (N_12124,N_10979,N_11820);
nor U12125 (N_12125,N_11296,N_11191);
nor U12126 (N_12126,N_11016,N_11231);
and U12127 (N_12127,N_11692,N_11762);
or U12128 (N_12128,N_11257,N_11099);
xor U12129 (N_12129,N_11776,N_10849);
nor U12130 (N_12130,N_11633,N_11582);
nand U12131 (N_12131,N_11339,N_11352);
nand U12132 (N_12132,N_11117,N_10878);
nand U12133 (N_12133,N_11895,N_10885);
nand U12134 (N_12134,N_10848,N_11148);
nand U12135 (N_12135,N_11402,N_11746);
and U12136 (N_12136,N_11326,N_11457);
or U12137 (N_12137,N_11304,N_11222);
or U12138 (N_12138,N_11398,N_10935);
and U12139 (N_12139,N_11628,N_11226);
nand U12140 (N_12140,N_11675,N_11254);
xor U12141 (N_12141,N_11399,N_11291);
nor U12142 (N_12142,N_10959,N_11999);
nor U12143 (N_12143,N_11918,N_11542);
nor U12144 (N_12144,N_11039,N_10872);
or U12145 (N_12145,N_11075,N_11274);
and U12146 (N_12146,N_11266,N_11033);
nand U12147 (N_12147,N_11113,N_11482);
xnor U12148 (N_12148,N_11705,N_10887);
nand U12149 (N_12149,N_11414,N_11671);
nand U12150 (N_12150,N_11463,N_11152);
and U12151 (N_12151,N_11810,N_11355);
or U12152 (N_12152,N_10932,N_11521);
and U12153 (N_12153,N_11914,N_11157);
nor U12154 (N_12154,N_11238,N_11353);
xor U12155 (N_12155,N_11459,N_11801);
xnor U12156 (N_12156,N_11269,N_11345);
nor U12157 (N_12157,N_11052,N_11816);
or U12158 (N_12158,N_11854,N_11825);
nand U12159 (N_12159,N_10836,N_11279);
nand U12160 (N_12160,N_10859,N_11522);
and U12161 (N_12161,N_11095,N_11130);
nor U12162 (N_12162,N_11173,N_11456);
and U12163 (N_12163,N_11541,N_11479);
xor U12164 (N_12164,N_11365,N_11719);
nor U12165 (N_12165,N_10981,N_10964);
and U12166 (N_12166,N_11546,N_11088);
nand U12167 (N_12167,N_11621,N_11048);
or U12168 (N_12168,N_10987,N_11829);
nor U12169 (N_12169,N_11437,N_11467);
and U12170 (N_12170,N_11484,N_11528);
and U12171 (N_12171,N_11878,N_10929);
nor U12172 (N_12172,N_10824,N_11270);
nor U12173 (N_12173,N_11193,N_11953);
nor U12174 (N_12174,N_11591,N_11424);
nand U12175 (N_12175,N_11128,N_11336);
or U12176 (N_12176,N_11893,N_11250);
or U12177 (N_12177,N_11518,N_11195);
nor U12178 (N_12178,N_11704,N_11782);
and U12179 (N_12179,N_11155,N_11904);
xor U12180 (N_12180,N_11883,N_11220);
and U12181 (N_12181,N_11178,N_11844);
or U12182 (N_12182,N_11485,N_11434);
and U12183 (N_12183,N_11190,N_11935);
nand U12184 (N_12184,N_10983,N_11216);
xnor U12185 (N_12185,N_11342,N_10850);
and U12186 (N_12186,N_11501,N_11791);
xnor U12187 (N_12187,N_11553,N_11393);
and U12188 (N_12188,N_11879,N_11912);
nor U12189 (N_12189,N_11356,N_11873);
or U12190 (N_12190,N_10907,N_11085);
or U12191 (N_12191,N_10922,N_11960);
or U12192 (N_12192,N_11941,N_11614);
or U12193 (N_12193,N_11752,N_10909);
and U12194 (N_12194,N_11619,N_10835);
xnor U12195 (N_12195,N_10996,N_11439);
nand U12196 (N_12196,N_11046,N_10893);
nand U12197 (N_12197,N_11389,N_11394);
and U12198 (N_12198,N_11391,N_11023);
xor U12199 (N_12199,N_11884,N_11742);
or U12200 (N_12200,N_11495,N_11395);
nand U12201 (N_12201,N_11122,N_11830);
and U12202 (N_12202,N_11221,N_10937);
or U12203 (N_12203,N_11234,N_11963);
nor U12204 (N_12204,N_11171,N_11600);
and U12205 (N_12205,N_10974,N_11529);
xor U12206 (N_12206,N_11772,N_11609);
nor U12207 (N_12207,N_11224,N_11855);
nor U12208 (N_12208,N_10811,N_11814);
nor U12209 (N_12209,N_11944,N_11452);
or U12210 (N_12210,N_11204,N_11134);
nand U12211 (N_12211,N_11835,N_11322);
nand U12212 (N_12212,N_10809,N_11505);
xnor U12213 (N_12213,N_11590,N_11416);
nand U12214 (N_12214,N_11951,N_11487);
nor U12215 (N_12215,N_11874,N_11599);
nor U12216 (N_12216,N_11903,N_11584);
and U12217 (N_12217,N_11785,N_10952);
xor U12218 (N_12218,N_11998,N_11470);
and U12219 (N_12219,N_10918,N_11610);
and U12220 (N_12220,N_10871,N_11201);
or U12221 (N_12221,N_11965,N_11379);
and U12222 (N_12222,N_10877,N_11346);
or U12223 (N_12223,N_11509,N_11841);
or U12224 (N_12224,N_11915,N_11710);
or U12225 (N_12225,N_11964,N_10942);
nor U12226 (N_12226,N_11858,N_10864);
or U12227 (N_12227,N_11956,N_11673);
xor U12228 (N_12228,N_11943,N_11255);
or U12229 (N_12229,N_10883,N_11554);
xor U12230 (N_12230,N_11127,N_11663);
nor U12231 (N_12231,N_10901,N_11335);
and U12232 (N_12232,N_11503,N_11278);
and U12233 (N_12233,N_11580,N_11133);
or U12234 (N_12234,N_11259,N_10803);
xor U12235 (N_12235,N_11905,N_11911);
xnor U12236 (N_12236,N_11205,N_11268);
or U12237 (N_12237,N_11775,N_11298);
or U12238 (N_12238,N_11795,N_11847);
and U12239 (N_12239,N_10863,N_11954);
xor U12240 (N_12240,N_11405,N_11177);
nor U12241 (N_12241,N_11531,N_11738);
xor U12242 (N_12242,N_10968,N_11068);
xor U12243 (N_12243,N_11442,N_10904);
xnor U12244 (N_12244,N_10912,N_11385);
and U12245 (N_12245,N_11071,N_11312);
xor U12246 (N_12246,N_11721,N_10874);
nor U12247 (N_12247,N_11277,N_11267);
and U12248 (N_12248,N_10905,N_11629);
or U12249 (N_12249,N_11454,N_11472);
nor U12250 (N_12250,N_11849,N_11490);
or U12251 (N_12251,N_11243,N_11575);
nor U12252 (N_12252,N_11035,N_11525);
nor U12253 (N_12253,N_11198,N_11626);
xnor U12254 (N_12254,N_11189,N_11215);
nand U12255 (N_12255,N_11512,N_11151);
and U12256 (N_12256,N_11061,N_11572);
nand U12257 (N_12257,N_11703,N_11210);
xor U12258 (N_12258,N_11135,N_11908);
xnor U12259 (N_12259,N_11831,N_11093);
nand U12260 (N_12260,N_11767,N_11299);
xor U12261 (N_12261,N_10896,N_11868);
xnor U12262 (N_12262,N_11916,N_11403);
nor U12263 (N_12263,N_11865,N_10965);
and U12264 (N_12264,N_11739,N_11038);
and U12265 (N_12265,N_11318,N_11496);
nand U12266 (N_12266,N_11996,N_11455);
nor U12267 (N_12267,N_10860,N_11668);
nor U12268 (N_12268,N_11981,N_10808);
nor U12269 (N_12269,N_11295,N_10880);
or U12270 (N_12270,N_11760,N_10839);
or U12271 (N_12271,N_11656,N_11929);
and U12272 (N_12272,N_11324,N_10967);
xnor U12273 (N_12273,N_10923,N_11053);
or U12274 (N_12274,N_11292,N_10889);
nand U12275 (N_12275,N_11514,N_11558);
or U12276 (N_12276,N_11720,N_11723);
xor U12277 (N_12277,N_11217,N_11073);
xor U12278 (N_12278,N_10927,N_11926);
or U12279 (N_12279,N_11889,N_10984);
xor U12280 (N_12280,N_11990,N_11372);
and U12281 (N_12281,N_10825,N_10948);
and U12282 (N_12282,N_10991,N_10842);
nor U12283 (N_12283,N_11561,N_11184);
nand U12284 (N_12284,N_10817,N_11833);
xor U12285 (N_12285,N_10828,N_11197);
nor U12286 (N_12286,N_11724,N_11149);
nor U12287 (N_12287,N_11842,N_11138);
xor U12288 (N_12288,N_11748,N_11550);
or U12289 (N_12289,N_11492,N_11202);
nor U12290 (N_12290,N_11764,N_11925);
or U12291 (N_12291,N_11991,N_10801);
and U12292 (N_12292,N_11771,N_11131);
nor U12293 (N_12293,N_11700,N_11694);
nand U12294 (N_12294,N_10816,N_11041);
nor U12295 (N_12295,N_11103,N_11586);
nor U12296 (N_12296,N_11169,N_11797);
nand U12297 (N_12297,N_11684,N_11350);
and U12298 (N_12298,N_11611,N_11285);
xor U12299 (N_12299,N_11294,N_11119);
xnor U12300 (N_12300,N_11949,N_11374);
xnor U12301 (N_12301,N_11364,N_11765);
nand U12302 (N_12302,N_11375,N_11527);
nor U12303 (N_12303,N_11034,N_11114);
nand U12304 (N_12304,N_11696,N_11624);
or U12305 (N_12305,N_11618,N_11761);
and U12306 (N_12306,N_11070,N_11986);
nand U12307 (N_12307,N_11713,N_10827);
nand U12308 (N_12308,N_11413,N_11699);
nand U12309 (N_12309,N_11281,N_11245);
and U12310 (N_12310,N_11175,N_11932);
and U12311 (N_12311,N_11688,N_11404);
or U12312 (N_12312,N_11661,N_11664);
nor U12313 (N_12313,N_11697,N_11731);
or U12314 (N_12314,N_11587,N_11877);
nand U12315 (N_12315,N_10969,N_10891);
nor U12316 (N_12316,N_11922,N_11930);
xnor U12317 (N_12317,N_10997,N_11017);
xor U12318 (N_12318,N_10899,N_11338);
xnor U12319 (N_12319,N_11106,N_11827);
and U12320 (N_12320,N_11623,N_11780);
nand U12321 (N_12321,N_11845,N_11881);
and U12322 (N_12322,N_10869,N_11120);
or U12323 (N_12323,N_11870,N_11716);
nand U12324 (N_12324,N_11517,N_11987);
or U12325 (N_12325,N_11176,N_11754);
xnor U12326 (N_12326,N_11907,N_11667);
or U12327 (N_12327,N_11863,N_11583);
xnor U12328 (N_12328,N_10813,N_11798);
nor U12329 (N_12329,N_10962,N_11594);
nor U12330 (N_12330,N_11265,N_11344);
or U12331 (N_12331,N_11826,N_11736);
or U12332 (N_12332,N_11427,N_11436);
nand U12333 (N_12333,N_11655,N_11062);
and U12334 (N_12334,N_11792,N_11971);
nor U12335 (N_12335,N_11010,N_11407);
and U12336 (N_12336,N_11107,N_11415);
or U12337 (N_12337,N_11851,N_11984);
xnor U12338 (N_12338,N_11024,N_11004);
and U12339 (N_12339,N_10818,N_11050);
nor U12340 (N_12340,N_11125,N_11773);
nand U12341 (N_12341,N_11275,N_11637);
or U12342 (N_12342,N_11605,N_11687);
xor U12343 (N_12343,N_10911,N_11838);
xor U12344 (N_12344,N_11237,N_11727);
or U12345 (N_12345,N_11223,N_10895);
xnor U12346 (N_12346,N_11834,N_11090);
nor U12347 (N_12347,N_11378,N_11464);
nor U12348 (N_12348,N_11293,N_11653);
xnor U12349 (N_12349,N_11241,N_11480);
and U12350 (N_12350,N_11411,N_11301);
xnor U12351 (N_12351,N_11779,N_11638);
or U12352 (N_12352,N_10945,N_11678);
and U12353 (N_12353,N_10876,N_11540);
nor U12354 (N_12354,N_11670,N_10971);
nand U12355 (N_12355,N_11567,N_11327);
nand U12356 (N_12356,N_11979,N_11581);
xnor U12357 (N_12357,N_10999,N_10833);
or U12358 (N_12358,N_11648,N_11140);
or U12359 (N_12359,N_10882,N_11632);
xnor U12360 (N_12360,N_11471,N_10916);
and U12361 (N_12361,N_11659,N_10822);
nand U12362 (N_12362,N_10838,N_11866);
nand U12363 (N_12363,N_11923,N_10994);
nand U12364 (N_12364,N_11498,N_11218);
nor U12365 (N_12365,N_11441,N_11737);
xnor U12366 (N_12366,N_11008,N_11317);
or U12367 (N_12367,N_11869,N_11937);
and U12368 (N_12368,N_11494,N_11462);
nor U12369 (N_12369,N_11387,N_11026);
xor U12370 (N_12370,N_11896,N_10947);
nor U12371 (N_12371,N_11186,N_11989);
or U12372 (N_12372,N_11853,N_11715);
nand U12373 (N_12373,N_11955,N_11019);
nor U12374 (N_12374,N_11566,N_10903);
nor U12375 (N_12375,N_11288,N_11511);
nor U12376 (N_12376,N_10820,N_11707);
nand U12377 (N_12377,N_10960,N_11030);
nand U12378 (N_12378,N_11640,N_10917);
xor U12379 (N_12379,N_11958,N_11947);
xor U12380 (N_12380,N_10931,N_11000);
and U12381 (N_12381,N_11132,N_11040);
or U12382 (N_12382,N_10840,N_11995);
nor U12383 (N_12383,N_11787,N_11630);
or U12384 (N_12384,N_11244,N_11804);
and U12385 (N_12385,N_11538,N_11662);
or U12386 (N_12386,N_11927,N_10915);
and U12387 (N_12387,N_11383,N_11332);
nand U12388 (N_12388,N_11565,N_11446);
nor U12389 (N_12389,N_11232,N_11280);
xnor U12390 (N_12390,N_11612,N_11473);
nand U12391 (N_12391,N_11840,N_11445);
xnor U12392 (N_12392,N_11077,N_11154);
nand U12393 (N_12393,N_11172,N_11848);
or U12394 (N_12394,N_11256,N_11945);
and U12395 (N_12395,N_10926,N_11952);
xor U12396 (N_12396,N_10875,N_11570);
or U12397 (N_12397,N_11913,N_11711);
or U12398 (N_12398,N_10857,N_11219);
nand U12399 (N_12399,N_11819,N_10845);
or U12400 (N_12400,N_10934,N_11613);
and U12401 (N_12401,N_11028,N_11812);
nand U12402 (N_12402,N_11082,N_11617);
xnor U12403 (N_12403,N_10807,N_11443);
nand U12404 (N_12404,N_11579,N_11015);
xor U12405 (N_12405,N_11083,N_11063);
nand U12406 (N_12406,N_10868,N_11568);
and U12407 (N_12407,N_11902,N_10930);
or U12408 (N_12408,N_11069,N_11481);
nor U12409 (N_12409,N_11183,N_10886);
nor U12410 (N_12410,N_10961,N_11060);
nand U12411 (N_12411,N_10940,N_11168);
or U12412 (N_12412,N_11516,N_11690);
nand U12413 (N_12413,N_11314,N_11145);
and U12414 (N_12414,N_11793,N_11111);
and U12415 (N_12415,N_11506,N_11563);
nor U12416 (N_12416,N_11328,N_11351);
xnor U12417 (N_12417,N_10921,N_11876);
nor U12418 (N_12418,N_11592,N_11763);
nor U12419 (N_12419,N_11919,N_11036);
and U12420 (N_12420,N_11702,N_10829);
xor U12421 (N_12421,N_11320,N_10861);
nand U12422 (N_12422,N_11802,N_11894);
nor U12423 (N_12423,N_11362,N_11284);
and U12424 (N_12424,N_10985,N_11520);
or U12425 (N_12425,N_11751,N_11282);
xor U12426 (N_12426,N_11593,N_11717);
and U12427 (N_12427,N_11272,N_11504);
and U12428 (N_12428,N_10975,N_11537);
or U12429 (N_12429,N_11377,N_11423);
nand U12430 (N_12430,N_11369,N_11722);
nand U12431 (N_12431,N_11044,N_10900);
or U12432 (N_12432,N_11229,N_10862);
xor U12433 (N_12433,N_11451,N_11658);
nor U12434 (N_12434,N_11199,N_11156);
nand U12435 (N_12435,N_11920,N_11212);
or U12436 (N_12436,N_11252,N_11021);
nor U12437 (N_12437,N_11311,N_11005);
nand U12438 (N_12438,N_11276,N_11321);
xor U12439 (N_12439,N_10955,N_11976);
xnor U12440 (N_12440,N_11882,N_11143);
nor U12441 (N_12441,N_11309,N_10957);
xor U12442 (N_12442,N_11100,N_11180);
and U12443 (N_12443,N_11139,N_11236);
or U12444 (N_12444,N_11530,N_11420);
and U12445 (N_12445,N_11153,N_11735);
or U12446 (N_12446,N_11213,N_11187);
or U12447 (N_12447,N_11701,N_11759);
nand U12448 (N_12448,N_11962,N_11806);
xor U12449 (N_12449,N_11349,N_11753);
nand U12450 (N_12450,N_11774,N_11817);
xor U12451 (N_12451,N_10943,N_11730);
nand U12452 (N_12452,N_11337,N_11058);
nor U12453 (N_12453,N_11489,N_11975);
xnor U12454 (N_12454,N_11588,N_11188);
or U12455 (N_12455,N_11794,N_11891);
nand U12456 (N_12456,N_11933,N_11569);
nor U12457 (N_12457,N_11233,N_11536);
nand U12458 (N_12458,N_11693,N_11022);
and U12459 (N_12459,N_11373,N_10972);
nor U12460 (N_12460,N_11646,N_11732);
or U12461 (N_12461,N_10800,N_11897);
nand U12462 (N_12462,N_11144,N_11150);
xnor U12463 (N_12463,N_11246,N_11200);
and U12464 (N_12464,N_10815,N_11784);
nand U12465 (N_12465,N_11392,N_10867);
xnor U12466 (N_12466,N_10894,N_10988);
and U12467 (N_12467,N_11287,N_11823);
xnor U12468 (N_12468,N_11636,N_11161);
nand U12469 (N_12469,N_11957,N_10837);
nor U12470 (N_12470,N_11750,N_11500);
nand U12471 (N_12471,N_10995,N_11329);
or U12472 (N_12472,N_11948,N_11167);
and U12473 (N_12473,N_10897,N_10844);
nor U12474 (N_12474,N_11564,N_10806);
or U12475 (N_12475,N_11340,N_11755);
and U12476 (N_12476,N_11089,N_11555);
and U12477 (N_12477,N_11994,N_11417);
nor U12478 (N_12478,N_10821,N_11253);
nand U12479 (N_12479,N_10958,N_11909);
nor U12480 (N_12480,N_11635,N_11808);
and U12481 (N_12481,N_11846,N_11871);
nor U12482 (N_12482,N_11032,N_11081);
nand U12483 (N_12483,N_11745,N_11042);
xnor U12484 (N_12484,N_11412,N_11576);
xnor U12485 (N_12485,N_11029,N_11747);
nor U12486 (N_12486,N_11037,N_11003);
nand U12487 (N_12487,N_11104,N_11726);
nor U12488 (N_12488,N_11080,N_11556);
xor U12489 (N_12489,N_10870,N_11733);
xor U12490 (N_12490,N_11856,N_11712);
nand U12491 (N_12491,N_11533,N_11777);
or U12492 (N_12492,N_10832,N_11162);
nor U12493 (N_12493,N_11890,N_11006);
and U12494 (N_12494,N_11969,N_11966);
nor U12495 (N_12495,N_11450,N_10856);
xnor U12496 (N_12496,N_11940,N_11985);
xor U12497 (N_12497,N_11086,N_11014);
and U12498 (N_12498,N_11698,N_11543);
nand U12499 (N_12499,N_11448,N_11654);
and U12500 (N_12500,N_10993,N_10980);
nand U12501 (N_12501,N_11980,N_11054);
xnor U12502 (N_12502,N_10951,N_11677);
and U12503 (N_12503,N_11799,N_11651);
or U12504 (N_12504,N_11388,N_11551);
xor U12505 (N_12505,N_11507,N_11939);
xor U12506 (N_12506,N_11419,N_11665);
and U12507 (N_12507,N_11892,N_11289);
xnor U12508 (N_12508,N_11428,N_11012);
xnor U12509 (N_12509,N_11354,N_11258);
nor U12510 (N_12510,N_11938,N_10939);
xnor U12511 (N_12511,N_11477,N_10892);
nand U12512 (N_12512,N_11136,N_11781);
or U12513 (N_12513,N_10986,N_11433);
nand U12514 (N_12514,N_11478,N_11027);
nor U12515 (N_12515,N_11660,N_11674);
xnor U12516 (N_12516,N_11867,N_10810);
and U12517 (N_12517,N_11396,N_11400);
nand U12518 (N_12518,N_11666,N_11620);
and U12519 (N_12519,N_10851,N_11627);
and U12520 (N_12520,N_11934,N_11714);
or U12521 (N_12521,N_10946,N_10914);
xor U12522 (N_12522,N_11872,N_11084);
xnor U12523 (N_12523,N_11602,N_11862);
nor U12524 (N_12524,N_11306,N_10855);
nor U12525 (N_12525,N_10919,N_11770);
or U12526 (N_12526,N_11087,N_11559);
and U12527 (N_12527,N_11532,N_11182);
or U12528 (N_12528,N_11545,N_11682);
nor U12529 (N_12529,N_10928,N_11789);
xnor U12530 (N_12530,N_11649,N_11622);
nand U12531 (N_12531,N_11766,N_10853);
xnor U12532 (N_12532,N_11013,N_11092);
nor U12533 (N_12533,N_10873,N_11163);
xnor U12534 (N_12534,N_11901,N_11483);
nand U12535 (N_12535,N_11435,N_11316);
or U12536 (N_12536,N_11822,N_11432);
or U12537 (N_12537,N_11604,N_11367);
xor U12538 (N_12538,N_11734,N_11978);
nand U12539 (N_12539,N_11603,N_11124);
or U12540 (N_12540,N_11768,N_11020);
nor U12541 (N_12541,N_11824,N_10884);
nor U12542 (N_12542,N_10843,N_11669);
nor U12543 (N_12543,N_11967,N_11641);
and U12544 (N_12544,N_10866,N_10847);
nor U12545 (N_12545,N_11474,N_10802);
or U12546 (N_12546,N_11691,N_11508);
nand U12547 (N_12547,N_11358,N_11548);
xor U12548 (N_12548,N_11018,N_11225);
and U12549 (N_12549,N_10956,N_11460);
or U12550 (N_12550,N_11740,N_11051);
xnor U12551 (N_12551,N_11809,N_11440);
or U12552 (N_12552,N_11685,N_11805);
and U12553 (N_12553,N_11181,N_11821);
nand U12554 (N_12554,N_11860,N_11709);
nor U12555 (N_12555,N_11997,N_11843);
nand U12556 (N_12556,N_11743,N_11011);
nor U12557 (N_12557,N_11248,N_11072);
nand U12558 (N_12558,N_11597,N_11126);
xnor U12559 (N_12559,N_10902,N_11366);
or U12560 (N_12560,N_11380,N_11461);
nor U12561 (N_12561,N_11408,N_11778);
nand U12562 (N_12562,N_11059,N_10989);
xnor U12563 (N_12563,N_11676,N_11264);
xnor U12564 (N_12564,N_11475,N_11300);
or U12565 (N_12565,N_11615,N_11526);
xor U12566 (N_12566,N_10982,N_11273);
nand U12567 (N_12567,N_11861,N_11261);
xnor U12568 (N_12568,N_11601,N_11447);
and U12569 (N_12569,N_11977,N_10953);
nand U12570 (N_12570,N_11519,N_11596);
or U12571 (N_12571,N_11361,N_11310);
and U12572 (N_12572,N_11097,N_11102);
xnor U12573 (N_12573,N_11249,N_11718);
and U12574 (N_12574,N_11859,N_11757);
xnor U12575 (N_12575,N_11547,N_11968);
or U12576 (N_12576,N_11196,N_11170);
nand U12577 (N_12577,N_11108,N_11179);
nand U12578 (N_12578,N_11357,N_11469);
and U12579 (N_12579,N_11129,N_11535);
nor U12580 (N_12580,N_11488,N_11887);
xor U12581 (N_12581,N_11192,N_11453);
nor U12582 (N_12582,N_11497,N_11214);
and U12583 (N_12583,N_11783,N_11422);
nor U12584 (N_12584,N_11544,N_11158);
xnor U12585 (N_12585,N_11302,N_10879);
nand U12586 (N_12586,N_11009,N_11098);
xnor U12587 (N_12587,N_11631,N_11607);
xor U12588 (N_12588,N_11290,N_10950);
and U12589 (N_12589,N_11888,N_11343);
xor U12590 (N_12590,N_11091,N_10966);
nand U12591 (N_12591,N_10805,N_11695);
nand U12592 (N_12592,N_11228,N_11319);
and U12593 (N_12593,N_11886,N_11910);
nand U12594 (N_12594,N_10819,N_11410);
and U12595 (N_12595,N_11360,N_11875);
nand U12596 (N_12596,N_11043,N_11906);
nor U12597 (N_12597,N_11147,N_11706);
and U12598 (N_12598,N_11652,N_10804);
and U12599 (N_12599,N_11686,N_11950);
xor U12600 (N_12600,N_11258,N_11955);
nor U12601 (N_12601,N_11400,N_11079);
or U12602 (N_12602,N_11408,N_10916);
and U12603 (N_12603,N_11529,N_11464);
nand U12604 (N_12604,N_11197,N_11196);
and U12605 (N_12605,N_11336,N_11339);
nand U12606 (N_12606,N_10988,N_11376);
or U12607 (N_12607,N_10850,N_10878);
or U12608 (N_12608,N_11172,N_11282);
nand U12609 (N_12609,N_10839,N_10869);
nor U12610 (N_12610,N_11954,N_11766);
and U12611 (N_12611,N_11502,N_11151);
and U12612 (N_12612,N_11144,N_11110);
or U12613 (N_12613,N_11957,N_11404);
or U12614 (N_12614,N_11668,N_11924);
and U12615 (N_12615,N_11020,N_11247);
and U12616 (N_12616,N_11113,N_10889);
xor U12617 (N_12617,N_11191,N_11901);
and U12618 (N_12618,N_11304,N_11857);
nand U12619 (N_12619,N_11049,N_10808);
and U12620 (N_12620,N_11106,N_11157);
and U12621 (N_12621,N_11395,N_11232);
and U12622 (N_12622,N_11044,N_11468);
and U12623 (N_12623,N_11266,N_10965);
or U12624 (N_12624,N_10942,N_11153);
nand U12625 (N_12625,N_11575,N_10801);
nand U12626 (N_12626,N_11798,N_11028);
and U12627 (N_12627,N_11587,N_11200);
xnor U12628 (N_12628,N_11741,N_11851);
and U12629 (N_12629,N_11080,N_11545);
and U12630 (N_12630,N_11394,N_11958);
or U12631 (N_12631,N_10914,N_11629);
and U12632 (N_12632,N_11591,N_11223);
nand U12633 (N_12633,N_11960,N_11704);
nor U12634 (N_12634,N_11868,N_11699);
nor U12635 (N_12635,N_11468,N_11959);
nand U12636 (N_12636,N_11546,N_11048);
and U12637 (N_12637,N_10870,N_11071);
nor U12638 (N_12638,N_11131,N_11297);
and U12639 (N_12639,N_11243,N_11203);
and U12640 (N_12640,N_11027,N_11259);
xnor U12641 (N_12641,N_11203,N_11849);
nor U12642 (N_12642,N_11235,N_10882);
nand U12643 (N_12643,N_11503,N_11297);
xnor U12644 (N_12644,N_10961,N_11412);
and U12645 (N_12645,N_11194,N_11741);
xor U12646 (N_12646,N_11611,N_11080);
or U12647 (N_12647,N_11443,N_11232);
and U12648 (N_12648,N_11055,N_10944);
xor U12649 (N_12649,N_11768,N_11872);
xor U12650 (N_12650,N_11105,N_11396);
nand U12651 (N_12651,N_11900,N_11295);
nor U12652 (N_12652,N_11940,N_10922);
xor U12653 (N_12653,N_11285,N_11090);
xor U12654 (N_12654,N_11343,N_11623);
nand U12655 (N_12655,N_10880,N_11385);
nor U12656 (N_12656,N_11137,N_10829);
or U12657 (N_12657,N_10919,N_11828);
xor U12658 (N_12658,N_11191,N_11397);
nor U12659 (N_12659,N_11902,N_11673);
xor U12660 (N_12660,N_10836,N_10808);
nor U12661 (N_12661,N_11613,N_11310);
nand U12662 (N_12662,N_11767,N_11691);
nand U12663 (N_12663,N_10926,N_11421);
nand U12664 (N_12664,N_11944,N_11306);
or U12665 (N_12665,N_11315,N_11615);
nor U12666 (N_12666,N_11121,N_11881);
and U12667 (N_12667,N_11864,N_10934);
nand U12668 (N_12668,N_11277,N_11263);
nor U12669 (N_12669,N_10874,N_11725);
and U12670 (N_12670,N_11925,N_11657);
and U12671 (N_12671,N_11406,N_11699);
xnor U12672 (N_12672,N_11269,N_11445);
xnor U12673 (N_12673,N_11738,N_11285);
and U12674 (N_12674,N_11172,N_11922);
or U12675 (N_12675,N_11272,N_11717);
and U12676 (N_12676,N_11057,N_11583);
or U12677 (N_12677,N_11334,N_11720);
or U12678 (N_12678,N_10807,N_11925);
and U12679 (N_12679,N_11949,N_11926);
nor U12680 (N_12680,N_11187,N_11126);
and U12681 (N_12681,N_10979,N_11141);
or U12682 (N_12682,N_11372,N_11424);
or U12683 (N_12683,N_11951,N_11544);
xnor U12684 (N_12684,N_11073,N_11686);
and U12685 (N_12685,N_11707,N_10976);
nand U12686 (N_12686,N_11260,N_11497);
or U12687 (N_12687,N_11866,N_10841);
or U12688 (N_12688,N_11897,N_11322);
nand U12689 (N_12689,N_11010,N_10879);
or U12690 (N_12690,N_11922,N_10805);
or U12691 (N_12691,N_11500,N_10916);
xnor U12692 (N_12692,N_10851,N_11032);
xnor U12693 (N_12693,N_11027,N_11335);
xor U12694 (N_12694,N_11469,N_11995);
and U12695 (N_12695,N_11115,N_11554);
nor U12696 (N_12696,N_11543,N_11221);
nor U12697 (N_12697,N_11089,N_11329);
and U12698 (N_12698,N_10836,N_11430);
nor U12699 (N_12699,N_11832,N_11213);
xnor U12700 (N_12700,N_11030,N_11345);
nand U12701 (N_12701,N_11863,N_11779);
nand U12702 (N_12702,N_11724,N_11968);
and U12703 (N_12703,N_10972,N_11419);
xnor U12704 (N_12704,N_10948,N_11404);
and U12705 (N_12705,N_11561,N_11031);
or U12706 (N_12706,N_11305,N_11101);
nand U12707 (N_12707,N_11930,N_10947);
nand U12708 (N_12708,N_11315,N_11322);
and U12709 (N_12709,N_10899,N_11499);
nor U12710 (N_12710,N_11186,N_11314);
nand U12711 (N_12711,N_11572,N_11926);
nor U12712 (N_12712,N_11518,N_11190);
nand U12713 (N_12713,N_11038,N_11274);
or U12714 (N_12714,N_10972,N_11429);
nand U12715 (N_12715,N_11537,N_11009);
or U12716 (N_12716,N_10868,N_11205);
and U12717 (N_12717,N_11480,N_11246);
nand U12718 (N_12718,N_10909,N_11862);
and U12719 (N_12719,N_11817,N_11882);
nand U12720 (N_12720,N_11002,N_11010);
and U12721 (N_12721,N_10888,N_11336);
and U12722 (N_12722,N_11797,N_11776);
nor U12723 (N_12723,N_11978,N_11943);
xnor U12724 (N_12724,N_11865,N_11909);
nand U12725 (N_12725,N_11212,N_11566);
or U12726 (N_12726,N_11174,N_11657);
nand U12727 (N_12727,N_11074,N_11393);
xnor U12728 (N_12728,N_11372,N_11455);
nor U12729 (N_12729,N_11057,N_11305);
nor U12730 (N_12730,N_11840,N_11408);
and U12731 (N_12731,N_11234,N_10824);
xnor U12732 (N_12732,N_11940,N_10870);
xnor U12733 (N_12733,N_10889,N_11866);
nand U12734 (N_12734,N_11863,N_10939);
nor U12735 (N_12735,N_11512,N_11141);
xor U12736 (N_12736,N_10825,N_10992);
nor U12737 (N_12737,N_11160,N_10814);
xor U12738 (N_12738,N_11344,N_11732);
nand U12739 (N_12739,N_10948,N_11364);
and U12740 (N_12740,N_10839,N_11949);
xnor U12741 (N_12741,N_11361,N_11153);
and U12742 (N_12742,N_10882,N_11090);
xor U12743 (N_12743,N_11788,N_11178);
or U12744 (N_12744,N_11627,N_11786);
xnor U12745 (N_12745,N_11593,N_10895);
nand U12746 (N_12746,N_11748,N_11302);
and U12747 (N_12747,N_11044,N_11505);
or U12748 (N_12748,N_11627,N_11529);
nand U12749 (N_12749,N_10928,N_11251);
or U12750 (N_12750,N_11291,N_11031);
nor U12751 (N_12751,N_11331,N_11067);
nand U12752 (N_12752,N_11798,N_11931);
and U12753 (N_12753,N_11611,N_11793);
and U12754 (N_12754,N_11809,N_11450);
xnor U12755 (N_12755,N_11086,N_10818);
xor U12756 (N_12756,N_11077,N_11026);
xor U12757 (N_12757,N_10939,N_11702);
xor U12758 (N_12758,N_11033,N_11010);
nor U12759 (N_12759,N_11030,N_11700);
and U12760 (N_12760,N_11179,N_11430);
and U12761 (N_12761,N_11620,N_11263);
xor U12762 (N_12762,N_10840,N_11094);
and U12763 (N_12763,N_11984,N_11495);
xnor U12764 (N_12764,N_11735,N_11373);
nor U12765 (N_12765,N_11060,N_10847);
nor U12766 (N_12766,N_11777,N_11409);
and U12767 (N_12767,N_11723,N_11258);
or U12768 (N_12768,N_11406,N_11447);
nand U12769 (N_12769,N_11528,N_11970);
and U12770 (N_12770,N_11461,N_11449);
or U12771 (N_12771,N_10829,N_11064);
nand U12772 (N_12772,N_11375,N_11917);
nor U12773 (N_12773,N_11247,N_11393);
or U12774 (N_12774,N_11869,N_11071);
nor U12775 (N_12775,N_11574,N_11293);
and U12776 (N_12776,N_11508,N_11214);
xor U12777 (N_12777,N_11208,N_11799);
nand U12778 (N_12778,N_11547,N_11755);
nor U12779 (N_12779,N_11017,N_11756);
xor U12780 (N_12780,N_11913,N_11601);
nor U12781 (N_12781,N_11489,N_11856);
nor U12782 (N_12782,N_10804,N_11186);
or U12783 (N_12783,N_10848,N_11573);
nand U12784 (N_12784,N_11078,N_11281);
and U12785 (N_12785,N_10865,N_11284);
and U12786 (N_12786,N_10961,N_11640);
or U12787 (N_12787,N_11192,N_11011);
nor U12788 (N_12788,N_11307,N_11947);
and U12789 (N_12789,N_10900,N_11431);
nor U12790 (N_12790,N_11349,N_11829);
and U12791 (N_12791,N_11981,N_11075);
or U12792 (N_12792,N_11630,N_11037);
nand U12793 (N_12793,N_11490,N_11963);
xor U12794 (N_12794,N_10901,N_11917);
or U12795 (N_12795,N_11391,N_11341);
nor U12796 (N_12796,N_11330,N_11570);
or U12797 (N_12797,N_11244,N_11451);
or U12798 (N_12798,N_11692,N_10922);
and U12799 (N_12799,N_11962,N_11618);
xor U12800 (N_12800,N_10905,N_11406);
nand U12801 (N_12801,N_11885,N_11679);
and U12802 (N_12802,N_11949,N_10814);
xor U12803 (N_12803,N_11959,N_11473);
nand U12804 (N_12804,N_11535,N_11481);
xor U12805 (N_12805,N_11431,N_11654);
xnor U12806 (N_12806,N_10990,N_10809);
nand U12807 (N_12807,N_11123,N_11567);
nor U12808 (N_12808,N_11240,N_11591);
xor U12809 (N_12809,N_11064,N_11884);
nor U12810 (N_12810,N_11386,N_11370);
and U12811 (N_12811,N_11079,N_11176);
xor U12812 (N_12812,N_11922,N_11650);
and U12813 (N_12813,N_11349,N_11192);
nand U12814 (N_12814,N_10828,N_11823);
nand U12815 (N_12815,N_11048,N_11298);
nand U12816 (N_12816,N_11193,N_11462);
nor U12817 (N_12817,N_11564,N_11165);
and U12818 (N_12818,N_11714,N_11183);
or U12819 (N_12819,N_11992,N_10880);
and U12820 (N_12820,N_11162,N_10941);
or U12821 (N_12821,N_11734,N_11224);
xor U12822 (N_12822,N_11724,N_10849);
or U12823 (N_12823,N_11792,N_11457);
and U12824 (N_12824,N_11016,N_11423);
nor U12825 (N_12825,N_11808,N_11871);
or U12826 (N_12826,N_11631,N_10951);
nor U12827 (N_12827,N_10971,N_11844);
nand U12828 (N_12828,N_11147,N_11163);
or U12829 (N_12829,N_10986,N_11046);
or U12830 (N_12830,N_11098,N_10854);
nand U12831 (N_12831,N_11349,N_11598);
nand U12832 (N_12832,N_11526,N_11370);
xor U12833 (N_12833,N_11894,N_11113);
and U12834 (N_12834,N_11504,N_11205);
or U12835 (N_12835,N_11536,N_10958);
nor U12836 (N_12836,N_11664,N_11481);
xor U12837 (N_12837,N_11155,N_11473);
xnor U12838 (N_12838,N_11258,N_11054);
and U12839 (N_12839,N_11583,N_11610);
and U12840 (N_12840,N_11406,N_11262);
xnor U12841 (N_12841,N_11270,N_11055);
nand U12842 (N_12842,N_11642,N_11753);
and U12843 (N_12843,N_11430,N_11038);
nand U12844 (N_12844,N_10964,N_11528);
xnor U12845 (N_12845,N_11291,N_11548);
or U12846 (N_12846,N_11759,N_11494);
xnor U12847 (N_12847,N_11235,N_10878);
nor U12848 (N_12848,N_10871,N_10815);
and U12849 (N_12849,N_10932,N_10801);
and U12850 (N_12850,N_11733,N_11904);
nand U12851 (N_12851,N_11923,N_11487);
and U12852 (N_12852,N_11311,N_11842);
or U12853 (N_12853,N_11988,N_11860);
or U12854 (N_12854,N_11724,N_11044);
and U12855 (N_12855,N_11430,N_10966);
xnor U12856 (N_12856,N_11003,N_11676);
and U12857 (N_12857,N_11390,N_11478);
nor U12858 (N_12858,N_11335,N_10816);
and U12859 (N_12859,N_11274,N_11205);
and U12860 (N_12860,N_11922,N_11709);
or U12861 (N_12861,N_11708,N_11497);
and U12862 (N_12862,N_10821,N_11529);
or U12863 (N_12863,N_10912,N_11115);
and U12864 (N_12864,N_11218,N_10954);
nand U12865 (N_12865,N_11189,N_11794);
and U12866 (N_12866,N_11284,N_11356);
xor U12867 (N_12867,N_11410,N_11203);
or U12868 (N_12868,N_11105,N_11016);
or U12869 (N_12869,N_11683,N_11194);
or U12870 (N_12870,N_11287,N_11118);
xnor U12871 (N_12871,N_11742,N_10911);
or U12872 (N_12872,N_11233,N_10957);
xnor U12873 (N_12873,N_11775,N_11068);
nand U12874 (N_12874,N_11936,N_11221);
and U12875 (N_12875,N_10829,N_10977);
and U12876 (N_12876,N_11555,N_11685);
nor U12877 (N_12877,N_11478,N_11816);
and U12878 (N_12878,N_11811,N_11474);
and U12879 (N_12879,N_11752,N_11123);
and U12880 (N_12880,N_11076,N_10838);
xnor U12881 (N_12881,N_11836,N_10812);
or U12882 (N_12882,N_11482,N_11625);
xnor U12883 (N_12883,N_11390,N_11530);
or U12884 (N_12884,N_11506,N_10898);
nor U12885 (N_12885,N_11415,N_11349);
xor U12886 (N_12886,N_11191,N_11567);
nor U12887 (N_12887,N_11119,N_11693);
xor U12888 (N_12888,N_11546,N_11729);
or U12889 (N_12889,N_11330,N_11405);
xnor U12890 (N_12890,N_11623,N_11302);
xnor U12891 (N_12891,N_10867,N_11539);
nor U12892 (N_12892,N_11600,N_10935);
and U12893 (N_12893,N_11855,N_11793);
or U12894 (N_12894,N_11129,N_11615);
nand U12895 (N_12895,N_10966,N_11086);
nand U12896 (N_12896,N_11121,N_11470);
nand U12897 (N_12897,N_11688,N_11427);
nor U12898 (N_12898,N_11400,N_10869);
nor U12899 (N_12899,N_11767,N_10835);
or U12900 (N_12900,N_11839,N_11341);
or U12901 (N_12901,N_10881,N_11964);
and U12902 (N_12902,N_10820,N_11135);
nor U12903 (N_12903,N_11241,N_11401);
nor U12904 (N_12904,N_11383,N_11925);
nand U12905 (N_12905,N_11015,N_11265);
and U12906 (N_12906,N_11497,N_11896);
nor U12907 (N_12907,N_11641,N_11248);
nor U12908 (N_12908,N_11255,N_11561);
nor U12909 (N_12909,N_11268,N_11430);
nor U12910 (N_12910,N_11259,N_11545);
or U12911 (N_12911,N_11141,N_10876);
and U12912 (N_12912,N_11164,N_11641);
xnor U12913 (N_12913,N_11987,N_11407);
xor U12914 (N_12914,N_11475,N_11611);
and U12915 (N_12915,N_11505,N_11231);
nor U12916 (N_12916,N_10808,N_11348);
or U12917 (N_12917,N_11420,N_11471);
xor U12918 (N_12918,N_11069,N_11210);
xnor U12919 (N_12919,N_11937,N_11482);
or U12920 (N_12920,N_10980,N_11439);
nor U12921 (N_12921,N_11363,N_11216);
and U12922 (N_12922,N_11308,N_11247);
xor U12923 (N_12923,N_11222,N_11722);
nor U12924 (N_12924,N_11108,N_10859);
and U12925 (N_12925,N_10830,N_11911);
nand U12926 (N_12926,N_11000,N_11590);
nor U12927 (N_12927,N_11658,N_11727);
nor U12928 (N_12928,N_11834,N_10972);
nor U12929 (N_12929,N_11875,N_11992);
nand U12930 (N_12930,N_11113,N_11135);
nand U12931 (N_12931,N_11778,N_11610);
and U12932 (N_12932,N_11730,N_11412);
and U12933 (N_12933,N_10952,N_10921);
xnor U12934 (N_12934,N_11942,N_11974);
xor U12935 (N_12935,N_11704,N_11773);
nand U12936 (N_12936,N_11356,N_11879);
or U12937 (N_12937,N_10967,N_11199);
or U12938 (N_12938,N_11889,N_10836);
and U12939 (N_12939,N_10921,N_11700);
and U12940 (N_12940,N_11876,N_10896);
or U12941 (N_12941,N_11178,N_11471);
and U12942 (N_12942,N_11011,N_11036);
nor U12943 (N_12943,N_11755,N_11771);
xor U12944 (N_12944,N_10874,N_11772);
and U12945 (N_12945,N_11524,N_11534);
and U12946 (N_12946,N_11040,N_11854);
nor U12947 (N_12947,N_11911,N_11621);
xnor U12948 (N_12948,N_11649,N_11189);
xor U12949 (N_12949,N_11738,N_11066);
xor U12950 (N_12950,N_11606,N_10814);
nor U12951 (N_12951,N_11905,N_11625);
xnor U12952 (N_12952,N_10866,N_10917);
or U12953 (N_12953,N_11062,N_11334);
nand U12954 (N_12954,N_10932,N_11085);
nand U12955 (N_12955,N_11141,N_11211);
and U12956 (N_12956,N_11766,N_11175);
nand U12957 (N_12957,N_11490,N_11836);
or U12958 (N_12958,N_11703,N_11898);
nor U12959 (N_12959,N_11713,N_10936);
and U12960 (N_12960,N_11560,N_11392);
nor U12961 (N_12961,N_11627,N_11788);
or U12962 (N_12962,N_11965,N_11216);
or U12963 (N_12963,N_11378,N_11703);
nand U12964 (N_12964,N_11412,N_11347);
xor U12965 (N_12965,N_11850,N_11861);
and U12966 (N_12966,N_11470,N_11789);
nand U12967 (N_12967,N_11283,N_11960);
nand U12968 (N_12968,N_11394,N_11640);
and U12969 (N_12969,N_11836,N_11240);
or U12970 (N_12970,N_11628,N_10958);
nor U12971 (N_12971,N_10852,N_11346);
or U12972 (N_12972,N_11412,N_11369);
or U12973 (N_12973,N_11893,N_11420);
and U12974 (N_12974,N_11531,N_11128);
xor U12975 (N_12975,N_10804,N_10814);
xnor U12976 (N_12976,N_11896,N_11647);
xnor U12977 (N_12977,N_11879,N_11830);
xnor U12978 (N_12978,N_11694,N_11600);
nor U12979 (N_12979,N_11631,N_10933);
or U12980 (N_12980,N_11156,N_11139);
xnor U12981 (N_12981,N_11911,N_10825);
nand U12982 (N_12982,N_11181,N_10849);
nand U12983 (N_12983,N_10945,N_11933);
xor U12984 (N_12984,N_11320,N_11091);
nand U12985 (N_12985,N_11967,N_10881);
or U12986 (N_12986,N_11079,N_10865);
xor U12987 (N_12987,N_11179,N_11742);
and U12988 (N_12988,N_11708,N_11634);
nor U12989 (N_12989,N_11203,N_11912);
xnor U12990 (N_12990,N_11811,N_11129);
xor U12991 (N_12991,N_11850,N_11923);
nand U12992 (N_12992,N_10810,N_11874);
or U12993 (N_12993,N_11765,N_11115);
or U12994 (N_12994,N_11168,N_11335);
or U12995 (N_12995,N_11987,N_11415);
nand U12996 (N_12996,N_11463,N_11624);
and U12997 (N_12997,N_11193,N_11082);
and U12998 (N_12998,N_11556,N_11502);
nand U12999 (N_12999,N_11384,N_11492);
xnor U13000 (N_13000,N_11443,N_11894);
nor U13001 (N_13001,N_11508,N_11433);
and U13002 (N_13002,N_11642,N_11933);
nor U13003 (N_13003,N_11708,N_11399);
and U13004 (N_13004,N_11079,N_11239);
or U13005 (N_13005,N_11615,N_11575);
nand U13006 (N_13006,N_11154,N_11132);
nand U13007 (N_13007,N_11401,N_11062);
nor U13008 (N_13008,N_10896,N_11124);
xnor U13009 (N_13009,N_11215,N_11971);
and U13010 (N_13010,N_11190,N_11412);
nand U13011 (N_13011,N_11349,N_11088);
xor U13012 (N_13012,N_10983,N_11857);
or U13013 (N_13013,N_11917,N_11946);
nand U13014 (N_13014,N_11995,N_10833);
or U13015 (N_13015,N_11091,N_11540);
nand U13016 (N_13016,N_11261,N_11013);
and U13017 (N_13017,N_11468,N_11484);
and U13018 (N_13018,N_11519,N_11937);
xnor U13019 (N_13019,N_10853,N_11136);
nand U13020 (N_13020,N_11670,N_10985);
nand U13021 (N_13021,N_11119,N_11092);
xnor U13022 (N_13022,N_11584,N_10825);
nor U13023 (N_13023,N_11810,N_11222);
xor U13024 (N_13024,N_11331,N_10987);
nand U13025 (N_13025,N_11869,N_11345);
and U13026 (N_13026,N_10844,N_11311);
and U13027 (N_13027,N_11508,N_11284);
xnor U13028 (N_13028,N_11301,N_10975);
or U13029 (N_13029,N_11098,N_11486);
xor U13030 (N_13030,N_11957,N_11962);
nor U13031 (N_13031,N_11640,N_11426);
xnor U13032 (N_13032,N_11161,N_11318);
and U13033 (N_13033,N_11184,N_11469);
xor U13034 (N_13034,N_11080,N_11886);
nand U13035 (N_13035,N_11946,N_11009);
xor U13036 (N_13036,N_10806,N_11683);
xnor U13037 (N_13037,N_11042,N_11748);
nor U13038 (N_13038,N_11837,N_11322);
nand U13039 (N_13039,N_11684,N_11433);
and U13040 (N_13040,N_11300,N_11262);
and U13041 (N_13041,N_10899,N_11549);
and U13042 (N_13042,N_11649,N_11360);
xnor U13043 (N_13043,N_11660,N_11603);
or U13044 (N_13044,N_11082,N_11501);
nand U13045 (N_13045,N_10930,N_10889);
or U13046 (N_13046,N_11849,N_11196);
or U13047 (N_13047,N_11325,N_11844);
xor U13048 (N_13048,N_10808,N_11373);
nand U13049 (N_13049,N_11144,N_11062);
xor U13050 (N_13050,N_10847,N_11093);
nand U13051 (N_13051,N_11134,N_10823);
nand U13052 (N_13052,N_10993,N_11747);
xnor U13053 (N_13053,N_11276,N_11121);
nand U13054 (N_13054,N_11376,N_10940);
and U13055 (N_13055,N_11981,N_11442);
nor U13056 (N_13056,N_11390,N_11041);
nand U13057 (N_13057,N_11543,N_11103);
xor U13058 (N_13058,N_10873,N_11558);
and U13059 (N_13059,N_11091,N_11746);
or U13060 (N_13060,N_11777,N_11473);
xor U13061 (N_13061,N_11406,N_10890);
nand U13062 (N_13062,N_11873,N_11763);
nand U13063 (N_13063,N_10851,N_10824);
xor U13064 (N_13064,N_10822,N_11708);
nand U13065 (N_13065,N_11699,N_10816);
and U13066 (N_13066,N_11162,N_11592);
nand U13067 (N_13067,N_10995,N_11046);
xnor U13068 (N_13068,N_11097,N_11750);
and U13069 (N_13069,N_11040,N_11976);
or U13070 (N_13070,N_11919,N_11228);
or U13071 (N_13071,N_11631,N_11516);
or U13072 (N_13072,N_11634,N_11090);
nor U13073 (N_13073,N_11292,N_11755);
or U13074 (N_13074,N_11556,N_11990);
nor U13075 (N_13075,N_11447,N_11817);
and U13076 (N_13076,N_11479,N_11083);
nor U13077 (N_13077,N_11489,N_10946);
or U13078 (N_13078,N_11782,N_11132);
nand U13079 (N_13079,N_11345,N_11885);
nor U13080 (N_13080,N_11319,N_11162);
and U13081 (N_13081,N_11882,N_10947);
nand U13082 (N_13082,N_10843,N_11986);
or U13083 (N_13083,N_11060,N_11790);
and U13084 (N_13084,N_11463,N_11391);
xnor U13085 (N_13085,N_11606,N_11077);
nand U13086 (N_13086,N_11779,N_11887);
or U13087 (N_13087,N_11491,N_10950);
nor U13088 (N_13088,N_11958,N_11991);
nand U13089 (N_13089,N_10897,N_10824);
or U13090 (N_13090,N_11183,N_10905);
xor U13091 (N_13091,N_11713,N_11123);
xnor U13092 (N_13092,N_11473,N_11644);
nor U13093 (N_13093,N_11575,N_11399);
xor U13094 (N_13094,N_10862,N_11883);
and U13095 (N_13095,N_11027,N_11441);
nand U13096 (N_13096,N_11204,N_11329);
nor U13097 (N_13097,N_11737,N_11689);
xnor U13098 (N_13098,N_11026,N_10896);
or U13099 (N_13099,N_10846,N_10838);
nand U13100 (N_13100,N_11132,N_11675);
xor U13101 (N_13101,N_11685,N_11500);
or U13102 (N_13102,N_11383,N_11977);
and U13103 (N_13103,N_11993,N_11896);
nor U13104 (N_13104,N_10814,N_11076);
nor U13105 (N_13105,N_11250,N_11685);
nor U13106 (N_13106,N_11581,N_11915);
xnor U13107 (N_13107,N_11985,N_11704);
and U13108 (N_13108,N_10993,N_11790);
and U13109 (N_13109,N_11966,N_11193);
nand U13110 (N_13110,N_10885,N_10862);
and U13111 (N_13111,N_11675,N_11289);
xor U13112 (N_13112,N_11368,N_11073);
or U13113 (N_13113,N_11592,N_11200);
and U13114 (N_13114,N_11946,N_11820);
and U13115 (N_13115,N_11541,N_11807);
and U13116 (N_13116,N_11544,N_11349);
or U13117 (N_13117,N_11794,N_11021);
and U13118 (N_13118,N_11995,N_11395);
or U13119 (N_13119,N_11882,N_11186);
nand U13120 (N_13120,N_11357,N_11901);
or U13121 (N_13121,N_11525,N_11475);
or U13122 (N_13122,N_11662,N_11234);
or U13123 (N_13123,N_11100,N_11050);
xnor U13124 (N_13124,N_11497,N_11937);
and U13125 (N_13125,N_11418,N_11004);
or U13126 (N_13126,N_11598,N_11425);
or U13127 (N_13127,N_11358,N_11603);
xor U13128 (N_13128,N_11921,N_11574);
and U13129 (N_13129,N_11385,N_11571);
or U13130 (N_13130,N_11041,N_11394);
or U13131 (N_13131,N_11026,N_11431);
xor U13132 (N_13132,N_11455,N_10876);
or U13133 (N_13133,N_11198,N_11262);
nand U13134 (N_13134,N_10806,N_11244);
xor U13135 (N_13135,N_11914,N_10884);
xnor U13136 (N_13136,N_11062,N_10971);
nor U13137 (N_13137,N_11677,N_10883);
nand U13138 (N_13138,N_11836,N_11237);
nor U13139 (N_13139,N_11248,N_11954);
xnor U13140 (N_13140,N_10929,N_11684);
or U13141 (N_13141,N_10845,N_11596);
or U13142 (N_13142,N_11289,N_11595);
and U13143 (N_13143,N_10832,N_11567);
nand U13144 (N_13144,N_11679,N_11690);
nor U13145 (N_13145,N_11553,N_11208);
and U13146 (N_13146,N_11958,N_11948);
xnor U13147 (N_13147,N_11835,N_11359);
nand U13148 (N_13148,N_11674,N_11507);
or U13149 (N_13149,N_11605,N_11761);
nand U13150 (N_13150,N_11971,N_11266);
nor U13151 (N_13151,N_11946,N_11734);
nand U13152 (N_13152,N_10860,N_11246);
or U13153 (N_13153,N_11526,N_11574);
nand U13154 (N_13154,N_11054,N_11373);
nand U13155 (N_13155,N_11013,N_10908);
and U13156 (N_13156,N_11098,N_10990);
and U13157 (N_13157,N_11817,N_11518);
xor U13158 (N_13158,N_10823,N_10986);
or U13159 (N_13159,N_11027,N_11876);
nand U13160 (N_13160,N_11469,N_11453);
xor U13161 (N_13161,N_10973,N_11785);
xor U13162 (N_13162,N_10947,N_10932);
xor U13163 (N_13163,N_10882,N_11279);
nor U13164 (N_13164,N_11044,N_11767);
and U13165 (N_13165,N_11478,N_11760);
nor U13166 (N_13166,N_10866,N_11120);
or U13167 (N_13167,N_11678,N_11929);
nor U13168 (N_13168,N_11227,N_11005);
or U13169 (N_13169,N_11844,N_11775);
xor U13170 (N_13170,N_11769,N_11157);
or U13171 (N_13171,N_11246,N_11403);
xor U13172 (N_13172,N_11273,N_11409);
or U13173 (N_13173,N_11710,N_11660);
xor U13174 (N_13174,N_11741,N_11358);
and U13175 (N_13175,N_11165,N_11510);
or U13176 (N_13176,N_10879,N_11844);
and U13177 (N_13177,N_11161,N_11774);
xor U13178 (N_13178,N_11904,N_11947);
or U13179 (N_13179,N_11436,N_11925);
xnor U13180 (N_13180,N_11377,N_11290);
and U13181 (N_13181,N_10804,N_11415);
and U13182 (N_13182,N_11431,N_11106);
nand U13183 (N_13183,N_11821,N_11127);
nor U13184 (N_13184,N_11255,N_11765);
nor U13185 (N_13185,N_11980,N_11951);
xnor U13186 (N_13186,N_11586,N_11114);
or U13187 (N_13187,N_10960,N_11907);
nor U13188 (N_13188,N_11947,N_11299);
xor U13189 (N_13189,N_11660,N_11447);
xor U13190 (N_13190,N_11602,N_11592);
or U13191 (N_13191,N_11070,N_11959);
or U13192 (N_13192,N_10928,N_11471);
and U13193 (N_13193,N_11397,N_10989);
or U13194 (N_13194,N_10825,N_11826);
xor U13195 (N_13195,N_11158,N_11440);
and U13196 (N_13196,N_11948,N_11115);
or U13197 (N_13197,N_11197,N_11828);
or U13198 (N_13198,N_11532,N_11814);
and U13199 (N_13199,N_11671,N_10987);
xor U13200 (N_13200,N_12666,N_12733);
and U13201 (N_13201,N_12320,N_12986);
nor U13202 (N_13202,N_12084,N_12579);
and U13203 (N_13203,N_12214,N_13197);
and U13204 (N_13204,N_12585,N_12086);
nand U13205 (N_13205,N_12736,N_12246);
and U13206 (N_13206,N_12847,N_12791);
nand U13207 (N_13207,N_12704,N_12687);
xor U13208 (N_13208,N_12096,N_12574);
nor U13209 (N_13209,N_12296,N_13164);
nor U13210 (N_13210,N_12748,N_12248);
nand U13211 (N_13211,N_12104,N_12247);
xnor U13212 (N_13212,N_13111,N_12173);
nor U13213 (N_13213,N_12934,N_12827);
nand U13214 (N_13214,N_12971,N_12257);
and U13215 (N_13215,N_12695,N_12450);
xnor U13216 (N_13216,N_12019,N_12680);
xor U13217 (N_13217,N_12905,N_12156);
nor U13218 (N_13218,N_12809,N_12872);
nor U13219 (N_13219,N_12756,N_12618);
and U13220 (N_13220,N_12366,N_12122);
and U13221 (N_13221,N_12755,N_12874);
nor U13222 (N_13222,N_12647,N_12497);
and U13223 (N_13223,N_12002,N_13057);
and U13224 (N_13224,N_13150,N_12235);
nor U13225 (N_13225,N_13098,N_12272);
nor U13226 (N_13226,N_12642,N_12726);
xor U13227 (N_13227,N_12991,N_12951);
and U13228 (N_13228,N_12038,N_12340);
nand U13229 (N_13229,N_13025,N_12598);
xor U13230 (N_13230,N_12977,N_12492);
and U13231 (N_13231,N_12500,N_12111);
nor U13232 (N_13232,N_12932,N_12651);
nor U13233 (N_13233,N_12863,N_12969);
nor U13234 (N_13234,N_12379,N_12152);
nand U13235 (N_13235,N_12982,N_13076);
xor U13236 (N_13236,N_13060,N_12107);
and U13237 (N_13237,N_12395,N_12443);
nand U13238 (N_13238,N_12974,N_12179);
nand U13239 (N_13239,N_12390,N_12828);
nor U13240 (N_13240,N_12790,N_12669);
or U13241 (N_13241,N_12775,N_12461);
nor U13242 (N_13242,N_12779,N_12685);
or U13243 (N_13243,N_12478,N_12462);
or U13244 (N_13244,N_12141,N_12402);
or U13245 (N_13245,N_12040,N_12885);
or U13246 (N_13246,N_13126,N_12313);
or U13247 (N_13247,N_12297,N_12533);
nor U13248 (N_13248,N_12020,N_12530);
and U13249 (N_13249,N_12489,N_13162);
nor U13250 (N_13250,N_13037,N_12523);
nor U13251 (N_13251,N_12621,N_12614);
xor U13252 (N_13252,N_12644,N_12865);
or U13253 (N_13253,N_12149,N_13066);
or U13254 (N_13254,N_12336,N_12090);
nand U13255 (N_13255,N_12317,N_12232);
nor U13256 (N_13256,N_12041,N_12854);
nor U13257 (N_13257,N_12023,N_13038);
nand U13258 (N_13258,N_12590,N_12761);
and U13259 (N_13259,N_13032,N_12507);
and U13260 (N_13260,N_12311,N_13187);
nand U13261 (N_13261,N_12147,N_12697);
nor U13262 (N_13262,N_12267,N_12278);
nor U13263 (N_13263,N_12605,N_12841);
xor U13264 (N_13264,N_12565,N_12945);
xor U13265 (N_13265,N_12251,N_12085);
and U13266 (N_13266,N_12337,N_13017);
and U13267 (N_13267,N_12470,N_12781);
nand U13268 (N_13268,N_12675,N_12958);
or U13269 (N_13269,N_12563,N_13147);
nor U13270 (N_13270,N_12004,N_12606);
nor U13271 (N_13271,N_12586,N_12712);
or U13272 (N_13272,N_13129,N_12617);
and U13273 (N_13273,N_12539,N_12205);
or U13274 (N_13274,N_12894,N_12202);
nor U13275 (N_13275,N_12245,N_12783);
and U13276 (N_13276,N_12562,N_12315);
nor U13277 (N_13277,N_12108,N_12200);
nand U13278 (N_13278,N_12576,N_13152);
and U13279 (N_13279,N_12482,N_12098);
xor U13280 (N_13280,N_13042,N_13026);
or U13281 (N_13281,N_13118,N_12966);
xor U13282 (N_13282,N_12520,N_13014);
nor U13283 (N_13283,N_12377,N_12913);
nor U13284 (N_13284,N_12476,N_13106);
and U13285 (N_13285,N_12678,N_12433);
xnor U13286 (N_13286,N_12030,N_13123);
or U13287 (N_13287,N_12125,N_12400);
nor U13288 (N_13288,N_12677,N_12062);
and U13289 (N_13289,N_12404,N_12509);
and U13290 (N_13290,N_13097,N_12029);
xnor U13291 (N_13291,N_12498,N_13137);
xor U13292 (N_13292,N_13143,N_12887);
nand U13293 (N_13293,N_12972,N_13193);
or U13294 (N_13294,N_12412,N_12198);
nand U13295 (N_13295,N_12649,N_12438);
and U13296 (N_13296,N_12472,N_12195);
or U13297 (N_13297,N_12143,N_12948);
nand U13298 (N_13298,N_12375,N_12082);
or U13299 (N_13299,N_12480,N_12962);
nor U13300 (N_13300,N_12166,N_12488);
nor U13301 (N_13301,N_12324,N_12508);
xnor U13302 (N_13302,N_12429,N_12778);
nand U13303 (N_13303,N_12998,N_12672);
or U13304 (N_13304,N_13086,N_12229);
xor U13305 (N_13305,N_12486,N_13179);
nand U13306 (N_13306,N_12128,N_13101);
and U13307 (N_13307,N_12116,N_12811);
and U13308 (N_13308,N_12866,N_12852);
or U13309 (N_13309,N_12832,N_12446);
nor U13310 (N_13310,N_12210,N_13074);
nand U13311 (N_13311,N_12342,N_12407);
nor U13312 (N_13312,N_12061,N_12236);
xor U13313 (N_13313,N_13173,N_12683);
nand U13314 (N_13314,N_12178,N_12580);
or U13315 (N_13315,N_12378,N_13168);
nor U13316 (N_13316,N_12220,N_13140);
nor U13317 (N_13317,N_12593,N_13044);
or U13318 (N_13318,N_12941,N_13093);
xor U13319 (N_13319,N_13139,N_12559);
and U13320 (N_13320,N_12522,N_12435);
nor U13321 (N_13321,N_13083,N_12109);
nand U13322 (N_13322,N_12224,N_12723);
and U13323 (N_13323,N_12701,N_12754);
and U13324 (N_13324,N_12535,N_12284);
xor U13325 (N_13325,N_12900,N_12949);
and U13326 (N_13326,N_12646,N_12601);
nand U13327 (N_13327,N_12158,N_12469);
nand U13328 (N_13328,N_12737,N_12273);
or U13329 (N_13329,N_12912,N_12279);
and U13330 (N_13330,N_12308,N_12613);
or U13331 (N_13331,N_12066,N_12627);
xor U13332 (N_13332,N_13069,N_12549);
xor U13333 (N_13333,N_12380,N_12068);
nor U13334 (N_13334,N_13102,N_12430);
xnor U13335 (N_13335,N_12421,N_12713);
nand U13336 (N_13336,N_12921,N_12801);
nand U13337 (N_13337,N_13163,N_12184);
nor U13338 (N_13338,N_12581,N_12557);
and U13339 (N_13339,N_12459,N_12304);
nor U13340 (N_13340,N_12561,N_13018);
xor U13341 (N_13341,N_12275,N_12506);
or U13342 (N_13342,N_12793,N_12639);
nor U13343 (N_13343,N_12097,N_12487);
nand U13344 (N_13344,N_12322,N_12786);
nand U13345 (N_13345,N_12410,N_12334);
and U13346 (N_13346,N_12578,N_12177);
xnor U13347 (N_13347,N_12861,N_13020);
nand U13348 (N_13348,N_12194,N_12431);
nand U13349 (N_13349,N_13136,N_13009);
nor U13350 (N_13350,N_12751,N_12025);
nor U13351 (N_13351,N_13181,N_13186);
and U13352 (N_13352,N_13189,N_12927);
nand U13353 (N_13353,N_13192,N_12458);
xor U13354 (N_13354,N_12667,N_12138);
or U13355 (N_13355,N_12261,N_12001);
nor U13356 (N_13356,N_12961,N_12519);
nand U13357 (N_13357,N_12353,N_12815);
xor U13358 (N_13358,N_13119,N_12831);
xor U13359 (N_13359,N_12069,N_13030);
nand U13360 (N_13360,N_12049,N_12764);
or U13361 (N_13361,N_12770,N_12075);
or U13362 (N_13362,N_12588,N_12645);
or U13363 (N_13363,N_12853,N_13115);
xnor U13364 (N_13364,N_12848,N_12219);
or U13365 (N_13365,N_12804,N_13013);
nand U13366 (N_13366,N_12978,N_12993);
or U13367 (N_13367,N_12189,N_12452);
nor U13368 (N_13368,N_12720,N_12243);
nand U13369 (N_13369,N_12682,N_12239);
nor U13370 (N_13370,N_12244,N_12483);
and U13371 (N_13371,N_12341,N_12759);
and U13372 (N_13372,N_12065,N_12323);
xor U13373 (N_13373,N_12213,N_12042);
nand U13374 (N_13374,N_13003,N_12873);
and U13375 (N_13375,N_12270,N_13155);
xnor U13376 (N_13376,N_12413,N_12940);
or U13377 (N_13377,N_12923,N_12017);
and U13378 (N_13378,N_12216,N_13134);
xor U13379 (N_13379,N_13114,N_12591);
nand U13380 (N_13380,N_12953,N_12782);
and U13381 (N_13381,N_12406,N_13156);
or U13382 (N_13382,N_12052,N_12369);
and U13383 (N_13383,N_12491,N_13148);
and U13384 (N_13384,N_12330,N_12131);
nand U13385 (N_13385,N_12602,N_12384);
xor U13386 (N_13386,N_12454,N_12348);
and U13387 (N_13387,N_12571,N_12551);
or U13388 (N_13388,N_12298,N_12037);
nand U13389 (N_13389,N_13177,N_12199);
and U13390 (N_13390,N_13127,N_12329);
or U13391 (N_13391,N_13068,N_12548);
and U13392 (N_13392,N_12876,N_13064);
or U13393 (N_13393,N_13169,N_12240);
and U13394 (N_13394,N_12925,N_12439);
or U13395 (N_13395,N_12481,N_12150);
xnor U13396 (N_13396,N_12997,N_13006);
nand U13397 (N_13397,N_12203,N_12599);
and U13398 (N_13398,N_12662,N_12884);
and U13399 (N_13399,N_12118,N_13167);
xor U13400 (N_13400,N_12027,N_12850);
or U13401 (N_13401,N_12475,N_12631);
and U13402 (N_13402,N_13048,N_13157);
or U13403 (N_13403,N_12079,N_12931);
xor U13404 (N_13404,N_12741,N_12758);
nor U13405 (N_13405,N_12544,N_12453);
xnor U13406 (N_13406,N_12295,N_12165);
xor U13407 (N_13407,N_12493,N_12302);
or U13408 (N_13408,N_12449,N_12021);
nor U13409 (N_13409,N_12399,N_12473);
xnor U13410 (N_13410,N_12608,N_12699);
xnor U13411 (N_13411,N_13055,N_12162);
or U13412 (N_13412,N_12309,N_13029);
nand U13413 (N_13413,N_12636,N_12738);
or U13414 (N_13414,N_13180,N_13121);
nor U13415 (N_13415,N_13109,N_12992);
nor U13416 (N_13416,N_12350,N_13063);
xnor U13417 (N_13417,N_12813,N_12707);
and U13418 (N_13418,N_12538,N_12996);
xnor U13419 (N_13419,N_12554,N_12879);
xor U13420 (N_13420,N_13034,N_12694);
nor U13421 (N_13421,N_12271,N_12359);
nand U13422 (N_13422,N_12420,N_12505);
or U13423 (N_13423,N_12423,N_12164);
nor U13424 (N_13424,N_12231,N_12929);
and U13425 (N_13425,N_12665,N_12318);
or U13426 (N_13426,N_13149,N_12663);
and U13427 (N_13427,N_13135,N_12233);
or U13428 (N_13428,N_12316,N_12467);
xnor U13429 (N_13429,N_12319,N_12514);
and U13430 (N_13430,N_12526,N_12656);
or U13431 (N_13431,N_12881,N_12875);
nor U13432 (N_13432,N_13094,N_12135);
xnor U13433 (N_13433,N_12388,N_13062);
nand U13434 (N_13434,N_12772,N_12566);
or U13435 (N_13435,N_12451,N_12227);
nand U13436 (N_13436,N_12136,N_13122);
and U13437 (N_13437,N_13012,N_12005);
nand U13438 (N_13438,N_12944,N_12626);
nand U13439 (N_13439,N_12600,N_13005);
nor U13440 (N_13440,N_12836,N_13046);
nand U13441 (N_13441,N_12902,N_12312);
and U13442 (N_13442,N_12363,N_12047);
xnor U13443 (N_13443,N_13056,N_12840);
nand U13444 (N_13444,N_12915,N_12950);
xnor U13445 (N_13445,N_12387,N_12742);
nand U13446 (N_13446,N_12930,N_12133);
nor U13447 (N_13447,N_12589,N_12364);
nor U13448 (N_13448,N_12101,N_12365);
or U13449 (N_13449,N_12440,N_12587);
and U13450 (N_13450,N_12174,N_12124);
xor U13451 (N_13451,N_12422,N_12358);
or U13452 (N_13452,N_13041,N_13050);
nor U13453 (N_13453,N_12425,N_12277);
nand U13454 (N_13454,N_12238,N_12067);
nand U13455 (N_13455,N_12305,N_13166);
xor U13456 (N_13456,N_12528,N_12797);
nor U13457 (N_13457,N_13031,N_12735);
nor U13458 (N_13458,N_12054,N_12749);
or U13459 (N_13459,N_12620,N_12258);
xor U13460 (N_13460,N_12140,N_12632);
nor U13461 (N_13461,N_12218,N_12835);
xor U13462 (N_13462,N_12294,N_13124);
nand U13463 (N_13463,N_13151,N_12946);
nor U13464 (N_13464,N_12008,N_13184);
xor U13465 (N_13465,N_12844,N_12686);
nand U13466 (N_13466,N_12269,N_13052);
and U13467 (N_13467,N_12223,N_12990);
and U13468 (N_13468,N_12968,N_12477);
xor U13469 (N_13469,N_12648,N_12743);
nand U13470 (N_13470,N_12664,N_12250);
or U13471 (N_13471,N_12468,N_12081);
or U13472 (N_13472,N_12970,N_12910);
nor U13473 (N_13473,N_13084,N_13195);
xor U13474 (N_13474,N_13183,N_12356);
nor U13475 (N_13475,N_12083,N_12711);
nor U13476 (N_13476,N_12728,N_12256);
and U13477 (N_13477,N_12221,N_12120);
and U13478 (N_13478,N_12112,N_12092);
xor U13479 (N_13479,N_12033,N_13082);
xnor U13480 (N_13480,N_12820,N_13144);
or U13481 (N_13481,N_12362,N_12954);
or U13482 (N_13482,N_13002,N_12655);
and U13483 (N_13483,N_12003,N_12918);
xnor U13484 (N_13484,N_12592,N_12012);
xor U13485 (N_13485,N_13045,N_12878);
xor U13486 (N_13486,N_12121,N_12570);
or U13487 (N_13487,N_12939,N_12842);
and U13488 (N_13488,N_12466,N_12288);
xnor U13489 (N_13489,N_13185,N_12331);
xnor U13490 (N_13490,N_12710,N_13194);
nor U13491 (N_13491,N_12994,N_13175);
xor U13492 (N_13492,N_12051,N_12792);
nand U13493 (N_13493,N_12151,N_12088);
nand U13494 (N_13494,N_12398,N_12619);
and U13495 (N_13495,N_13072,N_12928);
or U13496 (N_13496,N_12328,N_12237);
xor U13497 (N_13497,N_12280,N_12688);
xor U13498 (N_13498,N_13142,N_12834);
xnor U13499 (N_13499,N_12070,N_13079);
and U13500 (N_13500,N_12628,N_12386);
or U13501 (N_13501,N_12916,N_12583);
nor U13502 (N_13502,N_13059,N_12769);
nand U13503 (N_13503,N_12106,N_12965);
nand U13504 (N_13504,N_12914,N_12572);
xor U13505 (N_13505,N_12569,N_12973);
nand U13506 (N_13506,N_12846,N_12689);
nor U13507 (N_13507,N_13035,N_12015);
nand U13508 (N_13508,N_12609,N_13125);
or U13509 (N_13509,N_13176,N_12260);
and U13510 (N_13510,N_12394,N_12830);
nor U13511 (N_13511,N_12490,N_12408);
nand U13512 (N_13512,N_12053,N_13138);
nor U13513 (N_13513,N_12127,N_12253);
nor U13514 (N_13514,N_12335,N_12411);
nand U13515 (N_13515,N_12188,N_12654);
nand U13516 (N_13516,N_13188,N_12056);
nor U13517 (N_13517,N_13054,N_12734);
and U13518 (N_13518,N_13080,N_12729);
xnor U13519 (N_13519,N_13145,N_12933);
nor U13520 (N_13520,N_12767,N_12625);
xnor U13521 (N_13521,N_12981,N_12447);
xnor U13522 (N_13522,N_12903,N_12252);
nor U13523 (N_13523,N_12424,N_12623);
and U13524 (N_13524,N_12901,N_12091);
nor U13525 (N_13525,N_12543,N_12956);
xor U13526 (N_13526,N_12441,N_12740);
or U13527 (N_13527,N_12432,N_12739);
xor U13528 (N_13528,N_12393,N_12155);
nand U13529 (N_13529,N_12904,N_13027);
or U13530 (N_13530,N_12546,N_12206);
xor U13531 (N_13531,N_12889,N_13130);
or U13532 (N_13532,N_12676,N_12354);
nor U13533 (N_13533,N_12306,N_12185);
and U13534 (N_13534,N_12518,N_12537);
or U13535 (N_13535,N_12367,N_12693);
or U13536 (N_13536,N_12800,N_12485);
nor U13537 (N_13537,N_12168,N_12445);
xor U13538 (N_13538,N_12290,N_13096);
nand U13539 (N_13539,N_12016,N_12825);
or U13540 (N_13540,N_12196,N_12225);
xor U13541 (N_13541,N_12730,N_12045);
nor U13542 (N_13542,N_12525,N_13146);
nor U13543 (N_13543,N_12172,N_12014);
nand U13544 (N_13544,N_12262,N_12540);
or U13545 (N_13545,N_12952,N_12937);
xor U13546 (N_13546,N_12890,N_12504);
and U13547 (N_13547,N_12531,N_12170);
xor U13548 (N_13548,N_12268,N_12715);
xnor U13549 (N_13549,N_12094,N_12132);
nand U13550 (N_13550,N_13160,N_13001);
and U13551 (N_13551,N_12137,N_12989);
nor U13552 (N_13552,N_12534,N_13071);
nor U13553 (N_13553,N_12006,N_12129);
and U13554 (N_13554,N_13110,N_12936);
nor U13555 (N_13555,N_12692,N_12607);
nand U13556 (N_13556,N_12671,N_12899);
nand U13557 (N_13557,N_12716,N_12524);
and U13558 (N_13558,N_12513,N_12009);
xor U13559 (N_13559,N_12871,N_13172);
and U13560 (N_13560,N_12437,N_12794);
xor U13561 (N_13561,N_12119,N_12629);
xnor U13562 (N_13562,N_13015,N_12771);
nand U13563 (N_13563,N_12532,N_13095);
nor U13564 (N_13564,N_12024,N_12843);
xnor U13565 (N_13565,N_12113,N_12596);
nor U13566 (N_13566,N_12230,N_12870);
or U13567 (N_13567,N_12911,N_12352);
xnor U13568 (N_13568,N_12382,N_12060);
nor U13569 (N_13569,N_12197,N_13007);
and U13570 (N_13570,N_12063,N_12058);
xor U13571 (N_13571,N_12474,N_12264);
nand U13572 (N_13572,N_12935,N_13061);
nand U13573 (N_13573,N_12799,N_12321);
and U13574 (N_13574,N_12265,N_12773);
nor U13575 (N_13575,N_12471,N_12985);
xnor U13576 (N_13576,N_12074,N_12637);
nand U13577 (N_13577,N_12886,N_12762);
nor U13578 (N_13578,N_13011,N_12616);
nand U13579 (N_13579,N_12670,N_13040);
nand U13580 (N_13580,N_12983,N_12594);
nor U13581 (N_13581,N_12212,N_12681);
or U13582 (N_13582,N_12703,N_12612);
and U13583 (N_13583,N_12640,N_12457);
nand U13584 (N_13584,N_13120,N_13141);
nor U13585 (N_13585,N_12721,N_12922);
and U13586 (N_13586,N_13075,N_12146);
and U13587 (N_13587,N_12635,N_12057);
nor U13588 (N_13588,N_12810,N_12650);
and U13589 (N_13589,N_12000,N_12700);
and U13590 (N_13590,N_12126,N_12327);
nor U13591 (N_13591,N_12752,N_12154);
nor U13592 (N_13592,N_12089,N_12034);
nor U13593 (N_13593,N_12709,N_12959);
and U13594 (N_13594,N_12975,N_12976);
or U13595 (N_13595,N_12414,N_12285);
nand U13596 (N_13596,N_13023,N_12010);
nand U13597 (N_13597,N_12496,N_13088);
or U13598 (N_13598,N_12355,N_12845);
nor U13599 (N_13599,N_12207,N_12638);
nand U13600 (N_13600,N_13128,N_12283);
xor U13601 (N_13601,N_12299,N_12684);
xor U13602 (N_13602,N_12849,N_12332);
nor U13603 (N_13603,N_12209,N_12343);
and U13604 (N_13604,N_13021,N_12674);
nand U13605 (N_13605,N_12529,N_12955);
and U13606 (N_13606,N_13047,N_12888);
nor U13607 (N_13607,N_12719,N_12494);
and U13608 (N_13608,N_12383,N_12920);
and U13609 (N_13609,N_12360,N_12228);
nand U13610 (N_13610,N_12917,N_12679);
and U13611 (N_13611,N_12806,N_12691);
xor U13612 (N_13612,N_12597,N_12044);
and U13613 (N_13613,N_12727,N_13039);
and U13614 (N_13614,N_12812,N_12603);
or U13615 (N_13615,N_12892,N_13159);
nor U13616 (N_13616,N_12788,N_12032);
and U13617 (N_13617,N_12660,N_12784);
or U13618 (N_13618,N_12558,N_12823);
nor U13619 (N_13619,N_12255,N_12215);
nor U13620 (N_13620,N_12502,N_12157);
or U13621 (N_13621,N_12142,N_12409);
nor U13622 (N_13622,N_12731,N_13171);
nor U13623 (N_13623,N_12796,N_12732);
nor U13624 (N_13624,N_12071,N_12499);
and U13625 (N_13625,N_13131,N_12908);
nor U13626 (N_13626,N_12818,N_12419);
nand U13627 (N_13627,N_12139,N_12643);
or U13628 (N_13628,N_12717,N_12960);
nand U13629 (N_13629,N_12924,N_12301);
xnor U13630 (N_13630,N_12093,N_12036);
nor U13631 (N_13631,N_12768,N_12282);
nand U13632 (N_13632,N_12403,N_13067);
nor U13633 (N_13633,N_13073,N_12292);
or U13634 (N_13634,N_12837,N_12018);
nand U13635 (N_13635,N_12897,N_12787);
nand U13636 (N_13636,N_12464,N_12527);
xnor U13637 (N_13637,N_12102,N_12351);
and U13638 (N_13638,N_13161,N_12201);
xnor U13639 (N_13639,N_13049,N_13090);
or U13640 (N_13640,N_12624,N_12829);
xnor U13641 (N_13641,N_12757,N_12705);
and U13642 (N_13642,N_12289,N_12658);
nor U13643 (N_13643,N_13158,N_12226);
nand U13644 (N_13644,N_12059,N_12826);
or U13645 (N_13645,N_12349,N_12192);
xor U13646 (N_13646,N_12634,N_12622);
nand U13647 (N_13647,N_12964,N_12028);
xor U13648 (N_13648,N_12263,N_12515);
or U13649 (N_13649,N_13019,N_12747);
or U13650 (N_13650,N_12760,N_12855);
nand U13651 (N_13651,N_12392,N_13178);
nor U13652 (N_13652,N_12517,N_12160);
nand U13653 (N_13653,N_12405,N_12026);
nand U13654 (N_13654,N_12347,N_12610);
or U13655 (N_13655,N_12114,N_12187);
or U13656 (N_13656,N_12947,N_12303);
and U13657 (N_13657,N_13004,N_12661);
or U13658 (N_13658,N_12281,N_12746);
xnor U13659 (N_13659,N_12180,N_12479);
nor U13660 (N_13660,N_13010,N_12307);
nor U13661 (N_13661,N_12326,N_12795);
and U13662 (N_13662,N_12595,N_12159);
and U13663 (N_13663,N_13065,N_12211);
or U13664 (N_13664,N_13024,N_12753);
or U13665 (N_13665,N_13105,N_12161);
or U13666 (N_13666,N_12582,N_12943);
xnor U13667 (N_13667,N_12541,N_12547);
and U13668 (N_13668,N_12389,N_13153);
nor U13669 (N_13669,N_12011,N_12907);
nor U13670 (N_13670,N_12860,N_12095);
nand U13671 (N_13671,N_12984,N_13100);
nand U13672 (N_13672,N_12556,N_12851);
and U13673 (N_13673,N_12611,N_12442);
or U13674 (N_13674,N_12314,N_12417);
xor U13675 (N_13675,N_12300,N_12217);
or U13676 (N_13676,N_13103,N_12169);
or U13677 (N_13677,N_12696,N_12103);
xor U13678 (N_13678,N_12105,N_12208);
and U13679 (N_13679,N_12274,N_12807);
nand U13680 (N_13680,N_12980,N_12031);
and U13681 (N_13681,N_12495,N_13070);
and U13682 (N_13682,N_12630,N_13087);
and U13683 (N_13683,N_13033,N_12906);
and U13684 (N_13684,N_12153,N_12512);
nand U13685 (N_13685,N_12817,N_13081);
nor U13686 (N_13686,N_12987,N_12087);
nand U13687 (N_13687,N_12181,N_12926);
and U13688 (N_13688,N_12766,N_12368);
nand U13689 (N_13689,N_12864,N_12839);
and U13690 (N_13690,N_12553,N_13107);
xor U13691 (N_13691,N_13196,N_12344);
nand U13692 (N_13692,N_12444,N_12789);
or U13693 (N_13693,N_12190,N_12833);
or U13694 (N_13694,N_12171,N_12573);
nor U13695 (N_13695,N_12785,N_13170);
or U13696 (N_13696,N_12898,N_13116);
nor U13697 (N_13697,N_12338,N_12763);
nor U13698 (N_13698,N_13198,N_12072);
and U13699 (N_13699,N_12148,N_12373);
xnor U13700 (N_13700,N_12484,N_12774);
or U13701 (N_13701,N_12182,N_12145);
or U13702 (N_13702,N_12073,N_12536);
xnor U13703 (N_13703,N_12416,N_12550);
xnor U13704 (N_13704,N_12668,N_13117);
nor U13705 (N_13705,N_12722,N_12463);
xor U13706 (N_13706,N_12808,N_12204);
xor U13707 (N_13707,N_12659,N_12222);
nor U13708 (N_13708,N_12436,N_12714);
or U13709 (N_13709,N_12460,N_12882);
nand U13710 (N_13710,N_12371,N_12293);
or U13711 (N_13711,N_12708,N_12266);
nor U13712 (N_13712,N_12123,N_13108);
and U13713 (N_13713,N_12724,N_12287);
and U13714 (N_13714,N_12013,N_12893);
xor U13715 (N_13715,N_13091,N_13085);
or U13716 (N_13716,N_12745,N_12259);
and U13717 (N_13717,N_12501,N_13191);
or U13718 (N_13718,N_12465,N_12035);
nand U13719 (N_13719,N_12076,N_13077);
nor U13720 (N_13720,N_12193,N_12370);
nor U13721 (N_13721,N_12564,N_12869);
or U13722 (N_13722,N_12415,N_12391);
nor U13723 (N_13723,N_12183,N_12191);
xnor U13724 (N_13724,N_13104,N_12455);
nand U13725 (N_13725,N_12175,N_12652);
and U13726 (N_13726,N_12821,N_12765);
or U13727 (N_13727,N_12050,N_12242);
nor U13728 (N_13728,N_12896,N_12824);
xor U13729 (N_13729,N_12979,N_12856);
nor U13730 (N_13730,N_12857,N_12077);
nand U13731 (N_13731,N_12333,N_12568);
nor U13732 (N_13732,N_12859,N_12542);
and U13733 (N_13733,N_13113,N_12567);
nand U13734 (N_13734,N_12144,N_12988);
xnor U13735 (N_13735,N_13133,N_12064);
xnor U13736 (N_13736,N_12276,N_12117);
and U13737 (N_13737,N_12325,N_12750);
xnor U13738 (N_13738,N_12657,N_12776);
nor U13739 (N_13739,N_12339,N_12510);
nor U13740 (N_13740,N_13043,N_12456);
nand U13741 (N_13741,N_12427,N_12963);
and U13742 (N_13742,N_12374,N_12584);
nor U13743 (N_13743,N_13092,N_12919);
and U13744 (N_13744,N_12560,N_13022);
and U13745 (N_13745,N_12186,N_12883);
or U13746 (N_13746,N_12819,N_12673);
nor U13747 (N_13747,N_12346,N_12134);
and U13748 (N_13748,N_12516,N_13174);
and U13749 (N_13749,N_12434,N_13182);
xor U13750 (N_13750,N_12777,N_12381);
and U13751 (N_13751,N_12022,N_12867);
nand U13752 (N_13752,N_12254,N_13000);
or U13753 (N_13753,N_13199,N_12575);
xor U13754 (N_13754,N_12503,N_12718);
nand U13755 (N_13755,N_12895,N_12706);
or U13756 (N_13756,N_12345,N_12942);
or U13757 (N_13757,N_12397,N_12780);
xor U13758 (N_13758,N_12099,N_12698);
and U13759 (N_13759,N_12048,N_12448);
nand U13760 (N_13760,N_12361,N_12310);
and U13761 (N_13761,N_13190,N_12967);
and U13762 (N_13762,N_12802,N_12167);
xnor U13763 (N_13763,N_13028,N_12816);
and U13764 (N_13764,N_12080,N_12838);
and U13765 (N_13765,N_12385,N_12286);
xnor U13766 (N_13766,N_12055,N_12822);
and U13767 (N_13767,N_12418,N_12555);
and U13768 (N_13768,N_12110,N_12858);
or U13769 (N_13769,N_12130,N_12798);
xor U13770 (N_13770,N_13099,N_12653);
or U13771 (N_13771,N_12615,N_12241);
nor U13772 (N_13772,N_12744,N_12163);
and U13773 (N_13773,N_13154,N_12805);
nor U13774 (N_13774,N_12234,N_12891);
nor U13775 (N_13775,N_13078,N_12357);
nor U13776 (N_13776,N_13089,N_12046);
or U13777 (N_13777,N_12545,N_13165);
nand U13778 (N_13778,N_13053,N_13051);
nor U13779 (N_13779,N_12641,N_12552);
nand U13780 (N_13780,N_12100,N_12877);
and U13781 (N_13781,N_12868,N_12511);
or U13782 (N_13782,N_12372,N_13132);
and U13783 (N_13783,N_12814,N_12862);
nand U13784 (N_13784,N_12999,N_12995);
nor U13785 (N_13785,N_12957,N_12521);
nand U13786 (N_13786,N_12428,N_12426);
and U13787 (N_13787,N_12577,N_12078);
xor U13788 (N_13788,N_13008,N_12604);
xor U13789 (N_13789,N_12633,N_12007);
or U13790 (N_13790,N_12115,N_13112);
or U13791 (N_13791,N_13036,N_12401);
xnor U13792 (N_13792,N_12249,N_12725);
nor U13793 (N_13793,N_12039,N_13058);
and U13794 (N_13794,N_12043,N_12396);
xnor U13795 (N_13795,N_12803,N_12291);
nor U13796 (N_13796,N_12176,N_12376);
xor U13797 (N_13797,N_12938,N_12880);
or U13798 (N_13798,N_12690,N_12909);
and U13799 (N_13799,N_12702,N_13016);
and U13800 (N_13800,N_12569,N_12806);
nand U13801 (N_13801,N_13153,N_13108);
nor U13802 (N_13802,N_12390,N_12441);
nand U13803 (N_13803,N_12653,N_13117);
nor U13804 (N_13804,N_12278,N_12308);
nor U13805 (N_13805,N_12537,N_12621);
and U13806 (N_13806,N_12078,N_12625);
and U13807 (N_13807,N_12355,N_13070);
nor U13808 (N_13808,N_12009,N_12833);
xnor U13809 (N_13809,N_12135,N_12061);
xor U13810 (N_13810,N_12081,N_12339);
and U13811 (N_13811,N_12837,N_12963);
nand U13812 (N_13812,N_12651,N_13092);
and U13813 (N_13813,N_13150,N_12607);
nor U13814 (N_13814,N_12316,N_12027);
nor U13815 (N_13815,N_13060,N_12090);
xor U13816 (N_13816,N_12475,N_12726);
nand U13817 (N_13817,N_12288,N_13184);
and U13818 (N_13818,N_12304,N_12903);
xnor U13819 (N_13819,N_12611,N_12989);
nand U13820 (N_13820,N_12394,N_12556);
nor U13821 (N_13821,N_12395,N_12985);
nor U13822 (N_13822,N_13059,N_12079);
xor U13823 (N_13823,N_12098,N_12611);
nand U13824 (N_13824,N_12424,N_12449);
and U13825 (N_13825,N_12209,N_12949);
or U13826 (N_13826,N_12156,N_12487);
xnor U13827 (N_13827,N_12849,N_12385);
nor U13828 (N_13828,N_12736,N_12936);
nor U13829 (N_13829,N_12251,N_12303);
xnor U13830 (N_13830,N_12247,N_12733);
or U13831 (N_13831,N_12232,N_12591);
or U13832 (N_13832,N_12120,N_12946);
nand U13833 (N_13833,N_12199,N_12961);
or U13834 (N_13834,N_12751,N_12836);
xnor U13835 (N_13835,N_12235,N_12279);
nor U13836 (N_13836,N_13146,N_12975);
nand U13837 (N_13837,N_12774,N_12564);
nand U13838 (N_13838,N_12848,N_12896);
xnor U13839 (N_13839,N_12170,N_12368);
nor U13840 (N_13840,N_12920,N_12182);
and U13841 (N_13841,N_12346,N_13095);
and U13842 (N_13842,N_12140,N_12200);
nor U13843 (N_13843,N_12605,N_12225);
xnor U13844 (N_13844,N_12431,N_12527);
and U13845 (N_13845,N_12213,N_12944);
and U13846 (N_13846,N_13090,N_12657);
nand U13847 (N_13847,N_12275,N_12193);
nand U13848 (N_13848,N_12843,N_12741);
nand U13849 (N_13849,N_12598,N_13129);
and U13850 (N_13850,N_12471,N_12864);
or U13851 (N_13851,N_12709,N_12108);
or U13852 (N_13852,N_12321,N_12908);
xor U13853 (N_13853,N_13036,N_12593);
nand U13854 (N_13854,N_13173,N_12782);
or U13855 (N_13855,N_12081,N_12357);
or U13856 (N_13856,N_12447,N_12168);
nor U13857 (N_13857,N_12081,N_12681);
and U13858 (N_13858,N_12762,N_13005);
xnor U13859 (N_13859,N_12745,N_12092);
nor U13860 (N_13860,N_12591,N_12882);
or U13861 (N_13861,N_12723,N_12419);
or U13862 (N_13862,N_12006,N_13062);
and U13863 (N_13863,N_12660,N_12627);
and U13864 (N_13864,N_12121,N_13034);
nand U13865 (N_13865,N_12542,N_12233);
and U13866 (N_13866,N_13067,N_13020);
or U13867 (N_13867,N_12014,N_12640);
nor U13868 (N_13868,N_12551,N_12550);
and U13869 (N_13869,N_13053,N_12679);
xnor U13870 (N_13870,N_12018,N_12925);
and U13871 (N_13871,N_13089,N_12602);
or U13872 (N_13872,N_12934,N_12155);
nand U13873 (N_13873,N_12366,N_12440);
and U13874 (N_13874,N_12446,N_12960);
and U13875 (N_13875,N_12579,N_13068);
and U13876 (N_13876,N_12963,N_12495);
or U13877 (N_13877,N_12332,N_12555);
xnor U13878 (N_13878,N_12492,N_12800);
xor U13879 (N_13879,N_12040,N_12957);
xor U13880 (N_13880,N_13198,N_12343);
xor U13881 (N_13881,N_12453,N_13030);
nand U13882 (N_13882,N_12015,N_12333);
or U13883 (N_13883,N_12883,N_13055);
or U13884 (N_13884,N_12542,N_12945);
and U13885 (N_13885,N_12728,N_12368);
or U13886 (N_13886,N_13166,N_13111);
xnor U13887 (N_13887,N_12670,N_12126);
nand U13888 (N_13888,N_12335,N_13001);
and U13889 (N_13889,N_12588,N_12581);
or U13890 (N_13890,N_12478,N_12328);
nand U13891 (N_13891,N_12166,N_13164);
or U13892 (N_13892,N_12796,N_12611);
or U13893 (N_13893,N_13139,N_13046);
or U13894 (N_13894,N_12908,N_12810);
xor U13895 (N_13895,N_12644,N_12326);
and U13896 (N_13896,N_13072,N_13181);
nand U13897 (N_13897,N_12567,N_12284);
or U13898 (N_13898,N_12709,N_12132);
xor U13899 (N_13899,N_12649,N_12642);
nor U13900 (N_13900,N_13021,N_12379);
and U13901 (N_13901,N_12188,N_12825);
or U13902 (N_13902,N_12726,N_12804);
or U13903 (N_13903,N_12409,N_12124);
xnor U13904 (N_13904,N_12508,N_12966);
and U13905 (N_13905,N_12123,N_12863);
xor U13906 (N_13906,N_12750,N_12279);
or U13907 (N_13907,N_12914,N_12706);
and U13908 (N_13908,N_13000,N_12205);
and U13909 (N_13909,N_12012,N_12481);
nand U13910 (N_13910,N_12779,N_12131);
xor U13911 (N_13911,N_13103,N_12704);
nand U13912 (N_13912,N_12207,N_12566);
xnor U13913 (N_13913,N_12744,N_12699);
or U13914 (N_13914,N_12864,N_12438);
nand U13915 (N_13915,N_12097,N_12322);
or U13916 (N_13916,N_12599,N_12315);
xor U13917 (N_13917,N_12823,N_12649);
and U13918 (N_13918,N_12376,N_12013);
and U13919 (N_13919,N_12783,N_12730);
or U13920 (N_13920,N_13180,N_12842);
or U13921 (N_13921,N_12560,N_12155);
nor U13922 (N_13922,N_12452,N_12869);
and U13923 (N_13923,N_12696,N_12846);
or U13924 (N_13924,N_13150,N_12620);
and U13925 (N_13925,N_12022,N_12569);
nand U13926 (N_13926,N_12572,N_13138);
or U13927 (N_13927,N_12143,N_12657);
nor U13928 (N_13928,N_12840,N_12783);
or U13929 (N_13929,N_12560,N_13189);
or U13930 (N_13930,N_12606,N_12800);
or U13931 (N_13931,N_12969,N_13100);
xnor U13932 (N_13932,N_12581,N_13157);
or U13933 (N_13933,N_12060,N_12144);
and U13934 (N_13934,N_13041,N_12484);
or U13935 (N_13935,N_12362,N_12318);
nand U13936 (N_13936,N_12288,N_12218);
or U13937 (N_13937,N_12842,N_12124);
xnor U13938 (N_13938,N_13026,N_12998);
and U13939 (N_13939,N_12701,N_12780);
xnor U13940 (N_13940,N_12856,N_13045);
xnor U13941 (N_13941,N_13045,N_13089);
or U13942 (N_13942,N_12245,N_12829);
or U13943 (N_13943,N_12163,N_12757);
xor U13944 (N_13944,N_12588,N_12634);
and U13945 (N_13945,N_13152,N_12919);
and U13946 (N_13946,N_12337,N_12617);
xnor U13947 (N_13947,N_12154,N_12807);
nand U13948 (N_13948,N_13117,N_13181);
or U13949 (N_13949,N_13118,N_12845);
or U13950 (N_13950,N_12638,N_13118);
xor U13951 (N_13951,N_12528,N_12227);
nand U13952 (N_13952,N_12401,N_12078);
xor U13953 (N_13953,N_12622,N_12186);
nand U13954 (N_13954,N_12740,N_12947);
nand U13955 (N_13955,N_12386,N_13129);
or U13956 (N_13956,N_12749,N_13161);
xor U13957 (N_13957,N_12066,N_13096);
nand U13958 (N_13958,N_12195,N_12044);
nand U13959 (N_13959,N_12593,N_12321);
or U13960 (N_13960,N_12398,N_12695);
xnor U13961 (N_13961,N_12823,N_13174);
and U13962 (N_13962,N_12429,N_12913);
and U13963 (N_13963,N_12921,N_12741);
nor U13964 (N_13964,N_12948,N_12047);
xor U13965 (N_13965,N_12927,N_13076);
and U13966 (N_13966,N_12424,N_12628);
xor U13967 (N_13967,N_12202,N_12522);
nand U13968 (N_13968,N_13061,N_12589);
or U13969 (N_13969,N_12753,N_12489);
xor U13970 (N_13970,N_12173,N_12865);
and U13971 (N_13971,N_12480,N_12582);
nand U13972 (N_13972,N_12975,N_12349);
or U13973 (N_13973,N_13045,N_12928);
or U13974 (N_13974,N_13151,N_12886);
or U13975 (N_13975,N_13107,N_12668);
nor U13976 (N_13976,N_12368,N_12398);
and U13977 (N_13977,N_12595,N_13149);
or U13978 (N_13978,N_12435,N_12413);
xnor U13979 (N_13979,N_12813,N_12015);
and U13980 (N_13980,N_12055,N_12103);
nor U13981 (N_13981,N_12368,N_12273);
nand U13982 (N_13982,N_13066,N_13083);
nor U13983 (N_13983,N_12786,N_12226);
or U13984 (N_13984,N_12392,N_13153);
xor U13985 (N_13985,N_12409,N_12239);
or U13986 (N_13986,N_12172,N_13051);
nor U13987 (N_13987,N_12758,N_13063);
xnor U13988 (N_13988,N_12957,N_12315);
nor U13989 (N_13989,N_12124,N_12987);
and U13990 (N_13990,N_12954,N_12909);
xnor U13991 (N_13991,N_12975,N_12262);
nor U13992 (N_13992,N_12801,N_12674);
xnor U13993 (N_13993,N_12188,N_12479);
and U13994 (N_13994,N_12627,N_13034);
xor U13995 (N_13995,N_12472,N_12380);
or U13996 (N_13996,N_12243,N_12303);
xor U13997 (N_13997,N_12879,N_13076);
or U13998 (N_13998,N_13114,N_12002);
and U13999 (N_13999,N_12317,N_12646);
or U14000 (N_14000,N_12859,N_12405);
or U14001 (N_14001,N_12813,N_12763);
or U14002 (N_14002,N_12785,N_12183);
nand U14003 (N_14003,N_12903,N_13101);
or U14004 (N_14004,N_12756,N_12913);
xnor U14005 (N_14005,N_12903,N_12671);
or U14006 (N_14006,N_12842,N_12690);
or U14007 (N_14007,N_12330,N_12067);
or U14008 (N_14008,N_12747,N_12158);
nor U14009 (N_14009,N_12753,N_12082);
and U14010 (N_14010,N_12680,N_12071);
and U14011 (N_14011,N_12403,N_12258);
xnor U14012 (N_14012,N_13096,N_12885);
and U14013 (N_14013,N_12714,N_13109);
xor U14014 (N_14014,N_12306,N_12578);
nor U14015 (N_14015,N_12682,N_12330);
or U14016 (N_14016,N_12404,N_12613);
or U14017 (N_14017,N_13112,N_12831);
or U14018 (N_14018,N_12974,N_12026);
nor U14019 (N_14019,N_13051,N_12344);
nand U14020 (N_14020,N_13103,N_12833);
and U14021 (N_14021,N_13072,N_12722);
xor U14022 (N_14022,N_12626,N_12524);
and U14023 (N_14023,N_12866,N_13169);
nor U14024 (N_14024,N_13054,N_13167);
or U14025 (N_14025,N_12963,N_12553);
nand U14026 (N_14026,N_12629,N_12226);
and U14027 (N_14027,N_12473,N_12372);
xor U14028 (N_14028,N_12682,N_13082);
nand U14029 (N_14029,N_12969,N_12488);
and U14030 (N_14030,N_12763,N_12412);
xor U14031 (N_14031,N_12710,N_12212);
xnor U14032 (N_14032,N_12862,N_12145);
nand U14033 (N_14033,N_12951,N_12577);
nor U14034 (N_14034,N_13003,N_12313);
or U14035 (N_14035,N_13078,N_13063);
xnor U14036 (N_14036,N_12622,N_12484);
nand U14037 (N_14037,N_12352,N_12049);
nand U14038 (N_14038,N_12288,N_12126);
nand U14039 (N_14039,N_12811,N_12032);
nand U14040 (N_14040,N_12022,N_12368);
or U14041 (N_14041,N_12231,N_12479);
xnor U14042 (N_14042,N_12414,N_12912);
or U14043 (N_14043,N_13067,N_12535);
xor U14044 (N_14044,N_12573,N_12651);
xor U14045 (N_14045,N_12852,N_12887);
nor U14046 (N_14046,N_12136,N_12585);
and U14047 (N_14047,N_12863,N_13079);
and U14048 (N_14048,N_13087,N_13094);
xnor U14049 (N_14049,N_12861,N_12198);
nor U14050 (N_14050,N_13185,N_12330);
or U14051 (N_14051,N_12930,N_12928);
and U14052 (N_14052,N_13024,N_12235);
nor U14053 (N_14053,N_12527,N_12777);
or U14054 (N_14054,N_12147,N_12346);
xor U14055 (N_14055,N_13168,N_12906);
and U14056 (N_14056,N_12412,N_12116);
nand U14057 (N_14057,N_13076,N_12694);
and U14058 (N_14058,N_12377,N_12830);
xnor U14059 (N_14059,N_12947,N_12212);
nand U14060 (N_14060,N_12513,N_13038);
nor U14061 (N_14061,N_12486,N_13176);
or U14062 (N_14062,N_12935,N_13063);
nand U14063 (N_14063,N_12619,N_12662);
nand U14064 (N_14064,N_12141,N_12960);
or U14065 (N_14065,N_13110,N_12658);
nor U14066 (N_14066,N_12295,N_12419);
and U14067 (N_14067,N_12914,N_12986);
nand U14068 (N_14068,N_12897,N_12328);
or U14069 (N_14069,N_12739,N_12639);
xor U14070 (N_14070,N_12851,N_12770);
or U14071 (N_14071,N_12543,N_13145);
nor U14072 (N_14072,N_12330,N_13023);
nor U14073 (N_14073,N_12806,N_12338);
nor U14074 (N_14074,N_12954,N_12734);
xnor U14075 (N_14075,N_13011,N_13199);
nand U14076 (N_14076,N_13054,N_12422);
and U14077 (N_14077,N_13121,N_13139);
nor U14078 (N_14078,N_12003,N_12262);
or U14079 (N_14079,N_12730,N_12381);
and U14080 (N_14080,N_12588,N_13193);
nor U14081 (N_14081,N_12060,N_12593);
nor U14082 (N_14082,N_12824,N_12844);
and U14083 (N_14083,N_12232,N_12682);
xnor U14084 (N_14084,N_12286,N_12747);
nand U14085 (N_14085,N_13190,N_12113);
or U14086 (N_14086,N_13119,N_13029);
and U14087 (N_14087,N_12913,N_12880);
and U14088 (N_14088,N_12506,N_12222);
and U14089 (N_14089,N_12652,N_12453);
and U14090 (N_14090,N_12543,N_12000);
nor U14091 (N_14091,N_12319,N_12460);
xnor U14092 (N_14092,N_12083,N_13120);
nand U14093 (N_14093,N_13075,N_12276);
nand U14094 (N_14094,N_12949,N_12725);
xnor U14095 (N_14095,N_12059,N_12362);
nor U14096 (N_14096,N_13008,N_12048);
xnor U14097 (N_14097,N_12482,N_12181);
or U14098 (N_14098,N_12679,N_12109);
nor U14099 (N_14099,N_12011,N_12911);
nor U14100 (N_14100,N_12057,N_12459);
xor U14101 (N_14101,N_12336,N_12297);
and U14102 (N_14102,N_12096,N_12406);
xor U14103 (N_14103,N_12715,N_12378);
and U14104 (N_14104,N_13180,N_13163);
nand U14105 (N_14105,N_12107,N_12889);
nand U14106 (N_14106,N_12682,N_12406);
nand U14107 (N_14107,N_12436,N_12970);
and U14108 (N_14108,N_12679,N_12407);
xor U14109 (N_14109,N_12846,N_13067);
or U14110 (N_14110,N_12485,N_12739);
nand U14111 (N_14111,N_12945,N_12834);
or U14112 (N_14112,N_12676,N_12714);
nand U14113 (N_14113,N_12987,N_12293);
nor U14114 (N_14114,N_12113,N_12433);
nor U14115 (N_14115,N_12416,N_12974);
nor U14116 (N_14116,N_12707,N_12400);
nor U14117 (N_14117,N_12435,N_12829);
and U14118 (N_14118,N_13199,N_12303);
or U14119 (N_14119,N_12493,N_13092);
and U14120 (N_14120,N_12362,N_12543);
or U14121 (N_14121,N_12852,N_12501);
xor U14122 (N_14122,N_12263,N_12911);
nor U14123 (N_14123,N_13019,N_12596);
nand U14124 (N_14124,N_12272,N_12003);
xor U14125 (N_14125,N_12058,N_12947);
nand U14126 (N_14126,N_12753,N_12634);
xor U14127 (N_14127,N_12455,N_12478);
and U14128 (N_14128,N_12520,N_13169);
xor U14129 (N_14129,N_12728,N_13150);
nand U14130 (N_14130,N_12214,N_13098);
nor U14131 (N_14131,N_12605,N_12664);
and U14132 (N_14132,N_12710,N_12531);
or U14133 (N_14133,N_12811,N_12923);
and U14134 (N_14134,N_13074,N_13015);
xnor U14135 (N_14135,N_12281,N_12803);
xor U14136 (N_14136,N_12427,N_12798);
nor U14137 (N_14137,N_13150,N_12249);
and U14138 (N_14138,N_12209,N_12200);
nor U14139 (N_14139,N_13136,N_12463);
xor U14140 (N_14140,N_13030,N_12539);
xor U14141 (N_14141,N_12223,N_12364);
xor U14142 (N_14142,N_12763,N_12818);
nand U14143 (N_14143,N_12983,N_12584);
and U14144 (N_14144,N_12800,N_13172);
nand U14145 (N_14145,N_12618,N_12780);
xnor U14146 (N_14146,N_12396,N_12374);
nand U14147 (N_14147,N_12675,N_13138);
and U14148 (N_14148,N_12056,N_12223);
nor U14149 (N_14149,N_12789,N_12572);
and U14150 (N_14150,N_12731,N_12144);
nor U14151 (N_14151,N_12063,N_12435);
nand U14152 (N_14152,N_12394,N_13099);
nor U14153 (N_14153,N_13019,N_12349);
nand U14154 (N_14154,N_12856,N_12245);
and U14155 (N_14155,N_12582,N_12522);
or U14156 (N_14156,N_12547,N_13125);
nand U14157 (N_14157,N_12073,N_12377);
xnor U14158 (N_14158,N_12533,N_12938);
xor U14159 (N_14159,N_13079,N_12005);
nand U14160 (N_14160,N_12460,N_12060);
nand U14161 (N_14161,N_12062,N_12178);
and U14162 (N_14162,N_12678,N_12116);
nand U14163 (N_14163,N_12962,N_13171);
nand U14164 (N_14164,N_12126,N_12168);
xor U14165 (N_14165,N_12993,N_12603);
or U14166 (N_14166,N_12276,N_13178);
nand U14167 (N_14167,N_12205,N_13144);
nor U14168 (N_14168,N_12380,N_12035);
xnor U14169 (N_14169,N_12193,N_12523);
nand U14170 (N_14170,N_12932,N_12586);
nor U14171 (N_14171,N_12674,N_12861);
xnor U14172 (N_14172,N_12636,N_13114);
nand U14173 (N_14173,N_12119,N_12319);
xor U14174 (N_14174,N_12087,N_12228);
xnor U14175 (N_14175,N_12771,N_13119);
xnor U14176 (N_14176,N_12457,N_12037);
xor U14177 (N_14177,N_12472,N_13066);
xnor U14178 (N_14178,N_12568,N_13006);
nand U14179 (N_14179,N_13181,N_12739);
and U14180 (N_14180,N_12015,N_13144);
and U14181 (N_14181,N_13195,N_12877);
and U14182 (N_14182,N_12404,N_13057);
and U14183 (N_14183,N_12612,N_12280);
xor U14184 (N_14184,N_12382,N_12399);
and U14185 (N_14185,N_12700,N_12539);
and U14186 (N_14186,N_12888,N_12548);
nand U14187 (N_14187,N_12112,N_12559);
and U14188 (N_14188,N_12401,N_12097);
nor U14189 (N_14189,N_12094,N_12077);
xnor U14190 (N_14190,N_12550,N_12445);
or U14191 (N_14191,N_12730,N_12264);
and U14192 (N_14192,N_12681,N_12576);
nand U14193 (N_14193,N_12557,N_12726);
or U14194 (N_14194,N_12689,N_12156);
nor U14195 (N_14195,N_13015,N_13030);
nor U14196 (N_14196,N_12028,N_12609);
nand U14197 (N_14197,N_13076,N_12308);
and U14198 (N_14198,N_12139,N_12677);
xor U14199 (N_14199,N_12712,N_12950);
nor U14200 (N_14200,N_12705,N_12439);
nand U14201 (N_14201,N_12639,N_13086);
xnor U14202 (N_14202,N_12821,N_12502);
xnor U14203 (N_14203,N_12121,N_12342);
xnor U14204 (N_14204,N_12425,N_12842);
or U14205 (N_14205,N_12021,N_12802);
or U14206 (N_14206,N_12285,N_12874);
nand U14207 (N_14207,N_12940,N_12065);
nand U14208 (N_14208,N_13156,N_12848);
and U14209 (N_14209,N_12903,N_12431);
nand U14210 (N_14210,N_12375,N_13076);
nor U14211 (N_14211,N_13188,N_12128);
nand U14212 (N_14212,N_12060,N_12118);
or U14213 (N_14213,N_12402,N_12501);
xnor U14214 (N_14214,N_12968,N_12266);
or U14215 (N_14215,N_13154,N_12689);
and U14216 (N_14216,N_12348,N_12488);
nand U14217 (N_14217,N_13161,N_12917);
and U14218 (N_14218,N_13164,N_12428);
nand U14219 (N_14219,N_12663,N_12322);
nor U14220 (N_14220,N_12344,N_12854);
nor U14221 (N_14221,N_12972,N_12280);
nand U14222 (N_14222,N_12779,N_12817);
and U14223 (N_14223,N_12772,N_12701);
nand U14224 (N_14224,N_12561,N_13041);
or U14225 (N_14225,N_12349,N_13135);
xnor U14226 (N_14226,N_12559,N_12446);
or U14227 (N_14227,N_12183,N_12197);
nand U14228 (N_14228,N_12250,N_12497);
or U14229 (N_14229,N_12879,N_12176);
xor U14230 (N_14230,N_12580,N_12975);
nand U14231 (N_14231,N_12154,N_12261);
or U14232 (N_14232,N_12839,N_12499);
nand U14233 (N_14233,N_12330,N_12226);
and U14234 (N_14234,N_12581,N_13063);
nand U14235 (N_14235,N_12444,N_12700);
nand U14236 (N_14236,N_12226,N_12164);
nand U14237 (N_14237,N_12889,N_12711);
nand U14238 (N_14238,N_12142,N_12569);
nand U14239 (N_14239,N_12402,N_12737);
and U14240 (N_14240,N_12173,N_12156);
nand U14241 (N_14241,N_12508,N_13183);
nor U14242 (N_14242,N_12646,N_12309);
xor U14243 (N_14243,N_12283,N_13072);
nand U14244 (N_14244,N_12326,N_13137);
nor U14245 (N_14245,N_12313,N_12778);
or U14246 (N_14246,N_12307,N_12284);
nand U14247 (N_14247,N_12760,N_12868);
or U14248 (N_14248,N_13007,N_12548);
nand U14249 (N_14249,N_12599,N_12639);
xor U14250 (N_14250,N_12891,N_12039);
nand U14251 (N_14251,N_12114,N_12234);
and U14252 (N_14252,N_12462,N_12240);
xor U14253 (N_14253,N_12961,N_12378);
nor U14254 (N_14254,N_12228,N_13022);
xnor U14255 (N_14255,N_12268,N_12940);
xnor U14256 (N_14256,N_12742,N_12377);
nand U14257 (N_14257,N_12658,N_12699);
or U14258 (N_14258,N_13101,N_13038);
xor U14259 (N_14259,N_12313,N_12344);
xnor U14260 (N_14260,N_12223,N_13001);
xor U14261 (N_14261,N_12210,N_12085);
xor U14262 (N_14262,N_12536,N_12811);
nor U14263 (N_14263,N_12581,N_12413);
nor U14264 (N_14264,N_13110,N_12656);
or U14265 (N_14265,N_13068,N_13179);
nand U14266 (N_14266,N_12096,N_12009);
and U14267 (N_14267,N_12275,N_12132);
and U14268 (N_14268,N_12284,N_12396);
nor U14269 (N_14269,N_12582,N_12495);
and U14270 (N_14270,N_13079,N_12296);
nand U14271 (N_14271,N_13134,N_12905);
nand U14272 (N_14272,N_13086,N_12144);
nor U14273 (N_14273,N_12667,N_12070);
or U14274 (N_14274,N_12486,N_12047);
and U14275 (N_14275,N_12840,N_13177);
or U14276 (N_14276,N_13183,N_12433);
and U14277 (N_14277,N_13125,N_13004);
or U14278 (N_14278,N_12600,N_12385);
xor U14279 (N_14279,N_12514,N_13114);
or U14280 (N_14280,N_12241,N_12297);
nor U14281 (N_14281,N_13096,N_12285);
nor U14282 (N_14282,N_13185,N_12873);
and U14283 (N_14283,N_12767,N_12230);
and U14284 (N_14284,N_12625,N_12640);
nor U14285 (N_14285,N_13092,N_13036);
nor U14286 (N_14286,N_12038,N_12449);
and U14287 (N_14287,N_12287,N_12950);
nand U14288 (N_14288,N_12617,N_13134);
nor U14289 (N_14289,N_12223,N_13080);
nor U14290 (N_14290,N_13156,N_12163);
or U14291 (N_14291,N_12769,N_12687);
nor U14292 (N_14292,N_12834,N_12361);
nor U14293 (N_14293,N_12758,N_12450);
and U14294 (N_14294,N_13167,N_12068);
and U14295 (N_14295,N_12645,N_13028);
nor U14296 (N_14296,N_12895,N_12217);
xor U14297 (N_14297,N_12009,N_12328);
nand U14298 (N_14298,N_12633,N_12711);
nand U14299 (N_14299,N_13094,N_12617);
or U14300 (N_14300,N_12836,N_12510);
nor U14301 (N_14301,N_12888,N_12795);
xnor U14302 (N_14302,N_13028,N_12439);
nand U14303 (N_14303,N_13148,N_12162);
nor U14304 (N_14304,N_12060,N_13146);
and U14305 (N_14305,N_12293,N_12484);
and U14306 (N_14306,N_13102,N_12416);
and U14307 (N_14307,N_13093,N_12787);
nor U14308 (N_14308,N_12110,N_12084);
and U14309 (N_14309,N_12883,N_12156);
nor U14310 (N_14310,N_12817,N_12608);
nor U14311 (N_14311,N_12000,N_13177);
or U14312 (N_14312,N_12451,N_12038);
and U14313 (N_14313,N_13186,N_12832);
and U14314 (N_14314,N_12910,N_12854);
or U14315 (N_14315,N_12957,N_12246);
or U14316 (N_14316,N_12861,N_12920);
nand U14317 (N_14317,N_12772,N_12765);
nand U14318 (N_14318,N_12220,N_12751);
and U14319 (N_14319,N_13082,N_12259);
and U14320 (N_14320,N_12615,N_12688);
nor U14321 (N_14321,N_12292,N_12556);
xor U14322 (N_14322,N_12170,N_12932);
nor U14323 (N_14323,N_13051,N_12780);
nor U14324 (N_14324,N_12432,N_12272);
and U14325 (N_14325,N_12522,N_12385);
or U14326 (N_14326,N_12992,N_12748);
xnor U14327 (N_14327,N_13012,N_12057);
nor U14328 (N_14328,N_13183,N_12449);
xnor U14329 (N_14329,N_12802,N_12898);
or U14330 (N_14330,N_12640,N_12303);
nand U14331 (N_14331,N_12465,N_12600);
nand U14332 (N_14332,N_12852,N_13194);
nor U14333 (N_14333,N_12383,N_12021);
or U14334 (N_14334,N_13070,N_12213);
xor U14335 (N_14335,N_12116,N_12817);
or U14336 (N_14336,N_12032,N_12507);
and U14337 (N_14337,N_12305,N_12364);
and U14338 (N_14338,N_12028,N_13024);
xor U14339 (N_14339,N_12217,N_13173);
nor U14340 (N_14340,N_12170,N_12329);
nand U14341 (N_14341,N_12691,N_12502);
and U14342 (N_14342,N_12820,N_12816);
nor U14343 (N_14343,N_12822,N_13102);
nor U14344 (N_14344,N_12928,N_12485);
nor U14345 (N_14345,N_13064,N_13131);
nor U14346 (N_14346,N_12823,N_12619);
or U14347 (N_14347,N_12717,N_12835);
and U14348 (N_14348,N_12505,N_12579);
nor U14349 (N_14349,N_12454,N_12418);
or U14350 (N_14350,N_12935,N_12269);
nor U14351 (N_14351,N_13053,N_12098);
nor U14352 (N_14352,N_12601,N_12348);
and U14353 (N_14353,N_12796,N_12189);
xor U14354 (N_14354,N_12162,N_12518);
nor U14355 (N_14355,N_12466,N_13151);
or U14356 (N_14356,N_12862,N_12402);
nand U14357 (N_14357,N_13132,N_12446);
and U14358 (N_14358,N_13034,N_13041);
xor U14359 (N_14359,N_12515,N_12758);
and U14360 (N_14360,N_12507,N_12993);
xor U14361 (N_14361,N_12391,N_13055);
nor U14362 (N_14362,N_12390,N_13154);
nor U14363 (N_14363,N_12418,N_12532);
and U14364 (N_14364,N_12490,N_12865);
xnor U14365 (N_14365,N_12437,N_12992);
nor U14366 (N_14366,N_13016,N_12286);
xnor U14367 (N_14367,N_12200,N_12591);
nor U14368 (N_14368,N_12053,N_12307);
nor U14369 (N_14369,N_12857,N_12209);
nand U14370 (N_14370,N_12302,N_12564);
nor U14371 (N_14371,N_12319,N_13049);
nor U14372 (N_14372,N_12674,N_12124);
nor U14373 (N_14373,N_12007,N_12236);
nor U14374 (N_14374,N_13095,N_12629);
or U14375 (N_14375,N_12149,N_12591);
and U14376 (N_14376,N_13076,N_13020);
and U14377 (N_14377,N_12159,N_12253);
and U14378 (N_14378,N_12759,N_12007);
or U14379 (N_14379,N_12034,N_12917);
nor U14380 (N_14380,N_12731,N_12109);
xnor U14381 (N_14381,N_12892,N_13192);
nor U14382 (N_14382,N_12094,N_13040);
xor U14383 (N_14383,N_12712,N_12152);
and U14384 (N_14384,N_12374,N_12372);
nor U14385 (N_14385,N_12791,N_12581);
xor U14386 (N_14386,N_12220,N_12623);
or U14387 (N_14387,N_12370,N_12225);
xnor U14388 (N_14388,N_12178,N_12179);
or U14389 (N_14389,N_12517,N_12923);
xor U14390 (N_14390,N_12897,N_12293);
xor U14391 (N_14391,N_12049,N_12085);
xor U14392 (N_14392,N_12799,N_12094);
nor U14393 (N_14393,N_12114,N_13160);
and U14394 (N_14394,N_12977,N_12292);
nand U14395 (N_14395,N_12506,N_12135);
nor U14396 (N_14396,N_12203,N_12670);
nand U14397 (N_14397,N_12939,N_12000);
or U14398 (N_14398,N_12931,N_12790);
and U14399 (N_14399,N_13111,N_13080);
and U14400 (N_14400,N_13670,N_14384);
nor U14401 (N_14401,N_13437,N_13946);
xnor U14402 (N_14402,N_14185,N_14157);
and U14403 (N_14403,N_13264,N_13868);
or U14404 (N_14404,N_14213,N_13660);
and U14405 (N_14405,N_14329,N_13518);
nor U14406 (N_14406,N_13656,N_13385);
xor U14407 (N_14407,N_13335,N_14042);
or U14408 (N_14408,N_13635,N_13399);
nand U14409 (N_14409,N_13957,N_13807);
nand U14410 (N_14410,N_14046,N_13879);
and U14411 (N_14411,N_14214,N_14210);
nand U14412 (N_14412,N_14339,N_14179);
or U14413 (N_14413,N_14102,N_14393);
nand U14414 (N_14414,N_14034,N_14357);
nand U14415 (N_14415,N_13625,N_13228);
nor U14416 (N_14416,N_13482,N_13369);
or U14417 (N_14417,N_13241,N_13654);
and U14418 (N_14418,N_13966,N_13576);
nand U14419 (N_14419,N_13422,N_14212);
nor U14420 (N_14420,N_13700,N_13722);
or U14421 (N_14421,N_14387,N_13507);
xor U14422 (N_14422,N_13371,N_13711);
xnor U14423 (N_14423,N_13651,N_13444);
or U14424 (N_14424,N_13995,N_13843);
xnor U14425 (N_14425,N_14146,N_13740);
xor U14426 (N_14426,N_13780,N_13208);
xnor U14427 (N_14427,N_13569,N_14031);
nand U14428 (N_14428,N_13585,N_13752);
and U14429 (N_14429,N_13288,N_14094);
nand U14430 (N_14430,N_13909,N_14089);
nor U14431 (N_14431,N_13336,N_13624);
nand U14432 (N_14432,N_14278,N_14095);
nor U14433 (N_14433,N_14349,N_13827);
nand U14434 (N_14434,N_13748,N_13575);
and U14435 (N_14435,N_13767,N_14048);
xnor U14436 (N_14436,N_13499,N_13560);
nor U14437 (N_14437,N_13955,N_14172);
nor U14438 (N_14438,N_14373,N_13447);
nand U14439 (N_14439,N_13796,N_14336);
and U14440 (N_14440,N_13339,N_14334);
nor U14441 (N_14441,N_13936,N_13834);
nand U14442 (N_14442,N_13380,N_13875);
xnor U14443 (N_14443,N_13242,N_13856);
or U14444 (N_14444,N_13218,N_13914);
or U14445 (N_14445,N_13311,N_13268);
xnor U14446 (N_14446,N_13490,N_13532);
or U14447 (N_14447,N_13838,N_13452);
nor U14448 (N_14448,N_13564,N_13679);
or U14449 (N_14449,N_14242,N_14366);
nand U14450 (N_14450,N_14104,N_13605);
xnor U14451 (N_14451,N_13392,N_14251);
nand U14452 (N_14452,N_13446,N_13474);
or U14453 (N_14453,N_14144,N_13500);
or U14454 (N_14454,N_14309,N_13787);
or U14455 (N_14455,N_13915,N_14380);
nand U14456 (N_14456,N_13816,N_13309);
xnor U14457 (N_14457,N_13993,N_13982);
nand U14458 (N_14458,N_13769,N_13550);
nand U14459 (N_14459,N_13898,N_13960);
nor U14460 (N_14460,N_13599,N_14300);
and U14461 (N_14461,N_13561,N_14347);
and U14462 (N_14462,N_14346,N_13979);
or U14463 (N_14463,N_13928,N_13233);
and U14464 (N_14464,N_13299,N_13744);
and U14465 (N_14465,N_13871,N_14388);
or U14466 (N_14466,N_13483,N_13872);
nand U14467 (N_14467,N_14353,N_13249);
and U14468 (N_14468,N_13859,N_14039);
or U14469 (N_14469,N_14147,N_13959);
or U14470 (N_14470,N_13703,N_14083);
xnor U14471 (N_14471,N_13906,N_13847);
nand U14472 (N_14472,N_14078,N_13319);
nand U14473 (N_14473,N_13831,N_14047);
nand U14474 (N_14474,N_13940,N_13985);
nor U14475 (N_14475,N_14389,N_13534);
nand U14476 (N_14476,N_14090,N_13893);
and U14477 (N_14477,N_14071,N_14222);
nand U14478 (N_14478,N_13902,N_13676);
and U14479 (N_14479,N_14323,N_13211);
or U14480 (N_14480,N_13954,N_13461);
nand U14481 (N_14481,N_14020,N_13379);
nor U14482 (N_14482,N_14316,N_13892);
and U14483 (N_14483,N_13750,N_13301);
nand U14484 (N_14484,N_14112,N_14129);
nor U14485 (N_14485,N_13222,N_13629);
nand U14486 (N_14486,N_13376,N_13925);
and U14487 (N_14487,N_14010,N_14209);
nor U14488 (N_14488,N_13470,N_13227);
or U14489 (N_14489,N_13287,N_13328);
or U14490 (N_14490,N_14162,N_13590);
and U14491 (N_14491,N_14196,N_13214);
and U14492 (N_14492,N_14063,N_14062);
nor U14493 (N_14493,N_14092,N_13673);
or U14494 (N_14494,N_13506,N_13808);
nand U14495 (N_14495,N_13696,N_14365);
or U14496 (N_14496,N_13795,N_13741);
nand U14497 (N_14497,N_13855,N_13934);
xnor U14498 (N_14498,N_14355,N_14382);
or U14499 (N_14499,N_13354,N_13495);
nor U14500 (N_14500,N_13964,N_13640);
or U14501 (N_14501,N_13753,N_14392);
and U14502 (N_14502,N_13207,N_13937);
nand U14503 (N_14503,N_14176,N_13996);
xnor U14504 (N_14504,N_13873,N_14275);
or U14505 (N_14505,N_14325,N_13215);
or U14506 (N_14506,N_13688,N_14301);
xnor U14507 (N_14507,N_13861,N_14002);
or U14508 (N_14508,N_13201,N_13721);
and U14509 (N_14509,N_14120,N_14293);
nand U14510 (N_14510,N_14158,N_14226);
nand U14511 (N_14511,N_14398,N_13597);
nand U14512 (N_14512,N_14271,N_13373);
nand U14513 (N_14513,N_14198,N_14156);
nand U14514 (N_14514,N_13313,N_13323);
nor U14515 (N_14515,N_13607,N_13205);
xnor U14516 (N_14516,N_14169,N_13238);
or U14517 (N_14517,N_14109,N_13970);
nor U14518 (N_14518,N_13984,N_13403);
or U14519 (N_14519,N_14099,N_14183);
xnor U14520 (N_14520,N_13972,N_13848);
and U14521 (N_14521,N_13484,N_14247);
xnor U14522 (N_14522,N_13743,N_14007);
and U14523 (N_14523,N_13684,N_14065);
and U14524 (N_14524,N_14106,N_13219);
or U14525 (N_14525,N_14233,N_13917);
nand U14526 (N_14526,N_13273,N_13286);
nand U14527 (N_14527,N_13505,N_13952);
xor U14528 (N_14528,N_14283,N_13536);
nor U14529 (N_14529,N_13747,N_14148);
nand U14530 (N_14530,N_14320,N_13876);
nand U14531 (N_14531,N_13489,N_13388);
nand U14532 (N_14532,N_13347,N_14221);
or U14533 (N_14533,N_14391,N_14216);
or U14534 (N_14534,N_14311,N_14282);
or U14535 (N_14535,N_13239,N_13329);
and U14536 (N_14536,N_13920,N_13768);
and U14537 (N_14537,N_13641,N_13653);
and U14538 (N_14538,N_13551,N_13573);
nor U14539 (N_14539,N_13887,N_13820);
nor U14540 (N_14540,N_13366,N_13666);
nor U14541 (N_14541,N_14115,N_13368);
and U14542 (N_14542,N_14269,N_13874);
nand U14543 (N_14543,N_14361,N_13969);
and U14544 (N_14544,N_14004,N_13316);
nand U14545 (N_14545,N_13738,N_13886);
and U14546 (N_14546,N_14113,N_13298);
nor U14547 (N_14547,N_13200,N_14088);
xor U14548 (N_14548,N_13284,N_14091);
and U14549 (N_14549,N_13459,N_13511);
nand U14550 (N_14550,N_13720,N_13938);
and U14551 (N_14551,N_13812,N_14135);
xor U14552 (N_14552,N_14204,N_14367);
or U14553 (N_14553,N_13332,N_13804);
nand U14554 (N_14554,N_13870,N_13839);
nand U14555 (N_14555,N_13442,N_13468);
or U14556 (N_14556,N_14197,N_13357);
nand U14557 (N_14557,N_13932,N_13594);
and U14558 (N_14558,N_14175,N_14189);
or U14559 (N_14559,N_14273,N_13644);
and U14560 (N_14560,N_13562,N_13510);
nand U14561 (N_14561,N_13389,N_13983);
nand U14562 (N_14562,N_13626,N_14161);
nand U14563 (N_14563,N_13467,N_14333);
xor U14564 (N_14564,N_14246,N_13669);
xnor U14565 (N_14565,N_14376,N_13690);
nand U14566 (N_14566,N_14289,N_13846);
or U14567 (N_14567,N_14192,N_13707);
nor U14568 (N_14568,N_13694,N_13760);
nand U14569 (N_14569,N_13358,N_13714);
nor U14570 (N_14570,N_14082,N_13315);
and U14571 (N_14571,N_13776,N_13863);
xnor U14572 (N_14572,N_13458,N_14011);
nor U14573 (N_14573,N_14267,N_13210);
nor U14574 (N_14574,N_14338,N_13338);
xnor U14575 (N_14575,N_14314,N_13782);
nand U14576 (N_14576,N_13475,N_13553);
and U14577 (N_14577,N_13968,N_13614);
nand U14578 (N_14578,N_13430,N_13426);
or U14579 (N_14579,N_14304,N_13680);
or U14580 (N_14580,N_14170,N_13501);
nor U14581 (N_14581,N_14043,N_13926);
or U14582 (N_14582,N_13420,N_13988);
or U14583 (N_14583,N_13734,N_13465);
nor U14584 (N_14584,N_13897,N_13327);
and U14585 (N_14585,N_13685,N_13657);
and U14586 (N_14586,N_14307,N_14395);
or U14587 (N_14587,N_13334,N_13419);
or U14588 (N_14588,N_13726,N_13217);
nand U14589 (N_14589,N_13824,N_13253);
or U14590 (N_14590,N_13903,N_13931);
and U14591 (N_14591,N_14318,N_14239);
nand U14592 (N_14592,N_14023,N_13310);
nand U14593 (N_14593,N_14211,N_13942);
xnor U14594 (N_14594,N_13455,N_13882);
or U14595 (N_14595,N_14126,N_14305);
or U14596 (N_14596,N_14360,N_13727);
and U14597 (N_14597,N_14080,N_13302);
nor U14598 (N_14598,N_13849,N_13520);
nor U14599 (N_14599,N_13853,N_13477);
and U14600 (N_14600,N_14150,N_13255);
xnor U14601 (N_14601,N_13819,N_13337);
nand U14602 (N_14602,N_14060,N_14155);
or U14603 (N_14603,N_13735,N_13413);
nand U14604 (N_14604,N_13616,N_14397);
or U14605 (N_14605,N_13258,N_14036);
or U14606 (N_14606,N_14364,N_13981);
and U14607 (N_14607,N_13251,N_13826);
and U14608 (N_14608,N_13622,N_13770);
xor U14609 (N_14609,N_13320,N_13252);
xnor U14610 (N_14610,N_13331,N_13910);
nor U14611 (N_14611,N_13300,N_13877);
or U14612 (N_14612,N_13404,N_13757);
and U14613 (N_14613,N_13888,N_14041);
xor U14614 (N_14614,N_14245,N_13415);
and U14615 (N_14615,N_13372,N_13649);
xnor U14616 (N_14616,N_14055,N_14165);
nand U14617 (N_14617,N_13643,N_13204);
nor U14618 (N_14618,N_14243,N_13555);
nand U14619 (N_14619,N_14138,N_14000);
or U14620 (N_14620,N_14199,N_13999);
or U14621 (N_14621,N_13686,N_14324);
xor U14622 (N_14622,N_14027,N_13650);
xor U14623 (N_14623,N_13529,N_14200);
and U14624 (N_14624,N_14371,N_13850);
nand U14625 (N_14625,N_13527,N_13541);
and U14626 (N_14626,N_13783,N_13929);
nor U14627 (N_14627,N_13628,N_14014);
nor U14628 (N_14628,N_14280,N_13351);
xor U14629 (N_14629,N_13277,N_14114);
or U14630 (N_14630,N_13509,N_14327);
xor U14631 (N_14631,N_14375,N_13502);
nand U14632 (N_14632,N_13784,N_14345);
nor U14633 (N_14633,N_14348,N_13647);
or U14634 (N_14634,N_13836,N_13531);
and U14635 (N_14635,N_13278,N_13733);
nor U14636 (N_14636,N_13570,N_13689);
nand U14637 (N_14637,N_14117,N_13466);
nand U14638 (N_14638,N_13491,N_14313);
and U14639 (N_14639,N_13758,N_14064);
and U14640 (N_14640,N_13405,N_13237);
nor U14641 (N_14641,N_14040,N_14207);
and U14642 (N_14642,N_13709,N_13266);
or U14643 (N_14643,N_13588,N_13860);
nand U14644 (N_14644,N_13514,N_14296);
nor U14645 (N_14645,N_13678,N_13386);
or U14646 (N_14646,N_13451,N_13907);
xnor U14647 (N_14647,N_14359,N_13213);
or U14648 (N_14648,N_14342,N_13225);
or U14649 (N_14649,N_14033,N_13355);
xor U14650 (N_14650,N_13958,N_13718);
nor U14651 (N_14651,N_14107,N_13542);
nand U14652 (N_14652,N_14141,N_13481);
nor U14653 (N_14653,N_14369,N_14208);
xnor U14654 (N_14654,N_13828,N_13798);
or U14655 (N_14655,N_13270,N_14038);
and U14656 (N_14656,N_13785,N_13781);
xnor U14657 (N_14657,N_13280,N_14317);
and U14658 (N_14658,N_13504,N_14328);
and U14659 (N_14659,N_13851,N_13203);
and U14660 (N_14660,N_13971,N_13589);
nand U14661 (N_14661,N_13433,N_13818);
or U14662 (N_14662,N_13579,N_13558);
or U14663 (N_14663,N_14035,N_13674);
nand U14664 (N_14664,N_13540,N_14276);
nor U14665 (N_14665,N_14285,N_13441);
nand U14666 (N_14666,N_14250,N_13880);
nor U14667 (N_14667,N_13487,N_14291);
xnor U14668 (N_14668,N_14279,N_13279);
nor U14669 (N_14669,N_13580,N_14191);
or U14670 (N_14670,N_14193,N_14206);
nor U14671 (N_14671,N_13445,N_14101);
xor U14672 (N_14672,N_13609,N_13845);
and U14673 (N_14673,N_14153,N_14385);
nor U14674 (N_14674,N_13916,N_13240);
nor U14675 (N_14675,N_14234,N_13811);
and U14676 (N_14676,N_14337,N_13692);
xnor U14677 (N_14677,N_13236,N_13620);
and U14678 (N_14678,N_13608,N_13391);
and U14679 (N_14679,N_13256,N_14136);
or U14680 (N_14680,N_14264,N_14287);
and U14681 (N_14681,N_14259,N_14274);
or U14682 (N_14682,N_13432,N_14315);
nand U14683 (N_14683,N_13434,N_13598);
nor U14684 (N_14684,N_13535,N_14186);
or U14685 (N_14685,N_13746,N_14070);
and U14686 (N_14686,N_13209,N_13642);
xnor U14687 (N_14687,N_13751,N_13922);
xnor U14688 (N_14688,N_13923,N_13627);
or U14689 (N_14689,N_14378,N_13544);
and U14690 (N_14690,N_13905,N_13621);
nor U14691 (N_14691,N_13900,N_13263);
or U14692 (N_14692,N_14167,N_14330);
nand U14693 (N_14693,N_13944,N_14195);
or U14694 (N_14694,N_13293,N_13414);
xor U14695 (N_14695,N_13687,N_13763);
nand U14696 (N_14696,N_13844,N_13581);
xor U14697 (N_14697,N_14383,N_14030);
nor U14698 (N_14698,N_14119,N_13658);
and U14699 (N_14699,N_13591,N_13899);
nor U14700 (N_14700,N_13409,N_13927);
or U14701 (N_14701,N_13889,N_13739);
or U14702 (N_14702,N_13494,N_13584);
xor U14703 (N_14703,N_13832,N_14142);
nand U14704 (N_14704,N_13539,N_14252);
nand U14705 (N_14705,N_13633,N_14021);
nand U14706 (N_14706,N_13630,N_14025);
nor U14707 (N_14707,N_13664,N_14077);
nand U14708 (N_14708,N_13401,N_13717);
and U14709 (N_14709,N_13362,N_14261);
nor U14710 (N_14710,N_13411,N_13324);
nand U14711 (N_14711,N_13572,N_14132);
nor U14712 (N_14712,N_14128,N_14254);
or U14713 (N_14713,N_14232,N_13830);
and U14714 (N_14714,N_13712,N_14013);
and U14715 (N_14715,N_14032,N_13503);
xnor U14716 (N_14716,N_13681,N_13406);
nand U14717 (N_14717,N_13755,N_13704);
xor U14718 (N_14718,N_13476,N_14321);
and U14719 (N_14719,N_13947,N_14164);
and U14720 (N_14720,N_13350,N_13600);
nor U14721 (N_14721,N_13693,N_13454);
nand U14722 (N_14722,N_13883,N_14100);
or U14723 (N_14723,N_13563,N_13774);
nand U14724 (N_14724,N_13878,N_14220);
nor U14725 (N_14725,N_13691,N_13567);
or U14726 (N_14726,N_13314,N_14399);
or U14727 (N_14727,N_14236,N_13809);
and U14728 (N_14728,N_13728,N_14332);
nand U14729 (N_14729,N_14139,N_13276);
nand U14730 (N_14730,N_14093,N_13566);
or U14731 (N_14731,N_14056,N_13961);
or U14732 (N_14732,N_14306,N_13574);
nand U14733 (N_14733,N_14024,N_14137);
and U14734 (N_14734,N_13800,N_13416);
nor U14735 (N_14735,N_14012,N_13360);
and U14736 (N_14736,N_13202,N_13761);
nor U14737 (N_14737,N_13552,N_13854);
and U14738 (N_14738,N_13973,N_14066);
or U14739 (N_14739,N_13583,N_14096);
or U14740 (N_14740,N_13431,N_13423);
and U14741 (N_14741,N_13655,N_14168);
nand U14742 (N_14742,N_13516,N_13479);
nor U14743 (N_14743,N_13901,N_14086);
nand U14744 (N_14744,N_13904,N_13601);
or U14745 (N_14745,N_13815,N_14160);
or U14746 (N_14746,N_13517,N_13646);
nand U14747 (N_14747,N_13425,N_13261);
nand U14748 (N_14748,N_13639,N_13374);
nor U14749 (N_14749,N_14235,N_13648);
or U14750 (N_14750,N_13449,N_13364);
or U14751 (N_14751,N_14068,N_13464);
and U14752 (N_14752,N_13797,N_13443);
nor U14753 (N_14753,N_13636,N_13611);
nor U14754 (N_14754,N_13297,N_13408);
or U14755 (N_14755,N_13448,N_13226);
or U14756 (N_14756,N_13548,N_13559);
nor U14757 (N_14757,N_14044,N_14370);
xor U14758 (N_14758,N_14260,N_13867);
xnor U14759 (N_14759,N_14178,N_13356);
nor U14760 (N_14760,N_13488,N_14331);
and U14761 (N_14761,N_13440,N_14008);
and U14762 (N_14762,N_13330,N_14029);
nand U14763 (N_14763,N_14223,N_13813);
xnor U14764 (N_14764,N_13456,N_13948);
and U14765 (N_14765,N_14085,N_14069);
or U14766 (N_14766,N_13632,N_14340);
nor U14767 (N_14767,N_13305,N_13894);
or U14768 (N_14768,N_13393,N_13394);
and U14769 (N_14769,N_13450,N_13306);
or U14770 (N_14770,N_14270,N_14374);
or U14771 (N_14771,N_14202,N_13267);
and U14772 (N_14772,N_13715,N_13852);
nor U14773 (N_14773,N_14177,N_13260);
nor U14774 (N_14774,N_14182,N_13604);
or U14775 (N_14775,N_14268,N_13478);
nand U14776 (N_14776,N_14187,N_14238);
and U14777 (N_14777,N_14127,N_14072);
nor U14778 (N_14778,N_13810,N_13556);
nor U14779 (N_14779,N_13930,N_13990);
and U14780 (N_14780,N_13496,N_13821);
xor U14781 (N_14781,N_13592,N_13992);
nor U14782 (N_14782,N_14299,N_13775);
xnor U14783 (N_14783,N_13383,N_14103);
or U14784 (N_14784,N_14130,N_13732);
or U14785 (N_14785,N_13216,N_13571);
nor U14786 (N_14786,N_14005,N_13547);
xor U14787 (N_14787,N_13349,N_13671);
nand U14788 (N_14788,N_13515,N_14075);
or U14789 (N_14789,N_14231,N_13662);
xnor U14790 (N_14790,N_13453,N_14229);
xnor U14791 (N_14791,N_13759,N_13603);
and U14792 (N_14792,N_13956,N_13924);
xor U14793 (N_14793,N_14118,N_13220);
nand U14794 (N_14794,N_14341,N_13943);
or U14795 (N_14795,N_13949,N_13865);
or U14796 (N_14796,N_14108,N_13524);
or U14797 (N_14797,N_13976,N_13799);
xor U14798 (N_14798,N_13792,N_14131);
or U14799 (N_14799,N_13377,N_13471);
nor U14800 (N_14800,N_14372,N_13773);
xnor U14801 (N_14801,N_13619,N_14225);
and U14802 (N_14802,N_14001,N_13232);
nand U14803 (N_14803,N_13421,N_14003);
or U14804 (N_14804,N_13342,N_14263);
and U14805 (N_14805,N_13840,N_14110);
nor U14806 (N_14806,N_13699,N_13424);
or U14807 (N_14807,N_13869,N_14217);
and U14808 (N_14808,N_13989,N_13533);
nand U14809 (N_14809,N_13742,N_14352);
and U14810 (N_14810,N_13480,N_14351);
and U14811 (N_14811,N_13212,N_13730);
nand U14812 (N_14812,N_14277,N_13918);
nor U14813 (N_14813,N_13790,N_13397);
xor U14814 (N_14814,N_13719,N_13986);
or U14815 (N_14815,N_13912,N_14049);
xor U14816 (N_14816,N_13675,N_13708);
and U14817 (N_14817,N_13230,N_14362);
nor U14818 (N_14818,N_13457,N_14084);
nor U14819 (N_14819,N_13395,N_13530);
nand U14820 (N_14820,N_14019,N_13596);
or U14821 (N_14821,N_14149,N_13842);
and U14822 (N_14822,N_13396,N_14249);
nor U14823 (N_14823,N_14151,N_13295);
nor U14824 (N_14824,N_13638,N_14188);
nor U14825 (N_14825,N_13617,N_13521);
nor U14826 (N_14826,N_14016,N_13265);
nand U14827 (N_14827,N_14180,N_13921);
and U14828 (N_14828,N_13884,N_14116);
or U14829 (N_14829,N_13460,N_14363);
xor U14830 (N_14830,N_14152,N_14344);
xor U14831 (N_14831,N_13231,N_13363);
or U14832 (N_14832,N_13677,N_13724);
nor U14833 (N_14833,N_14262,N_13308);
nor U14834 (N_14834,N_13602,N_14097);
nand U14835 (N_14835,N_13762,N_14292);
nand U14836 (N_14836,N_13365,N_14163);
xor U14837 (N_14837,N_13289,N_14227);
and U14838 (N_14838,N_13885,N_14073);
nand U14839 (N_14839,N_14241,N_13428);
and U14840 (N_14840,N_13290,N_13593);
nand U14841 (N_14841,N_14054,N_14058);
xor U14842 (N_14842,N_14173,N_13485);
xor U14843 (N_14843,N_14244,N_14015);
xnor U14844 (N_14844,N_13340,N_14218);
nand U14845 (N_14845,N_13754,N_13522);
or U14846 (N_14846,N_13412,N_13435);
and U14847 (N_14847,N_13262,N_13987);
nand U14848 (N_14848,N_13294,N_14266);
xor U14849 (N_14849,N_13789,N_13244);
nor U14850 (N_14850,N_13367,N_13341);
nand U14851 (N_14851,N_14111,N_13493);
nand U14852 (N_14852,N_13224,N_13513);
nor U14853 (N_14853,N_13829,N_14154);
or U14854 (N_14854,N_13822,N_14051);
nor U14855 (N_14855,N_14052,N_13545);
nor U14856 (N_14856,N_14368,N_13398);
and U14857 (N_14857,N_13269,N_13805);
or U14858 (N_14858,N_13317,N_13361);
and U14859 (N_14859,N_14294,N_14074);
nand U14860 (N_14860,N_13587,N_13967);
xnor U14861 (N_14861,N_13418,N_14205);
nor U14862 (N_14862,N_13469,N_13407);
nor U14863 (N_14863,N_13462,N_13473);
nor U14864 (N_14864,N_13390,N_13292);
nor U14865 (N_14865,N_13312,N_13257);
nor U14866 (N_14866,N_14050,N_13282);
xnor U14867 (N_14867,N_13283,N_13526);
or U14868 (N_14868,N_13941,N_13565);
nor U14869 (N_14869,N_14297,N_13788);
nand U14870 (N_14870,N_13307,N_14272);
and U14871 (N_14871,N_13557,N_14295);
nand U14872 (N_14872,N_13582,N_13672);
nor U14873 (N_14873,N_13223,N_13765);
or U14874 (N_14874,N_13382,N_13538);
nor U14875 (N_14875,N_14286,N_13980);
or U14876 (N_14876,N_13497,N_14350);
nand U14877 (N_14877,N_13634,N_13243);
nand U14878 (N_14878,N_13359,N_13519);
xor U14879 (N_14879,N_13353,N_13695);
nor U14880 (N_14880,N_13325,N_13525);
or U14881 (N_14881,N_13766,N_14098);
xnor U14882 (N_14882,N_13977,N_14343);
and U14883 (N_14883,N_13343,N_13595);
xor U14884 (N_14884,N_14310,N_13777);
nor U14885 (N_14885,N_14134,N_13318);
or U14886 (N_14886,N_13304,N_14061);
nor U14887 (N_14887,N_13913,N_13381);
or U14888 (N_14888,N_13933,N_14240);
nor U14889 (N_14889,N_13793,N_14037);
xor U14890 (N_14890,N_14143,N_13771);
xor U14891 (N_14891,N_13322,N_13891);
xor U14892 (N_14892,N_14386,N_13661);
and U14893 (N_14893,N_13778,N_13417);
or U14894 (N_14894,N_13723,N_13206);
or U14895 (N_14895,N_14125,N_14045);
and U14896 (N_14896,N_13645,N_14123);
and U14897 (N_14897,N_13321,N_13919);
xnor U14898 (N_14898,N_14356,N_13498);
and U14899 (N_14899,N_13710,N_13974);
xnor U14900 (N_14900,N_13950,N_13281);
nor U14901 (N_14901,N_13333,N_13610);
nand U14902 (N_14902,N_13963,N_13814);
nand U14903 (N_14903,N_14105,N_13250);
nand U14904 (N_14904,N_13384,N_13697);
or U14905 (N_14905,N_13606,N_14009);
xor U14906 (N_14906,N_13794,N_13659);
xnor U14907 (N_14907,N_13400,N_14312);
and U14908 (N_14908,N_13348,N_14121);
and U14909 (N_14909,N_14057,N_14224);
nor U14910 (N_14910,N_13706,N_13817);
nor U14911 (N_14911,N_13271,N_13291);
or U14912 (N_14912,N_14284,N_13663);
xor U14913 (N_14913,N_14215,N_13864);
nor U14914 (N_14914,N_13945,N_14298);
nor U14915 (N_14915,N_14303,N_13492);
nand U14916 (N_14916,N_13402,N_13486);
or U14917 (N_14917,N_14203,N_14067);
nor U14918 (N_14918,N_14394,N_13375);
nor U14919 (N_14919,N_14308,N_13370);
nand U14920 (N_14920,N_13668,N_13438);
nand U14921 (N_14921,N_13352,N_13229);
nor U14922 (N_14922,N_13835,N_14265);
or U14923 (N_14923,N_13729,N_14124);
or U14924 (N_14924,N_14257,N_14190);
and U14925 (N_14925,N_13806,N_13296);
and U14926 (N_14926,N_13235,N_13508);
nor U14927 (N_14927,N_13890,N_14358);
or U14928 (N_14928,N_13725,N_13221);
xor U14929 (N_14929,N_13578,N_13427);
and U14930 (N_14930,N_13951,N_14322);
nor U14931 (N_14931,N_13248,N_13857);
or U14932 (N_14932,N_14017,N_13756);
and U14933 (N_14933,N_13246,N_14379);
nor U14934 (N_14934,N_13895,N_13802);
and U14935 (N_14935,N_13346,N_13786);
xor U14936 (N_14936,N_13837,N_13247);
or U14937 (N_14937,N_14248,N_14174);
and U14938 (N_14938,N_13234,N_13245);
nor U14939 (N_14939,N_13962,N_13991);
nand U14940 (N_14940,N_13858,N_13537);
nand U14941 (N_14941,N_13713,N_14059);
or U14942 (N_14942,N_14396,N_13546);
xor U14943 (N_14943,N_13745,N_13512);
and U14944 (N_14944,N_13436,N_13736);
nor U14945 (N_14945,N_13275,N_13637);
or U14946 (N_14946,N_14219,N_14228);
nor U14947 (N_14947,N_13705,N_14022);
xor U14948 (N_14948,N_14081,N_13254);
nand U14949 (N_14949,N_13965,N_13463);
and U14950 (N_14950,N_14122,N_13272);
or U14951 (N_14951,N_14006,N_13908);
xor U14952 (N_14952,N_13791,N_14354);
nor U14953 (N_14953,N_13975,N_14290);
nand U14954 (N_14954,N_14319,N_14390);
xor U14955 (N_14955,N_13439,N_13779);
or U14956 (N_14956,N_13833,N_13939);
or U14957 (N_14957,N_13303,N_13896);
nand U14958 (N_14958,N_13683,N_13823);
nor U14959 (N_14959,N_14133,N_13378);
and U14960 (N_14960,N_14256,N_13701);
nor U14961 (N_14961,N_13586,N_14079);
nor U14962 (N_14962,N_13978,N_14181);
or U14963 (N_14963,N_13387,N_13911);
or U14964 (N_14964,N_14166,N_13285);
nand U14965 (N_14965,N_14053,N_13716);
nand U14966 (N_14966,N_13344,N_13612);
nand U14967 (N_14967,N_13731,N_13801);
and U14968 (N_14968,N_14281,N_13543);
nor U14969 (N_14969,N_13549,N_14087);
xor U14970 (N_14970,N_14377,N_13764);
nand U14971 (N_14971,N_13429,N_13631);
nand U14972 (N_14972,N_14026,N_13749);
and U14973 (N_14973,N_13274,N_13682);
nor U14974 (N_14974,N_13410,N_14028);
xnor U14975 (N_14975,N_13345,N_13528);
nor U14976 (N_14976,N_13523,N_13935);
and U14977 (N_14977,N_13772,N_14237);
nor U14978 (N_14978,N_14335,N_13953);
and U14979 (N_14979,N_13472,N_13825);
nand U14980 (N_14980,N_14171,N_14326);
nand U14981 (N_14981,N_13577,N_14194);
or U14982 (N_14982,N_13613,N_14159);
nor U14983 (N_14983,N_13994,N_14018);
or U14984 (N_14984,N_13665,N_14184);
nand U14985 (N_14985,N_13866,N_14140);
and U14986 (N_14986,N_13702,N_13862);
xor U14987 (N_14987,N_14302,N_13618);
xor U14988 (N_14988,N_13698,N_14288);
or U14989 (N_14989,N_14258,N_13803);
or U14990 (N_14990,N_13881,N_13554);
and U14991 (N_14991,N_13737,N_14230);
nand U14992 (N_14992,N_13623,N_13568);
and U14993 (N_14993,N_13667,N_13615);
nand U14994 (N_14994,N_13997,N_14255);
or U14995 (N_14995,N_14381,N_13326);
nand U14996 (N_14996,N_13998,N_13259);
nand U14997 (N_14997,N_14201,N_13841);
and U14998 (N_14998,N_14145,N_13652);
nand U14999 (N_14999,N_14076,N_14253);
nand U15000 (N_15000,N_14336,N_13368);
nor U15001 (N_15001,N_13813,N_13332);
nor U15002 (N_15002,N_13626,N_13366);
nor U15003 (N_15003,N_14017,N_13407);
xnor U15004 (N_15004,N_13774,N_13624);
xnor U15005 (N_15005,N_13698,N_13990);
nor U15006 (N_15006,N_14255,N_13762);
xor U15007 (N_15007,N_14239,N_13639);
or U15008 (N_15008,N_13742,N_14098);
nor U15009 (N_15009,N_13863,N_14132);
and U15010 (N_15010,N_13436,N_13920);
nor U15011 (N_15011,N_13960,N_14176);
nand U15012 (N_15012,N_14033,N_13448);
nor U15013 (N_15013,N_13973,N_14053);
or U15014 (N_15014,N_13480,N_13580);
and U15015 (N_15015,N_14186,N_13886);
nand U15016 (N_15016,N_13372,N_13397);
nand U15017 (N_15017,N_13826,N_14245);
nor U15018 (N_15018,N_14360,N_14249);
and U15019 (N_15019,N_13488,N_14376);
or U15020 (N_15020,N_13855,N_13500);
xor U15021 (N_15021,N_13467,N_13718);
or U15022 (N_15022,N_14000,N_13779);
nand U15023 (N_15023,N_14172,N_14061);
or U15024 (N_15024,N_13430,N_13887);
or U15025 (N_15025,N_13206,N_13752);
or U15026 (N_15026,N_14153,N_14074);
or U15027 (N_15027,N_14063,N_14354);
xor U15028 (N_15028,N_13433,N_13810);
nand U15029 (N_15029,N_13214,N_14194);
or U15030 (N_15030,N_13308,N_13460);
xor U15031 (N_15031,N_14149,N_14364);
nor U15032 (N_15032,N_13208,N_14252);
nor U15033 (N_15033,N_13227,N_13695);
nand U15034 (N_15034,N_13557,N_14281);
nor U15035 (N_15035,N_13702,N_13951);
nor U15036 (N_15036,N_14206,N_13783);
nand U15037 (N_15037,N_13637,N_13882);
and U15038 (N_15038,N_13464,N_14147);
xnor U15039 (N_15039,N_13927,N_13262);
xnor U15040 (N_15040,N_13270,N_14383);
or U15041 (N_15041,N_13420,N_14081);
and U15042 (N_15042,N_13899,N_13459);
nand U15043 (N_15043,N_13624,N_14288);
or U15044 (N_15044,N_13699,N_14003);
or U15045 (N_15045,N_13413,N_14167);
and U15046 (N_15046,N_14375,N_14292);
and U15047 (N_15047,N_13948,N_13662);
nand U15048 (N_15048,N_13331,N_14101);
or U15049 (N_15049,N_14104,N_14263);
nand U15050 (N_15050,N_14025,N_13574);
nor U15051 (N_15051,N_13834,N_13212);
xor U15052 (N_15052,N_13331,N_13504);
and U15053 (N_15053,N_13695,N_13803);
nand U15054 (N_15054,N_14119,N_14134);
nor U15055 (N_15055,N_13809,N_13877);
xnor U15056 (N_15056,N_13898,N_13923);
nand U15057 (N_15057,N_14290,N_14014);
xor U15058 (N_15058,N_13862,N_13364);
nor U15059 (N_15059,N_13942,N_14138);
or U15060 (N_15060,N_13500,N_13360);
xnor U15061 (N_15061,N_13425,N_14046);
nor U15062 (N_15062,N_13904,N_13481);
or U15063 (N_15063,N_13810,N_13618);
nand U15064 (N_15064,N_13819,N_13582);
nor U15065 (N_15065,N_13755,N_13982);
and U15066 (N_15066,N_14172,N_13734);
and U15067 (N_15067,N_13741,N_14136);
and U15068 (N_15068,N_13915,N_14114);
nor U15069 (N_15069,N_14315,N_14378);
nor U15070 (N_15070,N_13749,N_13750);
nor U15071 (N_15071,N_13397,N_14166);
nand U15072 (N_15072,N_13655,N_13698);
or U15073 (N_15073,N_13667,N_14019);
or U15074 (N_15074,N_13685,N_13648);
and U15075 (N_15075,N_14211,N_13790);
nand U15076 (N_15076,N_13342,N_13260);
nor U15077 (N_15077,N_13571,N_13894);
nand U15078 (N_15078,N_14267,N_13977);
or U15079 (N_15079,N_13374,N_13876);
nor U15080 (N_15080,N_13503,N_13627);
xnor U15081 (N_15081,N_13924,N_13945);
or U15082 (N_15082,N_13553,N_14270);
or U15083 (N_15083,N_14378,N_14039);
xor U15084 (N_15084,N_13210,N_13382);
or U15085 (N_15085,N_13941,N_13530);
and U15086 (N_15086,N_14372,N_13670);
nand U15087 (N_15087,N_13581,N_13441);
and U15088 (N_15088,N_13728,N_13882);
nand U15089 (N_15089,N_14017,N_13801);
xnor U15090 (N_15090,N_13938,N_13492);
xnor U15091 (N_15091,N_13396,N_13572);
nand U15092 (N_15092,N_13391,N_13454);
or U15093 (N_15093,N_14070,N_13667);
nand U15094 (N_15094,N_13773,N_13271);
nand U15095 (N_15095,N_13575,N_13984);
nor U15096 (N_15096,N_13337,N_13492);
and U15097 (N_15097,N_13350,N_14272);
nor U15098 (N_15098,N_13954,N_13714);
and U15099 (N_15099,N_13253,N_13751);
nand U15100 (N_15100,N_14342,N_13318);
and U15101 (N_15101,N_13207,N_14350);
or U15102 (N_15102,N_14004,N_13326);
and U15103 (N_15103,N_13362,N_13982);
xor U15104 (N_15104,N_14372,N_13675);
and U15105 (N_15105,N_14277,N_14014);
nand U15106 (N_15106,N_13867,N_13883);
nor U15107 (N_15107,N_13463,N_13230);
and U15108 (N_15108,N_13536,N_13861);
and U15109 (N_15109,N_14057,N_14129);
or U15110 (N_15110,N_13771,N_13217);
nor U15111 (N_15111,N_13301,N_14253);
xor U15112 (N_15112,N_13511,N_14119);
or U15113 (N_15113,N_13282,N_13887);
or U15114 (N_15114,N_13788,N_13273);
xnor U15115 (N_15115,N_13761,N_13806);
xor U15116 (N_15116,N_14022,N_13302);
nor U15117 (N_15117,N_14276,N_13393);
and U15118 (N_15118,N_14138,N_13393);
xor U15119 (N_15119,N_13873,N_13953);
or U15120 (N_15120,N_13240,N_13687);
nand U15121 (N_15121,N_13990,N_13646);
nor U15122 (N_15122,N_14176,N_13865);
nor U15123 (N_15123,N_14246,N_13647);
nor U15124 (N_15124,N_14098,N_13842);
xnor U15125 (N_15125,N_14133,N_14227);
nor U15126 (N_15126,N_13233,N_14010);
or U15127 (N_15127,N_13300,N_13279);
nor U15128 (N_15128,N_13217,N_13311);
nor U15129 (N_15129,N_13779,N_13348);
nor U15130 (N_15130,N_14020,N_14103);
nor U15131 (N_15131,N_14291,N_13208);
xor U15132 (N_15132,N_13668,N_14219);
or U15133 (N_15133,N_13610,N_13575);
xnor U15134 (N_15134,N_13379,N_13797);
nor U15135 (N_15135,N_13358,N_13731);
xor U15136 (N_15136,N_13261,N_14188);
or U15137 (N_15137,N_14296,N_13544);
and U15138 (N_15138,N_14323,N_13789);
and U15139 (N_15139,N_13954,N_13533);
and U15140 (N_15140,N_13699,N_13836);
and U15141 (N_15141,N_13620,N_13571);
xor U15142 (N_15142,N_13241,N_14112);
or U15143 (N_15143,N_14320,N_13770);
xnor U15144 (N_15144,N_13996,N_13390);
xor U15145 (N_15145,N_14166,N_13522);
nor U15146 (N_15146,N_13940,N_13863);
xor U15147 (N_15147,N_13604,N_13873);
xor U15148 (N_15148,N_13902,N_13993);
or U15149 (N_15149,N_14300,N_13844);
or U15150 (N_15150,N_14089,N_13782);
nor U15151 (N_15151,N_13931,N_13378);
xor U15152 (N_15152,N_13635,N_13742);
nor U15153 (N_15153,N_13768,N_13615);
nor U15154 (N_15154,N_13514,N_14000);
and U15155 (N_15155,N_13667,N_13753);
and U15156 (N_15156,N_13256,N_13217);
xor U15157 (N_15157,N_13633,N_13911);
xor U15158 (N_15158,N_13990,N_14044);
or U15159 (N_15159,N_13797,N_13856);
nor U15160 (N_15160,N_13425,N_13899);
xnor U15161 (N_15161,N_13808,N_13393);
nand U15162 (N_15162,N_14052,N_13972);
and U15163 (N_15163,N_13799,N_13475);
and U15164 (N_15164,N_13312,N_13330);
xnor U15165 (N_15165,N_13265,N_14315);
nand U15166 (N_15166,N_13686,N_13804);
nand U15167 (N_15167,N_13737,N_13675);
or U15168 (N_15168,N_13202,N_13508);
and U15169 (N_15169,N_13288,N_14273);
xor U15170 (N_15170,N_14325,N_13528);
xor U15171 (N_15171,N_14253,N_13722);
or U15172 (N_15172,N_13355,N_13646);
xor U15173 (N_15173,N_13699,N_14023);
and U15174 (N_15174,N_14178,N_13856);
and U15175 (N_15175,N_13284,N_13525);
nor U15176 (N_15176,N_13560,N_13974);
or U15177 (N_15177,N_13640,N_14140);
xnor U15178 (N_15178,N_13993,N_14067);
xnor U15179 (N_15179,N_13966,N_13950);
nor U15180 (N_15180,N_13331,N_13484);
nor U15181 (N_15181,N_13281,N_14086);
or U15182 (N_15182,N_13859,N_13564);
or U15183 (N_15183,N_14041,N_13263);
and U15184 (N_15184,N_14187,N_13691);
and U15185 (N_15185,N_13328,N_13652);
and U15186 (N_15186,N_13564,N_13453);
and U15187 (N_15187,N_13494,N_13282);
xnor U15188 (N_15188,N_13683,N_13971);
or U15189 (N_15189,N_14259,N_13542);
or U15190 (N_15190,N_14106,N_13794);
xor U15191 (N_15191,N_14190,N_13716);
and U15192 (N_15192,N_13763,N_13430);
nand U15193 (N_15193,N_13274,N_14188);
or U15194 (N_15194,N_14327,N_13905);
nor U15195 (N_15195,N_14093,N_13521);
or U15196 (N_15196,N_14396,N_13457);
or U15197 (N_15197,N_13740,N_13412);
xnor U15198 (N_15198,N_13681,N_14251);
xor U15199 (N_15199,N_13214,N_13908);
and U15200 (N_15200,N_14241,N_14062);
nand U15201 (N_15201,N_13220,N_14366);
nand U15202 (N_15202,N_13991,N_13610);
xnor U15203 (N_15203,N_13273,N_13664);
xnor U15204 (N_15204,N_13931,N_13768);
xor U15205 (N_15205,N_14352,N_13882);
nand U15206 (N_15206,N_13305,N_13833);
nand U15207 (N_15207,N_13490,N_13626);
and U15208 (N_15208,N_13808,N_14201);
xor U15209 (N_15209,N_13768,N_14113);
nand U15210 (N_15210,N_14233,N_14132);
nand U15211 (N_15211,N_13592,N_13723);
or U15212 (N_15212,N_13392,N_13645);
and U15213 (N_15213,N_13488,N_13244);
xor U15214 (N_15214,N_14158,N_14178);
nor U15215 (N_15215,N_13642,N_14244);
nor U15216 (N_15216,N_13672,N_13795);
nor U15217 (N_15217,N_13752,N_14333);
xnor U15218 (N_15218,N_13233,N_13586);
nand U15219 (N_15219,N_13379,N_14209);
or U15220 (N_15220,N_14045,N_14077);
xnor U15221 (N_15221,N_14395,N_13285);
nor U15222 (N_15222,N_13916,N_14322);
nand U15223 (N_15223,N_14371,N_14227);
xnor U15224 (N_15224,N_14125,N_14155);
and U15225 (N_15225,N_13475,N_14074);
and U15226 (N_15226,N_13737,N_14219);
nor U15227 (N_15227,N_14125,N_14211);
and U15228 (N_15228,N_13904,N_13472);
xor U15229 (N_15229,N_13594,N_14300);
xnor U15230 (N_15230,N_14021,N_13210);
and U15231 (N_15231,N_13795,N_13478);
nand U15232 (N_15232,N_14099,N_14370);
and U15233 (N_15233,N_13384,N_13240);
nand U15234 (N_15234,N_13272,N_13253);
nand U15235 (N_15235,N_13278,N_13721);
xor U15236 (N_15236,N_13821,N_13737);
nor U15237 (N_15237,N_13247,N_14152);
nand U15238 (N_15238,N_13257,N_14325);
or U15239 (N_15239,N_13671,N_13787);
and U15240 (N_15240,N_13498,N_13203);
xor U15241 (N_15241,N_13453,N_13458);
or U15242 (N_15242,N_13725,N_13636);
nand U15243 (N_15243,N_13843,N_13298);
nor U15244 (N_15244,N_13331,N_13796);
xor U15245 (N_15245,N_13374,N_13273);
and U15246 (N_15246,N_14351,N_13854);
and U15247 (N_15247,N_13279,N_14252);
xnor U15248 (N_15248,N_14187,N_14058);
nand U15249 (N_15249,N_13494,N_13920);
nor U15250 (N_15250,N_13805,N_13381);
nand U15251 (N_15251,N_13992,N_13649);
xor U15252 (N_15252,N_13985,N_13773);
nor U15253 (N_15253,N_14159,N_13788);
and U15254 (N_15254,N_13353,N_14208);
nand U15255 (N_15255,N_14365,N_13215);
and U15256 (N_15256,N_13318,N_14215);
and U15257 (N_15257,N_13925,N_14167);
or U15258 (N_15258,N_14313,N_14284);
nor U15259 (N_15259,N_13839,N_13745);
and U15260 (N_15260,N_14118,N_14002);
nand U15261 (N_15261,N_13604,N_13508);
and U15262 (N_15262,N_14163,N_13928);
nand U15263 (N_15263,N_13711,N_13987);
and U15264 (N_15264,N_14371,N_14099);
nor U15265 (N_15265,N_13690,N_13549);
nor U15266 (N_15266,N_14253,N_13758);
xnor U15267 (N_15267,N_14153,N_13832);
nor U15268 (N_15268,N_13592,N_13525);
xnor U15269 (N_15269,N_13692,N_13359);
xor U15270 (N_15270,N_13665,N_14192);
nor U15271 (N_15271,N_13440,N_13713);
or U15272 (N_15272,N_14116,N_13897);
and U15273 (N_15273,N_13452,N_13966);
xnor U15274 (N_15274,N_13902,N_13947);
nand U15275 (N_15275,N_14339,N_14368);
xor U15276 (N_15276,N_14337,N_14127);
xor U15277 (N_15277,N_13637,N_13300);
nand U15278 (N_15278,N_13477,N_13952);
or U15279 (N_15279,N_13902,N_14144);
or U15280 (N_15280,N_13670,N_14145);
nand U15281 (N_15281,N_13437,N_13800);
or U15282 (N_15282,N_13411,N_13726);
xnor U15283 (N_15283,N_14345,N_13213);
nor U15284 (N_15284,N_13694,N_13892);
xor U15285 (N_15285,N_13997,N_13533);
nand U15286 (N_15286,N_14183,N_13333);
nor U15287 (N_15287,N_14252,N_13843);
nor U15288 (N_15288,N_13904,N_13894);
nand U15289 (N_15289,N_14036,N_13488);
and U15290 (N_15290,N_13596,N_14012);
xor U15291 (N_15291,N_13929,N_14076);
or U15292 (N_15292,N_13314,N_13445);
nand U15293 (N_15293,N_13416,N_13644);
and U15294 (N_15294,N_13388,N_13259);
xor U15295 (N_15295,N_14314,N_14232);
nand U15296 (N_15296,N_14262,N_13543);
nor U15297 (N_15297,N_13440,N_14197);
nor U15298 (N_15298,N_14083,N_13840);
nor U15299 (N_15299,N_13228,N_13380);
nand U15300 (N_15300,N_14382,N_14163);
or U15301 (N_15301,N_14383,N_13940);
nand U15302 (N_15302,N_13315,N_13538);
nor U15303 (N_15303,N_14335,N_14270);
nor U15304 (N_15304,N_14128,N_13944);
nor U15305 (N_15305,N_13703,N_13541);
nor U15306 (N_15306,N_13274,N_13420);
and U15307 (N_15307,N_13241,N_14320);
nor U15308 (N_15308,N_13289,N_14121);
or U15309 (N_15309,N_13485,N_14221);
xnor U15310 (N_15310,N_13293,N_13433);
nand U15311 (N_15311,N_14357,N_13910);
xnor U15312 (N_15312,N_14346,N_13914);
xor U15313 (N_15313,N_14396,N_13479);
nand U15314 (N_15314,N_14162,N_13936);
xor U15315 (N_15315,N_13674,N_13906);
or U15316 (N_15316,N_13601,N_13248);
or U15317 (N_15317,N_14228,N_13716);
and U15318 (N_15318,N_13390,N_13755);
or U15319 (N_15319,N_13317,N_13609);
and U15320 (N_15320,N_13762,N_14170);
nand U15321 (N_15321,N_13824,N_13605);
nand U15322 (N_15322,N_13302,N_13946);
xnor U15323 (N_15323,N_14201,N_13768);
or U15324 (N_15324,N_13481,N_13519);
nand U15325 (N_15325,N_13983,N_14371);
and U15326 (N_15326,N_14088,N_14328);
xnor U15327 (N_15327,N_13689,N_14369);
or U15328 (N_15328,N_14267,N_14340);
and U15329 (N_15329,N_13732,N_14165);
nand U15330 (N_15330,N_13381,N_13889);
nor U15331 (N_15331,N_13718,N_13491);
xor U15332 (N_15332,N_14200,N_13634);
or U15333 (N_15333,N_14158,N_13731);
xnor U15334 (N_15334,N_13996,N_14158);
xnor U15335 (N_15335,N_13844,N_13289);
xnor U15336 (N_15336,N_13947,N_13830);
and U15337 (N_15337,N_13806,N_14190);
xor U15338 (N_15338,N_14201,N_14067);
or U15339 (N_15339,N_14043,N_14353);
or U15340 (N_15340,N_14274,N_13443);
or U15341 (N_15341,N_13225,N_13570);
nor U15342 (N_15342,N_13559,N_13296);
nand U15343 (N_15343,N_14047,N_14122);
and U15344 (N_15344,N_14399,N_13834);
or U15345 (N_15345,N_13653,N_14152);
or U15346 (N_15346,N_13710,N_13818);
nand U15347 (N_15347,N_13583,N_13563);
nor U15348 (N_15348,N_13289,N_14040);
and U15349 (N_15349,N_13913,N_14108);
nand U15350 (N_15350,N_13736,N_14232);
and U15351 (N_15351,N_13823,N_13635);
xnor U15352 (N_15352,N_14365,N_14013);
or U15353 (N_15353,N_13484,N_14311);
and U15354 (N_15354,N_13253,N_14046);
or U15355 (N_15355,N_14291,N_14014);
nand U15356 (N_15356,N_13571,N_13816);
or U15357 (N_15357,N_14304,N_14358);
nor U15358 (N_15358,N_13566,N_14226);
and U15359 (N_15359,N_13403,N_13511);
and U15360 (N_15360,N_13704,N_13235);
or U15361 (N_15361,N_13856,N_14035);
nor U15362 (N_15362,N_13406,N_13410);
and U15363 (N_15363,N_13987,N_13270);
or U15364 (N_15364,N_13620,N_14099);
and U15365 (N_15365,N_14133,N_14084);
nand U15366 (N_15366,N_13859,N_13613);
or U15367 (N_15367,N_13990,N_13654);
nand U15368 (N_15368,N_14203,N_14086);
xor U15369 (N_15369,N_13676,N_14097);
or U15370 (N_15370,N_13302,N_14075);
xnor U15371 (N_15371,N_13663,N_13726);
or U15372 (N_15372,N_13750,N_13380);
xnor U15373 (N_15373,N_14384,N_13430);
and U15374 (N_15374,N_13312,N_13272);
or U15375 (N_15375,N_13905,N_13498);
or U15376 (N_15376,N_13609,N_13435);
xnor U15377 (N_15377,N_14383,N_13839);
xor U15378 (N_15378,N_13280,N_13931);
nand U15379 (N_15379,N_14190,N_14001);
and U15380 (N_15380,N_13915,N_13633);
and U15381 (N_15381,N_13981,N_13222);
nor U15382 (N_15382,N_14201,N_13207);
nor U15383 (N_15383,N_14381,N_13991);
nand U15384 (N_15384,N_14054,N_13923);
or U15385 (N_15385,N_13435,N_13816);
or U15386 (N_15386,N_13270,N_13618);
and U15387 (N_15387,N_13523,N_14366);
and U15388 (N_15388,N_14069,N_13970);
nor U15389 (N_15389,N_14367,N_14166);
or U15390 (N_15390,N_13820,N_13985);
and U15391 (N_15391,N_13764,N_14311);
or U15392 (N_15392,N_14342,N_13861);
or U15393 (N_15393,N_13395,N_14230);
xnor U15394 (N_15394,N_13273,N_14204);
and U15395 (N_15395,N_13335,N_14300);
xor U15396 (N_15396,N_13849,N_13602);
nand U15397 (N_15397,N_13676,N_13321);
or U15398 (N_15398,N_13232,N_13247);
or U15399 (N_15399,N_13863,N_13831);
nor U15400 (N_15400,N_13790,N_13393);
nor U15401 (N_15401,N_14076,N_14198);
nor U15402 (N_15402,N_13482,N_14027);
nand U15403 (N_15403,N_13859,N_14178);
or U15404 (N_15404,N_14306,N_14362);
xnor U15405 (N_15405,N_14185,N_14283);
nand U15406 (N_15406,N_13382,N_14044);
nor U15407 (N_15407,N_14139,N_13283);
and U15408 (N_15408,N_14232,N_13395);
and U15409 (N_15409,N_13969,N_13826);
nor U15410 (N_15410,N_14031,N_14319);
nand U15411 (N_15411,N_13951,N_14146);
nand U15412 (N_15412,N_13968,N_13737);
nor U15413 (N_15413,N_13695,N_13809);
nand U15414 (N_15414,N_13805,N_14394);
nand U15415 (N_15415,N_13811,N_14211);
nor U15416 (N_15416,N_13691,N_13767);
or U15417 (N_15417,N_13399,N_14065);
or U15418 (N_15418,N_13817,N_14047);
or U15419 (N_15419,N_13831,N_13955);
nor U15420 (N_15420,N_14326,N_13232);
or U15421 (N_15421,N_13760,N_13484);
nor U15422 (N_15422,N_13912,N_14000);
xor U15423 (N_15423,N_13422,N_13725);
and U15424 (N_15424,N_14389,N_13722);
nor U15425 (N_15425,N_14172,N_13652);
xnor U15426 (N_15426,N_13209,N_13307);
xor U15427 (N_15427,N_14278,N_13560);
nor U15428 (N_15428,N_13725,N_13697);
nand U15429 (N_15429,N_13369,N_13790);
xor U15430 (N_15430,N_13947,N_13758);
xnor U15431 (N_15431,N_14392,N_13323);
and U15432 (N_15432,N_14241,N_13551);
or U15433 (N_15433,N_14098,N_13215);
nand U15434 (N_15434,N_13944,N_13687);
nand U15435 (N_15435,N_13873,N_14249);
nor U15436 (N_15436,N_13511,N_13223);
xnor U15437 (N_15437,N_14103,N_14104);
or U15438 (N_15438,N_13247,N_14142);
xnor U15439 (N_15439,N_13906,N_14121);
and U15440 (N_15440,N_14274,N_14289);
nor U15441 (N_15441,N_13689,N_13819);
nand U15442 (N_15442,N_14170,N_13784);
or U15443 (N_15443,N_14316,N_14137);
or U15444 (N_15444,N_14322,N_13528);
xor U15445 (N_15445,N_13514,N_13634);
or U15446 (N_15446,N_13932,N_14266);
xnor U15447 (N_15447,N_13498,N_13583);
xor U15448 (N_15448,N_14249,N_13796);
nor U15449 (N_15449,N_13242,N_13759);
and U15450 (N_15450,N_13603,N_14347);
nor U15451 (N_15451,N_14267,N_13313);
nand U15452 (N_15452,N_13302,N_13408);
nand U15453 (N_15453,N_14218,N_13678);
or U15454 (N_15454,N_14038,N_13230);
nand U15455 (N_15455,N_13822,N_13356);
nand U15456 (N_15456,N_14308,N_13288);
nor U15457 (N_15457,N_14197,N_13619);
nand U15458 (N_15458,N_13400,N_14178);
xor U15459 (N_15459,N_13388,N_13429);
and U15460 (N_15460,N_14346,N_13261);
xnor U15461 (N_15461,N_14218,N_14106);
nand U15462 (N_15462,N_13254,N_14344);
nor U15463 (N_15463,N_14159,N_13813);
or U15464 (N_15464,N_14054,N_14219);
nand U15465 (N_15465,N_13695,N_14100);
nor U15466 (N_15466,N_13681,N_13749);
and U15467 (N_15467,N_13880,N_13627);
nand U15468 (N_15468,N_13980,N_13576);
xor U15469 (N_15469,N_13656,N_13786);
and U15470 (N_15470,N_13808,N_13383);
nor U15471 (N_15471,N_13718,N_13612);
or U15472 (N_15472,N_14178,N_13963);
nor U15473 (N_15473,N_13351,N_13900);
and U15474 (N_15474,N_14286,N_13576);
nor U15475 (N_15475,N_13309,N_14283);
nand U15476 (N_15476,N_14275,N_13458);
nand U15477 (N_15477,N_14139,N_13671);
and U15478 (N_15478,N_13464,N_13847);
or U15479 (N_15479,N_14259,N_14389);
nand U15480 (N_15480,N_13397,N_14031);
nand U15481 (N_15481,N_13909,N_14011);
xor U15482 (N_15482,N_13277,N_13377);
nand U15483 (N_15483,N_13526,N_13233);
or U15484 (N_15484,N_13947,N_13668);
or U15485 (N_15485,N_13760,N_13574);
nand U15486 (N_15486,N_13520,N_13902);
or U15487 (N_15487,N_13582,N_13719);
or U15488 (N_15488,N_13745,N_13845);
nor U15489 (N_15489,N_13242,N_13684);
or U15490 (N_15490,N_13329,N_13485);
xor U15491 (N_15491,N_13548,N_13925);
and U15492 (N_15492,N_14335,N_14201);
xor U15493 (N_15493,N_13787,N_13932);
xor U15494 (N_15494,N_14079,N_13416);
xor U15495 (N_15495,N_13323,N_13629);
or U15496 (N_15496,N_14138,N_14068);
nor U15497 (N_15497,N_14161,N_13454);
nand U15498 (N_15498,N_13710,N_14210);
nand U15499 (N_15499,N_14225,N_13612);
nor U15500 (N_15500,N_14365,N_14240);
or U15501 (N_15501,N_13377,N_14316);
or U15502 (N_15502,N_14175,N_13512);
xnor U15503 (N_15503,N_14243,N_13874);
nor U15504 (N_15504,N_13521,N_13512);
or U15505 (N_15505,N_13872,N_13628);
xor U15506 (N_15506,N_14319,N_14087);
xor U15507 (N_15507,N_13316,N_13702);
nor U15508 (N_15508,N_13231,N_13780);
or U15509 (N_15509,N_13529,N_14098);
nor U15510 (N_15510,N_14386,N_13920);
nand U15511 (N_15511,N_13205,N_13799);
or U15512 (N_15512,N_14014,N_13426);
nand U15513 (N_15513,N_13572,N_13980);
nor U15514 (N_15514,N_14188,N_13852);
nand U15515 (N_15515,N_13809,N_13980);
nand U15516 (N_15516,N_13554,N_13889);
or U15517 (N_15517,N_13963,N_13220);
nor U15518 (N_15518,N_13478,N_13618);
or U15519 (N_15519,N_13224,N_13255);
nor U15520 (N_15520,N_13783,N_13632);
nor U15521 (N_15521,N_13494,N_13817);
xnor U15522 (N_15522,N_13750,N_13780);
and U15523 (N_15523,N_13323,N_14054);
nor U15524 (N_15524,N_13620,N_14351);
nor U15525 (N_15525,N_13746,N_14267);
and U15526 (N_15526,N_13703,N_13244);
and U15527 (N_15527,N_14018,N_13892);
and U15528 (N_15528,N_14147,N_13975);
or U15529 (N_15529,N_13891,N_13281);
or U15530 (N_15530,N_14380,N_13741);
or U15531 (N_15531,N_13415,N_13743);
and U15532 (N_15532,N_13618,N_14288);
nand U15533 (N_15533,N_13698,N_13434);
or U15534 (N_15534,N_13293,N_14169);
or U15535 (N_15535,N_13667,N_13447);
xnor U15536 (N_15536,N_13924,N_13297);
xnor U15537 (N_15537,N_14078,N_14398);
or U15538 (N_15538,N_14266,N_13403);
nand U15539 (N_15539,N_14045,N_14144);
nand U15540 (N_15540,N_13214,N_13359);
nand U15541 (N_15541,N_14281,N_13678);
and U15542 (N_15542,N_13599,N_13959);
nor U15543 (N_15543,N_13377,N_13676);
or U15544 (N_15544,N_13610,N_13449);
xor U15545 (N_15545,N_13867,N_14120);
or U15546 (N_15546,N_13550,N_13408);
or U15547 (N_15547,N_13793,N_13739);
nand U15548 (N_15548,N_13688,N_14172);
nor U15549 (N_15549,N_14205,N_13336);
and U15550 (N_15550,N_13750,N_13340);
nor U15551 (N_15551,N_14294,N_13303);
nand U15552 (N_15552,N_13356,N_14015);
nor U15553 (N_15553,N_13837,N_13786);
or U15554 (N_15554,N_13498,N_13455);
or U15555 (N_15555,N_14395,N_14335);
nor U15556 (N_15556,N_13928,N_14076);
nor U15557 (N_15557,N_13543,N_13874);
and U15558 (N_15558,N_13784,N_14091);
and U15559 (N_15559,N_13956,N_14232);
nor U15560 (N_15560,N_13703,N_14398);
or U15561 (N_15561,N_13857,N_14062);
nand U15562 (N_15562,N_13596,N_13778);
nand U15563 (N_15563,N_13850,N_13715);
or U15564 (N_15564,N_13591,N_13724);
nand U15565 (N_15565,N_13666,N_14167);
xnor U15566 (N_15566,N_13871,N_13874);
xor U15567 (N_15567,N_13464,N_13250);
nor U15568 (N_15568,N_13829,N_13225);
nor U15569 (N_15569,N_14171,N_13696);
nand U15570 (N_15570,N_14044,N_14166);
nand U15571 (N_15571,N_13638,N_13981);
nor U15572 (N_15572,N_13679,N_14343);
or U15573 (N_15573,N_13602,N_13977);
and U15574 (N_15574,N_13766,N_13579);
xnor U15575 (N_15575,N_14222,N_13612);
nor U15576 (N_15576,N_13949,N_13642);
nand U15577 (N_15577,N_13793,N_13665);
and U15578 (N_15578,N_13652,N_13862);
or U15579 (N_15579,N_14265,N_13407);
and U15580 (N_15580,N_13709,N_13736);
nor U15581 (N_15581,N_13606,N_14394);
nand U15582 (N_15582,N_13347,N_14173);
nand U15583 (N_15583,N_13223,N_14102);
or U15584 (N_15584,N_13754,N_14115);
xor U15585 (N_15585,N_14299,N_13923);
xor U15586 (N_15586,N_13690,N_13975);
nor U15587 (N_15587,N_13514,N_13724);
nand U15588 (N_15588,N_13988,N_13804);
nor U15589 (N_15589,N_13308,N_13647);
xor U15590 (N_15590,N_14262,N_13218);
nor U15591 (N_15591,N_14048,N_14028);
and U15592 (N_15592,N_13647,N_13377);
and U15593 (N_15593,N_14195,N_13555);
xnor U15594 (N_15594,N_14189,N_13336);
and U15595 (N_15595,N_13442,N_13613);
and U15596 (N_15596,N_13510,N_13314);
nand U15597 (N_15597,N_13650,N_13570);
nand U15598 (N_15598,N_14246,N_14028);
and U15599 (N_15599,N_13310,N_14274);
nor U15600 (N_15600,N_14494,N_14432);
or U15601 (N_15601,N_14515,N_15030);
nor U15602 (N_15602,N_14595,N_15131);
xor U15603 (N_15603,N_15305,N_15277);
or U15604 (N_15604,N_14799,N_14987);
nor U15605 (N_15605,N_14623,N_14563);
xnor U15606 (N_15606,N_14628,N_14483);
nand U15607 (N_15607,N_15302,N_14589);
xor U15608 (N_15608,N_15429,N_14410);
nand U15609 (N_15609,N_14531,N_15406);
or U15610 (N_15610,N_15110,N_15402);
or U15611 (N_15611,N_14653,N_14562);
and U15612 (N_15612,N_15467,N_15171);
or U15613 (N_15613,N_15437,N_14754);
nor U15614 (N_15614,N_15368,N_15235);
and U15615 (N_15615,N_14619,N_14752);
or U15616 (N_15616,N_15136,N_15345);
or U15617 (N_15617,N_15569,N_15330);
and U15618 (N_15618,N_14618,N_14892);
nor U15619 (N_15619,N_15562,N_14724);
or U15620 (N_15620,N_14742,N_14681);
nand U15621 (N_15621,N_14818,N_14981);
xor U15622 (N_15622,N_14812,N_15064);
xor U15623 (N_15623,N_15481,N_15009);
nand U15624 (N_15624,N_15320,N_15108);
nor U15625 (N_15625,N_14471,N_14973);
xor U15626 (N_15626,N_14509,N_15249);
nand U15627 (N_15627,N_15439,N_15325);
or U15628 (N_15628,N_15570,N_14641);
xor U15629 (N_15629,N_15237,N_14974);
nor U15630 (N_15630,N_15113,N_14686);
and U15631 (N_15631,N_14517,N_14580);
nor U15632 (N_15632,N_15232,N_15291);
xor U15633 (N_15633,N_14729,N_14978);
and U15634 (N_15634,N_14878,N_14888);
nor U15635 (N_15635,N_14961,N_15251);
and U15636 (N_15636,N_14725,N_14648);
nand U15637 (N_15637,N_15520,N_14583);
xnor U15638 (N_15638,N_14427,N_15488);
and U15639 (N_15639,N_14841,N_15304);
or U15640 (N_15640,N_15287,N_15041);
nor U15641 (N_15641,N_15040,N_15264);
nor U15642 (N_15642,N_14667,N_15270);
or U15643 (N_15643,N_15262,N_15242);
xnor U15644 (N_15644,N_14672,N_15024);
and U15645 (N_15645,N_14863,N_15065);
or U15646 (N_15646,N_15054,N_14657);
and U15647 (N_15647,N_14663,N_14552);
and U15648 (N_15648,N_14920,N_14645);
nand U15649 (N_15649,N_15373,N_15124);
nand U15650 (N_15650,N_15244,N_14430);
xor U15651 (N_15651,N_15226,N_15410);
nor U15652 (N_15652,N_15346,N_15573);
xor U15653 (N_15653,N_15228,N_15576);
nand U15654 (N_15654,N_14451,N_15478);
nor U15655 (N_15655,N_15190,N_15128);
or U15656 (N_15656,N_15545,N_15407);
nand U15657 (N_15657,N_14976,N_15152);
or U15658 (N_15658,N_14727,N_14824);
nand U15659 (N_15659,N_14439,N_14424);
and U15660 (N_15660,N_14640,N_14798);
nand U15661 (N_15661,N_14450,N_14579);
nand U15662 (N_15662,N_14869,N_15279);
and U15663 (N_15663,N_14594,N_15227);
nor U15664 (N_15664,N_14567,N_14776);
and U15665 (N_15665,N_15428,N_14834);
xor U15666 (N_15666,N_15360,N_15380);
nor U15667 (N_15667,N_15038,N_14791);
xnor U15668 (N_15668,N_15435,N_15280);
and U15669 (N_15669,N_15087,N_15082);
xor U15670 (N_15670,N_14982,N_15352);
nand U15671 (N_15671,N_14990,N_15204);
nor U15672 (N_15672,N_15475,N_15013);
nand U15673 (N_15673,N_15103,N_15512);
and U15674 (N_15674,N_14960,N_15544);
nand U15675 (N_15675,N_14435,N_15284);
nand U15676 (N_15676,N_15229,N_15115);
or U15677 (N_15677,N_14484,N_15278);
or U15678 (N_15678,N_15460,N_15076);
nand U15679 (N_15679,N_15252,N_14576);
nor U15680 (N_15680,N_14661,N_15586);
nor U15681 (N_15681,N_14709,N_15462);
nor U15682 (N_15682,N_14921,N_15163);
xnor U15683 (N_15683,N_15028,N_15449);
nand U15684 (N_15684,N_14865,N_15247);
and U15685 (N_15685,N_14783,N_14941);
nor U15686 (N_15686,N_14429,N_14666);
and U15687 (N_15687,N_14704,N_15166);
nor U15688 (N_15688,N_14492,N_14900);
and U15689 (N_15689,N_15200,N_15133);
xor U15690 (N_15690,N_15090,N_14689);
or U15691 (N_15691,N_14482,N_14956);
nor U15692 (N_15692,N_14574,N_14795);
nand U15693 (N_15693,N_15299,N_14603);
nor U15694 (N_15694,N_14573,N_14440);
and U15695 (N_15695,N_14930,N_14587);
or U15696 (N_15696,N_14767,N_14968);
or U15697 (N_15697,N_15531,N_14692);
nand U15698 (N_15698,N_15057,N_14983);
and U15699 (N_15699,N_14551,N_15017);
xnor U15700 (N_15700,N_14986,N_14928);
nor U15701 (N_15701,N_14885,N_14873);
and U15702 (N_15702,N_14462,N_15491);
nand U15703 (N_15703,N_14621,N_15172);
or U15704 (N_15704,N_14805,N_15358);
xnor U15705 (N_15705,N_14717,N_14607);
nor U15706 (N_15706,N_14914,N_15507);
xnor U15707 (N_15707,N_14512,N_14601);
nand U15708 (N_15708,N_15384,N_15070);
and U15709 (N_15709,N_15575,N_14505);
xnor U15710 (N_15710,N_15315,N_14929);
xnor U15711 (N_15711,N_14957,N_14437);
and U15712 (N_15712,N_14516,N_15191);
and U15713 (N_15713,N_14459,N_15421);
or U15714 (N_15714,N_15175,N_14556);
and U15715 (N_15715,N_14665,N_15011);
xnor U15716 (N_15716,N_15071,N_14538);
nor U15717 (N_15717,N_14639,N_14544);
xor U15718 (N_15718,N_15132,N_14488);
nor U15719 (N_15719,N_15374,N_15514);
or U15720 (N_15720,N_14845,N_15186);
and U15721 (N_15721,N_14889,N_14520);
or U15722 (N_15722,N_15533,N_15340);
nand U15723 (N_15723,N_14720,N_15220);
xor U15724 (N_15724,N_14786,N_15463);
xor U15725 (N_15725,N_14477,N_14470);
and U15726 (N_15726,N_14909,N_14790);
nor U15727 (N_15727,N_14687,N_14696);
nor U15728 (N_15728,N_14655,N_15151);
xnor U15729 (N_15729,N_14846,N_15493);
and U15730 (N_15730,N_15121,N_15519);
and U15731 (N_15731,N_14454,N_15422);
and U15732 (N_15732,N_15430,N_14891);
xnor U15733 (N_15733,N_14995,N_15504);
and U15734 (N_15734,N_14887,N_15185);
and U15735 (N_15735,N_15149,N_14588);
xnor U15736 (N_15736,N_14948,N_14452);
or U15737 (N_15737,N_14691,N_15307);
nor U15738 (N_15738,N_14751,N_15513);
nand U15739 (N_15739,N_15031,N_14453);
and U15740 (N_15740,N_14646,N_14425);
or U15741 (N_15741,N_15221,N_15117);
nand U15742 (N_15742,N_14548,N_15215);
xor U15743 (N_15743,N_15357,N_15399);
and U15744 (N_15744,N_15119,N_15441);
xnor U15745 (N_15745,N_15045,N_15105);
xnor U15746 (N_15746,N_14649,N_14860);
nor U15747 (N_15747,N_14807,N_14936);
nor U15748 (N_15748,N_15564,N_15257);
nor U15749 (N_15749,N_14656,N_15096);
or U15750 (N_15750,N_15336,N_15012);
nor U15751 (N_15751,N_15294,N_14744);
nand U15752 (N_15752,N_15189,N_15183);
xnor U15753 (N_15753,N_14693,N_15505);
and U15754 (N_15754,N_15272,N_14823);
nor U15755 (N_15755,N_14545,N_14962);
or U15756 (N_15756,N_15196,N_15224);
nand U15757 (N_15757,N_14967,N_15197);
or U15758 (N_15758,N_14868,N_14448);
nand U15759 (N_15759,N_15243,N_14408);
nor U15760 (N_15760,N_15479,N_14716);
nor U15761 (N_15761,N_14654,N_15142);
nor U15762 (N_15762,N_14555,N_14474);
nand U15763 (N_15763,N_15334,N_15271);
and U15764 (N_15764,N_14970,N_14778);
or U15765 (N_15765,N_14486,N_15387);
xnor U15766 (N_15766,N_15008,N_14854);
nand U15767 (N_15767,N_15006,N_15318);
xor U15768 (N_15768,N_15035,N_15212);
nor U15769 (N_15769,N_15127,N_14937);
nor U15770 (N_15770,N_14966,N_14830);
xor U15771 (N_15771,N_14793,N_14570);
or U15772 (N_15772,N_15100,N_15506);
and U15773 (N_15773,N_15112,N_15195);
xnor U15774 (N_15774,N_14820,N_15495);
nand U15775 (N_15775,N_14682,N_15263);
and U15776 (N_15776,N_15459,N_14670);
xnor U15777 (N_15777,N_14964,N_15522);
xor U15778 (N_15778,N_15414,N_14910);
xnor U15779 (N_15779,N_15168,N_14418);
nor U15780 (N_15780,N_15555,N_14721);
nand U15781 (N_15781,N_15353,N_14747);
and U15782 (N_15782,N_15297,N_14765);
or U15783 (N_15783,N_14815,N_14536);
nand U15784 (N_15784,N_14722,N_14695);
and U15785 (N_15785,N_14822,N_14674);
nand U15786 (N_15786,N_15393,N_14750);
nor U15787 (N_15787,N_14762,N_14712);
nand U15788 (N_15788,N_15579,N_14614);
nor U15789 (N_15789,N_15388,N_14883);
nor U15790 (N_15790,N_14669,N_15301);
xnor U15791 (N_15791,N_14897,N_14532);
nor U15792 (N_15792,N_15217,N_15187);
xor U15793 (N_15793,N_15344,N_15007);
nand U15794 (N_15794,N_15558,N_15085);
xnor U15795 (N_15795,N_14547,N_14874);
and U15796 (N_15796,N_15559,N_14895);
or U15797 (N_15797,N_15295,N_15597);
or U15798 (N_15798,N_15198,N_14668);
and U15799 (N_15799,N_14612,N_15125);
nor U15800 (N_15800,N_14445,N_15370);
nand U15801 (N_15801,N_15206,N_15174);
xor U15802 (N_15802,N_14461,N_14675);
xnor U15803 (N_15803,N_15298,N_15079);
xor U15804 (N_15804,N_14839,N_15201);
xnor U15805 (N_15805,N_14705,N_15526);
nor U15806 (N_15806,N_14525,N_14902);
nor U15807 (N_15807,N_15044,N_15022);
xnor U15808 (N_15808,N_15192,N_14939);
nor U15809 (N_15809,N_14787,N_15069);
nand U15810 (N_15810,N_15068,N_15029);
and U15811 (N_15811,N_15102,N_15419);
and U15812 (N_15812,N_14504,N_15395);
and U15813 (N_15813,N_14749,N_15099);
xor U15814 (N_15814,N_14605,N_14800);
nand U15815 (N_15815,N_15123,N_15179);
and U15816 (N_15816,N_14502,N_15309);
nand U15817 (N_15817,N_15162,N_15319);
or U15818 (N_15818,N_15004,N_15154);
and U15819 (N_15819,N_15147,N_14527);
or U15820 (N_15820,N_14991,N_14679);
or U15821 (N_15821,N_15002,N_14879);
and U15822 (N_15822,N_15454,N_15234);
nor U15823 (N_15823,N_14485,N_15219);
xor U15824 (N_15824,N_14855,N_14513);
nor U15825 (N_15825,N_14899,N_15107);
nor U15826 (N_15826,N_14518,N_15415);
nand U15827 (N_15827,N_14926,N_15485);
nor U15828 (N_15828,N_14472,N_14444);
nor U15829 (N_15829,N_14908,N_14503);
nor U15830 (N_15830,N_15155,N_15581);
and U15831 (N_15831,N_14549,N_15335);
xnor U15832 (N_15832,N_15266,N_14741);
xnor U15833 (N_15833,N_14817,N_15489);
nor U15834 (N_15834,N_14495,N_15074);
xnor U15835 (N_15835,N_15134,N_15273);
nand U15836 (N_15836,N_14610,N_15472);
and U15837 (N_15837,N_14756,N_15039);
nor U15838 (N_15838,N_14867,N_14542);
nand U15839 (N_15839,N_15508,N_15239);
and U15840 (N_15840,N_15253,N_14616);
and U15841 (N_15841,N_15104,N_14647);
nor U15842 (N_15842,N_14530,N_14568);
xnor U15843 (N_15843,N_14489,N_14876);
nor U15844 (N_15844,N_14535,N_14519);
and U15845 (N_15845,N_15329,N_14739);
nor U15846 (N_15846,N_15033,N_15178);
and U15847 (N_15847,N_14458,N_15396);
and U15848 (N_15848,N_14412,N_14797);
nor U15849 (N_15849,N_14821,N_14803);
nor U15850 (N_15850,N_14738,N_15118);
and U15851 (N_15851,N_15106,N_15553);
nor U15852 (N_15852,N_15549,N_14529);
nand U15853 (N_15853,N_15473,N_14507);
or U15854 (N_15854,N_14652,N_15036);
nor U15855 (N_15855,N_15476,N_14890);
xor U15856 (N_15856,N_15408,N_15282);
or U15857 (N_15857,N_14441,N_15500);
nand U15858 (N_15858,N_14680,N_14735);
and U15859 (N_15859,N_15317,N_15116);
xor U15860 (N_15860,N_15445,N_14554);
nand U15861 (N_15861,N_14984,N_15356);
nand U15862 (N_15862,N_14996,N_15049);
xnor U15863 (N_15863,N_14950,N_15528);
xor U15864 (N_15864,N_14491,N_15177);
xor U15865 (N_15865,N_14758,N_15331);
nor U15866 (N_15866,N_14761,N_15416);
or U15867 (N_15867,N_15173,N_15432);
nand U15868 (N_15868,N_15497,N_15233);
and U15869 (N_15869,N_15268,N_15350);
nand U15870 (N_15870,N_14918,N_15450);
nand U15871 (N_15871,N_15438,N_14677);
xnor U15872 (N_15872,N_14882,N_15015);
and U15873 (N_15873,N_15523,N_14400);
or U15874 (N_15874,N_14479,N_15561);
nand U15875 (N_15875,N_15509,N_14596);
and U15876 (N_15876,N_14952,N_14760);
or U15877 (N_15877,N_14771,N_14620);
nand U15878 (N_15878,N_14825,N_14944);
xor U15879 (N_15879,N_14659,N_14602);
nor U15880 (N_15880,N_14958,N_14922);
or U15881 (N_15881,N_14469,N_15580);
and U15882 (N_15882,N_15452,N_15274);
xnor U15883 (N_15883,N_14755,N_15584);
nand U15884 (N_15884,N_15202,N_14784);
nor U15885 (N_15885,N_14780,N_15498);
xor U15886 (N_15886,N_15516,N_15541);
nor U15887 (N_15887,N_15499,N_14508);
or U15888 (N_15888,N_15349,N_14493);
and U15889 (N_15889,N_15086,N_14924);
or U15890 (N_15890,N_15312,N_15587);
and U15891 (N_15891,N_14476,N_14553);
and U15892 (N_15892,N_15019,N_15378);
and U15893 (N_15893,N_14660,N_15053);
and U15894 (N_15894,N_14730,N_15148);
nand U15895 (N_15895,N_15180,N_14420);
xnor U15896 (N_15896,N_15440,N_15546);
and U15897 (N_15897,N_15095,N_15169);
xor U15898 (N_15898,N_14714,N_15397);
nand U15899 (N_15899,N_15120,N_15381);
and U15900 (N_15900,N_14840,N_15333);
nor U15901 (N_15901,N_15027,N_15518);
or U15902 (N_15902,N_14759,N_14559);
and U15903 (N_15903,N_15595,N_14584);
nand U15904 (N_15904,N_15126,N_14615);
or U15905 (N_15905,N_14774,N_14487);
and U15906 (N_15906,N_15321,N_14731);
and U15907 (N_15907,N_15355,N_14606);
and U15908 (N_15908,N_14935,N_14627);
nand U15909 (N_15909,N_15451,N_15275);
or U15910 (N_15910,N_14764,N_15109);
or U15911 (N_15911,N_15391,N_15455);
nand U15912 (N_15912,N_15306,N_15572);
and U15913 (N_15913,N_15588,N_15135);
nand U15914 (N_15914,N_15223,N_15139);
nor U15915 (N_15915,N_15556,N_14599);
or U15916 (N_15916,N_15591,N_15529);
nor U15917 (N_15917,N_14775,N_14501);
and U15918 (N_15918,N_14979,N_15480);
nor U15919 (N_15919,N_14510,N_15083);
nand U15920 (N_15920,N_15348,N_15230);
xnor U15921 (N_15921,N_14480,N_14903);
or U15922 (N_15922,N_14772,N_14917);
or U15923 (N_15923,N_15260,N_15313);
nand U15924 (N_15924,N_15448,N_14683);
and U15925 (N_15925,N_14702,N_15524);
or U15926 (N_15926,N_14838,N_14844);
and U15927 (N_15927,N_14988,N_15574);
or U15928 (N_15928,N_15337,N_14806);
xor U15929 (N_15929,N_14710,N_14861);
nand U15930 (N_15930,N_15372,N_14638);
nand U15931 (N_15931,N_15401,N_14597);
nor U15932 (N_15932,N_14585,N_14965);
nand U15933 (N_15933,N_14951,N_15474);
and U15934 (N_15934,N_15300,N_14631);
nand U15935 (N_15935,N_15005,N_15383);
nor U15936 (N_15936,N_15088,N_15471);
or U15937 (N_15937,N_15503,N_15339);
nor U15938 (N_15938,N_14433,N_15483);
nand U15939 (N_15939,N_14658,N_14431);
and U15940 (N_15940,N_15554,N_15457);
and U15941 (N_15941,N_15411,N_15256);
xnor U15942 (N_15942,N_14972,N_15486);
xnor U15943 (N_15943,N_14801,N_14463);
and U15944 (N_15944,N_15021,N_15332);
xnor U15945 (N_15945,N_15303,N_14911);
nand U15946 (N_15946,N_14782,N_15308);
nor U15947 (N_15947,N_14651,N_14872);
and U15948 (N_15948,N_14526,N_14411);
xnor U15949 (N_15949,N_15547,N_14577);
nand U15950 (N_15950,N_14466,N_15160);
nand U15951 (N_15951,N_15066,N_14792);
or U15952 (N_15952,N_15293,N_15314);
or U15953 (N_15953,N_15400,N_15001);
and U15954 (N_15954,N_15578,N_14633);
xor U15955 (N_15955,N_15327,N_14572);
and U15956 (N_15956,N_15248,N_15567);
or U15957 (N_15957,N_15170,N_14954);
or U15958 (N_15958,N_14907,N_15369);
nand U15959 (N_15959,N_14881,N_15427);
or U15960 (N_15960,N_15181,N_14877);
and U15961 (N_15961,N_15324,N_14985);
xor U15962 (N_15962,N_14718,N_15594);
nand U15963 (N_15963,N_15061,N_15062);
nor U15964 (N_15964,N_14608,N_14947);
xor U15965 (N_15965,N_14955,N_14401);
and U15966 (N_15966,N_15537,N_15236);
nor U15967 (N_15967,N_15592,N_14736);
xnor U15968 (N_15968,N_14637,N_15392);
xnor U15969 (N_15969,N_14500,N_15003);
nor U15970 (N_15970,N_14423,N_15359);
or U15971 (N_15971,N_14849,N_14733);
xor U15972 (N_15972,N_14713,N_14706);
xor U15973 (N_15973,N_15246,N_14403);
or U15974 (N_15974,N_15081,N_15059);
or U15975 (N_15975,N_14419,N_15159);
nor U15976 (N_15976,N_14901,N_14794);
and U15977 (N_15977,N_14875,N_14852);
nand U15978 (N_15978,N_15176,N_14848);
nor U15979 (N_15979,N_14933,N_14523);
or U15980 (N_15980,N_14905,N_14886);
or U15981 (N_15981,N_14748,N_15585);
xor U15982 (N_15982,N_15515,N_15379);
and U15983 (N_15983,N_14737,N_14913);
nand U15984 (N_15984,N_14829,N_14723);
and U15985 (N_15985,N_15341,N_14975);
or U15986 (N_15986,N_15351,N_14407);
nand U15987 (N_15987,N_15240,N_15482);
xnor U15988 (N_15988,N_15161,N_15091);
nand U15989 (N_15989,N_14893,N_14769);
nor U15990 (N_15990,N_14814,N_14591);
and U15991 (N_15991,N_15361,N_15286);
xnor U15992 (N_15992,N_14862,N_15470);
xnor U15993 (N_15993,N_14634,N_15205);
and U15994 (N_15994,N_14578,N_15216);
nor U15995 (N_15995,N_14916,N_14455);
or U15996 (N_15996,N_14934,N_15389);
or U15997 (N_15997,N_14963,N_15484);
and U15998 (N_15998,N_14406,N_15490);
nor U15999 (N_15999,N_14582,N_14629);
and U16000 (N_16000,N_15153,N_15265);
or U16001 (N_16001,N_14630,N_15164);
xnor U16002 (N_16002,N_15214,N_15042);
and U16003 (N_16003,N_15141,N_15250);
nand U16004 (N_16004,N_15140,N_14711);
or U16005 (N_16005,N_14992,N_14728);
xnor U16006 (N_16006,N_14745,N_14497);
xnor U16007 (N_16007,N_14919,N_14866);
or U16008 (N_16008,N_15596,N_14590);
and U16009 (N_16009,N_14511,N_14942);
and U16010 (N_16010,N_15466,N_14715);
nand U16011 (N_16011,N_15311,N_14566);
nor U16012 (N_16012,N_15122,N_14571);
xor U16013 (N_16013,N_14528,N_14404);
nor U16014 (N_16014,N_15194,N_15590);
nor U16015 (N_16015,N_15538,N_15150);
xor U16016 (N_16016,N_14467,N_14673);
nand U16017 (N_16017,N_15014,N_15412);
and U16018 (N_16018,N_14833,N_14904);
nand U16019 (N_16019,N_14943,N_14898);
nor U16020 (N_16020,N_15550,N_15433);
nor U16021 (N_16021,N_15165,N_15468);
xnor U16022 (N_16022,N_15539,N_15075);
and U16023 (N_16023,N_14773,N_14442);
nor U16024 (N_16024,N_14923,N_15037);
or U16025 (N_16025,N_14785,N_15078);
nor U16026 (N_16026,N_15458,N_15292);
nand U16027 (N_16027,N_15310,N_15157);
xnor U16028 (N_16028,N_14457,N_14998);
or U16029 (N_16029,N_15056,N_15434);
xor U16030 (N_16030,N_14927,N_15034);
nand U16031 (N_16031,N_14997,N_15290);
nand U16032 (N_16032,N_14636,N_15326);
nand U16033 (N_16033,N_15425,N_14600);
and U16034 (N_16034,N_15211,N_15403);
and U16035 (N_16035,N_14449,N_15382);
and U16036 (N_16036,N_15067,N_14481);
xor U16037 (N_16037,N_14434,N_15409);
or U16038 (N_16038,N_14506,N_15338);
and U16039 (N_16039,N_14809,N_14413);
nand U16040 (N_16040,N_14931,N_14617);
nor U16041 (N_16041,N_14611,N_14732);
nor U16042 (N_16042,N_15111,N_15281);
nor U16043 (N_16043,N_14953,N_15000);
xor U16044 (N_16044,N_14626,N_14896);
or U16045 (N_16045,N_15530,N_15568);
and U16046 (N_16046,N_14609,N_15089);
nand U16047 (N_16047,N_14575,N_14490);
nor U16048 (N_16048,N_15209,N_14850);
and U16049 (N_16049,N_15548,N_14625);
xnor U16050 (N_16050,N_14856,N_14859);
or U16051 (N_16051,N_15080,N_15521);
and U16052 (N_16052,N_14810,N_15413);
xnor U16053 (N_16053,N_15101,N_14644);
or U16054 (N_16054,N_14541,N_15502);
and U16055 (N_16055,N_14586,N_15525);
or U16056 (N_16056,N_15577,N_15188);
and U16057 (N_16057,N_15444,N_14700);
nor U16058 (N_16058,N_15261,N_15496);
and U16059 (N_16059,N_14811,N_14642);
and U16060 (N_16060,N_14828,N_15048);
and U16061 (N_16061,N_14478,N_14804);
nand U16062 (N_16062,N_15589,N_15436);
xnor U16063 (N_16063,N_14436,N_14417);
nand U16064 (N_16064,N_15532,N_15543);
xnor U16065 (N_16065,N_14465,N_15032);
or U16066 (N_16066,N_15026,N_14938);
nand U16067 (N_16067,N_15465,N_14635);
xor U16068 (N_16068,N_14426,N_14560);
nor U16069 (N_16069,N_15182,N_15225);
or U16070 (N_16070,N_15510,N_15145);
xnor U16071 (N_16071,N_14753,N_14779);
nor U16072 (N_16072,N_14853,N_14808);
xor U16073 (N_16073,N_15084,N_15144);
nand U16074 (N_16074,N_15058,N_15501);
and U16075 (N_16075,N_15456,N_14593);
nor U16076 (N_16076,N_14915,N_14880);
xor U16077 (N_16077,N_14832,N_15447);
xnor U16078 (N_16078,N_15167,N_15405);
nor U16079 (N_16079,N_15593,N_15137);
xor U16080 (N_16080,N_14496,N_14409);
nand U16081 (N_16081,N_14837,N_15492);
nor U16082 (N_16082,N_14543,N_15285);
and U16083 (N_16083,N_14842,N_15365);
xor U16084 (N_16084,N_14422,N_14707);
or U16085 (N_16085,N_14977,N_14402);
nand U16086 (N_16086,N_14757,N_14550);
nor U16087 (N_16087,N_15536,N_14766);
and U16088 (N_16088,N_14763,N_14561);
nor U16089 (N_16089,N_15423,N_15025);
and U16090 (N_16090,N_14468,N_14604);
or U16091 (N_16091,N_15363,N_15583);
xnor U16092 (N_16092,N_15560,N_15203);
or U16093 (N_16093,N_14940,N_15362);
xor U16094 (N_16094,N_14613,N_15442);
nor U16095 (N_16095,N_14581,N_15077);
or U16096 (N_16096,N_14726,N_14688);
nand U16097 (N_16097,N_15051,N_14777);
or U16098 (N_16098,N_14522,N_14894);
and U16099 (N_16099,N_15542,N_14514);
xor U16100 (N_16100,N_14415,N_14565);
or U16101 (N_16101,N_15385,N_14499);
or U16102 (N_16102,N_14802,N_15146);
nand U16103 (N_16103,N_15130,N_15477);
nor U16104 (N_16104,N_14827,N_14836);
nand U16105 (N_16105,N_14945,N_15092);
nand U16106 (N_16106,N_15535,N_15207);
or U16107 (N_16107,N_15511,N_14796);
xor U16108 (N_16108,N_14498,N_15269);
nand U16109 (N_16109,N_15143,N_15129);
nor U16110 (N_16110,N_14421,N_15461);
nand U16111 (N_16111,N_14521,N_15367);
and U16112 (N_16112,N_14558,N_15342);
or U16113 (N_16113,N_15020,N_15043);
or U16114 (N_16114,N_15055,N_15047);
or U16115 (N_16115,N_15552,N_14851);
xor U16116 (N_16116,N_14446,N_14438);
xor U16117 (N_16117,N_15322,N_15060);
nor U16118 (N_16118,N_15376,N_15241);
xor U16119 (N_16119,N_15259,N_15418);
xnor U16120 (N_16120,N_15453,N_15046);
xnor U16121 (N_16121,N_15557,N_14871);
and U16122 (N_16122,N_14456,N_15010);
nor U16123 (N_16123,N_15231,N_15193);
nor U16124 (N_16124,N_14788,N_14664);
or U16125 (N_16125,N_15276,N_15267);
nor U16126 (N_16126,N_14546,N_14819);
nand U16127 (N_16127,N_15072,N_14690);
nor U16128 (N_16128,N_14662,N_14694);
nand U16129 (N_16129,N_14464,N_15323);
nand U16130 (N_16130,N_14671,N_15023);
nand U16131 (N_16131,N_14980,N_14557);
or U16132 (N_16132,N_15464,N_15156);
nor U16133 (N_16133,N_14460,N_14708);
xor U16134 (N_16134,N_14813,N_14699);
xnor U16135 (N_16135,N_14912,N_14746);
nand U16136 (N_16136,N_14971,N_15566);
and U16137 (N_16137,N_14443,N_14447);
and U16138 (N_16138,N_14685,N_14906);
and U16139 (N_16139,N_14676,N_15487);
nor U16140 (N_16140,N_15283,N_14428);
or U16141 (N_16141,N_15016,N_15364);
and U16142 (N_16142,N_15213,N_14537);
nand U16143 (N_16143,N_14946,N_15571);
xnor U16144 (N_16144,N_15093,N_14540);
or U16145 (N_16145,N_15258,N_14405);
nand U16146 (N_16146,N_15210,N_15254);
nor U16147 (N_16147,N_15375,N_14864);
or U16148 (N_16148,N_14994,N_15582);
nor U16149 (N_16149,N_15063,N_15018);
and U16150 (N_16150,N_15527,N_15420);
nand U16151 (N_16151,N_15255,N_14989);
nand U16152 (N_16152,N_14925,N_15347);
or U16153 (N_16153,N_14598,N_14524);
nand U16154 (N_16154,N_15094,N_14734);
xnor U16155 (N_16155,N_14959,N_15417);
xor U16156 (N_16156,N_15328,N_14592);
nor U16157 (N_16157,N_14843,N_15371);
xnor U16158 (N_16158,N_14643,N_15288);
xnor U16159 (N_16159,N_14533,N_15563);
and U16160 (N_16160,N_14993,N_15431);
and U16161 (N_16161,N_15551,N_14932);
and U16162 (N_16162,N_14475,N_14969);
and U16163 (N_16163,N_14949,N_15534);
nor U16164 (N_16164,N_14678,N_15050);
xnor U16165 (N_16165,N_15446,N_15222);
or U16166 (N_16166,N_15598,N_15098);
nand U16167 (N_16167,N_14835,N_15073);
nand U16168 (N_16168,N_14847,N_14831);
nor U16169 (N_16169,N_15289,N_14770);
nor U16170 (N_16170,N_14632,N_15377);
nor U16171 (N_16171,N_15097,N_15238);
and U16172 (N_16172,N_15424,N_14569);
xnor U16173 (N_16173,N_15494,N_15158);
xor U16174 (N_16174,N_15565,N_14703);
and U16175 (N_16175,N_14701,N_14789);
xnor U16176 (N_16176,N_15366,N_14564);
nand U16177 (N_16177,N_15296,N_14857);
xor U16178 (N_16178,N_14719,N_14684);
or U16179 (N_16179,N_14743,N_14697);
nor U16180 (N_16180,N_15138,N_14698);
xnor U16181 (N_16181,N_15199,N_15469);
nand U16182 (N_16182,N_15343,N_14781);
nor U16183 (N_16183,N_15540,N_14870);
nor U16184 (N_16184,N_15517,N_15316);
and U16185 (N_16185,N_14539,N_14884);
or U16186 (N_16186,N_15386,N_14768);
nor U16187 (N_16187,N_14999,N_15208);
nand U16188 (N_16188,N_15599,N_15390);
xor U16189 (N_16189,N_14414,N_14858);
and U16190 (N_16190,N_15404,N_14740);
xor U16191 (N_16191,N_15426,N_15245);
nand U16192 (N_16192,N_15184,N_14624);
or U16193 (N_16193,N_15052,N_14816);
and U16194 (N_16194,N_14416,N_14622);
xnor U16195 (N_16195,N_15443,N_15398);
xnor U16196 (N_16196,N_15354,N_15114);
nor U16197 (N_16197,N_15394,N_14650);
xnor U16198 (N_16198,N_14826,N_14473);
and U16199 (N_16199,N_14534,N_15218);
and U16200 (N_16200,N_14966,N_15049);
nand U16201 (N_16201,N_14814,N_15574);
xor U16202 (N_16202,N_15553,N_14436);
and U16203 (N_16203,N_14927,N_14541);
or U16204 (N_16204,N_15050,N_14783);
or U16205 (N_16205,N_14928,N_14961);
nand U16206 (N_16206,N_14987,N_15237);
nand U16207 (N_16207,N_15563,N_15137);
or U16208 (N_16208,N_14900,N_15054);
nand U16209 (N_16209,N_15020,N_14929);
xor U16210 (N_16210,N_14457,N_14493);
nor U16211 (N_16211,N_15173,N_14896);
or U16212 (N_16212,N_14954,N_14604);
and U16213 (N_16213,N_15309,N_15038);
nor U16214 (N_16214,N_15127,N_14829);
and U16215 (N_16215,N_14793,N_15527);
nand U16216 (N_16216,N_14962,N_15210);
nand U16217 (N_16217,N_14676,N_14712);
and U16218 (N_16218,N_15150,N_15446);
nand U16219 (N_16219,N_14998,N_14476);
nand U16220 (N_16220,N_15059,N_15307);
and U16221 (N_16221,N_14936,N_15528);
and U16222 (N_16222,N_15121,N_14713);
or U16223 (N_16223,N_15266,N_15376);
and U16224 (N_16224,N_14958,N_14576);
xor U16225 (N_16225,N_14665,N_14838);
nand U16226 (N_16226,N_15449,N_14657);
nor U16227 (N_16227,N_14479,N_15540);
nor U16228 (N_16228,N_15588,N_14634);
or U16229 (N_16229,N_15132,N_14997);
nor U16230 (N_16230,N_14674,N_14719);
nand U16231 (N_16231,N_14961,N_15387);
xor U16232 (N_16232,N_15428,N_14618);
xor U16233 (N_16233,N_14929,N_15223);
or U16234 (N_16234,N_14688,N_14471);
or U16235 (N_16235,N_14772,N_15425);
or U16236 (N_16236,N_15192,N_14698);
nor U16237 (N_16237,N_14842,N_15259);
xor U16238 (N_16238,N_15463,N_15200);
nor U16239 (N_16239,N_15020,N_15597);
nand U16240 (N_16240,N_15232,N_14576);
xnor U16241 (N_16241,N_15414,N_15537);
nor U16242 (N_16242,N_15592,N_14988);
nand U16243 (N_16243,N_14413,N_14541);
or U16244 (N_16244,N_14847,N_15002);
xnor U16245 (N_16245,N_15215,N_15537);
or U16246 (N_16246,N_15374,N_14800);
nor U16247 (N_16247,N_15528,N_15411);
xnor U16248 (N_16248,N_14883,N_14705);
and U16249 (N_16249,N_15179,N_14982);
and U16250 (N_16250,N_14787,N_14812);
xor U16251 (N_16251,N_14877,N_15013);
or U16252 (N_16252,N_15497,N_14499);
nor U16253 (N_16253,N_15503,N_14609);
or U16254 (N_16254,N_15576,N_14776);
and U16255 (N_16255,N_15309,N_14519);
xor U16256 (N_16256,N_15056,N_15278);
and U16257 (N_16257,N_15304,N_14751);
or U16258 (N_16258,N_14728,N_15549);
xor U16259 (N_16259,N_14586,N_14990);
nand U16260 (N_16260,N_15048,N_15357);
or U16261 (N_16261,N_15160,N_14543);
xnor U16262 (N_16262,N_14924,N_15436);
and U16263 (N_16263,N_14443,N_15290);
nor U16264 (N_16264,N_14676,N_14952);
xnor U16265 (N_16265,N_14835,N_14564);
and U16266 (N_16266,N_15270,N_15213);
nand U16267 (N_16267,N_15153,N_15022);
xnor U16268 (N_16268,N_15559,N_14817);
xnor U16269 (N_16269,N_14401,N_15554);
xnor U16270 (N_16270,N_15466,N_14679);
nand U16271 (N_16271,N_15454,N_14623);
or U16272 (N_16272,N_14908,N_14769);
nand U16273 (N_16273,N_15045,N_15314);
xnor U16274 (N_16274,N_15158,N_15030);
nor U16275 (N_16275,N_15334,N_15189);
and U16276 (N_16276,N_14934,N_14598);
nor U16277 (N_16277,N_14628,N_15576);
nand U16278 (N_16278,N_14562,N_14648);
and U16279 (N_16279,N_15057,N_15391);
xnor U16280 (N_16280,N_15219,N_14723);
and U16281 (N_16281,N_15167,N_14840);
nand U16282 (N_16282,N_14594,N_14905);
nor U16283 (N_16283,N_14959,N_15592);
and U16284 (N_16284,N_15179,N_15175);
or U16285 (N_16285,N_15370,N_14844);
or U16286 (N_16286,N_14549,N_14987);
nor U16287 (N_16287,N_14910,N_15079);
and U16288 (N_16288,N_15174,N_14436);
xor U16289 (N_16289,N_14495,N_15162);
and U16290 (N_16290,N_14763,N_14748);
xor U16291 (N_16291,N_14868,N_14440);
and U16292 (N_16292,N_14574,N_14923);
or U16293 (N_16293,N_15490,N_15543);
nand U16294 (N_16294,N_14982,N_15546);
nand U16295 (N_16295,N_15536,N_15472);
nor U16296 (N_16296,N_14818,N_14965);
or U16297 (N_16297,N_14751,N_14599);
xor U16298 (N_16298,N_15285,N_14498);
nor U16299 (N_16299,N_15200,N_15268);
or U16300 (N_16300,N_15289,N_14956);
nor U16301 (N_16301,N_14463,N_15247);
nand U16302 (N_16302,N_14400,N_14869);
nand U16303 (N_16303,N_15526,N_14814);
or U16304 (N_16304,N_15331,N_14854);
and U16305 (N_16305,N_15416,N_15129);
nor U16306 (N_16306,N_14754,N_14788);
xor U16307 (N_16307,N_14712,N_15551);
nor U16308 (N_16308,N_15132,N_15333);
and U16309 (N_16309,N_14415,N_14474);
xnor U16310 (N_16310,N_14883,N_14562);
nand U16311 (N_16311,N_15546,N_14600);
and U16312 (N_16312,N_15326,N_15208);
and U16313 (N_16313,N_14937,N_14636);
nand U16314 (N_16314,N_15249,N_14946);
xor U16315 (N_16315,N_14455,N_14807);
and U16316 (N_16316,N_14675,N_14746);
nor U16317 (N_16317,N_14929,N_14894);
or U16318 (N_16318,N_14824,N_15012);
nor U16319 (N_16319,N_15485,N_15070);
xnor U16320 (N_16320,N_15479,N_14416);
xor U16321 (N_16321,N_14873,N_14950);
xor U16322 (N_16322,N_15501,N_15162);
or U16323 (N_16323,N_15160,N_15470);
and U16324 (N_16324,N_15028,N_14597);
nor U16325 (N_16325,N_15479,N_14432);
nand U16326 (N_16326,N_14662,N_15210);
and U16327 (N_16327,N_15186,N_15322);
and U16328 (N_16328,N_15229,N_14400);
and U16329 (N_16329,N_15001,N_15029);
nor U16330 (N_16330,N_15179,N_15183);
nor U16331 (N_16331,N_15279,N_14424);
xnor U16332 (N_16332,N_15367,N_15321);
xnor U16333 (N_16333,N_14405,N_14903);
nor U16334 (N_16334,N_15402,N_14963);
nand U16335 (N_16335,N_14710,N_15056);
xnor U16336 (N_16336,N_15237,N_15057);
nand U16337 (N_16337,N_14459,N_14452);
xor U16338 (N_16338,N_15028,N_14420);
nor U16339 (N_16339,N_14593,N_15235);
or U16340 (N_16340,N_14649,N_15110);
or U16341 (N_16341,N_14471,N_14847);
or U16342 (N_16342,N_14756,N_14609);
and U16343 (N_16343,N_14457,N_15088);
xnor U16344 (N_16344,N_15114,N_15440);
or U16345 (N_16345,N_15054,N_15567);
nand U16346 (N_16346,N_15158,N_14429);
nand U16347 (N_16347,N_15286,N_15067);
nor U16348 (N_16348,N_14607,N_14652);
xor U16349 (N_16349,N_14955,N_15006);
and U16350 (N_16350,N_15191,N_15385);
and U16351 (N_16351,N_14696,N_15473);
xor U16352 (N_16352,N_14457,N_14769);
and U16353 (N_16353,N_14769,N_15063);
or U16354 (N_16354,N_15272,N_14527);
nand U16355 (N_16355,N_15487,N_14745);
or U16356 (N_16356,N_15418,N_15461);
nor U16357 (N_16357,N_14490,N_14802);
xnor U16358 (N_16358,N_15432,N_14748);
xor U16359 (N_16359,N_14432,N_14816);
nor U16360 (N_16360,N_15354,N_14809);
and U16361 (N_16361,N_15141,N_15273);
nand U16362 (N_16362,N_15110,N_14803);
nor U16363 (N_16363,N_14738,N_14726);
nor U16364 (N_16364,N_15474,N_14838);
nand U16365 (N_16365,N_14410,N_15115);
nand U16366 (N_16366,N_15502,N_14699);
or U16367 (N_16367,N_14444,N_14881);
and U16368 (N_16368,N_14567,N_15146);
and U16369 (N_16369,N_15231,N_14948);
nand U16370 (N_16370,N_14869,N_15219);
or U16371 (N_16371,N_14850,N_14620);
nor U16372 (N_16372,N_15118,N_15338);
and U16373 (N_16373,N_15337,N_15019);
and U16374 (N_16374,N_15205,N_14532);
or U16375 (N_16375,N_14943,N_15565);
and U16376 (N_16376,N_15504,N_14528);
and U16377 (N_16377,N_15473,N_15575);
and U16378 (N_16378,N_14571,N_15111);
and U16379 (N_16379,N_14655,N_15595);
or U16380 (N_16380,N_14451,N_15212);
xor U16381 (N_16381,N_14870,N_15577);
nor U16382 (N_16382,N_15401,N_15014);
nand U16383 (N_16383,N_14719,N_14972);
or U16384 (N_16384,N_15268,N_15271);
xor U16385 (N_16385,N_14691,N_14626);
nand U16386 (N_16386,N_15052,N_15577);
or U16387 (N_16387,N_15126,N_15270);
nand U16388 (N_16388,N_14814,N_15148);
or U16389 (N_16389,N_15374,N_15432);
or U16390 (N_16390,N_14731,N_14478);
and U16391 (N_16391,N_15155,N_14544);
xor U16392 (N_16392,N_15480,N_14544);
and U16393 (N_16393,N_14966,N_15194);
and U16394 (N_16394,N_15276,N_15574);
and U16395 (N_16395,N_15033,N_14987);
and U16396 (N_16396,N_14770,N_15424);
or U16397 (N_16397,N_14429,N_15091);
xor U16398 (N_16398,N_15252,N_14686);
nand U16399 (N_16399,N_14983,N_15129);
and U16400 (N_16400,N_15171,N_15432);
or U16401 (N_16401,N_15128,N_15167);
nor U16402 (N_16402,N_14950,N_14863);
nor U16403 (N_16403,N_15102,N_15374);
nand U16404 (N_16404,N_14658,N_14801);
or U16405 (N_16405,N_15155,N_15280);
and U16406 (N_16406,N_14535,N_14839);
and U16407 (N_16407,N_15017,N_15432);
xnor U16408 (N_16408,N_15345,N_15179);
and U16409 (N_16409,N_14581,N_15562);
and U16410 (N_16410,N_14925,N_14855);
and U16411 (N_16411,N_15481,N_15402);
or U16412 (N_16412,N_14500,N_14482);
nand U16413 (N_16413,N_15071,N_14412);
and U16414 (N_16414,N_14696,N_14503);
and U16415 (N_16415,N_14569,N_15123);
nor U16416 (N_16416,N_14674,N_15270);
and U16417 (N_16417,N_14755,N_15233);
or U16418 (N_16418,N_14445,N_15132);
and U16419 (N_16419,N_14910,N_14899);
nor U16420 (N_16420,N_15135,N_14782);
and U16421 (N_16421,N_14789,N_14656);
and U16422 (N_16422,N_14999,N_14737);
and U16423 (N_16423,N_14413,N_14508);
and U16424 (N_16424,N_15291,N_15155);
xor U16425 (N_16425,N_14456,N_14629);
and U16426 (N_16426,N_15322,N_14526);
and U16427 (N_16427,N_14749,N_15534);
nand U16428 (N_16428,N_15138,N_15115);
and U16429 (N_16429,N_14652,N_14729);
nor U16430 (N_16430,N_15218,N_15277);
or U16431 (N_16431,N_15504,N_15278);
nor U16432 (N_16432,N_14444,N_15012);
nor U16433 (N_16433,N_14950,N_15425);
xnor U16434 (N_16434,N_14590,N_14849);
xnor U16435 (N_16435,N_14881,N_15189);
and U16436 (N_16436,N_15260,N_15375);
or U16437 (N_16437,N_14618,N_14937);
nor U16438 (N_16438,N_14421,N_15163);
nand U16439 (N_16439,N_14462,N_15123);
nor U16440 (N_16440,N_14466,N_14752);
or U16441 (N_16441,N_14781,N_14749);
nor U16442 (N_16442,N_15454,N_15151);
and U16443 (N_16443,N_14712,N_14690);
nor U16444 (N_16444,N_14570,N_15167);
nor U16445 (N_16445,N_15422,N_14887);
xor U16446 (N_16446,N_15425,N_15232);
nor U16447 (N_16447,N_15509,N_15477);
or U16448 (N_16448,N_14608,N_15348);
xnor U16449 (N_16449,N_15481,N_15522);
nand U16450 (N_16450,N_14452,N_15563);
nand U16451 (N_16451,N_14747,N_15278);
and U16452 (N_16452,N_14631,N_14890);
or U16453 (N_16453,N_14627,N_15088);
nor U16454 (N_16454,N_14452,N_15038);
nor U16455 (N_16455,N_15396,N_15335);
and U16456 (N_16456,N_15304,N_14560);
nor U16457 (N_16457,N_14432,N_15403);
xor U16458 (N_16458,N_15325,N_15342);
nor U16459 (N_16459,N_14589,N_15010);
nor U16460 (N_16460,N_15505,N_15576);
and U16461 (N_16461,N_14498,N_15395);
nor U16462 (N_16462,N_14557,N_15329);
nand U16463 (N_16463,N_15176,N_15346);
nand U16464 (N_16464,N_14794,N_15357);
xor U16465 (N_16465,N_15165,N_14520);
or U16466 (N_16466,N_14485,N_14694);
nor U16467 (N_16467,N_14846,N_14952);
and U16468 (N_16468,N_14464,N_15540);
nand U16469 (N_16469,N_14678,N_15060);
nand U16470 (N_16470,N_14822,N_15328);
and U16471 (N_16471,N_14921,N_15077);
nand U16472 (N_16472,N_14560,N_15535);
and U16473 (N_16473,N_15025,N_15211);
nand U16474 (N_16474,N_15545,N_14795);
or U16475 (N_16475,N_14825,N_15480);
or U16476 (N_16476,N_15341,N_14713);
xnor U16477 (N_16477,N_15510,N_14722);
nor U16478 (N_16478,N_15529,N_15038);
nor U16479 (N_16479,N_15017,N_15142);
and U16480 (N_16480,N_14791,N_15386);
xor U16481 (N_16481,N_15441,N_14786);
nor U16482 (N_16482,N_15355,N_14641);
xnor U16483 (N_16483,N_14869,N_14694);
nor U16484 (N_16484,N_15497,N_14947);
or U16485 (N_16485,N_15368,N_15576);
or U16486 (N_16486,N_14683,N_14888);
or U16487 (N_16487,N_14732,N_14847);
xor U16488 (N_16488,N_15448,N_14784);
xnor U16489 (N_16489,N_15326,N_15407);
nor U16490 (N_16490,N_14845,N_14764);
nor U16491 (N_16491,N_15154,N_15030);
nand U16492 (N_16492,N_15157,N_14904);
nand U16493 (N_16493,N_15222,N_15074);
xor U16494 (N_16494,N_14456,N_14820);
or U16495 (N_16495,N_15355,N_15042);
nor U16496 (N_16496,N_14481,N_15576);
nor U16497 (N_16497,N_14674,N_14404);
nand U16498 (N_16498,N_14906,N_15297);
and U16499 (N_16499,N_14614,N_15454);
and U16500 (N_16500,N_15403,N_14457);
and U16501 (N_16501,N_14926,N_14918);
and U16502 (N_16502,N_15349,N_14764);
xor U16503 (N_16503,N_15177,N_14469);
and U16504 (N_16504,N_15461,N_14731);
or U16505 (N_16505,N_15006,N_15160);
xor U16506 (N_16506,N_15118,N_14525);
and U16507 (N_16507,N_14976,N_15521);
and U16508 (N_16508,N_15163,N_14695);
xor U16509 (N_16509,N_14962,N_14571);
xor U16510 (N_16510,N_15108,N_14894);
and U16511 (N_16511,N_15409,N_15062);
and U16512 (N_16512,N_14799,N_15454);
nand U16513 (N_16513,N_15584,N_14768);
and U16514 (N_16514,N_14606,N_15592);
or U16515 (N_16515,N_15284,N_15261);
or U16516 (N_16516,N_15030,N_14725);
or U16517 (N_16517,N_15153,N_15114);
nand U16518 (N_16518,N_15345,N_14675);
xor U16519 (N_16519,N_14626,N_15363);
xnor U16520 (N_16520,N_14661,N_15129);
xnor U16521 (N_16521,N_14857,N_14634);
and U16522 (N_16522,N_15315,N_15373);
xnor U16523 (N_16523,N_14733,N_14823);
nand U16524 (N_16524,N_15082,N_14609);
nand U16525 (N_16525,N_15144,N_14453);
or U16526 (N_16526,N_14548,N_15269);
nor U16527 (N_16527,N_14830,N_14997);
xor U16528 (N_16528,N_14829,N_14915);
or U16529 (N_16529,N_14561,N_14627);
nand U16530 (N_16530,N_14823,N_15401);
xor U16531 (N_16531,N_15464,N_14889);
nand U16532 (N_16532,N_14871,N_15323);
xor U16533 (N_16533,N_15192,N_14622);
nor U16534 (N_16534,N_15277,N_15479);
xor U16535 (N_16535,N_14867,N_14585);
nand U16536 (N_16536,N_15280,N_14760);
or U16537 (N_16537,N_15472,N_15067);
or U16538 (N_16538,N_15069,N_14464);
and U16539 (N_16539,N_14874,N_14543);
nand U16540 (N_16540,N_14510,N_14802);
nand U16541 (N_16541,N_15150,N_15009);
nand U16542 (N_16542,N_14545,N_14990);
xor U16543 (N_16543,N_15149,N_15198);
nand U16544 (N_16544,N_14880,N_15517);
nor U16545 (N_16545,N_14824,N_14610);
nor U16546 (N_16546,N_15573,N_15526);
xnor U16547 (N_16547,N_14678,N_14646);
or U16548 (N_16548,N_15290,N_15476);
xnor U16549 (N_16549,N_14818,N_15285);
or U16550 (N_16550,N_14807,N_15209);
or U16551 (N_16551,N_15051,N_15107);
or U16552 (N_16552,N_14760,N_15126);
and U16553 (N_16553,N_14621,N_14616);
or U16554 (N_16554,N_15105,N_15507);
nand U16555 (N_16555,N_15137,N_15599);
and U16556 (N_16556,N_15111,N_15143);
nor U16557 (N_16557,N_14609,N_14970);
nor U16558 (N_16558,N_14601,N_15426);
or U16559 (N_16559,N_14508,N_14877);
or U16560 (N_16560,N_14546,N_14957);
nor U16561 (N_16561,N_15579,N_15393);
nor U16562 (N_16562,N_14470,N_14559);
and U16563 (N_16563,N_14685,N_14830);
nor U16564 (N_16564,N_14473,N_14421);
nand U16565 (N_16565,N_14658,N_14656);
and U16566 (N_16566,N_14663,N_15100);
xor U16567 (N_16567,N_15532,N_15463);
xor U16568 (N_16568,N_14479,N_15376);
xnor U16569 (N_16569,N_14970,N_14791);
xnor U16570 (N_16570,N_14728,N_15441);
and U16571 (N_16571,N_15261,N_15167);
or U16572 (N_16572,N_14962,N_14504);
xnor U16573 (N_16573,N_14854,N_14989);
xor U16574 (N_16574,N_15446,N_14685);
xor U16575 (N_16575,N_15595,N_15582);
and U16576 (N_16576,N_14680,N_14592);
or U16577 (N_16577,N_14851,N_15193);
nand U16578 (N_16578,N_15537,N_14596);
nor U16579 (N_16579,N_15069,N_15438);
nand U16580 (N_16580,N_15530,N_15088);
nand U16581 (N_16581,N_14858,N_15222);
nand U16582 (N_16582,N_15451,N_14426);
or U16583 (N_16583,N_14773,N_15547);
nor U16584 (N_16584,N_14608,N_14456);
and U16585 (N_16585,N_14956,N_15102);
nor U16586 (N_16586,N_14894,N_14717);
nor U16587 (N_16587,N_15295,N_14475);
nand U16588 (N_16588,N_14734,N_15326);
xor U16589 (N_16589,N_14556,N_15031);
nand U16590 (N_16590,N_15305,N_14402);
nor U16591 (N_16591,N_15406,N_14897);
xnor U16592 (N_16592,N_14669,N_15547);
xor U16593 (N_16593,N_15539,N_15516);
nor U16594 (N_16594,N_14521,N_14499);
nor U16595 (N_16595,N_15006,N_14584);
and U16596 (N_16596,N_15023,N_15463);
nand U16597 (N_16597,N_14460,N_14737);
or U16598 (N_16598,N_14726,N_15292);
and U16599 (N_16599,N_15327,N_14558);
xor U16600 (N_16600,N_14962,N_14915);
nand U16601 (N_16601,N_14869,N_15518);
xor U16602 (N_16602,N_15218,N_15419);
and U16603 (N_16603,N_15179,N_14774);
or U16604 (N_16604,N_15132,N_15028);
nor U16605 (N_16605,N_15390,N_15320);
nand U16606 (N_16606,N_14418,N_15203);
nand U16607 (N_16607,N_15170,N_15069);
and U16608 (N_16608,N_14954,N_15258);
and U16609 (N_16609,N_14851,N_14723);
or U16610 (N_16610,N_14664,N_15031);
nor U16611 (N_16611,N_15451,N_14895);
nor U16612 (N_16612,N_14679,N_14891);
nor U16613 (N_16613,N_15534,N_14963);
nand U16614 (N_16614,N_14469,N_14681);
or U16615 (N_16615,N_15483,N_15070);
xnor U16616 (N_16616,N_15394,N_14758);
xnor U16617 (N_16617,N_15273,N_14624);
xnor U16618 (N_16618,N_14958,N_14847);
and U16619 (N_16619,N_15040,N_14761);
xnor U16620 (N_16620,N_15439,N_14624);
nand U16621 (N_16621,N_15355,N_14672);
or U16622 (N_16622,N_15336,N_15196);
or U16623 (N_16623,N_14465,N_15000);
nand U16624 (N_16624,N_14430,N_15354);
nor U16625 (N_16625,N_14812,N_15499);
and U16626 (N_16626,N_14537,N_14850);
or U16627 (N_16627,N_14777,N_15175);
xor U16628 (N_16628,N_14434,N_14909);
or U16629 (N_16629,N_15543,N_15341);
nand U16630 (N_16630,N_15114,N_14595);
nand U16631 (N_16631,N_14629,N_14410);
nand U16632 (N_16632,N_14547,N_15484);
nand U16633 (N_16633,N_14680,N_15424);
or U16634 (N_16634,N_15502,N_14440);
or U16635 (N_16635,N_14518,N_15479);
and U16636 (N_16636,N_15517,N_15214);
nor U16637 (N_16637,N_14528,N_14790);
and U16638 (N_16638,N_15510,N_14706);
xor U16639 (N_16639,N_14411,N_14519);
xor U16640 (N_16640,N_15247,N_14852);
xnor U16641 (N_16641,N_14939,N_15510);
and U16642 (N_16642,N_15558,N_15345);
xor U16643 (N_16643,N_14995,N_15420);
xor U16644 (N_16644,N_15348,N_14450);
or U16645 (N_16645,N_15291,N_15201);
xnor U16646 (N_16646,N_15561,N_14495);
xnor U16647 (N_16647,N_15211,N_14507);
nor U16648 (N_16648,N_15203,N_15536);
nor U16649 (N_16649,N_14856,N_14790);
nor U16650 (N_16650,N_15430,N_14675);
nor U16651 (N_16651,N_14600,N_15541);
xor U16652 (N_16652,N_15445,N_14583);
or U16653 (N_16653,N_14779,N_14441);
or U16654 (N_16654,N_15408,N_14490);
nor U16655 (N_16655,N_15287,N_14450);
and U16656 (N_16656,N_15582,N_15519);
nand U16657 (N_16657,N_14860,N_14554);
or U16658 (N_16658,N_15313,N_14709);
or U16659 (N_16659,N_15077,N_15217);
nand U16660 (N_16660,N_14661,N_15110);
and U16661 (N_16661,N_15252,N_14617);
and U16662 (N_16662,N_14429,N_15354);
xnor U16663 (N_16663,N_15194,N_15390);
xor U16664 (N_16664,N_14844,N_15481);
and U16665 (N_16665,N_14833,N_15143);
nor U16666 (N_16666,N_14877,N_14714);
nand U16667 (N_16667,N_15239,N_14669);
nor U16668 (N_16668,N_15135,N_15425);
nor U16669 (N_16669,N_15594,N_14544);
xnor U16670 (N_16670,N_15161,N_15400);
or U16671 (N_16671,N_15309,N_14750);
xor U16672 (N_16672,N_14689,N_14710);
xnor U16673 (N_16673,N_15085,N_14695);
nor U16674 (N_16674,N_14872,N_15462);
xnor U16675 (N_16675,N_14920,N_14440);
nand U16676 (N_16676,N_14884,N_15248);
or U16677 (N_16677,N_14952,N_15186);
nand U16678 (N_16678,N_14650,N_15599);
nor U16679 (N_16679,N_15370,N_15221);
and U16680 (N_16680,N_14833,N_15308);
xnor U16681 (N_16681,N_15563,N_14773);
and U16682 (N_16682,N_15039,N_14713);
nand U16683 (N_16683,N_15245,N_14659);
nor U16684 (N_16684,N_14946,N_14683);
xor U16685 (N_16685,N_14783,N_15237);
or U16686 (N_16686,N_14545,N_15066);
nand U16687 (N_16687,N_15539,N_14580);
xor U16688 (N_16688,N_14529,N_15225);
nand U16689 (N_16689,N_15244,N_14988);
or U16690 (N_16690,N_14531,N_15407);
and U16691 (N_16691,N_14640,N_15165);
or U16692 (N_16692,N_15099,N_15501);
and U16693 (N_16693,N_15517,N_15479);
or U16694 (N_16694,N_15228,N_14682);
and U16695 (N_16695,N_15401,N_15434);
nand U16696 (N_16696,N_14943,N_15549);
or U16697 (N_16697,N_14604,N_14744);
and U16698 (N_16698,N_15437,N_15501);
nor U16699 (N_16699,N_15183,N_15257);
nor U16700 (N_16700,N_15037,N_15048);
nor U16701 (N_16701,N_14863,N_15562);
xnor U16702 (N_16702,N_15027,N_15230);
nor U16703 (N_16703,N_14484,N_14682);
and U16704 (N_16704,N_15455,N_15026);
nand U16705 (N_16705,N_15293,N_14569);
xnor U16706 (N_16706,N_14694,N_14546);
xnor U16707 (N_16707,N_14440,N_14952);
and U16708 (N_16708,N_14649,N_15024);
or U16709 (N_16709,N_14928,N_15299);
or U16710 (N_16710,N_14404,N_14821);
xnor U16711 (N_16711,N_14657,N_14495);
and U16712 (N_16712,N_15169,N_14537);
xnor U16713 (N_16713,N_14989,N_15194);
nor U16714 (N_16714,N_15173,N_14826);
or U16715 (N_16715,N_15401,N_14827);
xor U16716 (N_16716,N_14649,N_15208);
or U16717 (N_16717,N_15330,N_15497);
nand U16718 (N_16718,N_15468,N_14401);
or U16719 (N_16719,N_14426,N_15233);
and U16720 (N_16720,N_15449,N_15039);
xor U16721 (N_16721,N_15237,N_15326);
xor U16722 (N_16722,N_15513,N_15008);
and U16723 (N_16723,N_15171,N_14664);
xnor U16724 (N_16724,N_15048,N_15562);
nand U16725 (N_16725,N_15297,N_14420);
nand U16726 (N_16726,N_15346,N_15282);
nor U16727 (N_16727,N_14570,N_14926);
nand U16728 (N_16728,N_15494,N_15144);
nor U16729 (N_16729,N_14714,N_15424);
nand U16730 (N_16730,N_15434,N_15037);
nand U16731 (N_16731,N_15422,N_15467);
and U16732 (N_16732,N_14465,N_14563);
nand U16733 (N_16733,N_15162,N_14715);
xor U16734 (N_16734,N_15453,N_15076);
nand U16735 (N_16735,N_14807,N_15293);
xnor U16736 (N_16736,N_14863,N_15546);
nand U16737 (N_16737,N_15010,N_14664);
xor U16738 (N_16738,N_15206,N_15205);
and U16739 (N_16739,N_14542,N_14970);
and U16740 (N_16740,N_15188,N_14429);
xnor U16741 (N_16741,N_14642,N_14665);
and U16742 (N_16742,N_15232,N_14675);
xor U16743 (N_16743,N_14926,N_15135);
nor U16744 (N_16744,N_14850,N_15248);
and U16745 (N_16745,N_15351,N_14423);
or U16746 (N_16746,N_14854,N_15033);
nand U16747 (N_16747,N_14924,N_15274);
nor U16748 (N_16748,N_14445,N_15423);
or U16749 (N_16749,N_14863,N_15372);
nand U16750 (N_16750,N_15051,N_15253);
or U16751 (N_16751,N_14657,N_15173);
nand U16752 (N_16752,N_14823,N_14651);
nor U16753 (N_16753,N_14751,N_15052);
nand U16754 (N_16754,N_15433,N_14671);
and U16755 (N_16755,N_15070,N_15555);
and U16756 (N_16756,N_15101,N_15243);
nor U16757 (N_16757,N_15368,N_15543);
nand U16758 (N_16758,N_14781,N_15481);
and U16759 (N_16759,N_15015,N_15394);
nor U16760 (N_16760,N_15155,N_14964);
nor U16761 (N_16761,N_14820,N_15054);
xor U16762 (N_16762,N_15451,N_14988);
xor U16763 (N_16763,N_15490,N_14835);
nor U16764 (N_16764,N_15214,N_14405);
or U16765 (N_16765,N_15279,N_15160);
xnor U16766 (N_16766,N_14677,N_15317);
or U16767 (N_16767,N_15492,N_14976);
nand U16768 (N_16768,N_14417,N_14702);
nor U16769 (N_16769,N_14727,N_14529);
or U16770 (N_16770,N_15068,N_15366);
or U16771 (N_16771,N_15208,N_15119);
xor U16772 (N_16772,N_15169,N_15432);
nor U16773 (N_16773,N_15188,N_14793);
xor U16774 (N_16774,N_15575,N_15568);
nor U16775 (N_16775,N_14816,N_15320);
and U16776 (N_16776,N_15496,N_15510);
nor U16777 (N_16777,N_15556,N_15226);
nor U16778 (N_16778,N_15002,N_15143);
nand U16779 (N_16779,N_14790,N_14795);
or U16780 (N_16780,N_15589,N_15484);
nand U16781 (N_16781,N_14984,N_14679);
nand U16782 (N_16782,N_15534,N_15381);
xor U16783 (N_16783,N_15561,N_14655);
xnor U16784 (N_16784,N_15498,N_15046);
nand U16785 (N_16785,N_14451,N_14932);
xor U16786 (N_16786,N_15483,N_15298);
or U16787 (N_16787,N_14553,N_15365);
nor U16788 (N_16788,N_15002,N_14501);
nand U16789 (N_16789,N_14672,N_15572);
or U16790 (N_16790,N_14681,N_15030);
or U16791 (N_16791,N_15035,N_15314);
and U16792 (N_16792,N_14911,N_15490);
nor U16793 (N_16793,N_14628,N_14774);
nor U16794 (N_16794,N_15161,N_15480);
nor U16795 (N_16795,N_14684,N_14655);
xor U16796 (N_16796,N_14502,N_14406);
and U16797 (N_16797,N_15589,N_14595);
xor U16798 (N_16798,N_15556,N_15066);
nor U16799 (N_16799,N_15083,N_14942);
nand U16800 (N_16800,N_16511,N_15888);
nor U16801 (N_16801,N_16151,N_15794);
or U16802 (N_16802,N_16787,N_16220);
xnor U16803 (N_16803,N_16117,N_15716);
and U16804 (N_16804,N_15873,N_16425);
or U16805 (N_16805,N_16556,N_15711);
nor U16806 (N_16806,N_16119,N_16644);
or U16807 (N_16807,N_15670,N_15789);
xor U16808 (N_16808,N_16346,N_15936);
or U16809 (N_16809,N_15967,N_16040);
nand U16810 (N_16810,N_16638,N_15862);
xor U16811 (N_16811,N_15790,N_16774);
xor U16812 (N_16812,N_16351,N_15774);
nand U16813 (N_16813,N_16369,N_15658);
and U16814 (N_16814,N_15831,N_15787);
xor U16815 (N_16815,N_16715,N_16669);
nand U16816 (N_16816,N_15767,N_16374);
xor U16817 (N_16817,N_16540,N_16334);
nand U16818 (N_16818,N_15786,N_15970);
nor U16819 (N_16819,N_16300,N_16409);
nor U16820 (N_16820,N_15760,N_15610);
nor U16821 (N_16821,N_16578,N_15900);
xnor U16822 (N_16822,N_16637,N_15602);
nand U16823 (N_16823,N_16587,N_16663);
nor U16824 (N_16824,N_16470,N_16252);
xnor U16825 (N_16825,N_15889,N_15800);
or U16826 (N_16826,N_16089,N_15751);
or U16827 (N_16827,N_15994,N_16665);
nand U16828 (N_16828,N_15841,N_15962);
and U16829 (N_16829,N_16388,N_16284);
or U16830 (N_16830,N_16130,N_16543);
or U16831 (N_16831,N_16611,N_15838);
nor U16832 (N_16832,N_15980,N_16491);
nand U16833 (N_16833,N_16473,N_16791);
xor U16834 (N_16834,N_16128,N_15777);
nand U16835 (N_16835,N_16070,N_16083);
nor U16836 (N_16836,N_16147,N_15818);
nand U16837 (N_16837,N_16347,N_15926);
and U16838 (N_16838,N_15948,N_16745);
or U16839 (N_16839,N_15852,N_15817);
nor U16840 (N_16840,N_16646,N_15915);
nor U16841 (N_16841,N_16521,N_16358);
nand U16842 (N_16842,N_16135,N_16269);
and U16843 (N_16843,N_16495,N_15807);
nor U16844 (N_16844,N_16559,N_16653);
xnor U16845 (N_16845,N_16797,N_15880);
nor U16846 (N_16846,N_16176,N_16315);
xor U16847 (N_16847,N_16144,N_15981);
and U16848 (N_16848,N_15690,N_15867);
and U16849 (N_16849,N_15848,N_16529);
nor U16850 (N_16850,N_16668,N_16282);
or U16851 (N_16851,N_16722,N_16615);
nor U16852 (N_16852,N_15735,N_15979);
nor U16853 (N_16853,N_16339,N_15605);
nand U16854 (N_16854,N_16353,N_15683);
and U16855 (N_16855,N_16519,N_15886);
and U16856 (N_16856,N_16008,N_16068);
nor U16857 (N_16857,N_15825,N_15982);
or U16858 (N_16858,N_16253,N_16601);
nor U16859 (N_16859,N_15755,N_16503);
or U16860 (N_16860,N_16768,N_16712);
nand U16861 (N_16861,N_15727,N_16410);
nand U16862 (N_16862,N_16380,N_16430);
or U16863 (N_16863,N_16769,N_16591);
and U16864 (N_16864,N_16683,N_16733);
xor U16865 (N_16865,N_15650,N_16467);
xnor U16866 (N_16866,N_16293,N_16407);
xnor U16867 (N_16867,N_15703,N_15903);
nand U16868 (N_16868,N_15847,N_15715);
xnor U16869 (N_16869,N_16061,N_16671);
nor U16870 (N_16870,N_16513,N_16568);
xnor U16871 (N_16871,N_15770,N_16654);
nor U16872 (N_16872,N_16699,N_16105);
or U16873 (N_16873,N_16342,N_16716);
and U16874 (N_16874,N_16209,N_16181);
nor U16875 (N_16875,N_16270,N_16041);
nor U16876 (N_16876,N_15977,N_15698);
nand U16877 (N_16877,N_16240,N_15608);
nand U16878 (N_16878,N_15953,N_15733);
nor U16879 (N_16879,N_16448,N_16444);
nand U16880 (N_16880,N_16561,N_16583);
or U16881 (N_16881,N_16263,N_16162);
or U16882 (N_16882,N_16596,N_16034);
and U16883 (N_16883,N_16206,N_16594);
or U16884 (N_16884,N_16799,N_16152);
nor U16885 (N_16885,N_16186,N_15671);
xnor U16886 (N_16886,N_16316,N_15674);
nor U16887 (N_16887,N_16365,N_16143);
and U16888 (N_16888,N_16303,N_15891);
nor U16889 (N_16889,N_16087,N_15828);
nor U16890 (N_16890,N_16394,N_16558);
nor U16891 (N_16891,N_16493,N_16438);
nor U16892 (N_16892,N_15944,N_16291);
nand U16893 (N_16893,N_16516,N_16554);
and U16894 (N_16894,N_16238,N_15637);
xnor U16895 (N_16895,N_16221,N_15945);
nor U16896 (N_16896,N_16798,N_15752);
and U16897 (N_16897,N_16602,N_15662);
xor U16898 (N_16898,N_16058,N_16341);
or U16899 (N_16899,N_15990,N_16681);
or U16900 (N_16900,N_16792,N_16292);
or U16901 (N_16901,N_15866,N_15611);
nor U16902 (N_16902,N_16782,N_16166);
or U16903 (N_16903,N_15647,N_16426);
xnor U16904 (N_16904,N_16728,N_16645);
nand U16905 (N_16905,N_16532,N_15809);
or U16906 (N_16906,N_16113,N_16533);
and U16907 (N_16907,N_16161,N_16667);
xnor U16908 (N_16908,N_16729,N_16406);
and U16909 (N_16909,N_16738,N_16599);
nor U16910 (N_16910,N_16753,N_15991);
nor U16911 (N_16911,N_16458,N_16078);
or U16912 (N_16912,N_16014,N_15890);
or U16913 (N_16913,N_16028,N_16154);
nand U16914 (N_16914,N_16188,N_15859);
nor U16915 (N_16915,N_16204,N_15988);
nand U16916 (N_16916,N_16329,N_15968);
or U16917 (N_16917,N_15917,N_16643);
nor U16918 (N_16918,N_16052,N_16377);
nand U16919 (N_16919,N_16544,N_16441);
xnor U16920 (N_16920,N_16384,N_15844);
xnor U16921 (N_16921,N_16035,N_16060);
xor U16922 (N_16922,N_16746,N_16603);
nor U16923 (N_16923,N_16067,N_16709);
and U16924 (N_16924,N_15628,N_15850);
nor U16925 (N_16925,N_16126,N_15802);
nand U16926 (N_16926,N_15748,N_16691);
nand U16927 (N_16927,N_15745,N_16632);
and U16928 (N_16928,N_15705,N_15797);
and U16929 (N_16929,N_15680,N_16042);
or U16930 (N_16930,N_15734,N_15899);
nor U16931 (N_16931,N_15849,N_16542);
nor U16932 (N_16932,N_16099,N_16283);
or U16933 (N_16933,N_16720,N_16436);
nor U16934 (N_16934,N_16069,N_15798);
nand U16935 (N_16935,N_15618,N_15927);
nand U16936 (N_16936,N_16247,N_16148);
nor U16937 (N_16937,N_16555,N_16451);
xnor U16938 (N_16938,N_16701,N_16621);
or U16939 (N_16939,N_16318,N_15972);
and U16940 (N_16940,N_15835,N_16497);
nor U16941 (N_16941,N_16224,N_15644);
or U16942 (N_16942,N_16666,N_15858);
nand U16943 (N_16943,N_15692,N_16640);
nand U16944 (N_16944,N_16138,N_16309);
and U16945 (N_16945,N_16331,N_15935);
nor U16946 (N_16946,N_16415,N_16423);
nor U16947 (N_16947,N_16313,N_15771);
nand U16948 (N_16948,N_15805,N_16338);
nand U16949 (N_16949,N_15998,N_15791);
nor U16950 (N_16950,N_15648,N_15973);
nand U16951 (N_16951,N_16676,N_15892);
nand U16952 (N_16952,N_16770,N_15877);
xnor U16953 (N_16953,N_16781,N_16299);
nor U16954 (N_16954,N_16534,N_16790);
nor U16955 (N_16955,N_16110,N_15766);
or U16956 (N_16956,N_16127,N_16043);
xor U16957 (N_16957,N_16305,N_16675);
nor U16958 (N_16958,N_16474,N_16362);
xnor U16959 (N_16959,N_16017,N_16368);
and U16960 (N_16960,N_16698,N_15782);
or U16961 (N_16961,N_15952,N_16589);
and U16962 (N_16962,N_16562,N_16477);
nor U16963 (N_16963,N_16490,N_16420);
nand U16964 (N_16964,N_16761,N_15969);
or U16965 (N_16965,N_16149,N_16226);
or U16966 (N_16966,N_16055,N_15642);
nor U16967 (N_16967,N_15960,N_16582);
nand U16968 (N_16968,N_16585,N_16475);
and U16969 (N_16969,N_15621,N_15775);
xor U16970 (N_16970,N_15939,N_16672);
or U16971 (N_16971,N_16708,N_15653);
nor U16972 (N_16972,N_15660,N_16635);
and U16973 (N_16973,N_16694,N_16429);
nor U16974 (N_16974,N_15761,N_16222);
nor U16975 (N_16975,N_16743,N_16704);
and U16976 (N_16976,N_15712,N_16661);
or U16977 (N_16977,N_16277,N_16446);
or U16978 (N_16978,N_16619,N_15676);
or U16979 (N_16979,N_15630,N_16000);
or U16980 (N_16980,N_15768,N_16169);
nand U16981 (N_16981,N_15870,N_16725);
xnor U16982 (N_16982,N_16378,N_16649);
nor U16983 (N_16983,N_15928,N_16785);
nand U16984 (N_16984,N_16695,N_15744);
and U16985 (N_16985,N_16245,N_16392);
xor U16986 (N_16986,N_15933,N_16595);
or U16987 (N_16987,N_16590,N_16766);
xnor U16988 (N_16988,N_15930,N_16518);
or U16989 (N_16989,N_15914,N_16314);
nor U16990 (N_16990,N_16376,N_16740);
nor U16991 (N_16991,N_16626,N_16742);
xnor U16992 (N_16992,N_15638,N_16167);
or U16993 (N_16993,N_16597,N_15978);
nand U16994 (N_16994,N_15736,N_15822);
nand U16995 (N_16995,N_16025,N_16622);
or U16996 (N_16996,N_16480,N_16525);
xor U16997 (N_16997,N_15836,N_15942);
xnor U16998 (N_16998,N_16697,N_16326);
xnor U16999 (N_16999,N_16756,N_16005);
and U17000 (N_17000,N_16074,N_16786);
and U17001 (N_17001,N_16294,N_16100);
xor U17002 (N_17002,N_16379,N_15613);
or U17003 (N_17003,N_15905,N_16348);
and U17004 (N_17004,N_16302,N_16572);
and U17005 (N_17005,N_16153,N_16400);
nand U17006 (N_17006,N_16610,N_16424);
nor U17007 (N_17007,N_16512,N_16483);
and U17008 (N_17008,N_16612,N_16553);
or U17009 (N_17009,N_16628,N_15937);
nor U17010 (N_17010,N_16469,N_16581);
nand U17011 (N_17011,N_15857,N_15719);
or U17012 (N_17012,N_16662,N_16627);
nand U17013 (N_17013,N_16327,N_16616);
nand U17014 (N_17014,N_16489,N_16445);
nand U17015 (N_17015,N_16031,N_16051);
and U17016 (N_17016,N_15754,N_16271);
or U17017 (N_17017,N_16350,N_16796);
or U17018 (N_17018,N_16349,N_15776);
nor U17019 (N_17019,N_15806,N_15943);
and U17020 (N_17020,N_16009,N_15781);
or U17021 (N_17021,N_15722,N_16393);
or U17022 (N_17022,N_16447,N_16386);
or U17023 (N_17023,N_16090,N_16752);
or U17024 (N_17024,N_16404,N_16232);
or U17025 (N_17025,N_15827,N_15656);
nand U17026 (N_17026,N_16208,N_15718);
or U17027 (N_17027,N_15645,N_15851);
nor U17028 (N_17028,N_15758,N_16579);
or U17029 (N_17029,N_16565,N_15996);
nor U17030 (N_17030,N_15646,N_15992);
and U17031 (N_17031,N_15750,N_16175);
nor U17032 (N_17032,N_15779,N_16098);
xor U17033 (N_17033,N_16793,N_15919);
or U17034 (N_17034,N_16223,N_16629);
nor U17035 (N_17035,N_15629,N_16026);
nor U17036 (N_17036,N_16333,N_15778);
xnor U17037 (N_17037,N_16093,N_15856);
xnor U17038 (N_17038,N_15985,N_16755);
and U17039 (N_17039,N_16703,N_16084);
and U17040 (N_17040,N_16256,N_16211);
xnor U17041 (N_17041,N_15834,N_15631);
and U17042 (N_17042,N_16268,N_15704);
and U17043 (N_17043,N_16094,N_16539);
or U17044 (N_17044,N_16145,N_16399);
xor U17045 (N_17045,N_16767,N_16449);
xor U17046 (N_17046,N_15976,N_15821);
or U17047 (N_17047,N_16260,N_16139);
nor U17048 (N_17048,N_16702,N_16021);
or U17049 (N_17049,N_16775,N_15708);
xor U17050 (N_17050,N_16039,N_15869);
nor U17051 (N_17051,N_16494,N_15863);
or U17052 (N_17052,N_15635,N_16788);
nor U17053 (N_17053,N_16107,N_16259);
or U17054 (N_17054,N_16434,N_16295);
xnor U17055 (N_17055,N_16308,N_16194);
nor U17056 (N_17056,N_16297,N_16502);
nand U17057 (N_17057,N_15672,N_16359);
nand U17058 (N_17058,N_16080,N_16484);
xor U17059 (N_17059,N_16749,N_16246);
and U17060 (N_17060,N_16375,N_16567);
nor U17061 (N_17061,N_15614,N_16112);
xor U17062 (N_17062,N_16296,N_15643);
and U17063 (N_17063,N_16046,N_16433);
nand U17064 (N_17064,N_15951,N_16273);
nor U17065 (N_17065,N_15986,N_16383);
nand U17066 (N_17066,N_16779,N_15709);
nor U17067 (N_17067,N_16225,N_15684);
nor U17068 (N_17068,N_15729,N_15904);
or U17069 (N_17069,N_15609,N_16759);
or U17070 (N_17070,N_15925,N_16789);
and U17071 (N_17071,N_16257,N_16281);
xor U17072 (N_17072,N_16170,N_15947);
nor U17073 (N_17073,N_16057,N_15804);
nor U17074 (N_17074,N_15941,N_16241);
xor U17075 (N_17075,N_15907,N_15659);
nor U17076 (N_17076,N_16064,N_15842);
nor U17077 (N_17077,N_16506,N_16537);
and U17078 (N_17078,N_16442,N_16372);
xnor U17079 (N_17079,N_15860,N_16421);
nand U17080 (N_17080,N_15607,N_16593);
nand U17081 (N_17081,N_16413,N_16317);
nor U17082 (N_17082,N_16048,N_15639);
and U17083 (N_17083,N_16478,N_16464);
nand U17084 (N_17084,N_16054,N_16213);
xor U17085 (N_17085,N_15966,N_16357);
xor U17086 (N_17086,N_16726,N_16011);
and U17087 (N_17087,N_16509,N_15932);
or U17088 (N_17088,N_15765,N_16403);
and U17089 (N_17089,N_16624,N_16250);
or U17090 (N_17090,N_16706,N_16229);
or U17091 (N_17091,N_16165,N_16411);
xor U17092 (N_17092,N_16732,N_16307);
or U17093 (N_17093,N_16015,N_16457);
or U17094 (N_17094,N_16625,N_16355);
and U17095 (N_17095,N_16140,N_15934);
and U17096 (N_17096,N_15693,N_16598);
nand U17097 (N_17097,N_16718,N_16711);
nor U17098 (N_17098,N_16180,N_16385);
nor U17099 (N_17099,N_15724,N_15897);
or U17100 (N_17100,N_16724,N_15713);
and U17101 (N_17101,N_16784,N_16685);
or U17102 (N_17102,N_15701,N_16101);
and U17103 (N_17103,N_15746,N_15792);
xnor U17104 (N_17104,N_16416,N_16007);
and U17105 (N_17105,N_16199,N_15922);
and U17106 (N_17106,N_15799,N_15987);
xnor U17107 (N_17107,N_15901,N_16501);
or U17108 (N_17108,N_15938,N_16546);
xnor U17109 (N_17109,N_15652,N_16700);
and U17110 (N_17110,N_16202,N_16574);
or U17111 (N_17111,N_16045,N_16195);
xnor U17112 (N_17112,N_15906,N_16103);
or U17113 (N_17113,N_16038,N_16686);
nand U17114 (N_17114,N_16343,N_16634);
nor U17115 (N_17115,N_15853,N_15695);
nor U17116 (N_17116,N_15689,N_15772);
nor U17117 (N_17117,N_16472,N_15895);
or U17118 (N_17118,N_16431,N_16736);
xor U17119 (N_17119,N_16228,N_15974);
nor U17120 (N_17120,N_15625,N_16677);
or U17121 (N_17121,N_16254,N_15661);
or U17122 (N_17122,N_15902,N_16563);
nor U17123 (N_17123,N_15833,N_16397);
xnor U17124 (N_17124,N_16573,N_16535);
nor U17125 (N_17125,N_15997,N_15739);
nor U17126 (N_17126,N_16575,N_16412);
nand U17127 (N_17127,N_15824,N_16456);
nor U17128 (N_17128,N_15819,N_16655);
nor U17129 (N_17129,N_15923,N_16122);
and U17130 (N_17130,N_15989,N_16751);
nor U17131 (N_17131,N_16301,N_16123);
xor U17132 (N_17132,N_15871,N_16033);
nor U17133 (N_17133,N_16298,N_16095);
and U17134 (N_17134,N_16737,N_16023);
xor U17135 (N_17135,N_16580,N_16750);
xor U17136 (N_17136,N_15959,N_16227);
or U17137 (N_17137,N_16030,N_15725);
nor U17138 (N_17138,N_16692,N_16003);
xor U17139 (N_17139,N_16547,N_16248);
nand U17140 (N_17140,N_16124,N_16747);
nand U17141 (N_17141,N_15756,N_16371);
or U17142 (N_17142,N_16586,N_16549);
and U17143 (N_17143,N_16133,N_16522);
nor U17144 (N_17144,N_16363,N_16288);
or U17145 (N_17145,N_16177,N_15881);
nand U17146 (N_17146,N_16408,N_16673);
or U17147 (N_17147,N_16557,N_15971);
xor U17148 (N_17148,N_16462,N_16022);
or U17149 (N_17149,N_16244,N_15893);
or U17150 (N_17150,N_16114,N_16013);
xnor U17151 (N_17151,N_16739,N_16432);
xor U17152 (N_17152,N_16461,N_16066);
and U17153 (N_17153,N_16510,N_15872);
xnor U17154 (N_17154,N_16193,N_16207);
xor U17155 (N_17155,N_16754,N_16658);
xor U17156 (N_17156,N_16053,N_16391);
xor U17157 (N_17157,N_15780,N_15949);
xnor U17158 (N_17158,N_16325,N_16182);
nand U17159 (N_17159,N_16163,N_16024);
nor U17160 (N_17160,N_15706,N_15688);
and U17161 (N_17161,N_16541,N_15950);
xnor U17162 (N_17162,N_15911,N_16443);
nor U17163 (N_17163,N_16530,N_16029);
nand U17164 (N_17164,N_16289,N_15728);
nand U17165 (N_17165,N_16748,N_15679);
nor U17166 (N_17166,N_16352,N_15633);
nand U17167 (N_17167,N_16641,N_15921);
and U17168 (N_17168,N_15908,N_16336);
nand U17169 (N_17169,N_16255,N_15975);
nor U17170 (N_17170,N_16092,N_15731);
nor U17171 (N_17171,N_16734,N_16659);
nor U17172 (N_17172,N_16146,N_15784);
or U17173 (N_17173,N_16526,N_15983);
nor U17174 (N_17174,N_16075,N_15634);
nand U17175 (N_17175,N_16648,N_16486);
nor U17176 (N_17176,N_15811,N_16111);
or U17177 (N_17177,N_15603,N_16552);
and U17178 (N_17178,N_16016,N_16500);
xnor U17179 (N_17179,N_15763,N_16536);
nand U17180 (N_17180,N_16142,N_16262);
xor U17181 (N_17181,N_16560,N_15940);
or U17182 (N_17182,N_16159,N_15649);
or U17183 (N_17183,N_15875,N_16620);
nand U17184 (N_17184,N_16687,N_15861);
nor U17185 (N_17185,N_16082,N_15846);
nor U17186 (N_17186,N_16717,N_16498);
xnor U17187 (N_17187,N_15796,N_16231);
xnor U17188 (N_17188,N_16488,N_16218);
or U17189 (N_17189,N_16319,N_16088);
xor U17190 (N_17190,N_16680,N_16056);
xnor U17191 (N_17191,N_15788,N_16592);
and U17192 (N_17192,N_16249,N_15874);
xnor U17193 (N_17193,N_16453,N_16304);
nand U17194 (N_17194,N_16427,N_16608);
or U17195 (N_17195,N_16481,N_16201);
or U17196 (N_17196,N_16335,N_16373);
nor U17197 (N_17197,N_16523,N_16214);
and U17198 (N_17198,N_15795,N_16631);
nor U17199 (N_17199,N_16689,N_16763);
nor U17200 (N_17200,N_16515,N_16600);
xor U17201 (N_17201,N_15606,N_16670);
nor U17202 (N_17202,N_16120,N_16485);
nor U17203 (N_17203,N_15954,N_16280);
or U17204 (N_17204,N_16002,N_15747);
nor U17205 (N_17205,N_15696,N_15843);
nor U17206 (N_17206,N_16566,N_16460);
and U17207 (N_17207,N_15909,N_16604);
nor U17208 (N_17208,N_16037,N_16109);
nand U17209 (N_17209,N_16636,N_15687);
xor U17210 (N_17210,N_16266,N_16310);
or U17211 (N_17211,N_16027,N_15616);
and U17212 (N_17212,N_15612,N_16577);
xor U17213 (N_17213,N_16131,N_16215);
nor U17214 (N_17214,N_16360,N_16794);
or U17215 (N_17215,N_15865,N_15812);
and U17216 (N_17216,N_16440,N_16356);
or U17217 (N_17217,N_15783,N_16340);
or U17218 (N_17218,N_16508,N_15686);
and U17219 (N_17219,N_15700,N_16168);
and U17220 (N_17220,N_16435,N_16465);
xor U17221 (N_17221,N_15667,N_15864);
nand U17222 (N_17222,N_15810,N_16234);
or U17223 (N_17223,N_15636,N_16062);
or U17224 (N_17224,N_15965,N_15876);
nand U17225 (N_17225,N_15839,N_15655);
xnor U17226 (N_17226,N_15678,N_16036);
xnor U17227 (N_17227,N_16150,N_16765);
nor U17228 (N_17228,N_15813,N_16191);
xor U17229 (N_17229,N_15657,N_16504);
xnor U17230 (N_17230,N_16450,N_16354);
nor U17231 (N_17231,N_16382,N_16778);
and U17232 (N_17232,N_16097,N_15762);
or U17233 (N_17233,N_16390,N_16306);
xor U17234 (N_17234,N_15855,N_16479);
nor U17235 (N_17235,N_15801,N_16387);
xnor U17236 (N_17236,N_15898,N_16564);
nand U17237 (N_17237,N_15816,N_16570);
nor U17238 (N_17238,N_16290,N_16471);
or U17239 (N_17239,N_15894,N_15918);
nor U17240 (N_17240,N_16267,N_16520);
or U17241 (N_17241,N_15741,N_15883);
or U17242 (N_17242,N_16455,N_16727);
or U17243 (N_17243,N_16311,N_16688);
nor U17244 (N_17244,N_16192,N_15623);
nand U17245 (N_17245,N_16320,N_16286);
and U17246 (N_17246,N_15759,N_16200);
nand U17247 (N_17247,N_15654,N_15619);
and U17248 (N_17248,N_16623,N_16004);
nand U17249 (N_17249,N_16719,N_16337);
nor U17250 (N_17250,N_16705,N_16660);
nor U17251 (N_17251,N_15685,N_16613);
or U17252 (N_17252,N_16414,N_15993);
or U17253 (N_17253,N_16132,N_16721);
and U17254 (N_17254,N_16762,N_15617);
nand U17255 (N_17255,N_15885,N_16428);
and U17256 (N_17256,N_16125,N_16714);
nor U17257 (N_17257,N_16272,N_15879);
xnor U17258 (N_17258,N_16696,N_16398);
nand U17259 (N_17259,N_16459,N_16609);
xor U17260 (N_17260,N_15730,N_16639);
xor U17261 (N_17261,N_15837,N_16012);
nor U17262 (N_17262,N_15720,N_16230);
nand U17263 (N_17263,N_16731,N_16776);
nand U17264 (N_17264,N_16183,N_16744);
and U17265 (N_17265,N_16439,N_16196);
or U17266 (N_17266,N_16548,N_15721);
xor U17267 (N_17267,N_16106,N_15984);
nand U17268 (N_17268,N_15913,N_16086);
nor U17269 (N_17269,N_16020,N_15626);
and U17270 (N_17270,N_16251,N_16179);
nand U17271 (N_17271,N_16287,N_16630);
nor U17272 (N_17272,N_16656,N_16370);
nor U17273 (N_17273,N_16584,N_15615);
xnor U17274 (N_17274,N_16452,N_15714);
xor U17275 (N_17275,N_16758,N_16187);
nand U17276 (N_17276,N_15632,N_15620);
nor U17277 (N_17277,N_15931,N_15995);
xnor U17278 (N_17278,N_15668,N_16032);
nor U17279 (N_17279,N_16773,N_16212);
xor U17280 (N_17280,N_15803,N_15920);
nand U17281 (N_17281,N_16157,N_16527);
or U17282 (N_17282,N_16321,N_16496);
and U17283 (N_17283,N_15929,N_16401);
nor U17284 (N_17284,N_15764,N_16047);
or U17285 (N_17285,N_16239,N_15664);
xnor U17286 (N_17286,N_15815,N_16072);
nor U17287 (N_17287,N_16185,N_16437);
or U17288 (N_17288,N_16102,N_16517);
nor U17289 (N_17289,N_16417,N_15673);
and U17290 (N_17290,N_15832,N_16076);
and U17291 (N_17291,N_16278,N_15749);
and U17292 (N_17292,N_16569,N_16419);
xor U17293 (N_17293,N_15830,N_16395);
nor U17294 (N_17294,N_16693,N_16402);
nand U17295 (N_17295,N_15878,N_16487);
nor U17296 (N_17296,N_16664,N_16236);
or U17297 (N_17297,N_16242,N_16044);
xnor U17298 (N_17298,N_16174,N_16233);
xor U17299 (N_17299,N_16108,N_15814);
or U17300 (N_17300,N_16279,N_16463);
or U17301 (N_17301,N_16531,N_16197);
nor U17302 (N_17302,N_15604,N_16418);
nor U17303 (N_17303,N_16019,N_15710);
or U17304 (N_17304,N_16617,N_16764);
xor U17305 (N_17305,N_15946,N_15743);
and U17306 (N_17306,N_16190,N_16361);
and U17307 (N_17307,N_16614,N_15682);
nand U17308 (N_17308,N_16216,N_16576);
nand U17309 (N_17309,N_16261,N_16650);
or U17310 (N_17310,N_16605,N_15702);
or U17311 (N_17311,N_15916,N_16482);
or U17312 (N_17312,N_16171,N_16757);
nor U17313 (N_17313,N_15666,N_15958);
nand U17314 (N_17314,N_16049,N_16328);
or U17315 (N_17315,N_16723,N_16674);
or U17316 (N_17316,N_15808,N_15726);
nand U17317 (N_17317,N_15912,N_15738);
nor U17318 (N_17318,N_15924,N_16760);
and U17319 (N_17319,N_15845,N_15707);
and U17320 (N_17320,N_16210,N_15961);
nand U17321 (N_17321,N_16073,N_16551);
xnor U17322 (N_17322,N_16505,N_15622);
xor U17323 (N_17323,N_16771,N_16780);
nand U17324 (N_17324,N_16071,N_15665);
and U17325 (N_17325,N_16312,N_16050);
or U17326 (N_17326,N_16006,N_16205);
nand U17327 (N_17327,N_16085,N_16079);
xor U17328 (N_17328,N_16237,N_16730);
nor U17329 (N_17329,N_16783,N_15742);
or U17330 (N_17330,N_16330,N_16466);
nand U17331 (N_17331,N_16366,N_15717);
nand U17332 (N_17332,N_16524,N_16063);
or U17333 (N_17333,N_16499,N_16710);
nor U17334 (N_17334,N_16275,N_15963);
xor U17335 (N_17335,N_16323,N_15840);
nor U17336 (N_17336,N_15854,N_15884);
nor U17337 (N_17337,N_16381,N_16684);
xnor U17338 (N_17338,N_15826,N_16454);
nand U17339 (N_17339,N_15957,N_16189);
or U17340 (N_17340,N_16538,N_16607);
nand U17341 (N_17341,N_16713,N_16476);
or U17342 (N_17342,N_16258,N_15823);
nor U17343 (N_17343,N_16096,N_16571);
or U17344 (N_17344,N_16690,N_16344);
and U17345 (N_17345,N_16345,N_16129);
nor U17346 (N_17346,N_16507,N_15641);
nand U17347 (N_17347,N_15677,N_16322);
nor U17348 (N_17348,N_15868,N_15600);
and U17349 (N_17349,N_15955,N_15740);
nand U17350 (N_17350,N_15640,N_16184);
and U17351 (N_17351,N_16618,N_16172);
or U17352 (N_17352,N_16118,N_15785);
xnor U17353 (N_17353,N_15699,N_15956);
or U17354 (N_17354,N_16115,N_16642);
or U17355 (N_17355,N_16155,N_16264);
nor U17356 (N_17356,N_16243,N_16550);
and U17357 (N_17357,N_16265,N_16652);
nand U17358 (N_17358,N_16158,N_15910);
or U17359 (N_17359,N_15964,N_15793);
xnor U17360 (N_17360,N_16777,N_16010);
xor U17361 (N_17361,N_15624,N_16678);
or U17362 (N_17362,N_16219,N_16682);
nand U17363 (N_17363,N_16178,N_16018);
and U17364 (N_17364,N_15601,N_16364);
xnor U17365 (N_17365,N_16528,N_16468);
and U17366 (N_17366,N_16203,N_16104);
or U17367 (N_17367,N_16741,N_16137);
or U17368 (N_17368,N_16707,N_16795);
nor U17369 (N_17369,N_16173,N_15773);
nor U17370 (N_17370,N_15887,N_16081);
xor U17371 (N_17371,N_15681,N_15669);
and U17372 (N_17372,N_15753,N_15675);
xor U17373 (N_17373,N_16235,N_16492);
and U17374 (N_17374,N_16651,N_16657);
nor U17375 (N_17375,N_15896,N_16091);
or U17376 (N_17376,N_16077,N_15829);
nand U17377 (N_17377,N_15651,N_16332);
nor U17378 (N_17378,N_16001,N_16141);
nand U17379 (N_17379,N_16059,N_15820);
xor U17380 (N_17380,N_16324,N_16285);
xor U17381 (N_17381,N_16389,N_15627);
or U17382 (N_17382,N_16276,N_16198);
and U17383 (N_17383,N_16679,N_16647);
or U17384 (N_17384,N_15757,N_16606);
or U17385 (N_17385,N_16405,N_15999);
or U17386 (N_17386,N_16545,N_16121);
or U17387 (N_17387,N_15769,N_16116);
or U17388 (N_17388,N_16588,N_16514);
xor U17389 (N_17389,N_16160,N_16396);
nand U17390 (N_17390,N_16633,N_16735);
nor U17391 (N_17391,N_15694,N_16217);
nand U17392 (N_17392,N_15732,N_15737);
and U17393 (N_17393,N_16422,N_15691);
or U17394 (N_17394,N_16164,N_16772);
xor U17395 (N_17395,N_16134,N_16274);
xnor U17396 (N_17396,N_15697,N_16156);
nor U17397 (N_17397,N_16136,N_16065);
nor U17398 (N_17398,N_15882,N_15663);
nor U17399 (N_17399,N_16367,N_15723);
nand U17400 (N_17400,N_16569,N_16380);
and U17401 (N_17401,N_16537,N_15856);
nand U17402 (N_17402,N_15655,N_15678);
or U17403 (N_17403,N_16315,N_15889);
xor U17404 (N_17404,N_15815,N_15926);
nor U17405 (N_17405,N_16622,N_16297);
nor U17406 (N_17406,N_15633,N_15936);
xnor U17407 (N_17407,N_16293,N_16041);
or U17408 (N_17408,N_16292,N_16189);
and U17409 (N_17409,N_15826,N_16465);
nand U17410 (N_17410,N_16461,N_15883);
or U17411 (N_17411,N_16042,N_16797);
nor U17412 (N_17412,N_16105,N_16173);
nor U17413 (N_17413,N_16480,N_16660);
and U17414 (N_17414,N_15875,N_16531);
or U17415 (N_17415,N_16222,N_16636);
and U17416 (N_17416,N_16159,N_16054);
xor U17417 (N_17417,N_15832,N_15909);
nor U17418 (N_17418,N_16780,N_16139);
or U17419 (N_17419,N_16364,N_15783);
and U17420 (N_17420,N_16270,N_16136);
xor U17421 (N_17421,N_16016,N_16220);
xnor U17422 (N_17422,N_15611,N_16508);
nand U17423 (N_17423,N_16759,N_15752);
or U17424 (N_17424,N_16277,N_15800);
or U17425 (N_17425,N_15882,N_16305);
xnor U17426 (N_17426,N_16054,N_16515);
or U17427 (N_17427,N_15760,N_16220);
nor U17428 (N_17428,N_16191,N_16629);
xnor U17429 (N_17429,N_16615,N_16432);
nor U17430 (N_17430,N_15863,N_15842);
and U17431 (N_17431,N_16429,N_16565);
xnor U17432 (N_17432,N_15847,N_15794);
nand U17433 (N_17433,N_16008,N_16771);
nor U17434 (N_17434,N_16423,N_16433);
or U17435 (N_17435,N_16350,N_16773);
xor U17436 (N_17436,N_15616,N_15716);
nor U17437 (N_17437,N_15768,N_16751);
nand U17438 (N_17438,N_16635,N_15908);
and U17439 (N_17439,N_15889,N_15900);
nor U17440 (N_17440,N_15606,N_15669);
nand U17441 (N_17441,N_16023,N_15930);
and U17442 (N_17442,N_16187,N_16121);
nor U17443 (N_17443,N_15649,N_16674);
nand U17444 (N_17444,N_16055,N_16694);
xor U17445 (N_17445,N_16659,N_16448);
xnor U17446 (N_17446,N_16712,N_16407);
nand U17447 (N_17447,N_15807,N_16694);
nor U17448 (N_17448,N_15684,N_16049);
and U17449 (N_17449,N_15923,N_16625);
xnor U17450 (N_17450,N_16674,N_16171);
xnor U17451 (N_17451,N_16243,N_16629);
nand U17452 (N_17452,N_15632,N_15847);
or U17453 (N_17453,N_15640,N_16107);
nand U17454 (N_17454,N_16166,N_15743);
and U17455 (N_17455,N_16546,N_16200);
nor U17456 (N_17456,N_16122,N_15655);
or U17457 (N_17457,N_16200,N_15661);
nor U17458 (N_17458,N_16598,N_16137);
and U17459 (N_17459,N_16364,N_16764);
nor U17460 (N_17460,N_16181,N_16675);
and U17461 (N_17461,N_16434,N_15765);
nand U17462 (N_17462,N_15849,N_15901);
nand U17463 (N_17463,N_16044,N_15656);
or U17464 (N_17464,N_16496,N_16561);
or U17465 (N_17465,N_16742,N_16625);
or U17466 (N_17466,N_16336,N_16088);
and U17467 (N_17467,N_16057,N_16330);
or U17468 (N_17468,N_15775,N_16060);
nand U17469 (N_17469,N_15914,N_16446);
or U17470 (N_17470,N_16441,N_16030);
xnor U17471 (N_17471,N_15810,N_16606);
and U17472 (N_17472,N_16259,N_16029);
nand U17473 (N_17473,N_15748,N_15900);
or U17474 (N_17474,N_16680,N_16315);
nor U17475 (N_17475,N_15924,N_15675);
nor U17476 (N_17476,N_16391,N_16374);
nor U17477 (N_17477,N_15711,N_16698);
nor U17478 (N_17478,N_16544,N_16096);
nor U17479 (N_17479,N_16138,N_16500);
and U17480 (N_17480,N_16172,N_16453);
or U17481 (N_17481,N_16503,N_15899);
xor U17482 (N_17482,N_16660,N_15835);
and U17483 (N_17483,N_16315,N_15867);
nor U17484 (N_17484,N_16687,N_16016);
nor U17485 (N_17485,N_16074,N_16622);
nor U17486 (N_17486,N_15717,N_15754);
or U17487 (N_17487,N_16374,N_15970);
nand U17488 (N_17488,N_16250,N_16315);
or U17489 (N_17489,N_15999,N_16005);
nand U17490 (N_17490,N_16142,N_16609);
nand U17491 (N_17491,N_15606,N_16077);
nor U17492 (N_17492,N_16688,N_15913);
or U17493 (N_17493,N_15847,N_15648);
or U17494 (N_17494,N_15754,N_15761);
nand U17495 (N_17495,N_16264,N_15772);
or U17496 (N_17496,N_15889,N_16188);
nand U17497 (N_17497,N_15709,N_16652);
or U17498 (N_17498,N_16230,N_15612);
or U17499 (N_17499,N_16354,N_15856);
nor U17500 (N_17500,N_16573,N_16174);
and U17501 (N_17501,N_16128,N_16562);
xor U17502 (N_17502,N_15945,N_16515);
xnor U17503 (N_17503,N_15634,N_15854);
xor U17504 (N_17504,N_16502,N_15608);
xor U17505 (N_17505,N_16674,N_16032);
nor U17506 (N_17506,N_16770,N_16632);
or U17507 (N_17507,N_16292,N_16503);
xnor U17508 (N_17508,N_16256,N_15933);
and U17509 (N_17509,N_16248,N_16739);
xnor U17510 (N_17510,N_16437,N_15841);
or U17511 (N_17511,N_16131,N_16565);
xnor U17512 (N_17512,N_16604,N_15771);
xor U17513 (N_17513,N_15777,N_16099);
nor U17514 (N_17514,N_16119,N_16571);
and U17515 (N_17515,N_16546,N_15864);
or U17516 (N_17516,N_16040,N_15703);
nor U17517 (N_17517,N_16178,N_16701);
xnor U17518 (N_17518,N_16365,N_16279);
and U17519 (N_17519,N_15796,N_15840);
or U17520 (N_17520,N_15949,N_15967);
xnor U17521 (N_17521,N_15914,N_16745);
nand U17522 (N_17522,N_16517,N_15726);
nor U17523 (N_17523,N_15817,N_16356);
nand U17524 (N_17524,N_15620,N_16716);
nand U17525 (N_17525,N_16642,N_16459);
nand U17526 (N_17526,N_16200,N_16051);
and U17527 (N_17527,N_16008,N_16326);
nand U17528 (N_17528,N_16745,N_15994);
nand U17529 (N_17529,N_15808,N_16406);
and U17530 (N_17530,N_15639,N_16320);
and U17531 (N_17531,N_16573,N_16144);
nand U17532 (N_17532,N_16176,N_16152);
xor U17533 (N_17533,N_16041,N_15823);
or U17534 (N_17534,N_15905,N_15990);
xnor U17535 (N_17535,N_16685,N_16529);
nand U17536 (N_17536,N_15924,N_16251);
or U17537 (N_17537,N_15949,N_16199);
and U17538 (N_17538,N_15992,N_15849);
xor U17539 (N_17539,N_16360,N_16685);
or U17540 (N_17540,N_15760,N_16551);
nand U17541 (N_17541,N_15759,N_16437);
xor U17542 (N_17542,N_16115,N_16372);
and U17543 (N_17543,N_15835,N_15799);
xnor U17544 (N_17544,N_16081,N_16210);
nand U17545 (N_17545,N_15600,N_16116);
or U17546 (N_17546,N_16137,N_15621);
or U17547 (N_17547,N_16304,N_15925);
nand U17548 (N_17548,N_16178,N_15662);
nand U17549 (N_17549,N_15962,N_16033);
nand U17550 (N_17550,N_16377,N_16109);
and U17551 (N_17551,N_15610,N_16457);
and U17552 (N_17552,N_16495,N_16662);
nor U17553 (N_17553,N_15920,N_15876);
or U17554 (N_17554,N_16468,N_15616);
or U17555 (N_17555,N_16758,N_16757);
and U17556 (N_17556,N_16186,N_16057);
nor U17557 (N_17557,N_15681,N_15946);
nand U17558 (N_17558,N_16334,N_16129);
or U17559 (N_17559,N_15839,N_15713);
xnor U17560 (N_17560,N_15976,N_16534);
nand U17561 (N_17561,N_16399,N_16628);
nand U17562 (N_17562,N_16433,N_16136);
nor U17563 (N_17563,N_15625,N_16194);
and U17564 (N_17564,N_15717,N_15968);
or U17565 (N_17565,N_16214,N_15685);
nand U17566 (N_17566,N_16061,N_15702);
and U17567 (N_17567,N_15928,N_16205);
nand U17568 (N_17568,N_16419,N_16531);
nor U17569 (N_17569,N_15752,N_15829);
nor U17570 (N_17570,N_15806,N_16057);
and U17571 (N_17571,N_15674,N_16767);
and U17572 (N_17572,N_16385,N_15701);
xor U17573 (N_17573,N_16336,N_16599);
xor U17574 (N_17574,N_16527,N_15696);
xnor U17575 (N_17575,N_15767,N_16652);
or U17576 (N_17576,N_16714,N_16479);
xor U17577 (N_17577,N_16078,N_16623);
or U17578 (N_17578,N_15964,N_16381);
xnor U17579 (N_17579,N_15618,N_16194);
or U17580 (N_17580,N_16628,N_16196);
nand U17581 (N_17581,N_16542,N_15824);
and U17582 (N_17582,N_16312,N_16434);
xor U17583 (N_17583,N_16267,N_16012);
xnor U17584 (N_17584,N_15812,N_15642);
nor U17585 (N_17585,N_16649,N_16482);
nand U17586 (N_17586,N_16473,N_15836);
nor U17587 (N_17587,N_15793,N_16581);
and U17588 (N_17588,N_16465,N_16422);
or U17589 (N_17589,N_16243,N_15887);
or U17590 (N_17590,N_16768,N_16195);
xnor U17591 (N_17591,N_16031,N_16671);
nor U17592 (N_17592,N_16359,N_16320);
or U17593 (N_17593,N_16090,N_16019);
or U17594 (N_17594,N_16602,N_15993);
nor U17595 (N_17595,N_15905,N_15902);
nand U17596 (N_17596,N_16280,N_16451);
nor U17597 (N_17597,N_16250,N_15655);
xor U17598 (N_17598,N_16038,N_16727);
nand U17599 (N_17599,N_16278,N_15946);
nand U17600 (N_17600,N_16345,N_16168);
or U17601 (N_17601,N_16596,N_16183);
and U17602 (N_17602,N_16553,N_16615);
xnor U17603 (N_17603,N_16164,N_16146);
and U17604 (N_17604,N_15863,N_16794);
and U17605 (N_17605,N_16025,N_15619);
nand U17606 (N_17606,N_16581,N_16129);
nor U17607 (N_17607,N_16590,N_16427);
and U17608 (N_17608,N_16126,N_16507);
and U17609 (N_17609,N_15676,N_16389);
or U17610 (N_17610,N_15644,N_16358);
nor U17611 (N_17611,N_16143,N_15835);
nor U17612 (N_17612,N_15775,N_16512);
nor U17613 (N_17613,N_16702,N_16014);
xor U17614 (N_17614,N_16693,N_16199);
nor U17615 (N_17615,N_15936,N_16348);
nor U17616 (N_17616,N_16120,N_16350);
nand U17617 (N_17617,N_16732,N_15699);
or U17618 (N_17618,N_15705,N_16511);
and U17619 (N_17619,N_15997,N_16134);
and U17620 (N_17620,N_15966,N_16524);
nor U17621 (N_17621,N_16257,N_16032);
nor U17622 (N_17622,N_16723,N_16196);
nand U17623 (N_17623,N_15859,N_16455);
and U17624 (N_17624,N_16294,N_15895);
and U17625 (N_17625,N_16388,N_16366);
or U17626 (N_17626,N_15856,N_16389);
or U17627 (N_17627,N_16435,N_15822);
xor U17628 (N_17628,N_15970,N_16294);
and U17629 (N_17629,N_15754,N_16777);
or U17630 (N_17630,N_16246,N_16542);
nand U17631 (N_17631,N_16223,N_15806);
and U17632 (N_17632,N_16150,N_16123);
nand U17633 (N_17633,N_16448,N_16554);
xnor U17634 (N_17634,N_16234,N_16303);
nand U17635 (N_17635,N_16687,N_16655);
nand U17636 (N_17636,N_16300,N_16624);
nand U17637 (N_17637,N_15847,N_16293);
or U17638 (N_17638,N_16710,N_15740);
nor U17639 (N_17639,N_16295,N_16271);
and U17640 (N_17640,N_15638,N_16797);
nand U17641 (N_17641,N_16481,N_16265);
or U17642 (N_17642,N_16616,N_16570);
nand U17643 (N_17643,N_15710,N_16334);
or U17644 (N_17644,N_15679,N_16596);
or U17645 (N_17645,N_16501,N_15816);
xnor U17646 (N_17646,N_16230,N_15683);
nor U17647 (N_17647,N_16064,N_15668);
nand U17648 (N_17648,N_15650,N_15902);
and U17649 (N_17649,N_16058,N_15902);
nor U17650 (N_17650,N_16186,N_16219);
nor U17651 (N_17651,N_15899,N_16111);
and U17652 (N_17652,N_16503,N_15857);
xor U17653 (N_17653,N_16156,N_15830);
xor U17654 (N_17654,N_16449,N_16102);
nand U17655 (N_17655,N_16363,N_15853);
or U17656 (N_17656,N_16564,N_16011);
or U17657 (N_17657,N_15894,N_16638);
nand U17658 (N_17658,N_16528,N_16013);
xor U17659 (N_17659,N_16696,N_15820);
or U17660 (N_17660,N_16720,N_15706);
and U17661 (N_17661,N_15705,N_15769);
or U17662 (N_17662,N_15940,N_15659);
or U17663 (N_17663,N_16017,N_16723);
xnor U17664 (N_17664,N_16413,N_16702);
nor U17665 (N_17665,N_16387,N_15939);
xor U17666 (N_17666,N_15905,N_16773);
nor U17667 (N_17667,N_15795,N_16448);
or U17668 (N_17668,N_15974,N_16731);
xor U17669 (N_17669,N_16057,N_16797);
xor U17670 (N_17670,N_16669,N_15846);
and U17671 (N_17671,N_16352,N_15749);
or U17672 (N_17672,N_16060,N_15718);
or U17673 (N_17673,N_16381,N_16211);
or U17674 (N_17674,N_15717,N_16736);
xnor U17675 (N_17675,N_15624,N_15627);
xor U17676 (N_17676,N_16492,N_16036);
xor U17677 (N_17677,N_16166,N_16234);
and U17678 (N_17678,N_16693,N_15818);
nor U17679 (N_17679,N_16728,N_16297);
nand U17680 (N_17680,N_16043,N_15846);
xnor U17681 (N_17681,N_16276,N_16635);
nor U17682 (N_17682,N_15758,N_15756);
xor U17683 (N_17683,N_15774,N_15793);
nor U17684 (N_17684,N_16440,N_15855);
and U17685 (N_17685,N_16095,N_16567);
or U17686 (N_17686,N_16706,N_16695);
or U17687 (N_17687,N_15807,N_15942);
nor U17688 (N_17688,N_16622,N_15726);
nand U17689 (N_17689,N_16508,N_15933);
and U17690 (N_17690,N_15996,N_16373);
and U17691 (N_17691,N_16337,N_16180);
xnor U17692 (N_17692,N_16169,N_15942);
nor U17693 (N_17693,N_16089,N_16541);
and U17694 (N_17694,N_16029,N_16210);
or U17695 (N_17695,N_16112,N_16243);
or U17696 (N_17696,N_15781,N_15863);
or U17697 (N_17697,N_15770,N_15826);
nor U17698 (N_17698,N_16598,N_16765);
and U17699 (N_17699,N_16677,N_16122);
nor U17700 (N_17700,N_16795,N_15678);
nand U17701 (N_17701,N_16726,N_15856);
nand U17702 (N_17702,N_16547,N_16491);
nand U17703 (N_17703,N_15889,N_16263);
xor U17704 (N_17704,N_16007,N_16606);
nor U17705 (N_17705,N_16148,N_16450);
nand U17706 (N_17706,N_16291,N_15784);
nand U17707 (N_17707,N_15944,N_16297);
nand U17708 (N_17708,N_16428,N_16667);
nor U17709 (N_17709,N_15772,N_16565);
nand U17710 (N_17710,N_15669,N_16027);
xor U17711 (N_17711,N_16216,N_15870);
xnor U17712 (N_17712,N_16396,N_16102);
xor U17713 (N_17713,N_15698,N_15773);
xnor U17714 (N_17714,N_16767,N_16410);
and U17715 (N_17715,N_15884,N_15819);
or U17716 (N_17716,N_16479,N_15998);
nand U17717 (N_17717,N_15756,N_16100);
nand U17718 (N_17718,N_16051,N_15702);
xor U17719 (N_17719,N_16509,N_16542);
or U17720 (N_17720,N_16313,N_16355);
nand U17721 (N_17721,N_15629,N_16374);
and U17722 (N_17722,N_16484,N_16034);
or U17723 (N_17723,N_16612,N_16577);
nand U17724 (N_17724,N_15725,N_15604);
nor U17725 (N_17725,N_16148,N_16490);
and U17726 (N_17726,N_16697,N_16245);
nand U17727 (N_17727,N_16594,N_15601);
or U17728 (N_17728,N_15939,N_16007);
nand U17729 (N_17729,N_15868,N_15931);
xnor U17730 (N_17730,N_16654,N_16161);
nand U17731 (N_17731,N_15912,N_16798);
or U17732 (N_17732,N_16703,N_15641);
or U17733 (N_17733,N_16234,N_16666);
and U17734 (N_17734,N_16206,N_16478);
nand U17735 (N_17735,N_16155,N_16670);
and U17736 (N_17736,N_16165,N_16343);
xor U17737 (N_17737,N_16038,N_16270);
or U17738 (N_17738,N_16555,N_16605);
and U17739 (N_17739,N_15678,N_16680);
or U17740 (N_17740,N_15859,N_16022);
nand U17741 (N_17741,N_16738,N_16789);
or U17742 (N_17742,N_16460,N_15624);
or U17743 (N_17743,N_15911,N_16798);
or U17744 (N_17744,N_16272,N_16030);
and U17745 (N_17745,N_15955,N_16500);
xor U17746 (N_17746,N_16093,N_16349);
and U17747 (N_17747,N_15770,N_16579);
xnor U17748 (N_17748,N_15972,N_16526);
and U17749 (N_17749,N_16673,N_15918);
nand U17750 (N_17750,N_15826,N_15724);
nor U17751 (N_17751,N_16593,N_16239);
and U17752 (N_17752,N_15943,N_16758);
or U17753 (N_17753,N_16156,N_16480);
or U17754 (N_17754,N_16185,N_16272);
or U17755 (N_17755,N_16545,N_16017);
or U17756 (N_17756,N_16394,N_16693);
nand U17757 (N_17757,N_15746,N_15692);
xnor U17758 (N_17758,N_16387,N_16458);
or U17759 (N_17759,N_16108,N_16260);
and U17760 (N_17760,N_15931,N_16620);
or U17761 (N_17761,N_16178,N_16385);
nand U17762 (N_17762,N_15971,N_16162);
xnor U17763 (N_17763,N_16101,N_15684);
or U17764 (N_17764,N_16201,N_15945);
nor U17765 (N_17765,N_16562,N_15692);
nand U17766 (N_17766,N_15793,N_16707);
and U17767 (N_17767,N_16408,N_15877);
and U17768 (N_17768,N_15872,N_15783);
nor U17769 (N_17769,N_16110,N_16625);
xor U17770 (N_17770,N_16647,N_16592);
nand U17771 (N_17771,N_16427,N_16776);
nor U17772 (N_17772,N_16454,N_16130);
or U17773 (N_17773,N_15618,N_16670);
nand U17774 (N_17774,N_15783,N_16572);
and U17775 (N_17775,N_16657,N_16101);
or U17776 (N_17776,N_16078,N_16470);
nand U17777 (N_17777,N_15677,N_16797);
nor U17778 (N_17778,N_15630,N_15905);
or U17779 (N_17779,N_15727,N_16523);
nor U17780 (N_17780,N_15936,N_16123);
or U17781 (N_17781,N_16757,N_16418);
xor U17782 (N_17782,N_16279,N_15683);
nor U17783 (N_17783,N_16462,N_16036);
nand U17784 (N_17784,N_16028,N_15646);
xor U17785 (N_17785,N_16141,N_16095);
nor U17786 (N_17786,N_16058,N_16452);
nand U17787 (N_17787,N_16656,N_15687);
and U17788 (N_17788,N_15935,N_16263);
nand U17789 (N_17789,N_15629,N_15663);
and U17790 (N_17790,N_16133,N_16254);
or U17791 (N_17791,N_15929,N_16127);
nand U17792 (N_17792,N_15904,N_15614);
or U17793 (N_17793,N_16310,N_16050);
nor U17794 (N_17794,N_16730,N_16634);
and U17795 (N_17795,N_16233,N_16182);
nor U17796 (N_17796,N_15842,N_15658);
and U17797 (N_17797,N_16264,N_16144);
and U17798 (N_17798,N_15795,N_15747);
xnor U17799 (N_17799,N_16402,N_15630);
and U17800 (N_17800,N_16749,N_16518);
and U17801 (N_17801,N_16124,N_16383);
and U17802 (N_17802,N_16709,N_16656);
xnor U17803 (N_17803,N_16221,N_16084);
nor U17804 (N_17804,N_16463,N_16595);
xnor U17805 (N_17805,N_16753,N_15780);
or U17806 (N_17806,N_15810,N_16779);
nor U17807 (N_17807,N_15966,N_15699);
or U17808 (N_17808,N_16084,N_16737);
or U17809 (N_17809,N_15850,N_16146);
xnor U17810 (N_17810,N_16325,N_16561);
nand U17811 (N_17811,N_15866,N_16112);
nor U17812 (N_17812,N_16001,N_16764);
and U17813 (N_17813,N_16357,N_16294);
or U17814 (N_17814,N_15653,N_16208);
xor U17815 (N_17815,N_16374,N_16715);
and U17816 (N_17816,N_16167,N_16408);
nor U17817 (N_17817,N_16013,N_15747);
xor U17818 (N_17818,N_15605,N_16437);
nand U17819 (N_17819,N_15859,N_16620);
nor U17820 (N_17820,N_16033,N_16345);
nand U17821 (N_17821,N_16743,N_15818);
nor U17822 (N_17822,N_16558,N_16543);
nor U17823 (N_17823,N_15697,N_16300);
and U17824 (N_17824,N_16374,N_16362);
nand U17825 (N_17825,N_16442,N_15867);
xor U17826 (N_17826,N_15652,N_15693);
xor U17827 (N_17827,N_16245,N_16009);
nor U17828 (N_17828,N_15716,N_16752);
nor U17829 (N_17829,N_16317,N_16227);
or U17830 (N_17830,N_16754,N_16302);
nand U17831 (N_17831,N_16224,N_15670);
and U17832 (N_17832,N_16776,N_16642);
and U17833 (N_17833,N_16795,N_15795);
xnor U17834 (N_17834,N_15927,N_15990);
or U17835 (N_17835,N_16064,N_15923);
and U17836 (N_17836,N_16385,N_15640);
or U17837 (N_17837,N_16784,N_16386);
and U17838 (N_17838,N_16528,N_15898);
nor U17839 (N_17839,N_15651,N_15861);
xor U17840 (N_17840,N_16093,N_16139);
xnor U17841 (N_17841,N_16404,N_16057);
and U17842 (N_17842,N_16269,N_16730);
xnor U17843 (N_17843,N_15924,N_15721);
nor U17844 (N_17844,N_15697,N_16347);
and U17845 (N_17845,N_16492,N_15763);
or U17846 (N_17846,N_15640,N_15965);
xor U17847 (N_17847,N_15987,N_16533);
nand U17848 (N_17848,N_15969,N_15756);
and U17849 (N_17849,N_15886,N_16391);
or U17850 (N_17850,N_15988,N_16616);
or U17851 (N_17851,N_16308,N_15957);
xor U17852 (N_17852,N_15635,N_16119);
and U17853 (N_17853,N_15855,N_15677);
xnor U17854 (N_17854,N_16157,N_16187);
nor U17855 (N_17855,N_15768,N_16513);
nor U17856 (N_17856,N_15743,N_16199);
and U17857 (N_17857,N_16224,N_15966);
nor U17858 (N_17858,N_16488,N_16502);
and U17859 (N_17859,N_16240,N_15639);
nor U17860 (N_17860,N_16747,N_15667);
nand U17861 (N_17861,N_15854,N_16033);
nor U17862 (N_17862,N_15661,N_16702);
xnor U17863 (N_17863,N_16496,N_16353);
nor U17864 (N_17864,N_15728,N_15804);
nand U17865 (N_17865,N_16029,N_16170);
or U17866 (N_17866,N_16543,N_15893);
nand U17867 (N_17867,N_16369,N_16307);
nor U17868 (N_17868,N_15897,N_15915);
or U17869 (N_17869,N_16202,N_15760);
and U17870 (N_17870,N_16076,N_15895);
xor U17871 (N_17871,N_16682,N_16763);
nor U17872 (N_17872,N_15871,N_16402);
nand U17873 (N_17873,N_15756,N_16398);
xor U17874 (N_17874,N_16318,N_15795);
nand U17875 (N_17875,N_16231,N_16421);
xnor U17876 (N_17876,N_16492,N_16758);
nand U17877 (N_17877,N_16634,N_15882);
nor U17878 (N_17878,N_16503,N_16016);
and U17879 (N_17879,N_16306,N_15916);
or U17880 (N_17880,N_16768,N_16570);
and U17881 (N_17881,N_16768,N_16313);
xnor U17882 (N_17882,N_16161,N_16391);
nor U17883 (N_17883,N_16554,N_16251);
and U17884 (N_17884,N_16569,N_15739);
nor U17885 (N_17885,N_16689,N_16612);
or U17886 (N_17886,N_16470,N_16644);
nor U17887 (N_17887,N_15907,N_15850);
and U17888 (N_17888,N_15670,N_15804);
and U17889 (N_17889,N_16605,N_16479);
nand U17890 (N_17890,N_16202,N_15874);
xor U17891 (N_17891,N_16408,N_16333);
and U17892 (N_17892,N_16627,N_16202);
xor U17893 (N_17893,N_16772,N_16608);
nand U17894 (N_17894,N_15778,N_16122);
and U17895 (N_17895,N_16268,N_16062);
or U17896 (N_17896,N_16726,N_15941);
or U17897 (N_17897,N_15685,N_16711);
and U17898 (N_17898,N_15965,N_16599);
nand U17899 (N_17899,N_16707,N_16767);
and U17900 (N_17900,N_15640,N_16762);
nand U17901 (N_17901,N_16572,N_16490);
or U17902 (N_17902,N_16016,N_16175);
xor U17903 (N_17903,N_15952,N_16110);
and U17904 (N_17904,N_16757,N_15663);
xor U17905 (N_17905,N_16413,N_16333);
nand U17906 (N_17906,N_16446,N_15719);
nand U17907 (N_17907,N_16733,N_16548);
nor U17908 (N_17908,N_16285,N_15677);
xor U17909 (N_17909,N_15885,N_16652);
nand U17910 (N_17910,N_16226,N_15788);
nand U17911 (N_17911,N_16767,N_16355);
nor U17912 (N_17912,N_16064,N_16327);
nor U17913 (N_17913,N_16521,N_15851);
nor U17914 (N_17914,N_15695,N_16427);
and U17915 (N_17915,N_16129,N_15943);
nor U17916 (N_17916,N_16657,N_16344);
or U17917 (N_17917,N_16452,N_16438);
nor U17918 (N_17918,N_16260,N_16053);
or U17919 (N_17919,N_15728,N_16441);
nor U17920 (N_17920,N_16164,N_16137);
xnor U17921 (N_17921,N_16007,N_16555);
and U17922 (N_17922,N_15687,N_16560);
or U17923 (N_17923,N_16429,N_16217);
nor U17924 (N_17924,N_16469,N_16018);
xor U17925 (N_17925,N_15934,N_16526);
nand U17926 (N_17926,N_16421,N_16100);
or U17927 (N_17927,N_16577,N_15792);
and U17928 (N_17928,N_16796,N_16765);
and U17929 (N_17929,N_15706,N_16223);
xor U17930 (N_17930,N_15961,N_15893);
and U17931 (N_17931,N_16163,N_15613);
nor U17932 (N_17932,N_15605,N_15883);
or U17933 (N_17933,N_16591,N_16786);
nand U17934 (N_17934,N_16553,N_16419);
xnor U17935 (N_17935,N_16207,N_16465);
xnor U17936 (N_17936,N_15707,N_16035);
nand U17937 (N_17937,N_15879,N_16407);
or U17938 (N_17938,N_15676,N_16173);
nor U17939 (N_17939,N_16579,N_16247);
and U17940 (N_17940,N_16051,N_16799);
and U17941 (N_17941,N_16381,N_16556);
nand U17942 (N_17942,N_15855,N_15940);
nor U17943 (N_17943,N_16240,N_15903);
nand U17944 (N_17944,N_16614,N_16294);
and U17945 (N_17945,N_16010,N_15904);
or U17946 (N_17946,N_15821,N_15693);
or U17947 (N_17947,N_15773,N_16507);
or U17948 (N_17948,N_16145,N_15738);
nand U17949 (N_17949,N_16753,N_16117);
nand U17950 (N_17950,N_15676,N_16005);
and U17951 (N_17951,N_15902,N_16094);
and U17952 (N_17952,N_16061,N_16318);
nand U17953 (N_17953,N_16569,N_16731);
xor U17954 (N_17954,N_15830,N_16732);
nor U17955 (N_17955,N_15909,N_16224);
nand U17956 (N_17956,N_16204,N_16686);
xnor U17957 (N_17957,N_16329,N_16260);
nor U17958 (N_17958,N_16623,N_16020);
xor U17959 (N_17959,N_15741,N_15695);
or U17960 (N_17960,N_15710,N_16607);
nand U17961 (N_17961,N_16166,N_16690);
xnor U17962 (N_17962,N_16632,N_15675);
nor U17963 (N_17963,N_16291,N_16564);
or U17964 (N_17964,N_15697,N_15975);
or U17965 (N_17965,N_15856,N_15728);
and U17966 (N_17966,N_15953,N_16303);
and U17967 (N_17967,N_16749,N_15987);
xor U17968 (N_17968,N_16279,N_16067);
and U17969 (N_17969,N_16451,N_15934);
nor U17970 (N_17970,N_16761,N_16031);
nor U17971 (N_17971,N_15996,N_16161);
and U17972 (N_17972,N_16341,N_16307);
and U17973 (N_17973,N_15687,N_16008);
and U17974 (N_17974,N_16360,N_16297);
or U17975 (N_17975,N_16012,N_16505);
nand U17976 (N_17976,N_16110,N_16503);
nor U17977 (N_17977,N_16115,N_16738);
xnor U17978 (N_17978,N_16479,N_16463);
and U17979 (N_17979,N_15789,N_16081);
xnor U17980 (N_17980,N_16195,N_16742);
xnor U17981 (N_17981,N_15650,N_15968);
or U17982 (N_17982,N_16547,N_16508);
xor U17983 (N_17983,N_16191,N_15787);
nand U17984 (N_17984,N_16335,N_16610);
and U17985 (N_17985,N_16383,N_15725);
nor U17986 (N_17986,N_15695,N_16008);
nand U17987 (N_17987,N_16253,N_16075);
xnor U17988 (N_17988,N_15665,N_16577);
and U17989 (N_17989,N_16098,N_15849);
xnor U17990 (N_17990,N_16799,N_16305);
nor U17991 (N_17991,N_16272,N_16349);
or U17992 (N_17992,N_16051,N_16513);
and U17993 (N_17993,N_16200,N_15782);
nor U17994 (N_17994,N_16310,N_16451);
or U17995 (N_17995,N_15859,N_16112);
xor U17996 (N_17996,N_16441,N_16121);
and U17997 (N_17997,N_16356,N_16676);
and U17998 (N_17998,N_16549,N_15717);
and U17999 (N_17999,N_15641,N_16777);
nand U18000 (N_18000,N_16888,N_17038);
and U18001 (N_18001,N_17719,N_17774);
or U18002 (N_18002,N_17622,N_17930);
xor U18003 (N_18003,N_17413,N_17028);
and U18004 (N_18004,N_16825,N_17547);
or U18005 (N_18005,N_17842,N_17192);
or U18006 (N_18006,N_17739,N_17744);
and U18007 (N_18007,N_17761,N_17806);
xnor U18008 (N_18008,N_16981,N_17232);
or U18009 (N_18009,N_17572,N_17974);
nand U18010 (N_18010,N_17627,N_17630);
nor U18011 (N_18011,N_17268,N_17057);
or U18012 (N_18012,N_17474,N_17479);
nor U18013 (N_18013,N_17001,N_17717);
or U18014 (N_18014,N_17395,N_16872);
nor U18015 (N_18015,N_17350,N_17080);
nand U18016 (N_18016,N_17410,N_16869);
xnor U18017 (N_18017,N_16838,N_17998);
nand U18018 (N_18018,N_17514,N_17582);
nor U18019 (N_18019,N_17706,N_17629);
and U18020 (N_18020,N_17989,N_17443);
nor U18021 (N_18021,N_16951,N_17423);
nor U18022 (N_18022,N_17228,N_16864);
nand U18023 (N_18023,N_17578,N_17773);
nor U18024 (N_18024,N_16975,N_17862);
and U18025 (N_18025,N_17369,N_17515);
nand U18026 (N_18026,N_17062,N_17651);
nor U18027 (N_18027,N_16910,N_17921);
nand U18028 (N_18028,N_16844,N_16887);
xnor U18029 (N_18029,N_17598,N_17800);
and U18030 (N_18030,N_17382,N_17991);
xor U18031 (N_18031,N_17576,N_17979);
nor U18032 (N_18032,N_17561,N_17472);
nor U18033 (N_18033,N_17289,N_16821);
xnor U18034 (N_18034,N_17043,N_17143);
and U18035 (N_18035,N_17463,N_17094);
nor U18036 (N_18036,N_17841,N_17705);
nor U18037 (N_18037,N_17840,N_17802);
xor U18038 (N_18038,N_17136,N_17511);
or U18039 (N_18039,N_17411,N_17000);
or U18040 (N_18040,N_17639,N_17073);
or U18041 (N_18041,N_17619,N_17297);
nor U18042 (N_18042,N_17678,N_17643);
nand U18043 (N_18043,N_17755,N_17075);
and U18044 (N_18044,N_17018,N_17559);
nand U18045 (N_18045,N_17091,N_17770);
or U18046 (N_18046,N_16976,N_17121);
nor U18047 (N_18047,N_17550,N_17579);
nor U18048 (N_18048,N_17556,N_16862);
and U18049 (N_18049,N_17432,N_17496);
nand U18050 (N_18050,N_17174,N_17200);
and U18051 (N_18051,N_17026,N_16858);
nand U18052 (N_18052,N_17918,N_17296);
or U18053 (N_18053,N_17263,N_17799);
xor U18054 (N_18054,N_17061,N_17784);
nor U18055 (N_18055,N_16898,N_16851);
or U18056 (N_18056,N_17925,N_17548);
and U18057 (N_18057,N_17653,N_17148);
nand U18058 (N_18058,N_17461,N_17015);
xor U18059 (N_18059,N_16897,N_17007);
nor U18060 (N_18060,N_17664,N_17449);
xor U18061 (N_18061,N_17788,N_17199);
or U18062 (N_18062,N_16867,N_17117);
nand U18063 (N_18063,N_17224,N_16841);
and U18064 (N_18064,N_16824,N_17845);
and U18065 (N_18065,N_17183,N_17795);
nand U18066 (N_18066,N_16892,N_16837);
xor U18067 (N_18067,N_16967,N_16938);
nand U18068 (N_18068,N_17282,N_17586);
xnor U18069 (N_18069,N_17856,N_17066);
nand U18070 (N_18070,N_17944,N_17217);
or U18071 (N_18071,N_17684,N_17415);
nor U18072 (N_18072,N_17114,N_17523);
or U18073 (N_18073,N_17725,N_17190);
nor U18074 (N_18074,N_17687,N_17343);
and U18075 (N_18075,N_16893,N_17754);
nor U18076 (N_18076,N_17670,N_16880);
and U18077 (N_18077,N_17099,N_17155);
nand U18078 (N_18078,N_17288,N_16885);
nand U18079 (N_18079,N_17628,N_17792);
nand U18080 (N_18080,N_16937,N_17607);
or U18081 (N_18081,N_17573,N_17527);
nand U18082 (N_18082,N_17145,N_16912);
or U18083 (N_18083,N_17539,N_17919);
and U18084 (N_18084,N_16947,N_17210);
nor U18085 (N_18085,N_17734,N_16816);
nor U18086 (N_18086,N_17286,N_17872);
and U18087 (N_18087,N_17823,N_17748);
xnor U18088 (N_18088,N_17491,N_17574);
and U18089 (N_18089,N_16996,N_17189);
and U18090 (N_18090,N_17131,N_17654);
nor U18091 (N_18091,N_16907,N_17722);
and U18092 (N_18092,N_17027,N_17635);
and U18093 (N_18093,N_16911,N_17924);
xnor U18094 (N_18094,N_16944,N_17960);
xnor U18095 (N_18095,N_17950,N_17170);
xnor U18096 (N_18096,N_17280,N_17877);
nor U18097 (N_18097,N_17588,N_17609);
or U18098 (N_18098,N_16913,N_17266);
and U18099 (N_18099,N_17728,N_17405);
nand U18100 (N_18100,N_17457,N_17434);
and U18101 (N_18101,N_17851,N_16991);
and U18102 (N_18102,N_17605,N_17377);
xnor U18103 (N_18103,N_17133,N_17655);
or U18104 (N_18104,N_17575,N_16860);
nand U18105 (N_18105,N_17737,N_17911);
nand U18106 (N_18106,N_17243,N_17898);
nand U18107 (N_18107,N_17513,N_17384);
xnor U18108 (N_18108,N_17260,N_17420);
xnor U18109 (N_18109,N_17969,N_16823);
and U18110 (N_18110,N_17928,N_17392);
and U18111 (N_18111,N_17486,N_17585);
or U18112 (N_18112,N_17014,N_17315);
xnor U18113 (N_18113,N_17682,N_16906);
xor U18114 (N_18114,N_16828,N_17180);
xor U18115 (N_18115,N_17864,N_16903);
nand U18116 (N_18116,N_17068,N_17339);
nand U18117 (N_18117,N_17204,N_17901);
nor U18118 (N_18118,N_17334,N_16997);
nand U18119 (N_18119,N_17163,N_17187);
or U18120 (N_18120,N_17487,N_17086);
or U18121 (N_18121,N_17084,N_17345);
nor U18122 (N_18122,N_17389,N_17050);
nor U18123 (N_18123,N_17211,N_17107);
and U18124 (N_18124,N_16900,N_17031);
nor U18125 (N_18125,N_17674,N_17450);
nand U18126 (N_18126,N_16980,N_17064);
xor U18127 (N_18127,N_16982,N_16859);
xor U18128 (N_18128,N_17939,N_17876);
nor U18129 (N_18129,N_17226,N_17947);
xor U18130 (N_18130,N_16843,N_16891);
nor U18131 (N_18131,N_16852,N_16865);
and U18132 (N_18132,N_17025,N_17277);
or U18133 (N_18133,N_16985,N_17081);
nand U18134 (N_18134,N_16835,N_17763);
nor U18135 (N_18135,N_17894,N_17490);
or U18136 (N_18136,N_17853,N_17600);
nor U18137 (N_18137,N_16886,N_17879);
xnor U18138 (N_18138,N_17510,N_17890);
nor U18139 (N_18139,N_17326,N_17359);
nor U18140 (N_18140,N_17839,N_17525);
or U18141 (N_18141,N_17042,N_17690);
and U18142 (N_18142,N_17887,N_17594);
nand U18143 (N_18143,N_17358,N_17022);
xnor U18144 (N_18144,N_17857,N_17252);
nor U18145 (N_18145,N_17045,N_17290);
nor U18146 (N_18146,N_16806,N_17441);
and U18147 (N_18147,N_17077,N_17203);
nor U18148 (N_18148,N_17135,N_17591);
nand U18149 (N_18149,N_17716,N_16882);
or U18150 (N_18150,N_17004,N_17162);
nor U18151 (N_18151,N_17568,N_16979);
or U18152 (N_18152,N_17023,N_17518);
or U18153 (N_18153,N_16876,N_16977);
nor U18154 (N_18154,N_17319,N_17381);
or U18155 (N_18155,N_17040,N_17172);
xor U18156 (N_18156,N_17418,N_16936);
nand U18157 (N_18157,N_17942,N_17938);
and U18158 (N_18158,N_17868,N_17348);
and U18159 (N_18159,N_17151,N_17880);
nand U18160 (N_18160,N_17673,N_16855);
and U18161 (N_18161,N_16942,N_17460);
nor U18162 (N_18162,N_17936,N_17652);
and U18163 (N_18163,N_16846,N_17354);
and U18164 (N_18164,N_17669,N_17355);
nand U18165 (N_18165,N_17372,N_16874);
and U18166 (N_18166,N_17079,N_17320);
xor U18167 (N_18167,N_17909,N_17067);
nor U18168 (N_18168,N_17738,N_17765);
nand U18169 (N_18169,N_17408,N_17910);
and U18170 (N_18170,N_17499,N_17127);
nand U18171 (N_18171,N_17956,N_16870);
or U18172 (N_18172,N_17419,N_17492);
and U18173 (N_18173,N_17191,N_17948);
or U18174 (N_18174,N_17255,N_17834);
and U18175 (N_18175,N_17325,N_17269);
or U18176 (N_18176,N_17656,N_17299);
xor U18177 (N_18177,N_17003,N_16971);
or U18178 (N_18178,N_17584,N_17915);
nor U18179 (N_18179,N_17169,N_16905);
and U18180 (N_18180,N_17336,N_17214);
nand U18181 (N_18181,N_17536,N_16963);
nand U18182 (N_18182,N_17822,N_17638);
and U18183 (N_18183,N_16930,N_17794);
nor U18184 (N_18184,N_17284,N_17665);
nor U18185 (N_18185,N_17850,N_17399);
and U18186 (N_18186,N_17453,N_17797);
or U18187 (N_18187,N_17751,N_16948);
or U18188 (N_18188,N_17830,N_17459);
xor U18189 (N_18189,N_17954,N_17274);
nor U18190 (N_18190,N_17955,N_17153);
nand U18191 (N_18191,N_17837,N_17863);
or U18192 (N_18192,N_17386,N_17436);
and U18193 (N_18193,N_17526,N_17060);
xor U18194 (N_18194,N_17475,N_17704);
nor U18195 (N_18195,N_17708,N_17707);
and U18196 (N_18196,N_17537,N_17686);
and U18197 (N_18197,N_17509,N_17963);
and U18198 (N_18198,N_17668,N_17304);
nor U18199 (N_18199,N_17197,N_16969);
or U18200 (N_18200,N_17235,N_17287);
and U18201 (N_18201,N_17820,N_17446);
or U18202 (N_18202,N_17959,N_17016);
and U18203 (N_18203,N_17156,N_17893);
nand U18204 (N_18204,N_17616,N_17636);
or U18205 (N_18205,N_17886,N_17604);
or U18206 (N_18206,N_17109,N_16994);
nand U18207 (N_18207,N_17730,N_17128);
and U18208 (N_18208,N_17516,N_17481);
nand U18209 (N_18209,N_17082,N_17660);
xnor U18210 (N_18210,N_17647,N_17519);
xor U18211 (N_18211,N_17165,N_17309);
nor U18212 (N_18212,N_17878,N_17614);
and U18213 (N_18213,N_17048,N_17058);
nand U18214 (N_18214,N_17859,N_16932);
or U18215 (N_18215,N_17056,N_16809);
and U18216 (N_18216,N_17120,N_17785);
nor U18217 (N_18217,N_17882,N_17379);
nand U18218 (N_18218,N_17819,N_16978);
or U18219 (N_18219,N_17118,N_17809);
or U18220 (N_18220,N_17789,N_17714);
and U18221 (N_18221,N_17726,N_17929);
nand U18222 (N_18222,N_17270,N_17502);
nor U18223 (N_18223,N_16939,N_17821);
nand U18224 (N_18224,N_17544,N_16956);
xnor U18225 (N_18225,N_17231,N_17914);
nand U18226 (N_18226,N_17373,N_16877);
nand U18227 (N_18227,N_17313,N_17658);
xor U18228 (N_18228,N_17769,N_16941);
xnor U18229 (N_18229,N_17213,N_17941);
or U18230 (N_18230,N_17733,N_17138);
and U18231 (N_18231,N_17494,N_17293);
or U18232 (N_18232,N_17597,N_17972);
nor U18233 (N_18233,N_17601,N_16878);
nor U18234 (N_18234,N_16883,N_17371);
nor U18235 (N_18235,N_17321,N_17039);
xor U18236 (N_18236,N_16839,N_17438);
nor U18237 (N_18237,N_17602,N_17680);
nand U18238 (N_18238,N_17508,N_17827);
or U18239 (N_18239,N_16868,N_17676);
xor U18240 (N_18240,N_17988,N_17689);
or U18241 (N_18241,N_17896,N_17913);
nand U18242 (N_18242,N_17849,N_17796);
nand U18243 (N_18243,N_17141,N_17916);
xnor U18244 (N_18244,N_17347,N_17986);
or U18245 (N_18245,N_17428,N_17873);
nor U18246 (N_18246,N_17565,N_17551);
nand U18247 (N_18247,N_16952,N_17444);
nand U18248 (N_18248,N_16989,N_17803);
nor U18249 (N_18249,N_17606,N_17216);
or U18250 (N_18250,N_17100,N_17292);
nor U18251 (N_18251,N_17393,N_17414);
nor U18252 (N_18252,N_17521,N_16802);
xor U18253 (N_18253,N_17926,N_17417);
and U18254 (N_18254,N_17810,N_17677);
and U18255 (N_18255,N_17771,N_17246);
nand U18256 (N_18256,N_17051,N_17152);
nor U18257 (N_18257,N_16814,N_17430);
and U18258 (N_18258,N_17363,N_16803);
or U18259 (N_18259,N_17889,N_17171);
nand U18260 (N_18260,N_17957,N_17173);
nor U18261 (N_18261,N_17892,N_17949);
nor U18262 (N_18262,N_17179,N_16848);
xor U18263 (N_18263,N_17225,N_17498);
nor U18264 (N_18264,N_17462,N_17365);
or U18265 (N_18265,N_17425,N_17899);
xor U18266 (N_18266,N_17698,N_17778);
nor U18267 (N_18267,N_16922,N_17710);
xnor U18268 (N_18268,N_16861,N_17495);
and U18269 (N_18269,N_17049,N_17768);
nand U18270 (N_18270,N_17257,N_16958);
nand U18271 (N_18271,N_17092,N_17251);
and U18272 (N_18272,N_16972,N_17541);
or U18273 (N_18273,N_16854,N_17168);
nand U18274 (N_18274,N_17520,N_17227);
nand U18275 (N_18275,N_17661,N_17825);
xnor U18276 (N_18276,N_17599,N_17375);
and U18277 (N_18277,N_16856,N_17999);
nand U18278 (N_18278,N_17908,N_17147);
xnor U18279 (N_18279,N_17037,N_17471);
xnor U18280 (N_18280,N_17781,N_17455);
and U18281 (N_18281,N_17531,N_17241);
nor U18282 (N_18282,N_17254,N_17249);
nor U18283 (N_18283,N_16889,N_17020);
xor U18284 (N_18284,N_16933,N_16801);
or U18285 (N_18285,N_16826,N_17570);
or U18286 (N_18286,N_17965,N_17528);
nor U18287 (N_18287,N_16987,N_17694);
xor U18288 (N_18288,N_17757,N_16850);
nor U18289 (N_18289,N_17433,N_17401);
xor U18290 (N_18290,N_17826,N_17223);
nand U18291 (N_18291,N_17218,N_17154);
and U18292 (N_18292,N_17236,N_17104);
nand U18293 (N_18293,N_16822,N_17110);
or U18294 (N_18294,N_17976,N_17620);
or U18295 (N_18295,N_17946,N_17995);
nand U18296 (N_18296,N_17558,N_17448);
xnor U18297 (N_18297,N_17657,N_17340);
or U18298 (N_18298,N_16902,N_17804);
and U18299 (N_18299,N_17116,N_17967);
or U18300 (N_18300,N_17701,N_17997);
nor U18301 (N_18301,N_17435,N_17283);
nor U18302 (N_18302,N_17904,N_17012);
xor U18303 (N_18303,N_17964,N_17076);
and U18304 (N_18304,N_16984,N_17762);
and U18305 (N_18305,N_17977,N_16817);
nand U18306 (N_18306,N_17119,N_17580);
and U18307 (N_18307,N_17202,N_17406);
xor U18308 (N_18308,N_16995,N_16908);
nor U18309 (N_18309,N_17617,N_17356);
nor U18310 (N_18310,N_17344,N_17747);
nor U18311 (N_18311,N_17779,N_17517);
nand U18312 (N_18312,N_17087,N_17613);
nand U18313 (N_18313,N_16950,N_17063);
xnor U18314 (N_18314,N_16921,N_17807);
or U18315 (N_18315,N_17990,N_16840);
and U18316 (N_18316,N_17564,N_17302);
and U18317 (N_18317,N_17146,N_17727);
and U18318 (N_18318,N_17212,N_16901);
nor U18319 (N_18319,N_17533,N_17782);
xor U18320 (N_18320,N_17920,N_17250);
nor U18321 (N_18321,N_17306,N_17846);
nor U18322 (N_18322,N_16815,N_17718);
and U18323 (N_18323,N_17703,N_17166);
nand U18324 (N_18324,N_17829,N_17805);
nand U18325 (N_18325,N_17019,N_17412);
nand U18326 (N_18326,N_17456,N_17029);
nor U18327 (N_18327,N_17149,N_16863);
and U18328 (N_18328,N_17832,N_16896);
or U18329 (N_18329,N_17278,N_17464);
or U18330 (N_18330,N_16879,N_17905);
and U18331 (N_18331,N_17489,N_17069);
xnor U18332 (N_18332,N_17175,N_17096);
xor U18333 (N_18333,N_17342,N_17370);
or U18334 (N_18334,N_16909,N_16820);
or U18335 (N_18335,N_17385,N_17507);
nand U18336 (N_18336,N_17993,N_16800);
xor U18337 (N_18337,N_17105,N_17875);
nand U18338 (N_18338,N_16915,N_17641);
and U18339 (N_18339,N_17072,N_17229);
nand U18340 (N_18340,N_17966,N_17318);
or U18341 (N_18341,N_17261,N_17011);
or U18342 (N_18342,N_16924,N_17996);
nor U18343 (N_18343,N_16949,N_16928);
nor U18344 (N_18344,N_17383,N_17137);
and U18345 (N_18345,N_17695,N_17186);
or U18346 (N_18346,N_17663,N_17407);
nor U18347 (N_18347,N_17222,N_17101);
or U18348 (N_18348,N_17790,N_16849);
xnor U18349 (N_18349,N_17477,N_17161);
nor U18350 (N_18350,N_17157,N_17767);
and U18351 (N_18351,N_17934,N_16904);
and U18352 (N_18352,N_16954,N_17812);
xor U18353 (N_18353,N_17248,N_17308);
and U18354 (N_18354,N_17017,N_17331);
nand U18355 (N_18355,N_16934,N_17953);
nor U18356 (N_18356,N_16973,N_16943);
and U18357 (N_18357,N_17828,N_17182);
nor U18358 (N_18358,N_17852,N_17555);
nand U18359 (N_18359,N_17300,N_17088);
xor U18360 (N_18360,N_17699,N_17562);
nand U18361 (N_18361,N_16804,N_16847);
and U18362 (N_18362,N_17264,N_17712);
and U18363 (N_18363,N_17860,N_17397);
or U18364 (N_18364,N_17485,N_17815);
or U18365 (N_18365,N_17237,N_17888);
or U18366 (N_18366,N_17696,N_17743);
nand U18367 (N_18367,N_16813,N_17824);
and U18368 (N_18368,N_17760,N_17335);
xor U18369 (N_18369,N_16884,N_17279);
xor U18370 (N_18370,N_17612,N_17380);
xnor U18371 (N_18371,N_17298,N_17766);
nand U18372 (N_18372,N_17621,N_17317);
xor U18373 (N_18373,N_16988,N_17566);
nand U18374 (N_18374,N_17046,N_17535);
or U18375 (N_18375,N_17409,N_17675);
nor U18376 (N_18376,N_17758,N_17814);
nor U18377 (N_18377,N_17451,N_17590);
nand U18378 (N_18378,N_17097,N_16992);
and U18379 (N_18379,N_17623,N_17650);
xnor U18380 (N_18380,N_17745,N_17740);
or U18381 (N_18381,N_17843,N_16881);
and U18382 (N_18382,N_16986,N_17980);
xor U18383 (N_18383,N_17587,N_17333);
xor U18384 (N_18384,N_17595,N_16831);
and U18385 (N_18385,N_16965,N_17233);
xnor U18386 (N_18386,N_17847,N_17030);
and U18387 (N_18387,N_17106,N_17330);
or U18388 (N_18388,N_17741,N_17102);
and U18389 (N_18389,N_16918,N_17078);
or U18390 (N_18390,N_17242,N_17265);
nor U18391 (N_18391,N_17497,N_17140);
nand U18392 (N_18392,N_17569,N_17387);
xor U18393 (N_18393,N_17129,N_17258);
and U18394 (N_18394,N_17624,N_17891);
or U18395 (N_18395,N_17488,N_17362);
xnor U18396 (N_18396,N_17071,N_17070);
or U18397 (N_18397,N_17835,N_17534);
nand U18398 (N_18398,N_17985,N_17390);
nor U18399 (N_18399,N_17530,N_17962);
nand U18400 (N_18400,N_17906,N_16953);
and U18401 (N_18401,N_16836,N_17922);
or U18402 (N_18402,N_17374,N_17262);
nor U18403 (N_18403,N_17524,N_17281);
and U18404 (N_18404,N_17500,N_17367);
and U18405 (N_18405,N_17732,N_17112);
and U18406 (N_18406,N_17178,N_17752);
nand U18407 (N_18407,N_17307,N_16830);
xor U18408 (N_18408,N_17338,N_17775);
nand U18409 (N_18409,N_17798,N_17167);
nand U18410 (N_18410,N_16926,N_17713);
nor U18411 (N_18411,N_17787,N_17400);
nand U18412 (N_18412,N_17403,N_17632);
or U18413 (N_18413,N_17777,N_17780);
or U18414 (N_18414,N_17074,N_17501);
nand U18415 (N_18415,N_16970,N_17396);
nand U18416 (N_18416,N_16842,N_17378);
or U18417 (N_18417,N_16871,N_17431);
xnor U18418 (N_18418,N_17329,N_17505);
xor U18419 (N_18419,N_17831,N_17059);
or U18420 (N_18420,N_17240,N_17907);
nor U18421 (N_18421,N_17388,N_16957);
xor U18422 (N_18422,N_17208,N_16811);
or U18423 (N_18423,N_17855,N_17791);
nor U18424 (N_18424,N_17253,N_17113);
or U18425 (N_18425,N_16818,N_17724);
nor U18426 (N_18426,N_17865,N_16974);
and U18427 (N_18427,N_17337,N_17238);
nor U18428 (N_18428,N_17546,N_17454);
and U18429 (N_18429,N_17368,N_17532);
and U18430 (N_18430,N_17793,N_17881);
and U18431 (N_18431,N_17275,N_17560);
and U18432 (N_18432,N_17637,N_16945);
nand U18433 (N_18433,N_17567,N_17736);
nor U18434 (N_18434,N_17422,N_17391);
nor U18435 (N_18435,N_16827,N_17111);
nand U18436 (N_18436,N_17185,N_17421);
xor U18437 (N_18437,N_17452,N_16916);
nand U18438 (N_18438,N_17981,N_17646);
nor U18439 (N_18439,N_17122,N_16955);
nand U18440 (N_18440,N_17642,N_17349);
or U18441 (N_18441,N_16917,N_17543);
nand U18442 (N_18442,N_17476,N_17036);
and U18443 (N_18443,N_17177,N_17054);
or U18444 (N_18444,N_17327,N_17158);
nor U18445 (N_18445,N_17596,N_17858);
xor U18446 (N_18446,N_17437,N_17808);
or U18447 (N_18447,N_17010,N_17310);
or U18448 (N_18448,N_17903,N_17429);
nand U18449 (N_18449,N_17402,N_17583);
nand U18450 (N_18450,N_17522,N_17756);
nor U18451 (N_18451,N_17215,N_16873);
nand U18452 (N_18452,N_17644,N_17968);
or U18453 (N_18453,N_17376,N_17483);
and U18454 (N_18454,N_17303,N_16993);
nor U18455 (N_18455,N_17816,N_17357);
and U18456 (N_18456,N_17470,N_17659);
and U18457 (N_18457,N_17353,N_17323);
nor U18458 (N_18458,N_17746,N_17783);
or U18459 (N_18459,N_17818,N_17512);
nand U18460 (N_18460,N_17801,N_17468);
xnor U18461 (N_18461,N_17244,N_17176);
xor U18462 (N_18462,N_17683,N_17398);
xor U18463 (N_18463,N_17667,N_16819);
nand U18464 (N_18464,N_17144,N_17720);
or U18465 (N_18465,N_17052,N_17259);
or U18466 (N_18466,N_17473,N_16894);
and U18467 (N_18467,N_17749,N_17553);
and U18468 (N_18468,N_17447,N_17314);
and U18469 (N_18469,N_17867,N_17721);
nor U18470 (N_18470,N_17671,N_17552);
or U18471 (N_18471,N_17978,N_17529);
or U18472 (N_18472,N_17610,N_16832);
or U18473 (N_18473,N_17294,N_17184);
or U18474 (N_18474,N_17503,N_17723);
or U18475 (N_18475,N_17142,N_17123);
and U18476 (N_18476,N_17902,N_17776);
or U18477 (N_18477,N_17927,N_17895);
nand U18478 (N_18478,N_16935,N_17478);
xor U18479 (N_18479,N_17193,N_17332);
or U18480 (N_18480,N_17709,N_16845);
xor U18481 (N_18481,N_17188,N_17394);
or U18482 (N_18482,N_17442,N_17130);
or U18483 (N_18483,N_17571,N_16983);
and U18484 (N_18484,N_17230,N_17742);
nor U18485 (N_18485,N_17885,N_17871);
nand U18486 (N_18486,N_17764,N_17083);
or U18487 (N_18487,N_17034,N_17631);
and U18488 (N_18488,N_17933,N_17093);
xor U18489 (N_18489,N_17685,N_17198);
and U18490 (N_18490,N_16920,N_17589);
or U18491 (N_18491,N_17861,N_17341);
xor U18492 (N_18492,N_16990,N_17611);
or U18493 (N_18493,N_16866,N_17206);
and U18494 (N_18494,N_17813,N_17540);
nand U18495 (N_18495,N_17205,N_17817);
and U18496 (N_18496,N_17945,N_16962);
xor U18497 (N_18497,N_17917,N_17065);
and U18498 (N_18498,N_17970,N_17884);
and U18499 (N_18499,N_17465,N_16959);
nand U18500 (N_18500,N_17932,N_17440);
or U18501 (N_18501,N_17869,N_17328);
and U18502 (N_18502,N_17150,N_17874);
nor U18503 (N_18503,N_17711,N_17366);
or U18504 (N_18504,N_17691,N_17006);
nand U18505 (N_18505,N_17458,N_17833);
and U18506 (N_18506,N_17542,N_17615);
and U18507 (N_18507,N_17469,N_17008);
nand U18508 (N_18508,N_17681,N_17692);
nand U18509 (N_18509,N_16964,N_17134);
or U18510 (N_18510,N_17992,N_17032);
xor U18511 (N_18511,N_17900,N_17445);
or U18512 (N_18512,N_17424,N_17272);
nor U18513 (N_18513,N_17159,N_17245);
nand U18514 (N_18514,N_17750,N_17640);
or U18515 (N_18515,N_16966,N_17592);
or U18516 (N_18516,N_17923,N_16999);
xor U18517 (N_18517,N_17098,N_17352);
nor U18518 (N_18518,N_17951,N_17480);
or U18519 (N_18519,N_16805,N_17089);
nand U18520 (N_18520,N_17194,N_17618);
and U18521 (N_18521,N_17554,N_17854);
or U18522 (N_18522,N_16829,N_17633);
or U18523 (N_18523,N_17033,N_16925);
nor U18524 (N_18524,N_17164,N_17625);
or U18525 (N_18525,N_17697,N_17053);
nor U18526 (N_18526,N_17883,N_17729);
and U18527 (N_18527,N_17772,N_16853);
nor U18528 (N_18528,N_17731,N_17009);
and U18529 (N_18529,N_17125,N_17952);
nand U18530 (N_18530,N_17645,N_16895);
or U18531 (N_18531,N_17426,N_17961);
or U18532 (N_18532,N_17276,N_17838);
or U18533 (N_18533,N_17973,N_17931);
nand U18534 (N_18534,N_16931,N_17295);
and U18535 (N_18535,N_17538,N_17549);
and U18536 (N_18536,N_17958,N_16998);
xor U18537 (N_18537,N_17836,N_17866);
and U18538 (N_18538,N_17201,N_17291);
xnor U18539 (N_18539,N_17940,N_16808);
xnor U18540 (N_18540,N_17975,N_17221);
xnor U18541 (N_18541,N_17439,N_17811);
xor U18542 (N_18542,N_17364,N_17024);
or U18543 (N_18543,N_17124,N_17679);
or U18544 (N_18544,N_17239,N_17090);
or U18545 (N_18545,N_17844,N_17672);
and U18546 (N_18546,N_16919,N_17181);
or U18547 (N_18547,N_16812,N_17666);
nand U18548 (N_18548,N_16890,N_17360);
nand U18549 (N_18549,N_17634,N_16875);
nor U18550 (N_18550,N_17506,N_17195);
or U18551 (N_18551,N_17700,N_16927);
or U18552 (N_18552,N_17047,N_17311);
nand U18553 (N_18553,N_17688,N_17603);
or U18554 (N_18554,N_17346,N_17115);
or U18555 (N_18555,N_16968,N_17753);
xnor U18556 (N_18556,N_17139,N_17103);
nand U18557 (N_18557,N_17005,N_17937);
xor U18558 (N_18558,N_16946,N_17504);
xor U18559 (N_18559,N_17013,N_17002);
nor U18560 (N_18560,N_16810,N_16960);
and U18561 (N_18561,N_17220,N_17095);
nand U18562 (N_18562,N_16834,N_17870);
and U18563 (N_18563,N_17316,N_17427);
nor U18564 (N_18564,N_17467,N_17035);
nor U18565 (N_18565,N_17648,N_17735);
and U18566 (N_18566,N_17563,N_17557);
or U18567 (N_18567,N_17484,N_17983);
nand U18568 (N_18568,N_17935,N_17271);
or U18569 (N_18569,N_17108,N_17715);
nor U18570 (N_18570,N_17085,N_17219);
xnor U18571 (N_18571,N_16899,N_17247);
xnor U18572 (N_18572,N_17987,N_17943);
xor U18573 (N_18573,N_17234,N_17285);
xnor U18574 (N_18574,N_17693,N_17466);
nor U18575 (N_18575,N_17196,N_17305);
xor U18576 (N_18576,N_17351,N_17055);
and U18577 (N_18577,N_17702,N_17577);
nor U18578 (N_18578,N_17848,N_17482);
and U18579 (N_18579,N_17312,N_16929);
nand U18580 (N_18580,N_17132,N_17044);
nand U18581 (N_18581,N_17759,N_17273);
nor U18582 (N_18582,N_17361,N_17662);
xnor U18583 (N_18583,N_16833,N_17971);
and U18584 (N_18584,N_17994,N_17404);
nor U18585 (N_18585,N_17256,N_17493);
and U18586 (N_18586,N_17416,N_17301);
nand U18587 (N_18587,N_17126,N_17207);
nor U18588 (N_18588,N_16807,N_17021);
nor U18589 (N_18589,N_17322,N_17608);
nor U18590 (N_18590,N_17581,N_17649);
or U18591 (N_18591,N_17160,N_17209);
and U18592 (N_18592,N_17912,N_16857);
xnor U18593 (N_18593,N_17897,N_17324);
nor U18594 (N_18594,N_17982,N_17626);
nand U18595 (N_18595,N_17593,N_17545);
nor U18596 (N_18596,N_16914,N_16940);
xor U18597 (N_18597,N_16961,N_16923);
xnor U18598 (N_18598,N_17984,N_17267);
xor U18599 (N_18599,N_17041,N_17786);
or U18600 (N_18600,N_17445,N_17933);
or U18601 (N_18601,N_17640,N_17070);
and U18602 (N_18602,N_17436,N_17495);
or U18603 (N_18603,N_17938,N_17519);
nand U18604 (N_18604,N_17320,N_17653);
and U18605 (N_18605,N_16961,N_17106);
and U18606 (N_18606,N_17457,N_16956);
nand U18607 (N_18607,N_17055,N_17023);
xnor U18608 (N_18608,N_17430,N_16824);
and U18609 (N_18609,N_16929,N_17974);
and U18610 (N_18610,N_17124,N_17104);
nand U18611 (N_18611,N_16851,N_17479);
xnor U18612 (N_18612,N_17668,N_17787);
and U18613 (N_18613,N_17266,N_17240);
nor U18614 (N_18614,N_17081,N_17247);
nor U18615 (N_18615,N_17718,N_17308);
and U18616 (N_18616,N_17732,N_17669);
nand U18617 (N_18617,N_17099,N_17996);
nand U18618 (N_18618,N_17854,N_17396);
xor U18619 (N_18619,N_16898,N_17097);
nor U18620 (N_18620,N_17877,N_17948);
xnor U18621 (N_18621,N_17088,N_17081);
xor U18622 (N_18622,N_17173,N_17606);
nor U18623 (N_18623,N_17631,N_17980);
and U18624 (N_18624,N_17695,N_17816);
nor U18625 (N_18625,N_17677,N_17179);
and U18626 (N_18626,N_17551,N_17239);
or U18627 (N_18627,N_17782,N_17382);
nor U18628 (N_18628,N_17104,N_17213);
nand U18629 (N_18629,N_17801,N_17826);
and U18630 (N_18630,N_17966,N_17920);
xnor U18631 (N_18631,N_17918,N_17015);
nand U18632 (N_18632,N_17631,N_17102);
and U18633 (N_18633,N_17466,N_17907);
xnor U18634 (N_18634,N_17936,N_17168);
and U18635 (N_18635,N_17064,N_17685);
or U18636 (N_18636,N_17356,N_17412);
and U18637 (N_18637,N_17821,N_16910);
nor U18638 (N_18638,N_17646,N_17935);
nor U18639 (N_18639,N_16862,N_17164);
and U18640 (N_18640,N_17133,N_17187);
xnor U18641 (N_18641,N_17727,N_16963);
xnor U18642 (N_18642,N_17273,N_17258);
xor U18643 (N_18643,N_17041,N_17080);
nand U18644 (N_18644,N_17493,N_16933);
nand U18645 (N_18645,N_17786,N_17345);
nor U18646 (N_18646,N_17768,N_17682);
nor U18647 (N_18647,N_17977,N_17855);
nand U18648 (N_18648,N_16938,N_16884);
nor U18649 (N_18649,N_16948,N_16994);
nor U18650 (N_18650,N_17954,N_17928);
xor U18651 (N_18651,N_17135,N_17373);
and U18652 (N_18652,N_17192,N_17996);
xor U18653 (N_18653,N_16927,N_17827);
xor U18654 (N_18654,N_17451,N_17243);
xor U18655 (N_18655,N_17248,N_17875);
or U18656 (N_18656,N_17197,N_17386);
xor U18657 (N_18657,N_16989,N_17481);
and U18658 (N_18658,N_17418,N_17404);
xnor U18659 (N_18659,N_17997,N_17915);
xnor U18660 (N_18660,N_17900,N_17751);
or U18661 (N_18661,N_16822,N_17461);
xor U18662 (N_18662,N_17634,N_17202);
nand U18663 (N_18663,N_16886,N_17333);
and U18664 (N_18664,N_17201,N_17341);
xnor U18665 (N_18665,N_17954,N_16910);
nor U18666 (N_18666,N_17021,N_16801);
nand U18667 (N_18667,N_17583,N_17085);
and U18668 (N_18668,N_17297,N_17505);
and U18669 (N_18669,N_17918,N_17268);
or U18670 (N_18670,N_17445,N_17607);
or U18671 (N_18671,N_16973,N_17706);
nor U18672 (N_18672,N_17142,N_16889);
nand U18673 (N_18673,N_17510,N_17417);
nand U18674 (N_18674,N_17658,N_16971);
nor U18675 (N_18675,N_17658,N_17470);
nor U18676 (N_18676,N_17185,N_17614);
xor U18677 (N_18677,N_17898,N_17371);
xor U18678 (N_18678,N_16951,N_17388);
or U18679 (N_18679,N_17157,N_17515);
and U18680 (N_18680,N_17421,N_17708);
or U18681 (N_18681,N_17369,N_17248);
and U18682 (N_18682,N_17057,N_17998);
and U18683 (N_18683,N_17953,N_17941);
xor U18684 (N_18684,N_17908,N_17295);
and U18685 (N_18685,N_17691,N_17655);
and U18686 (N_18686,N_16907,N_17573);
nand U18687 (N_18687,N_17440,N_17765);
and U18688 (N_18688,N_17504,N_17529);
nor U18689 (N_18689,N_16943,N_17397);
and U18690 (N_18690,N_17755,N_17114);
xor U18691 (N_18691,N_16972,N_17323);
and U18692 (N_18692,N_17171,N_17074);
nand U18693 (N_18693,N_17312,N_17692);
and U18694 (N_18694,N_17117,N_17411);
nand U18695 (N_18695,N_16954,N_17169);
nand U18696 (N_18696,N_17353,N_17677);
or U18697 (N_18697,N_17654,N_16853);
or U18698 (N_18698,N_17871,N_17977);
and U18699 (N_18699,N_17311,N_17739);
and U18700 (N_18700,N_16991,N_17524);
xnor U18701 (N_18701,N_16973,N_17157);
or U18702 (N_18702,N_17169,N_17954);
nand U18703 (N_18703,N_17594,N_17340);
xor U18704 (N_18704,N_17222,N_17772);
or U18705 (N_18705,N_16949,N_17845);
or U18706 (N_18706,N_17275,N_17110);
xnor U18707 (N_18707,N_17145,N_17141);
nor U18708 (N_18708,N_17141,N_17122);
nand U18709 (N_18709,N_16802,N_17328);
nor U18710 (N_18710,N_17448,N_17642);
xor U18711 (N_18711,N_17049,N_17749);
nand U18712 (N_18712,N_17000,N_17226);
xnor U18713 (N_18713,N_17251,N_16868);
nor U18714 (N_18714,N_17322,N_17357);
and U18715 (N_18715,N_17221,N_17315);
nand U18716 (N_18716,N_17112,N_17345);
nor U18717 (N_18717,N_17902,N_17725);
nand U18718 (N_18718,N_17536,N_16919);
nor U18719 (N_18719,N_17471,N_17652);
nand U18720 (N_18720,N_17534,N_17556);
and U18721 (N_18721,N_17788,N_16869);
or U18722 (N_18722,N_17573,N_17330);
and U18723 (N_18723,N_17889,N_17465);
or U18724 (N_18724,N_17161,N_17893);
nor U18725 (N_18725,N_17860,N_16921);
or U18726 (N_18726,N_17258,N_17661);
nand U18727 (N_18727,N_17009,N_17110);
and U18728 (N_18728,N_17449,N_17468);
and U18729 (N_18729,N_17886,N_16937);
nand U18730 (N_18730,N_17216,N_17312);
nor U18731 (N_18731,N_16964,N_17544);
nor U18732 (N_18732,N_16808,N_16938);
nand U18733 (N_18733,N_17571,N_17757);
nor U18734 (N_18734,N_17713,N_16975);
nor U18735 (N_18735,N_17396,N_17506);
xnor U18736 (N_18736,N_17667,N_17188);
xnor U18737 (N_18737,N_16953,N_17538);
nand U18738 (N_18738,N_17905,N_17796);
or U18739 (N_18739,N_17831,N_17275);
nor U18740 (N_18740,N_17953,N_17974);
xor U18741 (N_18741,N_17371,N_17342);
xor U18742 (N_18742,N_17478,N_17590);
or U18743 (N_18743,N_17033,N_17875);
or U18744 (N_18744,N_17519,N_17802);
nor U18745 (N_18745,N_17844,N_17526);
or U18746 (N_18746,N_17543,N_17987);
or U18747 (N_18747,N_17970,N_16840);
nor U18748 (N_18748,N_17325,N_17736);
xor U18749 (N_18749,N_17024,N_17329);
nand U18750 (N_18750,N_17253,N_16906);
or U18751 (N_18751,N_17837,N_17667);
nand U18752 (N_18752,N_17079,N_16893);
nand U18753 (N_18753,N_17640,N_16840);
nand U18754 (N_18754,N_17321,N_17058);
and U18755 (N_18755,N_17512,N_17050);
nand U18756 (N_18756,N_17537,N_17540);
and U18757 (N_18757,N_16879,N_17318);
nor U18758 (N_18758,N_17225,N_17710);
and U18759 (N_18759,N_17327,N_17205);
nor U18760 (N_18760,N_17760,N_17991);
or U18761 (N_18761,N_17834,N_17463);
nor U18762 (N_18762,N_17096,N_17413);
nor U18763 (N_18763,N_17802,N_17485);
or U18764 (N_18764,N_17153,N_17130);
xor U18765 (N_18765,N_17384,N_17271);
and U18766 (N_18766,N_17705,N_17034);
and U18767 (N_18767,N_17290,N_16904);
nor U18768 (N_18768,N_16926,N_17142);
and U18769 (N_18769,N_17577,N_17668);
nor U18770 (N_18770,N_17765,N_17775);
or U18771 (N_18771,N_17298,N_17938);
nor U18772 (N_18772,N_17795,N_16947);
or U18773 (N_18773,N_17157,N_17863);
and U18774 (N_18774,N_17725,N_17671);
xor U18775 (N_18775,N_16939,N_17720);
nand U18776 (N_18776,N_17399,N_17550);
nor U18777 (N_18777,N_17887,N_16810);
or U18778 (N_18778,N_17929,N_17393);
nand U18779 (N_18779,N_17838,N_17044);
or U18780 (N_18780,N_17955,N_17468);
and U18781 (N_18781,N_17990,N_17931);
or U18782 (N_18782,N_17786,N_17189);
xnor U18783 (N_18783,N_17392,N_17617);
nand U18784 (N_18784,N_17191,N_17503);
or U18785 (N_18785,N_17696,N_16980);
nor U18786 (N_18786,N_17572,N_17547);
and U18787 (N_18787,N_17108,N_17058);
and U18788 (N_18788,N_17501,N_17535);
xor U18789 (N_18789,N_17127,N_17508);
xnor U18790 (N_18790,N_17143,N_17963);
nor U18791 (N_18791,N_16880,N_17422);
nand U18792 (N_18792,N_17663,N_17648);
nand U18793 (N_18793,N_16835,N_17610);
or U18794 (N_18794,N_17516,N_17051);
nor U18795 (N_18795,N_17295,N_17887);
nor U18796 (N_18796,N_17594,N_17368);
and U18797 (N_18797,N_16922,N_17210);
nand U18798 (N_18798,N_17917,N_17967);
nor U18799 (N_18799,N_17670,N_16846);
nand U18800 (N_18800,N_16956,N_17479);
and U18801 (N_18801,N_17130,N_17860);
or U18802 (N_18802,N_17015,N_16820);
nand U18803 (N_18803,N_16890,N_16923);
nor U18804 (N_18804,N_17967,N_17364);
or U18805 (N_18805,N_17339,N_17884);
or U18806 (N_18806,N_17981,N_17268);
and U18807 (N_18807,N_17309,N_17816);
nor U18808 (N_18808,N_17685,N_16841);
and U18809 (N_18809,N_17510,N_17913);
nand U18810 (N_18810,N_17469,N_16937);
xnor U18811 (N_18811,N_17982,N_16963);
and U18812 (N_18812,N_17583,N_17719);
nand U18813 (N_18813,N_16834,N_17308);
or U18814 (N_18814,N_17239,N_17399);
nand U18815 (N_18815,N_17823,N_17086);
or U18816 (N_18816,N_17734,N_17623);
xor U18817 (N_18817,N_17526,N_17528);
xor U18818 (N_18818,N_17540,N_17590);
nor U18819 (N_18819,N_16801,N_17107);
and U18820 (N_18820,N_17628,N_17773);
nand U18821 (N_18821,N_17357,N_17059);
and U18822 (N_18822,N_16859,N_17125);
xor U18823 (N_18823,N_17928,N_17463);
nand U18824 (N_18824,N_17119,N_17312);
nor U18825 (N_18825,N_17822,N_17069);
or U18826 (N_18826,N_17036,N_17220);
nor U18827 (N_18827,N_17706,N_17044);
and U18828 (N_18828,N_17238,N_16863);
xnor U18829 (N_18829,N_16906,N_17423);
and U18830 (N_18830,N_16881,N_17865);
or U18831 (N_18831,N_17122,N_17233);
nand U18832 (N_18832,N_16805,N_17192);
nor U18833 (N_18833,N_17291,N_17199);
and U18834 (N_18834,N_17482,N_17761);
nand U18835 (N_18835,N_17874,N_17990);
or U18836 (N_18836,N_16876,N_17951);
xor U18837 (N_18837,N_17877,N_17007);
nand U18838 (N_18838,N_17421,N_17884);
and U18839 (N_18839,N_17635,N_17365);
xnor U18840 (N_18840,N_17744,N_16954);
xor U18841 (N_18841,N_17545,N_17008);
and U18842 (N_18842,N_17483,N_16864);
and U18843 (N_18843,N_17865,N_17306);
nor U18844 (N_18844,N_17424,N_17854);
nand U18845 (N_18845,N_17892,N_16915);
and U18846 (N_18846,N_17013,N_17858);
or U18847 (N_18847,N_17275,N_16826);
or U18848 (N_18848,N_17306,N_17941);
nor U18849 (N_18849,N_16829,N_17798);
nand U18850 (N_18850,N_17448,N_16838);
or U18851 (N_18851,N_17354,N_17605);
xnor U18852 (N_18852,N_17424,N_17321);
and U18853 (N_18853,N_17386,N_16927);
nand U18854 (N_18854,N_17478,N_16970);
nor U18855 (N_18855,N_17444,N_17730);
nor U18856 (N_18856,N_16881,N_17355);
nor U18857 (N_18857,N_17017,N_16932);
nand U18858 (N_18858,N_17125,N_17070);
nand U18859 (N_18859,N_17638,N_17755);
nand U18860 (N_18860,N_16901,N_17240);
nand U18861 (N_18861,N_17112,N_17532);
nor U18862 (N_18862,N_17476,N_17102);
and U18863 (N_18863,N_17262,N_17846);
nand U18864 (N_18864,N_16975,N_17249);
nor U18865 (N_18865,N_17849,N_17614);
xor U18866 (N_18866,N_17197,N_16955);
or U18867 (N_18867,N_17247,N_17074);
or U18868 (N_18868,N_17943,N_16927);
nor U18869 (N_18869,N_17403,N_16896);
and U18870 (N_18870,N_16831,N_17221);
and U18871 (N_18871,N_16843,N_16985);
xor U18872 (N_18872,N_17305,N_17966);
and U18873 (N_18873,N_17203,N_16930);
and U18874 (N_18874,N_17612,N_17067);
and U18875 (N_18875,N_17821,N_17543);
or U18876 (N_18876,N_16887,N_17514);
xor U18877 (N_18877,N_17120,N_17724);
and U18878 (N_18878,N_16882,N_17848);
and U18879 (N_18879,N_17366,N_17663);
and U18880 (N_18880,N_17285,N_17058);
and U18881 (N_18881,N_17303,N_17547);
and U18882 (N_18882,N_17572,N_17774);
or U18883 (N_18883,N_17426,N_17772);
nor U18884 (N_18884,N_17578,N_16879);
xnor U18885 (N_18885,N_17629,N_17053);
or U18886 (N_18886,N_17509,N_17534);
and U18887 (N_18887,N_17304,N_17590);
nor U18888 (N_18888,N_17195,N_17250);
and U18889 (N_18889,N_17745,N_17459);
or U18890 (N_18890,N_17036,N_16903);
nand U18891 (N_18891,N_17967,N_17605);
and U18892 (N_18892,N_17405,N_17988);
nor U18893 (N_18893,N_17126,N_17449);
or U18894 (N_18894,N_17414,N_16902);
nor U18895 (N_18895,N_17438,N_17116);
nand U18896 (N_18896,N_17315,N_17113);
or U18897 (N_18897,N_16801,N_17022);
nand U18898 (N_18898,N_17103,N_17045);
nand U18899 (N_18899,N_17052,N_16947);
or U18900 (N_18900,N_17623,N_16824);
nand U18901 (N_18901,N_16906,N_17774);
xnor U18902 (N_18902,N_17303,N_16947);
nor U18903 (N_18903,N_16888,N_17901);
or U18904 (N_18904,N_17470,N_16999);
nor U18905 (N_18905,N_17917,N_17673);
nand U18906 (N_18906,N_16869,N_17455);
nor U18907 (N_18907,N_17627,N_17341);
and U18908 (N_18908,N_17918,N_17382);
and U18909 (N_18909,N_17476,N_17559);
or U18910 (N_18910,N_17383,N_17066);
nand U18911 (N_18911,N_17387,N_17533);
or U18912 (N_18912,N_17907,N_17590);
nor U18913 (N_18913,N_16867,N_17705);
and U18914 (N_18914,N_17533,N_17296);
nor U18915 (N_18915,N_17245,N_17782);
nor U18916 (N_18916,N_17653,N_17809);
nand U18917 (N_18917,N_17387,N_17825);
nand U18918 (N_18918,N_17046,N_17498);
or U18919 (N_18919,N_16801,N_17360);
and U18920 (N_18920,N_16920,N_17126);
xnor U18921 (N_18921,N_17872,N_17772);
nor U18922 (N_18922,N_17911,N_17653);
nand U18923 (N_18923,N_17181,N_17997);
xor U18924 (N_18924,N_17735,N_17470);
xnor U18925 (N_18925,N_17524,N_17344);
nor U18926 (N_18926,N_17793,N_17758);
xnor U18927 (N_18927,N_17931,N_16877);
nand U18928 (N_18928,N_17831,N_17561);
or U18929 (N_18929,N_17083,N_17368);
or U18930 (N_18930,N_16821,N_17715);
nor U18931 (N_18931,N_17390,N_17539);
nand U18932 (N_18932,N_17937,N_17357);
nand U18933 (N_18933,N_16809,N_16930);
or U18934 (N_18934,N_17592,N_17570);
xor U18935 (N_18935,N_17105,N_17606);
nand U18936 (N_18936,N_16979,N_17605);
and U18937 (N_18937,N_17611,N_17301);
xor U18938 (N_18938,N_17521,N_17634);
and U18939 (N_18939,N_17382,N_17659);
xnor U18940 (N_18940,N_17833,N_17823);
nor U18941 (N_18941,N_16902,N_17221);
nor U18942 (N_18942,N_17523,N_16847);
xnor U18943 (N_18943,N_17812,N_17136);
or U18944 (N_18944,N_17122,N_17313);
and U18945 (N_18945,N_17334,N_17314);
or U18946 (N_18946,N_17700,N_17529);
xnor U18947 (N_18947,N_17826,N_17755);
xor U18948 (N_18948,N_17923,N_17254);
nand U18949 (N_18949,N_17386,N_17813);
nor U18950 (N_18950,N_17548,N_17912);
and U18951 (N_18951,N_17376,N_17968);
nor U18952 (N_18952,N_17705,N_17304);
nand U18953 (N_18953,N_17697,N_16842);
nor U18954 (N_18954,N_17402,N_17794);
or U18955 (N_18955,N_17911,N_16998);
nand U18956 (N_18956,N_17565,N_17460);
nor U18957 (N_18957,N_17944,N_17227);
or U18958 (N_18958,N_17888,N_17240);
nor U18959 (N_18959,N_17330,N_17792);
xor U18960 (N_18960,N_17986,N_17292);
nand U18961 (N_18961,N_17003,N_17034);
and U18962 (N_18962,N_17751,N_17281);
nand U18963 (N_18963,N_17389,N_17800);
nand U18964 (N_18964,N_16959,N_16837);
nor U18965 (N_18965,N_16849,N_17734);
xnor U18966 (N_18966,N_17438,N_17980);
and U18967 (N_18967,N_17749,N_17816);
and U18968 (N_18968,N_17759,N_17140);
or U18969 (N_18969,N_17872,N_17202);
nor U18970 (N_18970,N_17373,N_17986);
and U18971 (N_18971,N_17904,N_17381);
and U18972 (N_18972,N_17725,N_17402);
and U18973 (N_18973,N_16878,N_17159);
or U18974 (N_18974,N_17852,N_16866);
and U18975 (N_18975,N_17944,N_16910);
or U18976 (N_18976,N_17743,N_17132);
nor U18977 (N_18977,N_16851,N_17647);
or U18978 (N_18978,N_16842,N_17710);
xnor U18979 (N_18979,N_17996,N_17944);
nor U18980 (N_18980,N_17391,N_17354);
or U18981 (N_18981,N_16838,N_17069);
nand U18982 (N_18982,N_17877,N_17934);
xnor U18983 (N_18983,N_17196,N_16849);
or U18984 (N_18984,N_17627,N_16815);
nor U18985 (N_18985,N_17038,N_16912);
nor U18986 (N_18986,N_17492,N_17551);
nand U18987 (N_18987,N_17700,N_17556);
and U18988 (N_18988,N_17588,N_16975);
or U18989 (N_18989,N_16959,N_17432);
nand U18990 (N_18990,N_17267,N_17563);
xnor U18991 (N_18991,N_17220,N_17532);
and U18992 (N_18992,N_16880,N_17338);
nand U18993 (N_18993,N_17320,N_17795);
nor U18994 (N_18994,N_17319,N_17459);
and U18995 (N_18995,N_17192,N_17286);
nand U18996 (N_18996,N_16981,N_17151);
or U18997 (N_18997,N_17013,N_16911);
nand U18998 (N_18998,N_16880,N_17717);
or U18999 (N_18999,N_16970,N_17589);
nor U19000 (N_19000,N_17888,N_17273);
or U19001 (N_19001,N_17053,N_17344);
and U19002 (N_19002,N_17090,N_17859);
nor U19003 (N_19003,N_17051,N_17432);
or U19004 (N_19004,N_17262,N_17197);
xnor U19005 (N_19005,N_17147,N_17658);
or U19006 (N_19006,N_17204,N_17977);
xor U19007 (N_19007,N_17716,N_16851);
nand U19008 (N_19008,N_17534,N_17757);
or U19009 (N_19009,N_17796,N_17379);
nand U19010 (N_19010,N_17114,N_17909);
and U19011 (N_19011,N_17125,N_17408);
or U19012 (N_19012,N_17038,N_16933);
and U19013 (N_19013,N_17081,N_17216);
xor U19014 (N_19014,N_17486,N_17766);
nand U19015 (N_19015,N_16938,N_17991);
nand U19016 (N_19016,N_17977,N_17912);
or U19017 (N_19017,N_17120,N_17004);
nand U19018 (N_19018,N_17543,N_17247);
xor U19019 (N_19019,N_16830,N_17780);
nor U19020 (N_19020,N_17504,N_17401);
nor U19021 (N_19021,N_17950,N_17879);
nor U19022 (N_19022,N_17010,N_17100);
nor U19023 (N_19023,N_17763,N_17350);
and U19024 (N_19024,N_17124,N_17674);
and U19025 (N_19025,N_17756,N_17792);
and U19026 (N_19026,N_17069,N_17742);
nand U19027 (N_19027,N_17287,N_16947);
nor U19028 (N_19028,N_17132,N_17285);
and U19029 (N_19029,N_16876,N_17058);
nor U19030 (N_19030,N_17473,N_17774);
or U19031 (N_19031,N_17081,N_17943);
or U19032 (N_19032,N_17128,N_17869);
and U19033 (N_19033,N_16842,N_17417);
or U19034 (N_19034,N_17526,N_17136);
nand U19035 (N_19035,N_17545,N_17389);
and U19036 (N_19036,N_17454,N_17672);
or U19037 (N_19037,N_16897,N_17144);
nor U19038 (N_19038,N_16837,N_17991);
nor U19039 (N_19039,N_17363,N_16930);
and U19040 (N_19040,N_16937,N_17962);
xnor U19041 (N_19041,N_17396,N_17333);
and U19042 (N_19042,N_17649,N_17480);
or U19043 (N_19043,N_17939,N_17231);
xor U19044 (N_19044,N_17889,N_17994);
or U19045 (N_19045,N_17279,N_17360);
xor U19046 (N_19046,N_16944,N_16942);
or U19047 (N_19047,N_17067,N_17217);
xor U19048 (N_19048,N_17550,N_17751);
or U19049 (N_19049,N_17849,N_17982);
and U19050 (N_19050,N_17841,N_17969);
nand U19051 (N_19051,N_16980,N_17474);
or U19052 (N_19052,N_17173,N_17485);
or U19053 (N_19053,N_17809,N_17484);
or U19054 (N_19054,N_16913,N_17034);
nand U19055 (N_19055,N_17993,N_17454);
xnor U19056 (N_19056,N_16810,N_17280);
or U19057 (N_19057,N_17903,N_17898);
nor U19058 (N_19058,N_17920,N_17936);
and U19059 (N_19059,N_16870,N_17720);
nand U19060 (N_19060,N_17648,N_17243);
xnor U19061 (N_19061,N_17108,N_17599);
nand U19062 (N_19062,N_17517,N_17003);
or U19063 (N_19063,N_17111,N_17814);
xor U19064 (N_19064,N_17130,N_17441);
and U19065 (N_19065,N_17587,N_17364);
nor U19066 (N_19066,N_17426,N_17264);
nand U19067 (N_19067,N_17614,N_17799);
xnor U19068 (N_19068,N_17590,N_17668);
or U19069 (N_19069,N_16915,N_17715);
or U19070 (N_19070,N_17733,N_17960);
or U19071 (N_19071,N_17491,N_17531);
nor U19072 (N_19072,N_17494,N_17116);
xnor U19073 (N_19073,N_17313,N_17899);
or U19074 (N_19074,N_17632,N_17277);
and U19075 (N_19075,N_16969,N_17206);
nor U19076 (N_19076,N_17736,N_17424);
or U19077 (N_19077,N_17570,N_16817);
nand U19078 (N_19078,N_17030,N_17858);
nand U19079 (N_19079,N_17794,N_17857);
and U19080 (N_19080,N_17209,N_17328);
xnor U19081 (N_19081,N_17677,N_17456);
and U19082 (N_19082,N_17030,N_16847);
or U19083 (N_19083,N_17476,N_17607);
or U19084 (N_19084,N_17100,N_17473);
xnor U19085 (N_19085,N_17410,N_17568);
or U19086 (N_19086,N_17453,N_17505);
or U19087 (N_19087,N_17847,N_17082);
and U19088 (N_19088,N_17189,N_17461);
nor U19089 (N_19089,N_17794,N_17993);
nor U19090 (N_19090,N_17507,N_17537);
nand U19091 (N_19091,N_16829,N_17377);
and U19092 (N_19092,N_17824,N_16861);
or U19093 (N_19093,N_17030,N_17131);
or U19094 (N_19094,N_17987,N_17937);
or U19095 (N_19095,N_17325,N_17638);
nand U19096 (N_19096,N_17895,N_17833);
and U19097 (N_19097,N_17736,N_17252);
nor U19098 (N_19098,N_17425,N_17182);
nor U19099 (N_19099,N_17577,N_16956);
and U19100 (N_19100,N_17216,N_17381);
or U19101 (N_19101,N_17630,N_17026);
and U19102 (N_19102,N_17173,N_17497);
or U19103 (N_19103,N_16839,N_17541);
nor U19104 (N_19104,N_16944,N_17325);
xnor U19105 (N_19105,N_16922,N_17444);
and U19106 (N_19106,N_17143,N_17600);
nor U19107 (N_19107,N_17914,N_17225);
and U19108 (N_19108,N_17722,N_17012);
nor U19109 (N_19109,N_17372,N_17108);
nand U19110 (N_19110,N_17550,N_17302);
or U19111 (N_19111,N_17752,N_17720);
nand U19112 (N_19112,N_16991,N_17177);
and U19113 (N_19113,N_16850,N_17248);
and U19114 (N_19114,N_17632,N_16836);
and U19115 (N_19115,N_17664,N_16854);
nand U19116 (N_19116,N_17679,N_17643);
and U19117 (N_19117,N_16938,N_17978);
or U19118 (N_19118,N_17778,N_17223);
and U19119 (N_19119,N_17253,N_17989);
or U19120 (N_19120,N_17531,N_17185);
nand U19121 (N_19121,N_17823,N_17617);
or U19122 (N_19122,N_17462,N_17578);
and U19123 (N_19123,N_17771,N_17836);
xnor U19124 (N_19124,N_16802,N_16933);
nor U19125 (N_19125,N_16936,N_17670);
or U19126 (N_19126,N_17120,N_17013);
and U19127 (N_19127,N_17166,N_16864);
nor U19128 (N_19128,N_17285,N_17126);
and U19129 (N_19129,N_17936,N_17657);
nand U19130 (N_19130,N_17010,N_17874);
nand U19131 (N_19131,N_17360,N_17552);
or U19132 (N_19132,N_17732,N_17475);
xor U19133 (N_19133,N_16943,N_17698);
and U19134 (N_19134,N_16939,N_16965);
xor U19135 (N_19135,N_17794,N_17678);
nor U19136 (N_19136,N_17781,N_17682);
and U19137 (N_19137,N_17514,N_17356);
and U19138 (N_19138,N_16912,N_17796);
or U19139 (N_19139,N_17523,N_17704);
xnor U19140 (N_19140,N_17810,N_17540);
or U19141 (N_19141,N_16851,N_17123);
or U19142 (N_19142,N_16863,N_17845);
or U19143 (N_19143,N_17636,N_17908);
xnor U19144 (N_19144,N_17452,N_17969);
or U19145 (N_19145,N_16884,N_17925);
nand U19146 (N_19146,N_16986,N_16957);
nand U19147 (N_19147,N_17498,N_17129);
nand U19148 (N_19148,N_17852,N_17098);
and U19149 (N_19149,N_16965,N_17276);
nand U19150 (N_19150,N_17040,N_17183);
or U19151 (N_19151,N_16939,N_16960);
or U19152 (N_19152,N_17105,N_17008);
or U19153 (N_19153,N_16898,N_17137);
and U19154 (N_19154,N_17240,N_17795);
and U19155 (N_19155,N_17665,N_17759);
nor U19156 (N_19156,N_17153,N_17806);
xor U19157 (N_19157,N_16904,N_17047);
or U19158 (N_19158,N_17142,N_17803);
or U19159 (N_19159,N_17348,N_17672);
nor U19160 (N_19160,N_17303,N_17448);
xnor U19161 (N_19161,N_17738,N_17181);
nor U19162 (N_19162,N_16922,N_17934);
nand U19163 (N_19163,N_17201,N_17695);
nand U19164 (N_19164,N_17977,N_17968);
or U19165 (N_19165,N_16936,N_17892);
or U19166 (N_19166,N_17780,N_16870);
and U19167 (N_19167,N_17422,N_17291);
nand U19168 (N_19168,N_17313,N_16939);
or U19169 (N_19169,N_17740,N_17259);
xor U19170 (N_19170,N_17174,N_17955);
or U19171 (N_19171,N_17101,N_17025);
or U19172 (N_19172,N_16809,N_17537);
nor U19173 (N_19173,N_17187,N_17249);
nor U19174 (N_19174,N_17816,N_17160);
nor U19175 (N_19175,N_17183,N_17342);
and U19176 (N_19176,N_16804,N_16877);
nand U19177 (N_19177,N_17528,N_17926);
nand U19178 (N_19178,N_16815,N_16893);
and U19179 (N_19179,N_17539,N_17031);
and U19180 (N_19180,N_17785,N_17030);
and U19181 (N_19181,N_17404,N_17610);
and U19182 (N_19182,N_17242,N_17597);
nand U19183 (N_19183,N_17678,N_17056);
or U19184 (N_19184,N_17180,N_16915);
and U19185 (N_19185,N_16843,N_17537);
and U19186 (N_19186,N_17893,N_17923);
nor U19187 (N_19187,N_17048,N_17400);
nand U19188 (N_19188,N_17130,N_17692);
or U19189 (N_19189,N_17769,N_17934);
nor U19190 (N_19190,N_17850,N_17859);
nor U19191 (N_19191,N_16862,N_16948);
nand U19192 (N_19192,N_17378,N_17602);
or U19193 (N_19193,N_17583,N_17878);
and U19194 (N_19194,N_17560,N_16811);
and U19195 (N_19195,N_17418,N_17767);
nor U19196 (N_19196,N_17648,N_17748);
or U19197 (N_19197,N_17072,N_16928);
xnor U19198 (N_19198,N_17516,N_17533);
xor U19199 (N_19199,N_17706,N_17566);
or U19200 (N_19200,N_18334,N_18695);
and U19201 (N_19201,N_18245,N_18272);
and U19202 (N_19202,N_18857,N_18293);
xnor U19203 (N_19203,N_18543,N_18175);
xnor U19204 (N_19204,N_18410,N_18460);
nor U19205 (N_19205,N_18082,N_18495);
nor U19206 (N_19206,N_19167,N_18990);
nand U19207 (N_19207,N_18562,N_18934);
nand U19208 (N_19208,N_18653,N_18737);
or U19209 (N_19209,N_18763,N_19004);
or U19210 (N_19210,N_18076,N_18059);
xor U19211 (N_19211,N_18137,N_19165);
nand U19212 (N_19212,N_18729,N_19186);
nand U19213 (N_19213,N_18218,N_18777);
or U19214 (N_19214,N_18000,N_19093);
xor U19215 (N_19215,N_18336,N_18483);
or U19216 (N_19216,N_18269,N_18103);
nand U19217 (N_19217,N_18920,N_18735);
nand U19218 (N_19218,N_19045,N_18120);
xor U19219 (N_19219,N_18100,N_18459);
nor U19220 (N_19220,N_19001,N_18162);
nor U19221 (N_19221,N_18654,N_18692);
nor U19222 (N_19222,N_18865,N_18933);
nor U19223 (N_19223,N_18730,N_18590);
and U19224 (N_19224,N_18870,N_18343);
or U19225 (N_19225,N_18772,N_18111);
nor U19226 (N_19226,N_18889,N_18009);
nand U19227 (N_19227,N_19048,N_18637);
nor U19228 (N_19228,N_18922,N_18971);
or U19229 (N_19229,N_19156,N_18426);
nor U19230 (N_19230,N_19053,N_18458);
xnor U19231 (N_19231,N_18386,N_18455);
or U19232 (N_19232,N_18391,N_18212);
xor U19233 (N_19233,N_18174,N_19192);
nand U19234 (N_19234,N_18449,N_18157);
or U19235 (N_19235,N_18819,N_18936);
or U19236 (N_19236,N_18412,N_18315);
nand U19237 (N_19237,N_18324,N_18633);
or U19238 (N_19238,N_18658,N_18159);
xor U19239 (N_19239,N_18660,N_18504);
nand U19240 (N_19240,N_18206,N_18131);
nand U19241 (N_19241,N_19163,N_19194);
xor U19242 (N_19242,N_18479,N_18609);
and U19243 (N_19243,N_18327,N_18310);
nor U19244 (N_19244,N_18491,N_18707);
and U19245 (N_19245,N_18210,N_19063);
or U19246 (N_19246,N_18438,N_18568);
nor U19247 (N_19247,N_18330,N_18624);
or U19248 (N_19248,N_19034,N_18924);
and U19249 (N_19249,N_19160,N_18985);
and U19250 (N_19250,N_18615,N_18860);
and U19251 (N_19251,N_18115,N_18164);
and U19252 (N_19252,N_18112,N_18379);
nand U19253 (N_19253,N_18943,N_18283);
and U19254 (N_19254,N_18812,N_18055);
nand U19255 (N_19255,N_18868,N_18418);
nor U19256 (N_19256,N_19044,N_18625);
nor U19257 (N_19257,N_18632,N_19091);
xor U19258 (N_19258,N_18688,N_18205);
nor U19259 (N_19259,N_18058,N_18903);
nor U19260 (N_19260,N_19189,N_18592);
or U19261 (N_19261,N_18011,N_18533);
nand U19262 (N_19262,N_18344,N_18117);
nand U19263 (N_19263,N_18193,N_18908);
nor U19264 (N_19264,N_18430,N_18199);
xnor U19265 (N_19265,N_18361,N_19134);
xor U19266 (N_19266,N_18958,N_18671);
nor U19267 (N_19267,N_19110,N_18030);
nor U19268 (N_19268,N_18997,N_18496);
xor U19269 (N_19269,N_18298,N_18874);
or U19270 (N_19270,N_18196,N_18045);
nand U19271 (N_19271,N_18313,N_18542);
or U19272 (N_19272,N_18034,N_18537);
or U19273 (N_19273,N_18250,N_18176);
xnor U19274 (N_19274,N_18647,N_18099);
xor U19275 (N_19275,N_18947,N_18895);
nor U19276 (N_19276,N_19016,N_18130);
and U19277 (N_19277,N_18505,N_18022);
xnor U19278 (N_19278,N_18687,N_18492);
nor U19279 (N_19279,N_18377,N_19132);
or U19280 (N_19280,N_18876,N_18114);
nor U19281 (N_19281,N_18864,N_18887);
nand U19282 (N_19282,N_18536,N_18309);
or U19283 (N_19283,N_18754,N_18720);
nand U19284 (N_19284,N_18502,N_18926);
and U19285 (N_19285,N_18843,N_18626);
or U19286 (N_19286,N_18408,N_18335);
nand U19287 (N_19287,N_18078,N_18349);
xnor U19288 (N_19288,N_18200,N_18622);
nand U19289 (N_19289,N_19133,N_19083);
and U19290 (N_19290,N_18708,N_18833);
nor U19291 (N_19291,N_18643,N_18963);
nand U19292 (N_19292,N_18796,N_18136);
nor U19293 (N_19293,N_18840,N_19169);
nand U19294 (N_19294,N_18056,N_18716);
and U19295 (N_19295,N_18650,N_18888);
or U19296 (N_19296,N_18527,N_18564);
and U19297 (N_19297,N_18935,N_19006);
xnor U19298 (N_19298,N_18565,N_18029);
nand U19299 (N_19299,N_18785,N_18705);
xnor U19300 (N_19300,N_18149,N_18538);
or U19301 (N_19301,N_18567,N_18719);
xnor U19302 (N_19302,N_18163,N_18422);
nand U19303 (N_19303,N_18991,N_19164);
nand U19304 (N_19304,N_18823,N_18975);
and U19305 (N_19305,N_19028,N_18247);
xor U19306 (N_19306,N_19181,N_18064);
nand U19307 (N_19307,N_18147,N_18745);
nor U19308 (N_19308,N_19137,N_18614);
nor U19309 (N_19309,N_18608,N_19066);
nor U19310 (N_19310,N_18445,N_18101);
xor U19311 (N_19311,N_18976,N_19150);
nor U19312 (N_19312,N_18851,N_18603);
or U19313 (N_19313,N_18532,N_18656);
or U19314 (N_19314,N_18649,N_19199);
nor U19315 (N_19315,N_18073,N_18522);
or U19316 (N_19316,N_18311,N_18489);
nor U19317 (N_19317,N_18747,N_18437);
and U19318 (N_19318,N_18528,N_18487);
xor U19319 (N_19319,N_19022,N_18681);
or U19320 (N_19320,N_19090,N_18731);
and U19321 (N_19321,N_18993,N_18042);
or U19322 (N_19322,N_18519,N_19040);
xnor U19323 (N_19323,N_18146,N_18791);
nand U19324 (N_19324,N_18395,N_18712);
nand U19325 (N_19325,N_18139,N_19043);
and U19326 (N_19326,N_19007,N_18267);
nor U19327 (N_19327,N_18684,N_18113);
xnor U19328 (N_19328,N_18160,N_18914);
nor U19329 (N_19329,N_19099,N_18493);
or U19330 (N_19330,N_18301,N_18303);
xor U19331 (N_19331,N_18424,N_18655);
xnor U19332 (N_19332,N_18203,N_18127);
nand U19333 (N_19333,N_18524,N_18413);
and U19334 (N_19334,N_18017,N_18988);
and U19335 (N_19335,N_18704,N_18815);
xnor U19336 (N_19336,N_18185,N_18748);
xnor U19337 (N_19337,N_18454,N_18967);
nand U19338 (N_19338,N_18631,N_19180);
nand U19339 (N_19339,N_18371,N_19069);
nand U19340 (N_19340,N_18084,N_18883);
or U19341 (N_19341,N_19144,N_18043);
or U19342 (N_19342,N_18096,N_18217);
and U19343 (N_19343,N_18342,N_18404);
or U19344 (N_19344,N_19023,N_18921);
nand U19345 (N_19345,N_18167,N_18530);
or U19346 (N_19346,N_18784,N_18884);
or U19347 (N_19347,N_18599,N_19036);
nor U19348 (N_19348,N_19191,N_18387);
nor U19349 (N_19349,N_18144,N_18916);
nand U19350 (N_19350,N_18586,N_19088);
nand U19351 (N_19351,N_18578,N_18954);
nand U19352 (N_19352,N_18125,N_18415);
or U19353 (N_19353,N_18634,N_18831);
nor U19354 (N_19354,N_18501,N_18845);
or U19355 (N_19355,N_18825,N_18222);
nand U19356 (N_19356,N_18420,N_18786);
or U19357 (N_19357,N_19012,N_18558);
xor U19358 (N_19358,N_18589,N_18952);
xor U19359 (N_19359,N_18025,N_18927);
nand U19360 (N_19360,N_18587,N_19195);
nand U19361 (N_19361,N_18063,N_19080);
and U19362 (N_19362,N_18242,N_18028);
and U19363 (N_19363,N_18828,N_18286);
or U19364 (N_19364,N_18328,N_19139);
nand U19365 (N_19365,N_19153,N_18014);
xor U19366 (N_19366,N_18497,N_18102);
and U19367 (N_19367,N_18544,N_18427);
and U19368 (N_19368,N_18554,N_18620);
nor U19369 (N_19369,N_18238,N_18663);
xnor U19370 (N_19370,N_19136,N_19027);
or U19371 (N_19371,N_18559,N_19055);
or U19372 (N_19372,N_18472,N_18989);
and U19373 (N_19373,N_19096,N_18691);
or U19374 (N_19374,N_18667,N_18621);
nor U19375 (N_19375,N_18782,N_18094);
nor U19376 (N_19376,N_18674,N_18640);
and U19377 (N_19377,N_19135,N_19077);
xnor U19378 (N_19378,N_19021,N_18290);
or U19379 (N_19379,N_19094,N_18095);
nor U19380 (N_19380,N_18261,N_18573);
nor U19381 (N_19381,N_18075,N_18680);
nor U19382 (N_19382,N_18436,N_18141);
nand U19383 (N_19383,N_18246,N_18188);
nor U19384 (N_19384,N_19052,N_18722);
or U19385 (N_19385,N_19108,N_19073);
and U19386 (N_19386,N_18440,N_18428);
xor U19387 (N_19387,N_19057,N_18539);
nand U19388 (N_19388,N_18541,N_18570);
xnor U19389 (N_19389,N_18739,N_18992);
and U19390 (N_19390,N_18208,N_18638);
xnor U19391 (N_19391,N_18588,N_18824);
nand U19392 (N_19392,N_18251,N_18968);
and U19393 (N_19393,N_18790,N_18381);
xor U19394 (N_19394,N_18597,N_18257);
nand U19395 (N_19395,N_18662,N_18219);
nor U19396 (N_19396,N_18723,N_18288);
nand U19397 (N_19397,N_18521,N_18929);
or U19398 (N_19398,N_19020,N_18803);
and U19399 (N_19399,N_18186,N_19092);
or U19400 (N_19400,N_18995,N_18296);
nand U19401 (N_19401,N_18338,N_18134);
nand U19402 (N_19402,N_18154,N_18977);
nor U19403 (N_19403,N_18177,N_18611);
nand U19404 (N_19404,N_18123,N_18917);
and U19405 (N_19405,N_18444,N_18646);
or U19406 (N_19406,N_19079,N_18804);
nand U19407 (N_19407,N_18322,N_18223);
xor U19408 (N_19408,N_18086,N_18026);
nand U19409 (N_19409,N_18821,N_18902);
or U19410 (N_19410,N_18035,N_18792);
or U19411 (N_19411,N_18757,N_18023);
nor U19412 (N_19412,N_18983,N_18696);
xor U19413 (N_19413,N_18467,N_18572);
and U19414 (N_19414,N_18861,N_19041);
nor U19415 (N_19415,N_19078,N_18179);
nor U19416 (N_19416,N_18087,N_18666);
nor U19417 (N_19417,N_18469,N_19178);
and U19418 (N_19418,N_18192,N_18996);
or U19419 (N_19419,N_18582,N_18940);
or U19420 (N_19420,N_19114,N_19126);
nand U19421 (N_19421,N_18080,N_18260);
xnor U19422 (N_19422,N_18569,N_19015);
and U19423 (N_19423,N_19017,N_18018);
and U19424 (N_19424,N_18794,N_18979);
nand U19425 (N_19425,N_18189,N_19193);
nand U19426 (N_19426,N_18198,N_18826);
and U19427 (N_19427,N_18165,N_18394);
nand U19428 (N_19428,N_18751,N_18284);
xor U19429 (N_19429,N_18306,N_19119);
and U19430 (N_19430,N_18066,N_18523);
nor U19431 (N_19431,N_18004,N_18067);
or U19432 (N_19432,N_18312,N_18282);
or U19433 (N_19433,N_18686,N_18685);
and U19434 (N_19434,N_18512,N_19148);
or U19435 (N_19435,N_18836,N_18417);
and U19436 (N_19436,N_18446,N_18276);
nand U19437 (N_19437,N_18170,N_18919);
or U19438 (N_19438,N_19098,N_18697);
and U19439 (N_19439,N_18750,N_19087);
nor U19440 (N_19440,N_18002,N_19060);
nand U19441 (N_19441,N_18001,N_18959);
and U19442 (N_19442,N_19158,N_18098);
nor U19443 (N_19443,N_18248,N_19033);
xor U19444 (N_19444,N_18606,N_19118);
or U19445 (N_19445,N_18419,N_18333);
or U19446 (N_19446,N_19140,N_18859);
nor U19447 (N_19447,N_18846,N_18788);
or U19448 (N_19448,N_18510,N_18879);
nand U19449 (N_19449,N_18951,N_18116);
nand U19450 (N_19450,N_18345,N_19071);
and U19451 (N_19451,N_18725,N_18027);
nand U19452 (N_19452,N_19068,N_19086);
nor U19453 (N_19453,N_18768,N_19184);
and U19454 (N_19454,N_18822,N_19032);
nor U19455 (N_19455,N_18249,N_19177);
and U19456 (N_19456,N_18885,N_19176);
nand U19457 (N_19457,N_18365,N_18264);
or U19458 (N_19458,N_18357,N_18341);
and U19459 (N_19459,N_19011,N_19122);
nor U19460 (N_19460,N_19105,N_18867);
or U19461 (N_19461,N_18372,N_19005);
and U19462 (N_19462,N_19111,N_18271);
nor U19463 (N_19463,N_18853,N_18962);
or U19464 (N_19464,N_18468,N_18856);
and U19465 (N_19465,N_19190,N_19101);
and U19466 (N_19466,N_18659,N_18106);
nor U19467 (N_19467,N_18414,N_19138);
nor U19468 (N_19468,N_18299,N_18292);
or U19469 (N_19469,N_18928,N_18239);
nand U19470 (N_19470,N_19116,N_18183);
and U19471 (N_19471,N_18227,N_18596);
or U19472 (N_19472,N_18966,N_18911);
xor U19473 (N_19473,N_18266,N_19065);
nand U19474 (N_19474,N_18462,N_18944);
and U19475 (N_19475,N_18746,N_18555);
or U19476 (N_19476,N_18918,N_18132);
or U19477 (N_19477,N_18892,N_18254);
or U19478 (N_19478,N_18579,N_19143);
or U19479 (N_19479,N_18535,N_18253);
and U19480 (N_19480,N_18965,N_18442);
xnor U19481 (N_19481,N_19067,N_18820);
nand U19482 (N_19482,N_18482,N_18051);
and U19483 (N_19483,N_19076,N_19081);
or U19484 (N_19484,N_18678,N_18577);
nor U19485 (N_19485,N_18202,N_18566);
xor U19486 (N_19486,N_18774,N_18370);
nand U19487 (N_19487,N_18872,N_18268);
nand U19488 (N_19488,N_19051,N_18829);
nor U19489 (N_19489,N_19030,N_19100);
xor U19490 (N_19490,N_18133,N_18509);
xnor U19491 (N_19491,N_18600,N_19024);
nand U19492 (N_19492,N_18500,N_18848);
or U19493 (N_19493,N_18576,N_18121);
nor U19494 (N_19494,N_18710,N_18040);
nor U19495 (N_19495,N_18435,N_18337);
and U19496 (N_19496,N_18138,N_18648);
or U19497 (N_19497,N_18668,N_18973);
nor U19498 (N_19498,N_18129,N_18727);
nor U19499 (N_19499,N_19107,N_18092);
xnor U19500 (N_19500,N_18873,N_18899);
xnor U19501 (N_19501,N_19145,N_18863);
and U19502 (N_19502,N_18764,N_18946);
xnor U19503 (N_19503,N_18817,N_18854);
xor U19504 (N_19504,N_18407,N_19025);
nand U19505 (N_19505,N_18516,N_18097);
and U19506 (N_19506,N_18894,N_19154);
and U19507 (N_19507,N_18783,N_18109);
and U19508 (N_19508,N_18838,N_18358);
nor U19509 (N_19509,N_19149,N_18265);
and U19510 (N_19510,N_18463,N_18302);
nand U19511 (N_19511,N_19120,N_18964);
nand U19512 (N_19512,N_18583,N_18173);
nand U19513 (N_19513,N_18942,N_18229);
or U19514 (N_19514,N_18373,N_18484);
nand U19515 (N_19515,N_19141,N_18220);
xnor U19516 (N_19516,N_18755,N_18970);
and U19517 (N_19517,N_19046,N_18221);
or U19518 (N_19518,N_18999,N_18461);
and U19519 (N_19519,N_18024,N_19035);
nand U19520 (N_19520,N_18316,N_19026);
xor U19521 (N_19521,N_18912,N_18672);
xor U19522 (N_19522,N_18610,N_18474);
xor U19523 (N_19523,N_18485,N_19064);
nand U19524 (N_19524,N_18213,N_18925);
xnor U19525 (N_19525,N_18593,N_18477);
nor U19526 (N_19526,N_18340,N_18279);
xor U19527 (N_19527,N_18694,N_18012);
nor U19528 (N_19528,N_18057,N_18368);
xor U19529 (N_19529,N_18779,N_18955);
or U19530 (N_19530,N_19029,N_18464);
and U19531 (N_19531,N_18190,N_18156);
nand U19532 (N_19532,N_18581,N_18802);
nand U19533 (N_19533,N_19173,N_18256);
nand U19534 (N_19534,N_18211,N_18814);
nor U19535 (N_19535,N_18457,N_18923);
nor U19536 (N_19536,N_18007,N_18771);
xnor U19537 (N_19537,N_18617,N_18550);
nor U19538 (N_19538,N_18258,N_18367);
xor U19539 (N_19539,N_18711,N_18354);
and U19540 (N_19540,N_19103,N_19050);
nor U19541 (N_19541,N_18339,N_19059);
or U19542 (N_19542,N_18263,N_18978);
xor U19543 (N_19543,N_18201,N_18307);
or U19544 (N_19544,N_18932,N_19121);
or U19545 (N_19545,N_18397,N_18518);
or U19546 (N_19546,N_18050,N_19061);
nand U19547 (N_19547,N_18628,N_18741);
and U19548 (N_19548,N_18432,N_18937);
or U19549 (N_19549,N_18652,N_18321);
and U19550 (N_19550,N_18036,N_18886);
nand U19551 (N_19551,N_18305,N_18070);
nor U19552 (N_19552,N_18601,N_18753);
and U19553 (N_19553,N_19038,N_19159);
nand U19554 (N_19554,N_18724,N_18068);
nor U19555 (N_19555,N_18297,N_18388);
nor U19556 (N_19556,N_18475,N_18118);
nor U19557 (N_19557,N_19131,N_18734);
nor U19558 (N_19558,N_18618,N_18171);
or U19559 (N_19559,N_18945,N_18897);
nor U19560 (N_19560,N_18204,N_18182);
xnor U19561 (N_19561,N_18398,N_18252);
and U19562 (N_19562,N_18168,N_19072);
and U19563 (N_19563,N_18225,N_18645);
xor U19564 (N_19564,N_18178,N_18287);
xor U19565 (N_19565,N_18304,N_18557);
xor U19566 (N_19566,N_18805,N_18380);
xnor U19567 (N_19567,N_18441,N_18604);
nand U19568 (N_19568,N_18346,N_18285);
xor U19569 (N_19569,N_18244,N_18364);
xor U19570 (N_19570,N_19062,N_18061);
xor U19571 (N_19571,N_18800,N_18142);
and U19572 (N_19572,N_18866,N_18957);
or U19573 (N_19573,N_18049,N_18396);
or U19574 (N_19574,N_18547,N_18953);
xor U19575 (N_19575,N_18683,N_18355);
xor U19576 (N_19576,N_18350,N_18984);
xnor U19577 (N_19577,N_18682,N_18300);
or U19578 (N_19578,N_18161,N_19128);
xor U19579 (N_19579,N_18037,N_18780);
or U19580 (N_19580,N_18661,N_18675);
or U19581 (N_19581,N_18839,N_18237);
nor U19582 (N_19582,N_18871,N_19089);
xnor U19583 (N_19583,N_18689,N_18972);
nand U19584 (N_19584,N_18122,N_18020);
and U19585 (N_19585,N_18706,N_19019);
and U19586 (N_19586,N_18560,N_18291);
xnor U19587 (N_19587,N_18069,N_18773);
nand U19588 (N_19588,N_18882,N_18834);
xor U19589 (N_19589,N_18893,N_19102);
xor U19590 (N_19590,N_18273,N_18382);
xor U19591 (N_19591,N_18451,N_18015);
xnor U19592 (N_19592,N_18629,N_18531);
nor U19593 (N_19593,N_18770,N_18875);
or U19594 (N_19594,N_18644,N_18197);
xnor U19595 (N_19595,N_18664,N_18514);
and U19596 (N_19596,N_18209,N_18904);
nor U19597 (N_19597,N_18347,N_18801);
xnor U19598 (N_19598,N_18758,N_19000);
and U19599 (N_19599,N_18584,N_19185);
or U19600 (N_19600,N_18961,N_18478);
and U19601 (N_19601,N_18761,N_18053);
or U19602 (N_19602,N_18486,N_18466);
nor U19603 (N_19603,N_18690,N_18850);
or U19604 (N_19604,N_18191,N_18392);
or U19605 (N_19605,N_18383,N_18448);
nand U19606 (N_19606,N_18549,N_19146);
and U19607 (N_19607,N_18849,N_18752);
or U19608 (N_19608,N_18169,N_18808);
xor U19609 (N_19609,N_18013,N_18709);
nand U19610 (N_19610,N_18409,N_18797);
nand U19611 (N_19611,N_18974,N_18228);
nor U19612 (N_19612,N_18939,N_19174);
xnor U19613 (N_19613,N_18670,N_18736);
or U19614 (N_19614,N_18948,N_18135);
xor U19615 (N_19615,N_18702,N_18799);
xor U19616 (N_19616,N_18006,N_18548);
nand U19617 (N_19617,N_18830,N_18809);
nor U19618 (N_19618,N_18047,N_18280);
and U19619 (N_19619,N_19170,N_18403);
nand U19620 (N_19620,N_19009,N_19049);
and U19621 (N_19621,N_18835,N_18743);
and U19622 (N_19622,N_18390,N_18525);
nor U19623 (N_19623,N_18148,N_18226);
or U19624 (N_19624,N_18807,N_18465);
or U19625 (N_19625,N_18145,N_19039);
xnor U19626 (N_19626,N_18635,N_18806);
nor U19627 (N_19627,N_18529,N_18143);
nand U19628 (N_19628,N_19018,N_18540);
or U19629 (N_19629,N_18488,N_18278);
or U19630 (N_19630,N_18054,N_18910);
nand U19631 (N_19631,N_18032,N_18842);
nor U19632 (N_19632,N_19166,N_19113);
xnor U19633 (N_19633,N_18930,N_18277);
nor U19634 (N_19634,N_18520,N_18571);
and U19635 (N_19635,N_18423,N_19109);
xor U19636 (N_19636,N_19123,N_18270);
xnor U19637 (N_19637,N_18091,N_19162);
nor U19638 (N_19638,N_18490,N_18281);
nand U19639 (N_19639,N_18950,N_19196);
nor U19640 (N_19640,N_19168,N_18362);
nand U19641 (N_19641,N_19008,N_18595);
and U19642 (N_19642,N_18005,N_18766);
nor U19643 (N_19643,N_18642,N_19056);
nand U19644 (N_19644,N_18781,N_18447);
or U19645 (N_19645,N_18847,N_18443);
xor U19646 (N_19646,N_18890,N_18065);
nand U19647 (N_19647,N_18598,N_18259);
and U19648 (N_19648,N_18616,N_18008);
nor U19649 (N_19649,N_18869,N_19106);
nand U19650 (N_19650,N_18074,N_19198);
nand U19651 (N_19651,N_18207,N_18400);
xor U19652 (N_19652,N_18793,N_18378);
or U19653 (N_19653,N_18798,N_18733);
xnor U19654 (N_19654,N_18552,N_18233);
xnor U19655 (N_19655,N_18150,N_18240);
xnor U19656 (N_19656,N_18318,N_18314);
nand U19657 (N_19657,N_18375,N_19095);
nor U19658 (N_19658,N_18083,N_18982);
nand U19659 (N_19659,N_18698,N_18818);
xor U19660 (N_19660,N_18431,N_18471);
nand U19661 (N_19661,N_18406,N_18038);
nand U19662 (N_19662,N_18986,N_19082);
nor U19663 (N_19663,N_18760,N_18320);
nor U19664 (N_19664,N_18232,N_18881);
nor U19665 (N_19665,N_18813,N_18331);
and U19666 (N_19666,N_18255,N_18641);
nand U19667 (N_19667,N_18325,N_18651);
and U19668 (N_19668,N_18909,N_18717);
nor U19669 (N_19669,N_18639,N_19047);
or U19670 (N_19670,N_18900,N_18308);
or U19671 (N_19671,N_19183,N_18071);
or U19672 (N_19672,N_18898,N_19147);
nand U19673 (N_19673,N_18816,N_18960);
or U19674 (N_19674,N_18844,N_19115);
xor U19675 (N_19675,N_18969,N_18837);
nand U19676 (N_19676,N_18081,N_18128);
xor U19677 (N_19677,N_19182,N_18738);
xnor U19678 (N_19678,N_18810,N_18401);
xnor U19679 (N_19679,N_18031,N_18858);
or U19680 (N_19680,N_18107,N_18841);
nand U19681 (N_19681,N_18941,N_18498);
and U19682 (N_19682,N_18998,N_18494);
or U19683 (N_19683,N_18526,N_18714);
nor U19684 (N_19684,N_18236,N_18476);
nand U19685 (N_19685,N_18088,N_18319);
and U19686 (N_19686,N_19085,N_18429);
nor U19687 (N_19687,N_18701,N_18353);
nor U19688 (N_19688,N_19010,N_19070);
or U19689 (N_19689,N_18052,N_18105);
nand U19690 (N_19690,N_18677,N_18039);
or U19691 (N_19691,N_18938,N_18913);
or U19692 (N_19692,N_18158,N_19075);
nand U19693 (N_19693,N_19175,N_18534);
nand U19694 (N_19694,N_18778,N_18506);
or U19695 (N_19695,N_18274,N_18456);
or U19696 (N_19696,N_19003,N_18767);
or U19697 (N_19697,N_18376,N_18317);
or U19698 (N_19698,N_18421,N_18545);
nand U19699 (N_19699,N_18673,N_18194);
nand U19700 (N_19700,N_18195,N_18832);
and U19701 (N_19701,N_18366,N_18862);
nand U19702 (N_19702,N_19031,N_18553);
and U19703 (N_19703,N_18980,N_18855);
or U19704 (N_19704,N_18515,N_18905);
nor U19705 (N_19705,N_18789,N_18439);
and U19706 (N_19706,N_18332,N_18994);
or U19707 (N_19707,N_18956,N_18411);
nor U19708 (N_19708,N_18405,N_18511);
xor U19709 (N_19709,N_18187,N_18878);
nand U19710 (N_19710,N_18044,N_18369);
xor U19711 (N_19711,N_18021,N_18561);
or U19712 (N_19712,N_18389,N_18184);
nor U19713 (N_19713,N_18517,N_18636);
nand U19714 (N_19714,N_18329,N_18385);
xnor U19715 (N_19715,N_18585,N_18852);
nor U19716 (N_19716,N_18010,N_19112);
nand U19717 (N_19717,N_18759,N_19155);
and U19718 (N_19718,N_18499,N_18234);
nor U19719 (N_19719,N_18363,N_18749);
nor U19720 (N_19720,N_18289,N_18470);
and U19721 (N_19721,N_18987,N_19152);
nor U19722 (N_19722,N_18612,N_18416);
nand U19723 (N_19723,N_18480,N_18374);
nor U19724 (N_19724,N_19151,N_19157);
xor U19725 (N_19725,N_18575,N_19042);
nor U19726 (N_19726,N_18181,N_18718);
nand U19727 (N_19727,N_18155,N_18715);
and U19728 (N_19728,N_18356,N_18765);
nor U19729 (N_19729,N_18110,N_19097);
xor U19730 (N_19730,N_19058,N_18089);
nor U19731 (N_19731,N_18152,N_18453);
or U19732 (N_19732,N_19117,N_19161);
or U19733 (N_19733,N_18679,N_18877);
xnor U19734 (N_19734,N_18019,N_18700);
or U19735 (N_19735,N_18172,N_19084);
and U19736 (N_19736,N_18602,N_18048);
nand U19737 (N_19737,N_18732,N_18151);
nand U19738 (N_19738,N_19187,N_18551);
nor U19739 (N_19739,N_18473,N_18452);
xor U19740 (N_19740,N_19014,N_19124);
nand U19741 (N_19741,N_18399,N_18880);
nor U19742 (N_19742,N_19054,N_18896);
and U19743 (N_19743,N_18119,N_18665);
nor U19744 (N_19744,N_18090,N_18699);
xnor U19745 (N_19745,N_18352,N_19142);
xor U19746 (N_19746,N_18744,N_18180);
and U19747 (N_19747,N_18085,N_18224);
and U19748 (N_19748,N_18033,N_18901);
nand U19749 (N_19749,N_19130,N_18450);
xnor U19750 (N_19750,N_18166,N_18795);
and U19751 (N_19751,N_18915,N_18713);
nor U19752 (N_19752,N_18077,N_18126);
or U19753 (N_19753,N_18481,N_19002);
nand U19754 (N_19754,N_19104,N_19188);
or U19755 (N_19755,N_18359,N_19127);
and U19756 (N_19756,N_18762,N_18079);
or U19757 (N_19757,N_18262,N_18230);
nand U19758 (N_19758,N_18108,N_18235);
nor U19759 (N_19759,N_18931,N_18775);
nor U19760 (N_19760,N_19037,N_18891);
and U19761 (N_19761,N_18433,N_18384);
nor U19762 (N_19762,N_18016,N_18046);
xnor U19763 (N_19763,N_19179,N_18907);
or U19764 (N_19764,N_18756,N_18348);
nand U19765 (N_19765,N_18241,N_18231);
xor U19766 (N_19766,N_18906,N_18508);
xor U19767 (N_19767,N_18360,N_18124);
xnor U19768 (N_19768,N_19013,N_18594);
and U19769 (N_19769,N_18657,N_18563);
and U19770 (N_19770,N_18676,N_18556);
xnor U19771 (N_19771,N_18703,N_19171);
xor U19772 (N_19772,N_18104,N_19074);
nand U19773 (N_19773,N_18627,N_18580);
nand U19774 (N_19774,N_18072,N_18243);
nor U19775 (N_19775,N_18827,N_19172);
nor U19776 (N_19776,N_18216,N_18215);
nor U19777 (N_19777,N_18214,N_18623);
and U19778 (N_19778,N_18093,N_18351);
or U19779 (N_19779,N_18693,N_18613);
nand U19780 (N_19780,N_18574,N_18728);
and U19781 (N_19781,N_18326,N_19129);
xnor U19782 (N_19782,N_18769,N_18605);
nor U19783 (N_19783,N_18591,N_18949);
nand U19784 (N_19784,N_18294,N_18513);
nand U19785 (N_19785,N_18507,N_18393);
nand U19786 (N_19786,N_18434,N_18153);
or U19787 (N_19787,N_18776,N_18742);
and U19788 (N_19788,N_18402,N_18425);
or U19789 (N_19789,N_18041,N_19125);
and U19790 (N_19790,N_18619,N_18546);
nor U19791 (N_19791,N_18981,N_18740);
nor U19792 (N_19792,N_18060,N_19197);
or U19793 (N_19793,N_18003,N_18721);
xor U19794 (N_19794,N_18140,N_18062);
and U19795 (N_19795,N_18607,N_18503);
and U19796 (N_19796,N_18811,N_18323);
or U19797 (N_19797,N_18275,N_18295);
and U19798 (N_19798,N_18726,N_18669);
nor U19799 (N_19799,N_18787,N_18630);
nor U19800 (N_19800,N_18952,N_18445);
nand U19801 (N_19801,N_18353,N_18523);
nand U19802 (N_19802,N_18163,N_19063);
or U19803 (N_19803,N_19073,N_18021);
and U19804 (N_19804,N_19084,N_18992);
or U19805 (N_19805,N_18108,N_18845);
nor U19806 (N_19806,N_18232,N_18810);
or U19807 (N_19807,N_19050,N_18266);
nor U19808 (N_19808,N_18511,N_18177);
nor U19809 (N_19809,N_18947,N_18674);
xnor U19810 (N_19810,N_18059,N_19092);
or U19811 (N_19811,N_18339,N_18802);
xnor U19812 (N_19812,N_18168,N_18873);
or U19813 (N_19813,N_18770,N_18942);
xor U19814 (N_19814,N_18216,N_18314);
xor U19815 (N_19815,N_18341,N_19087);
nor U19816 (N_19816,N_18600,N_18496);
xnor U19817 (N_19817,N_18244,N_18299);
or U19818 (N_19818,N_18998,N_18290);
nor U19819 (N_19819,N_18100,N_18553);
xor U19820 (N_19820,N_18354,N_19132);
and U19821 (N_19821,N_19134,N_18619);
nor U19822 (N_19822,N_18678,N_18371);
nand U19823 (N_19823,N_18135,N_18625);
xor U19824 (N_19824,N_18881,N_18272);
nand U19825 (N_19825,N_18204,N_18893);
or U19826 (N_19826,N_18775,N_18237);
and U19827 (N_19827,N_19073,N_18787);
and U19828 (N_19828,N_18498,N_18729);
or U19829 (N_19829,N_18195,N_18301);
nand U19830 (N_19830,N_18200,N_18957);
nor U19831 (N_19831,N_18597,N_18974);
xnor U19832 (N_19832,N_18747,N_19047);
xnor U19833 (N_19833,N_18869,N_18250);
and U19834 (N_19834,N_18735,N_18754);
and U19835 (N_19835,N_19060,N_18494);
or U19836 (N_19836,N_18463,N_18024);
or U19837 (N_19837,N_19163,N_18082);
xnor U19838 (N_19838,N_18401,N_18021);
or U19839 (N_19839,N_18030,N_18893);
and U19840 (N_19840,N_18703,N_18167);
and U19841 (N_19841,N_18015,N_18628);
xnor U19842 (N_19842,N_19084,N_18150);
nor U19843 (N_19843,N_19004,N_19183);
or U19844 (N_19844,N_18220,N_18510);
and U19845 (N_19845,N_18538,N_18220);
xnor U19846 (N_19846,N_18610,N_18184);
nor U19847 (N_19847,N_18921,N_18514);
or U19848 (N_19848,N_18840,N_19170);
and U19849 (N_19849,N_18433,N_18147);
nand U19850 (N_19850,N_18182,N_18032);
xnor U19851 (N_19851,N_18421,N_18438);
nand U19852 (N_19852,N_19147,N_18952);
or U19853 (N_19853,N_18367,N_18105);
nor U19854 (N_19854,N_18898,N_18588);
nor U19855 (N_19855,N_18014,N_18146);
nand U19856 (N_19856,N_18178,N_18304);
and U19857 (N_19857,N_18509,N_18014);
xor U19858 (N_19858,N_19011,N_18124);
nor U19859 (N_19859,N_19145,N_18865);
nor U19860 (N_19860,N_18419,N_18258);
nor U19861 (N_19861,N_18758,N_18025);
nor U19862 (N_19862,N_18182,N_18153);
or U19863 (N_19863,N_18871,N_18064);
xor U19864 (N_19864,N_18733,N_18725);
nand U19865 (N_19865,N_18832,N_18407);
nand U19866 (N_19866,N_18911,N_18914);
or U19867 (N_19867,N_19170,N_18563);
nor U19868 (N_19868,N_18057,N_18767);
nor U19869 (N_19869,N_18565,N_18925);
xnor U19870 (N_19870,N_18899,N_18771);
and U19871 (N_19871,N_19183,N_18010);
xor U19872 (N_19872,N_18913,N_18922);
xor U19873 (N_19873,N_18353,N_19128);
nor U19874 (N_19874,N_18553,N_18185);
or U19875 (N_19875,N_18486,N_18566);
and U19876 (N_19876,N_18403,N_18087);
or U19877 (N_19877,N_18989,N_19091);
nand U19878 (N_19878,N_18764,N_18036);
or U19879 (N_19879,N_18805,N_18520);
nand U19880 (N_19880,N_18493,N_18243);
nand U19881 (N_19881,N_18525,N_18274);
nand U19882 (N_19882,N_18467,N_18532);
and U19883 (N_19883,N_18441,N_18365);
nand U19884 (N_19884,N_18050,N_18638);
xnor U19885 (N_19885,N_19193,N_18619);
xnor U19886 (N_19886,N_18672,N_18410);
xnor U19887 (N_19887,N_18636,N_18256);
xor U19888 (N_19888,N_19032,N_18435);
or U19889 (N_19889,N_18055,N_18196);
xor U19890 (N_19890,N_19114,N_18535);
nand U19891 (N_19891,N_18649,N_18522);
and U19892 (N_19892,N_18355,N_18368);
and U19893 (N_19893,N_18705,N_18992);
xor U19894 (N_19894,N_18449,N_18440);
and U19895 (N_19895,N_19020,N_18601);
and U19896 (N_19896,N_18272,N_18215);
nand U19897 (N_19897,N_18886,N_18910);
xnor U19898 (N_19898,N_18124,N_19183);
xor U19899 (N_19899,N_18888,N_19136);
nand U19900 (N_19900,N_18857,N_18840);
nand U19901 (N_19901,N_18170,N_18342);
or U19902 (N_19902,N_19142,N_18158);
and U19903 (N_19903,N_18979,N_18398);
xnor U19904 (N_19904,N_18700,N_18787);
or U19905 (N_19905,N_18389,N_18518);
nor U19906 (N_19906,N_18923,N_18960);
nand U19907 (N_19907,N_18993,N_19160);
xor U19908 (N_19908,N_18092,N_18003);
nand U19909 (N_19909,N_18482,N_18923);
and U19910 (N_19910,N_18119,N_18961);
and U19911 (N_19911,N_18176,N_18237);
nand U19912 (N_19912,N_18042,N_18498);
xor U19913 (N_19913,N_18150,N_18100);
or U19914 (N_19914,N_18289,N_18321);
nor U19915 (N_19915,N_18350,N_18049);
and U19916 (N_19916,N_18958,N_18511);
or U19917 (N_19917,N_18108,N_19169);
and U19918 (N_19918,N_18121,N_18903);
and U19919 (N_19919,N_18889,N_18210);
or U19920 (N_19920,N_18501,N_18910);
nor U19921 (N_19921,N_18013,N_18875);
nor U19922 (N_19922,N_18544,N_18219);
and U19923 (N_19923,N_18687,N_18617);
nor U19924 (N_19924,N_18992,N_18728);
and U19925 (N_19925,N_19189,N_19130);
nor U19926 (N_19926,N_19129,N_18997);
and U19927 (N_19927,N_19189,N_18269);
nor U19928 (N_19928,N_18775,N_18851);
and U19929 (N_19929,N_18734,N_18419);
and U19930 (N_19930,N_18108,N_18720);
and U19931 (N_19931,N_18833,N_18243);
and U19932 (N_19932,N_18618,N_18549);
nor U19933 (N_19933,N_18462,N_18530);
nand U19934 (N_19934,N_18859,N_18255);
xor U19935 (N_19935,N_18274,N_19117);
xnor U19936 (N_19936,N_18531,N_18880);
and U19937 (N_19937,N_18166,N_18658);
and U19938 (N_19938,N_18259,N_18173);
xnor U19939 (N_19939,N_19059,N_18676);
xor U19940 (N_19940,N_18884,N_18879);
and U19941 (N_19941,N_18682,N_18522);
nand U19942 (N_19942,N_18790,N_18997);
nand U19943 (N_19943,N_18508,N_18546);
or U19944 (N_19944,N_19093,N_19011);
nor U19945 (N_19945,N_18520,N_18290);
or U19946 (N_19946,N_18440,N_18175);
nand U19947 (N_19947,N_18866,N_19040);
nor U19948 (N_19948,N_18137,N_18092);
nand U19949 (N_19949,N_18002,N_18816);
nor U19950 (N_19950,N_18930,N_18495);
nor U19951 (N_19951,N_18945,N_18614);
nor U19952 (N_19952,N_19066,N_19093);
xor U19953 (N_19953,N_18633,N_18092);
and U19954 (N_19954,N_18239,N_18854);
nand U19955 (N_19955,N_18982,N_18056);
or U19956 (N_19956,N_19174,N_18413);
or U19957 (N_19957,N_18403,N_19190);
and U19958 (N_19958,N_18104,N_18565);
xnor U19959 (N_19959,N_18990,N_19114);
and U19960 (N_19960,N_18125,N_18696);
or U19961 (N_19961,N_19103,N_19040);
nor U19962 (N_19962,N_18000,N_18511);
or U19963 (N_19963,N_19019,N_18048);
or U19964 (N_19964,N_18763,N_18458);
nand U19965 (N_19965,N_18306,N_18862);
and U19966 (N_19966,N_19179,N_18256);
nand U19967 (N_19967,N_18829,N_19114);
and U19968 (N_19968,N_18468,N_18905);
nand U19969 (N_19969,N_18096,N_18597);
or U19970 (N_19970,N_18372,N_18590);
or U19971 (N_19971,N_18106,N_18980);
and U19972 (N_19972,N_18810,N_18372);
nor U19973 (N_19973,N_18017,N_18619);
nor U19974 (N_19974,N_18861,N_18930);
nand U19975 (N_19975,N_18750,N_18820);
nand U19976 (N_19976,N_18531,N_18476);
nor U19977 (N_19977,N_18088,N_18922);
nand U19978 (N_19978,N_18113,N_18225);
nor U19979 (N_19979,N_18835,N_19181);
nand U19980 (N_19980,N_18266,N_19157);
nand U19981 (N_19981,N_18892,N_19005);
nor U19982 (N_19982,N_18086,N_18250);
and U19983 (N_19983,N_18151,N_18261);
and U19984 (N_19984,N_19017,N_18555);
nor U19985 (N_19985,N_18494,N_18931);
xor U19986 (N_19986,N_18909,N_18036);
or U19987 (N_19987,N_18693,N_18628);
nand U19988 (N_19988,N_18688,N_18449);
xnor U19989 (N_19989,N_18979,N_18565);
nand U19990 (N_19990,N_18247,N_19156);
xor U19991 (N_19991,N_18512,N_18700);
xnor U19992 (N_19992,N_18022,N_18797);
nand U19993 (N_19993,N_18180,N_18681);
nand U19994 (N_19994,N_18055,N_18378);
nor U19995 (N_19995,N_18448,N_18482);
xor U19996 (N_19996,N_18599,N_19098);
and U19997 (N_19997,N_18231,N_19126);
xor U19998 (N_19998,N_18819,N_18472);
nand U19999 (N_19999,N_18526,N_18399);
and U20000 (N_20000,N_19126,N_18181);
and U20001 (N_20001,N_18545,N_18985);
nand U20002 (N_20002,N_18884,N_18438);
nand U20003 (N_20003,N_18484,N_18298);
and U20004 (N_20004,N_18011,N_18762);
and U20005 (N_20005,N_18024,N_18186);
or U20006 (N_20006,N_18804,N_19111);
nand U20007 (N_20007,N_18076,N_19071);
nor U20008 (N_20008,N_18046,N_18279);
and U20009 (N_20009,N_19174,N_18490);
or U20010 (N_20010,N_18303,N_18564);
xor U20011 (N_20011,N_18072,N_18151);
nand U20012 (N_20012,N_18578,N_18137);
nand U20013 (N_20013,N_18986,N_18935);
xor U20014 (N_20014,N_19124,N_19059);
and U20015 (N_20015,N_18622,N_18891);
xor U20016 (N_20016,N_18708,N_19037);
nand U20017 (N_20017,N_18528,N_18442);
nand U20018 (N_20018,N_19062,N_18830);
nand U20019 (N_20019,N_19114,N_18649);
nand U20020 (N_20020,N_19103,N_18136);
xnor U20021 (N_20021,N_19163,N_19188);
or U20022 (N_20022,N_18678,N_18388);
nand U20023 (N_20023,N_19150,N_18713);
and U20024 (N_20024,N_18181,N_18427);
and U20025 (N_20025,N_18242,N_18929);
and U20026 (N_20026,N_18561,N_18282);
nor U20027 (N_20027,N_18189,N_19016);
xor U20028 (N_20028,N_18440,N_18358);
nand U20029 (N_20029,N_18990,N_19094);
and U20030 (N_20030,N_18395,N_18656);
nor U20031 (N_20031,N_18624,N_18856);
nand U20032 (N_20032,N_18218,N_18029);
and U20033 (N_20033,N_18194,N_19034);
or U20034 (N_20034,N_18112,N_18424);
xor U20035 (N_20035,N_18609,N_19116);
nor U20036 (N_20036,N_18887,N_19188);
and U20037 (N_20037,N_18495,N_19049);
or U20038 (N_20038,N_18487,N_18849);
nor U20039 (N_20039,N_18093,N_18287);
nor U20040 (N_20040,N_18422,N_19107);
nand U20041 (N_20041,N_19066,N_18300);
or U20042 (N_20042,N_18886,N_18316);
nor U20043 (N_20043,N_19134,N_18224);
nor U20044 (N_20044,N_18045,N_18789);
nand U20045 (N_20045,N_18211,N_18663);
nor U20046 (N_20046,N_19123,N_19089);
and U20047 (N_20047,N_19155,N_19104);
nand U20048 (N_20048,N_18321,N_18166);
or U20049 (N_20049,N_18721,N_18233);
nand U20050 (N_20050,N_19050,N_18089);
nor U20051 (N_20051,N_18863,N_18311);
or U20052 (N_20052,N_18620,N_18928);
or U20053 (N_20053,N_18389,N_18194);
xor U20054 (N_20054,N_18968,N_18979);
or U20055 (N_20055,N_19043,N_18906);
xor U20056 (N_20056,N_18121,N_18068);
nand U20057 (N_20057,N_18004,N_19080);
or U20058 (N_20058,N_18856,N_18261);
or U20059 (N_20059,N_18287,N_18094);
and U20060 (N_20060,N_18699,N_18715);
nor U20061 (N_20061,N_18315,N_18740);
or U20062 (N_20062,N_18798,N_18446);
xnor U20063 (N_20063,N_18832,N_18363);
and U20064 (N_20064,N_18369,N_18047);
xnor U20065 (N_20065,N_18064,N_18127);
nand U20066 (N_20066,N_18221,N_19129);
and U20067 (N_20067,N_18866,N_19004);
and U20068 (N_20068,N_18033,N_18005);
or U20069 (N_20069,N_18008,N_18266);
and U20070 (N_20070,N_18956,N_18682);
and U20071 (N_20071,N_18287,N_18162);
or U20072 (N_20072,N_18985,N_19009);
xor U20073 (N_20073,N_18955,N_18525);
and U20074 (N_20074,N_18922,N_18034);
nor U20075 (N_20075,N_18253,N_18796);
or U20076 (N_20076,N_18999,N_18359);
or U20077 (N_20077,N_18783,N_18787);
nand U20078 (N_20078,N_18488,N_18612);
and U20079 (N_20079,N_18083,N_18101);
and U20080 (N_20080,N_18345,N_18671);
xor U20081 (N_20081,N_18019,N_18424);
nor U20082 (N_20082,N_18705,N_18140);
nor U20083 (N_20083,N_18171,N_18690);
nand U20084 (N_20084,N_18729,N_18573);
xor U20085 (N_20085,N_18126,N_18824);
nor U20086 (N_20086,N_18683,N_18604);
or U20087 (N_20087,N_18250,N_18381);
and U20088 (N_20088,N_18281,N_18866);
or U20089 (N_20089,N_18585,N_18341);
and U20090 (N_20090,N_18765,N_18647);
xor U20091 (N_20091,N_18865,N_18163);
and U20092 (N_20092,N_18602,N_19009);
or U20093 (N_20093,N_18531,N_19019);
nand U20094 (N_20094,N_18342,N_18809);
and U20095 (N_20095,N_18029,N_18062);
or U20096 (N_20096,N_18649,N_19095);
or U20097 (N_20097,N_18299,N_19086);
nand U20098 (N_20098,N_18739,N_18264);
and U20099 (N_20099,N_18008,N_18333);
xnor U20100 (N_20100,N_18647,N_18128);
or U20101 (N_20101,N_19080,N_18258);
xnor U20102 (N_20102,N_18046,N_18911);
and U20103 (N_20103,N_18778,N_18703);
nand U20104 (N_20104,N_18066,N_18797);
and U20105 (N_20105,N_18069,N_18402);
and U20106 (N_20106,N_18229,N_18721);
xnor U20107 (N_20107,N_18339,N_19160);
nand U20108 (N_20108,N_18379,N_19022);
nand U20109 (N_20109,N_18992,N_19053);
or U20110 (N_20110,N_18931,N_18381);
and U20111 (N_20111,N_18616,N_18176);
xor U20112 (N_20112,N_18612,N_18979);
nor U20113 (N_20113,N_18570,N_18485);
nor U20114 (N_20114,N_18787,N_18337);
xnor U20115 (N_20115,N_18103,N_18055);
or U20116 (N_20116,N_18401,N_18094);
nor U20117 (N_20117,N_18684,N_18514);
nor U20118 (N_20118,N_18234,N_18409);
xor U20119 (N_20119,N_18998,N_18186);
or U20120 (N_20120,N_18146,N_18711);
xor U20121 (N_20121,N_18520,N_18650);
nand U20122 (N_20122,N_18378,N_19078);
nor U20123 (N_20123,N_18954,N_18123);
nand U20124 (N_20124,N_19089,N_19147);
xnor U20125 (N_20125,N_19102,N_18514);
nand U20126 (N_20126,N_18525,N_18467);
or U20127 (N_20127,N_18161,N_18040);
or U20128 (N_20128,N_18785,N_18550);
nor U20129 (N_20129,N_18964,N_19151);
and U20130 (N_20130,N_18664,N_19120);
or U20131 (N_20131,N_19188,N_18110);
and U20132 (N_20132,N_18395,N_18905);
nor U20133 (N_20133,N_19074,N_18614);
nor U20134 (N_20134,N_19016,N_18052);
nor U20135 (N_20135,N_18707,N_18008);
xnor U20136 (N_20136,N_18125,N_18280);
nor U20137 (N_20137,N_18038,N_18659);
and U20138 (N_20138,N_18714,N_18825);
nor U20139 (N_20139,N_19078,N_18363);
nand U20140 (N_20140,N_18627,N_18008);
xor U20141 (N_20141,N_18068,N_18679);
nor U20142 (N_20142,N_18324,N_18856);
or U20143 (N_20143,N_18463,N_18816);
nor U20144 (N_20144,N_18173,N_18887);
xor U20145 (N_20145,N_19116,N_18714);
xnor U20146 (N_20146,N_18940,N_18153);
and U20147 (N_20147,N_18531,N_19122);
nor U20148 (N_20148,N_18775,N_18930);
or U20149 (N_20149,N_18935,N_18533);
nor U20150 (N_20150,N_18830,N_18337);
nor U20151 (N_20151,N_18340,N_18803);
nor U20152 (N_20152,N_18631,N_18277);
nor U20153 (N_20153,N_18504,N_18675);
nand U20154 (N_20154,N_18280,N_18052);
or U20155 (N_20155,N_18239,N_18913);
xor U20156 (N_20156,N_18558,N_18461);
or U20157 (N_20157,N_18294,N_19132);
or U20158 (N_20158,N_18322,N_18429);
xnor U20159 (N_20159,N_18933,N_18267);
or U20160 (N_20160,N_18214,N_18996);
or U20161 (N_20161,N_18270,N_19112);
xnor U20162 (N_20162,N_19173,N_18822);
nand U20163 (N_20163,N_18115,N_19099);
or U20164 (N_20164,N_19160,N_19161);
or U20165 (N_20165,N_18490,N_18692);
and U20166 (N_20166,N_19186,N_18000);
nand U20167 (N_20167,N_18151,N_18556);
and U20168 (N_20168,N_18850,N_18104);
nand U20169 (N_20169,N_18212,N_18287);
xor U20170 (N_20170,N_18099,N_19019);
nand U20171 (N_20171,N_19172,N_18037);
nor U20172 (N_20172,N_19131,N_18759);
nand U20173 (N_20173,N_18397,N_18548);
or U20174 (N_20174,N_18045,N_18374);
nor U20175 (N_20175,N_18409,N_18700);
or U20176 (N_20176,N_18681,N_18216);
or U20177 (N_20177,N_18653,N_18205);
and U20178 (N_20178,N_18755,N_18108);
nand U20179 (N_20179,N_18655,N_18038);
nor U20180 (N_20180,N_19171,N_18700);
xor U20181 (N_20181,N_18775,N_19136);
nand U20182 (N_20182,N_18791,N_19095);
and U20183 (N_20183,N_18107,N_18960);
or U20184 (N_20184,N_18330,N_19195);
and U20185 (N_20185,N_18452,N_18841);
xor U20186 (N_20186,N_19037,N_18058);
or U20187 (N_20187,N_19149,N_18590);
nand U20188 (N_20188,N_18000,N_19130);
nand U20189 (N_20189,N_18260,N_18852);
nand U20190 (N_20190,N_18621,N_19021);
xor U20191 (N_20191,N_18471,N_19190);
xor U20192 (N_20192,N_18290,N_18852);
nand U20193 (N_20193,N_18848,N_19116);
or U20194 (N_20194,N_18602,N_18311);
and U20195 (N_20195,N_18699,N_18042);
or U20196 (N_20196,N_18629,N_18778);
and U20197 (N_20197,N_18048,N_18872);
xnor U20198 (N_20198,N_18118,N_18145);
or U20199 (N_20199,N_18526,N_18691);
or U20200 (N_20200,N_18539,N_18854);
xnor U20201 (N_20201,N_19167,N_19199);
nor U20202 (N_20202,N_18514,N_18211);
nor U20203 (N_20203,N_18417,N_18472);
nor U20204 (N_20204,N_18667,N_18684);
xnor U20205 (N_20205,N_18093,N_18064);
nand U20206 (N_20206,N_18546,N_18992);
xor U20207 (N_20207,N_18849,N_18379);
nor U20208 (N_20208,N_18629,N_18649);
nor U20209 (N_20209,N_19123,N_18596);
nor U20210 (N_20210,N_18604,N_19070);
nor U20211 (N_20211,N_18765,N_18143);
and U20212 (N_20212,N_18931,N_18097);
nand U20213 (N_20213,N_19080,N_19077);
xor U20214 (N_20214,N_18007,N_18562);
or U20215 (N_20215,N_18118,N_18433);
nand U20216 (N_20216,N_19193,N_18782);
and U20217 (N_20217,N_18620,N_18883);
nand U20218 (N_20218,N_18774,N_18132);
nand U20219 (N_20219,N_18630,N_18531);
nand U20220 (N_20220,N_18487,N_18731);
nand U20221 (N_20221,N_19152,N_18595);
nand U20222 (N_20222,N_19128,N_18285);
nor U20223 (N_20223,N_18282,N_18122);
nand U20224 (N_20224,N_18749,N_18539);
nand U20225 (N_20225,N_18530,N_18303);
or U20226 (N_20226,N_18933,N_18377);
and U20227 (N_20227,N_18685,N_18956);
nand U20228 (N_20228,N_18378,N_18575);
nor U20229 (N_20229,N_18490,N_18252);
or U20230 (N_20230,N_19093,N_19143);
and U20231 (N_20231,N_18658,N_19134);
nand U20232 (N_20232,N_18215,N_18443);
nor U20233 (N_20233,N_18849,N_18396);
or U20234 (N_20234,N_18312,N_19025);
nand U20235 (N_20235,N_18281,N_18839);
or U20236 (N_20236,N_18260,N_18737);
or U20237 (N_20237,N_18153,N_18661);
nor U20238 (N_20238,N_18514,N_19147);
xor U20239 (N_20239,N_18276,N_18867);
or U20240 (N_20240,N_18198,N_18608);
and U20241 (N_20241,N_18689,N_18815);
and U20242 (N_20242,N_18102,N_18237);
and U20243 (N_20243,N_18246,N_18661);
nor U20244 (N_20244,N_18218,N_19110);
nand U20245 (N_20245,N_18911,N_18499);
xor U20246 (N_20246,N_18218,N_18628);
nor U20247 (N_20247,N_18649,N_18082);
or U20248 (N_20248,N_18614,N_18963);
or U20249 (N_20249,N_18214,N_18655);
or U20250 (N_20250,N_18985,N_19090);
nand U20251 (N_20251,N_18342,N_18110);
nor U20252 (N_20252,N_18266,N_19135);
or U20253 (N_20253,N_19007,N_18025);
and U20254 (N_20254,N_18033,N_18693);
nor U20255 (N_20255,N_18016,N_18846);
xor U20256 (N_20256,N_18206,N_19005);
nand U20257 (N_20257,N_18826,N_18380);
xnor U20258 (N_20258,N_18891,N_19038);
xnor U20259 (N_20259,N_18519,N_18748);
nand U20260 (N_20260,N_18994,N_18745);
xnor U20261 (N_20261,N_18802,N_18203);
xnor U20262 (N_20262,N_18998,N_18383);
nand U20263 (N_20263,N_19088,N_19170);
xor U20264 (N_20264,N_18930,N_18662);
or U20265 (N_20265,N_18639,N_18713);
nand U20266 (N_20266,N_18241,N_19004);
nor U20267 (N_20267,N_18811,N_19003);
xor U20268 (N_20268,N_18260,N_18919);
nand U20269 (N_20269,N_18171,N_19138);
nand U20270 (N_20270,N_18986,N_19060);
and U20271 (N_20271,N_18155,N_18878);
nor U20272 (N_20272,N_18551,N_19058);
nand U20273 (N_20273,N_18510,N_19098);
or U20274 (N_20274,N_18146,N_19152);
nand U20275 (N_20275,N_19159,N_19149);
xor U20276 (N_20276,N_18592,N_18161);
nor U20277 (N_20277,N_19043,N_19180);
nand U20278 (N_20278,N_18562,N_18737);
or U20279 (N_20279,N_19130,N_18104);
and U20280 (N_20280,N_18719,N_18108);
xor U20281 (N_20281,N_18633,N_18892);
nand U20282 (N_20282,N_18959,N_18759);
and U20283 (N_20283,N_18537,N_18208);
xor U20284 (N_20284,N_18135,N_18668);
nor U20285 (N_20285,N_18743,N_19187);
nor U20286 (N_20286,N_18295,N_19120);
nor U20287 (N_20287,N_19094,N_19091);
xnor U20288 (N_20288,N_18548,N_18358);
and U20289 (N_20289,N_19037,N_18706);
xor U20290 (N_20290,N_19008,N_18307);
nor U20291 (N_20291,N_18059,N_18573);
nor U20292 (N_20292,N_18978,N_18798);
xor U20293 (N_20293,N_18779,N_18864);
or U20294 (N_20294,N_18559,N_18094);
xnor U20295 (N_20295,N_18645,N_18786);
and U20296 (N_20296,N_18406,N_18464);
nand U20297 (N_20297,N_18587,N_18217);
and U20298 (N_20298,N_18410,N_18549);
and U20299 (N_20299,N_18592,N_18480);
nor U20300 (N_20300,N_18116,N_18060);
nand U20301 (N_20301,N_19038,N_18084);
or U20302 (N_20302,N_18786,N_18726);
or U20303 (N_20303,N_18890,N_18470);
nand U20304 (N_20304,N_19018,N_18755);
and U20305 (N_20305,N_18278,N_18480);
nand U20306 (N_20306,N_18724,N_18701);
and U20307 (N_20307,N_18332,N_18317);
nor U20308 (N_20308,N_18429,N_19097);
xnor U20309 (N_20309,N_18212,N_19044);
nor U20310 (N_20310,N_18479,N_18202);
xnor U20311 (N_20311,N_18241,N_18817);
xnor U20312 (N_20312,N_18678,N_18725);
nor U20313 (N_20313,N_18787,N_18446);
xnor U20314 (N_20314,N_18156,N_19120);
nor U20315 (N_20315,N_18307,N_19142);
nor U20316 (N_20316,N_18955,N_18960);
and U20317 (N_20317,N_18877,N_18968);
and U20318 (N_20318,N_18895,N_19034);
nor U20319 (N_20319,N_18565,N_18864);
nand U20320 (N_20320,N_19162,N_19045);
nand U20321 (N_20321,N_18415,N_18736);
and U20322 (N_20322,N_19160,N_18168);
or U20323 (N_20323,N_18784,N_18182);
or U20324 (N_20324,N_18503,N_18165);
xor U20325 (N_20325,N_18854,N_18229);
or U20326 (N_20326,N_18244,N_18819);
and U20327 (N_20327,N_18514,N_18101);
nor U20328 (N_20328,N_18102,N_18963);
nand U20329 (N_20329,N_19162,N_18570);
and U20330 (N_20330,N_18485,N_18904);
and U20331 (N_20331,N_19095,N_18740);
or U20332 (N_20332,N_18131,N_19175);
xor U20333 (N_20333,N_19027,N_18531);
xor U20334 (N_20334,N_18186,N_18373);
or U20335 (N_20335,N_18001,N_18386);
nor U20336 (N_20336,N_18632,N_18140);
or U20337 (N_20337,N_18889,N_18297);
and U20338 (N_20338,N_18274,N_18686);
xor U20339 (N_20339,N_18131,N_18708);
or U20340 (N_20340,N_18279,N_18063);
xnor U20341 (N_20341,N_18393,N_18232);
xnor U20342 (N_20342,N_18857,N_18202);
and U20343 (N_20343,N_18111,N_19001);
nor U20344 (N_20344,N_18621,N_18190);
or U20345 (N_20345,N_18729,N_18346);
nor U20346 (N_20346,N_18020,N_18837);
nand U20347 (N_20347,N_18362,N_18584);
or U20348 (N_20348,N_18683,N_18841);
xor U20349 (N_20349,N_19002,N_18754);
and U20350 (N_20350,N_18431,N_18985);
nand U20351 (N_20351,N_18575,N_18046);
and U20352 (N_20352,N_18605,N_18663);
and U20353 (N_20353,N_18704,N_18705);
and U20354 (N_20354,N_18495,N_18687);
nor U20355 (N_20355,N_18332,N_18930);
xnor U20356 (N_20356,N_18177,N_18017);
nor U20357 (N_20357,N_18478,N_18189);
xor U20358 (N_20358,N_18203,N_18944);
nand U20359 (N_20359,N_18058,N_18080);
nand U20360 (N_20360,N_18782,N_18684);
nand U20361 (N_20361,N_18352,N_18966);
nand U20362 (N_20362,N_18736,N_19001);
nand U20363 (N_20363,N_19186,N_19128);
nor U20364 (N_20364,N_18442,N_18674);
nor U20365 (N_20365,N_18458,N_18821);
or U20366 (N_20366,N_18323,N_18934);
nor U20367 (N_20367,N_18108,N_18335);
and U20368 (N_20368,N_18192,N_19035);
and U20369 (N_20369,N_18585,N_19182);
and U20370 (N_20370,N_19082,N_18121);
xor U20371 (N_20371,N_18390,N_19097);
nand U20372 (N_20372,N_18574,N_18122);
nor U20373 (N_20373,N_18710,N_18004);
nand U20374 (N_20374,N_18408,N_18742);
and U20375 (N_20375,N_18073,N_18685);
and U20376 (N_20376,N_18402,N_18730);
xnor U20377 (N_20377,N_18185,N_18509);
nand U20378 (N_20378,N_18091,N_18423);
nand U20379 (N_20379,N_18085,N_18288);
and U20380 (N_20380,N_18744,N_18838);
or U20381 (N_20381,N_18533,N_19018);
xor U20382 (N_20382,N_18393,N_18968);
or U20383 (N_20383,N_18669,N_18566);
nor U20384 (N_20384,N_19091,N_18510);
xor U20385 (N_20385,N_19147,N_18210);
nand U20386 (N_20386,N_18983,N_18598);
nand U20387 (N_20387,N_18237,N_18968);
nand U20388 (N_20388,N_18972,N_19122);
nand U20389 (N_20389,N_18371,N_18430);
xnor U20390 (N_20390,N_18458,N_18511);
xor U20391 (N_20391,N_18049,N_18999);
nor U20392 (N_20392,N_18638,N_18844);
or U20393 (N_20393,N_18899,N_18020);
xor U20394 (N_20394,N_18646,N_18246);
nor U20395 (N_20395,N_18302,N_19133);
xor U20396 (N_20396,N_18056,N_18205);
and U20397 (N_20397,N_19067,N_18683);
and U20398 (N_20398,N_18451,N_18090);
or U20399 (N_20399,N_19097,N_18296);
and U20400 (N_20400,N_19943,N_19227);
nand U20401 (N_20401,N_20267,N_19493);
and U20402 (N_20402,N_19257,N_20233);
nand U20403 (N_20403,N_20054,N_20129);
nand U20404 (N_20404,N_19276,N_19356);
xnor U20405 (N_20405,N_19357,N_20075);
xnor U20406 (N_20406,N_19427,N_19948);
xor U20407 (N_20407,N_20105,N_19919);
and U20408 (N_20408,N_19247,N_19502);
xor U20409 (N_20409,N_20310,N_20214);
or U20410 (N_20410,N_20254,N_19343);
and U20411 (N_20411,N_20038,N_20186);
nand U20412 (N_20412,N_19437,N_19882);
and U20413 (N_20413,N_20360,N_19658);
or U20414 (N_20414,N_20036,N_19536);
and U20415 (N_20415,N_19921,N_19679);
nand U20416 (N_20416,N_19593,N_19607);
nand U20417 (N_20417,N_19843,N_19232);
xnor U20418 (N_20418,N_19614,N_19602);
nor U20419 (N_20419,N_20340,N_19370);
or U20420 (N_20420,N_19916,N_19487);
nand U20421 (N_20421,N_20021,N_19307);
and U20422 (N_20422,N_20175,N_19692);
xnor U20423 (N_20423,N_20218,N_20355);
nor U20424 (N_20424,N_19443,N_19511);
nand U20425 (N_20425,N_19539,N_19394);
nor U20426 (N_20426,N_20224,N_19796);
and U20427 (N_20427,N_20270,N_19985);
and U20428 (N_20428,N_19258,N_19344);
nand U20429 (N_20429,N_19220,N_20101);
nand U20430 (N_20430,N_19832,N_19981);
nor U20431 (N_20431,N_19622,N_19219);
xnor U20432 (N_20432,N_19709,N_19317);
and U20433 (N_20433,N_20055,N_19619);
nor U20434 (N_20434,N_20091,N_19777);
or U20435 (N_20435,N_19830,N_20322);
xor U20436 (N_20436,N_19890,N_19996);
xor U20437 (N_20437,N_19668,N_20196);
nor U20438 (N_20438,N_19512,N_19503);
or U20439 (N_20439,N_19854,N_19953);
and U20440 (N_20440,N_19945,N_19620);
and U20441 (N_20441,N_20077,N_19407);
xor U20442 (N_20442,N_20093,N_20385);
or U20443 (N_20443,N_20000,N_19324);
and U20444 (N_20444,N_19972,N_19616);
xnor U20445 (N_20445,N_19974,N_20028);
and U20446 (N_20446,N_20380,N_20042);
nand U20447 (N_20447,N_19845,N_19809);
and U20448 (N_20448,N_19390,N_19630);
nand U20449 (N_20449,N_19995,N_20294);
xnor U20450 (N_20450,N_20122,N_19445);
or U20451 (N_20451,N_20159,N_19495);
nand U20452 (N_20452,N_20158,N_19413);
nor U20453 (N_20453,N_19705,N_19557);
and U20454 (N_20454,N_20389,N_19578);
nand U20455 (N_20455,N_20066,N_20127);
or U20456 (N_20456,N_20151,N_20229);
xor U20457 (N_20457,N_20349,N_20369);
nor U20458 (N_20458,N_19527,N_19310);
and U20459 (N_20459,N_19648,N_19775);
nand U20460 (N_20460,N_19449,N_19715);
nor U20461 (N_20461,N_19359,N_19336);
and U20462 (N_20462,N_20399,N_20307);
xor U20463 (N_20463,N_19788,N_19534);
or U20464 (N_20464,N_20298,N_20372);
and U20465 (N_20465,N_19636,N_19375);
nand U20466 (N_20466,N_20248,N_19200);
nand U20467 (N_20467,N_19711,N_19458);
or U20468 (N_20468,N_19713,N_20025);
nor U20469 (N_20469,N_19531,N_20020);
nand U20470 (N_20470,N_19421,N_20081);
nand U20471 (N_20471,N_19629,N_20098);
xnor U20472 (N_20472,N_20117,N_20219);
nor U20473 (N_20473,N_20222,N_20133);
xor U20474 (N_20474,N_19387,N_19889);
xnor U20475 (N_20475,N_19997,N_19723);
xor U20476 (N_20476,N_19254,N_19386);
xor U20477 (N_20477,N_20004,N_19484);
or U20478 (N_20478,N_19522,N_19934);
or U20479 (N_20479,N_20303,N_20246);
nor U20480 (N_20480,N_19561,N_20283);
nand U20481 (N_20481,N_20191,N_20276);
nand U20482 (N_20482,N_19416,N_19951);
or U20483 (N_20483,N_19291,N_19624);
xnor U20484 (N_20484,N_20162,N_19990);
and U20485 (N_20485,N_19391,N_19769);
nor U20486 (N_20486,N_19419,N_19682);
xnor U20487 (N_20487,N_20083,N_19385);
xnor U20488 (N_20488,N_19831,N_19499);
or U20489 (N_20489,N_19966,N_19929);
xnor U20490 (N_20490,N_19829,N_19450);
and U20491 (N_20491,N_19733,N_20046);
or U20492 (N_20492,N_20285,N_19982);
and U20493 (N_20493,N_20280,N_19672);
or U20494 (N_20494,N_19621,N_19861);
nor U20495 (N_20495,N_20286,N_20318);
xnor U20496 (N_20496,N_19615,N_20386);
xnor U20497 (N_20497,N_19700,N_19252);
xnor U20498 (N_20498,N_19609,N_20217);
nor U20499 (N_20499,N_19738,N_19563);
or U20500 (N_20500,N_19489,N_19970);
nand U20501 (N_20501,N_19737,N_20095);
xor U20502 (N_20502,N_19828,N_20250);
and U20503 (N_20503,N_19547,N_19497);
xnor U20504 (N_20504,N_20252,N_19286);
or U20505 (N_20505,N_19347,N_19538);
nor U20506 (N_20506,N_19496,N_19325);
nor U20507 (N_20507,N_20263,N_20266);
or U20508 (N_20508,N_19474,N_19920);
or U20509 (N_20509,N_19873,N_19428);
xor U20510 (N_20510,N_19400,N_19261);
xor U20511 (N_20511,N_19752,N_20144);
xnor U20512 (N_20512,N_20064,N_19786);
nand U20513 (N_20513,N_20113,N_19817);
and U20514 (N_20514,N_19410,N_20211);
nor U20515 (N_20515,N_20199,N_19521);
or U20516 (N_20516,N_19922,N_19839);
and U20517 (N_20517,N_19305,N_19653);
nand U20518 (N_20518,N_20381,N_19568);
nand U20519 (N_20519,N_20333,N_20163);
and U20520 (N_20520,N_19902,N_19936);
nor U20521 (N_20521,N_19265,N_19859);
and U20522 (N_20522,N_20157,N_19438);
nor U20523 (N_20523,N_19627,N_20154);
nand U20524 (N_20524,N_19581,N_19288);
or U20525 (N_20525,N_19423,N_19867);
xnor U20526 (N_20526,N_19248,N_19710);
nand U20527 (N_20527,N_19467,N_19403);
and U20528 (N_20528,N_19411,N_19454);
nand U20529 (N_20529,N_19937,N_19562);
nor U20530 (N_20530,N_20301,N_20176);
xor U20531 (N_20531,N_20178,N_19430);
nor U20532 (N_20532,N_19743,N_19695);
nand U20533 (N_20533,N_20051,N_19909);
xor U20534 (N_20534,N_19482,N_19354);
or U20535 (N_20535,N_20183,N_19941);
or U20536 (N_20536,N_19281,N_20257);
or U20537 (N_20537,N_20092,N_19456);
xnor U20538 (N_20538,N_19514,N_19631);
xor U20539 (N_20539,N_19967,N_19510);
or U20540 (N_20540,N_19462,N_20226);
nand U20541 (N_20541,N_19857,N_20053);
or U20542 (N_20542,N_20264,N_19238);
and U20543 (N_20543,N_19623,N_20079);
nand U20544 (N_20544,N_20330,N_20114);
nand U20545 (N_20545,N_19575,N_20203);
nand U20546 (N_20546,N_20164,N_19923);
nor U20547 (N_20547,N_20378,N_20251);
nand U20548 (N_20548,N_19225,N_19481);
or U20549 (N_20549,N_19478,N_19924);
nand U20550 (N_20550,N_19712,N_19825);
nor U20551 (N_20551,N_19224,N_20040);
or U20552 (N_20552,N_19422,N_19349);
or U20553 (N_20553,N_19960,N_20261);
xor U20554 (N_20554,N_20361,N_19681);
xnor U20555 (N_20555,N_19698,N_19202);
xor U20556 (N_20556,N_19229,N_20209);
nor U20557 (N_20557,N_20287,N_20230);
nor U20558 (N_20558,N_20106,N_20321);
or U20559 (N_20559,N_20259,N_20135);
and U20560 (N_20560,N_19442,N_20011);
nor U20561 (N_20561,N_19841,N_19840);
and U20562 (N_20562,N_19911,N_19472);
nor U20563 (N_20563,N_19954,N_19611);
or U20564 (N_20564,N_19315,N_20236);
nand U20565 (N_20565,N_19803,N_20161);
nor U20566 (N_20566,N_19235,N_20029);
nand U20567 (N_20567,N_19676,N_20047);
or U20568 (N_20568,N_19498,N_19504);
xor U20569 (N_20569,N_20234,N_20205);
nor U20570 (N_20570,N_20018,N_20136);
nor U20571 (N_20571,N_19935,N_19714);
or U20572 (N_20572,N_19983,N_20168);
xnor U20573 (N_20573,N_20060,N_19644);
or U20574 (N_20574,N_19665,N_20078);
and U20575 (N_20575,N_19880,N_19452);
and U20576 (N_20576,N_19598,N_20245);
nor U20577 (N_20577,N_20160,N_20323);
or U20578 (N_20578,N_19309,N_20185);
nor U20579 (N_20579,N_19515,N_20056);
or U20580 (N_20580,N_19677,N_19938);
or U20581 (N_20581,N_20034,N_20352);
nand U20582 (N_20582,N_20271,N_19519);
xor U20583 (N_20583,N_19824,N_20353);
nor U20584 (N_20584,N_19260,N_20367);
and U20585 (N_20585,N_20174,N_19654);
nand U20586 (N_20586,N_19206,N_19275);
nand U20587 (N_20587,N_19290,N_19747);
nand U20588 (N_20588,N_19469,N_19740);
nor U20589 (N_20589,N_19213,N_19696);
nand U20590 (N_20590,N_19708,N_19780);
xor U20591 (N_20591,N_19204,N_20304);
or U20592 (N_20592,N_19520,N_19337);
and U20593 (N_20593,N_19564,N_20290);
nor U20594 (N_20594,N_19264,N_20341);
nor U20595 (N_20595,N_19486,N_19603);
or U20596 (N_20596,N_19331,N_20273);
and U20597 (N_20597,N_19551,N_19548);
and U20598 (N_20598,N_20071,N_19781);
xor U20599 (N_20599,N_20343,N_20024);
nand U20600 (N_20600,N_19353,N_19274);
nor U20601 (N_20601,N_19931,N_19362);
nor U20602 (N_20602,N_19580,N_20103);
nand U20603 (N_20603,N_20096,N_19569);
nand U20604 (N_20604,N_19772,N_19397);
nor U20605 (N_20605,N_20379,N_20317);
nor U20606 (N_20606,N_19699,N_19640);
nand U20607 (N_20607,N_19874,N_19998);
nand U20608 (N_20608,N_19552,N_19932);
nor U20609 (N_20609,N_20382,N_20215);
xor U20610 (N_20610,N_19372,N_20086);
or U20611 (N_20611,N_19457,N_19366);
xor U20612 (N_20612,N_20324,N_19540);
or U20613 (N_20613,N_19476,N_19312);
or U20614 (N_20614,N_20244,N_19283);
xor U20615 (N_20615,N_19374,N_19446);
nand U20616 (N_20616,N_19858,N_19451);
xnor U20617 (N_20617,N_19673,N_19688);
and U20618 (N_20618,N_19866,N_20313);
or U20619 (N_20619,N_19808,N_19214);
nor U20620 (N_20620,N_19759,N_19358);
and U20621 (N_20621,N_20049,N_20362);
nand U20622 (N_20622,N_20019,N_20084);
or U20623 (N_20623,N_19895,N_19739);
or U20624 (N_20624,N_20366,N_20088);
xnor U20625 (N_20625,N_20013,N_19693);
or U20626 (N_20626,N_19761,N_19546);
or U20627 (N_20627,N_19933,N_19968);
nand U20628 (N_20628,N_19234,N_20332);
nor U20629 (N_20629,N_19279,N_20210);
or U20630 (N_20630,N_19987,N_20147);
nor U20631 (N_20631,N_19961,N_20044);
and U20632 (N_20632,N_19271,N_19466);
and U20633 (N_20633,N_19601,N_19787);
nand U20634 (N_20634,N_19877,N_19685);
and U20635 (N_20635,N_20311,N_20309);
or U20636 (N_20636,N_19392,N_20169);
xor U20637 (N_20637,N_19815,N_19844);
and U20638 (N_20638,N_19399,N_20354);
nor U20639 (N_20639,N_20134,N_20110);
xnor U20640 (N_20640,N_19577,N_20282);
xnor U20641 (N_20641,N_19718,N_19952);
xor U20642 (N_20642,N_19304,N_19251);
nor U20643 (N_20643,N_20239,N_19683);
or U20644 (N_20644,N_19804,N_19471);
or U20645 (N_20645,N_19383,N_20177);
or U20646 (N_20646,N_19748,N_19605);
and U20647 (N_20647,N_19277,N_19595);
xor U20648 (N_20648,N_19453,N_19555);
or U20649 (N_20649,N_19298,N_19822);
nand U20650 (N_20650,N_20052,N_20202);
nand U20651 (N_20651,N_19986,N_20195);
nor U20652 (N_20652,N_19635,N_19460);
xnor U20653 (N_20653,N_19565,N_20278);
or U20654 (N_20654,N_19907,N_19662);
or U20655 (N_20655,N_19240,N_19228);
nor U20656 (N_20656,N_19364,N_19367);
xnor U20657 (N_20657,N_19612,N_20231);
nand U20658 (N_20658,N_19899,N_19342);
and U20659 (N_20659,N_19613,N_20281);
or U20660 (N_20660,N_19826,N_20358);
nand U20661 (N_20661,N_19927,N_20089);
nor U20662 (N_20662,N_20291,N_19537);
xnor U20663 (N_20663,N_19402,N_19380);
xnor U20664 (N_20664,N_19618,N_20308);
or U20665 (N_20665,N_19862,N_19352);
or U20666 (N_20666,N_19517,N_20204);
or U20667 (N_20667,N_20145,N_19205);
xnor U20668 (N_20668,N_19282,N_20012);
and U20669 (N_20669,N_20082,N_19633);
nand U20670 (N_20670,N_19433,N_19939);
nand U20671 (N_20671,N_19868,N_20228);
or U20672 (N_20672,N_19638,N_19837);
nor U20673 (N_20673,N_19884,N_19384);
and U20674 (N_20674,N_19827,N_19914);
nand U20675 (N_20675,N_19295,N_20108);
or U20676 (N_20676,N_19355,N_19389);
nor U20677 (N_20677,N_19706,N_19691);
nor U20678 (N_20678,N_19323,N_19465);
nor U20679 (N_20679,N_20043,N_19860);
nand U20680 (N_20680,N_20058,N_19716);
nand U20681 (N_20681,N_20374,N_19795);
or U20682 (N_20682,N_19993,N_20201);
nand U20683 (N_20683,N_20100,N_19785);
and U20684 (N_20684,N_20015,N_19412);
or U20685 (N_20685,N_19838,N_20391);
or U20686 (N_20686,N_19221,N_20302);
and U20687 (N_20687,N_19382,N_19529);
xor U20688 (N_20688,N_19525,N_19915);
nand U20689 (N_20689,N_20395,N_19313);
or U20690 (N_20690,N_20260,N_19617);
xnor U20691 (N_20691,N_19984,N_20325);
or U20692 (N_20692,N_20027,N_20062);
xnor U20693 (N_20693,N_19946,N_19763);
or U20694 (N_20694,N_19925,N_20327);
nor U20695 (N_20695,N_19243,N_20388);
nor U20696 (N_20696,N_19209,N_19792);
xor U20697 (N_20697,N_20048,N_19294);
xnor U20698 (N_20698,N_19420,N_19244);
or U20699 (N_20699,N_20232,N_20335);
nand U20700 (N_20700,N_19226,N_19641);
xor U20701 (N_20701,N_19545,N_19401);
nor U20702 (N_20702,N_19724,N_20299);
xnor U20703 (N_20703,N_20009,N_19905);
nor U20704 (N_20704,N_20155,N_20397);
xor U20705 (N_20705,N_19249,N_19731);
xnor U20706 (N_20706,N_20387,N_19255);
or U20707 (N_20707,N_19208,N_20328);
or U20708 (N_20708,N_19550,N_19330);
xor U20709 (N_20709,N_20262,N_20139);
and U20710 (N_20710,N_19736,N_19798);
nand U20711 (N_20711,N_19814,N_20334);
and U20712 (N_20712,N_19216,N_20085);
nor U20713 (N_20713,N_19988,N_20141);
xor U20714 (N_20714,N_20193,N_19722);
nor U20715 (N_20715,N_20057,N_20272);
nor U20716 (N_20716,N_20293,N_20065);
nand U20717 (N_20717,N_20253,N_19599);
and U20718 (N_20718,N_20208,N_19944);
xor U20719 (N_20719,N_20140,N_19233);
nor U20720 (N_20720,N_19293,N_20045);
nor U20721 (N_20721,N_20143,N_20041);
nand U20722 (N_20722,N_20339,N_19892);
or U20723 (N_20723,N_19871,N_19878);
xnor U20724 (N_20724,N_20150,N_19346);
nand U20725 (N_20725,N_19758,N_19579);
xor U20726 (N_20726,N_19500,N_19376);
and U20727 (N_20727,N_19459,N_19774);
nand U20728 (N_20728,N_19897,N_19544);
xor U20729 (N_20729,N_19771,N_20316);
or U20730 (N_20730,N_19348,N_19339);
nor U20731 (N_20731,N_19746,N_19553);
and U20732 (N_20732,N_20375,N_19646);
xor U20733 (N_20733,N_19217,N_19405);
and U20734 (N_20734,N_19663,N_19797);
xnor U20735 (N_20735,N_19314,N_19231);
xnor U20736 (N_20736,N_20165,N_19778);
and U20737 (N_20737,N_20225,N_19686);
xnor U20738 (N_20738,N_19483,N_19779);
nand U20739 (N_20739,N_20120,N_19661);
nor U20740 (N_20740,N_19820,N_20347);
xor U20741 (N_20741,N_19721,N_19757);
xnor U20742 (N_20742,N_20300,N_19742);
or U20743 (N_20743,N_19373,N_19311);
or U20744 (N_20744,N_19628,N_19360);
and U20745 (N_20745,N_20297,N_19321);
nand U20746 (N_20746,N_19913,N_19856);
or U20747 (N_20747,N_19574,N_19791);
nand U20748 (N_20748,N_19490,N_19704);
xor U20749 (N_20749,N_20125,N_19879);
or U20750 (N_20750,N_19532,N_19992);
nand U20751 (N_20751,N_19643,N_19651);
nor U20752 (N_20752,N_20249,N_19729);
and U20753 (N_20753,N_19821,N_19765);
xnor U20754 (N_20754,N_20364,N_19908);
nor U20755 (N_20755,N_20398,N_19901);
nor U20756 (N_20756,N_20014,N_19678);
xnor U20757 (N_20757,N_20269,N_20173);
nor U20758 (N_20758,N_19414,N_19592);
or U20759 (N_20759,N_20390,N_20356);
and U20760 (N_20760,N_20296,N_20344);
nor U20761 (N_20761,N_19319,N_19789);
nand U20762 (N_20762,N_19659,N_19876);
or U20763 (N_20763,N_19211,N_19432);
nor U20764 (N_20764,N_19891,N_19223);
and U20765 (N_20765,N_19806,N_19583);
and U20766 (N_20766,N_19292,N_19448);
nor U20767 (N_20767,N_20132,N_19477);
nand U20768 (N_20768,N_19823,N_20138);
nor U20769 (N_20769,N_19872,N_19393);
nor U20770 (N_20770,N_20087,N_19381);
xor U20771 (N_20771,N_19964,N_19697);
nor U20772 (N_20772,N_20212,N_20109);
nand U20773 (N_20773,N_19671,N_19720);
and U20774 (N_20774,N_19894,N_19273);
xnor U20775 (N_20775,N_19299,N_20288);
nand U20776 (N_20776,N_20240,N_20142);
nand U20777 (N_20777,N_19239,N_19926);
nor U20778 (N_20778,N_19816,N_19530);
and U20779 (N_20779,N_19674,N_19201);
or U20780 (N_20780,N_19253,N_19980);
xor U20781 (N_20781,N_19215,N_19719);
and U20782 (N_20782,N_20166,N_19979);
or U20783 (N_20783,N_19567,N_20030);
xor U20784 (N_20784,N_20121,N_19689);
and U20785 (N_20785,N_19610,N_20094);
nand U20786 (N_20786,N_19218,N_19409);
xor U20787 (N_20787,N_19470,N_19368);
nor U20788 (N_20788,N_19764,N_19508);
or U20789 (N_20789,N_20119,N_20346);
and U20790 (N_20790,N_20050,N_19554);
and U20791 (N_20791,N_19755,N_20206);
and U20792 (N_20792,N_19756,N_19241);
or U20793 (N_20793,N_19694,N_20365);
nor U20794 (N_20794,N_19287,N_20111);
nand U20795 (N_20795,N_20104,N_19664);
nor U20796 (N_20796,N_20221,N_20123);
nor U20797 (N_20797,N_19904,N_19429);
and U20798 (N_20798,N_20067,N_20377);
or U20799 (N_20799,N_20006,N_20170);
or U20800 (N_20800,N_19475,N_19881);
xor U20801 (N_20801,N_19463,N_20396);
and U20802 (N_20802,N_20213,N_19975);
and U20803 (N_20803,N_19655,N_20080);
nor U20804 (N_20804,N_19702,N_19335);
or U20805 (N_20805,N_20235,N_19207);
or U20806 (N_20806,N_20200,N_19887);
nor U20807 (N_20807,N_20010,N_20180);
nor U20808 (N_20808,N_19851,N_20031);
xnor U20809 (N_20809,N_19263,N_19259);
nor U20810 (N_20810,N_20167,N_20072);
xnor U20811 (N_20811,N_19666,N_20116);
nor U20812 (N_20812,N_19363,N_20023);
nand U20813 (N_20813,N_20342,N_19268);
nand U20814 (N_20814,N_20189,N_19849);
or U20815 (N_20815,N_19505,N_19541);
or U20816 (N_20816,N_19917,N_20171);
and U20817 (N_20817,N_20350,N_19332);
nand U20818 (N_20818,N_19807,N_20295);
xnor U20819 (N_20819,N_19594,N_20258);
nand U20820 (N_20820,N_19800,N_19345);
or U20821 (N_20821,N_19833,N_19865);
nor U20822 (N_20822,N_19649,N_19918);
xor U20823 (N_20823,N_20005,N_19542);
or U20824 (N_20824,N_19669,N_20274);
nor U20825 (N_20825,N_19690,N_20265);
nand U20826 (N_20826,N_19883,N_19930);
or U20827 (N_20827,N_19371,N_19900);
xnor U20828 (N_20828,N_19435,N_19418);
or U20829 (N_20829,N_19464,N_19957);
xor U20830 (N_20830,N_19308,N_19888);
and U20831 (N_20831,N_19415,N_19770);
or U20832 (N_20832,N_19639,N_20351);
or U20833 (N_20833,N_20131,N_19794);
nor U20834 (N_20834,N_19842,N_19543);
xnor U20835 (N_20835,N_19745,N_19341);
xnor U20836 (N_20836,N_19625,N_20247);
or U20837 (N_20837,N_19242,N_20063);
xor U20838 (N_20838,N_19272,N_20194);
nand U20839 (N_20839,N_20130,N_20146);
and U20840 (N_20840,N_19994,N_20242);
and U20841 (N_20841,N_19398,N_19645);
xnor U20842 (N_20842,N_19289,N_19506);
nor U20843 (N_20843,N_19256,N_20376);
or U20844 (N_20844,N_19327,N_20070);
and U20845 (N_20845,N_19589,N_19439);
or U20846 (N_20846,N_19447,N_19766);
or U20847 (N_20847,N_19480,N_20188);
xnor U20848 (N_20848,N_20179,N_20182);
and U20849 (N_20849,N_19590,N_20068);
and U20850 (N_20850,N_20319,N_19810);
xor U20851 (N_20851,N_19834,N_19912);
nand U20852 (N_20852,N_19701,N_19657);
and U20853 (N_20853,N_19587,N_20112);
and U20854 (N_20854,N_19491,N_19212);
nor U20855 (N_20855,N_19378,N_19726);
nor U20856 (N_20856,N_19479,N_20149);
xnor U20857 (N_20857,N_19507,N_20115);
nand U20858 (N_20858,N_20284,N_20008);
or U20859 (N_20859,N_20007,N_19230);
and U20860 (N_20860,N_19431,N_19395);
or U20861 (N_20861,N_19846,N_19855);
nand U20862 (N_20862,N_20032,N_19976);
xnor U20863 (N_20863,N_19560,N_19513);
xor U20864 (N_20864,N_19991,N_20314);
and U20865 (N_20865,N_19535,N_20279);
or U20866 (N_20866,N_20359,N_19707);
and U20867 (N_20867,N_19734,N_20394);
and U20868 (N_20868,N_20102,N_19727);
and U20869 (N_20869,N_19969,N_19684);
xor U20870 (N_20870,N_19750,N_19494);
nor U20871 (N_20871,N_20255,N_19801);
nand U20872 (N_20872,N_19942,N_19528);
nand U20873 (N_20873,N_19338,N_20306);
xor U20874 (N_20874,N_19973,N_19455);
or U20875 (N_20875,N_19408,N_19893);
and U20876 (N_20876,N_19559,N_19351);
xnor U20877 (N_20877,N_20238,N_19642);
nor U20878 (N_20878,N_19526,N_19652);
and U20879 (N_20879,N_19572,N_19949);
xnor U20880 (N_20880,N_19776,N_20039);
and U20881 (N_20881,N_20148,N_20320);
and U20882 (N_20882,N_20035,N_20241);
nor U20883 (N_20883,N_19333,N_19903);
and U20884 (N_20884,N_20237,N_19269);
xor U20885 (N_20885,N_19863,N_19262);
nor U20886 (N_20886,N_19848,N_19285);
or U20887 (N_20887,N_19441,N_19571);
nor U20888 (N_20888,N_19637,N_19236);
nor U20889 (N_20889,N_19773,N_20118);
or U20890 (N_20890,N_19425,N_19524);
nor U20891 (N_20891,N_19284,N_19790);
xnor U20892 (N_20892,N_19647,N_19965);
nor U20893 (N_20893,N_19584,N_19805);
or U20894 (N_20894,N_19509,N_19989);
or U20895 (N_20895,N_19928,N_19434);
nor U20896 (N_20896,N_19328,N_20022);
nand U20897 (N_20897,N_19898,N_19793);
and U20898 (N_20898,N_20156,N_20393);
xor U20899 (N_20899,N_19818,N_20363);
or U20900 (N_20900,N_19799,N_19977);
nor U20901 (N_20901,N_20220,N_19753);
or U20902 (N_20902,N_19586,N_20016);
nand U20903 (N_20903,N_20370,N_19782);
xor U20904 (N_20904,N_19910,N_19573);
or U20905 (N_20905,N_19591,N_19847);
nor U20906 (N_20906,N_19300,N_20124);
or U20907 (N_20907,N_20315,N_19606);
nand U20908 (N_20908,N_19301,N_19852);
or U20909 (N_20909,N_19735,N_20277);
or U20910 (N_20910,N_19836,N_19426);
xor U20911 (N_20911,N_19516,N_19767);
xor U20912 (N_20912,N_20073,N_19361);
xnor U20913 (N_20913,N_19566,N_19501);
or U20914 (N_20914,N_20216,N_20037);
xor U20915 (N_20915,N_19303,N_19334);
nand U20916 (N_20916,N_19302,N_19340);
nand U20917 (N_20917,N_19875,N_20338);
xor U20918 (N_20918,N_19670,N_19296);
and U20919 (N_20919,N_20383,N_19885);
and U20920 (N_20920,N_19811,N_19377);
nand U20921 (N_20921,N_20373,N_19813);
nand U20922 (N_20922,N_19864,N_20292);
nor U20923 (N_20923,N_20268,N_20152);
nand U20924 (N_20924,N_19768,N_19582);
nand U20925 (N_20925,N_20026,N_19608);
nand U20926 (N_20926,N_19999,N_20184);
nor U20927 (N_20927,N_19237,N_20289);
xor U20928 (N_20928,N_20207,N_19963);
nand U20929 (N_20929,N_19436,N_20312);
nor U20930 (N_20930,N_19246,N_20003);
and U20931 (N_20931,N_19245,N_19906);
nand U20932 (N_20932,N_19667,N_20076);
xnor U20933 (N_20933,N_19958,N_19956);
or U20934 (N_20934,N_19869,N_19634);
nor U20935 (N_20935,N_19444,N_20090);
xnor U20936 (N_20936,N_19396,N_20001);
or U20937 (N_20937,N_19523,N_19556);
or U20938 (N_20938,N_20187,N_19728);
or U20939 (N_20939,N_19388,N_19576);
nor U20940 (N_20940,N_20128,N_20099);
and U20941 (N_20941,N_20033,N_20059);
nand U20942 (N_20942,N_19971,N_19492);
nor U20943 (N_20943,N_19597,N_20097);
and U20944 (N_20944,N_19297,N_19406);
nor U20945 (N_20945,N_20181,N_19626);
or U20946 (N_20946,N_20017,N_20074);
nor U20947 (N_20947,N_19404,N_20069);
nand U20948 (N_20948,N_20256,N_19379);
nor U20949 (N_20949,N_19488,N_19266);
or U20950 (N_20950,N_19680,N_19656);
or U20951 (N_20951,N_20275,N_19318);
and U20952 (N_20952,N_19326,N_19762);
nor U20953 (N_20953,N_20126,N_19675);
and U20954 (N_20954,N_19886,N_19417);
xnor U20955 (N_20955,N_19744,N_19660);
nor U20956 (N_20956,N_19650,N_19210);
nand U20957 (N_20957,N_19730,N_19604);
or U20958 (N_20958,N_20137,N_20305);
nand U20959 (N_20959,N_19250,N_19853);
or U20960 (N_20960,N_19760,N_20192);
and U20961 (N_20961,N_19585,N_20392);
or U20962 (N_20962,N_20331,N_19533);
nand U20963 (N_20963,N_19819,N_20329);
nand U20964 (N_20964,N_20357,N_19978);
nand U20965 (N_20965,N_20172,N_19725);
nand U20966 (N_20966,N_19812,N_20153);
nand U20967 (N_20967,N_20326,N_20371);
nand U20968 (N_20968,N_19322,N_19732);
nand U20969 (N_20969,N_19369,N_20198);
and U20970 (N_20970,N_19267,N_19588);
nand U20971 (N_20971,N_19870,N_19741);
xnor U20972 (N_20972,N_19440,N_19350);
nand U20973 (N_20973,N_20336,N_19947);
nand U20974 (N_20974,N_20348,N_19896);
xnor U20975 (N_20975,N_19802,N_20002);
or U20976 (N_20976,N_19203,N_20243);
xnor U20977 (N_20977,N_19329,N_19270);
nand U20978 (N_20978,N_19461,N_19280);
or U20979 (N_20979,N_20223,N_20061);
nand U20980 (N_20980,N_19717,N_19955);
nor U20981 (N_20981,N_20107,N_19278);
nor U20982 (N_20982,N_19365,N_19222);
and U20983 (N_20983,N_19320,N_19754);
and U20984 (N_20984,N_19783,N_19632);
xor U20985 (N_20985,N_20197,N_20368);
nand U20986 (N_20986,N_19940,N_20227);
and U20987 (N_20987,N_19570,N_19687);
nor U20988 (N_20988,N_19468,N_19518);
nand U20989 (N_20989,N_19316,N_20337);
or U20990 (N_20990,N_20384,N_19749);
or U20991 (N_20991,N_19703,N_19558);
and U20992 (N_20992,N_19473,N_19959);
and U20993 (N_20993,N_19485,N_19784);
and U20994 (N_20994,N_19950,N_19962);
or U20995 (N_20995,N_19600,N_19835);
xor U20996 (N_20996,N_19549,N_19850);
xor U20997 (N_20997,N_20190,N_19424);
nor U20998 (N_20998,N_19596,N_20345);
and U20999 (N_20999,N_19751,N_19306);
xnor U21000 (N_21000,N_19868,N_19226);
and U21001 (N_21001,N_19345,N_19371);
and U21002 (N_21002,N_20370,N_19555);
and U21003 (N_21003,N_19455,N_19216);
nor U21004 (N_21004,N_20039,N_19444);
or U21005 (N_21005,N_20167,N_20392);
nand U21006 (N_21006,N_20071,N_19269);
nor U21007 (N_21007,N_20080,N_20383);
nor U21008 (N_21008,N_19508,N_20252);
or U21009 (N_21009,N_20351,N_20233);
or U21010 (N_21010,N_20147,N_19655);
or U21011 (N_21011,N_20299,N_19892);
nor U21012 (N_21012,N_19476,N_19575);
and U21013 (N_21013,N_19664,N_19484);
or U21014 (N_21014,N_19477,N_19599);
xnor U21015 (N_21015,N_19731,N_20135);
or U21016 (N_21016,N_19857,N_19621);
and U21017 (N_21017,N_20170,N_19410);
nand U21018 (N_21018,N_19647,N_19480);
and U21019 (N_21019,N_19305,N_19375);
and U21020 (N_21020,N_20034,N_19949);
nand U21021 (N_21021,N_19411,N_20130);
or U21022 (N_21022,N_19541,N_19348);
or U21023 (N_21023,N_20016,N_19549);
or U21024 (N_21024,N_19950,N_20097);
nor U21025 (N_21025,N_19480,N_20363);
or U21026 (N_21026,N_19342,N_19916);
or U21027 (N_21027,N_19414,N_20208);
or U21028 (N_21028,N_19588,N_19602);
nor U21029 (N_21029,N_19521,N_20008);
or U21030 (N_21030,N_19625,N_20033);
xnor U21031 (N_21031,N_19614,N_20051);
or U21032 (N_21032,N_19707,N_20317);
or U21033 (N_21033,N_19411,N_19241);
nor U21034 (N_21034,N_20038,N_19367);
nor U21035 (N_21035,N_19562,N_19651);
nor U21036 (N_21036,N_19876,N_19325);
nand U21037 (N_21037,N_20204,N_19984);
and U21038 (N_21038,N_19403,N_20089);
nand U21039 (N_21039,N_19509,N_19976);
or U21040 (N_21040,N_20264,N_20000);
nand U21041 (N_21041,N_20340,N_20320);
xor U21042 (N_21042,N_20136,N_20373);
xor U21043 (N_21043,N_19246,N_19641);
nor U21044 (N_21044,N_20303,N_20235);
and U21045 (N_21045,N_19530,N_20217);
and U21046 (N_21046,N_19466,N_20102);
xnor U21047 (N_21047,N_19905,N_19738);
xor U21048 (N_21048,N_19698,N_20057);
or U21049 (N_21049,N_20295,N_20290);
nand U21050 (N_21050,N_20043,N_20272);
nor U21051 (N_21051,N_19359,N_19312);
and U21052 (N_21052,N_19460,N_20234);
nand U21053 (N_21053,N_19655,N_19344);
nor U21054 (N_21054,N_20155,N_19973);
or U21055 (N_21055,N_19773,N_20296);
and U21056 (N_21056,N_19514,N_19873);
nor U21057 (N_21057,N_19684,N_20020);
nand U21058 (N_21058,N_19793,N_19799);
nand U21059 (N_21059,N_19481,N_19219);
nand U21060 (N_21060,N_20010,N_19622);
xor U21061 (N_21061,N_20363,N_19795);
and U21062 (N_21062,N_19689,N_19856);
or U21063 (N_21063,N_19448,N_19532);
nand U21064 (N_21064,N_20037,N_19986);
or U21065 (N_21065,N_20312,N_19593);
nand U21066 (N_21066,N_19639,N_20050);
nand U21067 (N_21067,N_20332,N_19350);
nand U21068 (N_21068,N_19705,N_20136);
xor U21069 (N_21069,N_19666,N_19531);
xor U21070 (N_21070,N_19780,N_20305);
nand U21071 (N_21071,N_19439,N_19926);
nor U21072 (N_21072,N_20185,N_19600);
nor U21073 (N_21073,N_20174,N_19973);
and U21074 (N_21074,N_20193,N_19957);
nor U21075 (N_21075,N_19772,N_20258);
xor U21076 (N_21076,N_19444,N_19973);
nand U21077 (N_21077,N_19209,N_19401);
xnor U21078 (N_21078,N_19780,N_19219);
or U21079 (N_21079,N_19701,N_19956);
xor U21080 (N_21080,N_19986,N_20387);
xnor U21081 (N_21081,N_19579,N_19510);
and U21082 (N_21082,N_19419,N_19347);
or U21083 (N_21083,N_19719,N_20085);
nor U21084 (N_21084,N_20363,N_19443);
xnor U21085 (N_21085,N_19351,N_20056);
and U21086 (N_21086,N_20254,N_19852);
xnor U21087 (N_21087,N_19904,N_19958);
nor U21088 (N_21088,N_19492,N_19635);
and U21089 (N_21089,N_20128,N_20168);
and U21090 (N_21090,N_20371,N_19872);
or U21091 (N_21091,N_19745,N_19672);
and U21092 (N_21092,N_19508,N_19215);
xor U21093 (N_21093,N_19828,N_20027);
or U21094 (N_21094,N_19413,N_20279);
or U21095 (N_21095,N_19204,N_20160);
and U21096 (N_21096,N_19798,N_20200);
and U21097 (N_21097,N_19507,N_19664);
xor U21098 (N_21098,N_20295,N_19833);
nor U21099 (N_21099,N_20217,N_19877);
xnor U21100 (N_21100,N_19996,N_19205);
nor U21101 (N_21101,N_19586,N_19567);
xor U21102 (N_21102,N_19484,N_19891);
nor U21103 (N_21103,N_19634,N_20375);
nor U21104 (N_21104,N_19658,N_19750);
and U21105 (N_21105,N_19232,N_20321);
xnor U21106 (N_21106,N_20302,N_19818);
and U21107 (N_21107,N_20312,N_20149);
or U21108 (N_21108,N_19249,N_19260);
nand U21109 (N_21109,N_20268,N_19413);
nor U21110 (N_21110,N_19837,N_19746);
and U21111 (N_21111,N_20143,N_20270);
or U21112 (N_21112,N_20362,N_19433);
nand U21113 (N_21113,N_19991,N_19694);
nand U21114 (N_21114,N_19998,N_19672);
xnor U21115 (N_21115,N_19709,N_19834);
and U21116 (N_21116,N_19335,N_20115);
and U21117 (N_21117,N_19511,N_19514);
nor U21118 (N_21118,N_19759,N_19287);
nor U21119 (N_21119,N_19334,N_19284);
or U21120 (N_21120,N_20366,N_19355);
nand U21121 (N_21121,N_19410,N_19518);
and U21122 (N_21122,N_19896,N_19444);
and U21123 (N_21123,N_19432,N_19972);
and U21124 (N_21124,N_19483,N_19624);
nand U21125 (N_21125,N_19856,N_19845);
nand U21126 (N_21126,N_20266,N_19227);
xor U21127 (N_21127,N_19963,N_20240);
or U21128 (N_21128,N_19663,N_20208);
and U21129 (N_21129,N_19411,N_19763);
and U21130 (N_21130,N_20217,N_20260);
nand U21131 (N_21131,N_20380,N_19766);
or U21132 (N_21132,N_20061,N_20224);
or U21133 (N_21133,N_19263,N_19604);
and U21134 (N_21134,N_20143,N_19908);
nor U21135 (N_21135,N_19971,N_19830);
xor U21136 (N_21136,N_19921,N_19333);
and U21137 (N_21137,N_19489,N_19960);
nor U21138 (N_21138,N_19254,N_19320);
nand U21139 (N_21139,N_20210,N_20096);
or U21140 (N_21140,N_19973,N_19604);
and U21141 (N_21141,N_20047,N_19446);
nand U21142 (N_21142,N_19319,N_20079);
xnor U21143 (N_21143,N_20022,N_19308);
nand U21144 (N_21144,N_20354,N_19343);
nor U21145 (N_21145,N_19797,N_19616);
nand U21146 (N_21146,N_19767,N_19821);
nor U21147 (N_21147,N_20067,N_19340);
xnor U21148 (N_21148,N_20102,N_19755);
nor U21149 (N_21149,N_19820,N_19383);
xnor U21150 (N_21150,N_19683,N_19269);
nor U21151 (N_21151,N_19817,N_19446);
or U21152 (N_21152,N_20236,N_19666);
nand U21153 (N_21153,N_19434,N_19256);
nor U21154 (N_21154,N_20084,N_19752);
nand U21155 (N_21155,N_19433,N_19592);
or U21156 (N_21156,N_20346,N_19565);
and U21157 (N_21157,N_19296,N_19755);
or U21158 (N_21158,N_19368,N_19701);
nand U21159 (N_21159,N_19464,N_19444);
nor U21160 (N_21160,N_19348,N_19504);
and U21161 (N_21161,N_19210,N_19473);
nor U21162 (N_21162,N_19465,N_20234);
xnor U21163 (N_21163,N_19346,N_19218);
or U21164 (N_21164,N_20237,N_19689);
nand U21165 (N_21165,N_20191,N_19250);
nand U21166 (N_21166,N_20243,N_20048);
xnor U21167 (N_21167,N_19617,N_19364);
or U21168 (N_21168,N_20054,N_19745);
xnor U21169 (N_21169,N_20279,N_19652);
nor U21170 (N_21170,N_20069,N_20171);
and U21171 (N_21171,N_19591,N_20387);
and U21172 (N_21172,N_19593,N_19231);
nand U21173 (N_21173,N_19234,N_20266);
nor U21174 (N_21174,N_19869,N_19754);
xnor U21175 (N_21175,N_19519,N_19205);
or U21176 (N_21176,N_19728,N_19959);
or U21177 (N_21177,N_19886,N_19472);
and U21178 (N_21178,N_20316,N_19642);
nor U21179 (N_21179,N_20054,N_20284);
or U21180 (N_21180,N_20172,N_19473);
xor U21181 (N_21181,N_19361,N_20246);
or U21182 (N_21182,N_19288,N_19830);
nor U21183 (N_21183,N_20165,N_20033);
nand U21184 (N_21184,N_19698,N_19573);
or U21185 (N_21185,N_19395,N_20020);
nor U21186 (N_21186,N_20018,N_19922);
nor U21187 (N_21187,N_19614,N_19685);
nor U21188 (N_21188,N_19205,N_19874);
nand U21189 (N_21189,N_20211,N_19448);
or U21190 (N_21190,N_20106,N_20282);
nor U21191 (N_21191,N_19975,N_19607);
nand U21192 (N_21192,N_19481,N_19820);
or U21193 (N_21193,N_19763,N_20300);
or U21194 (N_21194,N_19622,N_19640);
or U21195 (N_21195,N_19365,N_20152);
and U21196 (N_21196,N_19367,N_20219);
nand U21197 (N_21197,N_19466,N_20360);
and U21198 (N_21198,N_20153,N_20188);
nand U21199 (N_21199,N_19445,N_19234);
nand U21200 (N_21200,N_19714,N_20341);
xnor U21201 (N_21201,N_20382,N_19424);
and U21202 (N_21202,N_19966,N_19642);
or U21203 (N_21203,N_20180,N_19349);
and U21204 (N_21204,N_19982,N_20359);
or U21205 (N_21205,N_19212,N_19551);
nor U21206 (N_21206,N_19306,N_20272);
and U21207 (N_21207,N_20309,N_19588);
nor U21208 (N_21208,N_19664,N_20299);
and U21209 (N_21209,N_20366,N_19789);
or U21210 (N_21210,N_19269,N_19723);
nand U21211 (N_21211,N_20153,N_19839);
nand U21212 (N_21212,N_20314,N_19912);
and U21213 (N_21213,N_19669,N_19754);
or U21214 (N_21214,N_19959,N_20022);
nand U21215 (N_21215,N_19770,N_19718);
or U21216 (N_21216,N_20173,N_20040);
and U21217 (N_21217,N_20255,N_19258);
and U21218 (N_21218,N_19640,N_19930);
nand U21219 (N_21219,N_20249,N_20254);
xnor U21220 (N_21220,N_19486,N_19282);
nand U21221 (N_21221,N_19388,N_19983);
and U21222 (N_21222,N_19830,N_19246);
or U21223 (N_21223,N_19461,N_19721);
nand U21224 (N_21224,N_20097,N_19822);
or U21225 (N_21225,N_19781,N_19307);
nand U21226 (N_21226,N_20189,N_19881);
nand U21227 (N_21227,N_19514,N_19986);
or U21228 (N_21228,N_20216,N_19303);
nor U21229 (N_21229,N_20282,N_20134);
and U21230 (N_21230,N_20059,N_19797);
and U21231 (N_21231,N_19828,N_19886);
or U21232 (N_21232,N_19720,N_19295);
nand U21233 (N_21233,N_20391,N_20088);
and U21234 (N_21234,N_19581,N_19348);
and U21235 (N_21235,N_19359,N_19544);
xnor U21236 (N_21236,N_19463,N_19345);
nand U21237 (N_21237,N_19629,N_19441);
nand U21238 (N_21238,N_19558,N_19463);
nand U21239 (N_21239,N_19673,N_20034);
and U21240 (N_21240,N_20164,N_20021);
nand U21241 (N_21241,N_19445,N_19593);
xor U21242 (N_21242,N_19622,N_19508);
and U21243 (N_21243,N_20316,N_20053);
xnor U21244 (N_21244,N_19467,N_19488);
or U21245 (N_21245,N_20076,N_19873);
nand U21246 (N_21246,N_19416,N_19888);
xnor U21247 (N_21247,N_20258,N_20040);
and U21248 (N_21248,N_19699,N_19208);
or U21249 (N_21249,N_20332,N_20314);
xnor U21250 (N_21250,N_19682,N_19888);
or U21251 (N_21251,N_20165,N_19968);
xor U21252 (N_21252,N_20398,N_19623);
xnor U21253 (N_21253,N_19940,N_20300);
xor U21254 (N_21254,N_19846,N_20352);
nand U21255 (N_21255,N_19250,N_20336);
and U21256 (N_21256,N_19451,N_19895);
and U21257 (N_21257,N_19490,N_20241);
nor U21258 (N_21258,N_19250,N_19286);
or U21259 (N_21259,N_20367,N_19716);
nand U21260 (N_21260,N_19919,N_20071);
and U21261 (N_21261,N_19977,N_19844);
or U21262 (N_21262,N_19396,N_19317);
xnor U21263 (N_21263,N_19390,N_19833);
nor U21264 (N_21264,N_19834,N_19485);
xnor U21265 (N_21265,N_19604,N_20182);
xnor U21266 (N_21266,N_20389,N_19712);
nor U21267 (N_21267,N_19779,N_19320);
xnor U21268 (N_21268,N_19880,N_19227);
xor U21269 (N_21269,N_19563,N_19228);
and U21270 (N_21270,N_20348,N_19893);
nor U21271 (N_21271,N_19797,N_19439);
xnor U21272 (N_21272,N_19722,N_19918);
xnor U21273 (N_21273,N_19787,N_20388);
nor U21274 (N_21274,N_20257,N_20046);
or U21275 (N_21275,N_19299,N_20136);
and U21276 (N_21276,N_20104,N_20332);
and U21277 (N_21277,N_20203,N_20390);
nand U21278 (N_21278,N_20030,N_19250);
or U21279 (N_21279,N_19633,N_20333);
xor U21280 (N_21280,N_19426,N_19457);
and U21281 (N_21281,N_19746,N_19551);
and U21282 (N_21282,N_20086,N_19924);
and U21283 (N_21283,N_19717,N_19417);
xor U21284 (N_21284,N_19488,N_19314);
xnor U21285 (N_21285,N_19545,N_19406);
or U21286 (N_21286,N_19637,N_20396);
xor U21287 (N_21287,N_19343,N_19920);
or U21288 (N_21288,N_20002,N_19381);
or U21289 (N_21289,N_19708,N_19748);
or U21290 (N_21290,N_20179,N_20229);
and U21291 (N_21291,N_19672,N_19764);
nor U21292 (N_21292,N_19611,N_19464);
or U21293 (N_21293,N_20026,N_20149);
nor U21294 (N_21294,N_20224,N_20205);
nand U21295 (N_21295,N_19235,N_20299);
nor U21296 (N_21296,N_19497,N_19324);
xor U21297 (N_21297,N_20019,N_20168);
nand U21298 (N_21298,N_19623,N_19387);
and U21299 (N_21299,N_19795,N_19225);
or U21300 (N_21300,N_19857,N_19934);
nand U21301 (N_21301,N_19878,N_20195);
xnor U21302 (N_21302,N_20140,N_19851);
nand U21303 (N_21303,N_19900,N_20043);
or U21304 (N_21304,N_20076,N_19900);
nand U21305 (N_21305,N_20160,N_19944);
or U21306 (N_21306,N_20352,N_19898);
nand U21307 (N_21307,N_19788,N_19792);
nor U21308 (N_21308,N_20135,N_20344);
and U21309 (N_21309,N_19924,N_20141);
nand U21310 (N_21310,N_19842,N_19624);
xnor U21311 (N_21311,N_20310,N_20260);
or U21312 (N_21312,N_20359,N_19824);
xor U21313 (N_21313,N_19372,N_19495);
and U21314 (N_21314,N_19324,N_19737);
nor U21315 (N_21315,N_19221,N_19722);
nand U21316 (N_21316,N_20347,N_20291);
or U21317 (N_21317,N_19676,N_19892);
xnor U21318 (N_21318,N_20254,N_20390);
and U21319 (N_21319,N_19604,N_20356);
nand U21320 (N_21320,N_19589,N_19733);
xnor U21321 (N_21321,N_20167,N_19568);
nand U21322 (N_21322,N_19641,N_19207);
or U21323 (N_21323,N_20001,N_19805);
nor U21324 (N_21324,N_20121,N_20146);
nor U21325 (N_21325,N_19618,N_19826);
and U21326 (N_21326,N_19314,N_19740);
or U21327 (N_21327,N_19758,N_19602);
or U21328 (N_21328,N_20253,N_20275);
or U21329 (N_21329,N_20379,N_19917);
and U21330 (N_21330,N_19205,N_19789);
or U21331 (N_21331,N_20151,N_20216);
nor U21332 (N_21332,N_19769,N_19323);
and U21333 (N_21333,N_20090,N_19761);
nor U21334 (N_21334,N_19859,N_19913);
nand U21335 (N_21335,N_19863,N_19365);
xnor U21336 (N_21336,N_19785,N_19890);
xor U21337 (N_21337,N_20358,N_19367);
nor U21338 (N_21338,N_19363,N_20227);
nor U21339 (N_21339,N_20256,N_20206);
nand U21340 (N_21340,N_20372,N_19566);
nand U21341 (N_21341,N_20221,N_20168);
and U21342 (N_21342,N_19894,N_20003);
and U21343 (N_21343,N_19295,N_20276);
and U21344 (N_21344,N_20320,N_20139);
nor U21345 (N_21345,N_19814,N_19920);
nand U21346 (N_21346,N_19405,N_19523);
xor U21347 (N_21347,N_20030,N_19244);
and U21348 (N_21348,N_19805,N_19355);
xor U21349 (N_21349,N_20197,N_19681);
xnor U21350 (N_21350,N_19771,N_20345);
nand U21351 (N_21351,N_19910,N_19790);
nor U21352 (N_21352,N_19339,N_19629);
xnor U21353 (N_21353,N_19628,N_19395);
nor U21354 (N_21354,N_20382,N_19692);
or U21355 (N_21355,N_19355,N_19743);
nor U21356 (N_21356,N_19534,N_19642);
nor U21357 (N_21357,N_19511,N_20044);
and U21358 (N_21358,N_19331,N_20177);
nand U21359 (N_21359,N_19237,N_19945);
and U21360 (N_21360,N_19645,N_19772);
or U21361 (N_21361,N_19701,N_19934);
nor U21362 (N_21362,N_20300,N_19648);
nor U21363 (N_21363,N_19605,N_19688);
or U21364 (N_21364,N_20205,N_20308);
nand U21365 (N_21365,N_20256,N_19816);
nor U21366 (N_21366,N_19661,N_19614);
nand U21367 (N_21367,N_20354,N_19510);
and U21368 (N_21368,N_19865,N_19507);
nand U21369 (N_21369,N_19641,N_19591);
xor U21370 (N_21370,N_19820,N_19613);
xnor U21371 (N_21371,N_19928,N_19273);
nor U21372 (N_21372,N_19941,N_19431);
or U21373 (N_21373,N_19674,N_19604);
nor U21374 (N_21374,N_19808,N_20239);
or U21375 (N_21375,N_20111,N_20337);
xnor U21376 (N_21376,N_19762,N_19338);
or U21377 (N_21377,N_19233,N_20237);
nand U21378 (N_21378,N_19620,N_19692);
nand U21379 (N_21379,N_19587,N_19760);
nand U21380 (N_21380,N_19441,N_19975);
and U21381 (N_21381,N_20387,N_20225);
or U21382 (N_21382,N_20069,N_19731);
or U21383 (N_21383,N_20004,N_19510);
nand U21384 (N_21384,N_19399,N_19606);
nor U21385 (N_21385,N_19719,N_19219);
or U21386 (N_21386,N_19384,N_20097);
or U21387 (N_21387,N_19879,N_19945);
and U21388 (N_21388,N_20355,N_19397);
and U21389 (N_21389,N_19354,N_20036);
nand U21390 (N_21390,N_19981,N_19945);
or U21391 (N_21391,N_20316,N_19478);
xor U21392 (N_21392,N_20159,N_19917);
or U21393 (N_21393,N_20387,N_20296);
xnor U21394 (N_21394,N_19880,N_20157);
xor U21395 (N_21395,N_19912,N_19444);
nand U21396 (N_21396,N_19230,N_19604);
and U21397 (N_21397,N_19287,N_20209);
xor U21398 (N_21398,N_20315,N_19883);
or U21399 (N_21399,N_20208,N_19434);
nand U21400 (N_21400,N_20295,N_19912);
and U21401 (N_21401,N_20198,N_20141);
xor U21402 (N_21402,N_19520,N_19659);
or U21403 (N_21403,N_19781,N_19257);
xnor U21404 (N_21404,N_20185,N_19847);
and U21405 (N_21405,N_20110,N_19693);
and U21406 (N_21406,N_20202,N_19845);
nand U21407 (N_21407,N_19432,N_19660);
xor U21408 (N_21408,N_20192,N_19558);
or U21409 (N_21409,N_20188,N_19942);
or U21410 (N_21410,N_19407,N_19863);
and U21411 (N_21411,N_19744,N_20346);
nand U21412 (N_21412,N_20271,N_19673);
nor U21413 (N_21413,N_19775,N_19442);
and U21414 (N_21414,N_19849,N_19802);
nor U21415 (N_21415,N_20256,N_19957);
nor U21416 (N_21416,N_19248,N_19323);
and U21417 (N_21417,N_19304,N_19919);
or U21418 (N_21418,N_19308,N_19775);
xor U21419 (N_21419,N_19609,N_20335);
and U21420 (N_21420,N_19941,N_19832);
and U21421 (N_21421,N_20294,N_19912);
xnor U21422 (N_21422,N_19275,N_20129);
and U21423 (N_21423,N_20024,N_19907);
xor U21424 (N_21424,N_19240,N_20377);
or U21425 (N_21425,N_19471,N_20038);
and U21426 (N_21426,N_19381,N_20000);
nor U21427 (N_21427,N_20152,N_19550);
and U21428 (N_21428,N_19450,N_20307);
or U21429 (N_21429,N_19636,N_19722);
nor U21430 (N_21430,N_20298,N_19636);
xor U21431 (N_21431,N_19861,N_19286);
and U21432 (N_21432,N_19896,N_19527);
nor U21433 (N_21433,N_19752,N_19351);
or U21434 (N_21434,N_19361,N_19645);
nand U21435 (N_21435,N_20151,N_19535);
and U21436 (N_21436,N_20174,N_19537);
nand U21437 (N_21437,N_19305,N_20035);
nand U21438 (N_21438,N_20313,N_19446);
xnor U21439 (N_21439,N_20230,N_20288);
nand U21440 (N_21440,N_19395,N_19979);
nand U21441 (N_21441,N_19769,N_20002);
and U21442 (N_21442,N_20351,N_19992);
or U21443 (N_21443,N_19923,N_19302);
nor U21444 (N_21444,N_20383,N_20138);
xor U21445 (N_21445,N_19866,N_19983);
xnor U21446 (N_21446,N_19983,N_19532);
xnor U21447 (N_21447,N_19483,N_19232);
nor U21448 (N_21448,N_19968,N_20013);
nor U21449 (N_21449,N_20310,N_19519);
nand U21450 (N_21450,N_19992,N_20145);
or U21451 (N_21451,N_19291,N_20061);
nor U21452 (N_21452,N_20118,N_19443);
nor U21453 (N_21453,N_20045,N_19808);
xnor U21454 (N_21454,N_20094,N_19378);
xnor U21455 (N_21455,N_19794,N_20079);
nand U21456 (N_21456,N_19715,N_19739);
and U21457 (N_21457,N_19330,N_20098);
or U21458 (N_21458,N_19885,N_19590);
nand U21459 (N_21459,N_19911,N_19632);
nor U21460 (N_21460,N_19211,N_20107);
or U21461 (N_21461,N_20232,N_19299);
nand U21462 (N_21462,N_19729,N_19926);
or U21463 (N_21463,N_19478,N_20365);
nand U21464 (N_21464,N_20019,N_19304);
nor U21465 (N_21465,N_20356,N_19549);
or U21466 (N_21466,N_20310,N_20302);
nand U21467 (N_21467,N_19386,N_20394);
and U21468 (N_21468,N_19420,N_20241);
xnor U21469 (N_21469,N_20147,N_19891);
nor U21470 (N_21470,N_20147,N_19976);
and U21471 (N_21471,N_20245,N_19885);
nor U21472 (N_21472,N_20068,N_20317);
and U21473 (N_21473,N_20150,N_20324);
nor U21474 (N_21474,N_19966,N_19514);
xor U21475 (N_21475,N_20273,N_19230);
and U21476 (N_21476,N_19767,N_19848);
xnor U21477 (N_21477,N_19708,N_19200);
and U21478 (N_21478,N_19635,N_19591);
and U21479 (N_21479,N_19879,N_19475);
nor U21480 (N_21480,N_19521,N_19308);
xnor U21481 (N_21481,N_20106,N_19901);
xor U21482 (N_21482,N_19412,N_20089);
nor U21483 (N_21483,N_19212,N_19871);
and U21484 (N_21484,N_20399,N_19752);
nor U21485 (N_21485,N_19941,N_19395);
nor U21486 (N_21486,N_20101,N_19466);
xor U21487 (N_21487,N_20001,N_20320);
xnor U21488 (N_21488,N_19917,N_19331);
and U21489 (N_21489,N_19987,N_19901);
nand U21490 (N_21490,N_20351,N_20027);
and U21491 (N_21491,N_20250,N_19628);
nand U21492 (N_21492,N_19570,N_20372);
xor U21493 (N_21493,N_19644,N_19323);
xor U21494 (N_21494,N_19431,N_19249);
nand U21495 (N_21495,N_19711,N_19890);
or U21496 (N_21496,N_19723,N_19863);
nor U21497 (N_21497,N_19638,N_19562);
nand U21498 (N_21498,N_20147,N_20186);
nor U21499 (N_21499,N_20029,N_20023);
or U21500 (N_21500,N_20151,N_19923);
and U21501 (N_21501,N_19397,N_20174);
or U21502 (N_21502,N_19521,N_19392);
and U21503 (N_21503,N_19528,N_20147);
nor U21504 (N_21504,N_20243,N_20265);
xnor U21505 (N_21505,N_19959,N_19879);
nor U21506 (N_21506,N_19653,N_19809);
or U21507 (N_21507,N_19768,N_19931);
or U21508 (N_21508,N_19788,N_20075);
nand U21509 (N_21509,N_20256,N_20166);
and U21510 (N_21510,N_19389,N_19661);
nor U21511 (N_21511,N_19421,N_19847);
xnor U21512 (N_21512,N_20057,N_19499);
and U21513 (N_21513,N_19300,N_19610);
or U21514 (N_21514,N_20163,N_19630);
xor U21515 (N_21515,N_19549,N_19365);
nand U21516 (N_21516,N_20355,N_19372);
xor U21517 (N_21517,N_20029,N_19399);
or U21518 (N_21518,N_19741,N_19237);
nand U21519 (N_21519,N_19949,N_19733);
or U21520 (N_21520,N_20249,N_19685);
nor U21521 (N_21521,N_20018,N_19345);
nand U21522 (N_21522,N_19640,N_19867);
nor U21523 (N_21523,N_20199,N_20069);
xnor U21524 (N_21524,N_20263,N_19758);
or U21525 (N_21525,N_19963,N_20242);
and U21526 (N_21526,N_19344,N_20056);
nand U21527 (N_21527,N_19662,N_19652);
and U21528 (N_21528,N_20323,N_19802);
and U21529 (N_21529,N_19542,N_19853);
nand U21530 (N_21530,N_20000,N_20275);
or U21531 (N_21531,N_19849,N_19751);
nand U21532 (N_21532,N_19226,N_19350);
and U21533 (N_21533,N_19214,N_19991);
and U21534 (N_21534,N_19623,N_19765);
nor U21535 (N_21535,N_20117,N_19777);
or U21536 (N_21536,N_19904,N_19485);
nand U21537 (N_21537,N_19742,N_20081);
and U21538 (N_21538,N_19577,N_19882);
or U21539 (N_21539,N_19247,N_19589);
and U21540 (N_21540,N_20001,N_19268);
nor U21541 (N_21541,N_20353,N_20211);
nor U21542 (N_21542,N_19269,N_20150);
or U21543 (N_21543,N_19276,N_19840);
or U21544 (N_21544,N_20240,N_19683);
nand U21545 (N_21545,N_19324,N_19447);
xor U21546 (N_21546,N_19746,N_19377);
nor U21547 (N_21547,N_20179,N_19529);
xnor U21548 (N_21548,N_20242,N_19328);
nand U21549 (N_21549,N_20015,N_19729);
nor U21550 (N_21550,N_20231,N_19984);
and U21551 (N_21551,N_19930,N_20250);
nand U21552 (N_21552,N_20380,N_19768);
and U21553 (N_21553,N_20366,N_19309);
xnor U21554 (N_21554,N_19445,N_20052);
or U21555 (N_21555,N_19371,N_20127);
xnor U21556 (N_21556,N_20348,N_19426);
nand U21557 (N_21557,N_19627,N_19875);
and U21558 (N_21558,N_20338,N_19929);
nor U21559 (N_21559,N_19498,N_19647);
nand U21560 (N_21560,N_19496,N_19535);
nor U21561 (N_21561,N_20305,N_20118);
xnor U21562 (N_21562,N_19447,N_20298);
or U21563 (N_21563,N_20202,N_20323);
nand U21564 (N_21564,N_19823,N_20096);
and U21565 (N_21565,N_19896,N_19839);
nor U21566 (N_21566,N_19462,N_19333);
nor U21567 (N_21567,N_20050,N_19225);
nor U21568 (N_21568,N_19556,N_19805);
nor U21569 (N_21569,N_19804,N_19529);
xor U21570 (N_21570,N_20256,N_19245);
or U21571 (N_21571,N_19296,N_19982);
nor U21572 (N_21572,N_19763,N_19400);
and U21573 (N_21573,N_20257,N_19853);
or U21574 (N_21574,N_20061,N_19602);
nand U21575 (N_21575,N_20179,N_19858);
and U21576 (N_21576,N_19856,N_19248);
nor U21577 (N_21577,N_19821,N_20149);
nand U21578 (N_21578,N_19461,N_19453);
and U21579 (N_21579,N_20350,N_19580);
nor U21580 (N_21580,N_20166,N_19851);
or U21581 (N_21581,N_19908,N_20155);
nor U21582 (N_21582,N_20116,N_20120);
or U21583 (N_21583,N_19904,N_19722);
nand U21584 (N_21584,N_20026,N_19580);
nand U21585 (N_21585,N_19372,N_19853);
and U21586 (N_21586,N_19775,N_19898);
nor U21587 (N_21587,N_19356,N_19905);
xor U21588 (N_21588,N_19574,N_20054);
nand U21589 (N_21589,N_19594,N_20367);
or U21590 (N_21590,N_19220,N_20198);
and U21591 (N_21591,N_20158,N_20196);
or U21592 (N_21592,N_19622,N_19647);
nor U21593 (N_21593,N_19700,N_19548);
xor U21594 (N_21594,N_20173,N_19496);
and U21595 (N_21595,N_19274,N_19487);
or U21596 (N_21596,N_19519,N_19618);
and U21597 (N_21597,N_20148,N_19747);
xor U21598 (N_21598,N_20292,N_19681);
nand U21599 (N_21599,N_19788,N_19451);
and U21600 (N_21600,N_20985,N_21596);
or U21601 (N_21601,N_20690,N_20776);
and U21602 (N_21602,N_21031,N_21183);
and U21603 (N_21603,N_20511,N_20525);
nor U21604 (N_21604,N_21045,N_20559);
xor U21605 (N_21605,N_21259,N_20713);
or U21606 (N_21606,N_20947,N_21281);
nor U21607 (N_21607,N_21148,N_21426);
nand U21608 (N_21608,N_21108,N_21368);
or U21609 (N_21609,N_20978,N_20876);
or U21610 (N_21610,N_21138,N_20849);
nand U21611 (N_21611,N_20793,N_21157);
and U21612 (N_21612,N_21057,N_21216);
and U21613 (N_21613,N_20722,N_21127);
nand U21614 (N_21614,N_21122,N_21382);
nor U21615 (N_21615,N_21350,N_20547);
or U21616 (N_21616,N_20660,N_21161);
nor U21617 (N_21617,N_20774,N_21001);
or U21618 (N_21618,N_21591,N_20972);
and U21619 (N_21619,N_21209,N_21405);
nor U21620 (N_21620,N_21218,N_21344);
nor U21621 (N_21621,N_21531,N_21552);
xnor U21622 (N_21622,N_21356,N_20931);
xnor U21623 (N_21623,N_21347,N_20500);
and U21624 (N_21624,N_20683,N_20451);
or U21625 (N_21625,N_20880,N_20457);
xor U21626 (N_21626,N_20494,N_21064);
xor U21627 (N_21627,N_21567,N_20838);
and U21628 (N_21628,N_21118,N_20517);
and U21629 (N_21629,N_21337,N_21149);
or U21630 (N_21630,N_20999,N_21571);
or U21631 (N_21631,N_20790,N_20484);
xor U21632 (N_21632,N_20897,N_20493);
nand U21633 (N_21633,N_20724,N_21162);
or U21634 (N_21634,N_21179,N_21354);
nor U21635 (N_21635,N_21065,N_21555);
xnor U21636 (N_21636,N_20618,N_21488);
and U21637 (N_21637,N_20888,N_20811);
and U21638 (N_21638,N_20946,N_20551);
or U21639 (N_21639,N_21137,N_21251);
xor U21640 (N_21640,N_21005,N_20856);
nand U21641 (N_21641,N_20651,N_20958);
nor U21642 (N_21642,N_20658,N_21314);
nand U21643 (N_21643,N_20430,N_20821);
nand U21644 (N_21644,N_21178,N_20804);
nand U21645 (N_21645,N_21074,N_20687);
and U21646 (N_21646,N_21007,N_20626);
or U21647 (N_21647,N_21482,N_21174);
and U21648 (N_21648,N_21070,N_20749);
or U21649 (N_21649,N_20772,N_21263);
or U21650 (N_21650,N_21252,N_21526);
and U21651 (N_21651,N_21111,N_21208);
nor U21652 (N_21652,N_20432,N_20934);
xor U21653 (N_21653,N_20413,N_20645);
nand U21654 (N_21654,N_20447,N_21379);
or U21655 (N_21655,N_20665,N_20684);
xor U21656 (N_21656,N_20602,N_20697);
xnor U21657 (N_21657,N_21246,N_20608);
xnor U21658 (N_21658,N_20536,N_21414);
or U21659 (N_21659,N_20682,N_21302);
nand U21660 (N_21660,N_21508,N_21581);
and U21661 (N_21661,N_20706,N_20438);
nand U21662 (N_21662,N_21052,N_21260);
xnor U21663 (N_21663,N_20435,N_21400);
or U21664 (N_21664,N_21398,N_20686);
or U21665 (N_21665,N_21120,N_21322);
or U21666 (N_21666,N_21325,N_20534);
xor U21667 (N_21667,N_20858,N_20747);
xor U21668 (N_21668,N_20795,N_20777);
or U21669 (N_21669,N_21242,N_21357);
or U21670 (N_21670,N_20540,N_21318);
or U21671 (N_21671,N_20431,N_20485);
or U21672 (N_21672,N_20553,N_21213);
nor U21673 (N_21673,N_20967,N_20615);
nand U21674 (N_21674,N_21087,N_21291);
xor U21675 (N_21675,N_21163,N_20845);
and U21676 (N_21676,N_20598,N_20567);
or U21677 (N_21677,N_21570,N_21239);
and U21678 (N_21678,N_20760,N_21572);
and U21679 (N_21679,N_21026,N_20533);
nand U21680 (N_21680,N_21060,N_20711);
and U21681 (N_21681,N_21305,N_21378);
xnor U21682 (N_21682,N_21447,N_20609);
nor U21683 (N_21683,N_21542,N_20703);
nand U21684 (N_21684,N_21459,N_21268);
or U21685 (N_21685,N_20418,N_20773);
and U21686 (N_21686,N_21222,N_20635);
xor U21687 (N_21687,N_20782,N_21470);
nor U21688 (N_21688,N_20864,N_20653);
nor U21689 (N_21689,N_21015,N_20745);
or U21690 (N_21690,N_20977,N_21128);
or U21691 (N_21691,N_20610,N_20810);
xnor U21692 (N_21692,N_21427,N_21227);
xnor U21693 (N_21693,N_21105,N_20943);
and U21694 (N_21694,N_20488,N_21384);
or U21695 (N_21695,N_20663,N_21022);
or U21696 (N_21696,N_21450,N_20583);
xor U21697 (N_21697,N_21495,N_21404);
and U21698 (N_21698,N_21143,N_21520);
nand U21699 (N_21699,N_21392,N_21264);
nor U21700 (N_21700,N_21433,N_20673);
or U21701 (N_21701,N_21309,N_21124);
and U21702 (N_21702,N_20969,N_21288);
nand U21703 (N_21703,N_21301,N_20719);
and U21704 (N_21704,N_20467,N_21593);
or U21705 (N_21705,N_20539,N_21468);
and U21706 (N_21706,N_20736,N_21525);
nor U21707 (N_21707,N_21096,N_20529);
or U21708 (N_21708,N_20407,N_21206);
nand U21709 (N_21709,N_20971,N_20521);
and U21710 (N_21710,N_20837,N_21412);
or U21711 (N_21711,N_20566,N_21235);
nand U21712 (N_21712,N_21294,N_20925);
xor U21713 (N_21713,N_21088,N_20465);
or U21714 (N_21714,N_20405,N_21093);
nand U21715 (N_21715,N_21519,N_20460);
or U21716 (N_21716,N_20855,N_21214);
or U21717 (N_21717,N_20800,N_21406);
nand U21718 (N_21718,N_20834,N_21123);
nand U21719 (N_21719,N_20680,N_21316);
nor U21720 (N_21720,N_21276,N_21456);
nor U21721 (N_21721,N_20427,N_21272);
xnor U21722 (N_21722,N_21377,N_20434);
or U21723 (N_21723,N_21097,N_21312);
and U21724 (N_21724,N_20735,N_20937);
nor U21725 (N_21725,N_21241,N_20481);
and U21726 (N_21726,N_20454,N_20667);
and U21727 (N_21727,N_20926,N_21478);
and U21728 (N_21728,N_20678,N_20759);
nand U21729 (N_21729,N_20846,N_20953);
or U21730 (N_21730,N_20998,N_21202);
or U21731 (N_21731,N_20576,N_21422);
xnor U21732 (N_21732,N_21550,N_21089);
nand U21733 (N_21733,N_20631,N_21223);
or U21734 (N_21734,N_20633,N_20798);
nor U21735 (N_21735,N_21373,N_20844);
nand U21736 (N_21736,N_21198,N_20813);
or U21737 (N_21737,N_20504,N_20780);
or U21738 (N_21738,N_21579,N_21467);
nand U21739 (N_21739,N_21011,N_21189);
nor U21740 (N_21740,N_21561,N_20718);
and U21741 (N_21741,N_20968,N_20535);
nor U21742 (N_21742,N_21393,N_21320);
xnor U21743 (N_21743,N_20650,N_20445);
nor U21744 (N_21744,N_20412,N_21187);
and U21745 (N_21745,N_21131,N_20916);
xnor U21746 (N_21746,N_21410,N_21522);
xor U21747 (N_21747,N_20738,N_21255);
or U21748 (N_21748,N_20505,N_20563);
nor U21749 (N_21749,N_20848,N_20612);
and U21750 (N_21750,N_21315,N_21076);
or U21751 (N_21751,N_20901,N_20872);
nor U21752 (N_21752,N_21154,N_21006);
or U21753 (N_21753,N_20879,N_20584);
xor U21754 (N_21754,N_21429,N_21201);
and U21755 (N_21755,N_21588,N_20955);
xor U21756 (N_21756,N_21020,N_20932);
xnor U21757 (N_21757,N_20816,N_21266);
nand U21758 (N_21758,N_21539,N_21498);
nor U21759 (N_21759,N_21566,N_21421);
and U21760 (N_21760,N_21224,N_21469);
and U21761 (N_21761,N_21132,N_21317);
nand U21762 (N_21762,N_20865,N_21051);
and U21763 (N_21763,N_21182,N_21510);
nor U21764 (N_21764,N_20588,N_20456);
xnor U21765 (N_21765,N_20919,N_21441);
nand U21766 (N_21766,N_20979,N_20582);
nand U21767 (N_21767,N_20662,N_21190);
and U21768 (N_21768,N_21086,N_21136);
nor U21769 (N_21769,N_21541,N_20996);
or U21770 (N_21770,N_20611,N_21518);
or U21771 (N_21771,N_20907,N_20409);
xor U21772 (N_21772,N_20619,N_21017);
nand U21773 (N_21773,N_21551,N_21129);
and U21774 (N_21774,N_21115,N_21340);
xnor U21775 (N_21775,N_20963,N_20519);
or U21776 (N_21776,N_20512,N_21328);
nand U21777 (N_21777,N_20538,N_20779);
nand U21778 (N_21778,N_21346,N_21121);
and U21779 (N_21779,N_20765,N_21409);
or U21780 (N_21780,N_20927,N_21166);
nor U21781 (N_21781,N_21059,N_21338);
or U21782 (N_21782,N_21509,N_20941);
nor U21783 (N_21783,N_21164,N_20993);
and U21784 (N_21784,N_20560,N_21430);
and U21785 (N_21785,N_20840,N_21298);
nand U21786 (N_21786,N_20905,N_20617);
xnor U21787 (N_21787,N_21432,N_20448);
nand U21788 (N_21788,N_20604,N_21025);
and U21789 (N_21789,N_20984,N_20516);
nor U21790 (N_21790,N_20439,N_20891);
xnor U21791 (N_21791,N_21032,N_21390);
or U21792 (N_21792,N_21528,N_21027);
and U21793 (N_21793,N_21130,N_20899);
and U21794 (N_21794,N_21363,N_21226);
and U21795 (N_21795,N_20752,N_20928);
nor U21796 (N_21796,N_21590,N_20699);
xnor U21797 (N_21797,N_21535,N_21313);
nor U21798 (N_21798,N_20642,N_21262);
nor U21799 (N_21799,N_20657,N_20903);
or U21800 (N_21800,N_20802,N_20961);
nor U21801 (N_21801,N_21273,N_21040);
nand U21802 (N_21802,N_21497,N_21104);
or U21803 (N_21803,N_21077,N_21361);
nand U21804 (N_21804,N_20557,N_21286);
and U21805 (N_21805,N_20898,N_21385);
xor U21806 (N_21806,N_21444,N_21355);
nor U21807 (N_21807,N_21293,N_20807);
xor U21808 (N_21808,N_21254,N_20601);
xor U21809 (N_21809,N_21362,N_20710);
or U21810 (N_21810,N_20863,N_20712);
and U21811 (N_21811,N_21503,N_20693);
nand U21812 (N_21812,N_20675,N_20704);
nor U21813 (N_21813,N_21496,N_20526);
or U21814 (N_21814,N_20750,N_21270);
xnor U21815 (N_21815,N_21543,N_20530);
or U21816 (N_21816,N_21343,N_21176);
nand U21817 (N_21817,N_20873,N_21376);
nand U21818 (N_21818,N_21290,N_21307);
nand U21819 (N_21819,N_20669,N_21577);
nand U21820 (N_21820,N_20606,N_20854);
and U21821 (N_21821,N_20918,N_20761);
xor U21822 (N_21822,N_20694,N_20778);
and U21823 (N_21823,N_21153,N_20733);
nor U21824 (N_21824,N_21391,N_20462);
or U21825 (N_21825,N_20769,N_21063);
or U21826 (N_21826,N_20952,N_21245);
or U21827 (N_21827,N_20988,N_20990);
xor U21828 (N_21828,N_20671,N_20823);
nand U21829 (N_21829,N_21003,N_20995);
xor U21830 (N_21830,N_21486,N_21387);
nor U21831 (N_21831,N_20513,N_21348);
nor U21832 (N_21832,N_21126,N_21173);
nand U21833 (N_21833,N_21574,N_20477);
xor U21834 (N_21834,N_21587,N_21184);
nand U21835 (N_21835,N_20991,N_21267);
nand U21836 (N_21836,N_20832,N_20755);
or U21837 (N_21837,N_20422,N_21479);
or U21838 (N_21838,N_21280,N_21169);
or U21839 (N_21839,N_21014,N_20746);
and U21840 (N_21840,N_21069,N_21553);
and U21841 (N_21841,N_21146,N_20753);
xnor U21842 (N_21842,N_20792,N_20835);
xnor U21843 (N_21843,N_20709,N_20981);
nor U21844 (N_21844,N_21461,N_20674);
or U21845 (N_21845,N_21407,N_20799);
or U21846 (N_21846,N_20417,N_21033);
and U21847 (N_21847,N_21297,N_21047);
or U21848 (N_21848,N_21194,N_20910);
and U21849 (N_21849,N_20767,N_21394);
nor U21850 (N_21850,N_20920,N_21053);
nor U21851 (N_21851,N_20809,N_20411);
nor U21852 (N_21852,N_21466,N_21156);
and U21853 (N_21853,N_21413,N_21342);
and U21854 (N_21854,N_20625,N_21329);
xnor U21855 (N_21855,N_21349,N_21172);
and U21856 (N_21856,N_21012,N_20442);
or U21857 (N_21857,N_20890,N_21514);
nor U21858 (N_21858,N_21303,N_20531);
nand U21859 (N_21859,N_21168,N_20831);
and U21860 (N_21860,N_20884,N_21283);
xor U21861 (N_21861,N_20497,N_20424);
nand U21862 (N_21862,N_20554,N_20572);
nand U21863 (N_21863,N_20702,N_21576);
or U21864 (N_21864,N_20957,N_21592);
nand U21865 (N_21865,N_20740,N_20900);
xnor U21866 (N_21866,N_21389,N_20624);
or U21867 (N_21867,N_20661,N_20692);
nor U21868 (N_21868,N_21358,N_20788);
or U21869 (N_21869,N_21352,N_20942);
nor U21870 (N_21870,N_20587,N_21490);
nor U21871 (N_21871,N_20593,N_21151);
xnor U21872 (N_21872,N_21499,N_21269);
xnor U21873 (N_21873,N_21304,N_20819);
nor U21874 (N_21874,N_21068,N_21489);
nor U21875 (N_21875,N_20695,N_20647);
and U21876 (N_21876,N_21049,N_20426);
xor U21877 (N_21877,N_21050,N_21544);
nand U21878 (N_21878,N_20577,N_20469);
xor U21879 (N_21879,N_20503,N_21037);
xor U21880 (N_21880,N_20830,N_20794);
and U21881 (N_21881,N_21275,N_21473);
nor U21882 (N_21882,N_21125,N_20817);
nand U21883 (N_21883,N_21249,N_21333);
nor U21884 (N_21884,N_20425,N_21370);
nand U21885 (N_21885,N_20524,N_20762);
and U21886 (N_21886,N_21464,N_21000);
or U21887 (N_21887,N_20781,N_21423);
nor U21888 (N_21888,N_21434,N_20970);
or U21889 (N_21889,N_21009,N_21028);
or U21890 (N_21890,N_20805,N_20532);
xnor U21891 (N_21891,N_20550,N_20537);
nor U21892 (N_21892,N_20616,N_21471);
or U21893 (N_21893,N_20771,N_21462);
xor U21894 (N_21894,N_21147,N_21487);
nor U21895 (N_21895,N_20664,N_21061);
nand U21896 (N_21896,N_20480,N_20851);
and U21897 (N_21897,N_20894,N_20744);
nand U21898 (N_21898,N_21475,N_21085);
nor U21899 (N_21899,N_21265,N_21103);
nand U21900 (N_21900,N_21079,N_20676);
nand U21901 (N_21901,N_21439,N_20476);
nor U21902 (N_21902,N_20466,N_20419);
nor U21903 (N_21903,N_21424,N_21282);
or U21904 (N_21904,N_21133,N_21181);
or U21905 (N_21905,N_20472,N_21081);
nor U21906 (N_21906,N_21196,N_20654);
nor U21907 (N_21907,N_21277,N_20886);
or U21908 (N_21908,N_21205,N_21021);
or U21909 (N_21909,N_21537,N_21300);
nand U21910 (N_21910,N_20763,N_21578);
and U21911 (N_21911,N_20887,N_21159);
or U21912 (N_21912,N_21199,N_20429);
nor U21913 (N_21913,N_21425,N_20965);
nand U21914 (N_21914,N_21231,N_20685);
or U21915 (N_21915,N_20428,N_21100);
nor U21916 (N_21916,N_20473,N_21521);
or U21917 (N_21917,N_21474,N_21372);
xnor U21918 (N_21918,N_20726,N_21106);
or U21919 (N_21919,N_20571,N_21369);
xor U21920 (N_21920,N_20789,N_21326);
nand U21921 (N_21921,N_20670,N_20406);
and U21922 (N_21922,N_20637,N_20549);
or U21923 (N_21923,N_20696,N_20591);
xor U21924 (N_21924,N_21236,N_20951);
or U21925 (N_21925,N_21257,N_20446);
nor U21926 (N_21926,N_20478,N_20461);
xnor U21927 (N_21927,N_21084,N_21397);
xor U21928 (N_21928,N_21460,N_21319);
xnor U21929 (N_21929,N_21080,N_20496);
nand U21930 (N_21930,N_21504,N_20677);
nor U21931 (N_21931,N_21371,N_21197);
nand U21932 (N_21932,N_20956,N_20708);
xnor U21933 (N_21933,N_21102,N_21072);
or U21934 (N_21934,N_20590,N_21442);
nor U21935 (N_21935,N_21465,N_20607);
nor U21936 (N_21936,N_20764,N_21284);
or U21937 (N_21937,N_21240,N_21054);
nor U21938 (N_21938,N_21062,N_20510);
xor U21939 (N_21939,N_21417,N_21203);
nand U21940 (N_21940,N_20518,N_21367);
nor U21941 (N_21941,N_21233,N_20785);
and U21942 (N_21942,N_20882,N_20911);
xnor U21943 (N_21943,N_20906,N_20597);
nor U21944 (N_21944,N_20909,N_20471);
or U21945 (N_21945,N_20786,N_21219);
nor U21946 (N_21946,N_20867,N_21436);
xor U21947 (N_21947,N_20975,N_20640);
nand U21948 (N_21948,N_21386,N_20976);
nand U21949 (N_21949,N_21380,N_21211);
nor U21950 (N_21950,N_21457,N_20861);
nor U21951 (N_21951,N_20555,N_21180);
and U21952 (N_21952,N_21285,N_21279);
or U21953 (N_21953,N_20543,N_20499);
and U21954 (N_21954,N_20935,N_21292);
xnor U21955 (N_21955,N_21110,N_21010);
and U21956 (N_21956,N_20948,N_20562);
xnor U21957 (N_21957,N_20679,N_21287);
nand U21958 (N_21958,N_20960,N_21098);
or U21959 (N_21959,N_21381,N_20623);
nand U21960 (N_21960,N_20648,N_20564);
or U21961 (N_21961,N_20644,N_21044);
nor U21962 (N_21962,N_21212,N_20475);
or U21963 (N_21963,N_21418,N_20402);
and U21964 (N_21964,N_21220,N_21402);
nor U21965 (N_21965,N_20453,N_21582);
or U21966 (N_21966,N_21472,N_20913);
xor U21967 (N_21967,N_21351,N_20627);
nor U21968 (N_21968,N_21152,N_21411);
and U21969 (N_21969,N_21034,N_20507);
and U21970 (N_21970,N_21278,N_20522);
nand U21971 (N_21971,N_20592,N_20812);
nor U21972 (N_21972,N_21042,N_21116);
nand U21973 (N_21973,N_20917,N_21586);
xor U21974 (N_21974,N_21135,N_20808);
nor U21975 (N_21975,N_20578,N_20889);
xor U21976 (N_21976,N_20659,N_21530);
nor U21977 (N_21977,N_21540,N_20720);
or U21978 (N_21978,N_21364,N_21589);
nor U21979 (N_21979,N_20742,N_21048);
nand U21980 (N_21980,N_21140,N_20820);
or U21981 (N_21981,N_20655,N_20758);
nand U21982 (N_21982,N_20885,N_20495);
and U21983 (N_21983,N_20721,N_21420);
nor U21984 (N_21984,N_20404,N_20930);
xnor U21985 (N_21985,N_20725,N_20570);
and U21986 (N_21986,N_20492,N_20575);
and U21987 (N_21987,N_20688,N_20847);
and U21988 (N_21988,N_20945,N_20878);
and U21989 (N_21989,N_21299,N_21177);
nand U21990 (N_21990,N_21568,N_21039);
nand U21991 (N_21991,N_21332,N_21500);
nand U21992 (N_21992,N_20556,N_21564);
and U21993 (N_21993,N_20803,N_21360);
nor U21994 (N_21994,N_21112,N_21056);
and U21995 (N_21995,N_21247,N_20666);
nand U21996 (N_21996,N_20613,N_20929);
and U21997 (N_21997,N_20768,N_21480);
nor U21998 (N_21998,N_20877,N_21075);
or U21999 (N_21999,N_20672,N_20715);
or U22000 (N_22000,N_20579,N_20681);
or U22001 (N_22001,N_21598,N_21237);
nand U22002 (N_22002,N_20544,N_21554);
and U22003 (N_22003,N_21454,N_20620);
nor U22004 (N_22004,N_20836,N_20638);
xnor U22005 (N_22005,N_21506,N_21455);
or U22006 (N_22006,N_20852,N_21271);
nor U22007 (N_22007,N_21533,N_21559);
or U22008 (N_22008,N_21557,N_20515);
and U22009 (N_22009,N_20401,N_20509);
and U22010 (N_22010,N_21018,N_20828);
and U22011 (N_22011,N_20641,N_21230);
xor U22012 (N_22012,N_21019,N_20770);
nand U22013 (N_22013,N_21101,N_20589);
xor U22014 (N_22014,N_20423,N_20866);
nand U22015 (N_22015,N_21517,N_20839);
and U22016 (N_22016,N_21435,N_21144);
nor U22017 (N_22017,N_20595,N_21335);
xnor U22018 (N_22018,N_21323,N_21584);
nor U22019 (N_22019,N_20548,N_21502);
xor U22020 (N_22020,N_20815,N_21583);
xor U22021 (N_22021,N_20403,N_21150);
nand U22022 (N_22022,N_21548,N_21538);
or U22023 (N_22023,N_21109,N_21244);
nand U22024 (N_22024,N_21563,N_20987);
or U22025 (N_22025,N_21331,N_20748);
nor U22026 (N_22026,N_21234,N_20490);
xnor U22027 (N_22027,N_21145,N_21243);
or U22028 (N_22028,N_21585,N_21494);
or U22029 (N_22029,N_20464,N_21256);
xnor U22030 (N_22030,N_20737,N_20646);
nand U22031 (N_22031,N_20986,N_21155);
or U22032 (N_22032,N_21296,N_20691);
xnor U22033 (N_22033,N_20717,N_20441);
xnor U22034 (N_22034,N_21141,N_20443);
or U22035 (N_22035,N_21477,N_21594);
nand U22036 (N_22036,N_21117,N_20791);
and U22037 (N_22037,N_21595,N_21092);
xnor U22038 (N_22038,N_21396,N_21458);
or U22039 (N_22039,N_21401,N_20966);
and U22040 (N_22040,N_21217,N_20483);
or U22041 (N_22041,N_20705,N_20621);
or U22042 (N_22042,N_20922,N_20860);
xnor U22043 (N_22043,N_21188,N_21523);
xnor U22044 (N_22044,N_21547,N_21339);
nor U22045 (N_22045,N_20751,N_20974);
xnor U22046 (N_22046,N_20586,N_21515);
nor U22047 (N_22047,N_20874,N_20896);
or U22048 (N_22048,N_21099,N_21185);
and U22049 (N_22049,N_21446,N_20787);
or U22050 (N_22050,N_21562,N_20580);
or U22051 (N_22051,N_21330,N_20639);
or U22052 (N_22052,N_20491,N_20936);
or U22053 (N_22053,N_21599,N_21082);
and U22054 (N_22054,N_21388,N_20833);
xor U22055 (N_22055,N_21200,N_20437);
xor U22056 (N_22056,N_20414,N_20853);
nand U22057 (N_22057,N_21492,N_21225);
xor U22058 (N_22058,N_21415,N_21556);
nand U22059 (N_22059,N_21359,N_21485);
nand U22060 (N_22060,N_20741,N_20452);
xnor U22061 (N_22061,N_20904,N_20632);
xor U22062 (N_22062,N_20992,N_21448);
and U22063 (N_22063,N_20871,N_21134);
or U22064 (N_22064,N_21483,N_20883);
and U22065 (N_22065,N_21501,N_21066);
nor U22066 (N_22066,N_21016,N_20797);
nand U22067 (N_22067,N_20546,N_20498);
nand U22068 (N_22068,N_21353,N_20950);
xnor U22069 (N_22069,N_21041,N_20714);
nor U22070 (N_22070,N_20870,N_20973);
or U22071 (N_22071,N_20508,N_21440);
or U22072 (N_22072,N_21558,N_21250);
xor U22073 (N_22073,N_21071,N_21170);
and U22074 (N_22074,N_20732,N_21516);
nor U22075 (N_22075,N_21167,N_20824);
and U22076 (N_22076,N_20989,N_21186);
nor U22077 (N_22077,N_21580,N_20433);
or U22078 (N_22078,N_20980,N_21324);
or U22079 (N_22079,N_20600,N_20421);
xor U22080 (N_22080,N_21215,N_20501);
or U22081 (N_22081,N_20528,N_21431);
nand U22082 (N_22082,N_21321,N_20698);
xor U22083 (N_22083,N_21416,N_20585);
and U22084 (N_22084,N_20908,N_21008);
or U22085 (N_22085,N_20482,N_20668);
nand U22086 (N_22086,N_20756,N_20545);
nor U22087 (N_22087,N_20734,N_21046);
nand U22088 (N_22088,N_20444,N_21345);
or U22089 (N_22089,N_20859,N_20757);
and U22090 (N_22090,N_20459,N_21507);
or U22091 (N_22091,N_20474,N_21549);
nand U22092 (N_22092,N_21090,N_21114);
nor U22093 (N_22093,N_20420,N_21073);
and U22094 (N_22094,N_20829,N_21171);
and U22095 (N_22095,N_21094,N_20881);
or U22096 (N_22096,N_21083,N_21204);
nand U22097 (N_22097,N_21043,N_20743);
nor U22098 (N_22098,N_20826,N_20458);
or U22099 (N_22099,N_21035,N_20506);
and U22100 (N_22100,N_20902,N_20410);
nand U22101 (N_22101,N_21036,N_21463);
nor U22102 (N_22102,N_21095,N_20574);
and U22103 (N_22103,N_21524,N_20869);
xor U22104 (N_22104,N_21437,N_21399);
nor U22105 (N_22105,N_20796,N_21536);
or U22106 (N_22106,N_21527,N_21248);
and U22107 (N_22107,N_21024,N_20822);
and U22108 (N_22108,N_21306,N_21565);
and U22109 (N_22109,N_20415,N_21452);
nand U22110 (N_22110,N_20622,N_20933);
or U22111 (N_22111,N_21512,N_21165);
nor U22112 (N_22112,N_20463,N_21513);
or U22113 (N_22113,N_21113,N_20487);
xor U22114 (N_22114,N_21569,N_20739);
xor U22115 (N_22115,N_20841,N_21311);
xnor U22116 (N_22116,N_21228,N_20568);
xnor U22117 (N_22117,N_21295,N_21038);
or U22118 (N_22118,N_20716,N_20416);
nor U22119 (N_22119,N_20440,N_20775);
or U22120 (N_22120,N_21484,N_20827);
and U22121 (N_22121,N_20964,N_20605);
and U22122 (N_22122,N_21195,N_20801);
or U22123 (N_22123,N_21419,N_21253);
nor U22124 (N_22124,N_20450,N_20701);
and U22125 (N_22125,N_20502,N_21573);
nand U22126 (N_22126,N_20949,N_20723);
nand U22127 (N_22127,N_20814,N_20923);
xnor U22128 (N_22128,N_20614,N_20552);
nor U22129 (N_22129,N_20542,N_21207);
nor U22130 (N_22130,N_21575,N_21308);
xnor U22131 (N_22131,N_21597,N_20629);
and U22132 (N_22132,N_21334,N_21374);
and U22133 (N_22133,N_21013,N_21451);
or U22134 (N_22134,N_20940,N_20924);
nor U22135 (N_22135,N_20599,N_20561);
and U22136 (N_22136,N_20983,N_21449);
nand U22137 (N_22137,N_20857,N_21408);
nand U22138 (N_22138,N_20892,N_21443);
nor U22139 (N_22139,N_21336,N_20523);
nand U22140 (N_22140,N_20628,N_21289);
nor U22141 (N_22141,N_21545,N_21091);
and U22142 (N_22142,N_20784,N_20581);
xnor U22143 (N_22143,N_20825,N_20921);
or U22144 (N_22144,N_20783,N_20558);
and U22145 (N_22145,N_21210,N_20729);
or U22146 (N_22146,N_20727,N_21192);
xnor U22147 (N_22147,N_21119,N_20850);
or U22148 (N_22148,N_20596,N_21493);
nand U22149 (N_22149,N_21365,N_21078);
or U22150 (N_22150,N_21534,N_20643);
or U22151 (N_22151,N_21191,N_20689);
or U22152 (N_22152,N_20565,N_20875);
nor U22153 (N_22153,N_20862,N_21310);
and U22154 (N_22154,N_21481,N_20994);
nor U22155 (N_22155,N_20730,N_21229);
nor U22156 (N_22156,N_20731,N_21261);
and U22157 (N_22157,N_21491,N_21238);
and U22158 (N_22158,N_21529,N_20806);
xnor U22159 (N_22159,N_20486,N_20400);
nand U22160 (N_22160,N_20470,N_21055);
xor U22161 (N_22161,N_21023,N_20868);
and U22162 (N_22162,N_20436,N_20915);
xor U22163 (N_22163,N_20939,N_21383);
xnor U22164 (N_22164,N_21029,N_21532);
nand U22165 (N_22165,N_21139,N_20728);
nor U22166 (N_22166,N_20895,N_21058);
or U22167 (N_22167,N_20912,N_21505);
or U22168 (N_22168,N_20489,N_20573);
or U22169 (N_22169,N_21546,N_20603);
nor U22170 (N_22170,N_21445,N_20893);
nor U22171 (N_22171,N_21258,N_20594);
xnor U22172 (N_22172,N_21366,N_20843);
nor U22173 (N_22173,N_20541,N_20754);
nand U22174 (N_22174,N_20766,N_21274);
xor U22175 (N_22175,N_20656,N_20842);
nand U22176 (N_22176,N_21560,N_20408);
nor U22177 (N_22177,N_21403,N_20997);
or U22178 (N_22178,N_21438,N_21030);
xnor U22179 (N_22179,N_21428,N_20634);
nand U22180 (N_22180,N_20954,N_21232);
nor U22181 (N_22181,N_20914,N_21067);
nor U22182 (N_22182,N_20982,N_21341);
nor U22183 (N_22183,N_21476,N_21193);
nor U22184 (N_22184,N_20818,N_21175);
or U22185 (N_22185,N_21158,N_21002);
or U22186 (N_22186,N_20479,N_21221);
or U22187 (N_22187,N_20700,N_20652);
and U22188 (N_22188,N_21160,N_20569);
or U22189 (N_22189,N_20630,N_21375);
nor U22190 (N_22190,N_20527,N_21511);
xnor U22191 (N_22191,N_20707,N_20938);
nand U22192 (N_22192,N_20455,N_21395);
or U22193 (N_22193,N_20520,N_21327);
and U22194 (N_22194,N_20944,N_20649);
xor U22195 (N_22195,N_20449,N_20636);
nor U22196 (N_22196,N_21004,N_20514);
nor U22197 (N_22197,N_20468,N_21107);
xnor U22198 (N_22198,N_21142,N_20959);
nor U22199 (N_22199,N_20962,N_21453);
nand U22200 (N_22200,N_20901,N_20815);
or U22201 (N_22201,N_20487,N_20775);
or U22202 (N_22202,N_21286,N_20894);
xor U22203 (N_22203,N_21506,N_21149);
nor U22204 (N_22204,N_21412,N_20418);
xor U22205 (N_22205,N_20806,N_20963);
xnor U22206 (N_22206,N_21281,N_21476);
nand U22207 (N_22207,N_21349,N_20797);
nor U22208 (N_22208,N_20804,N_20935);
nor U22209 (N_22209,N_20555,N_21366);
nand U22210 (N_22210,N_20607,N_21549);
xnor U22211 (N_22211,N_20619,N_21346);
nand U22212 (N_22212,N_21570,N_21140);
or U22213 (N_22213,N_20421,N_20737);
nand U22214 (N_22214,N_20771,N_21063);
xor U22215 (N_22215,N_20592,N_20660);
and U22216 (N_22216,N_21133,N_20423);
or U22217 (N_22217,N_21024,N_21229);
nor U22218 (N_22218,N_20450,N_21021);
or U22219 (N_22219,N_21410,N_21502);
nand U22220 (N_22220,N_20952,N_20827);
nor U22221 (N_22221,N_21531,N_20536);
nor U22222 (N_22222,N_21464,N_20783);
nor U22223 (N_22223,N_21455,N_21532);
nand U22224 (N_22224,N_21592,N_20487);
xnor U22225 (N_22225,N_20433,N_20603);
xnor U22226 (N_22226,N_20478,N_20563);
xnor U22227 (N_22227,N_21367,N_20686);
or U22228 (N_22228,N_20945,N_20863);
xor U22229 (N_22229,N_21294,N_21537);
or U22230 (N_22230,N_20547,N_21297);
nor U22231 (N_22231,N_21214,N_20633);
nor U22232 (N_22232,N_20437,N_20822);
and U22233 (N_22233,N_21349,N_21193);
or U22234 (N_22234,N_20862,N_21366);
xor U22235 (N_22235,N_21165,N_20921);
nor U22236 (N_22236,N_21452,N_21294);
and U22237 (N_22237,N_21013,N_20640);
or U22238 (N_22238,N_21106,N_21017);
nor U22239 (N_22239,N_20899,N_20864);
xor U22240 (N_22240,N_20741,N_20669);
and U22241 (N_22241,N_21533,N_20412);
nand U22242 (N_22242,N_21572,N_21167);
or U22243 (N_22243,N_21139,N_20587);
nand U22244 (N_22244,N_20896,N_21280);
nand U22245 (N_22245,N_20817,N_20960);
xor U22246 (N_22246,N_21433,N_21146);
and U22247 (N_22247,N_20991,N_20894);
and U22248 (N_22248,N_21487,N_20769);
or U22249 (N_22249,N_21328,N_21001);
and U22250 (N_22250,N_21176,N_20748);
and U22251 (N_22251,N_21277,N_20744);
nand U22252 (N_22252,N_21114,N_21454);
or U22253 (N_22253,N_20908,N_20854);
and U22254 (N_22254,N_21195,N_20806);
nand U22255 (N_22255,N_21309,N_21412);
nand U22256 (N_22256,N_21001,N_20613);
xor U22257 (N_22257,N_20925,N_21067);
nand U22258 (N_22258,N_20805,N_21276);
xnor U22259 (N_22259,N_21529,N_20638);
xnor U22260 (N_22260,N_20404,N_21289);
or U22261 (N_22261,N_20769,N_21309);
or U22262 (N_22262,N_20701,N_20967);
nor U22263 (N_22263,N_21145,N_20562);
xnor U22264 (N_22264,N_20811,N_20563);
and U22265 (N_22265,N_21176,N_21303);
xnor U22266 (N_22266,N_21403,N_21006);
and U22267 (N_22267,N_20488,N_21098);
nand U22268 (N_22268,N_21435,N_20422);
or U22269 (N_22269,N_21128,N_20906);
and U22270 (N_22270,N_20639,N_21263);
and U22271 (N_22271,N_21107,N_21139);
and U22272 (N_22272,N_20976,N_21541);
and U22273 (N_22273,N_20416,N_21286);
or U22274 (N_22274,N_21237,N_21055);
nor U22275 (N_22275,N_20597,N_20835);
or U22276 (N_22276,N_21139,N_20438);
or U22277 (N_22277,N_20869,N_21127);
nor U22278 (N_22278,N_21251,N_20927);
nor U22279 (N_22279,N_20518,N_20769);
nor U22280 (N_22280,N_21242,N_20717);
nand U22281 (N_22281,N_20787,N_21253);
or U22282 (N_22282,N_21040,N_21540);
nand U22283 (N_22283,N_21265,N_21355);
and U22284 (N_22284,N_21334,N_21151);
nor U22285 (N_22285,N_21020,N_20700);
nand U22286 (N_22286,N_21445,N_21008);
xor U22287 (N_22287,N_21584,N_21361);
nor U22288 (N_22288,N_21009,N_21197);
nor U22289 (N_22289,N_20741,N_20618);
and U22290 (N_22290,N_20433,N_21137);
or U22291 (N_22291,N_20937,N_21207);
nand U22292 (N_22292,N_21141,N_20913);
nand U22293 (N_22293,N_20485,N_21534);
nand U22294 (N_22294,N_21413,N_21264);
and U22295 (N_22295,N_21007,N_21477);
and U22296 (N_22296,N_20955,N_20825);
and U22297 (N_22297,N_20714,N_20489);
nand U22298 (N_22298,N_21433,N_20553);
or U22299 (N_22299,N_21429,N_20618);
nand U22300 (N_22300,N_20584,N_20508);
nor U22301 (N_22301,N_21383,N_21187);
or U22302 (N_22302,N_20850,N_20600);
nand U22303 (N_22303,N_20933,N_20537);
and U22304 (N_22304,N_20400,N_20845);
or U22305 (N_22305,N_20507,N_20999);
xnor U22306 (N_22306,N_21330,N_21285);
and U22307 (N_22307,N_21159,N_21145);
nand U22308 (N_22308,N_21395,N_21061);
nor U22309 (N_22309,N_20943,N_20783);
nor U22310 (N_22310,N_20900,N_21448);
and U22311 (N_22311,N_20954,N_20665);
or U22312 (N_22312,N_21237,N_20854);
or U22313 (N_22313,N_21270,N_21182);
or U22314 (N_22314,N_21581,N_20883);
and U22315 (N_22315,N_21017,N_20693);
nor U22316 (N_22316,N_21594,N_21575);
and U22317 (N_22317,N_21329,N_20899);
nor U22318 (N_22318,N_20512,N_20968);
nor U22319 (N_22319,N_20712,N_20504);
xnor U22320 (N_22320,N_20829,N_21283);
xnor U22321 (N_22321,N_21307,N_20617);
and U22322 (N_22322,N_20465,N_21105);
and U22323 (N_22323,N_21295,N_21051);
or U22324 (N_22324,N_20904,N_20768);
xnor U22325 (N_22325,N_20421,N_20941);
or U22326 (N_22326,N_21378,N_21521);
or U22327 (N_22327,N_20951,N_21257);
nor U22328 (N_22328,N_21282,N_20411);
nand U22329 (N_22329,N_21342,N_21150);
nor U22330 (N_22330,N_20634,N_20735);
nor U22331 (N_22331,N_20706,N_20949);
nor U22332 (N_22332,N_21574,N_20464);
or U22333 (N_22333,N_21012,N_20727);
or U22334 (N_22334,N_20724,N_20659);
xnor U22335 (N_22335,N_21049,N_20449);
nor U22336 (N_22336,N_20979,N_21403);
xnor U22337 (N_22337,N_21068,N_20533);
or U22338 (N_22338,N_21093,N_20604);
nor U22339 (N_22339,N_21456,N_21049);
nand U22340 (N_22340,N_20511,N_20758);
or U22341 (N_22341,N_20433,N_21052);
or U22342 (N_22342,N_21034,N_20964);
nand U22343 (N_22343,N_20459,N_21143);
nand U22344 (N_22344,N_21553,N_20668);
nand U22345 (N_22345,N_21122,N_20567);
or U22346 (N_22346,N_21035,N_20727);
nor U22347 (N_22347,N_21004,N_20511);
and U22348 (N_22348,N_20515,N_20858);
nor U22349 (N_22349,N_20978,N_21141);
xnor U22350 (N_22350,N_21221,N_20489);
nand U22351 (N_22351,N_21304,N_20405);
or U22352 (N_22352,N_20671,N_21233);
nor U22353 (N_22353,N_20487,N_20810);
or U22354 (N_22354,N_20609,N_21040);
nor U22355 (N_22355,N_21296,N_21181);
xnor U22356 (N_22356,N_21391,N_21057);
or U22357 (N_22357,N_21273,N_21235);
nor U22358 (N_22358,N_21234,N_20876);
nor U22359 (N_22359,N_20544,N_20786);
nand U22360 (N_22360,N_21064,N_20610);
or U22361 (N_22361,N_20560,N_20725);
and U22362 (N_22362,N_20727,N_21189);
or U22363 (N_22363,N_20419,N_20868);
nor U22364 (N_22364,N_20589,N_20634);
nor U22365 (N_22365,N_20984,N_21171);
xor U22366 (N_22366,N_20581,N_21221);
nand U22367 (N_22367,N_21148,N_21460);
nand U22368 (N_22368,N_20866,N_21533);
and U22369 (N_22369,N_20994,N_21063);
nand U22370 (N_22370,N_21273,N_20918);
or U22371 (N_22371,N_20806,N_21534);
nor U22372 (N_22372,N_20661,N_21214);
or U22373 (N_22373,N_21493,N_21498);
nor U22374 (N_22374,N_20650,N_21298);
nor U22375 (N_22375,N_21139,N_20786);
and U22376 (N_22376,N_20507,N_20553);
nor U22377 (N_22377,N_20436,N_21548);
nand U22378 (N_22378,N_21411,N_20885);
nor U22379 (N_22379,N_21415,N_20685);
nor U22380 (N_22380,N_21077,N_21576);
or U22381 (N_22381,N_21288,N_20889);
or U22382 (N_22382,N_21035,N_20949);
nor U22383 (N_22383,N_21258,N_21326);
or U22384 (N_22384,N_21596,N_21288);
xnor U22385 (N_22385,N_20600,N_20987);
xnor U22386 (N_22386,N_20570,N_20448);
nor U22387 (N_22387,N_20641,N_21352);
and U22388 (N_22388,N_21541,N_20815);
xnor U22389 (N_22389,N_20834,N_20886);
nand U22390 (N_22390,N_20905,N_20543);
xnor U22391 (N_22391,N_20591,N_20756);
xnor U22392 (N_22392,N_20765,N_21459);
or U22393 (N_22393,N_20739,N_20870);
xnor U22394 (N_22394,N_21076,N_21599);
nor U22395 (N_22395,N_21050,N_20930);
xor U22396 (N_22396,N_21482,N_21010);
xor U22397 (N_22397,N_21437,N_20499);
xor U22398 (N_22398,N_20462,N_20718);
xnor U22399 (N_22399,N_21287,N_20462);
xor U22400 (N_22400,N_20760,N_21339);
and U22401 (N_22401,N_21539,N_21429);
nand U22402 (N_22402,N_20859,N_20936);
xor U22403 (N_22403,N_21166,N_20607);
xnor U22404 (N_22404,N_20536,N_21156);
or U22405 (N_22405,N_21266,N_21421);
nor U22406 (N_22406,N_21371,N_20971);
nand U22407 (N_22407,N_21552,N_20468);
xor U22408 (N_22408,N_21058,N_20784);
nand U22409 (N_22409,N_21031,N_20422);
xor U22410 (N_22410,N_20446,N_21577);
xnor U22411 (N_22411,N_21480,N_21461);
nor U22412 (N_22412,N_21565,N_21298);
and U22413 (N_22413,N_20570,N_20650);
nand U22414 (N_22414,N_21037,N_20675);
xnor U22415 (N_22415,N_20758,N_21198);
nand U22416 (N_22416,N_21505,N_20643);
nor U22417 (N_22417,N_21226,N_21091);
nor U22418 (N_22418,N_21498,N_21122);
nand U22419 (N_22419,N_21355,N_20941);
xor U22420 (N_22420,N_21562,N_21500);
nor U22421 (N_22421,N_20771,N_21099);
and U22422 (N_22422,N_21091,N_20638);
nand U22423 (N_22423,N_21597,N_21583);
nor U22424 (N_22424,N_21369,N_20540);
xor U22425 (N_22425,N_21565,N_21229);
nor U22426 (N_22426,N_20758,N_20709);
xor U22427 (N_22427,N_20561,N_20943);
nand U22428 (N_22428,N_21418,N_21276);
xnor U22429 (N_22429,N_20808,N_20941);
and U22430 (N_22430,N_20538,N_20828);
or U22431 (N_22431,N_21202,N_20555);
xnor U22432 (N_22432,N_21423,N_21057);
nor U22433 (N_22433,N_21546,N_20696);
xor U22434 (N_22434,N_21549,N_21512);
nand U22435 (N_22435,N_20827,N_20699);
and U22436 (N_22436,N_20445,N_21125);
xor U22437 (N_22437,N_20462,N_20776);
nand U22438 (N_22438,N_20476,N_20612);
and U22439 (N_22439,N_20960,N_21216);
nand U22440 (N_22440,N_21337,N_20907);
nand U22441 (N_22441,N_21568,N_21220);
xnor U22442 (N_22442,N_21206,N_20533);
nand U22443 (N_22443,N_20801,N_21562);
nor U22444 (N_22444,N_20750,N_20787);
nand U22445 (N_22445,N_21578,N_20462);
nor U22446 (N_22446,N_20905,N_20619);
and U22447 (N_22447,N_20842,N_21270);
nand U22448 (N_22448,N_20930,N_21446);
or U22449 (N_22449,N_20979,N_20996);
nor U22450 (N_22450,N_20420,N_20929);
nor U22451 (N_22451,N_21366,N_21382);
nand U22452 (N_22452,N_20833,N_21392);
nand U22453 (N_22453,N_20683,N_20857);
xnor U22454 (N_22454,N_21529,N_20807);
nor U22455 (N_22455,N_20415,N_20960);
nor U22456 (N_22456,N_20935,N_20794);
or U22457 (N_22457,N_20992,N_20714);
and U22458 (N_22458,N_21575,N_21037);
or U22459 (N_22459,N_20622,N_20607);
or U22460 (N_22460,N_20848,N_21202);
nand U22461 (N_22461,N_21531,N_20707);
nand U22462 (N_22462,N_20606,N_21187);
nand U22463 (N_22463,N_21198,N_21267);
xnor U22464 (N_22464,N_21179,N_20928);
xnor U22465 (N_22465,N_20593,N_20762);
xor U22466 (N_22466,N_20999,N_20790);
or U22467 (N_22467,N_20757,N_20768);
nand U22468 (N_22468,N_21507,N_20747);
nor U22469 (N_22469,N_21428,N_21450);
nand U22470 (N_22470,N_20631,N_21305);
or U22471 (N_22471,N_21009,N_21104);
or U22472 (N_22472,N_20589,N_21309);
xor U22473 (N_22473,N_20566,N_21172);
or U22474 (N_22474,N_20914,N_20915);
nor U22475 (N_22475,N_20889,N_21434);
xnor U22476 (N_22476,N_20803,N_20915);
or U22477 (N_22477,N_21120,N_21203);
xor U22478 (N_22478,N_21268,N_20522);
nor U22479 (N_22479,N_20581,N_20802);
and U22480 (N_22480,N_21165,N_20439);
nand U22481 (N_22481,N_21052,N_20502);
or U22482 (N_22482,N_21404,N_21282);
or U22483 (N_22483,N_20757,N_20927);
nand U22484 (N_22484,N_20906,N_21261);
and U22485 (N_22485,N_20665,N_21385);
xnor U22486 (N_22486,N_20801,N_21592);
nor U22487 (N_22487,N_21007,N_20465);
or U22488 (N_22488,N_21355,N_20992);
nor U22489 (N_22489,N_21454,N_21266);
xnor U22490 (N_22490,N_21590,N_21075);
xor U22491 (N_22491,N_21328,N_21222);
nand U22492 (N_22492,N_20654,N_21555);
and U22493 (N_22493,N_21294,N_21163);
xnor U22494 (N_22494,N_21142,N_21061);
or U22495 (N_22495,N_21349,N_21508);
or U22496 (N_22496,N_20756,N_21521);
xnor U22497 (N_22497,N_20575,N_21415);
xnor U22498 (N_22498,N_21079,N_20892);
nor U22499 (N_22499,N_21299,N_21233);
or U22500 (N_22500,N_20726,N_20401);
nand U22501 (N_22501,N_21178,N_20604);
or U22502 (N_22502,N_20961,N_20474);
or U22503 (N_22503,N_20612,N_21125);
nand U22504 (N_22504,N_20707,N_21497);
and U22505 (N_22505,N_21290,N_20866);
nand U22506 (N_22506,N_21484,N_21300);
nand U22507 (N_22507,N_20428,N_21564);
xor U22508 (N_22508,N_21322,N_21477);
xnor U22509 (N_22509,N_21061,N_20909);
and U22510 (N_22510,N_20860,N_20479);
xor U22511 (N_22511,N_20490,N_21145);
xor U22512 (N_22512,N_20584,N_21559);
and U22513 (N_22513,N_21205,N_20545);
nor U22514 (N_22514,N_21323,N_21407);
and U22515 (N_22515,N_20691,N_21455);
xnor U22516 (N_22516,N_21117,N_21030);
nor U22517 (N_22517,N_20445,N_20413);
and U22518 (N_22518,N_20962,N_20799);
nor U22519 (N_22519,N_21511,N_20441);
or U22520 (N_22520,N_20591,N_20858);
xor U22521 (N_22521,N_21066,N_21116);
nand U22522 (N_22522,N_20811,N_20822);
and U22523 (N_22523,N_21199,N_20419);
or U22524 (N_22524,N_21045,N_21526);
or U22525 (N_22525,N_21213,N_21391);
xnor U22526 (N_22526,N_20618,N_20951);
xor U22527 (N_22527,N_20578,N_21377);
xor U22528 (N_22528,N_20872,N_21134);
nand U22529 (N_22529,N_21299,N_20835);
and U22530 (N_22530,N_20954,N_21149);
and U22531 (N_22531,N_21326,N_21304);
and U22532 (N_22532,N_20777,N_21176);
nor U22533 (N_22533,N_21443,N_20407);
nand U22534 (N_22534,N_20483,N_20896);
or U22535 (N_22535,N_20476,N_20848);
nor U22536 (N_22536,N_20743,N_20502);
and U22537 (N_22537,N_21042,N_21184);
nor U22538 (N_22538,N_21471,N_21120);
or U22539 (N_22539,N_20580,N_21554);
nor U22540 (N_22540,N_21444,N_20817);
nor U22541 (N_22541,N_21299,N_20637);
and U22542 (N_22542,N_20653,N_21047);
nor U22543 (N_22543,N_21556,N_20522);
or U22544 (N_22544,N_21353,N_21122);
or U22545 (N_22545,N_20564,N_21341);
and U22546 (N_22546,N_21005,N_20468);
xnor U22547 (N_22547,N_20646,N_20722);
and U22548 (N_22548,N_20543,N_20588);
xnor U22549 (N_22549,N_20665,N_21394);
nor U22550 (N_22550,N_20470,N_20618);
or U22551 (N_22551,N_21591,N_21190);
nor U22552 (N_22552,N_20829,N_20709);
xnor U22553 (N_22553,N_20635,N_21251);
xor U22554 (N_22554,N_20918,N_21144);
xor U22555 (N_22555,N_21288,N_20408);
nor U22556 (N_22556,N_20934,N_21247);
or U22557 (N_22557,N_20676,N_21223);
nand U22558 (N_22558,N_21296,N_21348);
or U22559 (N_22559,N_20968,N_20896);
and U22560 (N_22560,N_21481,N_21297);
nor U22561 (N_22561,N_20578,N_20760);
or U22562 (N_22562,N_20761,N_21592);
xnor U22563 (N_22563,N_20559,N_21120);
xnor U22564 (N_22564,N_20438,N_21021);
and U22565 (N_22565,N_20577,N_21513);
and U22566 (N_22566,N_21540,N_20840);
nor U22567 (N_22567,N_20595,N_20921);
nand U22568 (N_22568,N_20586,N_21045);
nor U22569 (N_22569,N_21010,N_20972);
xor U22570 (N_22570,N_20689,N_20447);
nand U22571 (N_22571,N_20625,N_20520);
and U22572 (N_22572,N_20989,N_20909);
nand U22573 (N_22573,N_21597,N_21485);
nand U22574 (N_22574,N_20726,N_21316);
nor U22575 (N_22575,N_21429,N_20886);
nand U22576 (N_22576,N_21502,N_21176);
or U22577 (N_22577,N_20569,N_21311);
and U22578 (N_22578,N_20856,N_21142);
and U22579 (N_22579,N_21220,N_21593);
nand U22580 (N_22580,N_20864,N_21211);
nand U22581 (N_22581,N_20759,N_20672);
nand U22582 (N_22582,N_21318,N_20494);
nand U22583 (N_22583,N_20605,N_21208);
nor U22584 (N_22584,N_20622,N_21237);
xor U22585 (N_22585,N_20844,N_21158);
or U22586 (N_22586,N_20653,N_20887);
or U22587 (N_22587,N_20424,N_20560);
nand U22588 (N_22588,N_20500,N_21396);
or U22589 (N_22589,N_20977,N_20532);
nor U22590 (N_22590,N_20847,N_20425);
and U22591 (N_22591,N_21200,N_21590);
nand U22592 (N_22592,N_21487,N_21515);
xnor U22593 (N_22593,N_21459,N_21134);
and U22594 (N_22594,N_20742,N_21369);
nor U22595 (N_22595,N_21166,N_21196);
xnor U22596 (N_22596,N_20862,N_21417);
and U22597 (N_22597,N_20791,N_21412);
or U22598 (N_22598,N_21186,N_20498);
nor U22599 (N_22599,N_20709,N_21246);
or U22600 (N_22600,N_21445,N_21429);
nand U22601 (N_22601,N_20402,N_21033);
nor U22602 (N_22602,N_21278,N_21365);
or U22603 (N_22603,N_21149,N_21189);
xnor U22604 (N_22604,N_20825,N_20929);
xnor U22605 (N_22605,N_20795,N_21104);
and U22606 (N_22606,N_20491,N_20769);
nor U22607 (N_22607,N_20835,N_21156);
and U22608 (N_22608,N_21007,N_21211);
or U22609 (N_22609,N_21594,N_21312);
nor U22610 (N_22610,N_20754,N_20464);
nand U22611 (N_22611,N_20575,N_21456);
xor U22612 (N_22612,N_20422,N_21373);
xor U22613 (N_22613,N_21375,N_21517);
and U22614 (N_22614,N_21297,N_21281);
nor U22615 (N_22615,N_21267,N_21294);
nand U22616 (N_22616,N_21497,N_21522);
or U22617 (N_22617,N_21371,N_21199);
and U22618 (N_22618,N_20756,N_20514);
nand U22619 (N_22619,N_20720,N_21127);
nand U22620 (N_22620,N_21292,N_21545);
or U22621 (N_22621,N_20961,N_21189);
or U22622 (N_22622,N_21295,N_20422);
xor U22623 (N_22623,N_20690,N_21019);
xnor U22624 (N_22624,N_21495,N_21308);
nand U22625 (N_22625,N_20749,N_20463);
nor U22626 (N_22626,N_20951,N_20459);
nand U22627 (N_22627,N_20819,N_20626);
and U22628 (N_22628,N_20493,N_21474);
nor U22629 (N_22629,N_20726,N_20722);
nand U22630 (N_22630,N_20559,N_20868);
and U22631 (N_22631,N_20848,N_21384);
and U22632 (N_22632,N_21577,N_20949);
nor U22633 (N_22633,N_20621,N_20997);
nand U22634 (N_22634,N_21485,N_21051);
or U22635 (N_22635,N_21528,N_20867);
and U22636 (N_22636,N_20677,N_21512);
and U22637 (N_22637,N_21361,N_21043);
and U22638 (N_22638,N_20930,N_21304);
xnor U22639 (N_22639,N_21376,N_20869);
nand U22640 (N_22640,N_21211,N_21048);
xnor U22641 (N_22641,N_20995,N_20973);
nand U22642 (N_22642,N_21149,N_21477);
nand U22643 (N_22643,N_21399,N_20865);
nand U22644 (N_22644,N_20694,N_21000);
or U22645 (N_22645,N_20554,N_21182);
or U22646 (N_22646,N_21404,N_20580);
or U22647 (N_22647,N_21124,N_20906);
nor U22648 (N_22648,N_21080,N_21049);
nor U22649 (N_22649,N_20731,N_20641);
nand U22650 (N_22650,N_20548,N_21139);
and U22651 (N_22651,N_21042,N_21066);
nor U22652 (N_22652,N_20726,N_21147);
or U22653 (N_22653,N_20701,N_20796);
nor U22654 (N_22654,N_21038,N_21560);
nand U22655 (N_22655,N_21577,N_21130);
and U22656 (N_22656,N_20668,N_21353);
nand U22657 (N_22657,N_20898,N_21330);
or U22658 (N_22658,N_21413,N_21572);
xnor U22659 (N_22659,N_20628,N_21516);
nor U22660 (N_22660,N_21262,N_21026);
and U22661 (N_22661,N_20716,N_20903);
nor U22662 (N_22662,N_21498,N_21438);
nand U22663 (N_22663,N_21378,N_20684);
nand U22664 (N_22664,N_20735,N_21114);
and U22665 (N_22665,N_20704,N_20822);
or U22666 (N_22666,N_20853,N_20766);
and U22667 (N_22667,N_21226,N_20686);
or U22668 (N_22668,N_21351,N_21414);
nand U22669 (N_22669,N_21037,N_20658);
nor U22670 (N_22670,N_20457,N_21543);
nand U22671 (N_22671,N_20616,N_20510);
nand U22672 (N_22672,N_20611,N_20470);
xor U22673 (N_22673,N_21137,N_21414);
nor U22674 (N_22674,N_20530,N_20737);
nor U22675 (N_22675,N_20752,N_21284);
nand U22676 (N_22676,N_21455,N_20879);
xnor U22677 (N_22677,N_21191,N_21425);
or U22678 (N_22678,N_20962,N_21338);
or U22679 (N_22679,N_21343,N_21324);
and U22680 (N_22680,N_21597,N_21564);
nand U22681 (N_22681,N_20425,N_21191);
and U22682 (N_22682,N_20610,N_21148);
xnor U22683 (N_22683,N_20664,N_21258);
nor U22684 (N_22684,N_20572,N_21117);
and U22685 (N_22685,N_20829,N_21059);
xor U22686 (N_22686,N_20482,N_20576);
and U22687 (N_22687,N_21364,N_21388);
and U22688 (N_22688,N_20913,N_20844);
nor U22689 (N_22689,N_21378,N_20808);
xnor U22690 (N_22690,N_20783,N_21154);
nor U22691 (N_22691,N_20771,N_21033);
and U22692 (N_22692,N_20997,N_21011);
nand U22693 (N_22693,N_21159,N_21421);
nand U22694 (N_22694,N_20474,N_21502);
and U22695 (N_22695,N_21194,N_20638);
nand U22696 (N_22696,N_21142,N_21054);
nor U22697 (N_22697,N_20443,N_20447);
or U22698 (N_22698,N_21111,N_21109);
xor U22699 (N_22699,N_20968,N_21101);
and U22700 (N_22700,N_21114,N_21598);
and U22701 (N_22701,N_20994,N_21052);
nand U22702 (N_22702,N_21047,N_20808);
nor U22703 (N_22703,N_20575,N_21584);
xnor U22704 (N_22704,N_20954,N_20969);
nand U22705 (N_22705,N_20669,N_21454);
nand U22706 (N_22706,N_21094,N_21219);
nor U22707 (N_22707,N_21137,N_20961);
and U22708 (N_22708,N_21384,N_20611);
xnor U22709 (N_22709,N_20930,N_21209);
or U22710 (N_22710,N_20645,N_20640);
and U22711 (N_22711,N_20964,N_21548);
nor U22712 (N_22712,N_20841,N_21386);
or U22713 (N_22713,N_20680,N_20475);
xor U22714 (N_22714,N_20583,N_21483);
and U22715 (N_22715,N_20728,N_20478);
xnor U22716 (N_22716,N_21086,N_21249);
and U22717 (N_22717,N_21364,N_21564);
or U22718 (N_22718,N_20703,N_21220);
and U22719 (N_22719,N_20630,N_21454);
xnor U22720 (N_22720,N_21360,N_21471);
and U22721 (N_22721,N_20969,N_21472);
and U22722 (N_22722,N_21432,N_20593);
and U22723 (N_22723,N_20615,N_21088);
nor U22724 (N_22724,N_20789,N_21288);
and U22725 (N_22725,N_20852,N_21203);
nor U22726 (N_22726,N_20931,N_21324);
nand U22727 (N_22727,N_20659,N_21225);
nand U22728 (N_22728,N_20912,N_21424);
nand U22729 (N_22729,N_21101,N_21008);
or U22730 (N_22730,N_21090,N_21358);
and U22731 (N_22731,N_20517,N_21470);
nand U22732 (N_22732,N_21201,N_21120);
nor U22733 (N_22733,N_20647,N_21259);
xor U22734 (N_22734,N_21392,N_20417);
nand U22735 (N_22735,N_20730,N_21452);
and U22736 (N_22736,N_20444,N_21091);
and U22737 (N_22737,N_20442,N_21443);
nor U22738 (N_22738,N_21139,N_21396);
xnor U22739 (N_22739,N_20522,N_20828);
and U22740 (N_22740,N_20489,N_21534);
nor U22741 (N_22741,N_21524,N_21363);
nor U22742 (N_22742,N_21415,N_21259);
xnor U22743 (N_22743,N_20820,N_21288);
and U22744 (N_22744,N_20632,N_21381);
nor U22745 (N_22745,N_20736,N_20773);
nor U22746 (N_22746,N_21124,N_20997);
nand U22747 (N_22747,N_21326,N_21558);
or U22748 (N_22748,N_20574,N_21323);
xnor U22749 (N_22749,N_21096,N_21065);
nor U22750 (N_22750,N_20846,N_20614);
or U22751 (N_22751,N_21024,N_21578);
xnor U22752 (N_22752,N_20879,N_20608);
or U22753 (N_22753,N_20755,N_20400);
nand U22754 (N_22754,N_20897,N_20800);
nor U22755 (N_22755,N_21117,N_21011);
nor U22756 (N_22756,N_20700,N_21081);
nor U22757 (N_22757,N_20837,N_20523);
nor U22758 (N_22758,N_20434,N_21224);
and U22759 (N_22759,N_21292,N_21024);
and U22760 (N_22760,N_21400,N_21044);
or U22761 (N_22761,N_20737,N_21465);
nor U22762 (N_22762,N_20486,N_20432);
xnor U22763 (N_22763,N_21422,N_20441);
nor U22764 (N_22764,N_21027,N_21427);
and U22765 (N_22765,N_20519,N_20835);
nor U22766 (N_22766,N_20477,N_21425);
and U22767 (N_22767,N_20540,N_21532);
nand U22768 (N_22768,N_20743,N_20429);
nor U22769 (N_22769,N_21125,N_21250);
nand U22770 (N_22770,N_20966,N_20631);
nor U22771 (N_22771,N_21006,N_20857);
nor U22772 (N_22772,N_21501,N_21489);
and U22773 (N_22773,N_20474,N_21224);
nor U22774 (N_22774,N_21363,N_21193);
or U22775 (N_22775,N_20507,N_21149);
nand U22776 (N_22776,N_20514,N_21207);
xnor U22777 (N_22777,N_21080,N_21287);
and U22778 (N_22778,N_20643,N_21209);
or U22779 (N_22779,N_21071,N_21290);
nor U22780 (N_22780,N_21350,N_20702);
and U22781 (N_22781,N_21240,N_20817);
nor U22782 (N_22782,N_20800,N_20408);
nand U22783 (N_22783,N_21502,N_20431);
and U22784 (N_22784,N_21569,N_21060);
nor U22785 (N_22785,N_20694,N_20936);
nor U22786 (N_22786,N_20581,N_21522);
nand U22787 (N_22787,N_20892,N_21182);
or U22788 (N_22788,N_20824,N_20435);
or U22789 (N_22789,N_21191,N_20485);
nor U22790 (N_22790,N_21538,N_20839);
xor U22791 (N_22791,N_21243,N_20469);
and U22792 (N_22792,N_21220,N_20518);
and U22793 (N_22793,N_21119,N_20611);
nor U22794 (N_22794,N_20948,N_20961);
nand U22795 (N_22795,N_21580,N_21174);
nand U22796 (N_22796,N_20856,N_21035);
nor U22797 (N_22797,N_21214,N_20895);
nand U22798 (N_22798,N_20902,N_21442);
and U22799 (N_22799,N_20430,N_21019);
nand U22800 (N_22800,N_21765,N_22299);
or U22801 (N_22801,N_22111,N_22118);
nand U22802 (N_22802,N_21608,N_22215);
nor U22803 (N_22803,N_22202,N_22098);
nor U22804 (N_22804,N_21768,N_22570);
xnor U22805 (N_22805,N_21607,N_22546);
and U22806 (N_22806,N_21813,N_22131);
nand U22807 (N_22807,N_22372,N_21628);
xor U22808 (N_22808,N_21746,N_22268);
nand U22809 (N_22809,N_22148,N_21759);
nand U22810 (N_22810,N_22719,N_21641);
nand U22811 (N_22811,N_22089,N_22124);
or U22812 (N_22812,N_22047,N_22500);
and U22813 (N_22813,N_22613,N_21685);
xnor U22814 (N_22814,N_22312,N_22244);
and U22815 (N_22815,N_22397,N_22537);
or U22816 (N_22816,N_22127,N_22316);
and U22817 (N_22817,N_22125,N_22555);
xor U22818 (N_22818,N_21664,N_21832);
and U22819 (N_22819,N_22723,N_22349);
and U22820 (N_22820,N_22661,N_22487);
or U22821 (N_22821,N_22416,N_22797);
nor U22822 (N_22822,N_21748,N_22001);
and U22823 (N_22823,N_22593,N_22757);
nand U22824 (N_22824,N_21842,N_21870);
or U22825 (N_22825,N_22647,N_22581);
or U22826 (N_22826,N_22144,N_22600);
xor U22827 (N_22827,N_22674,N_22366);
and U22828 (N_22828,N_22548,N_22446);
or U22829 (N_22829,N_22778,N_22524);
and U22830 (N_22830,N_22032,N_21899);
or U22831 (N_22831,N_22338,N_22146);
nand U22832 (N_22832,N_22550,N_22116);
xnor U22833 (N_22833,N_22174,N_22136);
xor U22834 (N_22834,N_21881,N_21882);
nand U22835 (N_22835,N_21939,N_22567);
nor U22836 (N_22836,N_21704,N_22642);
nor U22837 (N_22837,N_21979,N_22354);
xnor U22838 (N_22838,N_22405,N_21609);
nand U22839 (N_22839,N_22605,N_22790);
xor U22840 (N_22840,N_22568,N_22387);
and U22841 (N_22841,N_22679,N_22743);
nor U22842 (N_22842,N_21643,N_22308);
nand U22843 (N_22843,N_21820,N_21804);
or U22844 (N_22844,N_22603,N_21604);
nor U22845 (N_22845,N_22331,N_22523);
or U22846 (N_22846,N_22208,N_22761);
nand U22847 (N_22847,N_22102,N_21960);
xnor U22848 (N_22848,N_22415,N_21869);
and U22849 (N_22849,N_21717,N_22254);
and U22850 (N_22850,N_22715,N_21743);
or U22851 (N_22851,N_22334,N_22158);
xnor U22852 (N_22852,N_21922,N_22495);
nand U22853 (N_22853,N_22189,N_21896);
and U22854 (N_22854,N_21834,N_22027);
nand U22855 (N_22855,N_22077,N_22453);
nor U22856 (N_22856,N_22191,N_22310);
xnor U22857 (N_22857,N_22736,N_22403);
nand U22858 (N_22858,N_22211,N_22115);
xor U22859 (N_22859,N_21699,N_21790);
nand U22860 (N_22860,N_21634,N_22544);
or U22861 (N_22861,N_22237,N_21885);
nor U22862 (N_22862,N_22409,N_22141);
nor U22863 (N_22863,N_22344,N_22503);
nor U22864 (N_22864,N_21942,N_21655);
xor U22865 (N_22865,N_22720,N_22060);
xnor U22866 (N_22866,N_21758,N_22579);
or U22867 (N_22867,N_22440,N_21658);
and U22868 (N_22868,N_22765,N_22560);
and U22869 (N_22869,N_21889,N_22363);
nor U22870 (N_22870,N_21769,N_22439);
and U22871 (N_22871,N_22696,N_21721);
nor U22872 (N_22872,N_22175,N_21877);
nand U22873 (N_22873,N_22539,N_22396);
or U22874 (N_22874,N_21781,N_22669);
or U22875 (N_22875,N_22304,N_21990);
or U22876 (N_22876,N_21940,N_21991);
xnor U22877 (N_22877,N_22655,N_22004);
xnor U22878 (N_22878,N_22713,N_22701);
nor U22879 (N_22879,N_22194,N_22074);
and U22880 (N_22880,N_22041,N_22585);
nor U22881 (N_22881,N_21610,N_21989);
nand U22882 (N_22882,N_21849,N_22143);
xnor U22883 (N_22883,N_22418,N_22520);
nor U22884 (N_22884,N_21876,N_22261);
or U22885 (N_22885,N_21963,N_22139);
xor U22886 (N_22886,N_21716,N_21733);
xor U22887 (N_22887,N_22119,N_22658);
and U22888 (N_22888,N_22741,N_22172);
nand U22889 (N_22889,N_21841,N_22055);
xor U22890 (N_22890,N_22619,N_22085);
nor U22891 (N_22891,N_21632,N_21888);
xor U22892 (N_22892,N_21946,N_22109);
nand U22893 (N_22893,N_22219,N_22683);
and U22894 (N_22894,N_22775,N_21648);
or U22895 (N_22895,N_21647,N_22288);
or U22896 (N_22896,N_21949,N_21833);
and U22897 (N_22897,N_22725,N_22580);
nand U22898 (N_22898,N_22637,N_22161);
or U22899 (N_22899,N_22315,N_22514);
nand U22900 (N_22900,N_21915,N_22404);
nand U22901 (N_22901,N_22681,N_21660);
xor U22902 (N_22902,N_22362,N_22230);
nand U22903 (N_22903,N_22216,N_22650);
or U22904 (N_22904,N_22005,N_22267);
xor U22905 (N_22905,N_21958,N_21972);
and U22906 (N_22906,N_22424,N_22097);
xnor U22907 (N_22907,N_22430,N_21627);
xnor U22908 (N_22908,N_22527,N_22739);
nand U22909 (N_22909,N_21779,N_21677);
nand U22910 (N_22910,N_22648,N_22697);
or U22911 (N_22911,N_21747,N_22229);
nor U22912 (N_22912,N_22384,N_22760);
and U22913 (N_22913,N_21909,N_22086);
or U22914 (N_22914,N_22375,N_21763);
nor U22915 (N_22915,N_22153,N_21966);
or U22916 (N_22916,N_22785,N_22223);
nand U22917 (N_22917,N_22121,N_22263);
nand U22918 (N_22918,N_21858,N_21892);
or U22919 (N_22919,N_22457,N_22318);
and U22920 (N_22920,N_22103,N_21616);
and U22921 (N_22921,N_22100,N_22105);
nand U22922 (N_22922,N_22203,N_21734);
xor U22923 (N_22923,N_22638,N_21709);
and U22924 (N_22924,N_22058,N_22438);
nor U22925 (N_22925,N_22162,N_22793);
nand U22926 (N_22926,N_22134,N_21749);
and U22927 (N_22927,N_22664,N_21937);
nor U22928 (N_22928,N_22623,N_21667);
and U22929 (N_22929,N_21917,N_22649);
xor U22930 (N_22930,N_22682,N_21735);
nor U22931 (N_22931,N_22030,N_21726);
and U22932 (N_22932,N_22584,N_22531);
or U22933 (N_22933,N_22050,N_22536);
nand U22934 (N_22934,N_22122,N_21950);
xor U22935 (N_22935,N_22395,N_22678);
xor U22936 (N_22936,N_22467,N_21874);
nand U22937 (N_22937,N_22522,N_21819);
nor U22938 (N_22938,N_22505,N_22294);
xor U22939 (N_22939,N_22196,N_22615);
xor U22940 (N_22940,N_22573,N_22411);
nand U22941 (N_22941,N_22087,N_22535);
nor U22942 (N_22942,N_22571,N_22693);
nor U22943 (N_22943,N_21943,N_21902);
xnor U22944 (N_22944,N_21783,N_22708);
and U22945 (N_22945,N_22408,N_22456);
and U22946 (N_22946,N_22184,N_22703);
nand U22947 (N_22947,N_22167,N_21736);
and U22948 (N_22948,N_21812,N_22243);
nor U22949 (N_22949,N_22242,N_21645);
and U22950 (N_22950,N_21626,N_21875);
or U22951 (N_22951,N_22156,N_21934);
nor U22952 (N_22952,N_22322,N_22429);
or U22953 (N_22953,N_22225,N_22721);
and U22954 (N_22954,N_22663,N_22474);
or U22955 (N_22955,N_22553,N_22400);
nand U22956 (N_22956,N_22667,N_21983);
nand U22957 (N_22957,N_22788,N_22427);
nor U22958 (N_22958,N_22026,N_22513);
nor U22959 (N_22959,N_22508,N_22690);
or U22960 (N_22960,N_22258,N_21797);
or U22961 (N_22961,N_22099,N_22486);
and U22962 (N_22962,N_21775,N_21618);
and U22963 (N_22963,N_22677,N_21708);
nor U22964 (N_22964,N_21864,N_21811);
and U22965 (N_22965,N_22543,N_22231);
nand U22966 (N_22966,N_22149,N_22750);
nand U22967 (N_22967,N_22478,N_21690);
xnor U22968 (N_22968,N_21929,N_21800);
and U22969 (N_22969,N_22443,N_22067);
and U22970 (N_22970,N_21831,N_22330);
xnor U22971 (N_22971,N_21612,N_22120);
nor U22972 (N_22972,N_22779,N_21810);
xnor U22973 (N_22973,N_21851,N_22406);
or U22974 (N_22974,N_21984,N_21697);
xnor U22975 (N_22975,N_22364,N_22062);
nand U22976 (N_22976,N_21964,N_22606);
xor U22977 (N_22977,N_21745,N_22024);
nor U22978 (N_22978,N_22186,N_21906);
nand U22979 (N_22979,N_21682,N_22510);
nand U22980 (N_22980,N_21680,N_22738);
nor U22981 (N_22981,N_22042,N_22525);
nor U22982 (N_22982,N_21826,N_21818);
or U22983 (N_22983,N_22670,N_21706);
and U22984 (N_22984,N_22528,N_22783);
and U22985 (N_22985,N_21995,N_22489);
nor U22986 (N_22986,N_22079,N_21657);
nor U22987 (N_22987,N_22680,N_21982);
or U22988 (N_22988,N_22140,N_21794);
nand U22989 (N_22989,N_21844,N_22031);
nor U22990 (N_22990,N_22691,N_21924);
and U22991 (N_22991,N_22700,N_21956);
and U22992 (N_22992,N_22711,N_22176);
nor U22993 (N_22993,N_22755,N_22671);
nand U22994 (N_22994,N_21730,N_22620);
and U22995 (N_22995,N_21878,N_22376);
nor U22996 (N_22996,N_22442,N_22034);
and U22997 (N_22997,N_22730,N_22051);
and U22998 (N_22998,N_22594,N_22292);
nor U22999 (N_22999,N_22740,N_21622);
nand U23000 (N_23000,N_22183,N_21791);
and U23001 (N_23001,N_22534,N_22274);
or U23002 (N_23002,N_21640,N_22273);
nor U23003 (N_23003,N_22745,N_22130);
nor U23004 (N_23004,N_22044,N_21923);
nand U23005 (N_23005,N_22076,N_22325);
xor U23006 (N_23006,N_22236,N_21969);
or U23007 (N_23007,N_22106,N_21776);
nand U23008 (N_23008,N_22205,N_21911);
xnor U23009 (N_23009,N_22417,N_22306);
or U23010 (N_23010,N_22113,N_21705);
nand U23011 (N_23011,N_21980,N_22784);
or U23012 (N_23012,N_22652,N_22068);
xnor U23013 (N_23013,N_21862,N_22129);
and U23014 (N_23014,N_22504,N_21863);
nand U23015 (N_23015,N_22052,N_22643);
nor U23016 (N_23016,N_22083,N_22596);
or U23017 (N_23017,N_21649,N_22270);
and U23018 (N_23018,N_21836,N_21828);
xor U23019 (N_23019,N_22073,N_22455);
or U23020 (N_23020,N_22163,N_22179);
nand U23021 (N_23021,N_22588,N_22762);
nor U23022 (N_23022,N_22450,N_22475);
nor U23023 (N_23023,N_22393,N_22155);
xnor U23024 (N_23024,N_22187,N_22493);
xor U23025 (N_23025,N_21996,N_22590);
nand U23026 (N_23026,N_22591,N_21687);
and U23027 (N_23027,N_21968,N_22729);
or U23028 (N_23028,N_22684,N_22782);
nand U23029 (N_23029,N_22000,N_22481);
and U23030 (N_23030,N_22759,N_22198);
or U23031 (N_23031,N_22253,N_21739);
xnor U23032 (N_23032,N_21824,N_22688);
xor U23033 (N_23033,N_21865,N_22726);
or U23034 (N_23034,N_22469,N_22309);
xor U23035 (N_23035,N_22046,N_22718);
and U23036 (N_23036,N_22353,N_22252);
and U23037 (N_23037,N_22123,N_21886);
xor U23038 (N_23038,N_21668,N_22259);
and U23039 (N_23039,N_21852,N_22464);
and U23040 (N_23040,N_21676,N_22574);
or U23041 (N_23041,N_22488,N_21977);
nand U23042 (N_23042,N_22282,N_22399);
nand U23043 (N_23043,N_22559,N_22714);
or U23044 (N_23044,N_22329,N_21957);
xnor U23045 (N_23045,N_22337,N_21941);
and U23046 (N_23046,N_22777,N_22006);
nand U23047 (N_23047,N_21930,N_22297);
nor U23048 (N_23048,N_21861,N_22742);
nand U23049 (N_23049,N_22212,N_22275);
nor U23050 (N_23050,N_22063,N_22771);
nand U23051 (N_23051,N_21838,N_21859);
or U23052 (N_23052,N_22214,N_22343);
xor U23053 (N_23053,N_21952,N_21920);
nor U23054 (N_23054,N_22003,N_22114);
and U23055 (N_23055,N_21879,N_22151);
and U23056 (N_23056,N_21637,N_22040);
nand U23057 (N_23057,N_22561,N_22311);
nand U23058 (N_23058,N_22369,N_21827);
or U23059 (N_23059,N_22689,N_22358);
or U23060 (N_23060,N_22728,N_21808);
nor U23061 (N_23061,N_22350,N_22497);
xnor U23062 (N_23062,N_22694,N_22080);
xnor U23063 (N_23063,N_22698,N_21633);
and U23064 (N_23064,N_22445,N_21650);
or U23065 (N_23065,N_22007,N_22668);
nor U23066 (N_23066,N_22036,N_21893);
xor U23067 (N_23067,N_21900,N_21724);
or U23068 (N_23068,N_22356,N_21914);
nand U23069 (N_23069,N_22324,N_22220);
or U23070 (N_23070,N_22673,N_22084);
nor U23071 (N_23071,N_21830,N_22257);
xor U23072 (N_23072,N_21729,N_22029);
xnor U23073 (N_23073,N_22465,N_21789);
xnor U23074 (N_23074,N_21787,N_22626);
xor U23075 (N_23075,N_22152,N_22296);
or U23076 (N_23076,N_21688,N_22075);
and U23077 (N_23077,N_22507,N_22160);
nor U23078 (N_23078,N_22379,N_22323);
xnor U23079 (N_23079,N_22422,N_21727);
xnor U23080 (N_23080,N_21635,N_21883);
and U23081 (N_23081,N_21772,N_22232);
or U23082 (N_23082,N_22702,N_22289);
xor U23083 (N_23083,N_22468,N_22657);
or U23084 (N_23084,N_21713,N_22389);
and U23085 (N_23085,N_22346,N_22756);
nand U23086 (N_23086,N_21689,N_21796);
nor U23087 (N_23087,N_21998,N_22054);
or U23088 (N_23088,N_22284,N_22355);
nor U23089 (N_23089,N_21912,N_22451);
or U23090 (N_23090,N_21750,N_21661);
nor U23091 (N_23091,N_22227,N_21624);
nor U23092 (N_23092,N_22371,N_22053);
xor U23093 (N_23093,N_22727,N_21719);
and U23094 (N_23094,N_21809,N_21891);
nand U23095 (N_23095,N_22096,N_21976);
or U23096 (N_23096,N_22250,N_22342);
and U23097 (N_23097,N_22607,N_22582);
nand U23098 (N_23098,N_22472,N_22473);
nor U23099 (N_23099,N_22287,N_21997);
and U23100 (N_23100,N_22092,N_22586);
nand U23101 (N_23101,N_22529,N_22420);
and U23102 (N_23102,N_22066,N_22597);
nand U23103 (N_23103,N_22374,N_21988);
xnor U23104 (N_23104,N_21951,N_22479);
nor U23105 (N_23105,N_22731,N_22748);
and U23106 (N_23106,N_22672,N_22137);
or U23107 (N_23107,N_22370,N_21792);
nand U23108 (N_23108,N_22070,N_21760);
and U23109 (N_23109,N_22563,N_21620);
nor U23110 (N_23110,N_22313,N_22281);
or U23111 (N_23111,N_22218,N_22101);
or U23112 (N_23112,N_21918,N_22436);
and U23113 (N_23113,N_22578,N_22628);
or U23114 (N_23114,N_21701,N_22599);
nand U23115 (N_23115,N_22768,N_21938);
nor U23116 (N_23116,N_22666,N_22392);
nand U23117 (N_23117,N_21898,N_22247);
and U23118 (N_23118,N_22754,N_21670);
xor U23119 (N_23119,N_22644,N_21659);
xor U23120 (N_23120,N_22181,N_22769);
xnor U23121 (N_23121,N_22065,N_21994);
or U23122 (N_23122,N_21756,N_22716);
or U23123 (N_23123,N_22238,N_22314);
xor U23124 (N_23124,N_21803,N_22201);
xnor U23125 (N_23125,N_22751,N_21965);
nor U23126 (N_23126,N_21817,N_21718);
nor U23127 (N_23127,N_22608,N_22383);
nor U23128 (N_23128,N_22554,N_22509);
nor U23129 (N_23129,N_22059,N_22391);
xor U23130 (N_23130,N_21725,N_22733);
xor U23131 (N_23131,N_22180,N_22094);
and U23132 (N_23132,N_22357,N_22645);
xnor U23133 (N_23133,N_22251,N_21798);
xor U23134 (N_23134,N_21700,N_21927);
and U23135 (N_23135,N_22540,N_22248);
xor U23136 (N_23136,N_21778,N_21967);
nand U23137 (N_23137,N_22091,N_21987);
or U23138 (N_23138,N_22150,N_22199);
xor U23139 (N_23139,N_21646,N_22685);
nor U23140 (N_23140,N_21860,N_22767);
xor U23141 (N_23141,N_21880,N_22385);
xnor U23142 (N_23142,N_22210,N_22377);
and U23143 (N_23143,N_22138,N_21691);
nand U23144 (N_23144,N_22494,N_21944);
nor U23145 (N_23145,N_21777,N_22014);
or U23146 (N_23146,N_22037,N_22640);
xor U23147 (N_23147,N_21948,N_22071);
nor U23148 (N_23148,N_22410,N_22200);
and U23149 (N_23149,N_22461,N_22386);
nand U23150 (N_23150,N_21639,N_22002);
nand U23151 (N_23151,N_22627,N_21847);
nor U23152 (N_23152,N_22612,N_21986);
or U23153 (N_23153,N_22629,N_21829);
or U23154 (N_23154,N_22758,N_21815);
nor U23155 (N_23155,N_22081,N_22255);
or U23156 (N_23156,N_22394,N_22434);
nor U23157 (N_23157,N_22300,N_22516);
xor U23158 (N_23158,N_22633,N_21771);
xor U23159 (N_23159,N_22018,N_21905);
nand U23160 (N_23160,N_22382,N_21707);
and U23161 (N_23161,N_21731,N_22185);
xnor U23162 (N_23162,N_21953,N_22441);
or U23163 (N_23163,N_22381,N_21853);
and U23164 (N_23164,N_22463,N_22774);
nor U23165 (N_23165,N_22630,N_22492);
and U23166 (N_23166,N_22799,N_22722);
and U23167 (N_23167,N_22401,N_22448);
or U23168 (N_23168,N_21686,N_21623);
xnor U23169 (N_23169,N_21933,N_22038);
xor U23170 (N_23170,N_22246,N_21839);
and U23171 (N_23171,N_22336,N_22280);
or U23172 (N_23172,N_21606,N_22302);
nor U23173 (N_23173,N_21702,N_22499);
and U23174 (N_23174,N_22462,N_22228);
or U23175 (N_23175,N_22753,N_22631);
xnor U23176 (N_23176,N_22290,N_22159);
or U23177 (N_23177,N_22699,N_22646);
nor U23178 (N_23178,N_22351,N_22665);
xnor U23179 (N_23179,N_21959,N_22166);
and U23180 (N_23180,N_22625,N_21894);
and U23181 (N_23181,N_22234,N_22426);
or U23182 (N_23182,N_22425,N_22734);
or U23183 (N_23183,N_22112,N_21611);
nand U23184 (N_23184,N_22519,N_21757);
and U23185 (N_23185,N_22088,N_21931);
nand U23186 (N_23186,N_21681,N_21871);
and U23187 (N_23187,N_22482,N_22773);
nor U23188 (N_23188,N_22610,N_22695);
nor U23189 (N_23189,N_21692,N_21897);
nand U23190 (N_23190,N_21848,N_22541);
or U23191 (N_23191,N_21973,N_22435);
nand U23192 (N_23192,N_22576,N_22572);
nor U23193 (N_23193,N_22611,N_22518);
nand U23194 (N_23194,N_22241,N_21850);
nor U23195 (N_23195,N_21784,N_22617);
nor U23196 (N_23196,N_21814,N_22278);
nor U23197 (N_23197,N_22752,N_22008);
and U23198 (N_23198,N_22796,N_22705);
or U23199 (N_23199,N_22732,N_22093);
and U23200 (N_23200,N_22653,N_21974);
or U23201 (N_23201,N_22340,N_22209);
and U23202 (N_23202,N_21916,N_21962);
nor U23203 (N_23203,N_21617,N_21711);
or U23204 (N_23204,N_22169,N_21936);
xnor U23205 (N_23205,N_21656,N_22303);
and U23206 (N_23206,N_22786,N_22177);
and U23207 (N_23207,N_22295,N_22023);
nand U23208 (N_23208,N_22654,N_22746);
or U23209 (N_23209,N_21751,N_21955);
nor U23210 (N_23210,N_22319,N_22780);
or U23211 (N_23211,N_21837,N_22348);
or U23212 (N_23212,N_22190,N_22239);
xor U23213 (N_23213,N_22710,N_22636);
xnor U23214 (N_23214,N_22624,N_22021);
or U23215 (N_23215,N_22533,N_21928);
nor U23216 (N_23216,N_21753,N_22632);
or U23217 (N_23217,N_21665,N_22367);
nand U23218 (N_23218,N_22562,N_22173);
xor U23219 (N_23219,N_22557,N_22432);
nor U23220 (N_23220,N_22283,N_22592);
or U23221 (N_23221,N_22517,N_22431);
or U23222 (N_23222,N_21675,N_22776);
or U23223 (N_23223,N_22207,N_22795);
or U23224 (N_23224,N_21601,N_22260);
nor U23225 (N_23225,N_21737,N_21728);
nand U23226 (N_23226,N_21683,N_22045);
nor U23227 (N_23227,N_22360,N_21932);
and U23228 (N_23228,N_21868,N_22328);
and U23229 (N_23229,N_22011,N_22240);
or U23230 (N_23230,N_22327,N_22305);
nand U23231 (N_23231,N_21884,N_22022);
nor U23232 (N_23232,N_22095,N_22460);
or U23233 (N_23233,N_22542,N_22614);
xor U23234 (N_23234,N_21652,N_22117);
or U23235 (N_23235,N_21671,N_22458);
xnor U23236 (N_23236,N_21695,N_22110);
xnor U23237 (N_23237,N_21712,N_21764);
and U23238 (N_23238,N_22766,N_22423);
and U23239 (N_23239,N_21903,N_22249);
nand U23240 (N_23240,N_22072,N_21947);
nand U23241 (N_23241,N_22341,N_21954);
nor U23242 (N_23242,N_22686,N_21744);
and U23243 (N_23243,N_22675,N_22286);
and U23244 (N_23244,N_22498,N_21825);
and U23245 (N_23245,N_22569,N_22704);
xnor U23246 (N_23246,N_22433,N_22589);
nand U23247 (N_23247,N_22293,N_21970);
or U23248 (N_23248,N_22333,N_22764);
nor U23249 (N_23249,N_22737,N_22020);
and U23250 (N_23250,N_22794,N_21774);
or U23251 (N_23251,N_22706,N_22556);
nor U23252 (N_23252,N_22388,N_21694);
nor U23253 (N_23253,N_22502,N_21770);
nand U23254 (N_23254,N_22549,N_22749);
and U23255 (N_23255,N_22171,N_22279);
xor U23256 (N_23256,N_22466,N_22476);
and U23257 (N_23257,N_22558,N_21823);
or U23258 (N_23258,N_21975,N_22545);
nand U23259 (N_23259,N_22421,N_22378);
or U23260 (N_23260,N_22235,N_21710);
xor U23261 (N_23261,N_21921,N_22039);
or U23262 (N_23262,N_21754,N_22604);
nor U23263 (N_23263,N_22147,N_22651);
nand U23264 (N_23264,N_21715,N_22326);
nand U23265 (N_23265,N_22365,N_21723);
xnor U23266 (N_23266,N_21782,N_22712);
nand U23267 (N_23267,N_21602,N_22265);
or U23268 (N_23268,N_22407,N_22028);
xnor U23269 (N_23269,N_21678,N_21621);
or U23270 (N_23270,N_22168,N_21788);
and U23271 (N_23271,N_22598,N_21614);
or U23272 (N_23272,N_22188,N_22551);
nor U23273 (N_23273,N_22221,N_22616);
nor U23274 (N_23274,N_22477,N_22233);
and U23275 (N_23275,N_22213,N_22010);
nand U23276 (N_23276,N_22532,N_21845);
xnor U23277 (N_23277,N_22483,N_22332);
xor U23278 (N_23278,N_22262,N_21907);
or U23279 (N_23279,N_22035,N_22662);
and U23280 (N_23280,N_22126,N_22291);
or U23281 (N_23281,N_22583,N_22339);
or U23282 (N_23282,N_22145,N_21821);
and U23283 (N_23283,N_22142,N_21945);
xor U23284 (N_23284,N_21767,N_21722);
or U23285 (N_23285,N_21762,N_21855);
or U23286 (N_23286,N_21857,N_22390);
and U23287 (N_23287,N_22447,N_21971);
and U23288 (N_23288,N_22656,N_22565);
nand U23289 (N_23289,N_22547,N_22659);
xor U23290 (N_23290,N_21887,N_22484);
xnor U23291 (N_23291,N_22090,N_22515);
xor U23292 (N_23292,N_21890,N_22501);
and U23293 (N_23293,N_22043,N_21785);
and U23294 (N_23294,N_22772,N_21631);
or U23295 (N_23295,N_22226,N_22272);
nor U23296 (N_23296,N_21801,N_22017);
xnor U23297 (N_23297,N_22587,N_22015);
xor U23298 (N_23298,N_21684,N_21908);
or U23299 (N_23299,N_21901,N_22564);
and U23300 (N_23300,N_21786,N_22276);
nand U23301 (N_23301,N_21867,N_22133);
and U23302 (N_23302,N_22687,N_21714);
nor U23303 (N_23303,N_21799,N_21840);
xnor U23304 (N_23304,N_21630,N_21696);
nand U23305 (N_23305,N_21693,N_22056);
or U23306 (N_23306,N_21629,N_22526);
xnor U23307 (N_23307,N_22530,N_22459);
nand U23308 (N_23308,N_21600,N_22078);
and U23309 (N_23309,N_22621,N_22359);
nor U23310 (N_23310,N_21644,N_21846);
nand U23311 (N_23311,N_21673,N_22345);
nor U23312 (N_23312,N_21766,N_22763);
nor U23313 (N_23313,N_22048,N_22641);
xor U23314 (N_23314,N_22414,N_22285);
nor U23315 (N_23315,N_22245,N_22064);
nand U23316 (N_23316,N_22485,N_21742);
and U23317 (N_23317,N_22521,N_21662);
nand U23318 (N_23318,N_22082,N_22016);
nand U23319 (N_23319,N_22132,N_22108);
and U23320 (N_23320,N_22154,N_21795);
nand U23321 (N_23321,N_21913,N_22577);
nand U23322 (N_23322,N_22195,N_21615);
xnor U23323 (N_23323,N_22320,N_22798);
nand U23324 (N_23324,N_22618,N_22033);
and U23325 (N_23325,N_21992,N_22025);
nand U23326 (N_23326,N_21752,N_22437);
xor U23327 (N_23327,N_22595,N_21822);
and U23328 (N_23328,N_21755,N_22491);
nand U23329 (N_23329,N_21669,N_22635);
and U23330 (N_23330,N_22269,N_22135);
nor U23331 (N_23331,N_21619,N_22107);
and U23332 (N_23332,N_22128,N_22789);
nor U23333 (N_23333,N_22449,N_21773);
or U23334 (N_23334,N_22009,N_22182);
nor U23335 (N_23335,N_21981,N_22791);
xor U23336 (N_23336,N_21651,N_22511);
nor U23337 (N_23337,N_21961,N_21666);
or U23338 (N_23338,N_22178,N_21653);
nand U23339 (N_23339,N_21904,N_22506);
nor U23340 (N_23340,N_22471,N_21856);
nand U23341 (N_23341,N_21807,N_21802);
nor U23342 (N_23342,N_22538,N_21605);
and U23343 (N_23343,N_21866,N_21625);
xnor U23344 (N_23344,N_22622,N_22398);
xnor U23345 (N_23345,N_22164,N_22217);
and U23346 (N_23346,N_21603,N_21805);
nand U23347 (N_23347,N_21873,N_22361);
or U23348 (N_23348,N_22413,N_22428);
nand U23349 (N_23349,N_22069,N_22298);
xor U23350 (N_23350,N_22104,N_22368);
or U23351 (N_23351,N_22380,N_22204);
and U23352 (N_23352,N_22321,N_22347);
and U23353 (N_23353,N_21895,N_22444);
nand U23354 (N_23354,N_22552,N_21674);
xnor U23355 (N_23355,N_21816,N_22609);
nand U23356 (N_23356,N_21642,N_22222);
nand U23357 (N_23357,N_22747,N_21843);
nor U23358 (N_23358,N_22264,N_21638);
nor U23359 (N_23359,N_22707,N_22307);
xor U23360 (N_23360,N_21999,N_22224);
nand U23361 (N_23361,N_22061,N_21978);
or U23362 (N_23362,N_22709,N_22602);
nor U23363 (N_23363,N_21806,N_22452);
nand U23364 (N_23364,N_21910,N_22419);
or U23365 (N_23365,N_21919,N_22490);
and U23366 (N_23366,N_21835,N_22412);
and U23367 (N_23367,N_22744,N_22634);
nand U23368 (N_23368,N_21679,N_22170);
or U23369 (N_23369,N_22402,N_21732);
nor U23370 (N_23370,N_22717,N_21925);
nand U23371 (N_23371,N_22197,N_22193);
nor U23372 (N_23372,N_21935,N_21720);
nand U23373 (N_23373,N_21740,N_22256);
and U23374 (N_23374,N_22781,N_22512);
nand U23375 (N_23375,N_22792,N_21926);
nand U23376 (N_23376,N_22575,N_21636);
or U23377 (N_23377,N_22165,N_22012);
or U23378 (N_23378,N_22660,N_22566);
and U23379 (N_23379,N_22676,N_22373);
nand U23380 (N_23380,N_21663,N_22206);
nand U23381 (N_23381,N_22735,N_21872);
and U23382 (N_23382,N_22192,N_22470);
nand U23383 (N_23383,N_22770,N_21854);
nand U23384 (N_23384,N_21793,N_21672);
nor U23385 (N_23385,N_22601,N_22057);
or U23386 (N_23386,N_22266,N_22019);
nor U23387 (N_23387,N_22157,N_21741);
nand U23388 (N_23388,N_22317,N_22013);
nor U23389 (N_23389,N_21761,N_22277);
and U23390 (N_23390,N_22787,N_21703);
or U23391 (N_23391,N_22271,N_22692);
or U23392 (N_23392,N_21993,N_22480);
and U23393 (N_23393,N_22335,N_22352);
nand U23394 (N_23394,N_21613,N_21738);
and U23395 (N_23395,N_22496,N_22639);
or U23396 (N_23396,N_22454,N_21654);
nor U23397 (N_23397,N_21698,N_22049);
nor U23398 (N_23398,N_21985,N_22724);
or U23399 (N_23399,N_21780,N_22301);
nand U23400 (N_23400,N_21647,N_22359);
nand U23401 (N_23401,N_22538,N_21716);
xor U23402 (N_23402,N_22568,N_21937);
xnor U23403 (N_23403,N_22152,N_21810);
xor U23404 (N_23404,N_22356,N_21703);
xnor U23405 (N_23405,N_22132,N_22459);
xor U23406 (N_23406,N_21994,N_21712);
and U23407 (N_23407,N_22334,N_21721);
or U23408 (N_23408,N_22513,N_22069);
xnor U23409 (N_23409,N_21729,N_22290);
xor U23410 (N_23410,N_22039,N_22477);
or U23411 (N_23411,N_22441,N_21772);
nor U23412 (N_23412,N_21789,N_21961);
xor U23413 (N_23413,N_22576,N_22281);
or U23414 (N_23414,N_21913,N_21849);
or U23415 (N_23415,N_22421,N_21821);
xor U23416 (N_23416,N_22227,N_22734);
and U23417 (N_23417,N_22711,N_21877);
nand U23418 (N_23418,N_21648,N_22227);
and U23419 (N_23419,N_21922,N_22737);
nand U23420 (N_23420,N_21977,N_21661);
or U23421 (N_23421,N_21709,N_22327);
nor U23422 (N_23422,N_21711,N_21780);
xor U23423 (N_23423,N_21981,N_22198);
nand U23424 (N_23424,N_22000,N_21730);
nor U23425 (N_23425,N_22006,N_21609);
or U23426 (N_23426,N_22670,N_22031);
xor U23427 (N_23427,N_22415,N_22699);
nand U23428 (N_23428,N_21748,N_22004);
or U23429 (N_23429,N_21858,N_22510);
xnor U23430 (N_23430,N_21823,N_21729);
and U23431 (N_23431,N_22020,N_22313);
xnor U23432 (N_23432,N_21874,N_22528);
or U23433 (N_23433,N_22284,N_21866);
xnor U23434 (N_23434,N_21861,N_22526);
nand U23435 (N_23435,N_22518,N_21845);
xor U23436 (N_23436,N_21715,N_22169);
or U23437 (N_23437,N_22421,N_22225);
nand U23438 (N_23438,N_22568,N_21815);
xnor U23439 (N_23439,N_22081,N_22548);
nand U23440 (N_23440,N_22759,N_21941);
nor U23441 (N_23441,N_22174,N_21686);
xor U23442 (N_23442,N_22438,N_22427);
and U23443 (N_23443,N_22522,N_22709);
xor U23444 (N_23444,N_22419,N_22026);
nor U23445 (N_23445,N_22752,N_21815);
xnor U23446 (N_23446,N_22351,N_22458);
nand U23447 (N_23447,N_22481,N_22703);
nand U23448 (N_23448,N_22759,N_22435);
nand U23449 (N_23449,N_21770,N_22358);
nor U23450 (N_23450,N_22049,N_22285);
xnor U23451 (N_23451,N_21949,N_22203);
or U23452 (N_23452,N_22377,N_22108);
or U23453 (N_23453,N_22423,N_21926);
xor U23454 (N_23454,N_22694,N_22581);
and U23455 (N_23455,N_21630,N_21728);
xnor U23456 (N_23456,N_21764,N_22314);
nand U23457 (N_23457,N_22497,N_21697);
nand U23458 (N_23458,N_21956,N_22634);
nand U23459 (N_23459,N_22336,N_22221);
nor U23460 (N_23460,N_21700,N_22140);
or U23461 (N_23461,N_22769,N_22744);
xnor U23462 (N_23462,N_21974,N_22491);
nor U23463 (N_23463,N_21942,N_22592);
or U23464 (N_23464,N_22721,N_22203);
or U23465 (N_23465,N_21623,N_22588);
or U23466 (N_23466,N_22641,N_22441);
nor U23467 (N_23467,N_22226,N_22778);
or U23468 (N_23468,N_22553,N_22565);
and U23469 (N_23469,N_22294,N_22041);
nand U23470 (N_23470,N_22044,N_22270);
or U23471 (N_23471,N_21697,N_22143);
nor U23472 (N_23472,N_22377,N_21917);
nor U23473 (N_23473,N_22671,N_21843);
nor U23474 (N_23474,N_22314,N_22240);
xnor U23475 (N_23475,N_21918,N_22425);
xnor U23476 (N_23476,N_22369,N_21816);
nand U23477 (N_23477,N_21765,N_22263);
and U23478 (N_23478,N_22327,N_21708);
and U23479 (N_23479,N_22102,N_21890);
nor U23480 (N_23480,N_22440,N_22738);
or U23481 (N_23481,N_22072,N_21620);
and U23482 (N_23482,N_21641,N_22206);
nor U23483 (N_23483,N_21850,N_22477);
nand U23484 (N_23484,N_21982,N_21807);
nand U23485 (N_23485,N_21873,N_21685);
or U23486 (N_23486,N_22632,N_22710);
nor U23487 (N_23487,N_22727,N_22232);
nand U23488 (N_23488,N_22003,N_22577);
or U23489 (N_23489,N_22561,N_22400);
nand U23490 (N_23490,N_22213,N_21949);
nand U23491 (N_23491,N_22616,N_22761);
xnor U23492 (N_23492,N_21741,N_21886);
nand U23493 (N_23493,N_22647,N_22620);
nand U23494 (N_23494,N_22651,N_22011);
or U23495 (N_23495,N_21918,N_21700);
nor U23496 (N_23496,N_21849,N_22573);
and U23497 (N_23497,N_22151,N_21971);
or U23498 (N_23498,N_21956,N_22733);
nand U23499 (N_23499,N_22769,N_22606);
or U23500 (N_23500,N_21819,N_21822);
and U23501 (N_23501,N_22260,N_21656);
xor U23502 (N_23502,N_22618,N_22233);
and U23503 (N_23503,N_21865,N_22298);
and U23504 (N_23504,N_22512,N_22650);
or U23505 (N_23505,N_21818,N_22742);
and U23506 (N_23506,N_21983,N_21743);
or U23507 (N_23507,N_22632,N_22158);
and U23508 (N_23508,N_22635,N_22757);
nor U23509 (N_23509,N_21701,N_22419);
or U23510 (N_23510,N_21648,N_21922);
nand U23511 (N_23511,N_22225,N_22165);
and U23512 (N_23512,N_21802,N_22127);
nor U23513 (N_23513,N_22711,N_21823);
nand U23514 (N_23514,N_22058,N_22722);
or U23515 (N_23515,N_21786,N_22349);
or U23516 (N_23516,N_22323,N_22329);
xor U23517 (N_23517,N_22605,N_21976);
nor U23518 (N_23518,N_22391,N_22660);
nor U23519 (N_23519,N_21954,N_22765);
xnor U23520 (N_23520,N_22773,N_22062);
xnor U23521 (N_23521,N_22429,N_22763);
or U23522 (N_23522,N_22293,N_21831);
nor U23523 (N_23523,N_22626,N_22547);
nand U23524 (N_23524,N_22766,N_22205);
or U23525 (N_23525,N_22639,N_22614);
nand U23526 (N_23526,N_22456,N_22127);
nor U23527 (N_23527,N_21779,N_22068);
or U23528 (N_23528,N_22479,N_21939);
nand U23529 (N_23529,N_22007,N_22713);
xor U23530 (N_23530,N_22541,N_22539);
and U23531 (N_23531,N_21757,N_22701);
or U23532 (N_23532,N_21794,N_21927);
xor U23533 (N_23533,N_21848,N_22459);
and U23534 (N_23534,N_22177,N_22613);
or U23535 (N_23535,N_22699,N_22483);
nand U23536 (N_23536,N_21999,N_22222);
nand U23537 (N_23537,N_22490,N_22569);
xnor U23538 (N_23538,N_22580,N_21850);
xor U23539 (N_23539,N_21907,N_21942);
xnor U23540 (N_23540,N_22337,N_21661);
or U23541 (N_23541,N_22668,N_22266);
xnor U23542 (N_23542,N_22447,N_22307);
nand U23543 (N_23543,N_22285,N_22018);
nor U23544 (N_23544,N_21990,N_22719);
nand U23545 (N_23545,N_22774,N_21820);
xor U23546 (N_23546,N_21618,N_21714);
nor U23547 (N_23547,N_22227,N_22010);
or U23548 (N_23548,N_21781,N_22540);
xor U23549 (N_23549,N_21984,N_22248);
and U23550 (N_23550,N_21913,N_22359);
xor U23551 (N_23551,N_21653,N_21978);
and U23552 (N_23552,N_22026,N_21922);
nor U23553 (N_23553,N_22389,N_21994);
xor U23554 (N_23554,N_21691,N_22070);
and U23555 (N_23555,N_22571,N_21750);
and U23556 (N_23556,N_21812,N_22519);
xnor U23557 (N_23557,N_22118,N_22580);
nor U23558 (N_23558,N_22265,N_21679);
xnor U23559 (N_23559,N_21936,N_22478);
nand U23560 (N_23560,N_22015,N_22435);
xnor U23561 (N_23561,N_22037,N_22548);
and U23562 (N_23562,N_21813,N_22614);
or U23563 (N_23563,N_21787,N_21720);
and U23564 (N_23564,N_22080,N_21629);
and U23565 (N_23565,N_22159,N_22105);
nor U23566 (N_23566,N_21983,N_22119);
and U23567 (N_23567,N_21716,N_22225);
and U23568 (N_23568,N_22274,N_22144);
xnor U23569 (N_23569,N_21999,N_21842);
or U23570 (N_23570,N_22220,N_21710);
xor U23571 (N_23571,N_21664,N_22532);
or U23572 (N_23572,N_22165,N_22385);
or U23573 (N_23573,N_21760,N_22497);
nand U23574 (N_23574,N_22583,N_22334);
nor U23575 (N_23575,N_22006,N_21959);
or U23576 (N_23576,N_22388,N_21926);
nor U23577 (N_23577,N_22164,N_22137);
and U23578 (N_23578,N_22060,N_22381);
and U23579 (N_23579,N_22408,N_21928);
and U23580 (N_23580,N_22239,N_21904);
nor U23581 (N_23581,N_21617,N_22460);
nor U23582 (N_23582,N_21607,N_22073);
nor U23583 (N_23583,N_21928,N_22235);
or U23584 (N_23584,N_22349,N_21913);
nor U23585 (N_23585,N_21821,N_21863);
xnor U23586 (N_23586,N_22407,N_21904);
nor U23587 (N_23587,N_21610,N_21654);
nand U23588 (N_23588,N_21740,N_22502);
and U23589 (N_23589,N_21889,N_22768);
xnor U23590 (N_23590,N_22794,N_22228);
and U23591 (N_23591,N_22125,N_21676);
nand U23592 (N_23592,N_21733,N_22450);
and U23593 (N_23593,N_22733,N_22690);
and U23594 (N_23594,N_21667,N_22490);
nand U23595 (N_23595,N_21759,N_21873);
and U23596 (N_23596,N_22480,N_22412);
nor U23597 (N_23597,N_21782,N_22231);
xnor U23598 (N_23598,N_22641,N_22350);
nand U23599 (N_23599,N_21843,N_22528);
nand U23600 (N_23600,N_22757,N_22102);
nand U23601 (N_23601,N_22237,N_21632);
nand U23602 (N_23602,N_22077,N_22209);
nand U23603 (N_23603,N_22415,N_22595);
xor U23604 (N_23604,N_22309,N_21649);
or U23605 (N_23605,N_22136,N_22228);
and U23606 (N_23606,N_22450,N_22636);
or U23607 (N_23607,N_22716,N_22689);
or U23608 (N_23608,N_21972,N_22781);
and U23609 (N_23609,N_22424,N_22198);
or U23610 (N_23610,N_21976,N_22504);
and U23611 (N_23611,N_22746,N_22194);
nand U23612 (N_23612,N_22311,N_22420);
xnor U23613 (N_23613,N_22216,N_22224);
xor U23614 (N_23614,N_22488,N_22309);
nor U23615 (N_23615,N_22719,N_21704);
xnor U23616 (N_23616,N_22048,N_21779);
or U23617 (N_23617,N_22711,N_21927);
and U23618 (N_23618,N_22196,N_21865);
or U23619 (N_23619,N_21906,N_22429);
nand U23620 (N_23620,N_22408,N_22230);
and U23621 (N_23621,N_21892,N_21965);
nor U23622 (N_23622,N_21879,N_22708);
and U23623 (N_23623,N_22021,N_22731);
nand U23624 (N_23624,N_22372,N_22153);
and U23625 (N_23625,N_21860,N_22168);
nor U23626 (N_23626,N_22539,N_21907);
nor U23627 (N_23627,N_22554,N_22744);
nand U23628 (N_23628,N_22327,N_22197);
or U23629 (N_23629,N_21986,N_21753);
nor U23630 (N_23630,N_22636,N_21889);
and U23631 (N_23631,N_22687,N_21877);
nand U23632 (N_23632,N_22735,N_22286);
nand U23633 (N_23633,N_22025,N_22147);
nand U23634 (N_23634,N_22536,N_22057);
xor U23635 (N_23635,N_21939,N_22210);
nor U23636 (N_23636,N_21705,N_22409);
and U23637 (N_23637,N_22450,N_21626);
and U23638 (N_23638,N_22213,N_22173);
nor U23639 (N_23639,N_21620,N_22780);
nor U23640 (N_23640,N_22698,N_22702);
nand U23641 (N_23641,N_21765,N_22506);
xnor U23642 (N_23642,N_22640,N_21876);
or U23643 (N_23643,N_22262,N_21779);
nand U23644 (N_23644,N_21699,N_21934);
or U23645 (N_23645,N_22768,N_21951);
xnor U23646 (N_23646,N_22531,N_22384);
nor U23647 (N_23647,N_22216,N_21740);
and U23648 (N_23648,N_22454,N_22227);
xor U23649 (N_23649,N_21987,N_22270);
and U23650 (N_23650,N_21851,N_21814);
or U23651 (N_23651,N_22569,N_22542);
nor U23652 (N_23652,N_21828,N_21993);
and U23653 (N_23653,N_22113,N_22528);
or U23654 (N_23654,N_21795,N_21631);
and U23655 (N_23655,N_22276,N_22471);
nand U23656 (N_23656,N_22575,N_22211);
and U23657 (N_23657,N_21742,N_21785);
and U23658 (N_23658,N_22181,N_21946);
and U23659 (N_23659,N_22070,N_22531);
or U23660 (N_23660,N_22692,N_22618);
nand U23661 (N_23661,N_22453,N_21773);
nor U23662 (N_23662,N_22767,N_22624);
xnor U23663 (N_23663,N_22513,N_22417);
and U23664 (N_23664,N_22746,N_22795);
xor U23665 (N_23665,N_22352,N_22254);
nand U23666 (N_23666,N_22139,N_22019);
or U23667 (N_23667,N_21946,N_22278);
or U23668 (N_23668,N_22765,N_22347);
nand U23669 (N_23669,N_21773,N_22310);
or U23670 (N_23670,N_22443,N_22532);
or U23671 (N_23671,N_22327,N_21854);
nor U23672 (N_23672,N_22760,N_22269);
and U23673 (N_23673,N_21765,N_22670);
nand U23674 (N_23674,N_22195,N_22656);
nand U23675 (N_23675,N_22325,N_22237);
nand U23676 (N_23676,N_22237,N_22122);
nor U23677 (N_23677,N_21823,N_22134);
nand U23678 (N_23678,N_22288,N_21965);
and U23679 (N_23679,N_21755,N_22629);
xor U23680 (N_23680,N_22656,N_22563);
xor U23681 (N_23681,N_21749,N_22350);
xnor U23682 (N_23682,N_22653,N_22458);
xnor U23683 (N_23683,N_22355,N_21730);
and U23684 (N_23684,N_22749,N_22566);
and U23685 (N_23685,N_22548,N_21882);
and U23686 (N_23686,N_22194,N_21682);
xor U23687 (N_23687,N_21696,N_22247);
nand U23688 (N_23688,N_22194,N_22627);
or U23689 (N_23689,N_22399,N_22247);
xnor U23690 (N_23690,N_21756,N_21932);
nand U23691 (N_23691,N_22127,N_22730);
or U23692 (N_23692,N_22335,N_22653);
nand U23693 (N_23693,N_21994,N_22547);
nand U23694 (N_23694,N_22755,N_22027);
nand U23695 (N_23695,N_22291,N_22254);
or U23696 (N_23696,N_22410,N_22261);
xor U23697 (N_23697,N_21823,N_21878);
and U23698 (N_23698,N_21998,N_22234);
xnor U23699 (N_23699,N_22700,N_21651);
nor U23700 (N_23700,N_22645,N_22323);
nor U23701 (N_23701,N_22262,N_22243);
or U23702 (N_23702,N_22615,N_22406);
xor U23703 (N_23703,N_21801,N_21773);
or U23704 (N_23704,N_21607,N_22093);
nor U23705 (N_23705,N_22658,N_21955);
and U23706 (N_23706,N_22114,N_22372);
nand U23707 (N_23707,N_22412,N_22129);
nor U23708 (N_23708,N_22037,N_21752);
xnor U23709 (N_23709,N_22000,N_22734);
nand U23710 (N_23710,N_21903,N_22555);
and U23711 (N_23711,N_22553,N_21759);
nor U23712 (N_23712,N_22326,N_22063);
nand U23713 (N_23713,N_22286,N_22041);
and U23714 (N_23714,N_21617,N_22281);
or U23715 (N_23715,N_21709,N_22648);
and U23716 (N_23716,N_22363,N_22434);
nor U23717 (N_23717,N_21847,N_21761);
or U23718 (N_23718,N_22235,N_22595);
and U23719 (N_23719,N_21658,N_22679);
and U23720 (N_23720,N_22355,N_22038);
nand U23721 (N_23721,N_22597,N_21758);
and U23722 (N_23722,N_21910,N_22596);
and U23723 (N_23723,N_22418,N_22210);
nand U23724 (N_23724,N_22431,N_22531);
xnor U23725 (N_23725,N_21943,N_22152);
or U23726 (N_23726,N_21884,N_22512);
and U23727 (N_23727,N_22519,N_22036);
or U23728 (N_23728,N_22231,N_22790);
xor U23729 (N_23729,N_21690,N_22486);
and U23730 (N_23730,N_22363,N_21896);
nand U23731 (N_23731,N_22505,N_22330);
or U23732 (N_23732,N_22482,N_22790);
and U23733 (N_23733,N_22675,N_22366);
nand U23734 (N_23734,N_22310,N_21651);
nor U23735 (N_23735,N_22180,N_22671);
nand U23736 (N_23736,N_22304,N_22361);
xnor U23737 (N_23737,N_21993,N_22173);
nand U23738 (N_23738,N_21959,N_22059);
and U23739 (N_23739,N_22152,N_22650);
nand U23740 (N_23740,N_21960,N_22165);
or U23741 (N_23741,N_21645,N_22506);
and U23742 (N_23742,N_22627,N_22130);
and U23743 (N_23743,N_21707,N_22360);
and U23744 (N_23744,N_21996,N_22542);
and U23745 (N_23745,N_22304,N_22593);
or U23746 (N_23746,N_22062,N_22358);
or U23747 (N_23747,N_21858,N_22710);
nor U23748 (N_23748,N_22530,N_22376);
and U23749 (N_23749,N_21831,N_22121);
xnor U23750 (N_23750,N_22790,N_22531);
nor U23751 (N_23751,N_22726,N_22182);
nand U23752 (N_23752,N_21842,N_22598);
nor U23753 (N_23753,N_22172,N_22641);
nand U23754 (N_23754,N_21844,N_22060);
nand U23755 (N_23755,N_21671,N_22073);
nor U23756 (N_23756,N_22292,N_21603);
or U23757 (N_23757,N_21764,N_22229);
xor U23758 (N_23758,N_21607,N_22065);
nor U23759 (N_23759,N_21841,N_22607);
and U23760 (N_23760,N_22535,N_22046);
xor U23761 (N_23761,N_22735,N_22232);
or U23762 (N_23762,N_22420,N_22440);
nand U23763 (N_23763,N_22605,N_21870);
or U23764 (N_23764,N_21777,N_22138);
and U23765 (N_23765,N_22009,N_22371);
xor U23766 (N_23766,N_22784,N_21898);
and U23767 (N_23767,N_22778,N_22589);
nor U23768 (N_23768,N_22037,N_21688);
nand U23769 (N_23769,N_21612,N_22155);
nand U23770 (N_23770,N_22362,N_22475);
and U23771 (N_23771,N_21941,N_21615);
and U23772 (N_23772,N_22208,N_21838);
nor U23773 (N_23773,N_22350,N_21623);
nand U23774 (N_23774,N_21787,N_22792);
xor U23775 (N_23775,N_22407,N_22676);
xor U23776 (N_23776,N_22513,N_22205);
xnor U23777 (N_23777,N_21891,N_22761);
nand U23778 (N_23778,N_22053,N_21735);
nand U23779 (N_23779,N_22444,N_21934);
or U23780 (N_23780,N_22146,N_21642);
nor U23781 (N_23781,N_21922,N_21702);
or U23782 (N_23782,N_21743,N_21646);
nor U23783 (N_23783,N_22221,N_22608);
and U23784 (N_23784,N_21770,N_21624);
xor U23785 (N_23785,N_22788,N_22075);
nor U23786 (N_23786,N_22716,N_22555);
nand U23787 (N_23787,N_21904,N_22008);
nand U23788 (N_23788,N_22607,N_22301);
nor U23789 (N_23789,N_21864,N_22233);
and U23790 (N_23790,N_22744,N_21728);
nor U23791 (N_23791,N_22148,N_22262);
nand U23792 (N_23792,N_22397,N_21796);
xor U23793 (N_23793,N_21834,N_21603);
nor U23794 (N_23794,N_22083,N_21915);
nor U23795 (N_23795,N_21920,N_22294);
nor U23796 (N_23796,N_22087,N_22305);
or U23797 (N_23797,N_22681,N_22733);
or U23798 (N_23798,N_21638,N_22721);
xor U23799 (N_23799,N_22097,N_22587);
or U23800 (N_23800,N_22624,N_22425);
xor U23801 (N_23801,N_22547,N_22789);
and U23802 (N_23802,N_22060,N_22671);
nand U23803 (N_23803,N_21701,N_22570);
nand U23804 (N_23804,N_22640,N_21915);
or U23805 (N_23805,N_22071,N_21766);
xor U23806 (N_23806,N_22064,N_22128);
and U23807 (N_23807,N_22561,N_22654);
or U23808 (N_23808,N_22580,N_22043);
xnor U23809 (N_23809,N_22165,N_22518);
nor U23810 (N_23810,N_22579,N_21724);
xor U23811 (N_23811,N_22337,N_21992);
or U23812 (N_23812,N_22428,N_22617);
or U23813 (N_23813,N_22155,N_22499);
and U23814 (N_23814,N_22010,N_21745);
nand U23815 (N_23815,N_21617,N_21956);
nand U23816 (N_23816,N_22421,N_22791);
and U23817 (N_23817,N_22066,N_21684);
xor U23818 (N_23818,N_22410,N_22767);
nand U23819 (N_23819,N_22518,N_21646);
nor U23820 (N_23820,N_22490,N_22145);
or U23821 (N_23821,N_22138,N_21932);
nand U23822 (N_23822,N_22165,N_21974);
or U23823 (N_23823,N_22468,N_22739);
and U23824 (N_23824,N_22113,N_22765);
or U23825 (N_23825,N_22754,N_22060);
nor U23826 (N_23826,N_22224,N_21972);
xnor U23827 (N_23827,N_22397,N_21736);
nand U23828 (N_23828,N_22021,N_22201);
or U23829 (N_23829,N_22559,N_21602);
nand U23830 (N_23830,N_22664,N_22409);
and U23831 (N_23831,N_22536,N_22784);
nand U23832 (N_23832,N_22558,N_22366);
nand U23833 (N_23833,N_22331,N_22396);
or U23834 (N_23834,N_22485,N_22447);
nor U23835 (N_23835,N_21840,N_22569);
xnor U23836 (N_23836,N_21777,N_22041);
nor U23837 (N_23837,N_22407,N_21918);
xor U23838 (N_23838,N_22684,N_22764);
xor U23839 (N_23839,N_21639,N_22227);
xor U23840 (N_23840,N_22416,N_22662);
xor U23841 (N_23841,N_22730,N_21888);
and U23842 (N_23842,N_22204,N_22756);
or U23843 (N_23843,N_22341,N_21863);
and U23844 (N_23844,N_22623,N_22446);
nor U23845 (N_23845,N_21671,N_22241);
nand U23846 (N_23846,N_21902,N_22452);
or U23847 (N_23847,N_22179,N_21627);
xnor U23848 (N_23848,N_22269,N_21890);
and U23849 (N_23849,N_22210,N_21866);
nor U23850 (N_23850,N_21627,N_22273);
and U23851 (N_23851,N_22653,N_22229);
nand U23852 (N_23852,N_22526,N_21842);
and U23853 (N_23853,N_21932,N_21780);
or U23854 (N_23854,N_21750,N_22340);
xnor U23855 (N_23855,N_22542,N_21939);
or U23856 (N_23856,N_22748,N_22096);
nand U23857 (N_23857,N_22526,N_22431);
and U23858 (N_23858,N_21802,N_21753);
xnor U23859 (N_23859,N_22214,N_21909);
nand U23860 (N_23860,N_22738,N_21614);
nand U23861 (N_23861,N_21929,N_21733);
nand U23862 (N_23862,N_22598,N_21929);
and U23863 (N_23863,N_22189,N_22122);
nand U23864 (N_23864,N_22722,N_22667);
or U23865 (N_23865,N_22602,N_21684);
or U23866 (N_23866,N_21920,N_22442);
and U23867 (N_23867,N_21834,N_21864);
or U23868 (N_23868,N_22256,N_22293);
and U23869 (N_23869,N_22473,N_21975);
nor U23870 (N_23870,N_22030,N_22389);
nor U23871 (N_23871,N_22113,N_22290);
and U23872 (N_23872,N_21601,N_21860);
and U23873 (N_23873,N_21829,N_22305);
nand U23874 (N_23874,N_21876,N_22521);
and U23875 (N_23875,N_21720,N_21893);
xnor U23876 (N_23876,N_21908,N_22023);
or U23877 (N_23877,N_22405,N_22444);
nor U23878 (N_23878,N_21947,N_21603);
and U23879 (N_23879,N_22427,N_22326);
and U23880 (N_23880,N_22510,N_21616);
or U23881 (N_23881,N_22080,N_22102);
or U23882 (N_23882,N_22027,N_21778);
nand U23883 (N_23883,N_21852,N_22484);
and U23884 (N_23884,N_22617,N_22563);
nor U23885 (N_23885,N_21858,N_21811);
nor U23886 (N_23886,N_22600,N_22132);
and U23887 (N_23887,N_22334,N_21707);
xor U23888 (N_23888,N_21893,N_22522);
or U23889 (N_23889,N_21618,N_21846);
nor U23890 (N_23890,N_21786,N_22266);
nand U23891 (N_23891,N_22579,N_21605);
or U23892 (N_23892,N_22661,N_22167);
or U23893 (N_23893,N_22018,N_22533);
xor U23894 (N_23894,N_22166,N_22687);
or U23895 (N_23895,N_22759,N_22488);
xor U23896 (N_23896,N_22399,N_22107);
nor U23897 (N_23897,N_22260,N_21728);
nor U23898 (N_23898,N_22468,N_21620);
and U23899 (N_23899,N_22148,N_22736);
nand U23900 (N_23900,N_21799,N_22471);
nand U23901 (N_23901,N_21800,N_21645);
xor U23902 (N_23902,N_21939,N_22077);
or U23903 (N_23903,N_22017,N_22449);
nor U23904 (N_23904,N_22183,N_21709);
xnor U23905 (N_23905,N_21730,N_22194);
xor U23906 (N_23906,N_22400,N_21736);
xnor U23907 (N_23907,N_22164,N_21838);
nand U23908 (N_23908,N_22765,N_22702);
xnor U23909 (N_23909,N_22368,N_21982);
xnor U23910 (N_23910,N_22117,N_22461);
nor U23911 (N_23911,N_22207,N_21655);
nand U23912 (N_23912,N_22394,N_21877);
and U23913 (N_23913,N_22380,N_22403);
nand U23914 (N_23914,N_22351,N_22640);
nor U23915 (N_23915,N_22062,N_22350);
and U23916 (N_23916,N_21865,N_21658);
or U23917 (N_23917,N_21678,N_22738);
or U23918 (N_23918,N_21942,N_22459);
and U23919 (N_23919,N_22483,N_22614);
nand U23920 (N_23920,N_22603,N_21856);
nor U23921 (N_23921,N_21936,N_21968);
nand U23922 (N_23922,N_22399,N_21815);
and U23923 (N_23923,N_22012,N_21815);
nor U23924 (N_23924,N_21952,N_22792);
and U23925 (N_23925,N_21888,N_21805);
and U23926 (N_23926,N_21829,N_22246);
nor U23927 (N_23927,N_22529,N_22533);
nand U23928 (N_23928,N_21923,N_21945);
nor U23929 (N_23929,N_22440,N_22647);
or U23930 (N_23930,N_22158,N_21976);
and U23931 (N_23931,N_22115,N_21739);
or U23932 (N_23932,N_22472,N_22302);
and U23933 (N_23933,N_22200,N_22651);
nand U23934 (N_23934,N_21942,N_22699);
nand U23935 (N_23935,N_21975,N_22521);
nand U23936 (N_23936,N_22449,N_22508);
xor U23937 (N_23937,N_22541,N_21791);
and U23938 (N_23938,N_22272,N_22140);
or U23939 (N_23939,N_21680,N_22418);
nor U23940 (N_23940,N_22631,N_21854);
nand U23941 (N_23941,N_22233,N_21632);
nor U23942 (N_23942,N_22351,N_22035);
nand U23943 (N_23943,N_21608,N_22281);
and U23944 (N_23944,N_22561,N_22777);
xnor U23945 (N_23945,N_22087,N_22656);
nor U23946 (N_23946,N_22261,N_22786);
xor U23947 (N_23947,N_22413,N_22174);
nand U23948 (N_23948,N_21789,N_22484);
and U23949 (N_23949,N_22373,N_21603);
and U23950 (N_23950,N_22652,N_21932);
nor U23951 (N_23951,N_21919,N_22729);
xnor U23952 (N_23952,N_22370,N_22443);
nand U23953 (N_23953,N_22588,N_22696);
and U23954 (N_23954,N_21636,N_22075);
or U23955 (N_23955,N_21897,N_22268);
or U23956 (N_23956,N_21624,N_21682);
nor U23957 (N_23957,N_22125,N_22689);
nand U23958 (N_23958,N_22411,N_22127);
or U23959 (N_23959,N_21987,N_22532);
or U23960 (N_23960,N_22404,N_22656);
xnor U23961 (N_23961,N_22064,N_22597);
or U23962 (N_23962,N_22050,N_22095);
and U23963 (N_23963,N_21810,N_22026);
nor U23964 (N_23964,N_22387,N_22290);
xor U23965 (N_23965,N_22172,N_22592);
and U23966 (N_23966,N_22372,N_22532);
xor U23967 (N_23967,N_22466,N_22147);
nor U23968 (N_23968,N_22604,N_21988);
and U23969 (N_23969,N_22115,N_22559);
nand U23970 (N_23970,N_21628,N_21884);
nand U23971 (N_23971,N_21986,N_21678);
or U23972 (N_23972,N_21855,N_22230);
xnor U23973 (N_23973,N_22499,N_22208);
xnor U23974 (N_23974,N_21654,N_21721);
xor U23975 (N_23975,N_22386,N_22027);
nor U23976 (N_23976,N_22707,N_22505);
and U23977 (N_23977,N_21615,N_22153);
and U23978 (N_23978,N_21706,N_22408);
xnor U23979 (N_23979,N_21659,N_21651);
xor U23980 (N_23980,N_22001,N_21621);
nand U23981 (N_23981,N_21614,N_22749);
nand U23982 (N_23982,N_22433,N_22714);
and U23983 (N_23983,N_22334,N_21706);
or U23984 (N_23984,N_22168,N_21967);
nor U23985 (N_23985,N_21662,N_22174);
and U23986 (N_23986,N_21634,N_22438);
and U23987 (N_23987,N_22463,N_22712);
xnor U23988 (N_23988,N_22115,N_22106);
nand U23989 (N_23989,N_22115,N_22345);
nand U23990 (N_23990,N_21746,N_21828);
nand U23991 (N_23991,N_22702,N_22071);
xor U23992 (N_23992,N_22331,N_22769);
xor U23993 (N_23993,N_21871,N_22161);
xor U23994 (N_23994,N_22443,N_22005);
nor U23995 (N_23995,N_22761,N_22248);
xnor U23996 (N_23996,N_22489,N_22186);
nand U23997 (N_23997,N_21836,N_21853);
nand U23998 (N_23998,N_22729,N_21655);
and U23999 (N_23999,N_22367,N_22090);
xor U24000 (N_24000,N_22938,N_23377);
and U24001 (N_24001,N_23399,N_23323);
and U24002 (N_24002,N_23950,N_23178);
nor U24003 (N_24003,N_23917,N_23855);
or U24004 (N_24004,N_23970,N_22835);
or U24005 (N_24005,N_23436,N_23426);
nor U24006 (N_24006,N_23143,N_23908);
nand U24007 (N_24007,N_23918,N_23265);
and U24008 (N_24008,N_23315,N_23607);
and U24009 (N_24009,N_23296,N_23494);
nor U24010 (N_24010,N_23881,N_23184);
and U24011 (N_24011,N_23883,N_23878);
or U24012 (N_24012,N_23848,N_23980);
xor U24013 (N_24013,N_23927,N_23899);
or U24014 (N_24014,N_23404,N_22883);
nor U24015 (N_24015,N_23892,N_23843);
nor U24016 (N_24016,N_23553,N_23111);
xnor U24017 (N_24017,N_23104,N_22884);
and U24018 (N_24018,N_23421,N_23171);
and U24019 (N_24019,N_23569,N_23545);
and U24020 (N_24020,N_23055,N_23630);
and U24021 (N_24021,N_23175,N_23849);
nor U24022 (N_24022,N_23515,N_23413);
nor U24023 (N_24023,N_23228,N_22875);
nor U24024 (N_24024,N_23901,N_22828);
nor U24025 (N_24025,N_23435,N_23162);
and U24026 (N_24026,N_22879,N_23960);
nand U24027 (N_24027,N_23453,N_23028);
and U24028 (N_24028,N_22955,N_23967);
and U24029 (N_24029,N_23324,N_23745);
or U24030 (N_24030,N_23281,N_23423);
xnor U24031 (N_24031,N_23441,N_23839);
nor U24032 (N_24032,N_22885,N_22963);
xor U24033 (N_24033,N_23815,N_23699);
and U24034 (N_24034,N_23022,N_23663);
or U24035 (N_24035,N_23664,N_23505);
nor U24036 (N_24036,N_23149,N_22886);
nor U24037 (N_24037,N_22889,N_22950);
nor U24038 (N_24038,N_23065,N_22932);
nor U24039 (N_24039,N_23557,N_23806);
and U24040 (N_24040,N_23714,N_23734);
and U24041 (N_24041,N_23250,N_23944);
and U24042 (N_24042,N_23754,N_23290);
nor U24043 (N_24043,N_23235,N_23256);
nor U24044 (N_24044,N_23566,N_23858);
xor U24045 (N_24045,N_23314,N_23108);
nand U24046 (N_24046,N_23114,N_23694);
nor U24047 (N_24047,N_23197,N_23631);
nor U24048 (N_24048,N_23711,N_23373);
and U24049 (N_24049,N_23447,N_23466);
xnor U24050 (N_24050,N_23568,N_22990);
nand U24051 (N_24051,N_23186,N_22942);
nor U24052 (N_24052,N_23365,N_23695);
xnor U24053 (N_24053,N_23551,N_23069);
xnor U24054 (N_24054,N_23039,N_23808);
xnor U24055 (N_24055,N_23946,N_22925);
and U24056 (N_24056,N_22867,N_23122);
xor U24057 (N_24057,N_23168,N_22901);
xor U24058 (N_24058,N_23230,N_23217);
xnor U24059 (N_24059,N_22813,N_23123);
nor U24060 (N_24060,N_23564,N_23238);
nor U24061 (N_24061,N_23592,N_23925);
and U24062 (N_24062,N_23137,N_23752);
xnor U24063 (N_24063,N_23876,N_23759);
or U24064 (N_24064,N_23716,N_23442);
nand U24065 (N_24065,N_23945,N_22803);
nor U24066 (N_24066,N_23212,N_22912);
nor U24067 (N_24067,N_23612,N_23457);
and U24068 (N_24068,N_23510,N_23937);
and U24069 (N_24069,N_22838,N_23240);
nand U24070 (N_24070,N_23078,N_22849);
and U24071 (N_24071,N_23718,N_23509);
and U24072 (N_24072,N_23613,N_22975);
xor U24073 (N_24073,N_23420,N_22829);
nand U24074 (N_24074,N_23401,N_23142);
xnor U24075 (N_24075,N_23206,N_23748);
and U24076 (N_24076,N_22928,N_23850);
nand U24077 (N_24077,N_23629,N_23052);
or U24078 (N_24078,N_23319,N_23776);
nor U24079 (N_24079,N_23710,N_23374);
or U24080 (N_24080,N_23583,N_23357);
xor U24081 (N_24081,N_23253,N_22823);
nand U24082 (N_24082,N_23463,N_22863);
nor U24083 (N_24083,N_23412,N_23982);
nand U24084 (N_24084,N_23194,N_23913);
nand U24085 (N_24085,N_23784,N_23382);
nor U24086 (N_24086,N_22979,N_22880);
nand U24087 (N_24087,N_23458,N_23347);
or U24088 (N_24088,N_23796,N_22972);
xnor U24089 (N_24089,N_22987,N_23264);
and U24090 (N_24090,N_23474,N_22916);
or U24091 (N_24091,N_23339,N_23395);
and U24092 (N_24092,N_22831,N_23020);
nor U24093 (N_24093,N_23047,N_23657);
or U24094 (N_24094,N_23160,N_22826);
nor U24095 (N_24095,N_23174,N_23450);
or U24096 (N_24096,N_23169,N_23621);
nand U24097 (N_24097,N_23258,N_23965);
or U24098 (N_24098,N_23904,N_23666);
xor U24099 (N_24099,N_23827,N_23999);
xnor U24100 (N_24100,N_23011,N_23738);
nor U24101 (N_24101,N_23172,N_23124);
or U24102 (N_24102,N_22906,N_23573);
nand U24103 (N_24103,N_23118,N_23682);
and U24104 (N_24104,N_22900,N_22935);
nand U24105 (N_24105,N_23215,N_23529);
xor U24106 (N_24106,N_23139,N_23717);
nor U24107 (N_24107,N_23819,N_23179);
nand U24108 (N_24108,N_23517,N_23167);
and U24109 (N_24109,N_23688,N_22919);
nor U24110 (N_24110,N_23581,N_22986);
or U24111 (N_24111,N_23976,N_22802);
and U24112 (N_24112,N_23035,N_23594);
and U24113 (N_24113,N_22993,N_23454);
nor U24114 (N_24114,N_23222,N_23807);
nand U24115 (N_24115,N_23888,N_23452);
nand U24116 (N_24116,N_23226,N_23084);
xnor U24117 (N_24117,N_23622,N_23891);
or U24118 (N_24118,N_23645,N_23797);
nor U24119 (N_24119,N_23031,N_23107);
nand U24120 (N_24120,N_23391,N_23193);
xor U24121 (N_24121,N_23831,N_23476);
nand U24122 (N_24122,N_23351,N_22852);
and U24123 (N_24123,N_23853,N_23823);
and U24124 (N_24124,N_22821,N_23934);
or U24125 (N_24125,N_22944,N_23667);
nand U24126 (N_24126,N_23309,N_22968);
nor U24127 (N_24127,N_23531,N_23964);
nand U24128 (N_24128,N_22920,N_23761);
nor U24129 (N_24129,N_22865,N_23246);
and U24130 (N_24130,N_23541,N_23998);
or U24131 (N_24131,N_23959,N_23155);
nand U24132 (N_24132,N_22898,N_22805);
and U24133 (N_24133,N_23742,N_23251);
nand U24134 (N_24134,N_23081,N_23275);
nor U24135 (N_24135,N_23987,N_23894);
and U24136 (N_24136,N_23070,N_23241);
or U24137 (N_24137,N_22911,N_23292);
nor U24138 (N_24138,N_23709,N_22891);
nand U24139 (N_24139,N_23864,N_23129);
nor U24140 (N_24140,N_23414,N_23799);
and U24141 (N_24141,N_22801,N_23203);
nand U24142 (N_24142,N_23034,N_23417);
and U24143 (N_24143,N_23283,N_23130);
and U24144 (N_24144,N_23394,N_23978);
or U24145 (N_24145,N_22927,N_23003);
nor U24146 (N_24146,N_23680,N_23266);
xor U24147 (N_24147,N_23276,N_23201);
or U24148 (N_24148,N_23095,N_23434);
and U24149 (N_24149,N_23696,N_23521);
nor U24150 (N_24150,N_23947,N_23019);
nand U24151 (N_24151,N_23390,N_23771);
or U24152 (N_24152,N_23572,N_23958);
nand U24153 (N_24153,N_22832,N_23082);
and U24154 (N_24154,N_23774,N_23582);
and U24155 (N_24155,N_23735,N_23627);
nor U24156 (N_24156,N_23677,N_23671);
xor U24157 (N_24157,N_23781,N_23061);
nor U24158 (N_24158,N_23080,N_23712);
xnor U24159 (N_24159,N_23768,N_23791);
xor U24160 (N_24160,N_23669,N_23514);
or U24161 (N_24161,N_23715,N_23772);
nor U24162 (N_24162,N_23364,N_23218);
nand U24163 (N_24163,N_22862,N_23010);
and U24164 (N_24164,N_22854,N_23792);
nand U24165 (N_24165,N_22913,N_23961);
nand U24166 (N_24166,N_23642,N_23425);
xnor U24167 (N_24167,N_23816,N_23490);
or U24168 (N_24168,N_23623,N_23340);
nand U24169 (N_24169,N_23932,N_22868);
nor U24170 (N_24170,N_23409,N_23345);
nor U24171 (N_24171,N_23144,N_23731);
and U24172 (N_24172,N_22969,N_22872);
or U24173 (N_24173,N_23181,N_23448);
xor U24174 (N_24174,N_23896,N_22910);
xnor U24175 (N_24175,N_23350,N_22941);
xor U24176 (N_24176,N_23727,N_23170);
and U24177 (N_24177,N_22903,N_23620);
xor U24178 (N_24178,N_23334,N_23646);
and U24179 (N_24179,N_23587,N_23886);
and U24180 (N_24180,N_23018,N_23979);
or U24181 (N_24181,N_22847,N_23141);
nand U24182 (N_24182,N_23578,N_23654);
nand U24183 (N_24183,N_23879,N_23535);
and U24184 (N_24184,N_23159,N_23308);
nand U24185 (N_24185,N_23626,N_23873);
nand U24186 (N_24186,N_22807,N_23307);
and U24187 (N_24187,N_22976,N_23562);
nand U24188 (N_24188,N_23190,N_23121);
or U24189 (N_24189,N_23755,N_23237);
nor U24190 (N_24190,N_23056,N_23493);
and U24191 (N_24191,N_23239,N_23336);
or U24192 (N_24192,N_23182,N_22897);
nand U24193 (N_24193,N_23550,N_23528);
nand U24194 (N_24194,N_23204,N_22827);
or U24195 (N_24195,N_23972,N_23681);
xor U24196 (N_24196,N_23060,N_23931);
or U24197 (N_24197,N_23532,N_23530);
or U24198 (N_24198,N_23651,N_23851);
xor U24199 (N_24199,N_23984,N_22895);
and U24200 (N_24200,N_23547,N_23431);
nor U24201 (N_24201,N_23559,N_23996);
or U24202 (N_24202,N_23176,N_23331);
and U24203 (N_24203,N_23325,N_22943);
and U24204 (N_24204,N_23496,N_23322);
xor U24205 (N_24205,N_23208,N_23558);
and U24206 (N_24206,N_23973,N_23817);
nor U24207 (N_24207,N_23229,N_23471);
nor U24208 (N_24208,N_23865,N_23396);
and U24209 (N_24209,N_23313,N_23272);
nor U24210 (N_24210,N_23672,N_23188);
nor U24211 (N_24211,N_23634,N_23372);
xor U24212 (N_24212,N_23036,N_22991);
or U24213 (N_24213,N_23368,N_23180);
nand U24214 (N_24214,N_23492,N_23116);
nor U24215 (N_24215,N_23770,N_23628);
xor U24216 (N_24216,N_23381,N_23491);
or U24217 (N_24217,N_23075,N_23106);
xor U24218 (N_24218,N_23024,N_22978);
or U24219 (N_24219,N_23546,N_23262);
nand U24220 (N_24220,N_22856,N_23577);
nand U24221 (N_24221,N_23145,N_23683);
xnor U24222 (N_24222,N_23685,N_23571);
and U24223 (N_24223,N_23895,N_23502);
and U24224 (N_24224,N_23183,N_23067);
nand U24225 (N_24225,N_23100,N_23854);
nand U24226 (N_24226,N_23349,N_23333);
nor U24227 (N_24227,N_22989,N_23802);
nor U24228 (N_24228,N_22904,N_23473);
and U24229 (N_24229,N_23094,N_23989);
xor U24230 (N_24230,N_22834,N_23297);
and U24231 (N_24231,N_22921,N_23000);
xnor U24232 (N_24232,N_23495,N_23554);
or U24233 (N_24233,N_22957,N_22917);
nor U24234 (N_24234,N_22971,N_23643);
nor U24235 (N_24235,N_23909,N_22806);
xnor U24236 (N_24236,N_23522,N_23138);
nor U24237 (N_24237,N_23109,N_23543);
or U24238 (N_24238,N_23779,N_23914);
and U24239 (N_24239,N_23150,N_23942);
nand U24240 (N_24240,N_23605,N_23378);
xnor U24241 (N_24241,N_23273,N_23236);
nor U24242 (N_24242,N_23147,N_23595);
and U24243 (N_24243,N_23274,N_23117);
and U24244 (N_24244,N_23650,N_23406);
or U24245 (N_24245,N_23088,N_23430);
nor U24246 (N_24246,N_23140,N_23133);
or U24247 (N_24247,N_23460,N_22860);
or U24248 (N_24248,N_23638,N_23611);
nor U24249 (N_24249,N_23220,N_23511);
nand U24250 (N_24250,N_23811,N_23812);
or U24251 (N_24251,N_23438,N_23997);
nor U24252 (N_24252,N_23542,N_22970);
and U24253 (N_24253,N_22960,N_22840);
or U24254 (N_24254,N_23586,N_23798);
nor U24255 (N_24255,N_22914,N_23113);
xnor U24256 (N_24256,N_22893,N_23609);
nor U24257 (N_24257,N_23379,N_23990);
or U24258 (N_24258,N_23846,N_23187);
nand U24259 (N_24259,N_23834,N_23472);
and U24260 (N_24260,N_23384,N_23269);
and U24261 (N_24261,N_22873,N_22984);
nor U24262 (N_24262,N_23902,N_23825);
nand U24263 (N_24263,N_23437,N_22850);
or U24264 (N_24264,N_23675,N_23744);
and U24265 (N_24265,N_23722,N_23311);
nor U24266 (N_24266,N_23371,N_23086);
and U24267 (N_24267,N_23983,N_23418);
xnor U24268 (N_24268,N_22890,N_22858);
nor U24269 (N_24269,N_23750,N_23915);
nand U24270 (N_24270,N_23933,N_23889);
or U24271 (N_24271,N_23291,N_22995);
nand U24272 (N_24272,N_23062,N_23247);
or U24273 (N_24273,N_23775,N_22998);
and U24274 (N_24274,N_23321,N_23278);
and U24275 (N_24275,N_23156,N_23829);
xor U24276 (N_24276,N_23303,N_23552);
and U24277 (N_24277,N_23832,N_23690);
nor U24278 (N_24278,N_23845,N_23064);
and U24279 (N_24279,N_23513,N_23045);
or U24280 (N_24280,N_23590,N_23974);
nor U24281 (N_24281,N_23740,N_23344);
nand U24282 (N_24282,N_23177,N_22949);
xnor U24283 (N_24283,N_23469,N_23952);
nor U24284 (N_24284,N_23068,N_23110);
and U24285 (N_24285,N_23299,N_23730);
nor U24286 (N_24286,N_23207,N_23506);
and U24287 (N_24287,N_23570,N_23198);
or U24288 (N_24288,N_23488,N_23804);
xnor U24289 (N_24289,N_23337,N_23661);
and U24290 (N_24290,N_23173,N_23192);
or U24291 (N_24291,N_23739,N_23949);
nand U24292 (N_24292,N_23388,N_22837);
nor U24293 (N_24293,N_22818,N_22894);
nand U24294 (N_24294,N_23687,N_23591);
nand U24295 (N_24295,N_23993,N_23093);
and U24296 (N_24296,N_22965,N_22908);
or U24297 (N_24297,N_23248,N_23294);
nand U24298 (N_24298,N_23422,N_23809);
and U24299 (N_24299,N_23030,N_23830);
or U24300 (N_24300,N_23589,N_23223);
xor U24301 (N_24301,N_23359,N_22804);
nand U24302 (N_24302,N_23462,N_23099);
and U24303 (N_24303,N_23049,N_23882);
and U24304 (N_24304,N_22951,N_23508);
nand U24305 (N_24305,N_22861,N_22811);
nand U24306 (N_24306,N_23635,N_23119);
nor U24307 (N_24307,N_23044,N_23800);
and U24308 (N_24308,N_22812,N_23284);
xor U24309 (N_24309,N_23136,N_23219);
xor U24310 (N_24310,N_23158,N_23348);
nor U24311 (N_24311,N_23948,N_23601);
xor U24312 (N_24312,N_23903,N_23705);
nor U24313 (N_24313,N_23255,N_22905);
nor U24314 (N_24314,N_23789,N_23887);
or U24315 (N_24315,N_23402,N_23939);
nand U24316 (N_24316,N_22845,N_23090);
nor U24317 (N_24317,N_23610,N_23050);
or U24318 (N_24318,N_23487,N_23383);
and U24319 (N_24319,N_23969,N_22822);
or U24320 (N_24320,N_23489,N_23432);
and U24321 (N_24321,N_23465,N_23684);
nor U24322 (N_24322,N_23868,N_23154);
nand U24323 (N_24323,N_23877,N_23386);
nor U24324 (N_24324,N_23330,N_23126);
nand U24325 (N_24325,N_22977,N_23354);
xor U24326 (N_24326,N_23482,N_22902);
nor U24327 (N_24327,N_23665,N_22922);
nand U24328 (N_24328,N_23618,N_23793);
and U24329 (N_24329,N_23477,N_23310);
nor U24330 (N_24330,N_23046,N_23668);
nor U24331 (N_24331,N_23499,N_23701);
xor U24332 (N_24332,N_23102,N_22930);
or U24333 (N_24333,N_23353,N_23518);
and U24334 (N_24334,N_22877,N_23009);
nand U24335 (N_24335,N_23704,N_23467);
and U24336 (N_24336,N_23691,N_23478);
nor U24337 (N_24337,N_23824,N_23526);
xor U24338 (N_24338,N_23741,N_23822);
or U24339 (N_24339,N_23871,N_23317);
or U24340 (N_24340,N_23561,N_23385);
or U24341 (N_24341,N_23540,N_23794);
nand U24342 (N_24342,N_23370,N_23614);
or U24343 (N_24343,N_23747,N_23012);
xnor U24344 (N_24344,N_23298,N_23641);
nor U24345 (N_24345,N_23146,N_23091);
and U24346 (N_24346,N_22918,N_23128);
and U24347 (N_24347,N_23166,N_23924);
xnor U24348 (N_24348,N_23214,N_23814);
or U24349 (N_24349,N_22946,N_23416);
or U24350 (N_24350,N_23880,N_23455);
and U24351 (N_24351,N_22825,N_23185);
xnor U24352 (N_24352,N_23335,N_23870);
xor U24353 (N_24353,N_23254,N_22924);
nand U24354 (N_24354,N_23066,N_23096);
or U24355 (N_24355,N_23985,N_23721);
nand U24356 (N_24356,N_23988,N_23363);
xnor U24357 (N_24357,N_23639,N_23803);
and U24358 (N_24358,N_23596,N_23367);
and U24359 (N_24359,N_23007,N_23523);
xor U24360 (N_24360,N_23277,N_23548);
nor U24361 (N_24361,N_23617,N_23736);
xor U24362 (N_24362,N_23783,N_23538);
nand U24363 (N_24363,N_23503,N_23602);
nor U24364 (N_24364,N_23732,N_23837);
nand U24365 (N_24365,N_22882,N_23625);
or U24366 (N_24366,N_23689,N_22923);
nor U24367 (N_24367,N_23757,N_23928);
nor U24368 (N_24368,N_23749,N_23686);
or U24369 (N_24369,N_23676,N_23243);
nor U24370 (N_24370,N_23637,N_23282);
or U24371 (N_24371,N_23369,N_23200);
and U24372 (N_24372,N_23164,N_23662);
or U24373 (N_24373,N_22881,N_23257);
or U24374 (N_24374,N_22853,N_23719);
or U24375 (N_24375,N_23938,N_23245);
or U24376 (N_24376,N_22857,N_23464);
nand U24377 (N_24377,N_23856,N_22859);
nand U24378 (N_24378,N_22864,N_23507);
nor U24379 (N_24379,N_23318,N_23125);
or U24380 (N_24380,N_23633,N_23986);
or U24381 (N_24381,N_23782,N_23444);
or U24382 (N_24382,N_22954,N_23906);
or U24383 (N_24383,N_23097,N_22952);
nor U24384 (N_24384,N_23157,N_22892);
and U24385 (N_24385,N_23659,N_22809);
or U24386 (N_24386,N_23234,N_23267);
xor U24387 (N_24387,N_22876,N_23644);
nor U24388 (N_24388,N_23580,N_22992);
nand U24389 (N_24389,N_23089,N_23048);
and U24390 (N_24390,N_23014,N_23821);
xor U24391 (N_24391,N_23285,N_23762);
xnor U24392 (N_24392,N_23723,N_22966);
and U24393 (N_24393,N_23520,N_23941);
nor U24394 (N_24394,N_22848,N_23512);
or U24395 (N_24395,N_23196,N_23764);
nor U24396 (N_24396,N_22929,N_23603);
xor U24397 (N_24397,N_23015,N_23189);
nand U24398 (N_24398,N_23361,N_23346);
nand U24399 (N_24399,N_23073,N_22945);
xnor U24400 (N_24400,N_23640,N_22870);
and U24401 (N_24401,N_23820,N_23397);
or U24402 (N_24402,N_23836,N_23955);
and U24403 (N_24403,N_23624,N_23112);
or U24404 (N_24404,N_22981,N_23598);
nor U24405 (N_24405,N_23358,N_23790);
or U24406 (N_24406,N_23287,N_23424);
nand U24407 (N_24407,N_23936,N_23127);
and U24408 (N_24408,N_23940,N_22958);
or U24409 (N_24409,N_23801,N_23232);
or U24410 (N_24410,N_23866,N_23079);
and U24411 (N_24411,N_23579,N_23327);
nand U24412 (N_24412,N_23280,N_23405);
xnor U24413 (N_24413,N_23101,N_23295);
and U24414 (N_24414,N_23910,N_23838);
nor U24415 (N_24415,N_23649,N_23210);
and U24416 (N_24416,N_23930,N_23470);
nand U24417 (N_24417,N_23926,N_23884);
nand U24418 (N_24418,N_23053,N_23083);
and U24419 (N_24419,N_23037,N_23058);
nand U24420 (N_24420,N_23098,N_23338);
nand U24421 (N_24421,N_23679,N_23027);
nor U24422 (N_24422,N_22887,N_23259);
nor U24423 (N_24423,N_23737,N_23760);
xor U24424 (N_24424,N_22997,N_22844);
xnor U24425 (N_24425,N_23302,N_23588);
and U24426 (N_24426,N_23852,N_23534);
xor U24427 (N_24427,N_23599,N_23362);
nor U24428 (N_24428,N_23074,N_22878);
and U24429 (N_24429,N_23700,N_23847);
and U24430 (N_24430,N_23040,N_23753);
nand U24431 (N_24431,N_22866,N_23576);
xnor U24432 (N_24432,N_23400,N_23525);
nand U24433 (N_24433,N_23756,N_23951);
or U24434 (N_24434,N_23693,N_23475);
nand U24435 (N_24435,N_23316,N_23135);
nand U24436 (N_24436,N_23874,N_23131);
nor U24437 (N_24437,N_23954,N_23165);
and U24438 (N_24438,N_23428,N_23746);
nor U24439 (N_24439,N_23004,N_23698);
nor U24440 (N_24440,N_23403,N_22817);
xnor U24441 (N_24441,N_23305,N_23563);
and U24442 (N_24442,N_23163,N_23501);
nand U24443 (N_24443,N_23293,N_23519);
nand U24444 (N_24444,N_23813,N_22907);
xnor U24445 (N_24445,N_22816,N_23890);
nor U24446 (N_24446,N_22814,N_23483);
xnor U24447 (N_24447,N_23021,N_23244);
or U24448 (N_24448,N_23555,N_23544);
or U24449 (N_24449,N_23320,N_23619);
nand U24450 (N_24450,N_22936,N_23356);
nor U24451 (N_24451,N_23392,N_23252);
xnor U24452 (N_24452,N_22810,N_23260);
xor U24453 (N_24453,N_23907,N_23439);
or U24454 (N_24454,N_23268,N_23826);
xor U24455 (N_24455,N_23697,N_23632);
nor U24456 (N_24456,N_23151,N_22956);
and U24457 (N_24457,N_23872,N_23604);
or U24458 (N_24458,N_23841,N_23072);
nand U24459 (N_24459,N_23860,N_22820);
nor U24460 (N_24460,N_23778,N_23485);
or U24461 (N_24461,N_23205,N_23134);
nand U24462 (N_24462,N_23648,N_23161);
and U24463 (N_24463,N_23355,N_23560);
or U24464 (N_24464,N_23600,N_23713);
nor U24465 (N_24465,N_23326,N_23115);
or U24466 (N_24466,N_23673,N_23728);
and U24467 (N_24467,N_23398,N_23242);
or U24468 (N_24468,N_23833,N_23975);
xor U24469 (N_24469,N_23213,N_23527);
nand U24470 (N_24470,N_23893,N_23270);
nand U24471 (N_24471,N_23249,N_22836);
xor U24472 (N_24472,N_22839,N_23375);
and U24473 (N_24473,N_23033,N_23769);
or U24474 (N_24474,N_23922,N_23703);
xor U24475 (N_24475,N_23724,N_23863);
nor U24476 (N_24476,N_23702,N_22896);
xor U24477 (N_24477,N_23221,N_23433);
or U24478 (N_24478,N_23263,N_23862);
nor U24479 (N_24479,N_22819,N_23306);
and U24480 (N_24480,N_22931,N_23962);
or U24481 (N_24481,N_23584,N_23013);
or U24482 (N_24482,N_23057,N_22926);
and U24483 (N_24483,N_23380,N_23788);
xor U24484 (N_24484,N_23733,N_23504);
nor U24485 (N_24485,N_23516,N_22982);
xor U24486 (N_24486,N_23708,N_23929);
nor U24487 (N_24487,N_22874,N_23005);
nand U24488 (N_24488,N_23051,N_23461);
nor U24489 (N_24489,N_23231,N_22939);
nor U24490 (N_24490,N_22899,N_23897);
xnor U24491 (N_24491,N_23329,N_23981);
xor U24492 (N_24492,N_22999,N_22994);
or U24493 (N_24493,N_23498,N_23763);
and U24494 (N_24494,N_23593,N_23479);
and U24495 (N_24495,N_23289,N_23043);
xor U24496 (N_24496,N_23038,N_23446);
nand U24497 (N_24497,N_23953,N_23468);
nor U24498 (N_24498,N_23077,N_23966);
nand U24499 (N_24499,N_23842,N_23606);
xnor U24500 (N_24500,N_23332,N_22983);
or U24501 (N_24501,N_22915,N_22808);
or U24502 (N_24502,N_23225,N_23957);
nand U24503 (N_24503,N_23120,N_23328);
nand U24504 (N_24504,N_23916,N_23288);
and U24505 (N_24505,N_23016,N_23006);
and U24506 (N_24506,N_23261,N_22851);
and U24507 (N_24507,N_23919,N_23410);
and U24508 (N_24508,N_22830,N_23658);
nor U24509 (N_24509,N_23224,N_23911);
and U24510 (N_24510,N_23773,N_23616);
and U24511 (N_24511,N_23440,N_22962);
and U24512 (N_24512,N_23859,N_22933);
nor U24513 (N_24513,N_23991,N_23199);
nand U24514 (N_24514,N_23787,N_23805);
nand U24515 (N_24515,N_22967,N_23608);
nor U24516 (N_24516,N_23191,N_23148);
and U24517 (N_24517,N_23419,N_23810);
or U24518 (N_24518,N_23393,N_23449);
xnor U24519 (N_24519,N_23565,N_23720);
nor U24520 (N_24520,N_23153,N_23725);
or U24521 (N_24521,N_23574,N_22959);
xnor U24522 (N_24522,N_22996,N_23085);
and U24523 (N_24523,N_23536,N_23995);
and U24524 (N_24524,N_23216,N_23674);
or U24525 (N_24525,N_23670,N_23032);
and U24526 (N_24526,N_23647,N_23869);
and U24527 (N_24527,N_23767,N_23304);
xor U24528 (N_24528,N_22833,N_23857);
nor U24529 (N_24529,N_23835,N_23920);
nand U24530 (N_24530,N_23360,N_23481);
and U24531 (N_24531,N_22842,N_23556);
nor U24532 (N_24532,N_23484,N_23105);
nand U24533 (N_24533,N_23042,N_23152);
nor U24534 (N_24534,N_22973,N_23968);
or U24535 (N_24535,N_22953,N_23301);
nor U24536 (N_24536,N_22841,N_23786);
xor U24537 (N_24537,N_23524,N_22824);
nand U24538 (N_24538,N_22988,N_23971);
and U24539 (N_24539,N_23575,N_23905);
nand U24540 (N_24540,N_23343,N_23312);
xor U24541 (N_24541,N_23023,N_23977);
nand U24542 (N_24542,N_23211,N_23103);
xnor U24543 (N_24543,N_23286,N_22815);
nand U24544 (N_24544,N_23758,N_22909);
and U24545 (N_24545,N_23898,N_23387);
xnor U24546 (N_24546,N_23828,N_23427);
and U24547 (N_24547,N_23636,N_23408);
nand U24548 (N_24548,N_23956,N_23300);
nor U24549 (N_24549,N_22888,N_23706);
or U24550 (N_24550,N_23766,N_23411);
nor U24551 (N_24551,N_23071,N_23539);
or U24552 (N_24552,N_22948,N_22961);
nor U24553 (N_24553,N_23726,N_23652);
xor U24554 (N_24554,N_23840,N_22934);
nand U24555 (N_24555,N_23875,N_22843);
or U24556 (N_24556,N_23001,N_23537);
nand U24557 (N_24557,N_23389,N_23963);
or U24558 (N_24558,N_23429,N_23041);
xnor U24559 (N_24559,N_23867,N_23992);
xor U24560 (N_24560,N_23780,N_22947);
and U24561 (N_24561,N_23692,N_23678);
or U24562 (N_24562,N_23132,N_23795);
nand U24563 (N_24563,N_23935,N_23059);
xnor U24564 (N_24564,N_22964,N_23459);
nand U24565 (N_24565,N_22974,N_23054);
xor U24566 (N_24566,N_23549,N_23923);
or U24567 (N_24567,N_23376,N_23352);
nor U24568 (N_24568,N_23751,N_23497);
and U24569 (N_24569,N_23407,N_23445);
xor U24570 (N_24570,N_23567,N_23366);
nand U24571 (N_24571,N_23025,N_23443);
or U24572 (N_24572,N_23202,N_23195);
or U24573 (N_24573,N_23087,N_23943);
and U24574 (N_24574,N_23765,N_23451);
and U24575 (N_24575,N_23861,N_23921);
nor U24576 (N_24576,N_23660,N_23900);
nor U24577 (N_24577,N_23777,N_23017);
and U24578 (N_24578,N_23063,N_23656);
and U24579 (N_24579,N_23026,N_23885);
and U24580 (N_24580,N_22846,N_23341);
or U24581 (N_24581,N_23002,N_23707);
or U24582 (N_24582,N_23912,N_23415);
or U24583 (N_24583,N_23597,N_23994);
and U24584 (N_24584,N_23785,N_23092);
nand U24585 (N_24585,N_23271,N_22871);
or U24586 (N_24586,N_23480,N_23342);
xor U24587 (N_24587,N_23076,N_23655);
and U24588 (N_24588,N_23500,N_23743);
nand U24589 (N_24589,N_23008,N_23233);
or U24590 (N_24590,N_23209,N_23029);
xor U24591 (N_24591,N_22855,N_22869);
nor U24592 (N_24592,N_23653,N_23227);
nor U24593 (N_24593,N_22800,N_23456);
and U24594 (N_24594,N_23486,N_23533);
xor U24595 (N_24595,N_23615,N_23844);
nand U24596 (N_24596,N_23818,N_22937);
and U24597 (N_24597,N_22985,N_22980);
or U24598 (N_24598,N_23585,N_23729);
or U24599 (N_24599,N_22940,N_23279);
and U24600 (N_24600,N_23803,N_23906);
or U24601 (N_24601,N_23598,N_23517);
or U24602 (N_24602,N_22814,N_23304);
or U24603 (N_24603,N_22958,N_23830);
xor U24604 (N_24604,N_23156,N_23033);
nor U24605 (N_24605,N_23385,N_23776);
nand U24606 (N_24606,N_23082,N_23621);
or U24607 (N_24607,N_23742,N_23331);
nor U24608 (N_24608,N_23691,N_23592);
nor U24609 (N_24609,N_23072,N_23960);
or U24610 (N_24610,N_23982,N_23644);
or U24611 (N_24611,N_23264,N_23081);
nand U24612 (N_24612,N_22965,N_23108);
xnor U24613 (N_24613,N_23893,N_23281);
or U24614 (N_24614,N_23659,N_23036);
and U24615 (N_24615,N_23964,N_23230);
nor U24616 (N_24616,N_22847,N_23906);
and U24617 (N_24617,N_23095,N_22974);
xor U24618 (N_24618,N_23079,N_23257);
or U24619 (N_24619,N_22912,N_23507);
and U24620 (N_24620,N_23340,N_23907);
nand U24621 (N_24621,N_23441,N_23075);
nor U24622 (N_24622,N_22921,N_23847);
xnor U24623 (N_24623,N_23114,N_23268);
or U24624 (N_24624,N_23784,N_23283);
nor U24625 (N_24625,N_23035,N_22917);
nor U24626 (N_24626,N_23811,N_23661);
and U24627 (N_24627,N_23982,N_23781);
xor U24628 (N_24628,N_23595,N_23717);
nand U24629 (N_24629,N_23343,N_23881);
and U24630 (N_24630,N_23734,N_23985);
xor U24631 (N_24631,N_23967,N_23169);
and U24632 (N_24632,N_23132,N_23994);
xor U24633 (N_24633,N_23354,N_23910);
nand U24634 (N_24634,N_23987,N_23838);
and U24635 (N_24635,N_23438,N_23864);
nand U24636 (N_24636,N_23377,N_23441);
nand U24637 (N_24637,N_23317,N_23038);
or U24638 (N_24638,N_23145,N_23082);
xor U24639 (N_24639,N_23881,N_23912);
xnor U24640 (N_24640,N_23749,N_23388);
nand U24641 (N_24641,N_22988,N_23760);
and U24642 (N_24642,N_23319,N_23503);
and U24643 (N_24643,N_23411,N_23031);
or U24644 (N_24644,N_23308,N_23828);
xnor U24645 (N_24645,N_23481,N_23076);
xnor U24646 (N_24646,N_23862,N_23740);
xor U24647 (N_24647,N_23079,N_23023);
and U24648 (N_24648,N_23206,N_23725);
xor U24649 (N_24649,N_23471,N_23147);
nor U24650 (N_24650,N_22969,N_23420);
xor U24651 (N_24651,N_23172,N_22847);
xor U24652 (N_24652,N_23181,N_23109);
nor U24653 (N_24653,N_23514,N_23009);
and U24654 (N_24654,N_23578,N_23906);
xnor U24655 (N_24655,N_23347,N_23403);
xnor U24656 (N_24656,N_22913,N_23298);
nor U24657 (N_24657,N_23148,N_23719);
or U24658 (N_24658,N_22969,N_23077);
and U24659 (N_24659,N_23693,N_23545);
xor U24660 (N_24660,N_23360,N_22978);
or U24661 (N_24661,N_23128,N_22855);
or U24662 (N_24662,N_23864,N_23310);
or U24663 (N_24663,N_22892,N_23696);
and U24664 (N_24664,N_23470,N_23570);
and U24665 (N_24665,N_23592,N_23184);
or U24666 (N_24666,N_23781,N_23535);
nand U24667 (N_24667,N_23864,N_22840);
nand U24668 (N_24668,N_22881,N_23788);
nor U24669 (N_24669,N_23731,N_23215);
nand U24670 (N_24670,N_23466,N_23758);
nand U24671 (N_24671,N_23697,N_23086);
nor U24672 (N_24672,N_23205,N_23163);
nor U24673 (N_24673,N_22967,N_23471);
nor U24674 (N_24674,N_23519,N_23451);
xor U24675 (N_24675,N_23456,N_23523);
and U24676 (N_24676,N_23189,N_22980);
nor U24677 (N_24677,N_23688,N_23479);
and U24678 (N_24678,N_23878,N_23605);
and U24679 (N_24679,N_22872,N_23554);
nand U24680 (N_24680,N_23095,N_23114);
nor U24681 (N_24681,N_23903,N_23707);
and U24682 (N_24682,N_23218,N_22990);
and U24683 (N_24683,N_23332,N_23910);
xor U24684 (N_24684,N_23964,N_23956);
and U24685 (N_24685,N_23847,N_23064);
or U24686 (N_24686,N_23894,N_23252);
nand U24687 (N_24687,N_23980,N_23042);
nor U24688 (N_24688,N_23412,N_23950);
nor U24689 (N_24689,N_23844,N_22869);
xor U24690 (N_24690,N_23532,N_23498);
nor U24691 (N_24691,N_22936,N_23650);
and U24692 (N_24692,N_23737,N_23215);
and U24693 (N_24693,N_22993,N_23776);
and U24694 (N_24694,N_23313,N_23564);
or U24695 (N_24695,N_23728,N_23958);
nand U24696 (N_24696,N_23959,N_23288);
or U24697 (N_24697,N_23793,N_22920);
or U24698 (N_24698,N_23777,N_23131);
xor U24699 (N_24699,N_22995,N_23577);
and U24700 (N_24700,N_23383,N_23278);
xnor U24701 (N_24701,N_23193,N_23121);
and U24702 (N_24702,N_23907,N_23723);
nor U24703 (N_24703,N_23130,N_22986);
nor U24704 (N_24704,N_23326,N_23991);
or U24705 (N_24705,N_23081,N_23956);
or U24706 (N_24706,N_23586,N_23067);
or U24707 (N_24707,N_23747,N_22864);
and U24708 (N_24708,N_23596,N_23486);
nand U24709 (N_24709,N_22833,N_22871);
nor U24710 (N_24710,N_23822,N_23705);
nand U24711 (N_24711,N_23152,N_23673);
nand U24712 (N_24712,N_23916,N_23292);
xor U24713 (N_24713,N_23800,N_23414);
or U24714 (N_24714,N_23729,N_23350);
nand U24715 (N_24715,N_23466,N_23380);
xnor U24716 (N_24716,N_23056,N_22920);
xor U24717 (N_24717,N_23492,N_23202);
nor U24718 (N_24718,N_23210,N_23053);
or U24719 (N_24719,N_23801,N_23067);
xnor U24720 (N_24720,N_23702,N_23569);
or U24721 (N_24721,N_23091,N_23213);
and U24722 (N_24722,N_23534,N_23463);
or U24723 (N_24723,N_23910,N_23780);
or U24724 (N_24724,N_23198,N_22975);
xor U24725 (N_24725,N_23616,N_23810);
or U24726 (N_24726,N_22885,N_23595);
or U24727 (N_24727,N_23370,N_23634);
xnor U24728 (N_24728,N_23334,N_23338);
nor U24729 (N_24729,N_23229,N_22994);
and U24730 (N_24730,N_23531,N_23540);
or U24731 (N_24731,N_23431,N_23773);
nor U24732 (N_24732,N_23233,N_23205);
or U24733 (N_24733,N_22950,N_23863);
xor U24734 (N_24734,N_22815,N_23816);
and U24735 (N_24735,N_23988,N_22850);
xor U24736 (N_24736,N_23145,N_22901);
or U24737 (N_24737,N_22876,N_22842);
nand U24738 (N_24738,N_23069,N_23875);
xor U24739 (N_24739,N_23716,N_23017);
and U24740 (N_24740,N_22865,N_23629);
nand U24741 (N_24741,N_23230,N_23494);
nand U24742 (N_24742,N_23272,N_23185);
nand U24743 (N_24743,N_23872,N_22958);
or U24744 (N_24744,N_23227,N_23124);
xor U24745 (N_24745,N_23896,N_23399);
xnor U24746 (N_24746,N_23167,N_23750);
and U24747 (N_24747,N_23390,N_23423);
nand U24748 (N_24748,N_23071,N_23401);
and U24749 (N_24749,N_22813,N_23950);
nor U24750 (N_24750,N_23994,N_23631);
nor U24751 (N_24751,N_23551,N_23712);
nor U24752 (N_24752,N_23988,N_23688);
xor U24753 (N_24753,N_23902,N_23154);
or U24754 (N_24754,N_23801,N_23524);
and U24755 (N_24755,N_23538,N_23998);
nor U24756 (N_24756,N_23025,N_23469);
and U24757 (N_24757,N_23961,N_23182);
nand U24758 (N_24758,N_22928,N_23619);
nor U24759 (N_24759,N_23211,N_23872);
or U24760 (N_24760,N_22877,N_23762);
and U24761 (N_24761,N_23957,N_23627);
or U24762 (N_24762,N_23057,N_22979);
nor U24763 (N_24763,N_23136,N_23447);
nor U24764 (N_24764,N_23324,N_23368);
and U24765 (N_24765,N_23078,N_23510);
xnor U24766 (N_24766,N_23729,N_23448);
nand U24767 (N_24767,N_22855,N_23125);
nand U24768 (N_24768,N_23989,N_23134);
nand U24769 (N_24769,N_22827,N_23898);
xnor U24770 (N_24770,N_23561,N_23844);
nand U24771 (N_24771,N_23991,N_23197);
nor U24772 (N_24772,N_23867,N_23668);
xor U24773 (N_24773,N_23392,N_23824);
nand U24774 (N_24774,N_22809,N_23196);
or U24775 (N_24775,N_23990,N_23204);
nor U24776 (N_24776,N_23201,N_23819);
nor U24777 (N_24777,N_23953,N_23442);
nand U24778 (N_24778,N_23801,N_22919);
and U24779 (N_24779,N_23494,N_23093);
or U24780 (N_24780,N_23979,N_23135);
xor U24781 (N_24781,N_23465,N_23740);
or U24782 (N_24782,N_22885,N_22999);
xnor U24783 (N_24783,N_22864,N_23897);
xor U24784 (N_24784,N_22947,N_23323);
nand U24785 (N_24785,N_23124,N_23383);
and U24786 (N_24786,N_23759,N_23771);
nand U24787 (N_24787,N_23597,N_23323);
nand U24788 (N_24788,N_23140,N_23502);
nor U24789 (N_24789,N_23865,N_23696);
nor U24790 (N_24790,N_23423,N_23093);
or U24791 (N_24791,N_23688,N_22802);
nor U24792 (N_24792,N_23157,N_23231);
xor U24793 (N_24793,N_23891,N_23291);
or U24794 (N_24794,N_23585,N_23854);
and U24795 (N_24795,N_23075,N_22982);
xnor U24796 (N_24796,N_23516,N_23610);
nor U24797 (N_24797,N_22821,N_23824);
and U24798 (N_24798,N_23409,N_23919);
nand U24799 (N_24799,N_23440,N_23818);
nand U24800 (N_24800,N_23672,N_22918);
or U24801 (N_24801,N_23180,N_23459);
and U24802 (N_24802,N_23852,N_23491);
nand U24803 (N_24803,N_23853,N_23067);
nor U24804 (N_24804,N_23995,N_23793);
nand U24805 (N_24805,N_22805,N_23394);
nor U24806 (N_24806,N_22877,N_23793);
nand U24807 (N_24807,N_23359,N_23809);
nor U24808 (N_24808,N_23341,N_23576);
and U24809 (N_24809,N_23485,N_23027);
nor U24810 (N_24810,N_23909,N_23855);
or U24811 (N_24811,N_23620,N_23355);
nand U24812 (N_24812,N_23715,N_22871);
xnor U24813 (N_24813,N_23298,N_22847);
nand U24814 (N_24814,N_23232,N_23344);
nor U24815 (N_24815,N_23289,N_23522);
xnor U24816 (N_24816,N_23145,N_23486);
nor U24817 (N_24817,N_22869,N_23644);
or U24818 (N_24818,N_23115,N_23637);
or U24819 (N_24819,N_23449,N_23291);
or U24820 (N_24820,N_23942,N_23520);
nand U24821 (N_24821,N_23134,N_23704);
nor U24822 (N_24822,N_23706,N_22894);
or U24823 (N_24823,N_23622,N_23131);
or U24824 (N_24824,N_23965,N_23710);
or U24825 (N_24825,N_23996,N_22817);
xor U24826 (N_24826,N_22922,N_23668);
or U24827 (N_24827,N_23895,N_23935);
xnor U24828 (N_24828,N_23146,N_23443);
and U24829 (N_24829,N_23143,N_23614);
nand U24830 (N_24830,N_23536,N_23334);
nor U24831 (N_24831,N_23742,N_22809);
xor U24832 (N_24832,N_23684,N_23064);
and U24833 (N_24833,N_23515,N_22933);
or U24834 (N_24834,N_23221,N_23218);
or U24835 (N_24835,N_23623,N_23499);
and U24836 (N_24836,N_23578,N_23342);
and U24837 (N_24837,N_23659,N_23046);
and U24838 (N_24838,N_23129,N_23198);
and U24839 (N_24839,N_22912,N_23186);
nand U24840 (N_24840,N_22972,N_23499);
xnor U24841 (N_24841,N_23841,N_22949);
nor U24842 (N_24842,N_23277,N_23855);
xor U24843 (N_24843,N_23317,N_22912);
nor U24844 (N_24844,N_23312,N_23716);
and U24845 (N_24845,N_23913,N_22915);
and U24846 (N_24846,N_23039,N_23864);
nand U24847 (N_24847,N_23974,N_23998);
and U24848 (N_24848,N_22816,N_23356);
and U24849 (N_24849,N_23043,N_23113);
xor U24850 (N_24850,N_23842,N_23954);
and U24851 (N_24851,N_23618,N_23260);
xnor U24852 (N_24852,N_23127,N_23926);
and U24853 (N_24853,N_23281,N_23109);
or U24854 (N_24854,N_23203,N_22965);
nand U24855 (N_24855,N_23779,N_23929);
and U24856 (N_24856,N_23538,N_22943);
nand U24857 (N_24857,N_22944,N_23820);
xnor U24858 (N_24858,N_23298,N_23566);
xnor U24859 (N_24859,N_23238,N_22812);
or U24860 (N_24860,N_23891,N_22889);
and U24861 (N_24861,N_23737,N_23063);
and U24862 (N_24862,N_23276,N_23247);
nor U24863 (N_24863,N_23622,N_23406);
xnor U24864 (N_24864,N_22917,N_23978);
and U24865 (N_24865,N_22937,N_23113);
nor U24866 (N_24866,N_23187,N_23543);
nor U24867 (N_24867,N_23967,N_23269);
or U24868 (N_24868,N_23730,N_23569);
nor U24869 (N_24869,N_22997,N_23557);
and U24870 (N_24870,N_22918,N_23430);
nor U24871 (N_24871,N_23342,N_23527);
nand U24872 (N_24872,N_23812,N_23486);
or U24873 (N_24873,N_22820,N_23399);
and U24874 (N_24874,N_23182,N_23853);
and U24875 (N_24875,N_22804,N_23331);
and U24876 (N_24876,N_23587,N_23552);
nor U24877 (N_24877,N_23567,N_23978);
and U24878 (N_24878,N_23360,N_23873);
and U24879 (N_24879,N_22804,N_23546);
and U24880 (N_24880,N_23423,N_23631);
nand U24881 (N_24881,N_23548,N_23840);
and U24882 (N_24882,N_23543,N_23913);
nand U24883 (N_24883,N_22999,N_23645);
or U24884 (N_24884,N_23829,N_23010);
xnor U24885 (N_24885,N_22997,N_23129);
xor U24886 (N_24886,N_23116,N_23358);
nand U24887 (N_24887,N_23920,N_23763);
nand U24888 (N_24888,N_23081,N_22884);
or U24889 (N_24889,N_22897,N_23808);
and U24890 (N_24890,N_22922,N_23855);
and U24891 (N_24891,N_23296,N_23292);
and U24892 (N_24892,N_22833,N_23787);
or U24893 (N_24893,N_23466,N_23096);
xor U24894 (N_24894,N_23255,N_23546);
or U24895 (N_24895,N_23293,N_23963);
and U24896 (N_24896,N_23684,N_23156);
or U24897 (N_24897,N_23172,N_23440);
nor U24898 (N_24898,N_23258,N_23117);
or U24899 (N_24899,N_23141,N_23658);
nand U24900 (N_24900,N_23056,N_22836);
nor U24901 (N_24901,N_23983,N_23388);
or U24902 (N_24902,N_23540,N_23408);
xnor U24903 (N_24903,N_23123,N_22862);
xnor U24904 (N_24904,N_23428,N_23665);
nor U24905 (N_24905,N_23327,N_23133);
or U24906 (N_24906,N_23868,N_23299);
nor U24907 (N_24907,N_23456,N_23023);
nor U24908 (N_24908,N_23744,N_23614);
or U24909 (N_24909,N_23400,N_23109);
nor U24910 (N_24910,N_23116,N_23466);
or U24911 (N_24911,N_23537,N_23726);
nand U24912 (N_24912,N_23828,N_23589);
xor U24913 (N_24913,N_23173,N_22954);
or U24914 (N_24914,N_22947,N_23240);
nand U24915 (N_24915,N_23338,N_23557);
and U24916 (N_24916,N_23719,N_23129);
or U24917 (N_24917,N_23532,N_23788);
xnor U24918 (N_24918,N_23570,N_23416);
nand U24919 (N_24919,N_23829,N_23828);
nand U24920 (N_24920,N_23253,N_23005);
nor U24921 (N_24921,N_23754,N_23782);
nor U24922 (N_24922,N_23318,N_22933);
or U24923 (N_24923,N_23081,N_23315);
and U24924 (N_24924,N_23321,N_22822);
nor U24925 (N_24925,N_22867,N_23612);
nor U24926 (N_24926,N_23630,N_23869);
or U24927 (N_24927,N_22903,N_23480);
or U24928 (N_24928,N_22881,N_22941);
nand U24929 (N_24929,N_23683,N_23152);
nand U24930 (N_24930,N_23524,N_22917);
and U24931 (N_24931,N_23982,N_23242);
nor U24932 (N_24932,N_23540,N_22879);
nor U24933 (N_24933,N_23595,N_23307);
or U24934 (N_24934,N_23467,N_23300);
and U24935 (N_24935,N_22984,N_22917);
xor U24936 (N_24936,N_23755,N_23917);
xnor U24937 (N_24937,N_22952,N_23541);
xor U24938 (N_24938,N_23999,N_23339);
nand U24939 (N_24939,N_23153,N_23849);
nand U24940 (N_24940,N_23930,N_23255);
nor U24941 (N_24941,N_23757,N_23490);
and U24942 (N_24942,N_23331,N_23478);
and U24943 (N_24943,N_23087,N_23860);
xnor U24944 (N_24944,N_23433,N_23030);
xor U24945 (N_24945,N_22818,N_22884);
nor U24946 (N_24946,N_23360,N_23277);
nand U24947 (N_24947,N_23794,N_22900);
nor U24948 (N_24948,N_23537,N_23629);
and U24949 (N_24949,N_23581,N_23925);
and U24950 (N_24950,N_23509,N_23553);
nand U24951 (N_24951,N_22967,N_23040);
nor U24952 (N_24952,N_23844,N_23305);
xor U24953 (N_24953,N_23837,N_23145);
or U24954 (N_24954,N_23496,N_23753);
and U24955 (N_24955,N_23605,N_23505);
and U24956 (N_24956,N_23465,N_23223);
or U24957 (N_24957,N_23867,N_23567);
and U24958 (N_24958,N_23528,N_23997);
nand U24959 (N_24959,N_23082,N_23887);
and U24960 (N_24960,N_23731,N_23879);
or U24961 (N_24961,N_23265,N_22842);
nor U24962 (N_24962,N_23707,N_23323);
or U24963 (N_24963,N_22854,N_22826);
nand U24964 (N_24964,N_23984,N_22898);
xor U24965 (N_24965,N_22919,N_23044);
nor U24966 (N_24966,N_23033,N_23629);
and U24967 (N_24967,N_23431,N_23601);
xnor U24968 (N_24968,N_23245,N_23022);
and U24969 (N_24969,N_23202,N_22853);
xnor U24970 (N_24970,N_23081,N_23687);
nor U24971 (N_24971,N_23849,N_23537);
xnor U24972 (N_24972,N_23911,N_23908);
or U24973 (N_24973,N_23647,N_23811);
or U24974 (N_24974,N_23544,N_23831);
nor U24975 (N_24975,N_22917,N_23862);
xor U24976 (N_24976,N_23679,N_23536);
or U24977 (N_24977,N_23029,N_23092);
xnor U24978 (N_24978,N_23919,N_23166);
xor U24979 (N_24979,N_22827,N_23870);
or U24980 (N_24980,N_23019,N_23630);
nor U24981 (N_24981,N_23187,N_23618);
nor U24982 (N_24982,N_23064,N_22972);
or U24983 (N_24983,N_23318,N_23829);
nand U24984 (N_24984,N_23884,N_23741);
and U24985 (N_24985,N_23473,N_22855);
xnor U24986 (N_24986,N_22893,N_23086);
and U24987 (N_24987,N_23661,N_22978);
or U24988 (N_24988,N_23799,N_23581);
xnor U24989 (N_24989,N_23216,N_23130);
xor U24990 (N_24990,N_22926,N_23950);
and U24991 (N_24991,N_23649,N_23874);
xor U24992 (N_24992,N_23070,N_23727);
or U24993 (N_24993,N_23040,N_23259);
or U24994 (N_24994,N_23292,N_22909);
xnor U24995 (N_24995,N_23355,N_23153);
and U24996 (N_24996,N_23598,N_23021);
or U24997 (N_24997,N_23430,N_23264);
and U24998 (N_24998,N_23621,N_23050);
or U24999 (N_24999,N_23128,N_23293);
nand U25000 (N_25000,N_23060,N_23593);
nor U25001 (N_25001,N_22958,N_23699);
xor U25002 (N_25002,N_23168,N_23600);
nor U25003 (N_25003,N_22865,N_23012);
xnor U25004 (N_25004,N_23973,N_23830);
and U25005 (N_25005,N_23757,N_22975);
nand U25006 (N_25006,N_23210,N_23320);
and U25007 (N_25007,N_23812,N_23236);
or U25008 (N_25008,N_23756,N_23164);
and U25009 (N_25009,N_23413,N_23719);
nor U25010 (N_25010,N_23719,N_22969);
and U25011 (N_25011,N_23797,N_23398);
and U25012 (N_25012,N_23363,N_23534);
xor U25013 (N_25013,N_23640,N_23121);
nor U25014 (N_25014,N_23719,N_23116);
xnor U25015 (N_25015,N_23808,N_23146);
xor U25016 (N_25016,N_23275,N_23427);
xnor U25017 (N_25017,N_23024,N_23768);
xnor U25018 (N_25018,N_23207,N_23194);
or U25019 (N_25019,N_23212,N_23515);
or U25020 (N_25020,N_23831,N_23400);
nand U25021 (N_25021,N_23229,N_23033);
xnor U25022 (N_25022,N_23725,N_23008);
xnor U25023 (N_25023,N_23651,N_23329);
nand U25024 (N_25024,N_23288,N_23822);
nor U25025 (N_25025,N_23638,N_22963);
nor U25026 (N_25026,N_23486,N_23571);
or U25027 (N_25027,N_23529,N_23549);
xnor U25028 (N_25028,N_23548,N_23977);
nor U25029 (N_25029,N_22821,N_23851);
xnor U25030 (N_25030,N_23235,N_23212);
and U25031 (N_25031,N_23790,N_22963);
xnor U25032 (N_25032,N_23247,N_23069);
and U25033 (N_25033,N_23269,N_23875);
and U25034 (N_25034,N_23791,N_23723);
xor U25035 (N_25035,N_22952,N_23975);
and U25036 (N_25036,N_22994,N_23145);
xnor U25037 (N_25037,N_23452,N_23158);
and U25038 (N_25038,N_23269,N_23500);
or U25039 (N_25039,N_23235,N_23196);
or U25040 (N_25040,N_23041,N_23516);
nand U25041 (N_25041,N_23642,N_23181);
or U25042 (N_25042,N_23524,N_22886);
xnor U25043 (N_25043,N_23127,N_23247);
nor U25044 (N_25044,N_22937,N_23027);
and U25045 (N_25045,N_23173,N_23332);
and U25046 (N_25046,N_23544,N_23584);
or U25047 (N_25047,N_23080,N_23184);
or U25048 (N_25048,N_22949,N_23691);
nor U25049 (N_25049,N_23078,N_23827);
and U25050 (N_25050,N_23335,N_23965);
xor U25051 (N_25051,N_23507,N_23038);
or U25052 (N_25052,N_23437,N_23098);
xor U25053 (N_25053,N_23695,N_22819);
and U25054 (N_25054,N_23649,N_23889);
and U25055 (N_25055,N_22937,N_23268);
nand U25056 (N_25056,N_23157,N_23847);
or U25057 (N_25057,N_23731,N_23252);
xor U25058 (N_25058,N_23520,N_23126);
or U25059 (N_25059,N_22851,N_23228);
nand U25060 (N_25060,N_23760,N_23945);
nor U25061 (N_25061,N_22995,N_23661);
xor U25062 (N_25062,N_23678,N_23479);
and U25063 (N_25063,N_23298,N_23153);
and U25064 (N_25064,N_22838,N_23209);
or U25065 (N_25065,N_23496,N_23158);
or U25066 (N_25066,N_23983,N_23319);
xor U25067 (N_25067,N_23719,N_23642);
xnor U25068 (N_25068,N_23571,N_23930);
nor U25069 (N_25069,N_23268,N_23893);
xnor U25070 (N_25070,N_23473,N_23682);
and U25071 (N_25071,N_23107,N_23819);
xor U25072 (N_25072,N_22867,N_23945);
and U25073 (N_25073,N_22808,N_22811);
nor U25074 (N_25074,N_22839,N_23845);
or U25075 (N_25075,N_23536,N_23934);
xnor U25076 (N_25076,N_23688,N_23064);
nand U25077 (N_25077,N_23553,N_23377);
nand U25078 (N_25078,N_22876,N_23228);
nor U25079 (N_25079,N_23352,N_23137);
nand U25080 (N_25080,N_23008,N_23260);
xnor U25081 (N_25081,N_23354,N_23331);
or U25082 (N_25082,N_23265,N_23533);
xor U25083 (N_25083,N_22946,N_22868);
xnor U25084 (N_25084,N_23354,N_23852);
and U25085 (N_25085,N_23225,N_23207);
nor U25086 (N_25086,N_23579,N_23371);
nor U25087 (N_25087,N_23380,N_23683);
xor U25088 (N_25088,N_22952,N_23255);
nand U25089 (N_25089,N_22965,N_22830);
nand U25090 (N_25090,N_23162,N_23113);
and U25091 (N_25091,N_23366,N_23924);
nor U25092 (N_25092,N_23634,N_23545);
xnor U25093 (N_25093,N_22816,N_23088);
and U25094 (N_25094,N_23163,N_23431);
nand U25095 (N_25095,N_23964,N_23203);
and U25096 (N_25096,N_23511,N_23931);
and U25097 (N_25097,N_23386,N_23926);
xor U25098 (N_25098,N_23593,N_22959);
or U25099 (N_25099,N_23401,N_22904);
nor U25100 (N_25100,N_23525,N_23328);
nor U25101 (N_25101,N_23062,N_23498);
nor U25102 (N_25102,N_23270,N_23769);
xnor U25103 (N_25103,N_23700,N_23044);
xnor U25104 (N_25104,N_23442,N_23760);
nor U25105 (N_25105,N_23265,N_23835);
and U25106 (N_25106,N_23383,N_22906);
or U25107 (N_25107,N_22928,N_23155);
nand U25108 (N_25108,N_23993,N_23777);
nor U25109 (N_25109,N_23085,N_23662);
or U25110 (N_25110,N_23341,N_23207);
and U25111 (N_25111,N_23976,N_23679);
nor U25112 (N_25112,N_23861,N_22890);
xor U25113 (N_25113,N_23397,N_23124);
and U25114 (N_25114,N_23184,N_23270);
or U25115 (N_25115,N_23591,N_23825);
nor U25116 (N_25116,N_22826,N_23351);
nor U25117 (N_25117,N_23388,N_23408);
or U25118 (N_25118,N_23066,N_22904);
nand U25119 (N_25119,N_22813,N_23657);
nand U25120 (N_25120,N_23122,N_23859);
nand U25121 (N_25121,N_23244,N_23506);
or U25122 (N_25122,N_23112,N_23539);
nor U25123 (N_25123,N_23318,N_23057);
nand U25124 (N_25124,N_23296,N_22822);
nor U25125 (N_25125,N_23297,N_22982);
nand U25126 (N_25126,N_23035,N_23674);
nand U25127 (N_25127,N_23897,N_22839);
xnor U25128 (N_25128,N_23754,N_23881);
or U25129 (N_25129,N_23426,N_23404);
xor U25130 (N_25130,N_23143,N_23767);
or U25131 (N_25131,N_23800,N_23558);
or U25132 (N_25132,N_22834,N_23514);
and U25133 (N_25133,N_23308,N_23520);
xor U25134 (N_25134,N_23984,N_23117);
xnor U25135 (N_25135,N_23244,N_23573);
nand U25136 (N_25136,N_23014,N_23516);
nand U25137 (N_25137,N_23743,N_23338);
or U25138 (N_25138,N_23689,N_23744);
or U25139 (N_25139,N_23836,N_23321);
nand U25140 (N_25140,N_22975,N_23425);
nor U25141 (N_25141,N_23530,N_23266);
and U25142 (N_25142,N_23689,N_23012);
xor U25143 (N_25143,N_23282,N_23787);
nand U25144 (N_25144,N_23012,N_23578);
nand U25145 (N_25145,N_23086,N_23130);
nand U25146 (N_25146,N_22866,N_23116);
and U25147 (N_25147,N_23109,N_23927);
and U25148 (N_25148,N_23142,N_23828);
nand U25149 (N_25149,N_22817,N_23807);
nor U25150 (N_25150,N_23081,N_23435);
nand U25151 (N_25151,N_23672,N_23774);
or U25152 (N_25152,N_23995,N_23281);
or U25153 (N_25153,N_23069,N_23210);
nand U25154 (N_25154,N_22985,N_23228);
and U25155 (N_25155,N_23534,N_23715);
and U25156 (N_25156,N_22968,N_22891);
nor U25157 (N_25157,N_22859,N_23051);
or U25158 (N_25158,N_22897,N_23308);
nor U25159 (N_25159,N_23502,N_23035);
nand U25160 (N_25160,N_23564,N_23732);
xor U25161 (N_25161,N_23433,N_22885);
nand U25162 (N_25162,N_22888,N_23703);
nand U25163 (N_25163,N_23138,N_23947);
or U25164 (N_25164,N_23024,N_23376);
xor U25165 (N_25165,N_22912,N_23966);
or U25166 (N_25166,N_22930,N_23130);
xnor U25167 (N_25167,N_23940,N_23774);
nand U25168 (N_25168,N_23448,N_23458);
xnor U25169 (N_25169,N_22984,N_23420);
xnor U25170 (N_25170,N_23692,N_23926);
xor U25171 (N_25171,N_23711,N_23468);
or U25172 (N_25172,N_23727,N_23441);
or U25173 (N_25173,N_23843,N_23569);
nand U25174 (N_25174,N_23842,N_22811);
and U25175 (N_25175,N_23978,N_23948);
and U25176 (N_25176,N_22882,N_23825);
and U25177 (N_25177,N_23304,N_23114);
nor U25178 (N_25178,N_23849,N_23583);
and U25179 (N_25179,N_23583,N_23975);
nor U25180 (N_25180,N_23989,N_23550);
nor U25181 (N_25181,N_23132,N_23287);
nor U25182 (N_25182,N_23326,N_23869);
xor U25183 (N_25183,N_23952,N_23793);
or U25184 (N_25184,N_22814,N_22844);
and U25185 (N_25185,N_23258,N_23559);
or U25186 (N_25186,N_23842,N_23139);
xnor U25187 (N_25187,N_22900,N_23214);
xor U25188 (N_25188,N_23071,N_23001);
nand U25189 (N_25189,N_23988,N_23962);
xnor U25190 (N_25190,N_23317,N_23428);
nor U25191 (N_25191,N_23609,N_23919);
and U25192 (N_25192,N_23016,N_23814);
nor U25193 (N_25193,N_22931,N_22901);
nand U25194 (N_25194,N_23944,N_23946);
nor U25195 (N_25195,N_23143,N_23496);
nor U25196 (N_25196,N_23626,N_22987);
xnor U25197 (N_25197,N_22928,N_23345);
or U25198 (N_25198,N_23568,N_22960);
nand U25199 (N_25199,N_23322,N_23131);
or U25200 (N_25200,N_24953,N_24036);
nor U25201 (N_25201,N_24356,N_24924);
nand U25202 (N_25202,N_24778,N_25058);
and U25203 (N_25203,N_25196,N_25077);
nor U25204 (N_25204,N_24618,N_25093);
nand U25205 (N_25205,N_24718,N_25184);
or U25206 (N_25206,N_24745,N_24787);
xnor U25207 (N_25207,N_24721,N_25039);
nand U25208 (N_25208,N_25028,N_24774);
and U25209 (N_25209,N_24054,N_24420);
and U25210 (N_25210,N_24884,N_24030);
xnor U25211 (N_25211,N_24244,N_24888);
nand U25212 (N_25212,N_24915,N_24404);
and U25213 (N_25213,N_24962,N_25183);
and U25214 (N_25214,N_24109,N_24866);
xor U25215 (N_25215,N_24453,N_24832);
or U25216 (N_25216,N_24211,N_24765);
nand U25217 (N_25217,N_24084,N_24784);
xor U25218 (N_25218,N_24754,N_24677);
and U25219 (N_25219,N_24532,N_24679);
or U25220 (N_25220,N_24265,N_24753);
nor U25221 (N_25221,N_24583,N_24736);
nor U25222 (N_25222,N_24555,N_24249);
nand U25223 (N_25223,N_24992,N_24213);
nand U25224 (N_25224,N_24806,N_24327);
and U25225 (N_25225,N_24683,N_24966);
and U25226 (N_25226,N_24695,N_24986);
or U25227 (N_25227,N_24194,N_25123);
xnor U25228 (N_25228,N_24584,N_24430);
or U25229 (N_25229,N_24949,N_25131);
xor U25230 (N_25230,N_24398,N_24139);
and U25231 (N_25231,N_24990,N_24958);
or U25232 (N_25232,N_24926,N_24815);
or U25233 (N_25233,N_24569,N_24137);
nor U25234 (N_25234,N_24086,N_24066);
xnor U25235 (N_25235,N_24578,N_25163);
or U25236 (N_25236,N_24971,N_24002);
nor U25237 (N_25237,N_25153,N_25011);
and U25238 (N_25238,N_24014,N_24908);
or U25239 (N_25239,N_25113,N_24433);
xor U25240 (N_25240,N_24422,N_25103);
xor U25241 (N_25241,N_25197,N_24897);
nand U25242 (N_25242,N_24751,N_25137);
xor U25243 (N_25243,N_24538,N_24409);
nor U25244 (N_25244,N_24122,N_24709);
nand U25245 (N_25245,N_24456,N_24923);
nor U25246 (N_25246,N_24803,N_24837);
nand U25247 (N_25247,N_24065,N_24167);
and U25248 (N_25248,N_24808,N_24489);
nor U25249 (N_25249,N_24620,N_24196);
and U25250 (N_25250,N_24887,N_24401);
nand U25251 (N_25251,N_24667,N_24664);
xnor U25252 (N_25252,N_24617,N_24344);
or U25253 (N_25253,N_24389,N_24481);
and U25254 (N_25254,N_25005,N_24956);
xnor U25255 (N_25255,N_25016,N_24017);
nor U25256 (N_25256,N_24568,N_24841);
and U25257 (N_25257,N_24429,N_25146);
xor U25258 (N_25258,N_24171,N_24684);
nand U25259 (N_25259,N_24871,N_24214);
or U25260 (N_25260,N_24523,N_24308);
nand U25261 (N_25261,N_24177,N_24713);
nand U25262 (N_25262,N_24464,N_24282);
xnor U25263 (N_25263,N_24518,N_24854);
nor U25264 (N_25264,N_24499,N_24847);
and U25265 (N_25265,N_25185,N_24968);
nand U25266 (N_25266,N_24354,N_25106);
nand U25267 (N_25267,N_24925,N_24980);
nand U25268 (N_25268,N_24276,N_24314);
nand U25269 (N_25269,N_25177,N_24559);
nor U25270 (N_25270,N_24496,N_24197);
or U25271 (N_25271,N_24328,N_24991);
xor U25272 (N_25272,N_24904,N_25001);
or U25273 (N_25273,N_25045,N_24056);
xnor U25274 (N_25274,N_25190,N_24217);
nand U25275 (N_25275,N_24125,N_24190);
nand U25276 (N_25276,N_24243,N_25095);
xor U25277 (N_25277,N_24175,N_24416);
nor U25278 (N_25278,N_24468,N_24572);
nand U25279 (N_25279,N_24993,N_24642);
and U25280 (N_25280,N_24373,N_24647);
nand U25281 (N_25281,N_24027,N_25101);
and U25282 (N_25282,N_24406,N_24637);
xnor U25283 (N_25283,N_24042,N_24105);
nor U25284 (N_25284,N_24222,N_24154);
or U25285 (N_25285,N_24382,N_24530);
nand U25286 (N_25286,N_24948,N_24945);
xor U25287 (N_25287,N_24828,N_24432);
and U25288 (N_25288,N_25121,N_24255);
nor U25289 (N_25289,N_24431,N_24087);
or U25290 (N_25290,N_24223,N_24360);
and U25291 (N_25291,N_24207,N_25086);
xnor U25292 (N_25292,N_25186,N_24757);
or U25293 (N_25293,N_24394,N_24645);
nor U25294 (N_25294,N_24622,N_24500);
nor U25295 (N_25295,N_24567,N_24299);
nand U25296 (N_25296,N_24903,N_24598);
nand U25297 (N_25297,N_24610,N_24524);
or U25298 (N_25298,N_24155,N_24918);
nor U25299 (N_25299,N_24914,N_24296);
xnor U25300 (N_25300,N_24369,N_24070);
xor U25301 (N_25301,N_24452,N_24064);
or U25302 (N_25302,N_24073,N_24149);
xnor U25303 (N_25303,N_24690,N_24882);
nand U25304 (N_25304,N_24131,N_24018);
and U25305 (N_25305,N_25108,N_24839);
nand U25306 (N_25306,N_24459,N_24779);
xor U25307 (N_25307,N_25047,N_24534);
xor U25308 (N_25308,N_25164,N_25167);
nand U25309 (N_25309,N_24599,N_25090);
and U25310 (N_25310,N_24367,N_24232);
and U25311 (N_25311,N_24669,N_24902);
and U25312 (N_25312,N_24026,N_24362);
nand U25313 (N_25313,N_25053,N_24045);
nor U25314 (N_25314,N_24399,N_24205);
nor U25315 (N_25315,N_24863,N_24425);
and U25316 (N_25316,N_24655,N_24929);
or U25317 (N_25317,N_24979,N_24288);
and U25318 (N_25318,N_25174,N_24798);
xnor U25319 (N_25319,N_24741,N_24597);
or U25320 (N_25320,N_25176,N_25009);
and U25321 (N_25321,N_25088,N_24047);
xnor U25322 (N_25322,N_25084,N_24564);
nand U25323 (N_25323,N_24396,N_24016);
nand U25324 (N_25324,N_25055,N_25130);
or U25325 (N_25325,N_24785,N_24776);
or U25326 (N_25326,N_25160,N_24670);
nand U25327 (N_25327,N_24272,N_24032);
or U25328 (N_25328,N_24164,N_24686);
xor U25329 (N_25329,N_24883,N_24880);
or U25330 (N_25330,N_25120,N_24748);
nor U25331 (N_25331,N_24525,N_24558);
xnor U25332 (N_25332,N_24038,N_24147);
nor U25333 (N_25333,N_25169,N_24556);
xnor U25334 (N_25334,N_24768,N_24738);
xor U25335 (N_25335,N_24209,N_24068);
and U25336 (N_25336,N_24366,N_24769);
and U25337 (N_25337,N_24913,N_24941);
nor U25338 (N_25338,N_24117,N_24383);
and U25339 (N_25339,N_24478,N_24173);
xnor U25340 (N_25340,N_24917,N_25142);
nand U25341 (N_25341,N_24458,N_25073);
nor U25342 (N_25342,N_24157,N_24851);
nor U25343 (N_25343,N_24928,N_24102);
and U25344 (N_25344,N_24994,N_25014);
xnor U25345 (N_25345,N_24003,N_24615);
or U25346 (N_25346,N_24744,N_24881);
nand U25347 (N_25347,N_24384,N_24400);
xor U25348 (N_25348,N_24230,N_25178);
nand U25349 (N_25349,N_25119,N_24505);
nor U25350 (N_25350,N_24245,N_24722);
nor U25351 (N_25351,N_25135,N_24840);
nand U25352 (N_25352,N_24659,N_24535);
and U25353 (N_25353,N_24332,N_24020);
nor U25354 (N_25354,N_24822,N_25173);
or U25355 (N_25355,N_25063,N_24274);
nand U25356 (N_25356,N_24719,N_24187);
nand U25357 (N_25357,N_24504,N_24121);
and U25358 (N_25358,N_25117,N_24737);
nor U25359 (N_25359,N_24075,N_24942);
and U25360 (N_25360,N_24161,N_24920);
nand U25361 (N_25361,N_24674,N_24864);
and U25362 (N_25362,N_24685,N_24786);
xnor U25363 (N_25363,N_24596,N_25080);
xor U25364 (N_25364,N_24810,N_24707);
and U25365 (N_25365,N_24811,N_24100);
nor U25366 (N_25366,N_24077,N_24015);
or U25367 (N_25367,N_24860,N_24012);
nand U25368 (N_25368,N_24338,N_24735);
nor U25369 (N_25369,N_24997,N_24001);
and U25370 (N_25370,N_24633,N_25104);
and U25371 (N_25371,N_24310,N_24188);
or U25372 (N_25372,N_24104,N_24393);
or U25373 (N_25373,N_24701,N_24410);
nor U25374 (N_25374,N_24119,N_24443);
or U25375 (N_25375,N_24061,N_24444);
nand U25376 (N_25376,N_24069,N_24013);
and U25377 (N_25377,N_25036,N_24982);
and U25378 (N_25378,N_24340,N_24297);
or U25379 (N_25379,N_24879,N_24263);
nor U25380 (N_25380,N_24788,N_24589);
nand U25381 (N_25381,N_24570,N_24767);
and U25382 (N_25382,N_25064,N_25065);
or U25383 (N_25383,N_24044,N_24361);
xnor U25384 (N_25384,N_24442,N_24176);
nand U25385 (N_25385,N_24562,N_24083);
nor U25386 (N_25386,N_24629,N_24755);
nand U25387 (N_25387,N_24421,N_25157);
and U25388 (N_25388,N_25094,N_24698);
nand U25389 (N_25389,N_24235,N_24875);
nand U25390 (N_25390,N_24868,N_25021);
xor U25391 (N_25391,N_24358,N_24316);
nand U25392 (N_25392,N_24877,N_24483);
and U25393 (N_25393,N_25127,N_24529);
nand U25394 (N_25394,N_24264,N_24052);
or U25395 (N_25395,N_24665,N_25052);
or U25396 (N_25396,N_24726,N_24163);
or U25397 (N_25397,N_24388,N_24976);
nand U25398 (N_25398,N_24770,N_24543);
or U25399 (N_25399,N_24536,N_24099);
or U25400 (N_25400,N_24965,N_24635);
or U25401 (N_25401,N_24551,N_24470);
and U25402 (N_25402,N_24440,N_24640);
or U25403 (N_25403,N_24080,N_24309);
or U25404 (N_25404,N_24479,N_24174);
nand U25405 (N_25405,N_24715,N_24984);
or U25406 (N_25406,N_24566,N_25149);
and U25407 (N_25407,N_25099,N_24446);
and U25408 (N_25408,N_24493,N_25161);
and U25409 (N_25409,N_24236,N_25151);
xor U25410 (N_25410,N_25066,N_24258);
and U25411 (N_25411,N_25054,N_24096);
xor U25412 (N_25412,N_25031,N_24716);
xnor U25413 (N_25413,N_24780,N_24134);
nor U25414 (N_25414,N_24436,N_24818);
or U25415 (N_25415,N_24028,N_25141);
nor U25416 (N_25416,N_24675,N_24078);
xnor U25417 (N_25417,N_24368,N_24423);
or U25418 (N_25418,N_24856,N_24789);
xnor U25419 (N_25419,N_25118,N_25180);
and U25420 (N_25420,N_24239,N_24931);
nor U25421 (N_25421,N_25129,N_24341);
nand U25422 (N_25422,N_24725,N_24112);
xnor U25423 (N_25423,N_24040,N_25195);
nand U25424 (N_25424,N_24724,N_24700);
or U25425 (N_25425,N_24303,N_24079);
or U25426 (N_25426,N_24353,N_25139);
and U25427 (N_25427,N_25152,N_24812);
and U25428 (N_25428,N_24322,N_24513);
nand U25429 (N_25429,N_24873,N_24326);
nor U25430 (N_25430,N_24132,N_25044);
or U25431 (N_25431,N_24495,N_25092);
xnor U25432 (N_25432,N_25159,N_24606);
and U25433 (N_25433,N_25034,N_24870);
or U25434 (N_25434,N_25050,N_24821);
and U25435 (N_25435,N_24231,N_24202);
nand U25436 (N_25436,N_24266,N_24376);
or U25437 (N_25437,N_24295,N_24720);
nand U25438 (N_25438,N_24123,N_24932);
nand U25439 (N_25439,N_24571,N_24170);
nand U25440 (N_25440,N_24426,N_24350);
or U25441 (N_25441,N_24031,N_24413);
or U25442 (N_25442,N_24379,N_24336);
or U25443 (N_25443,N_24050,N_24792);
nor U25444 (N_25444,N_24581,N_24275);
xnor U25445 (N_25445,N_24397,N_24541);
and U25446 (N_25446,N_24939,N_25026);
nand U25447 (N_25447,N_24592,N_24427);
xnor U25448 (N_25448,N_24375,N_24981);
or U25449 (N_25449,N_24708,N_24944);
xor U25450 (N_25450,N_24643,N_24638);
nor U25451 (N_25451,N_25182,N_24899);
or U25452 (N_25452,N_24498,N_24447);
xnor U25453 (N_25453,N_25078,N_24702);
or U25454 (N_25454,N_24909,N_24503);
or U25455 (N_25455,N_24372,N_24219);
and U25456 (N_25456,N_25061,N_25075);
and U25457 (N_25457,N_24095,N_24989);
or U25458 (N_25458,N_24648,N_24819);
nor U25459 (N_25459,N_24657,N_24051);
nand U25460 (N_25460,N_24257,N_25147);
or U25461 (N_25461,N_24408,N_24260);
nand U25462 (N_25462,N_24355,N_24672);
xnor U25463 (N_25463,N_24251,N_24836);
nor U25464 (N_25464,N_24957,N_24461);
nand U25465 (N_25465,N_25126,N_24502);
xor U25466 (N_25466,N_25006,N_24717);
nor U25467 (N_25467,N_24311,N_25144);
and U25468 (N_25468,N_24723,N_24465);
xnor U25469 (N_25469,N_25111,N_24682);
or U25470 (N_25470,N_24290,N_25125);
nor U25471 (N_25471,N_24226,N_24557);
and U25472 (N_25472,N_24590,N_24653);
and U25473 (N_25473,N_24537,N_24273);
and U25474 (N_25474,N_24576,N_24681);
or U25475 (N_25475,N_24298,N_24604);
nor U25476 (N_25476,N_25033,N_24193);
or U25477 (N_25477,N_24621,N_24651);
or U25478 (N_25478,N_25171,N_24330);
xnor U25479 (N_25479,N_24654,N_24278);
and U25480 (N_25480,N_25070,N_24834);
or U25481 (N_25481,N_25166,N_24339);
nor U25482 (N_25482,N_25068,N_24762);
or U25483 (N_25483,N_24844,N_24062);
nor U25484 (N_25484,N_24545,N_25189);
or U25485 (N_25485,N_24363,N_24135);
and U25486 (N_25486,N_24693,N_25140);
xor U25487 (N_25487,N_24714,N_24547);
nand U25488 (N_25488,N_24024,N_24644);
nor U25489 (N_25489,N_24975,N_24697);
xor U25490 (N_25490,N_24224,N_24419);
and U25491 (N_25491,N_25194,N_24143);
or U25492 (N_25492,N_24973,N_24067);
nand U25493 (N_25493,N_25096,N_25091);
nor U25494 (N_25494,N_24855,N_24922);
and U25495 (N_25495,N_24593,N_25102);
and U25496 (N_25496,N_25037,N_24185);
or U25497 (N_25497,N_24761,N_24208);
xnor U25498 (N_25498,N_24858,N_24696);
xnor U25499 (N_25499,N_24000,N_24799);
nor U25500 (N_25500,N_25124,N_24094);
nand U25501 (N_25501,N_24838,N_24457);
xnor U25502 (N_25502,N_24110,N_24019);
xnor U25503 (N_25503,N_25133,N_24463);
nand U25504 (N_25504,N_24520,N_24800);
or U25505 (N_25505,N_24471,N_24935);
nand U25506 (N_25506,N_24029,N_24097);
and U25507 (N_25507,N_24248,N_24141);
and U25508 (N_25508,N_24403,N_24201);
nand U25509 (N_25509,N_25081,N_24861);
and U25510 (N_25510,N_24954,N_24750);
nand U25511 (N_25511,N_24092,N_24378);
xnor U25512 (N_25512,N_24473,N_24252);
nor U25513 (N_25513,N_24711,N_24699);
or U25514 (N_25514,N_25089,N_24631);
and U25515 (N_25515,N_25004,N_24692);
nand U25516 (N_25516,N_25145,N_24178);
xor U25517 (N_25517,N_24160,N_24955);
and U25518 (N_25518,N_24449,N_24111);
or U25519 (N_25519,N_24138,N_24668);
nor U25520 (N_25520,N_24307,N_24960);
xnor U25521 (N_25521,N_24867,N_24055);
nor U25522 (N_25522,N_24650,N_24514);
and U25523 (N_25523,N_24203,N_24445);
or U25524 (N_25524,N_24963,N_24414);
xor U25525 (N_25525,N_25082,N_24796);
and U25526 (N_25526,N_24005,N_24008);
or U25527 (N_25527,N_24417,N_24186);
nand U25528 (N_25528,N_24775,N_24085);
or U25529 (N_25529,N_24827,N_25132);
nor U25530 (N_25530,N_24907,N_24270);
nand U25531 (N_25531,N_24936,N_24120);
nand U25532 (N_25532,N_24034,N_24689);
and U25533 (N_25533,N_24329,N_24970);
nor U25534 (N_25534,N_24346,N_24752);
nand U25535 (N_25535,N_25041,N_24241);
nand U25536 (N_25536,N_24046,N_24424);
xnor U25537 (N_25537,N_24418,N_24352);
or U25538 (N_25538,N_24743,N_24512);
nor U25539 (N_25539,N_25154,N_24180);
or U25540 (N_25540,N_24706,N_24550);
nand U25541 (N_25541,N_24704,N_24023);
and U25542 (N_25542,N_24227,N_24335);
and U25543 (N_25543,N_24634,N_25158);
nor U25544 (N_25544,N_24485,N_24763);
or U25545 (N_25545,N_24626,N_24579);
nor U25546 (N_25546,N_25069,N_25029);
or U25547 (N_25547,N_24995,N_24183);
xnor U25548 (N_25548,N_24033,N_24961);
xor U25549 (N_25549,N_24233,N_24283);
xor U25550 (N_25550,N_24829,N_24850);
xnor U25551 (N_25551,N_24772,N_24324);
nand U25552 (N_25552,N_24561,N_24256);
nor U25553 (N_25553,N_24756,N_24168);
nor U25554 (N_25554,N_24043,N_25008);
xnor U25555 (N_25555,N_24742,N_24127);
nor U25556 (N_25556,N_24636,N_24126);
and U25557 (N_25557,N_24371,N_24294);
xnor U25558 (N_25558,N_24402,N_24891);
xor U25559 (N_25559,N_24377,N_25188);
nor U25560 (N_25560,N_24090,N_24660);
or U25561 (N_25561,N_24246,N_24025);
nand U25562 (N_25562,N_24688,N_24824);
nor U25563 (N_25563,N_24057,N_24846);
nor U25564 (N_25564,N_24730,N_24969);
and U25565 (N_25565,N_24781,N_24959);
and U25566 (N_25566,N_24106,N_24269);
or U25567 (N_25567,N_24254,N_24058);
xor U25568 (N_25568,N_24374,N_25143);
and U25569 (N_25569,N_25002,N_25192);
xnor U25570 (N_25570,N_24522,N_24115);
or U25571 (N_25571,N_24365,N_25175);
nor U25572 (N_25572,N_24951,N_24359);
or U25573 (N_25573,N_24200,N_24885);
and U25574 (N_25574,N_24395,N_24280);
nand U25575 (N_25575,N_24204,N_24927);
nand U25576 (N_25576,N_24943,N_24805);
nand U25577 (N_25577,N_24455,N_24337);
and U25578 (N_25578,N_25136,N_24490);
nand U25579 (N_25579,N_24041,N_24623);
nand U25580 (N_25580,N_24370,N_24542);
xnor U25581 (N_25581,N_24487,N_24676);
and U25582 (N_25582,N_24758,N_24206);
nand U25583 (N_25583,N_24588,N_24331);
or U25584 (N_25584,N_24347,N_25038);
or U25585 (N_25585,N_25022,N_24777);
or U25586 (N_25586,N_24428,N_24729);
and U25587 (N_25587,N_24516,N_24531);
nor U25588 (N_25588,N_24947,N_24220);
nor U25589 (N_25589,N_25027,N_24007);
xnor U25590 (N_25590,N_24292,N_24286);
or U25591 (N_25591,N_24950,N_24662);
and U25592 (N_25592,N_24921,N_24509);
nand U25593 (N_25593,N_24315,N_24862);
and U25594 (N_25594,N_24411,N_25040);
or U25595 (N_25595,N_24494,N_25168);
nand U25596 (N_25596,N_24783,N_25162);
xnor U25597 (N_25597,N_25187,N_24790);
nor U25598 (N_25598,N_24603,N_24519);
or U25599 (N_25599,N_24004,N_24601);
nor U25600 (N_25600,N_24237,N_24894);
and U25601 (N_25601,N_25042,N_24467);
nand U25602 (N_25602,N_24952,N_24749);
nand U25603 (N_25603,N_24825,N_24304);
nand U25604 (N_25604,N_25181,N_24876);
xor U25605 (N_25605,N_25051,N_24142);
nor U25606 (N_25606,N_25060,N_24482);
nor U25607 (N_25607,N_24439,N_24901);
and U25608 (N_25608,N_24527,N_24826);
nand U25609 (N_25609,N_24938,N_24540);
xnor U25610 (N_25610,N_24469,N_25115);
nand U25611 (N_25611,N_24351,N_24974);
xnor U25612 (N_25612,N_24037,N_24933);
and U25613 (N_25613,N_24852,N_24919);
nand U25614 (N_25614,N_24632,N_24462);
and U25615 (N_25615,N_24460,N_24228);
and U25616 (N_25616,N_24253,N_25198);
xor U25617 (N_25617,N_24987,N_24998);
nand U25618 (N_25618,N_24817,N_24694);
xnor U25619 (N_25619,N_24565,N_24434);
xnor U25620 (N_25620,N_24611,N_24148);
xnor U25621 (N_25621,N_24182,N_24114);
and U25622 (N_25622,N_24595,N_24144);
nor U25623 (N_25623,N_24247,N_25019);
or U25624 (N_25624,N_24271,N_24602);
or U25625 (N_25625,N_24088,N_24848);
xnor U25626 (N_25626,N_24898,N_24133);
and U25627 (N_25627,N_24472,N_24477);
nor U25628 (N_25628,N_24267,N_24548);
xor U25629 (N_25629,N_24607,N_24886);
xor U25630 (N_25630,N_25043,N_24608);
xor U25631 (N_25631,N_24978,N_25079);
nor U25632 (N_25632,N_24614,N_25085);
nor U25633 (N_25633,N_24150,N_24437);
nor U25634 (N_25634,N_25087,N_24747);
nor U25635 (N_25635,N_24585,N_24814);
nor U25636 (N_25636,N_24739,N_24343);
xor U25637 (N_25637,N_25172,N_24321);
and U25638 (N_25638,N_24391,N_24911);
xor U25639 (N_25639,N_24782,N_25128);
nand U25640 (N_25640,N_24546,N_24250);
and U25641 (N_25641,N_24656,N_24710);
or U25642 (N_25642,N_24063,N_25024);
nor U25643 (N_25643,N_24528,N_24625);
and U25644 (N_25644,N_24238,N_24628);
xnor U25645 (N_25645,N_24937,N_24641);
or U25646 (N_25646,N_24619,N_25110);
or U25647 (N_25647,N_25150,N_24830);
or U25648 (N_25648,N_25056,N_24159);
and U25649 (N_25649,N_24549,N_24405);
nand U25650 (N_25650,N_24195,N_24666);
nand U25651 (N_25651,N_24893,N_24996);
and U25652 (N_25652,N_25170,N_24151);
or U25653 (N_25653,N_24334,N_25097);
nand U25654 (N_25654,N_24731,N_24845);
nand U25655 (N_25655,N_24221,N_25148);
xor U25656 (N_25656,N_25062,N_24605);
nor U25657 (N_25657,N_24049,N_24021);
nand U25658 (N_25658,N_24039,N_24544);
or U25659 (N_25659,N_24554,N_24539);
nor U25660 (N_25660,N_24661,N_24771);
nand U25661 (N_25661,N_24890,N_24874);
and U25662 (N_25662,N_25012,N_25067);
nand U25663 (N_25663,N_24116,N_24809);
nand U25664 (N_25664,N_24794,N_24071);
and U25665 (N_25665,N_24128,N_25191);
or U25666 (N_25666,N_25048,N_24480);
nor U25667 (N_25667,N_24407,N_24306);
and U25668 (N_25668,N_24476,N_25199);
xnor U25669 (N_25669,N_24158,N_24577);
or U25670 (N_25670,N_24865,N_25018);
xnor U25671 (N_25671,N_24912,N_25017);
or U25672 (N_25672,N_24103,N_24515);
or U25673 (N_25673,N_24022,N_24760);
or U25674 (N_25674,N_24277,N_24076);
xnor U25675 (N_25675,N_24474,N_24198);
xor U25676 (N_25676,N_25112,N_25057);
nor U25677 (N_25677,N_25155,N_25035);
nand U25678 (N_25678,N_24318,N_24035);
nand U25679 (N_25679,N_24212,N_24074);
xnor U25680 (N_25680,N_25046,N_24441);
or U25681 (N_25681,N_24797,N_24181);
and U25682 (N_25682,N_24098,N_24082);
nand U25683 (N_25683,N_24009,N_24624);
nand U25684 (N_25684,N_24878,N_24613);
xor U25685 (N_25685,N_24988,N_24946);
and U25686 (N_25686,N_25083,N_24448);
or U25687 (N_25687,N_25049,N_24060);
or U25688 (N_25688,N_24189,N_25030);
xor U25689 (N_25689,N_24435,N_24563);
nand U25690 (N_25690,N_24746,N_24475);
nand U25691 (N_25691,N_24390,N_24072);
nand U25692 (N_25692,N_24801,N_24802);
nor U25693 (N_25693,N_24705,N_24108);
or U25694 (N_25694,N_24560,N_24011);
nand U25695 (N_25695,N_24733,N_24906);
nand U25696 (N_25696,N_24740,N_24342);
xnor U25697 (N_25697,N_24302,N_25165);
nor U25698 (N_25698,N_24594,N_24113);
and U25699 (N_25699,N_24807,N_24506);
nor U25700 (N_25700,N_24517,N_24118);
or U25701 (N_25701,N_24533,N_25007);
and U25702 (N_25702,N_24964,N_24392);
xnor U25703 (N_25703,N_24162,N_24703);
nor U25704 (N_25704,N_24240,N_25071);
nor U25705 (N_25705,N_24146,N_24609);
nor U25706 (N_25706,N_25072,N_24728);
and U25707 (N_25707,N_24415,N_25107);
nor U25708 (N_25708,N_24387,N_24831);
nor U25709 (N_25709,N_24289,N_24300);
nor U25710 (N_25710,N_24454,N_24268);
nand U25711 (N_25711,N_24313,N_24930);
and U25712 (N_25712,N_24859,N_24591);
or U25713 (N_25713,N_24156,N_24804);
nand U25714 (N_25714,N_24165,N_25138);
xnor U25715 (N_25715,N_24508,N_24301);
xor U25716 (N_25716,N_24140,N_24130);
nor U25717 (N_25717,N_24348,N_24816);
nor U25718 (N_25718,N_25105,N_24843);
and U25719 (N_25719,N_24323,N_24934);
xor U25720 (N_25720,N_24582,N_24259);
nand U25721 (N_25721,N_24172,N_24081);
nor U25722 (N_25722,N_24600,N_25156);
nand U25723 (N_25723,N_24521,N_24053);
nand U25724 (N_25724,N_24892,N_24191);
and U25725 (N_25725,N_24325,N_25109);
nand U25726 (N_25726,N_25179,N_24486);
nor U25727 (N_25727,N_24192,N_25025);
nor U25728 (N_25728,N_24630,N_24872);
nor U25729 (N_25729,N_24291,N_24317);
xnor U25730 (N_25730,N_24553,N_25003);
and U25731 (N_25731,N_24199,N_24385);
nor U25732 (N_25732,N_24438,N_24727);
xor U25733 (N_25733,N_24823,N_24734);
nand U25734 (N_25734,N_24833,N_25013);
nand U25735 (N_25735,N_24869,N_24484);
nor U25736 (N_25736,N_24820,N_25100);
xnor U25737 (N_25737,N_24451,N_25098);
or U25738 (N_25738,N_24732,N_24510);
nand U25739 (N_25739,N_24466,N_24639);
and U25740 (N_25740,N_24279,N_25000);
nand U25741 (N_25741,N_24225,N_24712);
and U25742 (N_25742,N_24059,N_24215);
or U25743 (N_25743,N_24900,N_24284);
and U25744 (N_25744,N_24916,N_24835);
or U25745 (N_25745,N_24587,N_24091);
xnor U25746 (N_25746,N_24983,N_24229);
and U25747 (N_25747,N_24575,N_24905);
xor U25748 (N_25748,N_24497,N_24492);
and U25749 (N_25749,N_25116,N_24349);
xor U25750 (N_25750,N_24759,N_24857);
nand U25751 (N_25751,N_25193,N_24216);
or U25752 (N_25752,N_24166,N_24242);
nor U25753 (N_25753,N_24849,N_24680);
xnor U25754 (N_25754,N_24573,N_24691);
or U25755 (N_25755,N_24658,N_24574);
and U25756 (N_25756,N_24580,N_24977);
or U25757 (N_25757,N_24319,N_24552);
nor U25758 (N_25758,N_24006,N_25059);
nor U25759 (N_25759,N_24766,N_25023);
nand U25760 (N_25760,N_24333,N_25020);
or U25761 (N_25761,N_24381,N_24262);
or U25762 (N_25762,N_24320,N_24152);
nand U25763 (N_25763,N_24364,N_24287);
or U25764 (N_25764,N_24010,N_24764);
nor U25765 (N_25765,N_24491,N_24795);
nor U25766 (N_25766,N_24293,N_25015);
xnor U25767 (N_25767,N_24842,N_24129);
and U25768 (N_25768,N_24791,N_24281);
nand U25769 (N_25769,N_24889,N_24813);
or U25770 (N_25770,N_24357,N_24627);
nand U25771 (N_25771,N_24910,N_25074);
nand U25772 (N_25772,N_24678,N_24136);
and U25773 (N_25773,N_24184,N_24089);
xnor U25774 (N_25774,N_24048,N_24511);
and U25775 (N_25775,N_24412,N_24652);
nand U25776 (N_25776,N_24616,N_24124);
xor U25777 (N_25777,N_25134,N_24649);
or U25778 (N_25778,N_24646,N_24101);
xor U25779 (N_25779,N_24793,N_24218);
or U25780 (N_25780,N_24093,N_24488);
xor U25781 (N_25781,N_24169,N_24285);
and U25782 (N_25782,N_24773,N_25032);
nand U25783 (N_25783,N_25114,N_25122);
and U25784 (N_25784,N_24305,N_24380);
and U25785 (N_25785,N_24261,N_24107);
xnor U25786 (N_25786,N_24501,N_24179);
xor U25787 (N_25787,N_24450,N_24145);
or U25788 (N_25788,N_24687,N_24940);
nand U25789 (N_25789,N_24345,N_24586);
xor U25790 (N_25790,N_24999,N_24895);
or U25791 (N_25791,N_24673,N_24967);
xnor U25792 (N_25792,N_24507,N_24985);
nor U25793 (N_25793,N_24312,N_25076);
nor U25794 (N_25794,N_24853,N_24671);
xor U25795 (N_25795,N_24386,N_24663);
or U25796 (N_25796,N_24153,N_24526);
xnor U25797 (N_25797,N_24896,N_24972);
nand U25798 (N_25798,N_24234,N_25010);
nand U25799 (N_25799,N_24612,N_24210);
or U25800 (N_25800,N_24375,N_24182);
and U25801 (N_25801,N_24557,N_24566);
nand U25802 (N_25802,N_24420,N_24524);
xnor U25803 (N_25803,N_24780,N_25037);
or U25804 (N_25804,N_24577,N_24610);
and U25805 (N_25805,N_24995,N_24273);
and U25806 (N_25806,N_24596,N_24489);
nor U25807 (N_25807,N_24567,N_25014);
and U25808 (N_25808,N_25185,N_24740);
nand U25809 (N_25809,N_24737,N_24031);
xor U25810 (N_25810,N_24147,N_24142);
and U25811 (N_25811,N_24834,N_24863);
nand U25812 (N_25812,N_24281,N_24075);
nor U25813 (N_25813,N_24789,N_24675);
xor U25814 (N_25814,N_24974,N_25086);
or U25815 (N_25815,N_24709,N_24657);
nand U25816 (N_25816,N_24845,N_24070);
and U25817 (N_25817,N_24085,N_24398);
nand U25818 (N_25818,N_24161,N_24026);
and U25819 (N_25819,N_24083,N_24760);
and U25820 (N_25820,N_24433,N_24387);
or U25821 (N_25821,N_24098,N_24995);
or U25822 (N_25822,N_25134,N_24456);
xnor U25823 (N_25823,N_24440,N_25092);
nor U25824 (N_25824,N_24878,N_24473);
or U25825 (N_25825,N_24425,N_24169);
or U25826 (N_25826,N_24239,N_24460);
nand U25827 (N_25827,N_25167,N_24789);
or U25828 (N_25828,N_24860,N_24299);
xnor U25829 (N_25829,N_25039,N_24823);
and U25830 (N_25830,N_24584,N_25068);
nor U25831 (N_25831,N_24359,N_24639);
and U25832 (N_25832,N_24307,N_24105);
and U25833 (N_25833,N_24775,N_24572);
and U25834 (N_25834,N_24839,N_24402);
and U25835 (N_25835,N_25003,N_24836);
or U25836 (N_25836,N_25111,N_24548);
xnor U25837 (N_25837,N_25063,N_24930);
or U25838 (N_25838,N_24917,N_24629);
or U25839 (N_25839,N_24412,N_25173);
or U25840 (N_25840,N_24150,N_25180);
nor U25841 (N_25841,N_24738,N_24147);
xnor U25842 (N_25842,N_24110,N_24391);
xor U25843 (N_25843,N_24841,N_24393);
and U25844 (N_25844,N_24906,N_24415);
and U25845 (N_25845,N_25136,N_24220);
nor U25846 (N_25846,N_24099,N_25142);
nand U25847 (N_25847,N_24355,N_24422);
nand U25848 (N_25848,N_24734,N_24169);
xnor U25849 (N_25849,N_25113,N_24598);
and U25850 (N_25850,N_25141,N_24924);
nor U25851 (N_25851,N_24108,N_24429);
and U25852 (N_25852,N_24490,N_24421);
or U25853 (N_25853,N_24767,N_24041);
and U25854 (N_25854,N_24539,N_24079);
or U25855 (N_25855,N_24368,N_24085);
nor U25856 (N_25856,N_24629,N_24226);
and U25857 (N_25857,N_24450,N_25133);
nand U25858 (N_25858,N_24581,N_24389);
and U25859 (N_25859,N_24213,N_24600);
nand U25860 (N_25860,N_24614,N_25195);
nor U25861 (N_25861,N_24346,N_24341);
xor U25862 (N_25862,N_24503,N_24517);
or U25863 (N_25863,N_24804,N_24964);
or U25864 (N_25864,N_25128,N_24394);
or U25865 (N_25865,N_24130,N_24604);
nand U25866 (N_25866,N_24715,N_24607);
xnor U25867 (N_25867,N_24359,N_24848);
xnor U25868 (N_25868,N_25161,N_24121);
and U25869 (N_25869,N_24796,N_24486);
xor U25870 (N_25870,N_24503,N_24031);
nor U25871 (N_25871,N_25007,N_24355);
or U25872 (N_25872,N_24378,N_24572);
and U25873 (N_25873,N_25076,N_24178);
nor U25874 (N_25874,N_24395,N_24194);
xor U25875 (N_25875,N_24393,N_25011);
and U25876 (N_25876,N_24504,N_24793);
xor U25877 (N_25877,N_24395,N_24678);
nand U25878 (N_25878,N_24134,N_24682);
and U25879 (N_25879,N_24851,N_24440);
and U25880 (N_25880,N_24184,N_24865);
nand U25881 (N_25881,N_24568,N_24907);
nor U25882 (N_25882,N_24620,N_24023);
nor U25883 (N_25883,N_24949,N_24849);
nand U25884 (N_25884,N_24226,N_24476);
and U25885 (N_25885,N_24277,N_24572);
nand U25886 (N_25886,N_24979,N_24181);
nand U25887 (N_25887,N_24437,N_24903);
xor U25888 (N_25888,N_25075,N_25149);
and U25889 (N_25889,N_24691,N_24185);
xnor U25890 (N_25890,N_24565,N_25148);
xnor U25891 (N_25891,N_24807,N_25108);
xor U25892 (N_25892,N_25019,N_24287);
nor U25893 (N_25893,N_24931,N_24168);
nor U25894 (N_25894,N_24197,N_24474);
nand U25895 (N_25895,N_24788,N_24383);
and U25896 (N_25896,N_24801,N_24252);
xor U25897 (N_25897,N_24658,N_24481);
nor U25898 (N_25898,N_25107,N_24151);
nor U25899 (N_25899,N_24025,N_25167);
nand U25900 (N_25900,N_24250,N_24698);
xnor U25901 (N_25901,N_24696,N_24320);
nand U25902 (N_25902,N_24869,N_24560);
nor U25903 (N_25903,N_24736,N_24158);
xor U25904 (N_25904,N_24577,N_24013);
or U25905 (N_25905,N_24307,N_24500);
nor U25906 (N_25906,N_24123,N_24526);
nor U25907 (N_25907,N_24735,N_24136);
nand U25908 (N_25908,N_24104,N_24064);
nor U25909 (N_25909,N_24727,N_25068);
nand U25910 (N_25910,N_24932,N_24722);
and U25911 (N_25911,N_24846,N_24354);
and U25912 (N_25912,N_24888,N_25153);
nand U25913 (N_25913,N_24506,N_24194);
or U25914 (N_25914,N_24589,N_24172);
nand U25915 (N_25915,N_24799,N_25093);
nor U25916 (N_25916,N_24254,N_24962);
or U25917 (N_25917,N_25048,N_24165);
nand U25918 (N_25918,N_24970,N_24537);
nand U25919 (N_25919,N_24611,N_24733);
and U25920 (N_25920,N_24795,N_24092);
xnor U25921 (N_25921,N_24782,N_24833);
or U25922 (N_25922,N_24546,N_24299);
nand U25923 (N_25923,N_24413,N_24992);
and U25924 (N_25924,N_24599,N_24301);
xnor U25925 (N_25925,N_24689,N_25188);
or U25926 (N_25926,N_24311,N_24183);
and U25927 (N_25927,N_25114,N_24281);
or U25928 (N_25928,N_25021,N_24377);
nor U25929 (N_25929,N_24101,N_24557);
and U25930 (N_25930,N_24631,N_24811);
and U25931 (N_25931,N_24277,N_25054);
and U25932 (N_25932,N_24168,N_24744);
or U25933 (N_25933,N_24942,N_24599);
and U25934 (N_25934,N_24865,N_25154);
or U25935 (N_25935,N_25126,N_24353);
nor U25936 (N_25936,N_24091,N_25122);
nor U25937 (N_25937,N_24101,N_24539);
xnor U25938 (N_25938,N_24300,N_25063);
or U25939 (N_25939,N_24125,N_25003);
xor U25940 (N_25940,N_24608,N_24964);
nor U25941 (N_25941,N_25037,N_25177);
nand U25942 (N_25942,N_24851,N_24312);
nand U25943 (N_25943,N_24582,N_24894);
and U25944 (N_25944,N_24144,N_24773);
nand U25945 (N_25945,N_24601,N_24640);
nor U25946 (N_25946,N_24256,N_25128);
nand U25947 (N_25947,N_24808,N_24522);
nor U25948 (N_25948,N_24546,N_24439);
nand U25949 (N_25949,N_24113,N_24439);
xnor U25950 (N_25950,N_24732,N_25069);
or U25951 (N_25951,N_24366,N_24550);
or U25952 (N_25952,N_24330,N_24310);
xor U25953 (N_25953,N_24629,N_24575);
or U25954 (N_25954,N_25027,N_24831);
or U25955 (N_25955,N_24022,N_24290);
nor U25956 (N_25956,N_24437,N_24941);
nand U25957 (N_25957,N_24480,N_24947);
xnor U25958 (N_25958,N_24796,N_24771);
nand U25959 (N_25959,N_24694,N_24220);
or U25960 (N_25960,N_24672,N_24233);
and U25961 (N_25961,N_25086,N_24235);
nor U25962 (N_25962,N_24833,N_24196);
nand U25963 (N_25963,N_24548,N_25003);
or U25964 (N_25964,N_24196,N_24430);
or U25965 (N_25965,N_25147,N_24750);
xnor U25966 (N_25966,N_24440,N_24469);
xnor U25967 (N_25967,N_25001,N_24434);
nand U25968 (N_25968,N_24185,N_24957);
and U25969 (N_25969,N_24397,N_24499);
or U25970 (N_25970,N_24877,N_24858);
nor U25971 (N_25971,N_24269,N_24313);
or U25972 (N_25972,N_25057,N_24059);
xnor U25973 (N_25973,N_24206,N_24619);
and U25974 (N_25974,N_24531,N_25024);
or U25975 (N_25975,N_24262,N_24417);
xor U25976 (N_25976,N_24781,N_24878);
or U25977 (N_25977,N_25108,N_24452);
nand U25978 (N_25978,N_24602,N_25174);
xnor U25979 (N_25979,N_24878,N_24138);
nand U25980 (N_25980,N_24409,N_24145);
and U25981 (N_25981,N_24255,N_24606);
nor U25982 (N_25982,N_24144,N_25039);
and U25983 (N_25983,N_24958,N_24105);
nand U25984 (N_25984,N_24871,N_24579);
and U25985 (N_25985,N_24253,N_24779);
xor U25986 (N_25986,N_24015,N_24528);
and U25987 (N_25987,N_24756,N_24698);
nand U25988 (N_25988,N_24949,N_24475);
or U25989 (N_25989,N_25021,N_24333);
or U25990 (N_25990,N_24255,N_24593);
nand U25991 (N_25991,N_24015,N_24371);
and U25992 (N_25992,N_25116,N_24252);
and U25993 (N_25993,N_24576,N_24447);
and U25994 (N_25994,N_25055,N_24087);
or U25995 (N_25995,N_24145,N_24621);
or U25996 (N_25996,N_25108,N_24444);
nor U25997 (N_25997,N_24331,N_24093);
nor U25998 (N_25998,N_24735,N_25056);
xor U25999 (N_25999,N_24700,N_25055);
xnor U26000 (N_26000,N_24121,N_24902);
or U26001 (N_26001,N_24968,N_24935);
or U26002 (N_26002,N_24136,N_25029);
or U26003 (N_26003,N_24657,N_24098);
nor U26004 (N_26004,N_25002,N_24417);
or U26005 (N_26005,N_24405,N_24257);
nand U26006 (N_26006,N_24063,N_24951);
or U26007 (N_26007,N_24055,N_24394);
and U26008 (N_26008,N_24970,N_25049);
nor U26009 (N_26009,N_24719,N_24745);
xor U26010 (N_26010,N_24447,N_24816);
xnor U26011 (N_26011,N_25165,N_24877);
xor U26012 (N_26012,N_24502,N_25038);
nand U26013 (N_26013,N_24363,N_25062);
and U26014 (N_26014,N_24091,N_24002);
or U26015 (N_26015,N_24027,N_24484);
xor U26016 (N_26016,N_24803,N_24802);
nor U26017 (N_26017,N_24173,N_24038);
nor U26018 (N_26018,N_24168,N_24739);
and U26019 (N_26019,N_24964,N_24594);
nor U26020 (N_26020,N_24570,N_24172);
or U26021 (N_26021,N_24854,N_25188);
nand U26022 (N_26022,N_24348,N_24265);
nor U26023 (N_26023,N_24008,N_24149);
or U26024 (N_26024,N_24734,N_25034);
and U26025 (N_26025,N_25075,N_25017);
nand U26026 (N_26026,N_24792,N_24292);
nor U26027 (N_26027,N_24933,N_24848);
or U26028 (N_26028,N_24544,N_24755);
and U26029 (N_26029,N_24258,N_24888);
xnor U26030 (N_26030,N_24889,N_24749);
and U26031 (N_26031,N_24104,N_24311);
xor U26032 (N_26032,N_24703,N_24898);
xor U26033 (N_26033,N_24220,N_24979);
or U26034 (N_26034,N_24489,N_24297);
nand U26035 (N_26035,N_24196,N_24167);
and U26036 (N_26036,N_24382,N_24166);
and U26037 (N_26037,N_24227,N_24482);
or U26038 (N_26038,N_24384,N_24623);
and U26039 (N_26039,N_24924,N_24719);
xor U26040 (N_26040,N_24939,N_24890);
nor U26041 (N_26041,N_24062,N_24631);
and U26042 (N_26042,N_24211,N_24240);
or U26043 (N_26043,N_24258,N_24158);
or U26044 (N_26044,N_24524,N_25015);
xor U26045 (N_26045,N_24436,N_24055);
or U26046 (N_26046,N_24398,N_24675);
xor U26047 (N_26047,N_24594,N_25019);
or U26048 (N_26048,N_24688,N_24509);
nor U26049 (N_26049,N_24652,N_25054);
and U26050 (N_26050,N_25180,N_25080);
nor U26051 (N_26051,N_24932,N_24957);
or U26052 (N_26052,N_24823,N_25038);
or U26053 (N_26053,N_25140,N_24015);
nand U26054 (N_26054,N_24689,N_25003);
or U26055 (N_26055,N_24328,N_24327);
nor U26056 (N_26056,N_24286,N_24739);
nand U26057 (N_26057,N_24864,N_24354);
xnor U26058 (N_26058,N_24719,N_24306);
or U26059 (N_26059,N_24349,N_24023);
nand U26060 (N_26060,N_24380,N_24617);
or U26061 (N_26061,N_25102,N_24658);
nand U26062 (N_26062,N_25187,N_24600);
xor U26063 (N_26063,N_24432,N_24377);
and U26064 (N_26064,N_24304,N_24051);
nor U26065 (N_26065,N_24679,N_24208);
or U26066 (N_26066,N_24690,N_24027);
nand U26067 (N_26067,N_24827,N_24491);
and U26068 (N_26068,N_24223,N_24520);
and U26069 (N_26069,N_24558,N_24587);
nor U26070 (N_26070,N_24313,N_24426);
nand U26071 (N_26071,N_24993,N_24787);
or U26072 (N_26072,N_24161,N_24429);
or U26073 (N_26073,N_25013,N_24457);
and U26074 (N_26074,N_24159,N_25072);
nor U26075 (N_26075,N_25071,N_24293);
and U26076 (N_26076,N_24587,N_24782);
or U26077 (N_26077,N_24769,N_24279);
nor U26078 (N_26078,N_25040,N_24276);
nor U26079 (N_26079,N_24895,N_24479);
nor U26080 (N_26080,N_24328,N_24456);
xnor U26081 (N_26081,N_24901,N_24980);
xnor U26082 (N_26082,N_25072,N_24241);
or U26083 (N_26083,N_25096,N_24486);
and U26084 (N_26084,N_25089,N_24870);
and U26085 (N_26085,N_24698,N_24700);
xnor U26086 (N_26086,N_24684,N_24155);
xnor U26087 (N_26087,N_24386,N_24894);
and U26088 (N_26088,N_24591,N_25094);
xnor U26089 (N_26089,N_24566,N_24673);
and U26090 (N_26090,N_24980,N_24265);
nor U26091 (N_26091,N_24116,N_24926);
and U26092 (N_26092,N_24213,N_24089);
xnor U26093 (N_26093,N_24526,N_24088);
nor U26094 (N_26094,N_24173,N_24598);
and U26095 (N_26095,N_24098,N_24237);
nand U26096 (N_26096,N_25056,N_24229);
or U26097 (N_26097,N_24717,N_24527);
nand U26098 (N_26098,N_24556,N_24896);
and U26099 (N_26099,N_25099,N_24371);
xnor U26100 (N_26100,N_24593,N_24757);
and U26101 (N_26101,N_24532,N_24283);
and U26102 (N_26102,N_24272,N_24792);
and U26103 (N_26103,N_24495,N_24662);
xor U26104 (N_26104,N_24376,N_24898);
or U26105 (N_26105,N_24941,N_24950);
xor U26106 (N_26106,N_25163,N_24673);
xor U26107 (N_26107,N_24037,N_24356);
nand U26108 (N_26108,N_24669,N_24492);
nand U26109 (N_26109,N_25197,N_24653);
xnor U26110 (N_26110,N_25146,N_24629);
and U26111 (N_26111,N_24281,N_24599);
nand U26112 (N_26112,N_24901,N_24876);
and U26113 (N_26113,N_24321,N_25068);
nor U26114 (N_26114,N_24908,N_25024);
and U26115 (N_26115,N_25135,N_24784);
and U26116 (N_26116,N_24093,N_24413);
and U26117 (N_26117,N_24930,N_24211);
and U26118 (N_26118,N_24918,N_24049);
or U26119 (N_26119,N_24609,N_25088);
nand U26120 (N_26120,N_25042,N_24657);
xor U26121 (N_26121,N_24913,N_24030);
or U26122 (N_26122,N_24094,N_24818);
xor U26123 (N_26123,N_24821,N_24052);
nand U26124 (N_26124,N_24148,N_24706);
or U26125 (N_26125,N_24169,N_24378);
xor U26126 (N_26126,N_24614,N_24450);
or U26127 (N_26127,N_24249,N_24237);
nor U26128 (N_26128,N_24239,N_24191);
xor U26129 (N_26129,N_24286,N_24326);
or U26130 (N_26130,N_25177,N_24303);
nand U26131 (N_26131,N_24106,N_24562);
xor U26132 (N_26132,N_25155,N_24695);
and U26133 (N_26133,N_24270,N_25034);
nor U26134 (N_26134,N_24996,N_24981);
nand U26135 (N_26135,N_24395,N_24403);
or U26136 (N_26136,N_24500,N_24011);
or U26137 (N_26137,N_24952,N_24960);
nor U26138 (N_26138,N_24558,N_24806);
xnor U26139 (N_26139,N_24218,N_24102);
and U26140 (N_26140,N_25023,N_24774);
or U26141 (N_26141,N_24220,N_25131);
xnor U26142 (N_26142,N_24116,N_24800);
and U26143 (N_26143,N_24499,N_24494);
xor U26144 (N_26144,N_24428,N_25186);
and U26145 (N_26145,N_25191,N_24849);
nor U26146 (N_26146,N_24854,N_25013);
nand U26147 (N_26147,N_24793,N_24749);
or U26148 (N_26148,N_24434,N_25122);
nor U26149 (N_26149,N_24201,N_24775);
xnor U26150 (N_26150,N_24206,N_25144);
nand U26151 (N_26151,N_24062,N_24987);
and U26152 (N_26152,N_24496,N_24662);
xnor U26153 (N_26153,N_24693,N_24692);
xor U26154 (N_26154,N_24807,N_24929);
and U26155 (N_26155,N_24068,N_24945);
or U26156 (N_26156,N_24666,N_25168);
xnor U26157 (N_26157,N_24719,N_24143);
xnor U26158 (N_26158,N_24606,N_24074);
and U26159 (N_26159,N_24541,N_25053);
xnor U26160 (N_26160,N_25138,N_25182);
xnor U26161 (N_26161,N_24607,N_24410);
and U26162 (N_26162,N_24198,N_25109);
or U26163 (N_26163,N_24237,N_24325);
nor U26164 (N_26164,N_24210,N_24670);
and U26165 (N_26165,N_24492,N_25144);
and U26166 (N_26166,N_25018,N_24887);
nand U26167 (N_26167,N_24926,N_24447);
or U26168 (N_26168,N_25165,N_24770);
xnor U26169 (N_26169,N_25067,N_24806);
nor U26170 (N_26170,N_24025,N_24124);
xor U26171 (N_26171,N_24276,N_24691);
or U26172 (N_26172,N_24475,N_24049);
nand U26173 (N_26173,N_24492,N_24958);
or U26174 (N_26174,N_24261,N_24063);
nand U26175 (N_26175,N_25127,N_24022);
and U26176 (N_26176,N_24349,N_24968);
xor U26177 (N_26177,N_25149,N_24773);
and U26178 (N_26178,N_24909,N_24070);
nand U26179 (N_26179,N_24098,N_24919);
nand U26180 (N_26180,N_24663,N_24774);
xor U26181 (N_26181,N_24092,N_24100);
nand U26182 (N_26182,N_24040,N_24766);
nor U26183 (N_26183,N_24930,N_24022);
and U26184 (N_26184,N_24324,N_24753);
and U26185 (N_26185,N_24167,N_24056);
xor U26186 (N_26186,N_25031,N_25082);
and U26187 (N_26187,N_24255,N_24028);
nand U26188 (N_26188,N_24501,N_25121);
nor U26189 (N_26189,N_24305,N_24721);
or U26190 (N_26190,N_25075,N_25195);
or U26191 (N_26191,N_24324,N_24623);
xnor U26192 (N_26192,N_24127,N_24030);
nor U26193 (N_26193,N_24492,N_24836);
and U26194 (N_26194,N_24543,N_24117);
xnor U26195 (N_26195,N_24409,N_24963);
or U26196 (N_26196,N_24127,N_24658);
and U26197 (N_26197,N_24476,N_24139);
and U26198 (N_26198,N_24278,N_24892);
and U26199 (N_26199,N_24373,N_24724);
xnor U26200 (N_26200,N_24701,N_24497);
nor U26201 (N_26201,N_24971,N_24486);
nor U26202 (N_26202,N_24838,N_24047);
nand U26203 (N_26203,N_24306,N_24469);
nand U26204 (N_26204,N_25067,N_24208);
xor U26205 (N_26205,N_24728,N_25071);
and U26206 (N_26206,N_25060,N_25070);
xnor U26207 (N_26207,N_24143,N_24104);
or U26208 (N_26208,N_24905,N_24101);
nand U26209 (N_26209,N_24476,N_24533);
nand U26210 (N_26210,N_24093,N_24453);
or U26211 (N_26211,N_24047,N_24519);
and U26212 (N_26212,N_24797,N_24513);
nor U26213 (N_26213,N_24549,N_25014);
or U26214 (N_26214,N_24933,N_24025);
nand U26215 (N_26215,N_24115,N_24271);
nand U26216 (N_26216,N_24787,N_24180);
nor U26217 (N_26217,N_24533,N_25198);
xnor U26218 (N_26218,N_24070,N_24584);
nor U26219 (N_26219,N_24958,N_24053);
and U26220 (N_26220,N_24291,N_24916);
nor U26221 (N_26221,N_24114,N_25080);
or U26222 (N_26222,N_24307,N_24808);
xor U26223 (N_26223,N_24136,N_24296);
or U26224 (N_26224,N_24679,N_24804);
nand U26225 (N_26225,N_25088,N_25073);
or U26226 (N_26226,N_24852,N_24496);
nor U26227 (N_26227,N_24314,N_24882);
or U26228 (N_26228,N_24596,N_24061);
and U26229 (N_26229,N_24607,N_25117);
nand U26230 (N_26230,N_25111,N_24071);
and U26231 (N_26231,N_24042,N_24184);
and U26232 (N_26232,N_24004,N_24783);
nor U26233 (N_26233,N_25198,N_24427);
nand U26234 (N_26234,N_24076,N_24620);
and U26235 (N_26235,N_24756,N_24315);
or U26236 (N_26236,N_24852,N_24179);
nor U26237 (N_26237,N_25078,N_24819);
or U26238 (N_26238,N_24916,N_24037);
and U26239 (N_26239,N_24245,N_25080);
nand U26240 (N_26240,N_24156,N_25093);
xnor U26241 (N_26241,N_24363,N_24153);
and U26242 (N_26242,N_24520,N_24047);
or U26243 (N_26243,N_24077,N_25028);
and U26244 (N_26244,N_24694,N_24590);
and U26245 (N_26245,N_24760,N_24881);
or U26246 (N_26246,N_24427,N_24076);
nand U26247 (N_26247,N_24946,N_24836);
nand U26248 (N_26248,N_24811,N_24360);
and U26249 (N_26249,N_24895,N_24697);
nand U26250 (N_26250,N_24988,N_24199);
or U26251 (N_26251,N_24944,N_24122);
xnor U26252 (N_26252,N_24983,N_24697);
nand U26253 (N_26253,N_24481,N_24903);
nand U26254 (N_26254,N_24330,N_25009);
nor U26255 (N_26255,N_24564,N_24301);
xor U26256 (N_26256,N_25051,N_24904);
xor U26257 (N_26257,N_25141,N_24699);
and U26258 (N_26258,N_24824,N_24949);
or U26259 (N_26259,N_24268,N_24717);
nor U26260 (N_26260,N_24157,N_24370);
xor U26261 (N_26261,N_24133,N_24296);
and U26262 (N_26262,N_24908,N_25091);
nand U26263 (N_26263,N_24076,N_24704);
nand U26264 (N_26264,N_25111,N_24488);
nor U26265 (N_26265,N_24683,N_24815);
and U26266 (N_26266,N_24723,N_25106);
xnor U26267 (N_26267,N_25196,N_24021);
or U26268 (N_26268,N_24077,N_24160);
nand U26269 (N_26269,N_24708,N_24328);
xor U26270 (N_26270,N_25151,N_24686);
and U26271 (N_26271,N_24190,N_25162);
and U26272 (N_26272,N_24162,N_24287);
nor U26273 (N_26273,N_24444,N_24603);
or U26274 (N_26274,N_24163,N_24294);
or U26275 (N_26275,N_24690,N_24917);
nand U26276 (N_26276,N_25137,N_24822);
xnor U26277 (N_26277,N_24075,N_24099);
nand U26278 (N_26278,N_25141,N_24840);
nor U26279 (N_26279,N_24475,N_24015);
or U26280 (N_26280,N_25167,N_24539);
nor U26281 (N_26281,N_24213,N_24490);
xor U26282 (N_26282,N_24185,N_24746);
and U26283 (N_26283,N_25114,N_24826);
and U26284 (N_26284,N_24135,N_25120);
and U26285 (N_26285,N_24953,N_25171);
and U26286 (N_26286,N_24990,N_24692);
nor U26287 (N_26287,N_24055,N_25143);
or U26288 (N_26288,N_24542,N_24456);
nand U26289 (N_26289,N_24746,N_24725);
and U26290 (N_26290,N_25153,N_24199);
xnor U26291 (N_26291,N_24979,N_24611);
and U26292 (N_26292,N_24234,N_24538);
xnor U26293 (N_26293,N_24313,N_24591);
or U26294 (N_26294,N_24909,N_25012);
or U26295 (N_26295,N_24511,N_24670);
nand U26296 (N_26296,N_24063,N_24402);
and U26297 (N_26297,N_24986,N_25191);
xor U26298 (N_26298,N_24732,N_25035);
or U26299 (N_26299,N_24415,N_24774);
nor U26300 (N_26300,N_24982,N_24285);
or U26301 (N_26301,N_24963,N_25186);
nor U26302 (N_26302,N_24046,N_24378);
or U26303 (N_26303,N_24820,N_24606);
and U26304 (N_26304,N_24283,N_24136);
and U26305 (N_26305,N_24825,N_25001);
or U26306 (N_26306,N_24919,N_24642);
or U26307 (N_26307,N_24901,N_24334);
xnor U26308 (N_26308,N_24824,N_25158);
xnor U26309 (N_26309,N_24857,N_24109);
or U26310 (N_26310,N_24021,N_24420);
and U26311 (N_26311,N_24545,N_24965);
or U26312 (N_26312,N_25101,N_24494);
nor U26313 (N_26313,N_24212,N_24087);
and U26314 (N_26314,N_24418,N_24535);
nor U26315 (N_26315,N_24129,N_24546);
and U26316 (N_26316,N_25091,N_24630);
and U26317 (N_26317,N_24118,N_25084);
or U26318 (N_26318,N_24409,N_24386);
nand U26319 (N_26319,N_24748,N_24000);
nor U26320 (N_26320,N_24669,N_25134);
xnor U26321 (N_26321,N_24803,N_24403);
and U26322 (N_26322,N_25167,N_24479);
xnor U26323 (N_26323,N_25108,N_24334);
and U26324 (N_26324,N_25039,N_24216);
nand U26325 (N_26325,N_24423,N_24153);
nor U26326 (N_26326,N_24822,N_25081);
nor U26327 (N_26327,N_24378,N_25115);
xnor U26328 (N_26328,N_24674,N_24364);
and U26329 (N_26329,N_24242,N_24650);
nor U26330 (N_26330,N_24394,N_25197);
or U26331 (N_26331,N_24571,N_24082);
nor U26332 (N_26332,N_24032,N_24867);
or U26333 (N_26333,N_24914,N_24020);
nand U26334 (N_26334,N_25130,N_24840);
or U26335 (N_26335,N_24594,N_24988);
and U26336 (N_26336,N_25141,N_25171);
or U26337 (N_26337,N_24444,N_25181);
or U26338 (N_26338,N_24046,N_24959);
and U26339 (N_26339,N_24691,N_24693);
nand U26340 (N_26340,N_24588,N_24152);
or U26341 (N_26341,N_24784,N_24765);
and U26342 (N_26342,N_24183,N_24256);
and U26343 (N_26343,N_24173,N_24729);
xnor U26344 (N_26344,N_25002,N_24516);
nand U26345 (N_26345,N_24415,N_25155);
nand U26346 (N_26346,N_24019,N_25167);
nand U26347 (N_26347,N_25167,N_24145);
and U26348 (N_26348,N_25064,N_24639);
nand U26349 (N_26349,N_24823,N_25195);
or U26350 (N_26350,N_25034,N_24961);
nand U26351 (N_26351,N_24622,N_25190);
and U26352 (N_26352,N_24771,N_25028);
nand U26353 (N_26353,N_25083,N_24951);
nand U26354 (N_26354,N_24035,N_24192);
nor U26355 (N_26355,N_24567,N_24132);
and U26356 (N_26356,N_24932,N_24621);
and U26357 (N_26357,N_24268,N_25129);
and U26358 (N_26358,N_24223,N_24990);
nor U26359 (N_26359,N_24880,N_24376);
nand U26360 (N_26360,N_24573,N_24670);
xnor U26361 (N_26361,N_24768,N_24046);
or U26362 (N_26362,N_24112,N_25192);
or U26363 (N_26363,N_24695,N_24171);
nor U26364 (N_26364,N_25085,N_24594);
xnor U26365 (N_26365,N_24136,N_24337);
and U26366 (N_26366,N_24028,N_25050);
and U26367 (N_26367,N_24706,N_25135);
and U26368 (N_26368,N_24667,N_24637);
nand U26369 (N_26369,N_24039,N_24913);
nand U26370 (N_26370,N_24324,N_24577);
nor U26371 (N_26371,N_24159,N_24818);
nor U26372 (N_26372,N_24213,N_24060);
and U26373 (N_26373,N_24868,N_24989);
or U26374 (N_26374,N_24088,N_24265);
or U26375 (N_26375,N_24170,N_24815);
nor U26376 (N_26376,N_24564,N_24290);
xnor U26377 (N_26377,N_24488,N_25076);
or U26378 (N_26378,N_24556,N_24265);
xor U26379 (N_26379,N_24269,N_24188);
or U26380 (N_26380,N_24534,N_25141);
nand U26381 (N_26381,N_24578,N_24538);
and U26382 (N_26382,N_25142,N_24010);
nor U26383 (N_26383,N_24930,N_24186);
and U26384 (N_26384,N_24533,N_24123);
nand U26385 (N_26385,N_24180,N_24497);
nand U26386 (N_26386,N_24737,N_24938);
and U26387 (N_26387,N_24409,N_24380);
nand U26388 (N_26388,N_24003,N_25196);
nor U26389 (N_26389,N_24754,N_24321);
or U26390 (N_26390,N_25071,N_24893);
and U26391 (N_26391,N_24439,N_25179);
or U26392 (N_26392,N_24570,N_25164);
or U26393 (N_26393,N_24820,N_24025);
and U26394 (N_26394,N_24905,N_24401);
nand U26395 (N_26395,N_24442,N_24077);
xor U26396 (N_26396,N_24628,N_24733);
nor U26397 (N_26397,N_25140,N_24000);
xor U26398 (N_26398,N_24673,N_24849);
and U26399 (N_26399,N_24131,N_24954);
nor U26400 (N_26400,N_26337,N_25287);
or U26401 (N_26401,N_26323,N_26386);
or U26402 (N_26402,N_25668,N_26085);
nand U26403 (N_26403,N_25670,N_25643);
and U26404 (N_26404,N_25737,N_26032);
and U26405 (N_26405,N_25797,N_25838);
or U26406 (N_26406,N_25993,N_26017);
or U26407 (N_26407,N_25404,N_25754);
nor U26408 (N_26408,N_25834,N_25261);
or U26409 (N_26409,N_25704,N_25305);
nand U26410 (N_26410,N_26345,N_25269);
nor U26411 (N_26411,N_26223,N_25259);
xnor U26412 (N_26412,N_26182,N_26068);
xnor U26413 (N_26413,N_25553,N_25784);
xnor U26414 (N_26414,N_25612,N_25680);
and U26415 (N_26415,N_25381,N_26153);
nor U26416 (N_26416,N_26269,N_25209);
or U26417 (N_26417,N_25473,N_25839);
nor U26418 (N_26418,N_25501,N_25689);
or U26419 (N_26419,N_26061,N_26309);
nand U26420 (N_26420,N_25225,N_25367);
or U26421 (N_26421,N_26237,N_26366);
nand U26422 (N_26422,N_25571,N_25953);
or U26423 (N_26423,N_26267,N_26272);
nor U26424 (N_26424,N_26106,N_25851);
and U26425 (N_26425,N_26236,N_25540);
xor U26426 (N_26426,N_26071,N_25429);
or U26427 (N_26427,N_26308,N_25384);
or U26428 (N_26428,N_25854,N_26358);
nand U26429 (N_26429,N_26095,N_26203);
and U26430 (N_26430,N_25949,N_26098);
nor U26431 (N_26431,N_26190,N_25943);
and U26432 (N_26432,N_25349,N_26086);
nand U26433 (N_26433,N_26041,N_25685);
xor U26434 (N_26434,N_25466,N_26245);
xor U26435 (N_26435,N_26283,N_25999);
and U26436 (N_26436,N_25471,N_25246);
or U26437 (N_26437,N_25371,N_25551);
xnor U26438 (N_26438,N_26076,N_26087);
nor U26439 (N_26439,N_25502,N_25911);
or U26440 (N_26440,N_26066,N_26026);
or U26441 (N_26441,N_26208,N_25430);
and U26442 (N_26442,N_25897,N_26325);
or U26443 (N_26443,N_25334,N_26290);
xor U26444 (N_26444,N_25354,N_25324);
nor U26445 (N_26445,N_25688,N_26158);
xor U26446 (N_26446,N_25453,N_26392);
or U26447 (N_26447,N_25475,N_25550);
nor U26448 (N_26448,N_26051,N_26150);
xnor U26449 (N_26449,N_25974,N_26177);
and U26450 (N_26450,N_25344,N_25713);
or U26451 (N_26451,N_25403,N_25593);
nor U26452 (N_26452,N_25657,N_25989);
or U26453 (N_26453,N_25443,N_26099);
nand U26454 (N_26454,N_25478,N_25452);
nor U26455 (N_26455,N_26039,N_26151);
nor U26456 (N_26456,N_26102,N_26138);
or U26457 (N_26457,N_25929,N_25574);
nor U26458 (N_26458,N_25888,N_25458);
and U26459 (N_26459,N_25484,N_26217);
and U26460 (N_26460,N_25616,N_25948);
nor U26461 (N_26461,N_25772,N_26189);
or U26462 (N_26462,N_25849,N_26354);
or U26463 (N_26463,N_25856,N_25708);
nor U26464 (N_26464,N_26344,N_25927);
or U26465 (N_26465,N_26300,N_26214);
or U26466 (N_26466,N_25242,N_26383);
nand U26467 (N_26467,N_26378,N_25624);
nor U26468 (N_26468,N_25581,N_25207);
nand U26469 (N_26469,N_25614,N_26398);
and U26470 (N_26470,N_25248,N_25432);
nor U26471 (N_26471,N_26112,N_26002);
or U26472 (N_26472,N_25442,N_25707);
nor U26473 (N_26473,N_25237,N_25281);
xor U26474 (N_26474,N_25967,N_25831);
xnor U26475 (N_26475,N_25773,N_25961);
nand U26476 (N_26476,N_25303,N_25215);
xnor U26477 (N_26477,N_26265,N_26315);
nor U26478 (N_26478,N_25229,N_25279);
and U26479 (N_26479,N_25998,N_26012);
nor U26480 (N_26480,N_26389,N_26382);
nand U26481 (N_26481,N_25919,N_25687);
nand U26482 (N_26482,N_25480,N_26119);
xor U26483 (N_26483,N_26371,N_25368);
nand U26484 (N_26484,N_26171,N_26218);
and U26485 (N_26485,N_26063,N_26010);
nor U26486 (N_26486,N_25313,N_26376);
or U26487 (N_26487,N_25597,N_26336);
or U26488 (N_26488,N_25272,N_25992);
xnor U26489 (N_26489,N_25703,N_25861);
nand U26490 (N_26490,N_25330,N_25756);
or U26491 (N_26491,N_25232,N_25625);
xnor U26492 (N_26492,N_25814,N_26199);
nor U26493 (N_26493,N_26126,N_26259);
xor U26494 (N_26494,N_25759,N_25984);
xnor U26495 (N_26495,N_26205,N_26357);
or U26496 (N_26496,N_25309,N_25885);
xor U26497 (N_26497,N_25498,N_26155);
and U26498 (N_26498,N_25477,N_25348);
or U26499 (N_26499,N_25627,N_25677);
nand U26500 (N_26500,N_26121,N_25202);
xnor U26501 (N_26501,N_25629,N_25900);
and U26502 (N_26502,N_25801,N_26194);
xnor U26503 (N_26503,N_26341,N_26113);
and U26504 (N_26504,N_25321,N_25940);
xor U26505 (N_26505,N_25433,N_25291);
or U26506 (N_26506,N_25230,N_25813);
nand U26507 (N_26507,N_25251,N_25516);
and U26508 (N_26508,N_25370,N_26215);
or U26509 (N_26509,N_26221,N_25544);
nand U26510 (N_26510,N_25275,N_25575);
and U26511 (N_26511,N_25267,N_26124);
and U26512 (N_26512,N_25537,N_25561);
or U26513 (N_26513,N_25679,N_25996);
or U26514 (N_26514,N_25818,N_26100);
nor U26515 (N_26515,N_25448,N_26104);
and U26516 (N_26516,N_25892,N_25794);
and U26517 (N_26517,N_26249,N_25848);
nor U26518 (N_26518,N_26204,N_25988);
and U26519 (N_26519,N_26274,N_25307);
xor U26520 (N_26520,N_25363,N_25328);
or U26521 (N_26521,N_25735,N_25306);
nor U26522 (N_26522,N_25699,N_26110);
nand U26523 (N_26523,N_26390,N_26391);
nor U26524 (N_26524,N_26243,N_25422);
or U26525 (N_26525,N_25767,N_26096);
and U26526 (N_26526,N_25950,N_25636);
or U26527 (N_26527,N_25714,N_26050);
and U26528 (N_26528,N_25428,N_25592);
xnor U26529 (N_26529,N_25263,N_25669);
nor U26530 (N_26530,N_25378,N_26168);
nand U26531 (N_26531,N_25835,N_25775);
xnor U26532 (N_26532,N_25843,N_26052);
nor U26533 (N_26533,N_26288,N_26185);
and U26534 (N_26534,N_25506,N_25726);
and U26535 (N_26535,N_25341,N_25997);
nor U26536 (N_26536,N_25722,N_25783);
xnor U26537 (N_26537,N_26188,N_26084);
xor U26538 (N_26538,N_26338,N_26141);
and U26539 (N_26539,N_26340,N_25308);
nand U26540 (N_26540,N_26180,N_25605);
and U26541 (N_26541,N_26235,N_26228);
nand U26542 (N_26542,N_26329,N_26310);
xor U26543 (N_26543,N_25470,N_25810);
nand U26544 (N_26544,N_26263,N_25619);
xnor U26545 (N_26545,N_25638,N_25832);
or U26546 (N_26546,N_25730,N_26319);
or U26547 (N_26547,N_26014,N_26364);
nor U26548 (N_26548,N_25400,N_25690);
nor U26549 (N_26549,N_25678,N_25760);
or U26550 (N_26550,N_25734,N_26081);
or U26551 (N_26551,N_25482,N_25720);
nand U26552 (N_26552,N_25304,N_26388);
and U26553 (N_26553,N_25782,N_25650);
or U26554 (N_26554,N_26024,N_25938);
xor U26555 (N_26555,N_25695,N_26139);
nor U26556 (N_26556,N_25513,N_26307);
or U26557 (N_26557,N_25807,N_26143);
nor U26558 (N_26558,N_26105,N_26373);
nand U26559 (N_26559,N_26006,N_25828);
and U26560 (N_26560,N_26030,N_25790);
nor U26561 (N_26561,N_25414,N_26278);
and U26562 (N_26562,N_26036,N_25408);
and U26563 (N_26563,N_26046,N_25211);
nand U26564 (N_26564,N_25282,N_25770);
nor U26565 (N_26565,N_25978,N_26294);
or U26566 (N_26566,N_26266,N_26167);
nand U26567 (N_26567,N_26174,N_25745);
nor U26568 (N_26568,N_25504,N_25380);
or U26569 (N_26569,N_26367,N_25682);
and U26570 (N_26570,N_26216,N_25672);
or U26571 (N_26571,N_25904,N_26054);
and U26572 (N_26572,N_26231,N_25800);
xor U26573 (N_26573,N_25869,N_25623);
xnor U26574 (N_26574,N_25547,N_26077);
or U26575 (N_26575,N_25976,N_25542);
nor U26576 (N_26576,N_25977,N_25931);
nand U26577 (N_26577,N_25254,N_25583);
nor U26578 (N_26578,N_25595,N_25821);
nand U26579 (N_26579,N_26240,N_26239);
or U26580 (N_26580,N_25427,N_25965);
xor U26581 (N_26581,N_25910,N_26043);
nand U26582 (N_26582,N_25434,N_25902);
nand U26583 (N_26583,N_25509,N_25539);
nand U26584 (N_26584,N_25780,N_25260);
and U26585 (N_26585,N_26232,N_26279);
nand U26586 (N_26586,N_25994,N_26207);
or U26587 (N_26587,N_25683,N_25865);
or U26588 (N_26588,N_25360,N_26275);
nor U26589 (N_26589,N_26005,N_25765);
or U26590 (N_26590,N_25449,N_25359);
or U26591 (N_26591,N_25750,N_26169);
nand U26592 (N_26592,N_25289,N_25294);
or U26593 (N_26593,N_25858,N_26175);
nor U26594 (N_26594,N_26314,N_26202);
and U26595 (N_26595,N_25573,N_25546);
and U26596 (N_26596,N_26089,N_25985);
nand U26597 (N_26597,N_26109,N_26355);
xor U26598 (N_26598,N_26230,N_25292);
or U26599 (N_26599,N_25419,N_26082);
xor U26600 (N_26600,N_25374,N_25375);
xor U26601 (N_26601,N_26132,N_26332);
xor U26602 (N_26602,N_25552,N_25957);
nor U26603 (N_26603,N_26211,N_25694);
nor U26604 (N_26604,N_26331,N_25920);
and U26605 (N_26605,N_25918,N_25755);
or U26606 (N_26606,N_25369,N_25671);
and U26607 (N_26607,N_26136,N_25764);
and U26608 (N_26608,N_26114,N_26342);
or U26609 (N_26609,N_25883,N_25447);
nor U26610 (N_26610,N_26281,N_26326);
nand U26611 (N_26611,N_26349,N_25325);
nand U26612 (N_26612,N_25709,N_25317);
or U26613 (N_26613,N_25778,N_25589);
nand U26614 (N_26614,N_25836,N_25667);
nand U26615 (N_26615,N_26312,N_25896);
or U26616 (N_26616,N_26353,N_26397);
or U26617 (N_26617,N_26261,N_25675);
nand U26618 (N_26618,N_25200,N_25492);
nor U26619 (N_26619,N_26187,N_25523);
nor U26620 (N_26620,N_25223,N_26317);
nand U26621 (N_26621,N_25594,N_25364);
and U26622 (N_26622,N_26250,N_25837);
nand U26623 (N_26623,N_25362,N_26111);
and U26624 (N_26624,N_25298,N_25356);
and U26625 (N_26625,N_26343,N_25796);
xnor U26626 (N_26626,N_25580,N_25365);
and U26627 (N_26627,N_26154,N_26387);
nor U26628 (N_26628,N_25852,N_25468);
nand U26629 (N_26629,N_25728,N_26303);
xnor U26630 (N_26630,N_25236,N_25457);
xnor U26631 (N_26631,N_25895,N_26131);
nand U26632 (N_26632,N_25941,N_26293);
xor U26633 (N_26633,N_25626,N_26271);
and U26634 (N_26634,N_25867,N_25340);
xor U26635 (N_26635,N_25717,N_25959);
and U26636 (N_26636,N_25405,N_25226);
or U26637 (N_26637,N_25534,N_25841);
xnor U26638 (N_26638,N_25995,N_25829);
xor U26639 (N_26639,N_25411,N_26328);
xnor U26640 (N_26640,N_25753,N_25500);
nand U26641 (N_26641,N_26396,N_26226);
and U26642 (N_26642,N_25339,N_25859);
nand U26643 (N_26643,N_25766,N_25535);
xor U26644 (N_26644,N_25273,N_26322);
and U26645 (N_26645,N_25747,N_26210);
nor U26646 (N_26646,N_26011,N_25373);
xnor U26647 (N_26647,N_25845,N_25617);
and U26648 (N_26648,N_25227,N_26127);
nor U26649 (N_26649,N_25877,N_26140);
xnor U26650 (N_26650,N_26000,N_25438);
or U26651 (N_26651,N_26304,N_26257);
and U26652 (N_26652,N_25460,N_25873);
nor U26653 (N_26653,N_25548,N_26037);
and U26654 (N_26654,N_25576,N_25630);
and U26655 (N_26655,N_26393,N_25761);
and U26656 (N_26656,N_26248,N_26351);
xnor U26657 (N_26657,N_26365,N_25257);
and U26658 (N_26658,N_26166,N_25798);
nand U26659 (N_26659,N_26260,N_25803);
xnor U26660 (N_26660,N_25450,N_25284);
and U26661 (N_26661,N_25295,N_26198);
xnor U26662 (N_26662,N_25712,N_25811);
and U26663 (N_26663,N_26003,N_26135);
and U26664 (N_26664,N_26380,N_25206);
nand U26665 (N_26665,N_25244,N_25774);
nor U26666 (N_26666,N_26254,N_25543);
and U26667 (N_26667,N_25386,N_26262);
nor U26668 (N_26668,N_26056,N_25673);
nand U26669 (N_26669,N_25203,N_26035);
or U26670 (N_26670,N_25799,N_25596);
and U26671 (N_26671,N_25632,N_26146);
xnor U26672 (N_26672,N_25771,N_25610);
xnor U26673 (N_26673,N_25916,N_25401);
nand U26674 (N_26674,N_26381,N_25345);
or U26675 (N_26675,N_25567,N_25210);
nor U26676 (N_26676,N_25607,N_25701);
and U26677 (N_26677,N_25744,N_26137);
nand U26678 (N_26678,N_25748,N_25486);
xnor U26679 (N_26679,N_25641,N_25319);
nand U26680 (N_26680,N_26055,N_26350);
nand U26681 (N_26681,N_25901,N_25969);
and U26682 (N_26682,N_25216,N_25817);
nand U26683 (N_26683,N_26129,N_25991);
xnor U26684 (N_26684,N_25266,N_25819);
or U26685 (N_26685,N_25599,N_25826);
xor U26686 (N_26686,N_26133,N_26399);
xor U26687 (N_26687,N_26369,N_25739);
nand U26688 (N_26688,N_25644,N_25742);
xor U26689 (N_26689,N_26040,N_26222);
or U26690 (N_26690,N_25928,N_25436);
and U26691 (N_26691,N_25461,N_25326);
xor U26692 (N_26692,N_25662,N_25327);
xnor U26693 (N_26693,N_25472,N_26144);
and U26694 (N_26694,N_25337,N_26333);
nor U26695 (N_26695,N_26027,N_25440);
nor U26696 (N_26696,N_25923,N_26128);
xor U26697 (N_26697,N_25822,N_26280);
xnor U26698 (N_26698,N_25201,N_25787);
nand U26699 (N_26699,N_25417,N_25406);
and U26700 (N_26700,N_25323,N_25347);
xor U26701 (N_26701,N_25474,N_25591);
nand U26702 (N_26702,N_25299,N_26092);
nor U26703 (N_26703,N_25875,N_25924);
or U26704 (N_26704,N_25585,N_25280);
and U26705 (N_26705,N_25329,N_26339);
and U26706 (N_26706,N_26394,N_25914);
xnor U26707 (N_26707,N_25857,N_25389);
and U26708 (N_26708,N_25481,N_26184);
nor U26709 (N_26709,N_25264,N_25270);
nor U26710 (N_26710,N_25749,N_26117);
nor U26711 (N_26711,N_26251,N_25970);
or U26712 (N_26712,N_26224,N_26286);
xor U26713 (N_26713,N_25973,N_25862);
nor U26714 (N_26714,N_25318,N_25986);
and U26715 (N_26715,N_25681,N_26079);
or U26716 (N_26716,N_26247,N_25524);
nand U26717 (N_26717,N_26330,N_26276);
or U26718 (N_26718,N_25606,N_25410);
or U26719 (N_26719,N_25391,N_25558);
or U26720 (N_26720,N_25247,N_26074);
xnor U26721 (N_26721,N_25250,N_25532);
xnor U26722 (N_26722,N_26318,N_25954);
xnor U26723 (N_26723,N_25565,N_25265);
nor U26724 (N_26724,N_26152,N_26384);
or U26725 (N_26725,N_25850,N_25934);
xnor U26726 (N_26726,N_25972,N_25424);
nor U26727 (N_26727,N_25881,N_26327);
xnor U26728 (N_26728,N_25249,N_25520);
or U26729 (N_26729,N_26229,N_25393);
nor U26730 (N_26730,N_25785,N_26324);
or U26731 (N_26731,N_25646,N_25412);
xor U26732 (N_26732,N_25820,N_25510);
and U26733 (N_26733,N_25651,N_25512);
and U26734 (N_26734,N_25912,N_26164);
xor U26735 (N_26735,N_25431,N_25635);
or U26736 (N_26736,N_25331,N_25398);
xor U26737 (N_26737,N_26062,N_25878);
nor U26738 (N_26738,N_25971,N_26159);
or U26739 (N_26739,N_25377,N_25531);
xor U26740 (N_26740,N_25777,N_26334);
or U26741 (N_26741,N_25816,N_25301);
nor U26742 (N_26742,N_25894,N_25312);
nand U26743 (N_26743,N_25219,N_26372);
and U26744 (N_26744,N_25715,N_25732);
or U26745 (N_26745,N_25930,N_25666);
nor U26746 (N_26746,N_25598,N_25926);
xor U26747 (N_26747,N_25587,N_25383);
nand U26748 (N_26748,N_25618,N_25351);
nand U26749 (N_26749,N_25958,N_26277);
nand U26750 (N_26750,N_26157,N_26118);
and U26751 (N_26751,N_25889,N_26219);
or U26752 (N_26752,N_25469,N_25310);
or U26753 (N_26753,N_26311,N_26346);
xnor U26754 (N_26754,N_25654,N_25743);
or U26755 (N_26755,N_25917,N_25653);
nand U26756 (N_26756,N_25352,N_26108);
nand U26757 (N_26757,N_25376,N_26255);
or U26758 (N_26758,N_25674,N_26073);
and U26759 (N_26759,N_25494,N_26170);
or U26760 (N_26760,N_26178,N_25659);
nand U26761 (N_26761,N_25982,N_25420);
or U26762 (N_26762,N_25533,N_25256);
and U26763 (N_26763,N_26183,N_25724);
and U26764 (N_26764,N_25647,N_26197);
nor U26765 (N_26765,N_25692,N_25907);
and U26766 (N_26766,N_25827,N_26088);
nor U26767 (N_26767,N_26091,N_25763);
xnor U26768 (N_26768,N_26292,N_26008);
and U26769 (N_26769,N_25621,N_26161);
nor U26770 (N_26770,N_25932,N_26045);
nand U26771 (N_26771,N_26298,N_25416);
or U26772 (N_26772,N_25757,N_25719);
xnor U26773 (N_26773,N_25795,N_25566);
xnor U26774 (N_26774,N_25615,N_25824);
nor U26775 (N_26775,N_25963,N_25684);
nand U26776 (N_26776,N_26356,N_25898);
or U26777 (N_26777,N_25538,N_25385);
nand U26778 (N_26778,N_26352,N_25268);
xor U26779 (N_26779,N_26241,N_25517);
nor U26780 (N_26780,N_25915,N_25245);
or U26781 (N_26781,N_26107,N_25353);
xnor U26782 (N_26782,N_26044,N_25947);
and U26783 (N_26783,N_25569,N_25788);
or U26784 (N_26784,N_25333,N_26284);
xnor U26785 (N_26785,N_25676,N_25490);
xnor U26786 (N_26786,N_25893,N_25476);
xnor U26787 (N_26787,N_26209,N_25577);
nor U26788 (N_26788,N_25456,N_25925);
nor U26789 (N_26789,N_26148,N_25559);
nor U26790 (N_26790,N_25903,N_25554);
nand U26791 (N_26791,N_25343,N_25387);
xor U26792 (N_26792,N_25527,N_25487);
nand U26793 (N_26793,N_25846,N_25608);
nor U26794 (N_26794,N_25979,N_25628);
xor U26795 (N_26795,N_25570,N_26165);
xor U26796 (N_26796,N_25741,N_25296);
and U26797 (N_26797,N_25253,N_26201);
nand U26798 (N_26798,N_25239,N_25224);
xnor U26799 (N_26799,N_25939,N_25241);
nand U26800 (N_26800,N_26029,N_25485);
nor U26801 (N_26801,N_25696,N_25886);
xor U26802 (N_26802,N_25658,N_25497);
and U26803 (N_26803,N_25437,N_25913);
xnor U26804 (N_26804,N_25853,N_26022);
or U26805 (N_26805,N_25395,N_26234);
nor U26806 (N_26806,N_25418,N_25711);
or U26807 (N_26807,N_26080,N_25705);
or U26808 (N_26808,N_25514,N_25981);
or U26809 (N_26809,N_25871,N_25840);
xnor U26810 (N_26810,N_25402,N_25451);
and U26811 (N_26811,N_26238,N_26038);
and U26812 (N_26812,N_25311,N_25776);
or U26813 (N_26813,N_26075,N_25952);
xor U26814 (N_26814,N_25718,N_26048);
or U26815 (N_26815,N_25283,N_26244);
or U26816 (N_26816,N_26034,N_25661);
nand U26817 (N_26817,N_25231,N_25293);
and U26818 (N_26818,N_25505,N_26149);
xnor U26819 (N_26819,N_25611,N_25951);
and U26820 (N_26820,N_26285,N_25738);
and U26821 (N_26821,N_26060,N_25483);
nor U26822 (N_26822,N_25459,N_26142);
and U26823 (N_26823,N_26007,N_25648);
nand U26824 (N_26824,N_25302,N_25413);
xor U26825 (N_26825,N_25721,N_26227);
nand U26826 (N_26826,N_26072,N_25208);
and U26827 (N_26827,N_25604,N_25495);
xor U26828 (N_26828,N_25518,N_25415);
nand U26829 (N_26829,N_25511,N_25652);
nand U26830 (N_26830,N_26302,N_25697);
xor U26831 (N_26831,N_25812,N_25286);
or U26832 (N_26832,N_25716,N_25698);
xor U26833 (N_26833,N_26374,N_25663);
or U26834 (N_26834,N_25602,N_26359);
and U26835 (N_26835,N_26147,N_25786);
or U26836 (N_26836,N_25921,N_25880);
or U26837 (N_26837,N_25465,N_25507);
or U26838 (N_26838,N_25631,N_25613);
or U26839 (N_26839,N_25276,N_25751);
nor U26840 (N_26840,N_25278,N_26120);
nor U26841 (N_26841,N_25664,N_26009);
nand U26842 (N_26842,N_26375,N_25536);
nand U26843 (N_26843,N_25693,N_25758);
xor U26844 (N_26844,N_25884,N_25467);
and U26845 (N_26845,N_26206,N_26134);
xnor U26846 (N_26846,N_25221,N_25503);
nor U26847 (N_26847,N_25445,N_26103);
or U26848 (N_26848,N_25691,N_26173);
nor U26849 (N_26849,N_26116,N_26016);
or U26850 (N_26850,N_25409,N_25937);
nor U26851 (N_26851,N_26145,N_25590);
nor U26852 (N_26852,N_25336,N_25423);
and U26853 (N_26853,N_26273,N_25700);
or U26854 (N_26854,N_25463,N_25545);
nor U26855 (N_26855,N_26053,N_25962);
nand U26856 (N_26856,N_25521,N_25966);
nor U26857 (N_26857,N_25252,N_25665);
nor U26858 (N_26858,N_26023,N_26196);
nor U26859 (N_26859,N_25656,N_25890);
nand U26860 (N_26860,N_25499,N_25358);
and U26861 (N_26861,N_25355,N_25218);
or U26862 (N_26862,N_26160,N_25866);
and U26863 (N_26863,N_25600,N_25342);
xor U26864 (N_26864,N_25955,N_25335);
xnor U26865 (N_26865,N_26242,N_26335);
and U26866 (N_26866,N_26191,N_25842);
xnor U26867 (N_26867,N_25922,N_25882);
and U26868 (N_26868,N_25562,N_25396);
or U26869 (N_26869,N_25568,N_25825);
nor U26870 (N_26870,N_25488,N_25390);
and U26871 (N_26871,N_25235,N_25909);
xnor U26872 (N_26872,N_26019,N_26057);
or U26873 (N_26873,N_26093,N_25238);
xor U26874 (N_26874,N_26395,N_25815);
and U26875 (N_26875,N_25526,N_26094);
nand U26876 (N_26876,N_25529,N_26186);
nand U26877 (N_26877,N_25762,N_26172);
and U26878 (N_26878,N_25563,N_25556);
and U26879 (N_26879,N_25781,N_26291);
or U26880 (N_26880,N_25425,N_26101);
nor U26881 (N_26881,N_25315,N_25946);
nand U26882 (N_26882,N_25746,N_25833);
and U26883 (N_26883,N_26047,N_26301);
nor U26884 (N_26884,N_26069,N_25601);
or U26885 (N_26885,N_25805,N_25723);
and U26886 (N_26886,N_25320,N_25258);
nand U26887 (N_26887,N_26233,N_26049);
and U26888 (N_26888,N_25768,N_26316);
xor U26889 (N_26889,N_25655,N_25397);
and U26890 (N_26890,N_26031,N_26252);
and U26891 (N_26891,N_26122,N_26195);
nand U26892 (N_26892,N_25809,N_25462);
and U26893 (N_26893,N_26001,N_25528);
and U26894 (N_26894,N_25454,N_26287);
xor U26895 (N_26895,N_25964,N_25769);
nor U26896 (N_26896,N_26033,N_26320);
xnor U26897 (N_26897,N_25300,N_25564);
nor U26898 (N_26898,N_25297,N_25572);
or U26899 (N_26899,N_26156,N_26018);
or U26900 (N_26900,N_26313,N_26021);
xor U26901 (N_26901,N_26212,N_25285);
and U26902 (N_26902,N_25891,N_25727);
nor U26903 (N_26903,N_26299,N_25515);
xnor U26904 (N_26904,N_25372,N_25455);
xnor U26905 (N_26905,N_25983,N_25530);
or U26906 (N_26906,N_25622,N_25361);
xnor U26907 (N_26907,N_25779,N_25649);
or U26908 (N_26908,N_25508,N_25640);
and U26909 (N_26909,N_25860,N_25710);
nor U26910 (N_26910,N_25350,N_25394);
nor U26911 (N_26911,N_25870,N_25525);
nand U26912 (N_26912,N_26306,N_25578);
and U26913 (N_26913,N_25464,N_26379);
and U26914 (N_26914,N_25634,N_25322);
and U26915 (N_26915,N_26163,N_25560);
and U26916 (N_26916,N_26282,N_25586);
and U26917 (N_26917,N_25990,N_26065);
and U26918 (N_26918,N_25868,N_25582);
nor U26919 (N_26919,N_25942,N_25314);
nor U26920 (N_26920,N_25399,N_25332);
or U26921 (N_26921,N_25555,N_25435);
nand U26922 (N_26922,N_25346,N_25729);
or U26923 (N_26923,N_26078,N_25855);
nor U26924 (N_26924,N_25935,N_25639);
and U26925 (N_26925,N_25802,N_26361);
nand U26926 (N_26926,N_25887,N_26295);
xnor U26927 (N_26927,N_26115,N_25493);
xor U26928 (N_26928,N_26015,N_26246);
nor U26929 (N_26929,N_25980,N_26362);
or U26930 (N_26930,N_26348,N_25357);
xor U26931 (N_26931,N_25222,N_25686);
or U26932 (N_26932,N_26130,N_25905);
and U26933 (N_26933,N_25220,N_25876);
or U26934 (N_26934,N_25584,N_26025);
nor U26935 (N_26935,N_25933,N_26058);
or U26936 (N_26936,N_25874,N_25706);
xnor U26937 (N_26937,N_26004,N_25379);
and U26938 (N_26938,N_26347,N_26225);
or U26939 (N_26939,N_25491,N_25213);
nand U26940 (N_26940,N_25872,N_26377);
or U26941 (N_26941,N_26253,N_25863);
or U26942 (N_26942,N_25603,N_26028);
nand U26943 (N_26943,N_25906,N_25262);
or U26944 (N_26944,N_25725,N_25702);
nand U26945 (N_26945,N_25228,N_25444);
nor U26946 (N_26946,N_26360,N_25944);
nor U26947 (N_26947,N_25233,N_25366);
and U26948 (N_26948,N_25271,N_25960);
xnor U26949 (N_26949,N_25733,N_25426);
nand U26950 (N_26950,N_25620,N_25288);
nor U26951 (N_26951,N_25255,N_25240);
nand U26952 (N_26952,N_25234,N_26370);
nor U26953 (N_26953,N_26305,N_26268);
and U26954 (N_26954,N_25806,N_25290);
or U26955 (N_26955,N_26179,N_25316);
xor U26956 (N_26956,N_25945,N_26193);
or U26957 (N_26957,N_26270,N_25645);
nand U26958 (N_26958,N_25899,N_25879);
xnor U26959 (N_26959,N_26125,N_26097);
or U26960 (N_26960,N_26297,N_26200);
xnor U26961 (N_26961,N_25987,N_26296);
xor U26962 (N_26962,N_25864,N_25736);
nor U26963 (N_26963,N_25633,N_26162);
or U26964 (N_26964,N_26368,N_25479);
and U26965 (N_26965,N_25792,N_25217);
and U26966 (N_26966,N_25908,N_25274);
nand U26967 (N_26967,N_26220,N_26070);
nor U26968 (N_26968,N_25731,N_25847);
or U26969 (N_26969,N_26264,N_25496);
and U26970 (N_26970,N_25205,N_26181);
or U26971 (N_26971,N_25557,N_25382);
nor U26972 (N_26972,N_25637,N_26090);
nand U26973 (N_26973,N_26013,N_25642);
nor U26974 (N_26974,N_26385,N_25441);
nand U26975 (N_26975,N_25522,N_25214);
or U26976 (N_26976,N_25609,N_25956);
nand U26977 (N_26977,N_26064,N_26256);
xnor U26978 (N_26978,N_25579,N_25243);
or U26979 (N_26979,N_26123,N_25277);
or U26980 (N_26980,N_25789,N_25968);
and U26981 (N_26981,N_26020,N_26059);
xnor U26982 (N_26982,N_25549,N_25740);
nand U26983 (N_26983,N_25204,N_26192);
or U26984 (N_26984,N_25793,N_25975);
nand U26985 (N_26985,N_26042,N_25212);
nand U26986 (N_26986,N_26289,N_25407);
or U26987 (N_26987,N_26363,N_25388);
nor U26988 (N_26988,N_25541,N_25752);
xor U26989 (N_26989,N_25936,N_26258);
or U26990 (N_26990,N_25421,N_25823);
nor U26991 (N_26991,N_25439,N_25338);
or U26992 (N_26992,N_26083,N_25588);
or U26993 (N_26993,N_25392,N_26176);
xor U26994 (N_26994,N_25519,N_25808);
nor U26995 (N_26995,N_25446,N_25804);
nor U26996 (N_26996,N_25791,N_26321);
and U26997 (N_26997,N_26213,N_25844);
nor U26998 (N_26998,N_26067,N_25660);
nor U26999 (N_26999,N_25489,N_25830);
and U27000 (N_27000,N_25630,N_26232);
xnor U27001 (N_27001,N_25611,N_26294);
nand U27002 (N_27002,N_26284,N_26112);
nand U27003 (N_27003,N_26080,N_25202);
or U27004 (N_27004,N_26345,N_25677);
nor U27005 (N_27005,N_25836,N_26330);
or U27006 (N_27006,N_26236,N_25558);
and U27007 (N_27007,N_25923,N_25773);
or U27008 (N_27008,N_25460,N_25843);
xor U27009 (N_27009,N_25948,N_25708);
and U27010 (N_27010,N_26045,N_25570);
nand U27011 (N_27011,N_25596,N_25534);
and U27012 (N_27012,N_26025,N_25911);
and U27013 (N_27013,N_25373,N_25371);
or U27014 (N_27014,N_26131,N_25269);
xor U27015 (N_27015,N_26380,N_25762);
xnor U27016 (N_27016,N_25296,N_25801);
xor U27017 (N_27017,N_26390,N_25309);
nand U27018 (N_27018,N_25237,N_26382);
nor U27019 (N_27019,N_25852,N_26362);
xor U27020 (N_27020,N_25521,N_26226);
nand U27021 (N_27021,N_25393,N_25705);
or U27022 (N_27022,N_26238,N_25660);
and U27023 (N_27023,N_25200,N_25747);
and U27024 (N_27024,N_26345,N_25787);
xnor U27025 (N_27025,N_25727,N_25247);
xnor U27026 (N_27026,N_26055,N_25454);
nor U27027 (N_27027,N_26039,N_25980);
and U27028 (N_27028,N_25756,N_26046);
or U27029 (N_27029,N_25850,N_25266);
nand U27030 (N_27030,N_25584,N_25366);
or U27031 (N_27031,N_25854,N_26230);
nand U27032 (N_27032,N_25852,N_25260);
nor U27033 (N_27033,N_25588,N_25657);
xnor U27034 (N_27034,N_26348,N_25367);
or U27035 (N_27035,N_26392,N_25950);
xnor U27036 (N_27036,N_25203,N_25357);
nor U27037 (N_27037,N_25893,N_25498);
xor U27038 (N_27038,N_25520,N_25655);
nand U27039 (N_27039,N_25573,N_26072);
or U27040 (N_27040,N_26194,N_26192);
or U27041 (N_27041,N_25929,N_26261);
and U27042 (N_27042,N_25952,N_26069);
nor U27043 (N_27043,N_26012,N_25952);
nor U27044 (N_27044,N_25524,N_25418);
xnor U27045 (N_27045,N_26102,N_25539);
and U27046 (N_27046,N_25890,N_26267);
xnor U27047 (N_27047,N_26374,N_26028);
or U27048 (N_27048,N_25230,N_26265);
nand U27049 (N_27049,N_26235,N_25747);
or U27050 (N_27050,N_25482,N_26066);
nor U27051 (N_27051,N_26157,N_25942);
nand U27052 (N_27052,N_25394,N_26209);
nor U27053 (N_27053,N_25743,N_26394);
or U27054 (N_27054,N_26343,N_25473);
nor U27055 (N_27055,N_26237,N_25414);
xnor U27056 (N_27056,N_26243,N_25636);
or U27057 (N_27057,N_25406,N_26194);
nor U27058 (N_27058,N_26314,N_26328);
and U27059 (N_27059,N_25509,N_25902);
nand U27060 (N_27060,N_25643,N_26207);
nor U27061 (N_27061,N_25944,N_25258);
and U27062 (N_27062,N_26310,N_25482);
or U27063 (N_27063,N_26143,N_25760);
nor U27064 (N_27064,N_25555,N_25972);
nor U27065 (N_27065,N_25649,N_26354);
nor U27066 (N_27066,N_25944,N_25378);
and U27067 (N_27067,N_26281,N_26324);
or U27068 (N_27068,N_26343,N_25716);
nand U27069 (N_27069,N_25940,N_25828);
and U27070 (N_27070,N_25806,N_25887);
nand U27071 (N_27071,N_26196,N_26174);
or U27072 (N_27072,N_25881,N_25617);
or U27073 (N_27073,N_26104,N_26194);
nand U27074 (N_27074,N_25398,N_25736);
nor U27075 (N_27075,N_25754,N_25745);
nor U27076 (N_27076,N_25906,N_26323);
xnor U27077 (N_27077,N_25257,N_26160);
nand U27078 (N_27078,N_25816,N_25686);
or U27079 (N_27079,N_25931,N_26026);
or U27080 (N_27080,N_26017,N_25202);
nor U27081 (N_27081,N_26031,N_26229);
nand U27082 (N_27082,N_25306,N_25890);
nor U27083 (N_27083,N_25586,N_26351);
or U27084 (N_27084,N_25881,N_25401);
nor U27085 (N_27085,N_26070,N_25670);
nor U27086 (N_27086,N_25607,N_26317);
nand U27087 (N_27087,N_25824,N_26121);
nor U27088 (N_27088,N_26210,N_25679);
nor U27089 (N_27089,N_26190,N_26272);
and U27090 (N_27090,N_25662,N_25448);
or U27091 (N_27091,N_26350,N_26304);
or U27092 (N_27092,N_26015,N_26224);
and U27093 (N_27093,N_25339,N_25242);
or U27094 (N_27094,N_25775,N_25666);
xnor U27095 (N_27095,N_25345,N_25595);
nor U27096 (N_27096,N_26332,N_26060);
nor U27097 (N_27097,N_26048,N_26022);
nand U27098 (N_27098,N_26220,N_26035);
or U27099 (N_27099,N_26300,N_25322);
and U27100 (N_27100,N_25912,N_25275);
xor U27101 (N_27101,N_25955,N_25502);
nor U27102 (N_27102,N_26237,N_26024);
xnor U27103 (N_27103,N_25825,N_26008);
or U27104 (N_27104,N_25468,N_26154);
and U27105 (N_27105,N_25380,N_26281);
nand U27106 (N_27106,N_25612,N_25440);
nand U27107 (N_27107,N_25637,N_25434);
or U27108 (N_27108,N_25696,N_25222);
xnor U27109 (N_27109,N_26083,N_25224);
or U27110 (N_27110,N_25316,N_25973);
nor U27111 (N_27111,N_25705,N_26203);
or U27112 (N_27112,N_26213,N_26239);
nor U27113 (N_27113,N_26347,N_25618);
nand U27114 (N_27114,N_26359,N_25316);
or U27115 (N_27115,N_25996,N_25253);
nor U27116 (N_27116,N_26161,N_26054);
nand U27117 (N_27117,N_25938,N_25591);
xor U27118 (N_27118,N_25757,N_26320);
xor U27119 (N_27119,N_26108,N_25566);
xnor U27120 (N_27120,N_26327,N_25669);
or U27121 (N_27121,N_25571,N_25798);
or U27122 (N_27122,N_26192,N_26281);
xor U27123 (N_27123,N_26045,N_26149);
nor U27124 (N_27124,N_26131,N_26020);
nor U27125 (N_27125,N_25364,N_25906);
nand U27126 (N_27126,N_25644,N_26226);
nor U27127 (N_27127,N_25799,N_25822);
or U27128 (N_27128,N_25905,N_26171);
nand U27129 (N_27129,N_26191,N_25424);
nand U27130 (N_27130,N_26035,N_25723);
and U27131 (N_27131,N_25961,N_25237);
and U27132 (N_27132,N_25249,N_26304);
nand U27133 (N_27133,N_25223,N_25420);
and U27134 (N_27134,N_25726,N_25975);
nor U27135 (N_27135,N_25750,N_25667);
or U27136 (N_27136,N_26156,N_26073);
and U27137 (N_27137,N_26378,N_26127);
or U27138 (N_27138,N_26180,N_26259);
nor U27139 (N_27139,N_25653,N_25923);
and U27140 (N_27140,N_25519,N_26052);
nor U27141 (N_27141,N_25879,N_26171);
or U27142 (N_27142,N_26345,N_25805);
nand U27143 (N_27143,N_25563,N_26085);
or U27144 (N_27144,N_26341,N_25261);
nand U27145 (N_27145,N_25532,N_25282);
nor U27146 (N_27146,N_26029,N_25368);
xnor U27147 (N_27147,N_26342,N_26100);
and U27148 (N_27148,N_25577,N_26328);
and U27149 (N_27149,N_25290,N_26172);
xor U27150 (N_27150,N_26326,N_26214);
and U27151 (N_27151,N_26091,N_26252);
and U27152 (N_27152,N_26281,N_25305);
nor U27153 (N_27153,N_26392,N_26154);
nand U27154 (N_27154,N_25559,N_25366);
nand U27155 (N_27155,N_26277,N_25254);
xnor U27156 (N_27156,N_25702,N_25349);
or U27157 (N_27157,N_26333,N_25827);
nor U27158 (N_27158,N_25330,N_25226);
nor U27159 (N_27159,N_25866,N_25688);
or U27160 (N_27160,N_26262,N_26360);
nor U27161 (N_27161,N_26267,N_26353);
nand U27162 (N_27162,N_26257,N_26184);
and U27163 (N_27163,N_26075,N_25420);
nor U27164 (N_27164,N_26350,N_26193);
nand U27165 (N_27165,N_26183,N_25415);
and U27166 (N_27166,N_25765,N_26136);
xor U27167 (N_27167,N_25414,N_25221);
xor U27168 (N_27168,N_26156,N_25650);
nor U27169 (N_27169,N_25322,N_26228);
or U27170 (N_27170,N_26220,N_25526);
or U27171 (N_27171,N_25309,N_25308);
nand U27172 (N_27172,N_25719,N_25608);
and U27173 (N_27173,N_25929,N_25265);
nand U27174 (N_27174,N_26251,N_25226);
or U27175 (N_27175,N_25396,N_25805);
xnor U27176 (N_27176,N_25842,N_25996);
or U27177 (N_27177,N_26356,N_26381);
or U27178 (N_27178,N_25331,N_26169);
nand U27179 (N_27179,N_25893,N_25612);
nor U27180 (N_27180,N_25532,N_25577);
nand U27181 (N_27181,N_25453,N_26126);
or U27182 (N_27182,N_26152,N_25696);
or U27183 (N_27183,N_25636,N_25432);
xnor U27184 (N_27184,N_25858,N_25696);
nand U27185 (N_27185,N_25813,N_25760);
or U27186 (N_27186,N_25497,N_26011);
xnor U27187 (N_27187,N_25687,N_25643);
or U27188 (N_27188,N_26133,N_25474);
nand U27189 (N_27189,N_26323,N_25202);
xnor U27190 (N_27190,N_25478,N_25473);
or U27191 (N_27191,N_25330,N_25703);
nand U27192 (N_27192,N_26275,N_26121);
nor U27193 (N_27193,N_26334,N_25993);
nor U27194 (N_27194,N_26363,N_25242);
xnor U27195 (N_27195,N_25646,N_25274);
or U27196 (N_27196,N_25521,N_25801);
nand U27197 (N_27197,N_26234,N_25647);
nand U27198 (N_27198,N_26157,N_25541);
and U27199 (N_27199,N_25580,N_26270);
nand U27200 (N_27200,N_25517,N_25978);
and U27201 (N_27201,N_25512,N_26180);
nor U27202 (N_27202,N_25299,N_25789);
xnor U27203 (N_27203,N_25559,N_25806);
xor U27204 (N_27204,N_25514,N_26122);
or U27205 (N_27205,N_25260,N_25882);
or U27206 (N_27206,N_26147,N_25502);
or U27207 (N_27207,N_26102,N_25207);
nand U27208 (N_27208,N_26370,N_25470);
nand U27209 (N_27209,N_26032,N_25342);
nand U27210 (N_27210,N_26150,N_25572);
and U27211 (N_27211,N_25352,N_25791);
nand U27212 (N_27212,N_25204,N_25884);
xnor U27213 (N_27213,N_26207,N_26080);
nor U27214 (N_27214,N_25725,N_26182);
or U27215 (N_27215,N_25907,N_25454);
and U27216 (N_27216,N_25603,N_25333);
xnor U27217 (N_27217,N_25253,N_25436);
or U27218 (N_27218,N_26100,N_25334);
and U27219 (N_27219,N_25976,N_25726);
nand U27220 (N_27220,N_26017,N_25297);
or U27221 (N_27221,N_25634,N_26374);
nor U27222 (N_27222,N_26001,N_26168);
and U27223 (N_27223,N_26001,N_25303);
xor U27224 (N_27224,N_25384,N_25677);
nor U27225 (N_27225,N_25271,N_26203);
xnor U27226 (N_27226,N_25925,N_25823);
or U27227 (N_27227,N_26319,N_26245);
nand U27228 (N_27228,N_25501,N_26396);
and U27229 (N_27229,N_26173,N_25356);
and U27230 (N_27230,N_25425,N_26318);
nand U27231 (N_27231,N_26035,N_25291);
or U27232 (N_27232,N_25919,N_25886);
nor U27233 (N_27233,N_26060,N_25280);
xnor U27234 (N_27234,N_25944,N_26130);
and U27235 (N_27235,N_26136,N_26128);
nand U27236 (N_27236,N_26378,N_25404);
nor U27237 (N_27237,N_25728,N_25296);
nand U27238 (N_27238,N_25951,N_26144);
or U27239 (N_27239,N_25380,N_26186);
nor U27240 (N_27240,N_25209,N_25974);
or U27241 (N_27241,N_25361,N_25878);
nor U27242 (N_27242,N_26311,N_25241);
nor U27243 (N_27243,N_25777,N_26275);
nand U27244 (N_27244,N_26111,N_25440);
nor U27245 (N_27245,N_25905,N_25430);
or U27246 (N_27246,N_25748,N_25749);
nand U27247 (N_27247,N_25394,N_25482);
xnor U27248 (N_27248,N_25324,N_25225);
or U27249 (N_27249,N_25592,N_25937);
or U27250 (N_27250,N_26210,N_26000);
nor U27251 (N_27251,N_25676,N_25923);
nor U27252 (N_27252,N_25890,N_26121);
or U27253 (N_27253,N_25212,N_25703);
and U27254 (N_27254,N_25507,N_25254);
or U27255 (N_27255,N_25805,N_25616);
xnor U27256 (N_27256,N_25217,N_26176);
or U27257 (N_27257,N_25900,N_26000);
xnor U27258 (N_27258,N_25646,N_25896);
or U27259 (N_27259,N_25648,N_25686);
nor U27260 (N_27260,N_26114,N_25714);
and U27261 (N_27261,N_26387,N_26145);
and U27262 (N_27262,N_26083,N_25360);
and U27263 (N_27263,N_26207,N_25713);
xnor U27264 (N_27264,N_26198,N_26383);
xor U27265 (N_27265,N_25855,N_25696);
nand U27266 (N_27266,N_25458,N_26039);
nor U27267 (N_27267,N_26100,N_25439);
xor U27268 (N_27268,N_25215,N_25572);
nand U27269 (N_27269,N_25766,N_25708);
or U27270 (N_27270,N_25815,N_25823);
nor U27271 (N_27271,N_25808,N_25610);
xnor U27272 (N_27272,N_26391,N_26073);
and U27273 (N_27273,N_25852,N_26070);
and U27274 (N_27274,N_26243,N_26377);
or U27275 (N_27275,N_26233,N_25287);
nor U27276 (N_27276,N_26149,N_25654);
nor U27277 (N_27277,N_25288,N_26386);
nor U27278 (N_27278,N_26103,N_25216);
nor U27279 (N_27279,N_25225,N_25416);
or U27280 (N_27280,N_26169,N_25827);
or U27281 (N_27281,N_25907,N_25301);
nand U27282 (N_27282,N_25225,N_25612);
xnor U27283 (N_27283,N_26381,N_25502);
xnor U27284 (N_27284,N_25254,N_25342);
or U27285 (N_27285,N_25496,N_26360);
or U27286 (N_27286,N_26120,N_25920);
nand U27287 (N_27287,N_25879,N_26265);
or U27288 (N_27288,N_25649,N_26278);
nor U27289 (N_27289,N_26181,N_25463);
nand U27290 (N_27290,N_25990,N_25729);
nand U27291 (N_27291,N_25550,N_26357);
xor U27292 (N_27292,N_25873,N_25912);
or U27293 (N_27293,N_26135,N_25509);
xor U27294 (N_27294,N_25625,N_25273);
nor U27295 (N_27295,N_25291,N_25438);
and U27296 (N_27296,N_26371,N_25854);
or U27297 (N_27297,N_25611,N_26330);
or U27298 (N_27298,N_25574,N_26165);
and U27299 (N_27299,N_25458,N_25319);
and U27300 (N_27300,N_26271,N_25932);
nor U27301 (N_27301,N_26132,N_26341);
or U27302 (N_27302,N_25629,N_26144);
nand U27303 (N_27303,N_26318,N_25902);
and U27304 (N_27304,N_26382,N_26167);
and U27305 (N_27305,N_25252,N_25845);
nor U27306 (N_27306,N_26114,N_25593);
nand U27307 (N_27307,N_25621,N_25718);
nand U27308 (N_27308,N_25651,N_26256);
and U27309 (N_27309,N_25241,N_25793);
xnor U27310 (N_27310,N_25244,N_25627);
nand U27311 (N_27311,N_25574,N_26151);
or U27312 (N_27312,N_25679,N_26234);
nand U27313 (N_27313,N_25969,N_25748);
or U27314 (N_27314,N_25967,N_26074);
and U27315 (N_27315,N_26168,N_25464);
nor U27316 (N_27316,N_26129,N_25276);
nand U27317 (N_27317,N_26304,N_25422);
xor U27318 (N_27318,N_25216,N_26392);
nand U27319 (N_27319,N_25694,N_25446);
or U27320 (N_27320,N_25552,N_26135);
nor U27321 (N_27321,N_25321,N_26328);
nand U27322 (N_27322,N_26337,N_25720);
xor U27323 (N_27323,N_26146,N_25505);
or U27324 (N_27324,N_25596,N_26363);
nor U27325 (N_27325,N_25453,N_26104);
and U27326 (N_27326,N_25691,N_25905);
and U27327 (N_27327,N_26027,N_25422);
nor U27328 (N_27328,N_26169,N_25816);
nand U27329 (N_27329,N_25333,N_25622);
and U27330 (N_27330,N_25286,N_25544);
xor U27331 (N_27331,N_25989,N_26388);
nand U27332 (N_27332,N_26394,N_25964);
xnor U27333 (N_27333,N_25424,N_25276);
and U27334 (N_27334,N_26381,N_26223);
nand U27335 (N_27335,N_25788,N_26246);
nand U27336 (N_27336,N_25576,N_25523);
nor U27337 (N_27337,N_26359,N_26251);
or U27338 (N_27338,N_25693,N_26030);
or U27339 (N_27339,N_26114,N_26168);
xor U27340 (N_27340,N_26386,N_25281);
and U27341 (N_27341,N_25635,N_25456);
nor U27342 (N_27342,N_25258,N_25370);
and U27343 (N_27343,N_25287,N_26017);
and U27344 (N_27344,N_25900,N_25874);
and U27345 (N_27345,N_25770,N_25251);
nand U27346 (N_27346,N_25794,N_25644);
and U27347 (N_27347,N_26399,N_25288);
xor U27348 (N_27348,N_25967,N_25426);
nor U27349 (N_27349,N_25323,N_25246);
or U27350 (N_27350,N_25791,N_25319);
nor U27351 (N_27351,N_25880,N_25236);
nand U27352 (N_27352,N_25481,N_26166);
and U27353 (N_27353,N_26342,N_26130);
xor U27354 (N_27354,N_26046,N_25977);
and U27355 (N_27355,N_26232,N_25295);
nand U27356 (N_27356,N_26226,N_25667);
and U27357 (N_27357,N_25949,N_26123);
nand U27358 (N_27358,N_25216,N_25694);
and U27359 (N_27359,N_25686,N_25972);
nor U27360 (N_27360,N_25909,N_26005);
xnor U27361 (N_27361,N_25951,N_25487);
xor U27362 (N_27362,N_25969,N_25553);
or U27363 (N_27363,N_25750,N_25402);
xor U27364 (N_27364,N_25707,N_25879);
and U27365 (N_27365,N_25712,N_25972);
nand U27366 (N_27366,N_25415,N_25660);
and U27367 (N_27367,N_25367,N_26050);
nand U27368 (N_27368,N_25378,N_26114);
nand U27369 (N_27369,N_25498,N_26103);
and U27370 (N_27370,N_26322,N_25394);
and U27371 (N_27371,N_25370,N_26383);
xor U27372 (N_27372,N_26261,N_26037);
or U27373 (N_27373,N_26010,N_25316);
nor U27374 (N_27374,N_26018,N_26145);
nand U27375 (N_27375,N_26324,N_26369);
or U27376 (N_27376,N_25720,N_25443);
nor U27377 (N_27377,N_26004,N_25726);
or U27378 (N_27378,N_26139,N_25848);
xor U27379 (N_27379,N_25743,N_26344);
nand U27380 (N_27380,N_25548,N_25543);
nor U27381 (N_27381,N_26134,N_26097);
nand U27382 (N_27382,N_25791,N_25655);
and U27383 (N_27383,N_25592,N_25467);
nor U27384 (N_27384,N_25372,N_25471);
or U27385 (N_27385,N_26315,N_25724);
or U27386 (N_27386,N_25945,N_25776);
and U27387 (N_27387,N_25206,N_26301);
xor U27388 (N_27388,N_25526,N_25825);
and U27389 (N_27389,N_26003,N_25767);
nor U27390 (N_27390,N_25881,N_25200);
nor U27391 (N_27391,N_26213,N_25993);
or U27392 (N_27392,N_25368,N_25857);
or U27393 (N_27393,N_26249,N_26085);
and U27394 (N_27394,N_25919,N_25883);
or U27395 (N_27395,N_25600,N_26175);
and U27396 (N_27396,N_25239,N_26389);
nor U27397 (N_27397,N_25478,N_26301);
nand U27398 (N_27398,N_26114,N_25740);
and U27399 (N_27399,N_26389,N_25558);
nor U27400 (N_27400,N_25535,N_25813);
or U27401 (N_27401,N_26101,N_26207);
or U27402 (N_27402,N_25465,N_25569);
nand U27403 (N_27403,N_25790,N_26241);
nor U27404 (N_27404,N_26074,N_25849);
or U27405 (N_27405,N_25384,N_25823);
nand U27406 (N_27406,N_25982,N_25501);
xor U27407 (N_27407,N_25490,N_26248);
or U27408 (N_27408,N_25962,N_25667);
or U27409 (N_27409,N_26201,N_25570);
nand U27410 (N_27410,N_25807,N_25296);
nand U27411 (N_27411,N_26388,N_25535);
or U27412 (N_27412,N_25277,N_26054);
xnor U27413 (N_27413,N_25200,N_26269);
nand U27414 (N_27414,N_25738,N_25866);
nand U27415 (N_27415,N_25308,N_26057);
and U27416 (N_27416,N_26193,N_25578);
or U27417 (N_27417,N_26218,N_25523);
nand U27418 (N_27418,N_26079,N_25471);
xor U27419 (N_27419,N_25417,N_25920);
and U27420 (N_27420,N_26097,N_26169);
nand U27421 (N_27421,N_26096,N_26367);
and U27422 (N_27422,N_25945,N_25494);
nor U27423 (N_27423,N_25752,N_25781);
nand U27424 (N_27424,N_25530,N_25741);
or U27425 (N_27425,N_25868,N_26140);
nor U27426 (N_27426,N_25297,N_25525);
xor U27427 (N_27427,N_25686,N_25876);
xor U27428 (N_27428,N_25342,N_25498);
and U27429 (N_27429,N_25277,N_26232);
and U27430 (N_27430,N_25632,N_26397);
nand U27431 (N_27431,N_25305,N_25752);
or U27432 (N_27432,N_25711,N_26397);
xor U27433 (N_27433,N_25214,N_26247);
or U27434 (N_27434,N_26286,N_25303);
xor U27435 (N_27435,N_26158,N_25277);
and U27436 (N_27436,N_25852,N_26113);
nor U27437 (N_27437,N_25829,N_25536);
nor U27438 (N_27438,N_25650,N_25787);
nand U27439 (N_27439,N_25607,N_26319);
and U27440 (N_27440,N_26364,N_25448);
nand U27441 (N_27441,N_26398,N_26006);
nand U27442 (N_27442,N_25722,N_25669);
nand U27443 (N_27443,N_25758,N_25349);
xnor U27444 (N_27444,N_25279,N_25689);
nand U27445 (N_27445,N_26105,N_26039);
and U27446 (N_27446,N_26342,N_25471);
or U27447 (N_27447,N_25885,N_25652);
nor U27448 (N_27448,N_25555,N_25262);
and U27449 (N_27449,N_26196,N_25644);
xor U27450 (N_27450,N_25334,N_25567);
and U27451 (N_27451,N_25665,N_25727);
or U27452 (N_27452,N_25457,N_26087);
nor U27453 (N_27453,N_25306,N_26332);
nor U27454 (N_27454,N_25657,N_26288);
or U27455 (N_27455,N_25593,N_25801);
and U27456 (N_27456,N_25351,N_26389);
nand U27457 (N_27457,N_25986,N_25536);
or U27458 (N_27458,N_25207,N_26059);
and U27459 (N_27459,N_26068,N_26090);
and U27460 (N_27460,N_25756,N_26059);
and U27461 (N_27461,N_25791,N_25807);
or U27462 (N_27462,N_26304,N_25646);
or U27463 (N_27463,N_25821,N_26014);
and U27464 (N_27464,N_25857,N_25810);
xor U27465 (N_27465,N_26302,N_26157);
xor U27466 (N_27466,N_25824,N_25889);
xnor U27467 (N_27467,N_26348,N_26047);
nor U27468 (N_27468,N_25654,N_25653);
nor U27469 (N_27469,N_25384,N_25746);
xor U27470 (N_27470,N_26088,N_25494);
and U27471 (N_27471,N_25891,N_25385);
nand U27472 (N_27472,N_25746,N_26347);
nand U27473 (N_27473,N_26085,N_25794);
and U27474 (N_27474,N_26362,N_25907);
and U27475 (N_27475,N_25635,N_26368);
xnor U27476 (N_27476,N_25355,N_25991);
nor U27477 (N_27477,N_25727,N_25404);
xnor U27478 (N_27478,N_25710,N_25773);
or U27479 (N_27479,N_25204,N_25443);
xor U27480 (N_27480,N_25369,N_25523);
nand U27481 (N_27481,N_25241,N_25221);
nor U27482 (N_27482,N_25999,N_26238);
nand U27483 (N_27483,N_26328,N_25509);
xor U27484 (N_27484,N_26243,N_25491);
nand U27485 (N_27485,N_26393,N_25705);
nor U27486 (N_27486,N_25472,N_26381);
nor U27487 (N_27487,N_25369,N_25912);
nor U27488 (N_27488,N_25365,N_25684);
and U27489 (N_27489,N_25368,N_25873);
nand U27490 (N_27490,N_26044,N_26222);
or U27491 (N_27491,N_25305,N_25526);
nor U27492 (N_27492,N_26262,N_25212);
xor U27493 (N_27493,N_26391,N_26104);
nand U27494 (N_27494,N_25441,N_26201);
or U27495 (N_27495,N_25969,N_25998);
and U27496 (N_27496,N_25313,N_26358);
xor U27497 (N_27497,N_25567,N_26159);
nand U27498 (N_27498,N_25593,N_25857);
nor U27499 (N_27499,N_26296,N_25540);
xnor U27500 (N_27500,N_25580,N_25596);
nand U27501 (N_27501,N_25409,N_25720);
nor U27502 (N_27502,N_26157,N_26309);
or U27503 (N_27503,N_25380,N_25962);
nor U27504 (N_27504,N_25378,N_26211);
nand U27505 (N_27505,N_25708,N_25983);
or U27506 (N_27506,N_25236,N_26123);
and U27507 (N_27507,N_25819,N_26199);
xor U27508 (N_27508,N_25214,N_25845);
or U27509 (N_27509,N_25318,N_25719);
nand U27510 (N_27510,N_25333,N_25649);
and U27511 (N_27511,N_25300,N_25447);
and U27512 (N_27512,N_26143,N_26365);
and U27513 (N_27513,N_25481,N_26198);
or U27514 (N_27514,N_26160,N_25601);
nand U27515 (N_27515,N_26225,N_25598);
nor U27516 (N_27516,N_26273,N_25328);
and U27517 (N_27517,N_26380,N_25995);
xnor U27518 (N_27518,N_25284,N_26173);
xor U27519 (N_27519,N_26179,N_25938);
nand U27520 (N_27520,N_25220,N_25519);
nand U27521 (N_27521,N_25838,N_26304);
nor U27522 (N_27522,N_26001,N_25732);
nand U27523 (N_27523,N_25797,N_26189);
or U27524 (N_27524,N_26200,N_26049);
xor U27525 (N_27525,N_26095,N_25415);
and U27526 (N_27526,N_26002,N_25476);
and U27527 (N_27527,N_25243,N_25934);
and U27528 (N_27528,N_25899,N_26262);
xnor U27529 (N_27529,N_25860,N_25447);
and U27530 (N_27530,N_26293,N_26038);
and U27531 (N_27531,N_26396,N_26074);
xor U27532 (N_27532,N_25946,N_25685);
and U27533 (N_27533,N_25525,N_25301);
nor U27534 (N_27534,N_25942,N_26292);
nand U27535 (N_27535,N_26052,N_26356);
nor U27536 (N_27536,N_25935,N_26331);
nand U27537 (N_27537,N_25310,N_26113);
and U27538 (N_27538,N_26175,N_25231);
nand U27539 (N_27539,N_25757,N_25733);
and U27540 (N_27540,N_25239,N_25799);
nand U27541 (N_27541,N_25319,N_25630);
xnor U27542 (N_27542,N_26066,N_26061);
and U27543 (N_27543,N_25433,N_25711);
or U27544 (N_27544,N_25235,N_26258);
xnor U27545 (N_27545,N_25445,N_26094);
xnor U27546 (N_27546,N_26195,N_25219);
or U27547 (N_27547,N_26283,N_25420);
xor U27548 (N_27548,N_26226,N_25626);
or U27549 (N_27549,N_25541,N_25574);
nand U27550 (N_27550,N_26086,N_25437);
nand U27551 (N_27551,N_25599,N_26130);
xor U27552 (N_27552,N_25470,N_25323);
nor U27553 (N_27553,N_26312,N_25854);
nand U27554 (N_27554,N_25627,N_26062);
or U27555 (N_27555,N_26391,N_25331);
xnor U27556 (N_27556,N_26228,N_25892);
or U27557 (N_27557,N_25416,N_25685);
nor U27558 (N_27558,N_25363,N_25566);
nor U27559 (N_27559,N_26079,N_26139);
nor U27560 (N_27560,N_25568,N_25735);
xnor U27561 (N_27561,N_25850,N_25785);
or U27562 (N_27562,N_25872,N_25679);
nor U27563 (N_27563,N_25670,N_25578);
nand U27564 (N_27564,N_26139,N_26390);
nand U27565 (N_27565,N_25506,N_26073);
or U27566 (N_27566,N_25583,N_25889);
or U27567 (N_27567,N_25781,N_25502);
and U27568 (N_27568,N_25785,N_25627);
or U27569 (N_27569,N_26068,N_25504);
or U27570 (N_27570,N_25473,N_25529);
or U27571 (N_27571,N_25422,N_26154);
nand U27572 (N_27572,N_25648,N_25264);
or U27573 (N_27573,N_25751,N_26061);
xnor U27574 (N_27574,N_25728,N_25355);
and U27575 (N_27575,N_25536,N_25641);
or U27576 (N_27576,N_25429,N_25863);
xor U27577 (N_27577,N_25773,N_26219);
nand U27578 (N_27578,N_25915,N_25413);
or U27579 (N_27579,N_26146,N_25959);
nand U27580 (N_27580,N_25543,N_25365);
nor U27581 (N_27581,N_25614,N_25861);
and U27582 (N_27582,N_25941,N_25266);
and U27583 (N_27583,N_25281,N_25509);
nand U27584 (N_27584,N_25744,N_26142);
nor U27585 (N_27585,N_25905,N_26253);
xnor U27586 (N_27586,N_25619,N_25562);
nor U27587 (N_27587,N_25904,N_25216);
and U27588 (N_27588,N_25743,N_25749);
or U27589 (N_27589,N_25604,N_26214);
nor U27590 (N_27590,N_25918,N_25793);
xnor U27591 (N_27591,N_26174,N_25998);
nand U27592 (N_27592,N_25652,N_25697);
and U27593 (N_27593,N_25769,N_25957);
and U27594 (N_27594,N_25445,N_26018);
or U27595 (N_27595,N_25210,N_25756);
and U27596 (N_27596,N_26026,N_25402);
and U27597 (N_27597,N_25882,N_26055);
and U27598 (N_27598,N_25922,N_25316);
and U27599 (N_27599,N_26040,N_25226);
and U27600 (N_27600,N_27169,N_27473);
nand U27601 (N_27601,N_26561,N_27131);
nor U27602 (N_27602,N_27234,N_27322);
nand U27603 (N_27603,N_26755,N_27578);
nor U27604 (N_27604,N_26441,N_26552);
and U27605 (N_27605,N_26558,N_26538);
nand U27606 (N_27606,N_27583,N_27317);
or U27607 (N_27607,N_26432,N_26532);
xor U27608 (N_27608,N_27468,N_26696);
or U27609 (N_27609,N_26550,N_26946);
nand U27610 (N_27610,N_26433,N_26999);
nor U27611 (N_27611,N_27487,N_27018);
or U27612 (N_27612,N_27100,N_27107);
nor U27613 (N_27613,N_26882,N_26542);
or U27614 (N_27614,N_27055,N_27428);
xor U27615 (N_27615,N_27476,N_26661);
or U27616 (N_27616,N_27188,N_26651);
and U27617 (N_27617,N_26994,N_26872);
nand U27618 (N_27618,N_27464,N_27365);
nand U27619 (N_27619,N_27060,N_27096);
nand U27620 (N_27620,N_26940,N_26977);
and U27621 (N_27621,N_27565,N_27435);
xnor U27622 (N_27622,N_26916,N_27210);
nand U27623 (N_27623,N_26417,N_27048);
nand U27624 (N_27624,N_26584,N_26492);
nand U27625 (N_27625,N_26511,N_26683);
or U27626 (N_27626,N_27184,N_27352);
nor U27627 (N_27627,N_26470,N_27488);
xnor U27628 (N_27628,N_27074,N_27548);
xor U27629 (N_27629,N_26408,N_27293);
or U27630 (N_27630,N_27148,N_26873);
nor U27631 (N_27631,N_26857,N_27196);
or U27632 (N_27632,N_27389,N_27008);
nand U27633 (N_27633,N_26845,N_27002);
or U27634 (N_27634,N_26874,N_27553);
xor U27635 (N_27635,N_27089,N_26896);
nand U27636 (N_27636,N_27495,N_26621);
and U27637 (N_27637,N_27297,N_27400);
and U27638 (N_27638,N_27153,N_26768);
and U27639 (N_27639,N_27178,N_26478);
or U27640 (N_27640,N_26497,N_26700);
nor U27641 (N_27641,N_26838,N_27031);
xnor U27642 (N_27642,N_27205,N_27462);
nand U27643 (N_27643,N_27315,N_27544);
or U27644 (N_27644,N_27115,N_27432);
or U27645 (N_27645,N_27429,N_27512);
or U27646 (N_27646,N_26949,N_26580);
xor U27647 (N_27647,N_27445,N_26843);
and U27648 (N_27648,N_26713,N_26719);
nor U27649 (N_27649,N_26596,N_27149);
or U27650 (N_27650,N_26503,N_27095);
xor U27651 (N_27651,N_26615,N_26565);
nor U27652 (N_27652,N_27254,N_26603);
and U27653 (N_27653,N_27189,N_27146);
nor U27654 (N_27654,N_27434,N_27246);
and U27655 (N_27655,N_27356,N_27391);
and U27656 (N_27656,N_26498,N_26460);
nand U27657 (N_27657,N_26834,N_26657);
or U27658 (N_27658,N_27067,N_27291);
and U27659 (N_27659,N_26490,N_26436);
nand U27660 (N_27660,N_26588,N_27374);
and U27661 (N_27661,N_26599,N_26846);
nand U27662 (N_27662,N_27326,N_26763);
and U27663 (N_27663,N_26793,N_26427);
xnor U27664 (N_27664,N_27073,N_27342);
nand U27665 (N_27665,N_27243,N_26413);
nor U27666 (N_27666,N_26777,N_26812);
or U27667 (N_27667,N_26508,N_26664);
and U27668 (N_27668,N_27005,N_27227);
and U27669 (N_27669,N_27394,N_27537);
and U27670 (N_27670,N_26677,N_26574);
nor U27671 (N_27671,N_27047,N_27579);
xor U27672 (N_27672,N_27284,N_26626);
nor U27673 (N_27673,N_27397,N_26414);
nand U27674 (N_27674,N_27581,N_27217);
nand U27675 (N_27675,N_27013,N_26566);
xnor U27676 (N_27676,N_26480,N_27329);
nor U27677 (N_27677,N_27318,N_26516);
nand U27678 (N_27678,N_27170,N_26948);
xor U27679 (N_27679,N_26646,N_26644);
or U27680 (N_27680,N_26469,N_27511);
nand U27681 (N_27681,N_26530,N_27162);
xnor U27682 (N_27682,N_26461,N_27139);
nor U27683 (N_27683,N_26544,N_27088);
and U27684 (N_27684,N_27395,N_26681);
and U27685 (N_27685,N_26870,N_27305);
nor U27686 (N_27686,N_27050,N_27549);
nand U27687 (N_27687,N_26638,N_26903);
xnor U27688 (N_27688,N_27026,N_26613);
nor U27689 (N_27689,N_27304,N_26703);
xnor U27690 (N_27690,N_27515,N_27194);
nand U27691 (N_27691,N_27382,N_26444);
nand U27692 (N_27692,N_27150,N_27152);
or U27693 (N_27693,N_26745,N_26947);
nor U27694 (N_27694,N_26850,N_27599);
and U27695 (N_27695,N_26964,N_26546);
nand U27696 (N_27696,N_26496,N_27235);
nor U27697 (N_27697,N_27399,N_26835);
xnor U27698 (N_27698,N_26955,N_27283);
or U27699 (N_27699,N_26652,N_26821);
nor U27700 (N_27700,N_26760,N_27257);
nor U27701 (N_27701,N_26918,N_26617);
nand U27702 (N_27702,N_26888,N_26879);
nand U27703 (N_27703,N_26930,N_27481);
xnor U27704 (N_27704,N_26649,N_27555);
xnor U27705 (N_27705,N_27396,N_26869);
or U27706 (N_27706,N_27522,N_27489);
nand U27707 (N_27707,N_26634,N_26686);
or U27708 (N_27708,N_26409,N_26782);
or U27709 (N_27709,N_27255,N_27423);
and U27710 (N_27710,N_26911,N_26709);
or U27711 (N_27711,N_26883,N_26775);
nor U27712 (N_27712,N_26692,N_26894);
and U27713 (N_27713,N_26820,N_26688);
and U27714 (N_27714,N_27054,N_26773);
nor U27715 (N_27715,N_26829,N_27193);
and U27716 (N_27716,N_26961,N_26789);
and U27717 (N_27717,N_26774,N_27556);
and U27718 (N_27718,N_27427,N_27408);
nor U27719 (N_27719,N_27559,N_26984);
and U27720 (N_27720,N_27083,N_27064);
xnor U27721 (N_27721,N_27500,N_26972);
nand U27722 (N_27722,N_26989,N_27388);
and U27723 (N_27723,N_26886,N_26998);
or U27724 (N_27724,N_26722,N_27024);
xnor U27725 (N_27725,N_27593,N_26906);
and U27726 (N_27726,N_27053,N_26919);
nand U27727 (N_27727,N_27081,N_27454);
xnor U27728 (N_27728,N_27068,N_26996);
nand U27729 (N_27729,N_27531,N_26744);
or U27730 (N_27730,N_26437,N_27174);
and U27731 (N_27731,N_27456,N_27425);
nor U27732 (N_27732,N_27300,N_27136);
and U27733 (N_27733,N_26974,N_27204);
xnor U27734 (N_27734,N_27233,N_26482);
and U27735 (N_27735,N_27044,N_27350);
nand U27736 (N_27736,N_26485,N_26855);
or U27737 (N_27737,N_27279,N_26985);
nand U27738 (N_27738,N_26741,N_26702);
or U27739 (N_27739,N_27239,N_26951);
and U27740 (N_27740,N_27087,N_27041);
and U27741 (N_27741,N_27258,N_27175);
xnor U27742 (N_27742,N_26628,N_27465);
and U27743 (N_27743,N_26594,N_26770);
nand U27744 (N_27744,N_27539,N_27290);
or U27745 (N_27745,N_27527,N_26660);
or U27746 (N_27746,N_26993,N_27373);
or U27747 (N_27747,N_26553,N_26711);
or U27748 (N_27748,N_26808,N_27316);
nor U27749 (N_27749,N_27085,N_26509);
and U27750 (N_27750,N_26578,N_27142);
nor U27751 (N_27751,N_27173,N_26786);
or U27752 (N_27752,N_26790,N_27192);
or U27753 (N_27753,N_26904,N_26841);
nor U27754 (N_27754,N_26738,N_27438);
xor U27755 (N_27755,N_26592,N_26945);
and U27756 (N_27756,N_27528,N_26758);
or U27757 (N_27757,N_27514,N_27541);
or U27758 (N_27758,N_26818,N_27477);
nand U27759 (N_27759,N_27001,N_26495);
nor U27760 (N_27760,N_27348,N_26524);
nor U27761 (N_27761,N_26701,N_27166);
nand U27762 (N_27762,N_27209,N_27224);
and U27763 (N_27763,N_26699,N_26784);
or U27764 (N_27764,N_27450,N_26783);
or U27765 (N_27765,N_27075,N_26670);
nand U27766 (N_27766,N_27575,N_27530);
nand U27767 (N_27767,N_27057,N_27406);
xor U27768 (N_27768,N_26969,N_26513);
nor U27769 (N_27769,N_27120,N_27498);
or U27770 (N_27770,N_26965,N_26865);
xnor U27771 (N_27771,N_27510,N_26848);
nand U27772 (N_27772,N_26415,N_27598);
and U27773 (N_27773,N_26863,N_27499);
nor U27774 (N_27774,N_26800,N_26929);
nand U27775 (N_27775,N_26765,N_26840);
xor U27776 (N_27776,N_26551,N_27179);
or U27777 (N_27777,N_27289,N_26605);
nand U27778 (N_27778,N_27281,N_26693);
or U27779 (N_27779,N_26725,N_26942);
and U27780 (N_27780,N_26801,N_26598);
or U27781 (N_27781,N_26915,N_26844);
nand U27782 (N_27782,N_26604,N_26512);
nand U27783 (N_27783,N_26807,N_27584);
xnor U27784 (N_27784,N_26875,N_26867);
and U27785 (N_27785,N_26860,N_26514);
xnor U27786 (N_27786,N_27410,N_26987);
nor U27787 (N_27787,N_27138,N_26575);
nand U27788 (N_27788,N_26629,N_26849);
nand U27789 (N_27789,N_26953,N_27165);
nor U27790 (N_27790,N_26715,N_27051);
and U27791 (N_27791,N_27383,N_27122);
xor U27792 (N_27792,N_26522,N_26486);
or U27793 (N_27793,N_27301,N_27480);
and U27794 (N_27794,N_27197,N_26827);
and U27795 (N_27795,N_26406,N_26619);
nand U27796 (N_27796,N_27216,N_27469);
or U27797 (N_27797,N_27437,N_26650);
or U27798 (N_27798,N_26891,N_27546);
or U27799 (N_27799,N_26721,N_26412);
and U27800 (N_27800,N_26585,N_26749);
and U27801 (N_27801,N_26536,N_26407);
or U27802 (N_27802,N_27452,N_26724);
xor U27803 (N_27803,N_26442,N_27478);
xor U27804 (N_27804,N_26577,N_26813);
nor U27805 (N_27805,N_27533,N_27124);
xnor U27806 (N_27806,N_26854,N_27474);
xor U27807 (N_27807,N_26796,N_26581);
nor U27808 (N_27808,N_27167,N_27133);
and U27809 (N_27809,N_27127,N_27347);
xnor U27810 (N_27810,N_26554,N_26501);
or U27811 (N_27811,N_26739,N_27463);
xor U27812 (N_27812,N_27341,N_26515);
or U27813 (N_27813,N_27418,N_27069);
or U27814 (N_27814,N_27004,N_27278);
nor U27815 (N_27815,N_26909,N_26457);
xnor U27816 (N_27816,N_26440,N_26979);
or U27817 (N_27817,N_27415,N_27385);
xnor U27818 (N_27818,N_26549,N_27339);
nor U27819 (N_27819,N_27595,N_27331);
xnor U27820 (N_27820,N_27103,N_26928);
nand U27821 (N_27821,N_26426,N_27168);
and U27822 (N_27822,N_26571,N_27245);
and U27823 (N_27823,N_26557,N_27422);
nand U27824 (N_27824,N_26640,N_27486);
xor U27825 (N_27825,N_27158,N_27379);
and U27826 (N_27826,N_26729,N_26662);
nor U27827 (N_27827,N_27307,N_27591);
or U27828 (N_27828,N_27276,N_26932);
nand U27829 (N_27829,N_27490,N_26454);
and U27830 (N_27830,N_27020,N_26676);
nand U27831 (N_27831,N_26809,N_27125);
or U27832 (N_27832,N_27517,N_27572);
or U27833 (N_27833,N_27111,N_26806);
and U27834 (N_27834,N_27263,N_26714);
xnor U27835 (N_27835,N_26448,N_26614);
and U27836 (N_27836,N_27470,N_27264);
xor U27837 (N_27837,N_27377,N_27065);
and U27838 (N_27838,N_27409,N_27232);
or U27839 (N_27839,N_26502,N_27497);
xnor U27840 (N_27840,N_27560,N_26505);
and U27841 (N_27841,N_27154,N_27424);
nand U27842 (N_27842,N_27414,N_27349);
and U27843 (N_27843,N_27229,N_26569);
xnor U27844 (N_27844,N_27206,N_27298);
xnor U27845 (N_27845,N_26787,N_26525);
and U27846 (N_27846,N_27187,N_26752);
or U27847 (N_27847,N_27567,N_27505);
or U27848 (N_27848,N_27368,N_26772);
nand U27849 (N_27849,N_26941,N_26420);
and U27850 (N_27850,N_26506,N_27504);
nor U27851 (N_27851,N_26507,N_27426);
xor U27852 (N_27852,N_27538,N_26885);
xor U27853 (N_27853,N_26901,N_27061);
or U27854 (N_27854,N_27401,N_27145);
nand U27855 (N_27855,N_27453,N_26567);
or U27856 (N_27856,N_27569,N_27431);
xnor U27857 (N_27857,N_27355,N_26656);
nor U27858 (N_27858,N_26517,N_27485);
and U27859 (N_27859,N_26622,N_26762);
or U27860 (N_27860,N_26535,N_26658);
nor U27861 (N_27861,N_26451,N_27092);
or U27862 (N_27862,N_27540,N_26707);
nor U27863 (N_27863,N_27015,N_27256);
nor U27864 (N_27864,N_27525,N_26632);
nor U27865 (N_27865,N_27413,N_26421);
nor U27866 (N_27866,N_26689,N_26543);
or U27867 (N_27867,N_26952,N_27526);
nor U27868 (N_27868,N_27220,N_27439);
nor U27869 (N_27869,N_27340,N_27303);
nor U27870 (N_27870,N_26842,N_27455);
xor U27871 (N_27871,N_27286,N_27573);
or U27872 (N_27872,N_27249,N_26685);
xor U27873 (N_27873,N_26464,N_26913);
and U27874 (N_27874,N_26935,N_26499);
xnor U27875 (N_27875,N_27277,N_27117);
xnor U27876 (N_27876,N_27223,N_26611);
xor U27877 (N_27877,N_27010,N_27324);
nand U27878 (N_27878,N_26810,N_26589);
nand U27879 (N_27879,N_26859,N_27346);
xnor U27880 (N_27880,N_27585,N_26852);
xor U27881 (N_27881,N_26927,N_27237);
and U27882 (N_27882,N_27457,N_27271);
nand U27883 (N_27883,N_26912,N_26489);
or U27884 (N_27884,N_27101,N_27518);
or U27885 (N_27885,N_26582,N_27274);
and U27886 (N_27886,N_26527,N_26630);
or U27887 (N_27887,N_27272,N_27180);
xor U27888 (N_27888,N_27513,N_27144);
and U27889 (N_27889,N_26892,N_26862);
and U27890 (N_27890,N_26443,N_27359);
xor U27891 (N_27891,N_27507,N_27362);
and U27892 (N_27892,N_27587,N_26923);
nand U27893 (N_27893,N_26736,N_26449);
nor U27894 (N_27894,N_27268,N_27104);
and U27895 (N_27895,N_27135,N_27059);
nand U27896 (N_27896,N_26743,N_27156);
or U27897 (N_27897,N_26612,N_26430);
xor U27898 (N_27898,N_27536,N_26471);
nor U27899 (N_27899,N_26794,N_26423);
and U27900 (N_27900,N_26521,N_27444);
nand U27901 (N_27901,N_27151,N_27099);
and U27902 (N_27902,N_27482,N_27366);
xnor U27903 (N_27903,N_27370,N_27308);
xnor U27904 (N_27904,N_26541,N_26731);
and U27905 (N_27905,N_26742,N_26769);
and U27906 (N_27906,N_26697,N_26908);
or U27907 (N_27907,N_27551,N_26944);
xor U27908 (N_27908,N_27267,N_27292);
and U27909 (N_27909,N_27282,N_27046);
or U27910 (N_27910,N_26753,N_26483);
or U27911 (N_27911,N_27022,N_27491);
nand U27912 (N_27912,N_26730,N_27521);
xor U27913 (N_27913,N_26897,N_27171);
nor U27914 (N_27914,N_26601,N_27492);
nand U27915 (N_27915,N_27344,N_27405);
or U27916 (N_27916,N_27387,N_27320);
nor U27917 (N_27917,N_27484,N_26833);
nor U27918 (N_27918,N_26695,N_27404);
nand U27919 (N_27919,N_27098,N_27345);
nand U27920 (N_27920,N_26917,N_26710);
or U27921 (N_27921,N_26455,N_27000);
nand U27922 (N_27922,N_27384,N_27381);
xor U27923 (N_27923,N_26520,N_26708);
and U27924 (N_27924,N_27147,N_27052);
or U27925 (N_27925,N_27269,N_26439);
nor U27926 (N_27926,N_27161,N_27011);
nor U27927 (N_27927,N_26537,N_26559);
xor U27928 (N_27928,N_26826,N_26799);
xor U27929 (N_27929,N_27200,N_26816);
xor U27930 (N_27930,N_27181,N_27260);
nand U27931 (N_27931,N_27328,N_27443);
nand U27932 (N_27932,N_26518,N_27248);
nor U27933 (N_27933,N_27312,N_27412);
nand U27934 (N_27934,N_27006,N_26411);
or U27935 (N_27935,N_26548,N_26531);
or U27936 (N_27936,N_26756,N_26720);
xor U27937 (N_27937,N_27313,N_27529);
nor U27938 (N_27938,N_26832,N_26402);
nand U27939 (N_27939,N_26572,N_26428);
or U27940 (N_27940,N_27577,N_26616);
or U27941 (N_27941,N_27212,N_27371);
nand U27942 (N_27942,N_26805,N_27072);
xnor U27943 (N_27943,N_26960,N_27336);
or U27944 (N_27944,N_26494,N_26705);
nor U27945 (N_27945,N_27333,N_26950);
xnor U27946 (N_27946,N_26479,N_26597);
nand U27947 (N_27947,N_27545,N_26804);
and U27948 (N_27948,N_27358,N_26624);
or U27949 (N_27949,N_27208,N_27532);
or U27950 (N_27950,N_26583,N_26864);
nor U27951 (N_27951,N_27523,N_27078);
xor U27952 (N_27952,N_26510,N_27494);
nor U27953 (N_27953,N_27032,N_27369);
and U27954 (N_27954,N_27203,N_26447);
nor U27955 (N_27955,N_26422,N_26654);
xnor U27956 (N_27956,N_27112,N_26938);
nand U27957 (N_27957,N_26450,N_26887);
and U27958 (N_27958,N_26956,N_26878);
and U27959 (N_27959,N_27009,N_27442);
and U27960 (N_27960,N_26687,N_27108);
xnor U27961 (N_27961,N_27590,N_26665);
nor U27962 (N_27962,N_26853,N_26416);
nand U27963 (N_27963,N_26839,N_27119);
nand U27964 (N_27964,N_27177,N_27580);
nand U27965 (N_27965,N_27576,N_26452);
or U27966 (N_27966,N_27325,N_26602);
and U27967 (N_27967,N_26750,N_26748);
nor U27968 (N_27968,N_26943,N_26682);
nor U27969 (N_27969,N_27123,N_27589);
or U27970 (N_27970,N_27080,N_26523);
xnor U27971 (N_27971,N_27091,N_26746);
or U27972 (N_27972,N_26610,N_27077);
and U27973 (N_27973,N_27376,N_27028);
nand U27974 (N_27974,N_27393,N_27299);
nand U27975 (N_27975,N_27129,N_27343);
nor U27976 (N_27976,N_26905,N_26671);
xor U27977 (N_27977,N_27519,N_27386);
nor U27978 (N_27978,N_26732,N_26933);
or U27979 (N_27979,N_26727,N_27471);
nor U27980 (N_27980,N_26830,N_26642);
xnor U27981 (N_27981,N_27594,N_26576);
nand U27982 (N_27982,N_27155,N_27163);
xnor U27983 (N_27983,N_27126,N_26868);
and U27984 (N_27984,N_27109,N_27114);
nor U27985 (N_27985,N_27524,N_27066);
nor U27986 (N_27986,N_26716,N_26636);
or U27987 (N_27987,N_27570,N_27475);
or U27988 (N_27988,N_26895,N_26831);
or U27989 (N_27989,N_27084,N_27357);
nand U27990 (N_27990,N_27520,N_27242);
xor U27991 (N_27991,N_27458,N_27140);
and U27992 (N_27992,N_26545,N_27398);
xnor U27993 (N_27993,N_26771,N_26500);
or U27994 (N_27994,N_27390,N_26971);
nor U27995 (N_27995,N_26757,N_27071);
nand U27996 (N_27996,N_27294,N_27199);
nor U27997 (N_27997,N_26988,N_27319);
xnor U27998 (N_27998,N_26620,N_27436);
or U27999 (N_27999,N_27063,N_26898);
or U28000 (N_28000,N_27007,N_26690);
nor U28001 (N_28001,N_26925,N_27550);
nand U28002 (N_28002,N_26811,N_26675);
and U28003 (N_28003,N_27222,N_27118);
nor U28004 (N_28004,N_26963,N_27261);
nand U28005 (N_28005,N_27157,N_26893);
or U28006 (N_28006,N_26476,N_26992);
xnor U28007 (N_28007,N_27448,N_27561);
nor U28008 (N_28008,N_27097,N_27190);
and U28009 (N_28009,N_27247,N_27016);
or U28010 (N_28010,N_27266,N_26631);
and U28011 (N_28011,N_26803,N_26679);
nand U28012 (N_28012,N_26600,N_26639);
nor U28013 (N_28013,N_26717,N_26973);
nand U28014 (N_28014,N_26907,N_26410);
and U28015 (N_28015,N_27558,N_26990);
and U28016 (N_28016,N_26997,N_26627);
nor U28017 (N_28017,N_27003,N_26766);
nor U28018 (N_28018,N_27211,N_26698);
nor U28019 (N_28019,N_27449,N_27288);
xor U28020 (N_28020,N_27421,N_27265);
nand U28021 (N_28021,N_27262,N_26900);
xnor U28022 (N_28022,N_27037,N_27023);
nand U28023 (N_28023,N_26824,N_26740);
nor U28024 (N_28024,N_26761,N_26435);
xor U28025 (N_28025,N_27040,N_26563);
xnor U28026 (N_28026,N_27547,N_27094);
xnor U28027 (N_28027,N_27207,N_27106);
or U28028 (N_28028,N_26814,N_27451);
or U28029 (N_28029,N_26400,N_26890);
and U28030 (N_28030,N_27296,N_26466);
and U28031 (N_28031,N_26481,N_26637);
and U28032 (N_28032,N_27597,N_27502);
nand U28033 (N_28033,N_26962,N_26529);
or U28034 (N_28034,N_26534,N_26866);
nand U28035 (N_28035,N_27093,N_27564);
xor U28036 (N_28036,N_27172,N_27466);
or U28037 (N_28037,N_27407,N_27186);
xnor U28038 (N_28038,N_26718,N_27433);
xnor U28039 (N_28039,N_26607,N_27542);
and U28040 (N_28040,N_26791,N_26815);
or U28041 (N_28041,N_27554,N_27353);
xor U28042 (N_28042,N_27334,N_26593);
or U28043 (N_28043,N_27230,N_26822);
nor U28044 (N_28044,N_27259,N_26767);
nand U28045 (N_28045,N_27082,N_26877);
or U28046 (N_28046,N_26934,N_27164);
nor U28047 (N_28047,N_27049,N_26780);
nor U28048 (N_28048,N_26493,N_27375);
and U28049 (N_28049,N_26587,N_27360);
nor U28050 (N_28050,N_27116,N_27461);
and U28051 (N_28051,N_27250,N_26474);
nor U28052 (N_28052,N_27191,N_26954);
nand U28053 (N_28053,N_26666,N_27440);
nand U28054 (N_28054,N_26609,N_26463);
nand U28055 (N_28055,N_26591,N_27185);
nor U28056 (N_28056,N_26881,N_27506);
nor U28057 (N_28057,N_26728,N_26528);
xnor U28058 (N_28058,N_26425,N_26568);
and U28059 (N_28059,N_27218,N_27159);
and U28060 (N_28060,N_26733,N_26655);
and U28061 (N_28061,N_27563,N_26737);
nand U28062 (N_28062,N_27105,N_26547);
nor U28063 (N_28063,N_27574,N_27496);
nor U28064 (N_28064,N_26484,N_26723);
nand U28065 (N_28065,N_27330,N_27090);
nand U28066 (N_28066,N_26876,N_27035);
nand U28067 (N_28067,N_26462,N_26764);
and U28068 (N_28068,N_26668,N_26459);
and U28069 (N_28069,N_26817,N_27535);
nand U28070 (N_28070,N_26920,N_26936);
nor U28071 (N_28071,N_26976,N_27483);
nand U28072 (N_28072,N_27302,N_26473);
and U28073 (N_28073,N_27586,N_26564);
xnor U28074 (N_28074,N_27056,N_27420);
and U28075 (N_28075,N_26641,N_26788);
nand U28076 (N_28076,N_27568,N_26431);
nand U28077 (N_28077,N_27493,N_26526);
nor U28078 (N_28078,N_27447,N_26623);
xnor U28079 (N_28079,N_27417,N_26643);
xor U28080 (N_28080,N_26798,N_27034);
or U28081 (N_28081,N_27198,N_26959);
nand U28082 (N_28082,N_26982,N_26590);
and U28083 (N_28083,N_27273,N_27596);
nand U28084 (N_28084,N_26467,N_26751);
nand U28085 (N_28085,N_27446,N_26403);
nand U28086 (N_28086,N_26663,N_26776);
xor U28087 (N_28087,N_26851,N_27311);
or U28088 (N_28088,N_26975,N_27592);
or U28089 (N_28089,N_27351,N_26735);
xnor U28090 (N_28090,N_26570,N_26968);
xor U28091 (N_28091,N_27176,N_27562);
nor U28092 (N_28092,N_27557,N_27309);
and U28093 (N_28093,N_27402,N_27042);
and U28094 (N_28094,N_26465,N_26635);
xnor U28095 (N_28095,N_27086,N_26924);
nor U28096 (N_28096,N_26606,N_26475);
nor U28097 (N_28097,N_26704,N_27025);
nor U28098 (N_28098,N_26673,N_26647);
xor U28099 (N_28099,N_26659,N_27215);
nand U28100 (N_28100,N_26967,N_27030);
xor U28101 (N_28101,N_26684,N_26648);
nor U28102 (N_28102,N_27403,N_27231);
xnor U28103 (N_28103,N_26778,N_27552);
xor U28104 (N_28104,N_26653,N_27017);
nor U28105 (N_28105,N_26405,N_26983);
and U28106 (N_28106,N_26472,N_26836);
and U28107 (N_28107,N_27411,N_26401);
xnor U28108 (N_28108,N_27043,N_27582);
nor U28109 (N_28109,N_27058,N_26922);
xnor U28110 (N_28110,N_26734,N_27295);
nand U28111 (N_28111,N_26560,N_27503);
and U28112 (N_28112,N_27228,N_26539);
and U28113 (N_28113,N_27021,N_27076);
and U28114 (N_28114,N_26533,N_26889);
nor U28115 (N_28115,N_27225,N_27240);
nor U28116 (N_28116,N_26424,N_26595);
and U28117 (N_28117,N_26837,N_26823);
and U28118 (N_28118,N_27033,N_27110);
nand U28119 (N_28119,N_26446,N_26910);
nor U28120 (N_28120,N_27201,N_26966);
or U28121 (N_28121,N_27202,N_27285);
nand U28122 (N_28122,N_26504,N_26487);
nand U28123 (N_28123,N_27014,N_27226);
or U28124 (N_28124,N_27195,N_27363);
nor U28125 (N_28125,N_26556,N_26754);
nor U28126 (N_28126,N_27275,N_27141);
nand U28127 (N_28127,N_27029,N_27338);
nand U28128 (N_28128,N_26645,N_26795);
nor U28129 (N_28129,N_26555,N_27566);
and U28130 (N_28130,N_26981,N_26667);
nor U28131 (N_28131,N_27236,N_27102);
nor U28132 (N_28132,N_27430,N_27321);
nor U28133 (N_28133,N_26939,N_26453);
nor U28134 (N_28134,N_26871,N_26759);
xnor U28135 (N_28135,N_26706,N_27062);
nor U28136 (N_28136,N_27472,N_27354);
xnor U28137 (N_28137,N_27323,N_27214);
nor U28138 (N_28138,N_26858,N_27441);
nor U28139 (N_28139,N_27460,N_27508);
and U28140 (N_28140,N_27314,N_27253);
and U28141 (N_28141,N_26477,N_27244);
nand U28142 (N_28142,N_27335,N_27337);
and U28143 (N_28143,N_27310,N_26579);
nand U28144 (N_28144,N_26519,N_27182);
and U28145 (N_28145,N_26861,N_27038);
xnor U28146 (N_28146,N_26625,N_26995);
xor U28147 (N_28147,N_27270,N_27143);
xnor U28148 (N_28148,N_26779,N_26958);
or U28149 (N_28149,N_26691,N_27364);
and U28150 (N_28150,N_27213,N_27479);
nand U28151 (N_28151,N_27534,N_27130);
nand U28152 (N_28152,N_27012,N_27571);
and U28153 (N_28153,N_27392,N_27027);
nor U28154 (N_28154,N_27183,N_27036);
xor U28155 (N_28155,N_26672,N_26418);
and U28156 (N_28156,N_26438,N_27306);
or U28157 (N_28157,N_26847,N_27137);
xnor U28158 (N_28158,N_26468,N_26674);
xor U28159 (N_28159,N_27467,N_26902);
xnor U28160 (N_28160,N_27419,N_27516);
and U28161 (N_28161,N_26931,N_27113);
and U28162 (N_28162,N_26456,N_27287);
xor U28163 (N_28163,N_27252,N_26404);
or U28164 (N_28164,N_26921,N_26608);
and U28165 (N_28165,N_26445,N_26491);
nand U28166 (N_28166,N_27361,N_27380);
nand U28167 (N_28167,N_27134,N_26991);
and U28168 (N_28168,N_26488,N_27039);
xor U28169 (N_28169,N_26458,N_26434);
nand U28170 (N_28170,N_27121,N_26562);
nand U28171 (N_28171,N_26540,N_27332);
or U28172 (N_28172,N_26586,N_27543);
and U28173 (N_28173,N_26792,N_27280);
nand U28174 (N_28174,N_26747,N_27501);
or U28175 (N_28175,N_27327,N_27378);
nand U28176 (N_28176,N_26970,N_26781);
and U28177 (N_28177,N_26712,N_26899);
nor U28178 (N_28178,N_26937,N_27070);
nor U28179 (N_28179,N_27079,N_26694);
or U28180 (N_28180,N_27588,N_26633);
or U28181 (N_28181,N_26980,N_26819);
nor U28182 (N_28182,N_26986,N_26678);
nand U28183 (N_28183,N_27251,N_27221);
or U28184 (N_28184,N_27160,N_27367);
nor U28185 (N_28185,N_26884,N_26669);
nor U28186 (N_28186,N_26429,N_26914);
nor U28187 (N_28187,N_26802,N_26573);
or U28188 (N_28188,N_26726,N_26785);
or U28189 (N_28189,N_26880,N_26797);
nor U28190 (N_28190,N_26618,N_26856);
or U28191 (N_28191,N_27219,N_27045);
xor U28192 (N_28192,N_27459,N_27128);
xnor U28193 (N_28193,N_26828,N_26978);
and U28194 (N_28194,N_27238,N_27132);
and U28195 (N_28195,N_27509,N_27241);
nand U28196 (N_28196,N_27019,N_26825);
xor U28197 (N_28197,N_27372,N_26419);
xor U28198 (N_28198,N_26957,N_26680);
nor U28199 (N_28199,N_26926,N_27416);
xor U28200 (N_28200,N_26873,N_26692);
nor U28201 (N_28201,N_27047,N_26491);
and U28202 (N_28202,N_27018,N_27085);
nor U28203 (N_28203,N_26589,N_26627);
nand U28204 (N_28204,N_26428,N_27215);
nor U28205 (N_28205,N_27519,N_26950);
nor U28206 (N_28206,N_27159,N_26784);
nand U28207 (N_28207,N_27583,N_26900);
nand U28208 (N_28208,N_26668,N_27411);
xor U28209 (N_28209,N_26892,N_26675);
nor U28210 (N_28210,N_27448,N_26746);
nand U28211 (N_28211,N_27286,N_27415);
xnor U28212 (N_28212,N_27068,N_26527);
nand U28213 (N_28213,N_26896,N_27222);
and U28214 (N_28214,N_27584,N_26743);
nor U28215 (N_28215,N_27134,N_27251);
xor U28216 (N_28216,N_27125,N_27170);
or U28217 (N_28217,N_26525,N_26572);
nand U28218 (N_28218,N_26943,N_27486);
xor U28219 (N_28219,N_26549,N_26833);
nor U28220 (N_28220,N_26811,N_27250);
or U28221 (N_28221,N_26721,N_27140);
and U28222 (N_28222,N_26659,N_26883);
and U28223 (N_28223,N_27423,N_27299);
nor U28224 (N_28224,N_27034,N_27001);
nand U28225 (N_28225,N_26783,N_26791);
and U28226 (N_28226,N_27428,N_26701);
or U28227 (N_28227,N_27124,N_27232);
or U28228 (N_28228,N_26980,N_27483);
and U28229 (N_28229,N_26527,N_26810);
or U28230 (N_28230,N_27173,N_27542);
and U28231 (N_28231,N_27296,N_26527);
and U28232 (N_28232,N_27173,N_27452);
nand U28233 (N_28233,N_26881,N_27283);
nor U28234 (N_28234,N_27116,N_27589);
and U28235 (N_28235,N_27159,N_26773);
or U28236 (N_28236,N_27241,N_26585);
xnor U28237 (N_28237,N_27594,N_27010);
nand U28238 (N_28238,N_27291,N_27364);
nor U28239 (N_28239,N_26869,N_26831);
or U28240 (N_28240,N_26407,N_27044);
nand U28241 (N_28241,N_27037,N_27220);
nor U28242 (N_28242,N_27105,N_26534);
xnor U28243 (N_28243,N_26889,N_27405);
or U28244 (N_28244,N_26834,N_27448);
nor U28245 (N_28245,N_27019,N_27241);
xor U28246 (N_28246,N_26846,N_26536);
and U28247 (N_28247,N_26564,N_26732);
nor U28248 (N_28248,N_27409,N_26989);
nor U28249 (N_28249,N_27378,N_26521);
nand U28250 (N_28250,N_26565,N_27013);
nor U28251 (N_28251,N_26818,N_27079);
nand U28252 (N_28252,N_26722,N_26492);
or U28253 (N_28253,N_26839,N_27465);
xor U28254 (N_28254,N_27270,N_27421);
xnor U28255 (N_28255,N_26525,N_26524);
and U28256 (N_28256,N_27100,N_27324);
nand U28257 (N_28257,N_26706,N_26783);
and U28258 (N_28258,N_26880,N_27033);
xnor U28259 (N_28259,N_26812,N_26684);
xnor U28260 (N_28260,N_27064,N_26570);
and U28261 (N_28261,N_27454,N_27103);
or U28262 (N_28262,N_27376,N_26981);
and U28263 (N_28263,N_26982,N_27496);
and U28264 (N_28264,N_26549,N_27189);
xor U28265 (N_28265,N_26883,N_27043);
nor U28266 (N_28266,N_27004,N_27563);
nand U28267 (N_28267,N_26643,N_26503);
xor U28268 (N_28268,N_27592,N_27350);
nor U28269 (N_28269,N_26598,N_26933);
or U28270 (N_28270,N_26820,N_27196);
xor U28271 (N_28271,N_27274,N_26831);
nand U28272 (N_28272,N_27481,N_26429);
nand U28273 (N_28273,N_26783,N_27265);
and U28274 (N_28274,N_26418,N_26950);
nor U28275 (N_28275,N_27022,N_27527);
nand U28276 (N_28276,N_26991,N_26648);
nand U28277 (N_28277,N_26880,N_27144);
nor U28278 (N_28278,N_26774,N_26819);
nand U28279 (N_28279,N_27208,N_27051);
and U28280 (N_28280,N_27581,N_27483);
nand U28281 (N_28281,N_27096,N_27533);
or U28282 (N_28282,N_26801,N_26947);
xnor U28283 (N_28283,N_27200,N_26561);
nor U28284 (N_28284,N_26932,N_26643);
or U28285 (N_28285,N_26982,N_26598);
or U28286 (N_28286,N_27592,N_27189);
and U28287 (N_28287,N_27227,N_26488);
nor U28288 (N_28288,N_26742,N_27388);
nor U28289 (N_28289,N_27012,N_27559);
xor U28290 (N_28290,N_27032,N_26787);
and U28291 (N_28291,N_27482,N_26440);
nor U28292 (N_28292,N_27551,N_27545);
or U28293 (N_28293,N_27126,N_26671);
nand U28294 (N_28294,N_27274,N_26804);
xor U28295 (N_28295,N_26559,N_26671);
xnor U28296 (N_28296,N_26428,N_27361);
nor U28297 (N_28297,N_27262,N_26953);
nor U28298 (N_28298,N_26771,N_27313);
nor U28299 (N_28299,N_26492,N_26442);
xor U28300 (N_28300,N_26717,N_27529);
and U28301 (N_28301,N_26822,N_27287);
nor U28302 (N_28302,N_26620,N_27539);
nor U28303 (N_28303,N_27367,N_27303);
nand U28304 (N_28304,N_26691,N_26536);
and U28305 (N_28305,N_26428,N_26922);
and U28306 (N_28306,N_26406,N_27536);
and U28307 (N_28307,N_26635,N_27556);
or U28308 (N_28308,N_26531,N_26607);
or U28309 (N_28309,N_26943,N_26607);
xnor U28310 (N_28310,N_27200,N_27594);
nor U28311 (N_28311,N_26660,N_26984);
xnor U28312 (N_28312,N_27342,N_26552);
or U28313 (N_28313,N_27438,N_27373);
and U28314 (N_28314,N_27376,N_27430);
or U28315 (N_28315,N_26812,N_27261);
or U28316 (N_28316,N_27006,N_27365);
or U28317 (N_28317,N_26499,N_26954);
nand U28318 (N_28318,N_26975,N_26739);
or U28319 (N_28319,N_27099,N_26473);
nand U28320 (N_28320,N_26860,N_27149);
or U28321 (N_28321,N_27358,N_26923);
or U28322 (N_28322,N_26651,N_27029);
xnor U28323 (N_28323,N_27043,N_27542);
and U28324 (N_28324,N_27006,N_26694);
and U28325 (N_28325,N_26452,N_26841);
and U28326 (N_28326,N_26895,N_26750);
nand U28327 (N_28327,N_26765,N_26918);
nor U28328 (N_28328,N_27193,N_27429);
nand U28329 (N_28329,N_27189,N_26486);
xor U28330 (N_28330,N_26443,N_27471);
and U28331 (N_28331,N_26799,N_27502);
xnor U28332 (N_28332,N_26647,N_27047);
nand U28333 (N_28333,N_26582,N_27263);
and U28334 (N_28334,N_27305,N_27013);
nor U28335 (N_28335,N_26924,N_26913);
nor U28336 (N_28336,N_27322,N_27024);
or U28337 (N_28337,N_26499,N_27496);
or U28338 (N_28338,N_27168,N_27479);
nor U28339 (N_28339,N_26875,N_27049);
nand U28340 (N_28340,N_26484,N_26508);
xor U28341 (N_28341,N_27141,N_27353);
nand U28342 (N_28342,N_27509,N_26775);
and U28343 (N_28343,N_26888,N_27273);
and U28344 (N_28344,N_27360,N_27460);
nand U28345 (N_28345,N_27081,N_26649);
and U28346 (N_28346,N_27129,N_27426);
or U28347 (N_28347,N_27162,N_26570);
nand U28348 (N_28348,N_26634,N_26946);
xnor U28349 (N_28349,N_27259,N_27320);
or U28350 (N_28350,N_27548,N_26502);
and U28351 (N_28351,N_26635,N_26582);
xnor U28352 (N_28352,N_27399,N_27253);
xor U28353 (N_28353,N_27036,N_26507);
and U28354 (N_28354,N_26632,N_27560);
or U28355 (N_28355,N_26649,N_27322);
nand U28356 (N_28356,N_26722,N_27019);
nand U28357 (N_28357,N_27260,N_26479);
xnor U28358 (N_28358,N_27305,N_26788);
xnor U28359 (N_28359,N_26620,N_27430);
and U28360 (N_28360,N_26770,N_27317);
nor U28361 (N_28361,N_26542,N_26756);
xnor U28362 (N_28362,N_26589,N_27348);
and U28363 (N_28363,N_26562,N_27294);
nand U28364 (N_28364,N_27286,N_26777);
xnor U28365 (N_28365,N_27579,N_27359);
nand U28366 (N_28366,N_27495,N_27398);
nor U28367 (N_28367,N_27342,N_26415);
nor U28368 (N_28368,N_27137,N_27564);
nand U28369 (N_28369,N_27550,N_26624);
xnor U28370 (N_28370,N_27334,N_26595);
and U28371 (N_28371,N_27372,N_27433);
nor U28372 (N_28372,N_26742,N_26747);
nand U28373 (N_28373,N_27155,N_26512);
nor U28374 (N_28374,N_26871,N_26714);
nor U28375 (N_28375,N_26906,N_27368);
or U28376 (N_28376,N_26452,N_26940);
nand U28377 (N_28377,N_27541,N_26592);
or U28378 (N_28378,N_27328,N_26993);
xnor U28379 (N_28379,N_27126,N_26897);
nor U28380 (N_28380,N_27320,N_26555);
or U28381 (N_28381,N_26877,N_26586);
xnor U28382 (N_28382,N_26868,N_27092);
or U28383 (N_28383,N_27543,N_27407);
xnor U28384 (N_28384,N_26622,N_26732);
and U28385 (N_28385,N_27377,N_27374);
or U28386 (N_28386,N_27118,N_26735);
or U28387 (N_28387,N_27240,N_27524);
xnor U28388 (N_28388,N_27005,N_27378);
nor U28389 (N_28389,N_26992,N_27141);
nor U28390 (N_28390,N_27331,N_27471);
and U28391 (N_28391,N_26601,N_27305);
nand U28392 (N_28392,N_27467,N_27356);
nor U28393 (N_28393,N_26626,N_27447);
or U28394 (N_28394,N_27580,N_27285);
xnor U28395 (N_28395,N_27394,N_27261);
or U28396 (N_28396,N_26981,N_26448);
xor U28397 (N_28397,N_27169,N_27151);
and U28398 (N_28398,N_26869,N_26676);
or U28399 (N_28399,N_27525,N_27094);
or U28400 (N_28400,N_27009,N_26873);
nor U28401 (N_28401,N_27359,N_27196);
xnor U28402 (N_28402,N_26658,N_26890);
and U28403 (N_28403,N_27044,N_26414);
or U28404 (N_28404,N_27108,N_26892);
or U28405 (N_28405,N_26508,N_27274);
or U28406 (N_28406,N_27232,N_27091);
nor U28407 (N_28407,N_26404,N_26742);
xor U28408 (N_28408,N_27589,N_26961);
and U28409 (N_28409,N_26642,N_27223);
nand U28410 (N_28410,N_27000,N_26826);
or U28411 (N_28411,N_27551,N_27380);
xnor U28412 (N_28412,N_27047,N_27268);
nor U28413 (N_28413,N_27487,N_26553);
and U28414 (N_28414,N_27050,N_27427);
or U28415 (N_28415,N_26897,N_27356);
nor U28416 (N_28416,N_27132,N_27193);
or U28417 (N_28417,N_27336,N_27583);
nand U28418 (N_28418,N_27211,N_27071);
nand U28419 (N_28419,N_27510,N_26600);
or U28420 (N_28420,N_27024,N_27585);
xor U28421 (N_28421,N_26408,N_27000);
nor U28422 (N_28422,N_26427,N_27110);
xnor U28423 (N_28423,N_27067,N_26599);
xnor U28424 (N_28424,N_27559,N_27593);
and U28425 (N_28425,N_26639,N_27307);
nand U28426 (N_28426,N_27293,N_27527);
xnor U28427 (N_28427,N_27175,N_27012);
and U28428 (N_28428,N_27530,N_26540);
nor U28429 (N_28429,N_26547,N_27362);
and U28430 (N_28430,N_27098,N_26947);
nor U28431 (N_28431,N_26934,N_26902);
and U28432 (N_28432,N_27283,N_26663);
or U28433 (N_28433,N_26966,N_27339);
nand U28434 (N_28434,N_27195,N_27229);
or U28435 (N_28435,N_27226,N_27503);
and U28436 (N_28436,N_27011,N_26996);
or U28437 (N_28437,N_27058,N_26467);
nand U28438 (N_28438,N_27280,N_27182);
nand U28439 (N_28439,N_26419,N_27336);
nand U28440 (N_28440,N_26865,N_26518);
xnor U28441 (N_28441,N_26511,N_26470);
and U28442 (N_28442,N_27412,N_26533);
xor U28443 (N_28443,N_27599,N_27470);
and U28444 (N_28444,N_26727,N_27266);
or U28445 (N_28445,N_27298,N_27203);
nand U28446 (N_28446,N_27500,N_26443);
nor U28447 (N_28447,N_26882,N_26842);
nand U28448 (N_28448,N_26831,N_27590);
nand U28449 (N_28449,N_27352,N_26990);
xor U28450 (N_28450,N_26951,N_26982);
nand U28451 (N_28451,N_26415,N_26432);
nor U28452 (N_28452,N_26811,N_26604);
and U28453 (N_28453,N_26591,N_27588);
xor U28454 (N_28454,N_27027,N_27500);
nand U28455 (N_28455,N_27198,N_27411);
nor U28456 (N_28456,N_26859,N_27123);
nor U28457 (N_28457,N_26524,N_27080);
nor U28458 (N_28458,N_27410,N_26467);
nand U28459 (N_28459,N_27463,N_27040);
nand U28460 (N_28460,N_27014,N_27142);
and U28461 (N_28461,N_27548,N_27017);
or U28462 (N_28462,N_26962,N_26619);
nor U28463 (N_28463,N_26717,N_26475);
and U28464 (N_28464,N_26504,N_27134);
or U28465 (N_28465,N_26786,N_27423);
xor U28466 (N_28466,N_26509,N_27482);
or U28467 (N_28467,N_26503,N_27306);
or U28468 (N_28468,N_27265,N_27167);
or U28469 (N_28469,N_26963,N_27479);
or U28470 (N_28470,N_27287,N_26847);
xor U28471 (N_28471,N_27351,N_27048);
nor U28472 (N_28472,N_26479,N_27288);
and U28473 (N_28473,N_27282,N_27524);
xor U28474 (N_28474,N_27374,N_26858);
xnor U28475 (N_28475,N_27106,N_27496);
or U28476 (N_28476,N_27465,N_27067);
or U28477 (N_28477,N_26538,N_27127);
xnor U28478 (N_28478,N_26451,N_27341);
nor U28479 (N_28479,N_27526,N_26597);
nand U28480 (N_28480,N_26509,N_26717);
xnor U28481 (N_28481,N_26586,N_27160);
xor U28482 (N_28482,N_26684,N_27575);
and U28483 (N_28483,N_26528,N_26732);
xor U28484 (N_28484,N_27090,N_27510);
and U28485 (N_28485,N_26748,N_26477);
and U28486 (N_28486,N_27016,N_26815);
nand U28487 (N_28487,N_26618,N_27372);
and U28488 (N_28488,N_26481,N_26646);
xor U28489 (N_28489,N_27594,N_26947);
nand U28490 (N_28490,N_26640,N_26547);
xnor U28491 (N_28491,N_27218,N_26992);
nor U28492 (N_28492,N_27539,N_27273);
nor U28493 (N_28493,N_27191,N_27233);
and U28494 (N_28494,N_27274,N_26482);
nand U28495 (N_28495,N_27004,N_26952);
xor U28496 (N_28496,N_26828,N_27241);
and U28497 (N_28497,N_27343,N_27344);
xor U28498 (N_28498,N_27263,N_27275);
nand U28499 (N_28499,N_27047,N_27041);
and U28500 (N_28500,N_27436,N_26723);
nor U28501 (N_28501,N_26540,N_26639);
nor U28502 (N_28502,N_26849,N_26864);
or U28503 (N_28503,N_27575,N_26655);
nand U28504 (N_28504,N_27598,N_27204);
nor U28505 (N_28505,N_26951,N_27107);
and U28506 (N_28506,N_27453,N_26829);
or U28507 (N_28507,N_26884,N_26812);
xnor U28508 (N_28508,N_26848,N_27379);
xor U28509 (N_28509,N_27021,N_26531);
xnor U28510 (N_28510,N_26438,N_26988);
nand U28511 (N_28511,N_26796,N_26480);
nand U28512 (N_28512,N_26479,N_26483);
nor U28513 (N_28513,N_27555,N_26970);
xnor U28514 (N_28514,N_27314,N_26950);
xnor U28515 (N_28515,N_27279,N_26722);
nor U28516 (N_28516,N_26754,N_27130);
nor U28517 (N_28517,N_27295,N_26554);
and U28518 (N_28518,N_26779,N_27474);
xnor U28519 (N_28519,N_27056,N_27276);
nand U28520 (N_28520,N_26621,N_27140);
nand U28521 (N_28521,N_26455,N_27552);
and U28522 (N_28522,N_26819,N_27298);
xor U28523 (N_28523,N_27228,N_27242);
or U28524 (N_28524,N_26421,N_27013);
and U28525 (N_28525,N_26401,N_27004);
and U28526 (N_28526,N_26882,N_27421);
xor U28527 (N_28527,N_26983,N_27394);
and U28528 (N_28528,N_26637,N_26771);
xnor U28529 (N_28529,N_26828,N_27509);
and U28530 (N_28530,N_26823,N_27012);
or U28531 (N_28531,N_27415,N_26996);
nand U28532 (N_28532,N_27160,N_27068);
or U28533 (N_28533,N_26995,N_26403);
nand U28534 (N_28534,N_26434,N_26951);
or U28535 (N_28535,N_27055,N_26630);
nor U28536 (N_28536,N_27236,N_26422);
nor U28537 (N_28537,N_26456,N_27248);
and U28538 (N_28538,N_26431,N_26795);
or U28539 (N_28539,N_26699,N_27385);
or U28540 (N_28540,N_27297,N_26465);
nand U28541 (N_28541,N_27048,N_27108);
nand U28542 (N_28542,N_26951,N_27137);
and U28543 (N_28543,N_27112,N_26820);
xnor U28544 (N_28544,N_26451,N_27018);
or U28545 (N_28545,N_27107,N_26650);
nor U28546 (N_28546,N_27477,N_26929);
and U28547 (N_28547,N_27123,N_27146);
or U28548 (N_28548,N_26734,N_26528);
xor U28549 (N_28549,N_26416,N_26941);
nor U28550 (N_28550,N_26941,N_26714);
nand U28551 (N_28551,N_26951,N_27207);
nor U28552 (N_28552,N_26855,N_27327);
xor U28553 (N_28553,N_27591,N_26508);
and U28554 (N_28554,N_27266,N_26656);
nand U28555 (N_28555,N_26468,N_26768);
xnor U28556 (N_28556,N_27438,N_26518);
nand U28557 (N_28557,N_26651,N_27031);
or U28558 (N_28558,N_27157,N_27393);
or U28559 (N_28559,N_26911,N_27090);
nand U28560 (N_28560,N_26473,N_27323);
nand U28561 (N_28561,N_26751,N_27260);
nor U28562 (N_28562,N_26850,N_27553);
nand U28563 (N_28563,N_26840,N_26829);
or U28564 (N_28564,N_26736,N_26811);
xor U28565 (N_28565,N_27365,N_26783);
or U28566 (N_28566,N_26466,N_26863);
or U28567 (N_28567,N_27322,N_26914);
and U28568 (N_28568,N_27105,N_27463);
nor U28569 (N_28569,N_27285,N_27529);
nor U28570 (N_28570,N_26511,N_26719);
nor U28571 (N_28571,N_27359,N_27190);
or U28572 (N_28572,N_26883,N_27245);
nor U28573 (N_28573,N_27213,N_26806);
nor U28574 (N_28574,N_26690,N_27506);
nor U28575 (N_28575,N_27048,N_26662);
nand U28576 (N_28576,N_26961,N_27138);
xnor U28577 (N_28577,N_26580,N_26769);
nand U28578 (N_28578,N_27247,N_27261);
and U28579 (N_28579,N_26967,N_27334);
and U28580 (N_28580,N_27384,N_26683);
nand U28581 (N_28581,N_27193,N_26621);
xor U28582 (N_28582,N_27112,N_26578);
and U28583 (N_28583,N_26587,N_26761);
nor U28584 (N_28584,N_26802,N_27405);
nand U28585 (N_28585,N_26825,N_26654);
nor U28586 (N_28586,N_26965,N_26427);
nor U28587 (N_28587,N_26924,N_26535);
xnor U28588 (N_28588,N_26663,N_27516);
nand U28589 (N_28589,N_27590,N_27204);
nand U28590 (N_28590,N_26894,N_27447);
nand U28591 (N_28591,N_26483,N_27247);
nand U28592 (N_28592,N_27411,N_26829);
nor U28593 (N_28593,N_27065,N_26491);
xor U28594 (N_28594,N_27096,N_27363);
nor U28595 (N_28595,N_27057,N_26997);
and U28596 (N_28596,N_27491,N_27248);
or U28597 (N_28597,N_26788,N_27387);
and U28598 (N_28598,N_26866,N_27413);
xnor U28599 (N_28599,N_27138,N_27496);
or U28600 (N_28600,N_26528,N_26435);
or U28601 (N_28601,N_26987,N_26450);
xor U28602 (N_28602,N_26992,N_27010);
and U28603 (N_28603,N_26504,N_27114);
nor U28604 (N_28604,N_26853,N_26515);
xor U28605 (N_28605,N_27243,N_26545);
xor U28606 (N_28606,N_27550,N_26933);
and U28607 (N_28607,N_26431,N_27415);
nor U28608 (N_28608,N_27175,N_27148);
and U28609 (N_28609,N_26977,N_27574);
xnor U28610 (N_28610,N_26734,N_26983);
xnor U28611 (N_28611,N_27132,N_27121);
nand U28612 (N_28612,N_26931,N_27123);
or U28613 (N_28613,N_27587,N_26634);
nor U28614 (N_28614,N_27488,N_27492);
or U28615 (N_28615,N_26895,N_26798);
and U28616 (N_28616,N_27218,N_27422);
xor U28617 (N_28617,N_26726,N_26612);
xnor U28618 (N_28618,N_26665,N_27112);
xnor U28619 (N_28619,N_26891,N_27278);
and U28620 (N_28620,N_27472,N_27599);
or U28621 (N_28621,N_27376,N_26820);
and U28622 (N_28622,N_27082,N_26591);
nand U28623 (N_28623,N_26552,N_27260);
nor U28624 (N_28624,N_26428,N_26577);
nand U28625 (N_28625,N_27051,N_26977);
nor U28626 (N_28626,N_26703,N_27198);
nand U28627 (N_28627,N_27113,N_27222);
and U28628 (N_28628,N_27315,N_26666);
or U28629 (N_28629,N_27333,N_27586);
or U28630 (N_28630,N_27506,N_26519);
or U28631 (N_28631,N_26583,N_27463);
nor U28632 (N_28632,N_27265,N_26540);
nor U28633 (N_28633,N_27358,N_27270);
nand U28634 (N_28634,N_27138,N_26683);
and U28635 (N_28635,N_26812,N_26437);
and U28636 (N_28636,N_27224,N_26485);
or U28637 (N_28637,N_26432,N_27512);
and U28638 (N_28638,N_26524,N_27010);
nand U28639 (N_28639,N_26462,N_26973);
xor U28640 (N_28640,N_26423,N_27070);
nor U28641 (N_28641,N_26530,N_26473);
nand U28642 (N_28642,N_26683,N_26649);
or U28643 (N_28643,N_27377,N_26456);
nor U28644 (N_28644,N_27415,N_27391);
nand U28645 (N_28645,N_26421,N_27447);
nand U28646 (N_28646,N_26958,N_26417);
nand U28647 (N_28647,N_27378,N_27170);
and U28648 (N_28648,N_27297,N_26940);
or U28649 (N_28649,N_26985,N_27548);
and U28650 (N_28650,N_26577,N_26618);
nor U28651 (N_28651,N_26610,N_27487);
nor U28652 (N_28652,N_26894,N_26861);
xnor U28653 (N_28653,N_26760,N_27058);
nand U28654 (N_28654,N_27164,N_27364);
or U28655 (N_28655,N_26627,N_27544);
or U28656 (N_28656,N_26859,N_26417);
nor U28657 (N_28657,N_26942,N_26477);
nand U28658 (N_28658,N_26751,N_27172);
nor U28659 (N_28659,N_27221,N_27225);
and U28660 (N_28660,N_26724,N_26867);
xor U28661 (N_28661,N_26715,N_27368);
or U28662 (N_28662,N_26769,N_27474);
xor U28663 (N_28663,N_26515,N_26671);
nand U28664 (N_28664,N_26459,N_27111);
or U28665 (N_28665,N_26979,N_26608);
nor U28666 (N_28666,N_26511,N_26640);
xnor U28667 (N_28667,N_26891,N_27375);
or U28668 (N_28668,N_27368,N_27259);
nand U28669 (N_28669,N_27528,N_26827);
nor U28670 (N_28670,N_27482,N_27207);
or U28671 (N_28671,N_27100,N_27158);
nor U28672 (N_28672,N_27539,N_26825);
xnor U28673 (N_28673,N_26977,N_27358);
xnor U28674 (N_28674,N_27396,N_26649);
xor U28675 (N_28675,N_26437,N_26778);
and U28676 (N_28676,N_26491,N_26544);
nor U28677 (N_28677,N_27066,N_27491);
xnor U28678 (N_28678,N_26739,N_26650);
nand U28679 (N_28679,N_27240,N_26607);
or U28680 (N_28680,N_26933,N_26488);
nand U28681 (N_28681,N_26988,N_26831);
or U28682 (N_28682,N_27426,N_27332);
or U28683 (N_28683,N_26793,N_26552);
and U28684 (N_28684,N_27039,N_26688);
nor U28685 (N_28685,N_26890,N_26438);
xnor U28686 (N_28686,N_27047,N_26683);
nand U28687 (N_28687,N_27171,N_26690);
nor U28688 (N_28688,N_27463,N_26828);
and U28689 (N_28689,N_27229,N_27221);
nand U28690 (N_28690,N_27480,N_27162);
or U28691 (N_28691,N_27025,N_26809);
nor U28692 (N_28692,N_26808,N_26974);
and U28693 (N_28693,N_26844,N_26536);
or U28694 (N_28694,N_26816,N_27410);
nor U28695 (N_28695,N_27396,N_27220);
nor U28696 (N_28696,N_27191,N_27303);
or U28697 (N_28697,N_27153,N_27571);
or U28698 (N_28698,N_27428,N_26764);
or U28699 (N_28699,N_27230,N_27441);
and U28700 (N_28700,N_26503,N_26731);
and U28701 (N_28701,N_26536,N_26773);
nand U28702 (N_28702,N_27146,N_27131);
or U28703 (N_28703,N_27177,N_26979);
nand U28704 (N_28704,N_27553,N_26841);
nand U28705 (N_28705,N_27146,N_26597);
and U28706 (N_28706,N_27579,N_26743);
and U28707 (N_28707,N_26495,N_27161);
or U28708 (N_28708,N_26819,N_27513);
or U28709 (N_28709,N_26880,N_27557);
nor U28710 (N_28710,N_27038,N_27236);
nor U28711 (N_28711,N_27271,N_26457);
nand U28712 (N_28712,N_27199,N_26417);
nor U28713 (N_28713,N_26690,N_26951);
and U28714 (N_28714,N_27456,N_27562);
xor U28715 (N_28715,N_27283,N_26773);
nor U28716 (N_28716,N_26860,N_27554);
or U28717 (N_28717,N_26971,N_27505);
nand U28718 (N_28718,N_27069,N_26788);
nand U28719 (N_28719,N_26685,N_26736);
nand U28720 (N_28720,N_26780,N_27028);
nor U28721 (N_28721,N_26693,N_26976);
nand U28722 (N_28722,N_26425,N_26918);
or U28723 (N_28723,N_27069,N_27099);
and U28724 (N_28724,N_26924,N_26545);
nand U28725 (N_28725,N_26770,N_27050);
or U28726 (N_28726,N_27377,N_27450);
xnor U28727 (N_28727,N_27203,N_26541);
nand U28728 (N_28728,N_27466,N_27292);
xor U28729 (N_28729,N_27529,N_27383);
or U28730 (N_28730,N_27580,N_27005);
or U28731 (N_28731,N_27315,N_27505);
and U28732 (N_28732,N_27351,N_27586);
nand U28733 (N_28733,N_26536,N_27554);
nand U28734 (N_28734,N_27411,N_26877);
nor U28735 (N_28735,N_26736,N_27553);
nand U28736 (N_28736,N_26424,N_27377);
xor U28737 (N_28737,N_27090,N_26955);
nand U28738 (N_28738,N_26535,N_26500);
nor U28739 (N_28739,N_27456,N_26572);
xnor U28740 (N_28740,N_26455,N_26694);
or U28741 (N_28741,N_26495,N_27233);
and U28742 (N_28742,N_26705,N_26825);
xnor U28743 (N_28743,N_27455,N_27268);
nand U28744 (N_28744,N_27055,N_26775);
nand U28745 (N_28745,N_26821,N_27315);
or U28746 (N_28746,N_26486,N_27157);
nor U28747 (N_28747,N_26716,N_26862);
xor U28748 (N_28748,N_27213,N_26421);
and U28749 (N_28749,N_27003,N_26826);
xnor U28750 (N_28750,N_27286,N_27207);
nand U28751 (N_28751,N_26972,N_26743);
nand U28752 (N_28752,N_27063,N_27131);
nand U28753 (N_28753,N_26607,N_26973);
xnor U28754 (N_28754,N_26776,N_26876);
nor U28755 (N_28755,N_27223,N_27415);
nor U28756 (N_28756,N_27329,N_27007);
xnor U28757 (N_28757,N_26774,N_26472);
and U28758 (N_28758,N_27203,N_27024);
and U28759 (N_28759,N_27019,N_26491);
xor U28760 (N_28760,N_27268,N_27093);
and U28761 (N_28761,N_27060,N_27290);
nand U28762 (N_28762,N_27493,N_27550);
xnor U28763 (N_28763,N_27074,N_26981);
xor U28764 (N_28764,N_26418,N_26635);
and U28765 (N_28765,N_26660,N_26963);
nor U28766 (N_28766,N_26794,N_26624);
nor U28767 (N_28767,N_26545,N_27151);
or U28768 (N_28768,N_27223,N_27457);
and U28769 (N_28769,N_26537,N_26878);
nand U28770 (N_28770,N_27023,N_26453);
nor U28771 (N_28771,N_27592,N_27073);
xnor U28772 (N_28772,N_27278,N_26969);
nor U28773 (N_28773,N_27555,N_26866);
and U28774 (N_28774,N_27325,N_26745);
and U28775 (N_28775,N_26769,N_27072);
xnor U28776 (N_28776,N_27046,N_26520);
and U28777 (N_28777,N_26552,N_26592);
nor U28778 (N_28778,N_27397,N_26878);
and U28779 (N_28779,N_26509,N_27093);
and U28780 (N_28780,N_26894,N_26727);
nand U28781 (N_28781,N_27182,N_26877);
nand U28782 (N_28782,N_27580,N_26400);
xor U28783 (N_28783,N_27134,N_27182);
and U28784 (N_28784,N_27091,N_26879);
nand U28785 (N_28785,N_27036,N_26787);
or U28786 (N_28786,N_26716,N_26912);
or U28787 (N_28787,N_26599,N_27186);
or U28788 (N_28788,N_27124,N_27523);
and U28789 (N_28789,N_27576,N_27103);
xnor U28790 (N_28790,N_27128,N_27280);
or U28791 (N_28791,N_27449,N_27335);
or U28792 (N_28792,N_26455,N_27572);
nand U28793 (N_28793,N_27304,N_27214);
nor U28794 (N_28794,N_26965,N_26617);
and U28795 (N_28795,N_26847,N_27174);
nor U28796 (N_28796,N_26949,N_26611);
nand U28797 (N_28797,N_26482,N_26851);
nor U28798 (N_28798,N_26870,N_27571);
nand U28799 (N_28799,N_27525,N_26692);
xnor U28800 (N_28800,N_28411,N_27887);
or U28801 (N_28801,N_27975,N_28401);
nand U28802 (N_28802,N_28356,N_28440);
or U28803 (N_28803,N_27996,N_28350);
and U28804 (N_28804,N_28735,N_27639);
and U28805 (N_28805,N_28711,N_27811);
and U28806 (N_28806,N_27621,N_27979);
xor U28807 (N_28807,N_27623,N_27720);
nand U28808 (N_28808,N_28265,N_28017);
xnor U28809 (N_28809,N_28639,N_28743);
or U28810 (N_28810,N_27840,N_28488);
nand U28811 (N_28811,N_28293,N_27873);
or U28812 (N_28812,N_28039,N_27907);
nand U28813 (N_28813,N_28114,N_27947);
nor U28814 (N_28814,N_28789,N_27966);
nor U28815 (N_28815,N_27831,N_28042);
xor U28816 (N_28816,N_28694,N_27763);
or U28817 (N_28817,N_28489,N_28018);
nand U28818 (N_28818,N_28438,N_27883);
nor U28819 (N_28819,N_28298,N_28523);
xnor U28820 (N_28820,N_27861,N_28797);
and U28821 (N_28821,N_28455,N_28349);
nand U28822 (N_28822,N_27889,N_28552);
nand U28823 (N_28823,N_28103,N_28062);
or U28824 (N_28824,N_28340,N_28315);
or U28825 (N_28825,N_28270,N_27886);
nand U28826 (N_28826,N_28646,N_27788);
or U28827 (N_28827,N_28511,N_27854);
or U28828 (N_28828,N_27839,N_28447);
and U28829 (N_28829,N_28628,N_28359);
and U28830 (N_28830,N_27875,N_27827);
and U28831 (N_28831,N_28212,N_28543);
and U28832 (N_28832,N_28519,N_28645);
and U28833 (N_28833,N_28445,N_28760);
nand U28834 (N_28834,N_28416,N_28613);
or U28835 (N_28835,N_27712,N_27882);
nand U28836 (N_28836,N_28490,N_28703);
and U28837 (N_28837,N_28091,N_28081);
xnor U28838 (N_28838,N_28547,N_28339);
and U28839 (N_28839,N_27704,N_28650);
or U28840 (N_28840,N_27800,N_27798);
or U28841 (N_28841,N_28742,N_27904);
nor U28842 (N_28842,N_28205,N_28408);
nand U28843 (N_28843,N_28257,N_28381);
xnor U28844 (N_28844,N_28412,N_28510);
nor U28845 (N_28845,N_28560,N_28219);
nand U28846 (N_28846,N_28341,N_28175);
nor U28847 (N_28847,N_28579,N_28693);
nand U28848 (N_28848,N_27717,N_28286);
nor U28849 (N_28849,N_27685,N_28058);
xor U28850 (N_28850,N_28558,N_28136);
nand U28851 (N_28851,N_28528,N_27863);
nor U28852 (N_28852,N_27986,N_28569);
or U28853 (N_28853,N_28435,N_27707);
nor U28854 (N_28854,N_27933,N_28718);
and U28855 (N_28855,N_28413,N_28477);
nand U28856 (N_28856,N_28451,N_28657);
nor U28857 (N_28857,N_28456,N_28141);
nand U28858 (N_28858,N_27995,N_28326);
or U28859 (N_28859,N_27965,N_28085);
or U28860 (N_28860,N_28464,N_27708);
xor U28861 (N_28861,N_27999,N_28061);
nor U28862 (N_28862,N_27769,N_28223);
and U28863 (N_28863,N_27761,N_28037);
and U28864 (N_28864,N_28502,N_28565);
nand U28865 (N_28865,N_28596,N_27692);
or U28866 (N_28866,N_28330,N_28758);
xnor U28867 (N_28867,N_28163,N_27984);
xnor U28868 (N_28868,N_28788,N_27964);
nor U28869 (N_28869,N_28000,N_28222);
nor U28870 (N_28870,N_28483,N_28656);
and U28871 (N_28871,N_28513,N_27749);
or U28872 (N_28872,N_27968,N_28666);
and U28873 (N_28873,N_27916,N_28331);
and U28874 (N_28874,N_28497,N_27684);
nor U28875 (N_28875,N_28779,N_27715);
and U28876 (N_28876,N_28710,N_28673);
nor U28877 (N_28877,N_28151,N_28618);
nand U28878 (N_28878,N_28199,N_27668);
xnor U28879 (N_28879,N_27696,N_28626);
or U28880 (N_28880,N_28550,N_28010);
nand U28881 (N_28881,N_28736,N_28679);
and U28882 (N_28882,N_28759,N_27772);
xnor U28883 (N_28883,N_28778,N_28684);
nor U28884 (N_28884,N_28159,N_28140);
or U28885 (N_28885,N_28194,N_27655);
nand U28886 (N_28886,N_27843,N_28697);
xor U28887 (N_28887,N_28516,N_28250);
nand U28888 (N_28888,N_28690,N_27688);
and U28889 (N_28889,N_28745,N_28486);
nor U28890 (N_28890,N_28067,N_28252);
or U28891 (N_28891,N_27961,N_28491);
nand U28892 (N_28892,N_27697,N_28109);
nor U28893 (N_28893,N_27837,N_27726);
and U28894 (N_28894,N_28299,N_27755);
or U28895 (N_28895,N_28083,N_28229);
and U28896 (N_28896,N_28709,N_28344);
nand U28897 (N_28897,N_28323,N_28009);
xnor U28898 (N_28898,N_27991,N_28783);
and U28899 (N_28899,N_28170,N_28167);
xnor U28900 (N_28900,N_28303,N_28734);
and U28901 (N_28901,N_28134,N_27799);
or U28902 (N_28902,N_28021,N_28052);
xor U28903 (N_28903,N_28110,N_28430);
nor U28904 (N_28904,N_28393,N_27808);
nor U28905 (N_28905,N_27943,N_27906);
nor U28906 (N_28906,N_27691,N_27862);
xor U28907 (N_28907,N_28396,N_28769);
or U28908 (N_28908,N_28441,N_28634);
xor U28909 (N_28909,N_28149,N_27924);
or U28910 (N_28910,N_27928,N_27758);
nand U28911 (N_28911,N_28678,N_28544);
and U28912 (N_28912,N_28568,N_27821);
or U28913 (N_28913,N_27624,N_28708);
nor U28914 (N_28914,N_27713,N_28095);
or U28915 (N_28915,N_28255,N_28145);
nand U28916 (N_28916,N_28672,N_28115);
xnor U28917 (N_28917,N_28600,N_27678);
and U28918 (N_28918,N_27665,N_28328);
nor U28919 (N_28919,N_28006,N_28147);
nand U28920 (N_28920,N_28705,N_27909);
or U28921 (N_28921,N_28732,N_27675);
or U28922 (N_28922,N_27662,N_28234);
xnor U28923 (N_28923,N_28403,N_27884);
xnor U28924 (N_28924,N_28587,N_28774);
nand U28925 (N_28925,N_28022,N_28125);
nand U28926 (N_28926,N_28518,N_28087);
or U28927 (N_28927,N_28271,N_28740);
nand U28928 (N_28928,N_27780,N_28480);
nor U28929 (N_28929,N_28195,N_28231);
nand U28930 (N_28930,N_28545,N_27954);
xor U28931 (N_28931,N_28176,N_27676);
nand U28932 (N_28932,N_27718,N_27736);
and U28933 (N_28933,N_28570,N_27743);
nor U28934 (N_28934,N_28251,N_28549);
or U28935 (N_28935,N_28644,N_27617);
and U28936 (N_28936,N_28319,N_28578);
xor U28937 (N_28937,N_28417,N_28671);
and U28938 (N_28938,N_28047,N_28571);
xor U28939 (N_28939,N_28691,N_28036);
nor U28940 (N_28940,N_28476,N_28425);
xor U28941 (N_28941,N_28075,N_27638);
xnor U28942 (N_28942,N_28505,N_28386);
xor U28943 (N_28943,N_28046,N_28700);
xnor U28944 (N_28944,N_28316,N_28226);
nand U28945 (N_28945,N_27950,N_28228);
nor U28946 (N_28946,N_27709,N_28224);
and U28947 (N_28947,N_28437,N_28675);
and U28948 (N_28948,N_28765,N_28215);
or U28949 (N_28949,N_28495,N_27997);
or U28950 (N_28950,N_27871,N_28757);
xor U28951 (N_28951,N_28637,N_28238);
and U28952 (N_28952,N_27880,N_27728);
or U28953 (N_28953,N_27642,N_27716);
nor U28954 (N_28954,N_28164,N_28111);
or U28955 (N_28955,N_28439,N_28272);
and U28956 (N_28956,N_28135,N_27687);
nand U28957 (N_28957,N_28730,N_27838);
or U28958 (N_28958,N_28374,N_28460);
xnor U28959 (N_28959,N_28669,N_28168);
or U28960 (N_28960,N_28603,N_28706);
and U28961 (N_28961,N_27876,N_28245);
and U28962 (N_28962,N_27711,N_27795);
nor U28963 (N_28963,N_27633,N_28492);
and U28964 (N_28964,N_27867,N_27959);
or U28965 (N_28965,N_28107,N_28443);
nand U28966 (N_28966,N_28225,N_28246);
nand U28967 (N_28967,N_28643,N_28457);
nand U28968 (N_28968,N_28232,N_28373);
nand U28969 (N_28969,N_28296,N_27865);
nand U28970 (N_28970,N_27751,N_28343);
and U28971 (N_28971,N_28053,N_28621);
nor U28972 (N_28972,N_28243,N_28566);
and U28973 (N_28973,N_27686,N_27955);
xnor U28974 (N_28974,N_28239,N_28512);
nor U28975 (N_28975,N_28715,N_28398);
nand U28976 (N_28976,N_27657,N_27990);
nor U28977 (N_28977,N_27829,N_27896);
xor U28978 (N_28978,N_28410,N_28065);
nor U28979 (N_28979,N_28770,N_28099);
xnor U28980 (N_28980,N_27635,N_27608);
nor U28981 (N_28981,N_28415,N_28470);
nor U28982 (N_28982,N_28612,N_28129);
xor U28983 (N_28983,N_28186,N_27866);
nor U28984 (N_28984,N_28450,N_28355);
or U28985 (N_28985,N_28572,N_28153);
nor U28986 (N_28986,N_28027,N_27819);
nor U28987 (N_28987,N_27872,N_27976);
nand U28988 (N_28988,N_27836,N_27745);
or U28989 (N_28989,N_28309,N_28409);
nand U28990 (N_28990,N_27994,N_27849);
or U28991 (N_28991,N_27698,N_28414);
and U28992 (N_28992,N_27683,N_28794);
or U28993 (N_28993,N_28764,N_28320);
nor U28994 (N_28994,N_28102,N_27905);
and U28995 (N_28995,N_28761,N_28367);
nand U28996 (N_28996,N_28122,N_27803);
or U28997 (N_28997,N_27703,N_28419);
and U28998 (N_28998,N_28210,N_28586);
nor U28999 (N_28999,N_28216,N_28487);
xnor U29000 (N_29000,N_27774,N_27792);
xnor U29001 (N_29001,N_27952,N_27693);
and U29002 (N_29002,N_28244,N_27659);
and U29003 (N_29003,N_27941,N_28683);
xnor U29004 (N_29004,N_27851,N_27796);
xnor U29005 (N_29005,N_27768,N_28448);
or U29006 (N_29006,N_28559,N_28092);
nand U29007 (N_29007,N_27636,N_28322);
nor U29008 (N_29008,N_28484,N_28206);
nand U29009 (N_29009,N_28124,N_28235);
or U29010 (N_29010,N_28689,N_28466);
nor U29011 (N_29011,N_28695,N_27765);
or U29012 (N_29012,N_28201,N_28467);
nand U29013 (N_29013,N_27742,N_28337);
nand U29014 (N_29014,N_28647,N_27852);
xnor U29015 (N_29015,N_28627,N_27900);
nor U29016 (N_29016,N_28591,N_28629);
and U29017 (N_29017,N_28190,N_28453);
nand U29018 (N_29018,N_27998,N_28539);
or U29019 (N_29019,N_28066,N_28658);
or U29020 (N_29020,N_27634,N_27701);
nand U29021 (N_29021,N_28527,N_27985);
nor U29022 (N_29022,N_28722,N_27978);
nor U29023 (N_29023,N_28059,N_28481);
nand U29024 (N_29024,N_28790,N_27787);
xnor U29025 (N_29025,N_27694,N_28659);
or U29026 (N_29026,N_28332,N_27641);
and U29027 (N_29027,N_27982,N_28529);
nand U29028 (N_29028,N_27897,N_28288);
nand U29029 (N_29029,N_28432,N_27719);
nand U29030 (N_29030,N_28653,N_28280);
and U29031 (N_29031,N_28593,N_28585);
nand U29032 (N_29032,N_27894,N_27784);
nor U29033 (N_29033,N_28589,N_28729);
and U29034 (N_29034,N_28763,N_28236);
xor U29035 (N_29035,N_28617,N_28093);
nor U29036 (N_29036,N_28055,N_28424);
nand U29037 (N_29037,N_28044,N_27877);
xnor U29038 (N_29038,N_28353,N_27680);
xnor U29039 (N_29039,N_27644,N_28638);
nor U29040 (N_29040,N_27814,N_28670);
nor U29041 (N_29041,N_28040,N_28173);
xor U29042 (N_29042,N_27935,N_28562);
nor U29043 (N_29043,N_28015,N_27731);
xnor U29044 (N_29044,N_27818,N_28597);
nand U29045 (N_29045,N_28325,N_27927);
nand U29046 (N_29046,N_27972,N_27604);
and U29047 (N_29047,N_28258,N_28172);
nor U29048 (N_29048,N_28407,N_28594);
xor U29049 (N_29049,N_28090,N_28079);
xor U29050 (N_29050,N_28035,N_28610);
nor U29051 (N_29051,N_27930,N_28792);
nand U29052 (N_29052,N_28204,N_28793);
nand U29053 (N_29053,N_28625,N_28713);
nand U29054 (N_29054,N_28171,N_28786);
nand U29055 (N_29055,N_28148,N_28121);
or U29056 (N_29056,N_28050,N_28459);
nor U29057 (N_29057,N_27932,N_28567);
nor U29058 (N_29058,N_27806,N_27901);
nor U29059 (N_29059,N_27674,N_28588);
and U29060 (N_29060,N_28064,N_27936);
xnor U29061 (N_29061,N_28318,N_28423);
nor U29062 (N_29062,N_28573,N_28247);
and U29063 (N_29063,N_28772,N_28023);
xnor U29064 (N_29064,N_27670,N_28139);
nor U29065 (N_29065,N_28514,N_27681);
nand U29066 (N_29066,N_27810,N_28184);
and U29067 (N_29067,N_27812,N_28198);
nand U29068 (N_29068,N_28422,N_28004);
xor U29069 (N_29069,N_27611,N_28192);
nand U29070 (N_29070,N_27620,N_28601);
or U29071 (N_29071,N_27918,N_28752);
xor U29072 (N_29072,N_27614,N_28185);
nand U29073 (N_29073,N_28074,N_27885);
or U29074 (N_29074,N_27922,N_27816);
and U29075 (N_29075,N_27741,N_27962);
xnor U29076 (N_29076,N_28369,N_28775);
nor U29077 (N_29077,N_28312,N_28724);
or U29078 (N_29078,N_28463,N_28418);
and U29079 (N_29079,N_28507,N_28582);
nor U29080 (N_29080,N_28631,N_28624);
nand U29081 (N_29081,N_28755,N_28385);
nand U29082 (N_29082,N_28282,N_27898);
nand U29083 (N_29083,N_27789,N_27949);
nand U29084 (N_29084,N_27878,N_28276);
and U29085 (N_29085,N_28060,N_28378);
or U29086 (N_29086,N_27729,N_27738);
nor U29087 (N_29087,N_28317,N_28520);
or U29088 (N_29088,N_27673,N_28329);
and U29089 (N_29089,N_28746,N_28465);
nand U29090 (N_29090,N_27753,N_28214);
or U29091 (N_29091,N_28599,N_28458);
xor U29092 (N_29092,N_28056,N_28782);
xor U29093 (N_29093,N_28461,N_28426);
nor U29094 (N_29094,N_28032,N_28576);
nand U29095 (N_29095,N_27627,N_28592);
and U29096 (N_29096,N_28712,N_28605);
nor U29097 (N_29097,N_28595,N_27615);
nor U29098 (N_29098,N_28651,N_27920);
xor U29099 (N_29099,N_28479,N_28564);
nor U29100 (N_29100,N_28632,N_28640);
and U29101 (N_29101,N_27946,N_28554);
nand U29102 (N_29102,N_28581,N_28105);
xor U29103 (N_29103,N_27942,N_28749);
nand U29104 (N_29104,N_27605,N_27859);
and U29105 (N_29105,N_28274,N_28155);
nand U29106 (N_29106,N_28086,N_28157);
xor U29107 (N_29107,N_28498,N_28721);
or U29108 (N_29108,N_27853,N_28364);
xnor U29109 (N_29109,N_28311,N_28744);
nand U29110 (N_29110,N_28767,N_28241);
nor U29111 (N_29111,N_27759,N_28748);
nor U29112 (N_29112,N_27649,N_27899);
xor U29113 (N_29113,N_28150,N_27770);
xnor U29114 (N_29114,N_28473,N_28382);
and U29115 (N_29115,N_28324,N_27663);
xnor U29116 (N_29116,N_28394,N_27864);
nor U29117 (N_29117,N_28526,N_28667);
nand U29118 (N_29118,N_27915,N_27848);
nand U29119 (N_29119,N_28619,N_27817);
or U29120 (N_29120,N_28371,N_27804);
nor U29121 (N_29121,N_28716,N_27855);
nor U29122 (N_29122,N_27622,N_27970);
or U29123 (N_29123,N_28183,N_28063);
nor U29124 (N_29124,N_27791,N_28030);
nand U29125 (N_29125,N_27654,N_28029);
xnor U29126 (N_29126,N_27912,N_27782);
xnor U29127 (N_29127,N_28402,N_28073);
xnor U29128 (N_29128,N_28256,N_28146);
nand U29129 (N_29129,N_27793,N_27895);
or U29130 (N_29130,N_27705,N_28723);
and U29131 (N_29131,N_28444,N_28387);
nor U29132 (N_29132,N_28663,N_28284);
or U29133 (N_29133,N_28446,N_27797);
xor U29134 (N_29134,N_28652,N_27706);
or U29135 (N_29135,N_28266,N_27747);
or U29136 (N_29136,N_28674,N_27777);
nand U29137 (N_29137,N_28692,N_28242);
xnor U29138 (N_29138,N_27746,N_28395);
nor U29139 (N_29139,N_28714,N_28113);
and U29140 (N_29140,N_28676,N_27893);
or U29141 (N_29141,N_28524,N_28662);
and U29142 (N_29142,N_28379,N_27771);
nand U29143 (N_29143,N_28048,N_28208);
nor U29144 (N_29144,N_28025,N_27656);
nand U29145 (N_29145,N_27903,N_28162);
nor U29146 (N_29146,N_27667,N_27658);
nand U29147 (N_29147,N_27606,N_28376);
and U29148 (N_29148,N_28682,N_28737);
nor U29149 (N_29149,N_28200,N_27891);
and U29150 (N_29150,N_28260,N_28001);
xnor U29151 (N_29151,N_28615,N_28160);
nor U29152 (N_29152,N_27648,N_27723);
nor U29153 (N_29153,N_28421,N_28211);
nor U29154 (N_29154,N_28360,N_28751);
nor U29155 (N_29155,N_27881,N_28454);
nand U29156 (N_29156,N_27913,N_27987);
and U29157 (N_29157,N_28154,N_28361);
nor U29158 (N_29158,N_28471,N_27664);
xnor U29159 (N_29159,N_28144,N_27923);
nand U29160 (N_29160,N_28633,N_28281);
nor U29161 (N_29161,N_27825,N_27646);
nand U29162 (N_29162,N_28166,N_27980);
nor U29163 (N_29163,N_27695,N_28301);
nor U29164 (N_29164,N_27993,N_27842);
nor U29165 (N_29165,N_28556,N_28366);
nor U29166 (N_29166,N_28370,N_27779);
nand U29167 (N_29167,N_27600,N_28537);
nor U29168 (N_29168,N_27815,N_28704);
nor U29169 (N_29169,N_27832,N_27910);
or U29170 (N_29170,N_28462,N_28762);
xor U29171 (N_29171,N_28494,N_28687);
and U29172 (N_29172,N_27757,N_27937);
and U29173 (N_29173,N_27939,N_28305);
nand U29174 (N_29174,N_27822,N_27677);
nor U29175 (N_29175,N_28026,N_28531);
nor U29176 (N_29176,N_28623,N_27764);
and U29177 (N_29177,N_28133,N_27874);
nand U29178 (N_29178,N_28750,N_27858);
and U29179 (N_29179,N_28654,N_28449);
or U29180 (N_29180,N_28614,N_28089);
nand U29181 (N_29181,N_28493,N_27888);
nor U29182 (N_29182,N_28269,N_28606);
nand U29183 (N_29183,N_28277,N_28038);
or U29184 (N_29184,N_28636,N_28431);
xnor U29185 (N_29185,N_27739,N_28043);
nor U29186 (N_29186,N_28268,N_28118);
nand U29187 (N_29187,N_27992,N_28563);
nand U29188 (N_29188,N_28391,N_28347);
xnor U29189 (N_29189,N_27630,N_28327);
and U29190 (N_29190,N_27834,N_27653);
nand U29191 (N_29191,N_27748,N_28207);
xnor U29192 (N_29192,N_28005,N_28427);
nor U29193 (N_29193,N_27981,N_28616);
or U29194 (N_29194,N_28094,N_27690);
nor U29195 (N_29195,N_27652,N_27989);
xnor U29196 (N_29196,N_27781,N_28611);
and U29197 (N_29197,N_27805,N_28002);
nand U29198 (N_29198,N_28680,N_28101);
xnor U29199 (N_29199,N_28011,N_28525);
xnor U29200 (N_29200,N_27661,N_28719);
and U29201 (N_29201,N_28368,N_28177);
nand U29202 (N_29202,N_28538,N_27682);
nand U29203 (N_29203,N_27601,N_27754);
nand U29204 (N_29204,N_28070,N_28203);
nand U29205 (N_29205,N_28738,N_28100);
nand U29206 (N_29206,N_28338,N_28574);
and U29207 (N_29207,N_27846,N_28237);
or U29208 (N_29208,N_27809,N_28024);
xor U29209 (N_29209,N_27737,N_28182);
or U29210 (N_29210,N_28012,N_27647);
nand U29211 (N_29211,N_28434,N_27724);
nor U29212 (N_29212,N_27645,N_28187);
nor U29213 (N_29213,N_27650,N_28076);
or U29214 (N_29214,N_27689,N_27926);
xnor U29215 (N_29215,N_28165,N_28112);
xnor U29216 (N_29216,N_28766,N_27857);
or U29217 (N_29217,N_28791,N_27786);
and U29218 (N_29218,N_28088,N_28590);
nand U29219 (N_29219,N_28197,N_28196);
or U29220 (N_29220,N_28688,N_28096);
and U29221 (N_29221,N_28661,N_28346);
xor U29222 (N_29222,N_28399,N_27890);
or U29223 (N_29223,N_28137,N_28003);
and U29224 (N_29224,N_27813,N_28392);
or U29225 (N_29225,N_28209,N_28054);
nor U29226 (N_29226,N_27640,N_27917);
nor U29227 (N_29227,N_28390,N_28362);
xnor U29228 (N_29228,N_27613,N_28278);
and U29229 (N_29229,N_28358,N_28248);
xnor U29230 (N_29230,N_28383,N_27734);
and U29231 (N_29231,N_27977,N_27628);
nand U29232 (N_29232,N_28377,N_28283);
nand U29233 (N_29233,N_27612,N_28655);
or U29234 (N_29234,N_28178,N_27660);
nor U29235 (N_29235,N_28668,N_27725);
nor U29236 (N_29236,N_28754,N_28375);
nor U29237 (N_29237,N_28138,N_28607);
xor U29238 (N_29238,N_27618,N_27752);
nor U29239 (N_29239,N_28253,N_28785);
and U29240 (N_29240,N_28007,N_28726);
or U29241 (N_29241,N_28077,N_27826);
xnor U29242 (N_29242,N_28230,N_27609);
xor U29243 (N_29243,N_27960,N_28433);
nor U29244 (N_29244,N_27762,N_28336);
or U29245 (N_29245,N_28189,N_27672);
nor U29246 (N_29246,N_27776,N_28174);
and U29247 (N_29247,N_28262,N_28097);
and U29248 (N_29248,N_28126,N_28254);
xor U29249 (N_29249,N_28045,N_28583);
or U29250 (N_29250,N_27974,N_28249);
nor U29251 (N_29251,N_28041,N_28532);
or U29252 (N_29252,N_28686,N_28795);
nor U29253 (N_29253,N_28108,N_28302);
nand U29254 (N_29254,N_27794,N_27911);
nor U29255 (N_29255,N_28546,N_27969);
nor U29256 (N_29256,N_28753,N_27919);
xnor U29257 (N_29257,N_28389,N_28580);
nor U29258 (N_29258,N_28279,N_28648);
and U29259 (N_29259,N_27957,N_28221);
xnor U29260 (N_29260,N_28130,N_28622);
nand U29261 (N_29261,N_27807,N_28406);
xnor U29262 (N_29262,N_28474,N_28259);
and U29263 (N_29263,N_28768,N_27948);
nand U29264 (N_29264,N_28798,N_28741);
nand U29265 (N_29265,N_28188,N_28291);
or U29266 (N_29266,N_27730,N_27938);
nor U29267 (N_29267,N_28584,N_27956);
nand U29268 (N_29268,N_28120,N_27740);
nor U29269 (N_29269,N_27610,N_28404);
or U29270 (N_29270,N_28530,N_28747);
nor U29271 (N_29271,N_28142,N_28127);
and U29272 (N_29272,N_28515,N_28452);
nor U29273 (N_29273,N_28784,N_27845);
nand U29274 (N_29274,N_27631,N_28739);
and U29275 (N_29275,N_28776,N_28796);
or U29276 (N_29276,N_28504,N_28069);
nor U29277 (N_29277,N_27679,N_27951);
or U29278 (N_29278,N_28131,N_27651);
xor U29279 (N_29279,N_28780,N_28609);
nand U29280 (N_29280,N_28436,N_28314);
nand U29281 (N_29281,N_28123,N_28169);
xnor U29282 (N_29282,N_28553,N_28264);
nand U29283 (N_29283,N_27744,N_27778);
nor U29284 (N_29284,N_28106,N_28152);
xnor U29285 (N_29285,N_27727,N_27790);
or U29286 (N_29286,N_28468,N_28348);
xnor U29287 (N_29287,N_28240,N_28482);
nand U29288 (N_29288,N_28304,N_28540);
xnor U29289 (N_29289,N_27844,N_27637);
nor U29290 (N_29290,N_28143,N_28517);
nor U29291 (N_29291,N_27988,N_28313);
nand U29292 (N_29292,N_27940,N_28275);
xor U29293 (N_29293,N_28365,N_28084);
xnor U29294 (N_29294,N_28536,N_28664);
nand U29295 (N_29295,N_27945,N_28698);
xnor U29296 (N_29296,N_27616,N_28263);
and U29297 (N_29297,N_28400,N_28202);
or U29298 (N_29298,N_28104,N_27931);
nand U29299 (N_29299,N_28478,N_28509);
and U29300 (N_29300,N_28227,N_28561);
xnor U29301 (N_29301,N_28577,N_28707);
nand U29302 (N_29302,N_28608,N_28308);
or U29303 (N_29303,N_27775,N_27953);
and U29304 (N_29304,N_28181,N_28078);
and U29305 (N_29305,N_28384,N_27783);
nand U29306 (N_29306,N_28420,N_28620);
xor U29307 (N_29307,N_27892,N_28685);
nand U29308 (N_29308,N_27830,N_27625);
xor U29309 (N_29309,N_28380,N_28472);
nor U29310 (N_29310,N_27925,N_27735);
nand U29311 (N_29311,N_28397,N_27733);
xnor U29312 (N_29312,N_28496,N_27967);
xor U29313 (N_29313,N_28117,N_28604);
nor U29314 (N_29314,N_27802,N_28213);
xor U29315 (N_29315,N_28521,N_27671);
nor U29316 (N_29316,N_28082,N_28548);
nor U29317 (N_29317,N_28500,N_27721);
or U29318 (N_29318,N_28728,N_28049);
nand U29319 (N_29319,N_27921,N_27766);
and U29320 (N_29320,N_28442,N_28068);
or U29321 (N_29321,N_28499,N_27823);
nor U29322 (N_29322,N_28014,N_28342);
xnor U29323 (N_29323,N_27801,N_28660);
nor U29324 (N_29324,N_27958,N_27944);
and U29325 (N_29325,N_28363,N_28522);
nor U29326 (N_29326,N_27824,N_27833);
xnor U29327 (N_29327,N_28267,N_28731);
nor U29328 (N_29328,N_27722,N_27629);
nor U29329 (N_29329,N_28310,N_28727);
and U29330 (N_29330,N_28295,N_28233);
nand U29331 (N_29331,N_27710,N_28051);
or U29332 (N_29332,N_28701,N_28475);
or U29333 (N_29333,N_28080,N_28773);
nand U29334 (N_29334,N_28428,N_28720);
and U29335 (N_29335,N_28033,N_28191);
nand U29336 (N_29336,N_27785,N_28777);
and U29337 (N_29337,N_28469,N_28535);
nand U29338 (N_29338,N_28071,N_28630);
or U29339 (N_29339,N_27756,N_28297);
xnor U29340 (N_29340,N_28193,N_28575);
nand U29341 (N_29341,N_28098,N_28034);
or U29342 (N_29342,N_27626,N_28008);
or U29343 (N_29343,N_28218,N_28335);
nand U29344 (N_29344,N_28156,N_28354);
xor U29345 (N_29345,N_28013,N_28031);
and U29346 (N_29346,N_27669,N_27847);
or U29347 (N_29347,N_28287,N_28649);
nor U29348 (N_29348,N_28602,N_27700);
and U29349 (N_29349,N_27963,N_27699);
xnor U29350 (N_29350,N_27732,N_27860);
nand U29351 (N_29351,N_27632,N_28696);
nor U29352 (N_29352,N_28220,N_27820);
xor U29353 (N_29353,N_28699,N_28733);
nor U29354 (N_29354,N_28285,N_28294);
nand U29355 (N_29355,N_28405,N_28503);
xnor U29356 (N_29356,N_27850,N_28725);
and U29357 (N_29357,N_27767,N_27828);
and U29358 (N_29358,N_28357,N_28508);
and U29359 (N_29359,N_28717,N_28217);
nand U29360 (N_29360,N_28665,N_28019);
nor U29361 (N_29361,N_28542,N_27643);
nand U29362 (N_29362,N_27602,N_28681);
and U29363 (N_29363,N_28161,N_28261);
or U29364 (N_29364,N_28020,N_28756);
and U29365 (N_29365,N_27868,N_27619);
xor U29366 (N_29366,N_27666,N_27702);
nand U29367 (N_29367,N_28551,N_28388);
and U29368 (N_29368,N_28787,N_28641);
nor U29369 (N_29369,N_28345,N_28352);
or U29370 (N_29370,N_27714,N_28799);
and U29371 (N_29371,N_28016,N_28290);
nor U29372 (N_29372,N_28179,N_28300);
nand U29373 (N_29373,N_28307,N_27870);
nor U29374 (N_29374,N_28292,N_27750);
nand U29375 (N_29375,N_28677,N_28506);
nand U29376 (N_29376,N_27908,N_28334);
xor U29377 (N_29377,N_28771,N_28057);
xnor U29378 (N_29378,N_28702,N_27841);
and U29379 (N_29379,N_27879,N_28485);
nor U29380 (N_29380,N_28598,N_27607);
xnor U29381 (N_29381,N_27835,N_27869);
xnor U29382 (N_29382,N_28557,N_27914);
nor U29383 (N_29383,N_28372,N_28132);
xnor U29384 (N_29384,N_28158,N_28116);
nor U29385 (N_29385,N_27929,N_27760);
nor U29386 (N_29386,N_28306,N_28273);
nor U29387 (N_29387,N_28180,N_28128);
or U29388 (N_29388,N_28119,N_27973);
nor U29389 (N_29389,N_27603,N_28289);
xor U29390 (N_29390,N_28028,N_28534);
nor U29391 (N_29391,N_28501,N_28333);
xor U29392 (N_29392,N_27971,N_28321);
and U29393 (N_29393,N_28533,N_28541);
nor U29394 (N_29394,N_28555,N_27902);
and U29395 (N_29395,N_28635,N_28642);
nand U29396 (N_29396,N_27856,N_27983);
or U29397 (N_29397,N_27773,N_28072);
xor U29398 (N_29398,N_28351,N_27934);
and U29399 (N_29399,N_28429,N_28781);
xnor U29400 (N_29400,N_28261,N_28547);
and U29401 (N_29401,N_28746,N_27685);
and U29402 (N_29402,N_28270,N_27840);
nor U29403 (N_29403,N_28057,N_28779);
and U29404 (N_29404,N_27790,N_28240);
or U29405 (N_29405,N_27617,N_27782);
or U29406 (N_29406,N_28660,N_27641);
and U29407 (N_29407,N_28396,N_28578);
nand U29408 (N_29408,N_28085,N_28458);
nand U29409 (N_29409,N_27888,N_28288);
xnor U29410 (N_29410,N_28263,N_28018);
or U29411 (N_29411,N_27866,N_28161);
nand U29412 (N_29412,N_27616,N_28686);
or U29413 (N_29413,N_28678,N_28113);
nand U29414 (N_29414,N_27977,N_28240);
or U29415 (N_29415,N_27714,N_28761);
nand U29416 (N_29416,N_28645,N_27617);
and U29417 (N_29417,N_28682,N_28255);
nand U29418 (N_29418,N_28298,N_27709);
nor U29419 (N_29419,N_27739,N_28276);
nand U29420 (N_29420,N_27948,N_28789);
or U29421 (N_29421,N_27604,N_27900);
or U29422 (N_29422,N_28319,N_28735);
xnor U29423 (N_29423,N_27945,N_28387);
nor U29424 (N_29424,N_28611,N_27752);
or U29425 (N_29425,N_28618,N_27626);
and U29426 (N_29426,N_27711,N_28014);
or U29427 (N_29427,N_28609,N_28470);
and U29428 (N_29428,N_28045,N_28128);
and U29429 (N_29429,N_28214,N_27724);
nand U29430 (N_29430,N_28053,N_28204);
and U29431 (N_29431,N_28242,N_27878);
xor U29432 (N_29432,N_27824,N_28661);
nor U29433 (N_29433,N_28609,N_28583);
and U29434 (N_29434,N_27805,N_27843);
nor U29435 (N_29435,N_28081,N_28270);
xnor U29436 (N_29436,N_27884,N_28733);
nor U29437 (N_29437,N_28287,N_27878);
xnor U29438 (N_29438,N_27975,N_28066);
xnor U29439 (N_29439,N_28395,N_28132);
nor U29440 (N_29440,N_28357,N_28433);
nand U29441 (N_29441,N_28324,N_28555);
nand U29442 (N_29442,N_28026,N_28336);
or U29443 (N_29443,N_28280,N_27831);
nor U29444 (N_29444,N_28780,N_27966);
or U29445 (N_29445,N_27683,N_27740);
and U29446 (N_29446,N_27976,N_28663);
nand U29447 (N_29447,N_28527,N_27627);
xor U29448 (N_29448,N_28144,N_27926);
or U29449 (N_29449,N_28180,N_28386);
or U29450 (N_29450,N_27969,N_28310);
nor U29451 (N_29451,N_27633,N_28273);
xnor U29452 (N_29452,N_27815,N_27931);
and U29453 (N_29453,N_27954,N_27754);
or U29454 (N_29454,N_28135,N_28646);
nand U29455 (N_29455,N_28764,N_27892);
nor U29456 (N_29456,N_28225,N_27800);
nor U29457 (N_29457,N_27991,N_28105);
and U29458 (N_29458,N_27959,N_27703);
or U29459 (N_29459,N_28613,N_28349);
xnor U29460 (N_29460,N_28236,N_28385);
or U29461 (N_29461,N_28743,N_28787);
nor U29462 (N_29462,N_28545,N_28054);
xor U29463 (N_29463,N_28190,N_28726);
xor U29464 (N_29464,N_28661,N_28231);
xnor U29465 (N_29465,N_28391,N_28070);
nor U29466 (N_29466,N_27933,N_28562);
or U29467 (N_29467,N_27748,N_27747);
nor U29468 (N_29468,N_28086,N_28659);
and U29469 (N_29469,N_27611,N_28615);
nor U29470 (N_29470,N_27737,N_28751);
xor U29471 (N_29471,N_28489,N_27618);
and U29472 (N_29472,N_27725,N_27665);
and U29473 (N_29473,N_27742,N_27994);
nor U29474 (N_29474,N_27769,N_28328);
xnor U29475 (N_29475,N_27846,N_28530);
or U29476 (N_29476,N_28000,N_28376);
nand U29477 (N_29477,N_28042,N_28440);
nand U29478 (N_29478,N_27863,N_28707);
nor U29479 (N_29479,N_28683,N_28402);
or U29480 (N_29480,N_28599,N_27742);
and U29481 (N_29481,N_28703,N_28142);
and U29482 (N_29482,N_28370,N_27725);
and U29483 (N_29483,N_28517,N_27905);
nor U29484 (N_29484,N_28533,N_27788);
and U29485 (N_29485,N_28505,N_28610);
nand U29486 (N_29486,N_27900,N_27867);
or U29487 (N_29487,N_28539,N_28364);
nand U29488 (N_29488,N_27929,N_28010);
or U29489 (N_29489,N_28061,N_27745);
or U29490 (N_29490,N_27718,N_28391);
or U29491 (N_29491,N_27829,N_28630);
nand U29492 (N_29492,N_27634,N_28481);
and U29493 (N_29493,N_28750,N_28452);
nor U29494 (N_29494,N_28158,N_27660);
and U29495 (N_29495,N_27660,N_27949);
or U29496 (N_29496,N_28370,N_28186);
nor U29497 (N_29497,N_28449,N_28511);
xnor U29498 (N_29498,N_27660,N_27809);
nand U29499 (N_29499,N_27741,N_28084);
nand U29500 (N_29500,N_28193,N_28478);
or U29501 (N_29501,N_28552,N_28799);
or U29502 (N_29502,N_27691,N_27929);
nor U29503 (N_29503,N_28775,N_28428);
xnor U29504 (N_29504,N_28008,N_28662);
or U29505 (N_29505,N_28276,N_27876);
nand U29506 (N_29506,N_28401,N_28793);
nor U29507 (N_29507,N_28595,N_28658);
nor U29508 (N_29508,N_28322,N_28672);
nor U29509 (N_29509,N_28421,N_28578);
nor U29510 (N_29510,N_28241,N_28672);
and U29511 (N_29511,N_27844,N_28426);
and U29512 (N_29512,N_27835,N_28713);
and U29513 (N_29513,N_28424,N_28012);
nor U29514 (N_29514,N_28543,N_28651);
or U29515 (N_29515,N_28706,N_27640);
and U29516 (N_29516,N_27915,N_28361);
and U29517 (N_29517,N_27989,N_28204);
nor U29518 (N_29518,N_28347,N_27785);
or U29519 (N_29519,N_28175,N_27739);
nor U29520 (N_29520,N_28377,N_27963);
nand U29521 (N_29521,N_28424,N_28535);
or U29522 (N_29522,N_28758,N_27624);
or U29523 (N_29523,N_28347,N_28669);
xnor U29524 (N_29524,N_28379,N_27797);
and U29525 (N_29525,N_28749,N_28280);
and U29526 (N_29526,N_27777,N_28421);
nor U29527 (N_29527,N_28181,N_28774);
nand U29528 (N_29528,N_28530,N_28094);
xor U29529 (N_29529,N_28679,N_28796);
nor U29530 (N_29530,N_28717,N_27819);
and U29531 (N_29531,N_28077,N_27679);
and U29532 (N_29532,N_28259,N_28645);
and U29533 (N_29533,N_28390,N_28481);
and U29534 (N_29534,N_28576,N_27821);
nand U29535 (N_29535,N_28587,N_28128);
nor U29536 (N_29536,N_28492,N_27718);
and U29537 (N_29537,N_28502,N_28032);
nand U29538 (N_29538,N_27938,N_27637);
and U29539 (N_29539,N_27720,N_28174);
xnor U29540 (N_29540,N_28417,N_27902);
nand U29541 (N_29541,N_28459,N_27976);
and U29542 (N_29542,N_28241,N_28748);
xnor U29543 (N_29543,N_27882,N_28056);
and U29544 (N_29544,N_28789,N_27810);
nor U29545 (N_29545,N_27634,N_27887);
xor U29546 (N_29546,N_27612,N_28682);
nor U29547 (N_29547,N_28690,N_28794);
and U29548 (N_29548,N_27678,N_28522);
nor U29549 (N_29549,N_28269,N_28724);
nor U29550 (N_29550,N_28057,N_27708);
nand U29551 (N_29551,N_28088,N_28451);
or U29552 (N_29552,N_28681,N_28776);
xor U29553 (N_29553,N_28472,N_28560);
or U29554 (N_29554,N_28694,N_27610);
nor U29555 (N_29555,N_28265,N_27613);
and U29556 (N_29556,N_28007,N_28365);
nor U29557 (N_29557,N_27664,N_27611);
nand U29558 (N_29558,N_28004,N_28229);
nand U29559 (N_29559,N_27988,N_28294);
or U29560 (N_29560,N_28062,N_27846);
nand U29561 (N_29561,N_27631,N_28799);
or U29562 (N_29562,N_27601,N_27956);
nor U29563 (N_29563,N_27873,N_27772);
and U29564 (N_29564,N_28763,N_28459);
nor U29565 (N_29565,N_28002,N_28147);
nand U29566 (N_29566,N_27723,N_27796);
or U29567 (N_29567,N_28139,N_27700);
and U29568 (N_29568,N_28337,N_28032);
or U29569 (N_29569,N_27930,N_27868);
xor U29570 (N_29570,N_28546,N_28207);
and U29571 (N_29571,N_28393,N_27923);
or U29572 (N_29572,N_28379,N_27858);
nor U29573 (N_29573,N_28755,N_27674);
xor U29574 (N_29574,N_28784,N_28072);
nor U29575 (N_29575,N_28248,N_28429);
or U29576 (N_29576,N_28659,N_28411);
nand U29577 (N_29577,N_27828,N_28308);
xor U29578 (N_29578,N_27938,N_28123);
xor U29579 (N_29579,N_28717,N_28620);
or U29580 (N_29580,N_27685,N_28526);
or U29581 (N_29581,N_27633,N_28568);
nand U29582 (N_29582,N_28050,N_27887);
nand U29583 (N_29583,N_27963,N_28359);
nor U29584 (N_29584,N_28290,N_28303);
nand U29585 (N_29585,N_27620,N_28799);
and U29586 (N_29586,N_28101,N_27910);
nor U29587 (N_29587,N_27605,N_27948);
and U29588 (N_29588,N_28670,N_28744);
nor U29589 (N_29589,N_27992,N_27982);
nor U29590 (N_29590,N_28628,N_27628);
nor U29591 (N_29591,N_28722,N_28781);
nand U29592 (N_29592,N_27869,N_27986);
nor U29593 (N_29593,N_28784,N_28684);
xnor U29594 (N_29594,N_28594,N_27608);
xor U29595 (N_29595,N_27652,N_27720);
or U29596 (N_29596,N_28384,N_27642);
or U29597 (N_29597,N_28071,N_28255);
and U29598 (N_29598,N_28404,N_28150);
nand U29599 (N_29599,N_28404,N_28613);
xor U29600 (N_29600,N_28521,N_27919);
nand U29601 (N_29601,N_27607,N_28005);
and U29602 (N_29602,N_27730,N_27744);
nand U29603 (N_29603,N_28648,N_28312);
nor U29604 (N_29604,N_28095,N_28665);
and U29605 (N_29605,N_28079,N_27702);
and U29606 (N_29606,N_28190,N_27790);
xnor U29607 (N_29607,N_28172,N_27607);
or U29608 (N_29608,N_28095,N_28635);
or U29609 (N_29609,N_27879,N_28677);
xnor U29610 (N_29610,N_28088,N_28703);
or U29611 (N_29611,N_28688,N_28764);
nor U29612 (N_29612,N_27705,N_28219);
nand U29613 (N_29613,N_28209,N_27625);
xor U29614 (N_29614,N_28056,N_28245);
or U29615 (N_29615,N_27720,N_28480);
and U29616 (N_29616,N_28701,N_28426);
and U29617 (N_29617,N_27846,N_28137);
and U29618 (N_29618,N_27834,N_28663);
xnor U29619 (N_29619,N_28442,N_28484);
xnor U29620 (N_29620,N_28543,N_27957);
nor U29621 (N_29621,N_28172,N_28388);
xnor U29622 (N_29622,N_28690,N_27854);
nor U29623 (N_29623,N_28201,N_28601);
nor U29624 (N_29624,N_28014,N_27985);
nand U29625 (N_29625,N_28433,N_28463);
nand U29626 (N_29626,N_28415,N_28607);
nand U29627 (N_29627,N_27931,N_28224);
nor U29628 (N_29628,N_28790,N_28430);
or U29629 (N_29629,N_28490,N_27754);
or U29630 (N_29630,N_27907,N_28361);
and U29631 (N_29631,N_28597,N_27873);
and U29632 (N_29632,N_27639,N_27651);
xor U29633 (N_29633,N_28298,N_28023);
nand U29634 (N_29634,N_27863,N_27833);
or U29635 (N_29635,N_28235,N_28713);
nor U29636 (N_29636,N_28053,N_28762);
nor U29637 (N_29637,N_28248,N_27779);
nor U29638 (N_29638,N_27863,N_27705);
nor U29639 (N_29639,N_28698,N_28275);
and U29640 (N_29640,N_28157,N_28275);
or U29641 (N_29641,N_28544,N_28411);
nor U29642 (N_29642,N_28193,N_28146);
xnor U29643 (N_29643,N_28039,N_28682);
nand U29644 (N_29644,N_28329,N_28771);
nand U29645 (N_29645,N_28608,N_28208);
and U29646 (N_29646,N_27967,N_28106);
or U29647 (N_29647,N_28062,N_27904);
and U29648 (N_29648,N_27752,N_27625);
nand U29649 (N_29649,N_28120,N_27865);
nand U29650 (N_29650,N_28795,N_27853);
or U29651 (N_29651,N_27789,N_28695);
xor U29652 (N_29652,N_28208,N_27727);
and U29653 (N_29653,N_27659,N_27788);
nor U29654 (N_29654,N_28694,N_28668);
or U29655 (N_29655,N_28491,N_27932);
and U29656 (N_29656,N_28786,N_27779);
and U29657 (N_29657,N_28406,N_27972);
nand U29658 (N_29658,N_27859,N_28356);
nor U29659 (N_29659,N_28764,N_28398);
and U29660 (N_29660,N_27609,N_28043);
xnor U29661 (N_29661,N_27970,N_28017);
nor U29662 (N_29662,N_27711,N_27719);
or U29663 (N_29663,N_28289,N_27869);
and U29664 (N_29664,N_27980,N_27964);
and U29665 (N_29665,N_28036,N_28653);
nand U29666 (N_29666,N_27935,N_27609);
nand U29667 (N_29667,N_28523,N_28376);
nor U29668 (N_29668,N_28113,N_27807);
or U29669 (N_29669,N_28262,N_28686);
xnor U29670 (N_29670,N_28352,N_28630);
and U29671 (N_29671,N_28366,N_28573);
nor U29672 (N_29672,N_28103,N_28033);
nor U29673 (N_29673,N_28325,N_28386);
or U29674 (N_29674,N_27697,N_27911);
and U29675 (N_29675,N_28348,N_28546);
and U29676 (N_29676,N_28357,N_28527);
nor U29677 (N_29677,N_28294,N_28721);
xor U29678 (N_29678,N_27997,N_28769);
or U29679 (N_29679,N_28066,N_28663);
and U29680 (N_29680,N_28104,N_27921);
and U29681 (N_29681,N_28590,N_28049);
and U29682 (N_29682,N_28319,N_28731);
nand U29683 (N_29683,N_27745,N_28364);
xor U29684 (N_29684,N_27984,N_27602);
xnor U29685 (N_29685,N_28077,N_28644);
xnor U29686 (N_29686,N_28439,N_28489);
or U29687 (N_29687,N_28455,N_28359);
nor U29688 (N_29688,N_27714,N_27685);
or U29689 (N_29689,N_27770,N_28286);
and U29690 (N_29690,N_28539,N_28717);
nand U29691 (N_29691,N_27949,N_28385);
or U29692 (N_29692,N_27908,N_27912);
nand U29693 (N_29693,N_27631,N_28169);
nor U29694 (N_29694,N_28020,N_28116);
or U29695 (N_29695,N_27662,N_27918);
or U29696 (N_29696,N_27670,N_28501);
or U29697 (N_29697,N_28348,N_27828);
and U29698 (N_29698,N_27819,N_27742);
or U29699 (N_29699,N_28699,N_27868);
and U29700 (N_29700,N_28282,N_28336);
xor U29701 (N_29701,N_27778,N_27919);
or U29702 (N_29702,N_28709,N_27962);
xnor U29703 (N_29703,N_28266,N_27977);
nand U29704 (N_29704,N_27701,N_27613);
or U29705 (N_29705,N_28265,N_28225);
and U29706 (N_29706,N_28354,N_28064);
nand U29707 (N_29707,N_28133,N_27786);
nor U29708 (N_29708,N_28090,N_28064);
and U29709 (N_29709,N_28440,N_28712);
and U29710 (N_29710,N_28242,N_28106);
xnor U29711 (N_29711,N_27628,N_28055);
xor U29712 (N_29712,N_27836,N_28598);
or U29713 (N_29713,N_28040,N_27640);
nor U29714 (N_29714,N_27707,N_28555);
xor U29715 (N_29715,N_28794,N_28605);
and U29716 (N_29716,N_28158,N_27621);
xnor U29717 (N_29717,N_28685,N_28630);
xor U29718 (N_29718,N_27888,N_27672);
or U29719 (N_29719,N_27822,N_28013);
xnor U29720 (N_29720,N_27920,N_28361);
or U29721 (N_29721,N_28717,N_28418);
nor U29722 (N_29722,N_28077,N_28262);
xnor U29723 (N_29723,N_27780,N_28028);
nor U29724 (N_29724,N_28695,N_27913);
xor U29725 (N_29725,N_28663,N_28436);
xnor U29726 (N_29726,N_28137,N_27840);
xor U29727 (N_29727,N_28718,N_27707);
xnor U29728 (N_29728,N_28587,N_28345);
nand U29729 (N_29729,N_28723,N_28555);
nor U29730 (N_29730,N_27684,N_28672);
nand U29731 (N_29731,N_28055,N_27901);
nor U29732 (N_29732,N_28129,N_28025);
nor U29733 (N_29733,N_27879,N_27777);
or U29734 (N_29734,N_28235,N_27898);
and U29735 (N_29735,N_28531,N_28546);
nor U29736 (N_29736,N_27831,N_27689);
nand U29737 (N_29737,N_28297,N_28509);
and U29738 (N_29738,N_27789,N_28739);
nand U29739 (N_29739,N_27910,N_28718);
nor U29740 (N_29740,N_28689,N_28779);
or U29741 (N_29741,N_28075,N_28380);
nand U29742 (N_29742,N_28187,N_27816);
nand U29743 (N_29743,N_28282,N_28322);
nand U29744 (N_29744,N_28410,N_27765);
or U29745 (N_29745,N_27974,N_28351);
and U29746 (N_29746,N_28350,N_27834);
or U29747 (N_29747,N_28602,N_27808);
nand U29748 (N_29748,N_27941,N_27692);
xor U29749 (N_29749,N_27781,N_27915);
and U29750 (N_29750,N_27890,N_28713);
or U29751 (N_29751,N_28482,N_27850);
nand U29752 (N_29752,N_28734,N_28030);
nor U29753 (N_29753,N_28292,N_28662);
nor U29754 (N_29754,N_28679,N_28254);
nor U29755 (N_29755,N_28606,N_27659);
nor U29756 (N_29756,N_27809,N_27865);
nand U29757 (N_29757,N_28780,N_28301);
nand U29758 (N_29758,N_28788,N_27674);
and U29759 (N_29759,N_27668,N_27627);
nand U29760 (N_29760,N_27775,N_27674);
nand U29761 (N_29761,N_28040,N_28659);
xnor U29762 (N_29762,N_28048,N_28293);
nor U29763 (N_29763,N_28470,N_27866);
xor U29764 (N_29764,N_27670,N_27687);
xor U29765 (N_29765,N_27683,N_28695);
xnor U29766 (N_29766,N_28394,N_28352);
nand U29767 (N_29767,N_27681,N_28351);
or U29768 (N_29768,N_27959,N_28173);
nor U29769 (N_29769,N_28188,N_27787);
xor U29770 (N_29770,N_28424,N_28761);
xnor U29771 (N_29771,N_27896,N_27750);
nor U29772 (N_29772,N_28152,N_27819);
nand U29773 (N_29773,N_28149,N_28501);
or U29774 (N_29774,N_28503,N_28067);
or U29775 (N_29775,N_28056,N_27910);
nand U29776 (N_29776,N_28087,N_28503);
and U29777 (N_29777,N_28631,N_28436);
xor U29778 (N_29778,N_28358,N_28131);
nand U29779 (N_29779,N_28163,N_28107);
and U29780 (N_29780,N_28477,N_28609);
or U29781 (N_29781,N_28201,N_27938);
and U29782 (N_29782,N_27820,N_27947);
xor U29783 (N_29783,N_28487,N_28153);
and U29784 (N_29784,N_27880,N_27810);
and U29785 (N_29785,N_28774,N_28172);
or U29786 (N_29786,N_28323,N_27642);
or U29787 (N_29787,N_28437,N_28304);
or U29788 (N_29788,N_28430,N_27964);
or U29789 (N_29789,N_28579,N_27929);
nand U29790 (N_29790,N_28107,N_28619);
and U29791 (N_29791,N_28140,N_28736);
nor U29792 (N_29792,N_28381,N_28439);
xnor U29793 (N_29793,N_27915,N_27772);
and U29794 (N_29794,N_27681,N_28642);
and U29795 (N_29795,N_27636,N_27958);
and U29796 (N_29796,N_28511,N_27914);
and U29797 (N_29797,N_28685,N_28452);
xnor U29798 (N_29798,N_27756,N_28584);
and U29799 (N_29799,N_28656,N_28713);
nor U29800 (N_29800,N_28637,N_28372);
xor U29801 (N_29801,N_28531,N_28699);
nand U29802 (N_29802,N_27687,N_28122);
nor U29803 (N_29803,N_28786,N_28323);
nor U29804 (N_29804,N_28097,N_27709);
and U29805 (N_29805,N_27678,N_27673);
or U29806 (N_29806,N_28347,N_27794);
nand U29807 (N_29807,N_27688,N_28070);
and U29808 (N_29808,N_28086,N_28740);
and U29809 (N_29809,N_28024,N_28775);
xnor U29810 (N_29810,N_27872,N_27827);
or U29811 (N_29811,N_28380,N_27986);
nor U29812 (N_29812,N_28565,N_28410);
nand U29813 (N_29813,N_28167,N_28147);
nor U29814 (N_29814,N_28297,N_28784);
and U29815 (N_29815,N_27916,N_27621);
nand U29816 (N_29816,N_28516,N_28357);
or U29817 (N_29817,N_28566,N_28117);
nand U29818 (N_29818,N_28103,N_28024);
xnor U29819 (N_29819,N_28162,N_28434);
or U29820 (N_29820,N_27999,N_28378);
xor U29821 (N_29821,N_28357,N_27790);
xnor U29822 (N_29822,N_28319,N_28231);
nand U29823 (N_29823,N_28236,N_28185);
nand U29824 (N_29824,N_27806,N_28516);
and U29825 (N_29825,N_28684,N_28793);
nor U29826 (N_29826,N_27754,N_28423);
or U29827 (N_29827,N_28117,N_28056);
xnor U29828 (N_29828,N_28714,N_28777);
and U29829 (N_29829,N_28385,N_28747);
nand U29830 (N_29830,N_27998,N_27913);
xor U29831 (N_29831,N_28421,N_28727);
xnor U29832 (N_29832,N_27653,N_28725);
nand U29833 (N_29833,N_28167,N_28511);
or U29834 (N_29834,N_27653,N_28015);
or U29835 (N_29835,N_28406,N_27601);
nor U29836 (N_29836,N_28588,N_28501);
and U29837 (N_29837,N_28113,N_28284);
nor U29838 (N_29838,N_27659,N_27776);
xor U29839 (N_29839,N_28224,N_27605);
xor U29840 (N_29840,N_28040,N_27938);
and U29841 (N_29841,N_27747,N_28272);
nor U29842 (N_29842,N_27778,N_28287);
and U29843 (N_29843,N_28462,N_27617);
and U29844 (N_29844,N_28677,N_28478);
nor U29845 (N_29845,N_27714,N_27859);
nand U29846 (N_29846,N_28127,N_28384);
nand U29847 (N_29847,N_28770,N_27712);
nand U29848 (N_29848,N_28107,N_27667);
nor U29849 (N_29849,N_28244,N_28600);
xnor U29850 (N_29850,N_27739,N_28068);
or U29851 (N_29851,N_28393,N_27937);
or U29852 (N_29852,N_28439,N_28284);
nand U29853 (N_29853,N_28203,N_28121);
nor U29854 (N_29854,N_28735,N_28366);
nor U29855 (N_29855,N_28409,N_28559);
nor U29856 (N_29856,N_28050,N_28065);
xnor U29857 (N_29857,N_28160,N_27844);
nor U29858 (N_29858,N_28113,N_27834);
xor U29859 (N_29859,N_27763,N_28535);
nor U29860 (N_29860,N_28141,N_27746);
xnor U29861 (N_29861,N_28725,N_27819);
nor U29862 (N_29862,N_27841,N_28687);
nor U29863 (N_29863,N_28015,N_27768);
or U29864 (N_29864,N_28446,N_27967);
or U29865 (N_29865,N_28798,N_27982);
xor U29866 (N_29866,N_28688,N_28046);
xor U29867 (N_29867,N_27857,N_28507);
and U29868 (N_29868,N_28794,N_27626);
or U29869 (N_29869,N_28438,N_27820);
xnor U29870 (N_29870,N_27749,N_27743);
or U29871 (N_29871,N_28091,N_28494);
nor U29872 (N_29872,N_27903,N_27736);
and U29873 (N_29873,N_28713,N_27927);
and U29874 (N_29874,N_28330,N_28449);
nor U29875 (N_29875,N_28400,N_27722);
xor U29876 (N_29876,N_28185,N_28600);
and U29877 (N_29877,N_28185,N_27715);
nor U29878 (N_29878,N_28254,N_27772);
and U29879 (N_29879,N_28597,N_28117);
or U29880 (N_29880,N_28599,N_27995);
xnor U29881 (N_29881,N_28095,N_27636);
nand U29882 (N_29882,N_28000,N_27687);
and U29883 (N_29883,N_28213,N_28357);
nand U29884 (N_29884,N_27899,N_27754);
or U29885 (N_29885,N_28138,N_27899);
xnor U29886 (N_29886,N_28249,N_28662);
and U29887 (N_29887,N_28271,N_27648);
nor U29888 (N_29888,N_27849,N_28532);
xnor U29889 (N_29889,N_27648,N_28434);
nor U29890 (N_29890,N_28723,N_28119);
xnor U29891 (N_29891,N_28635,N_28063);
or U29892 (N_29892,N_28560,N_28392);
xnor U29893 (N_29893,N_28192,N_27636);
nor U29894 (N_29894,N_28009,N_28398);
and U29895 (N_29895,N_28452,N_28009);
nor U29896 (N_29896,N_28204,N_27847);
nand U29897 (N_29897,N_27875,N_28642);
nor U29898 (N_29898,N_27768,N_28128);
nand U29899 (N_29899,N_27924,N_28423);
nor U29900 (N_29900,N_28596,N_28746);
xnor U29901 (N_29901,N_28449,N_27804);
or U29902 (N_29902,N_27890,N_28551);
xor U29903 (N_29903,N_28281,N_28254);
xor U29904 (N_29904,N_28258,N_27623);
xnor U29905 (N_29905,N_28617,N_28132);
xor U29906 (N_29906,N_28436,N_28767);
xnor U29907 (N_29907,N_28213,N_28764);
xnor U29908 (N_29908,N_28531,N_27828);
and U29909 (N_29909,N_27880,N_28604);
or U29910 (N_29910,N_27729,N_28387);
nand U29911 (N_29911,N_27661,N_28108);
and U29912 (N_29912,N_28420,N_28377);
xor U29913 (N_29913,N_28770,N_28237);
nor U29914 (N_29914,N_28696,N_27857);
or U29915 (N_29915,N_28228,N_28712);
nor U29916 (N_29916,N_28469,N_28302);
and U29917 (N_29917,N_28296,N_28021);
nand U29918 (N_29918,N_28608,N_28553);
nand U29919 (N_29919,N_28582,N_28310);
nand U29920 (N_29920,N_27749,N_27684);
and U29921 (N_29921,N_28036,N_28510);
or U29922 (N_29922,N_27883,N_28677);
nand U29923 (N_29923,N_28689,N_28008);
nor U29924 (N_29924,N_28241,N_28319);
nor U29925 (N_29925,N_28773,N_27730);
xor U29926 (N_29926,N_27618,N_28663);
or U29927 (N_29927,N_27812,N_28772);
nand U29928 (N_29928,N_28364,N_27950);
nor U29929 (N_29929,N_28752,N_28736);
nand U29930 (N_29930,N_28548,N_28345);
or U29931 (N_29931,N_27848,N_28167);
or U29932 (N_29932,N_28336,N_27626);
nor U29933 (N_29933,N_28654,N_28253);
or U29934 (N_29934,N_28152,N_27718);
nor U29935 (N_29935,N_27807,N_27747);
nand U29936 (N_29936,N_28545,N_27821);
xnor U29937 (N_29937,N_27612,N_28746);
and U29938 (N_29938,N_28316,N_27733);
nor U29939 (N_29939,N_27658,N_28482);
nand U29940 (N_29940,N_27779,N_27802);
nor U29941 (N_29941,N_28285,N_28547);
and U29942 (N_29942,N_27750,N_28091);
and U29943 (N_29943,N_28114,N_27912);
nor U29944 (N_29944,N_28399,N_28559);
or U29945 (N_29945,N_27801,N_28670);
xor U29946 (N_29946,N_28460,N_28661);
nand U29947 (N_29947,N_28164,N_27655);
xnor U29948 (N_29948,N_27738,N_28549);
nor U29949 (N_29949,N_28139,N_27844);
or U29950 (N_29950,N_27718,N_27888);
xor U29951 (N_29951,N_28048,N_27660);
and U29952 (N_29952,N_28045,N_28760);
xnor U29953 (N_29953,N_28347,N_28298);
and U29954 (N_29954,N_28327,N_28548);
xor U29955 (N_29955,N_27974,N_28550);
nand U29956 (N_29956,N_28142,N_28182);
nand U29957 (N_29957,N_27925,N_28552);
nand U29958 (N_29958,N_28279,N_28281);
or U29959 (N_29959,N_27845,N_28542);
nand U29960 (N_29960,N_28652,N_27842);
or U29961 (N_29961,N_28535,N_28063);
and U29962 (N_29962,N_27911,N_28391);
nor U29963 (N_29963,N_28170,N_28041);
nand U29964 (N_29964,N_28095,N_27714);
xor U29965 (N_29965,N_28019,N_28243);
xor U29966 (N_29966,N_28518,N_27616);
nand U29967 (N_29967,N_28514,N_27887);
or U29968 (N_29968,N_28796,N_28031);
or U29969 (N_29969,N_28120,N_28787);
and U29970 (N_29970,N_28422,N_28318);
nor U29971 (N_29971,N_28076,N_28263);
nand U29972 (N_29972,N_27713,N_28799);
and U29973 (N_29973,N_28026,N_27991);
nor U29974 (N_29974,N_28463,N_28371);
xnor U29975 (N_29975,N_28770,N_28631);
nor U29976 (N_29976,N_28130,N_28314);
and U29977 (N_29977,N_28737,N_28722);
xor U29978 (N_29978,N_28257,N_28456);
nand U29979 (N_29979,N_27628,N_28468);
or U29980 (N_29980,N_27997,N_28300);
or U29981 (N_29981,N_28025,N_27849);
nor U29982 (N_29982,N_27911,N_28452);
nor U29983 (N_29983,N_28156,N_28394);
xor U29984 (N_29984,N_28363,N_27964);
or U29985 (N_29985,N_28719,N_28569);
xnor U29986 (N_29986,N_28594,N_27778);
nor U29987 (N_29987,N_28593,N_27628);
nand U29988 (N_29988,N_28013,N_28678);
and U29989 (N_29989,N_27797,N_28742);
or U29990 (N_29990,N_28164,N_27872);
xor U29991 (N_29991,N_28031,N_28133);
nor U29992 (N_29992,N_27893,N_28313);
nor U29993 (N_29993,N_28176,N_28775);
xor U29994 (N_29994,N_27896,N_27997);
or U29995 (N_29995,N_28536,N_27715);
nand U29996 (N_29996,N_27848,N_27847);
or U29997 (N_29997,N_27927,N_27935);
and U29998 (N_29998,N_28614,N_28751);
or U29999 (N_29999,N_28013,N_27601);
xnor UO_0 (O_0,N_29022,N_29904);
nand UO_1 (O_1,N_29076,N_29687);
xor UO_2 (O_2,N_29034,N_28886);
xnor UO_3 (O_3,N_29423,N_29221);
nor UO_4 (O_4,N_28931,N_28838);
nand UO_5 (O_5,N_29421,N_29878);
nand UO_6 (O_6,N_28858,N_29734);
nor UO_7 (O_7,N_29648,N_29325);
nor UO_8 (O_8,N_29066,N_29260);
and UO_9 (O_9,N_28817,N_29144);
nor UO_10 (O_10,N_29282,N_28910);
nand UO_11 (O_11,N_29104,N_29015);
and UO_12 (O_12,N_29250,N_28881);
nand UO_13 (O_13,N_29661,N_29458);
nor UO_14 (O_14,N_29120,N_29197);
nor UO_15 (O_15,N_29431,N_29061);
nor UO_16 (O_16,N_29702,N_29227);
or UO_17 (O_17,N_29683,N_28875);
nor UO_18 (O_18,N_28959,N_29566);
and UO_19 (O_19,N_29241,N_29742);
nor UO_20 (O_20,N_29289,N_29910);
xor UO_21 (O_21,N_28861,N_29259);
or UO_22 (O_22,N_28946,N_28936);
and UO_23 (O_23,N_29943,N_29272);
nor UO_24 (O_24,N_29396,N_29494);
or UO_25 (O_25,N_29643,N_29845);
nand UO_26 (O_26,N_28970,N_29997);
nor UO_27 (O_27,N_29003,N_29575);
and UO_28 (O_28,N_29803,N_29715);
nand UO_29 (O_29,N_28884,N_28960);
nor UO_30 (O_30,N_29211,N_29814);
and UO_31 (O_31,N_29758,N_29453);
xnor UO_32 (O_32,N_28808,N_29649);
xor UO_33 (O_33,N_29491,N_29021);
and UO_34 (O_34,N_29417,N_28978);
and UO_35 (O_35,N_29657,N_29085);
xnor UO_36 (O_36,N_28816,N_29502);
or UO_37 (O_37,N_29306,N_29794);
and UO_38 (O_38,N_28991,N_29834);
xor UO_39 (O_39,N_29969,N_29437);
and UO_40 (O_40,N_28871,N_29865);
and UO_41 (O_41,N_29596,N_28963);
xor UO_42 (O_42,N_29757,N_29674);
xnor UO_43 (O_43,N_29372,N_29941);
and UO_44 (O_44,N_29179,N_29716);
or UO_45 (O_45,N_29462,N_29040);
nor UO_46 (O_46,N_29949,N_29217);
nand UO_47 (O_47,N_29778,N_29813);
nand UO_48 (O_48,N_29083,N_29070);
nor UO_49 (O_49,N_29473,N_29956);
and UO_50 (O_50,N_29307,N_29212);
nor UO_51 (O_51,N_29351,N_29882);
xnor UO_52 (O_52,N_29712,N_29979);
nand UO_53 (O_53,N_29917,N_29350);
nor UO_54 (O_54,N_29189,N_29831);
nand UO_55 (O_55,N_29750,N_29441);
and UO_56 (O_56,N_29428,N_29369);
or UO_57 (O_57,N_29493,N_29581);
or UO_58 (O_58,N_29014,N_28919);
and UO_59 (O_59,N_29490,N_29515);
and UO_60 (O_60,N_29989,N_29311);
and UO_61 (O_61,N_29435,N_29377);
nand UO_62 (O_62,N_29353,N_29746);
nand UO_63 (O_63,N_29592,N_29165);
nor UO_64 (O_64,N_29568,N_29467);
nor UO_65 (O_65,N_29129,N_29113);
xnor UO_66 (O_66,N_28865,N_28958);
nor UO_67 (O_67,N_29169,N_29535);
nor UO_68 (O_68,N_29001,N_29516);
and UO_69 (O_69,N_28940,N_29761);
or UO_70 (O_70,N_29864,N_29608);
xnor UO_71 (O_71,N_29810,N_29247);
nand UO_72 (O_72,N_29151,N_29457);
or UO_73 (O_73,N_29265,N_29549);
and UO_74 (O_74,N_29118,N_29704);
and UO_75 (O_75,N_29237,N_29642);
and UO_76 (O_76,N_29853,N_29578);
xnor UO_77 (O_77,N_29287,N_29090);
nor UO_78 (O_78,N_29631,N_29593);
and UO_79 (O_79,N_29496,N_29769);
or UO_80 (O_80,N_29278,N_29116);
xnor UO_81 (O_81,N_29006,N_29470);
nor UO_82 (O_82,N_29330,N_29536);
or UO_83 (O_83,N_29112,N_29459);
nor UO_84 (O_84,N_29286,N_29824);
nand UO_85 (O_85,N_29662,N_29400);
nor UO_86 (O_86,N_29986,N_29929);
and UO_87 (O_87,N_29542,N_29737);
nor UO_88 (O_88,N_29889,N_29861);
or UO_89 (O_89,N_28918,N_29655);
or UO_90 (O_90,N_29206,N_29921);
xnor UO_91 (O_91,N_29092,N_29378);
xnor UO_92 (O_92,N_29362,N_29345);
and UO_93 (O_93,N_29302,N_29646);
or UO_94 (O_94,N_29045,N_29869);
xnor UO_95 (O_95,N_29572,N_29830);
nand UO_96 (O_96,N_29589,N_29177);
and UO_97 (O_97,N_28802,N_29952);
nand UO_98 (O_98,N_29360,N_29105);
nor UO_99 (O_99,N_29859,N_29768);
and UO_100 (O_100,N_29042,N_29312);
nor UO_101 (O_101,N_29366,N_29276);
and UO_102 (O_102,N_29140,N_28995);
and UO_103 (O_103,N_29897,N_28899);
nor UO_104 (O_104,N_29298,N_29318);
or UO_105 (O_105,N_29765,N_28992);
nor UO_106 (O_106,N_29053,N_28925);
and UO_107 (O_107,N_29398,N_29392);
and UO_108 (O_108,N_28880,N_29275);
or UO_109 (O_109,N_29624,N_29680);
nand UO_110 (O_110,N_29681,N_28862);
nand UO_111 (O_111,N_29843,N_29590);
and UO_112 (O_112,N_28806,N_29797);
or UO_113 (O_113,N_29444,N_29770);
nor UO_114 (O_114,N_29044,N_29163);
xnor UO_115 (O_115,N_29072,N_29766);
and UO_116 (O_116,N_29503,N_28869);
nor UO_117 (O_117,N_29037,N_29464);
nand UO_118 (O_118,N_29628,N_29297);
or UO_119 (O_119,N_29841,N_29429);
nand UO_120 (O_120,N_28945,N_29415);
or UO_121 (O_121,N_28801,N_29786);
nand UO_122 (O_122,N_29548,N_29709);
or UO_123 (O_123,N_29605,N_29847);
xor UO_124 (O_124,N_29139,N_29574);
or UO_125 (O_125,N_29625,N_29263);
nand UO_126 (O_126,N_29973,N_29356);
nand UO_127 (O_127,N_29521,N_29051);
nand UO_128 (O_128,N_29594,N_29495);
and UO_129 (O_129,N_28850,N_29501);
nand UO_130 (O_130,N_29075,N_29907);
or UO_131 (O_131,N_29915,N_28812);
xor UO_132 (O_132,N_29065,N_29252);
and UO_133 (O_133,N_29448,N_29077);
nor UO_134 (O_134,N_29736,N_29422);
or UO_135 (O_135,N_28965,N_29887);
nand UO_136 (O_136,N_28878,N_29695);
xor UO_137 (O_137,N_28897,N_29000);
xnor UO_138 (O_138,N_28906,N_29122);
xor UO_139 (O_139,N_28944,N_29023);
nand UO_140 (O_140,N_29980,N_29520);
nor UO_141 (O_141,N_29955,N_28926);
or UO_142 (O_142,N_29762,N_29792);
xnor UO_143 (O_143,N_29425,N_29328);
or UO_144 (O_144,N_28819,N_29175);
nor UO_145 (O_145,N_29722,N_29050);
xnor UO_146 (O_146,N_28962,N_29101);
xnor UO_147 (O_147,N_29771,N_28939);
nand UO_148 (O_148,N_29898,N_28997);
nor UO_149 (O_149,N_29570,N_29086);
or UO_150 (O_150,N_29799,N_29998);
or UO_151 (O_151,N_28948,N_29508);
or UO_152 (O_152,N_28905,N_29403);
and UO_153 (O_153,N_29653,N_29229);
and UO_154 (O_154,N_29127,N_29760);
xor UO_155 (O_155,N_29303,N_28985);
nand UO_156 (O_156,N_29759,N_29510);
xor UO_157 (O_157,N_29947,N_29942);
nor UO_158 (O_158,N_29851,N_29296);
or UO_159 (O_159,N_29767,N_29513);
or UO_160 (O_160,N_29675,N_29945);
nand UO_161 (O_161,N_29685,N_29056);
and UO_162 (O_162,N_28996,N_29957);
nand UO_163 (O_163,N_29093,N_29048);
nor UO_164 (O_164,N_29486,N_29407);
or UO_165 (O_165,N_29204,N_29848);
nand UO_166 (O_166,N_29043,N_29811);
nand UO_167 (O_167,N_29809,N_28974);
or UO_168 (O_168,N_29310,N_29717);
and UO_169 (O_169,N_28845,N_29235);
and UO_170 (O_170,N_29497,N_29283);
and UO_171 (O_171,N_29103,N_29599);
or UO_172 (O_172,N_29180,N_29886);
nor UO_173 (O_173,N_28832,N_29613);
and UO_174 (O_174,N_29245,N_28934);
or UO_175 (O_175,N_29035,N_29481);
or UO_176 (O_176,N_29883,N_29530);
nor UO_177 (O_177,N_29741,N_29747);
nand UO_178 (O_178,N_29959,N_29963);
and UO_179 (O_179,N_29082,N_29013);
nor UO_180 (O_180,N_29927,N_29162);
or UO_181 (O_181,N_29452,N_29560);
and UO_182 (O_182,N_29440,N_29751);
nor UO_183 (O_183,N_29840,N_29384);
or UO_184 (O_184,N_29138,N_29091);
nand UO_185 (O_185,N_29798,N_29595);
nor UO_186 (O_186,N_29564,N_29524);
nor UO_187 (O_187,N_29902,N_29807);
nor UO_188 (O_188,N_29281,N_29096);
xnor UO_189 (O_189,N_29996,N_29382);
nor UO_190 (O_190,N_29256,N_28969);
nor UO_191 (O_191,N_29923,N_29132);
nand UO_192 (O_192,N_28907,N_29801);
xnor UO_193 (O_193,N_29063,N_29055);
or UO_194 (O_194,N_29069,N_29783);
and UO_195 (O_195,N_29912,N_28955);
xor UO_196 (O_196,N_28800,N_29446);
nor UO_197 (O_197,N_29506,N_29111);
or UO_198 (O_198,N_29196,N_29614);
nand UO_199 (O_199,N_29379,N_29500);
and UO_200 (O_200,N_29877,N_29777);
nand UO_201 (O_201,N_29802,N_29395);
and UO_202 (O_202,N_29089,N_29846);
or UO_203 (O_203,N_29461,N_29167);
xor UO_204 (O_204,N_29436,N_29479);
nand UO_205 (O_205,N_29413,N_29094);
xor UO_206 (O_206,N_29805,N_28855);
or UO_207 (O_207,N_28930,N_29744);
and UO_208 (O_208,N_28859,N_28929);
xnor UO_209 (O_209,N_29556,N_29133);
or UO_210 (O_210,N_28987,N_29552);
and UO_211 (O_211,N_29620,N_29779);
or UO_212 (O_212,N_29067,N_29532);
and UO_213 (O_213,N_29514,N_28831);
xor UO_214 (O_214,N_29465,N_29414);
nor UO_215 (O_215,N_28823,N_29143);
nand UO_216 (O_216,N_29266,N_29836);
or UO_217 (O_217,N_29219,N_29693);
and UO_218 (O_218,N_29389,N_29203);
nand UO_219 (O_219,N_29255,N_29031);
nand UO_220 (O_220,N_28885,N_29667);
nor UO_221 (O_221,N_29125,N_29157);
nor UO_222 (O_222,N_29191,N_29823);
nor UO_223 (O_223,N_29107,N_29844);
nor UO_224 (O_224,N_29058,N_29126);
xor UO_225 (O_225,N_29208,N_29254);
xnor UO_226 (O_226,N_29367,N_28856);
or UO_227 (O_227,N_29121,N_28889);
nand UO_228 (O_228,N_29012,N_29027);
nand UO_229 (O_229,N_29602,N_29612);
nor UO_230 (O_230,N_29174,N_29504);
or UO_231 (O_231,N_28847,N_29890);
nor UO_232 (O_232,N_29349,N_29701);
nor UO_233 (O_233,N_29874,N_28986);
nor UO_234 (O_234,N_29993,N_29478);
nand UO_235 (O_235,N_29321,N_29363);
or UO_236 (O_236,N_29273,N_29764);
xnor UO_237 (O_237,N_28851,N_29885);
nor UO_238 (O_238,N_29079,N_29198);
nor UO_239 (O_239,N_29939,N_29210);
xor UO_240 (O_240,N_28879,N_29074);
xnor UO_241 (O_241,N_29397,N_29563);
nand UO_242 (O_242,N_29626,N_28935);
and UO_243 (O_243,N_29753,N_29019);
xnor UO_244 (O_244,N_29011,N_29527);
and UO_245 (O_245,N_29352,N_29616);
xnor UO_246 (O_246,N_29238,N_29916);
nor UO_247 (O_247,N_29110,N_29267);
and UO_248 (O_248,N_29732,N_29243);
nand UO_249 (O_249,N_29324,N_28868);
or UO_250 (O_250,N_29867,N_28813);
nor UO_251 (O_251,N_28814,N_29322);
nor UO_252 (O_252,N_29388,N_28972);
xor UO_253 (O_253,N_29991,N_29698);
xnor UO_254 (O_254,N_29474,N_29948);
nor UO_255 (O_255,N_29894,N_28891);
nor UO_256 (O_256,N_29009,N_29336);
or UO_257 (O_257,N_29134,N_29842);
and UO_258 (O_258,N_29825,N_29374);
or UO_259 (O_259,N_29466,N_29804);
nand UO_260 (O_260,N_28921,N_29720);
or UO_261 (O_261,N_29394,N_29308);
nor UO_262 (O_262,N_29543,N_29936);
xnor UO_263 (O_263,N_28933,N_29185);
xor UO_264 (O_264,N_29137,N_28901);
xnor UO_265 (O_265,N_28887,N_28951);
or UO_266 (O_266,N_29966,N_29489);
nand UO_267 (O_267,N_29512,N_29450);
xor UO_268 (O_268,N_29224,N_29052);
xnor UO_269 (O_269,N_28998,N_29730);
nor UO_270 (O_270,N_29933,N_29926);
nand UO_271 (O_271,N_29985,N_29600);
or UO_272 (O_272,N_28888,N_29983);
or UO_273 (O_273,N_29684,N_29906);
nand UO_274 (O_274,N_29641,N_29977);
nor UO_275 (O_275,N_29551,N_29547);
xor UO_276 (O_276,N_29326,N_28843);
xnor UO_277 (O_277,N_28857,N_29222);
nor UO_278 (O_278,N_29226,N_29689);
or UO_279 (O_279,N_29875,N_29334);
nand UO_280 (O_280,N_29344,N_29299);
nand UO_281 (O_281,N_29978,N_29253);
and UO_282 (O_282,N_28961,N_29156);
xor UO_283 (O_283,N_29635,N_28999);
xor UO_284 (O_284,N_29323,N_29230);
nor UO_285 (O_285,N_29630,N_29451);
nor UO_286 (O_286,N_28911,N_29519);
or UO_287 (O_287,N_29725,N_29895);
and UO_288 (O_288,N_29270,N_28988);
nor UO_289 (O_289,N_29533,N_29617);
or UO_290 (O_290,N_29348,N_29558);
nand UO_291 (O_291,N_29577,N_29782);
or UO_292 (O_292,N_29449,N_28898);
or UO_293 (O_293,N_29430,N_29611);
nor UO_294 (O_294,N_29333,N_29119);
nand UO_295 (O_295,N_28914,N_29406);
or UO_296 (O_296,N_29723,N_29432);
or UO_297 (O_297,N_29188,N_29220);
or UO_298 (O_298,N_29438,N_29607);
and UO_299 (O_299,N_29025,N_29246);
nor UO_300 (O_300,N_29335,N_29492);
or UO_301 (O_301,N_29239,N_28920);
nor UO_302 (O_302,N_29383,N_29148);
xor UO_303 (O_303,N_29309,N_29901);
or UO_304 (O_304,N_29586,N_29331);
nor UO_305 (O_305,N_29534,N_29488);
and UO_306 (O_306,N_29068,N_29733);
xnor UO_307 (O_307,N_29472,N_29920);
xor UO_308 (O_308,N_29932,N_29905);
and UO_309 (O_309,N_29772,N_28942);
and UO_310 (O_310,N_28968,N_29528);
nand UO_311 (O_311,N_29944,N_29080);
nor UO_312 (O_312,N_29410,N_29062);
and UO_313 (O_313,N_29338,N_29295);
xnor UO_314 (O_314,N_29900,N_29161);
nor UO_315 (O_315,N_29688,N_29573);
and UO_316 (O_316,N_29817,N_29863);
nor UO_317 (O_317,N_29756,N_29639);
xor UO_318 (O_318,N_29584,N_29455);
and UO_319 (O_319,N_29205,N_28964);
or UO_320 (O_320,N_29540,N_28874);
and UO_321 (O_321,N_29029,N_29142);
nand UO_322 (O_322,N_29005,N_28928);
or UO_323 (O_323,N_29790,N_29509);
nand UO_324 (O_324,N_29195,N_29827);
nor UO_325 (O_325,N_29731,N_29475);
nand UO_326 (O_326,N_29539,N_29419);
nor UO_327 (O_327,N_29938,N_29412);
nand UO_328 (O_328,N_29829,N_29629);
nor UO_329 (O_329,N_28894,N_29168);
or UO_330 (O_330,N_28864,N_29598);
or UO_331 (O_331,N_29313,N_28912);
nor UO_332 (O_332,N_29114,N_29522);
nor UO_333 (O_333,N_29291,N_29327);
nand UO_334 (O_334,N_29187,N_29544);
xnor UO_335 (O_335,N_29903,N_29248);
or UO_336 (O_336,N_29049,N_29580);
or UO_337 (O_337,N_28848,N_29781);
nand UO_338 (O_338,N_29269,N_29236);
and UO_339 (O_339,N_28837,N_29748);
nand UO_340 (O_340,N_29499,N_29373);
nor UO_341 (O_341,N_28873,N_29565);
or UO_342 (O_342,N_29555,N_28803);
nand UO_343 (O_343,N_29922,N_29320);
nor UO_344 (O_344,N_29697,N_29855);
xnor UO_345 (O_345,N_29637,N_28815);
xor UO_346 (O_346,N_29773,N_29958);
or UO_347 (O_347,N_29718,N_29057);
nor UO_348 (O_348,N_29002,N_29972);
xor UO_349 (O_349,N_28954,N_28818);
and UO_350 (O_350,N_29487,N_29918);
xor UO_351 (O_351,N_29445,N_29036);
nor UO_352 (O_352,N_29658,N_29365);
xor UO_353 (O_353,N_29870,N_28896);
nor UO_354 (O_354,N_28833,N_29100);
nand UO_355 (O_355,N_29583,N_29340);
xnor UO_356 (O_356,N_29405,N_29482);
nor UO_357 (O_357,N_29812,N_29705);
nor UO_358 (O_358,N_29582,N_29319);
or UO_359 (O_359,N_29385,N_29970);
or UO_360 (O_360,N_29806,N_29135);
xnor UO_361 (O_361,N_29416,N_28976);
or UO_362 (O_362,N_29816,N_28904);
xor UO_363 (O_363,N_29136,N_29961);
nor UO_364 (O_364,N_29652,N_29007);
and UO_365 (O_365,N_28849,N_29749);
or UO_366 (O_366,N_29277,N_29017);
nor UO_367 (O_367,N_29891,N_29604);
xnor UO_368 (O_368,N_28826,N_29257);
nand UO_369 (O_369,N_29884,N_29154);
nor UO_370 (O_370,N_29087,N_28824);
and UO_371 (O_371,N_29686,N_29856);
xnor UO_372 (O_372,N_29951,N_29186);
and UO_373 (O_373,N_29391,N_29665);
nand UO_374 (O_374,N_29707,N_28971);
xnor UO_375 (O_375,N_29788,N_29357);
or UO_376 (O_376,N_29288,N_29627);
or UO_377 (O_377,N_28883,N_28980);
or UO_378 (O_378,N_28893,N_29131);
xor UO_379 (O_379,N_29182,N_29699);
or UO_380 (O_380,N_29868,N_29442);
nor UO_381 (O_381,N_29839,N_28863);
and UO_382 (O_382,N_29673,N_29214);
nand UO_383 (O_383,N_29164,N_29526);
and UO_384 (O_384,N_29738,N_29171);
xor UO_385 (O_385,N_29633,N_28830);
nor UO_386 (O_386,N_28956,N_29571);
and UO_387 (O_387,N_29975,N_29974);
nand UO_388 (O_388,N_28872,N_29930);
xnor UO_389 (O_389,N_29776,N_29651);
nand UO_390 (O_390,N_29477,N_28966);
and UO_391 (O_391,N_29919,N_29147);
or UO_392 (O_392,N_28829,N_29439);
nand UO_393 (O_393,N_29468,N_29071);
or UO_394 (O_394,N_29632,N_29517);
or UO_395 (O_395,N_28908,N_29740);
nand UO_396 (O_396,N_29207,N_29190);
and UO_397 (O_397,N_29361,N_29787);
and UO_398 (O_398,N_29264,N_29332);
nand UO_399 (O_399,N_29914,N_29343);
nor UO_400 (O_400,N_28828,N_28842);
and UO_401 (O_401,N_29393,N_29850);
nor UO_402 (O_402,N_29404,N_29420);
xnor UO_403 (O_403,N_29928,N_29251);
xor UO_404 (O_404,N_29106,N_29523);
xor UO_405 (O_405,N_29692,N_28902);
xor UO_406 (O_406,N_29010,N_29800);
or UO_407 (O_407,N_29304,N_28866);
nand UO_408 (O_408,N_28938,N_29896);
and UO_409 (O_409,N_29622,N_29682);
nand UO_410 (O_410,N_29576,N_28984);
or UO_411 (O_411,N_29359,N_29588);
or UO_412 (O_412,N_29215,N_29078);
nor UO_413 (O_413,N_29178,N_29409);
and UO_414 (O_414,N_29562,N_29279);
xor UO_415 (O_415,N_29644,N_29988);
and UO_416 (O_416,N_28839,N_29399);
nor UO_417 (O_417,N_29780,N_29666);
and UO_418 (O_418,N_28805,N_29060);
nor UO_419 (O_419,N_29200,N_29739);
and UO_420 (O_420,N_29621,N_29108);
and UO_421 (O_421,N_29567,N_29833);
nand UO_422 (O_422,N_29480,N_29244);
nor UO_423 (O_423,N_28913,N_29550);
nor UO_424 (O_424,N_29808,N_29888);
xnor UO_425 (O_425,N_28975,N_29992);
and UO_426 (O_426,N_29199,N_28981);
and UO_427 (O_427,N_29004,N_29370);
nor UO_428 (O_428,N_29899,N_29341);
or UO_429 (O_429,N_29483,N_29376);
nand UO_430 (O_430,N_29030,N_29016);
or UO_431 (O_431,N_29940,N_29554);
or UO_432 (O_432,N_29854,N_28820);
and UO_433 (O_433,N_29173,N_29694);
nor UO_434 (O_434,N_28882,N_29640);
and UO_435 (O_435,N_29587,N_29176);
and UO_436 (O_436,N_28953,N_28917);
or UO_437 (O_437,N_28870,N_28982);
xnor UO_438 (O_438,N_28977,N_29218);
xor UO_439 (O_439,N_29380,N_29285);
nand UO_440 (O_440,N_29424,N_29231);
nand UO_441 (O_441,N_29347,N_29881);
and UO_442 (O_442,N_29858,N_28916);
or UO_443 (O_443,N_29202,N_29946);
and UO_444 (O_444,N_29028,N_29791);
xor UO_445 (O_445,N_29690,N_28979);
or UO_446 (O_446,N_29866,N_29981);
xor UO_447 (O_447,N_29819,N_29654);
nor UO_448 (O_448,N_29498,N_29460);
xnor UO_449 (O_449,N_29821,N_29893);
xor UO_450 (O_450,N_29838,N_29619);
xnor UO_451 (O_451,N_29559,N_29234);
xnor UO_452 (O_452,N_29953,N_28844);
xnor UO_453 (O_453,N_28821,N_29342);
or UO_454 (O_454,N_29358,N_29967);
and UO_455 (O_455,N_29908,N_29911);
xor UO_456 (O_456,N_29636,N_29982);
and UO_457 (O_457,N_28973,N_29700);
or UO_458 (O_458,N_28943,N_29386);
nor UO_459 (O_459,N_29081,N_29909);
nand UO_460 (O_460,N_29280,N_28895);
nand UO_461 (O_461,N_29775,N_29039);
and UO_462 (O_462,N_29390,N_28822);
nand UO_463 (O_463,N_29201,N_29109);
or UO_464 (O_464,N_28836,N_29754);
nor UO_465 (O_465,N_28950,N_29262);
xor UO_466 (O_466,N_29124,N_28993);
nor UO_467 (O_467,N_29857,N_29041);
xor UO_468 (O_468,N_29346,N_29871);
nor UO_469 (O_469,N_29965,N_29184);
or UO_470 (O_470,N_29678,N_29609);
or UO_471 (O_471,N_28860,N_29145);
nand UO_472 (O_472,N_29228,N_29098);
nand UO_473 (O_473,N_28923,N_29354);
nand UO_474 (O_474,N_29597,N_29294);
or UO_475 (O_475,N_29317,N_29954);
nand UO_476 (O_476,N_29258,N_29024);
xnor UO_477 (O_477,N_28990,N_29976);
nand UO_478 (O_478,N_29401,N_29669);
xor UO_479 (O_479,N_29618,N_29117);
xor UO_480 (O_480,N_28876,N_29995);
nand UO_481 (O_481,N_29149,N_29454);
nor UO_482 (O_482,N_29170,N_28854);
nand UO_483 (O_483,N_29815,N_29115);
nand UO_484 (O_484,N_28915,N_29507);
xnor UO_485 (O_485,N_29233,N_29292);
nor UO_486 (O_486,N_29463,N_29879);
nor UO_487 (O_487,N_29402,N_29443);
and UO_488 (O_488,N_29315,N_28890);
xnor UO_489 (O_489,N_29476,N_29691);
nor UO_490 (O_490,N_29375,N_29579);
nand UO_491 (O_491,N_29677,N_29670);
or UO_492 (O_492,N_29194,N_29033);
or UO_493 (O_493,N_28840,N_29159);
or UO_494 (O_494,N_29822,N_29102);
nand UO_495 (O_495,N_29913,N_28949);
nor UO_496 (O_496,N_29880,N_29721);
xnor UO_497 (O_497,N_29659,N_29925);
nor UO_498 (O_498,N_29064,N_29650);
xnor UO_499 (O_499,N_29427,N_28994);
or UO_500 (O_500,N_29032,N_29796);
or UO_501 (O_501,N_28846,N_29545);
xor UO_502 (O_502,N_29511,N_29706);
or UO_503 (O_503,N_28827,N_29860);
xor UO_504 (O_504,N_29793,N_29828);
or UO_505 (O_505,N_29727,N_28809);
or UO_506 (O_506,N_29054,N_29752);
nor UO_507 (O_507,N_29610,N_29964);
nor UO_508 (O_508,N_29059,N_29789);
xor UO_509 (O_509,N_29676,N_29268);
and UO_510 (O_510,N_29316,N_28957);
xor UO_511 (O_511,N_28877,N_29505);
or UO_512 (O_512,N_29183,N_29216);
nor UO_513 (O_513,N_29931,N_28983);
xor UO_514 (O_514,N_29301,N_29745);
nor UO_515 (O_515,N_29529,N_29950);
xor UO_516 (O_516,N_29987,N_29962);
nor UO_517 (O_517,N_28811,N_29647);
or UO_518 (O_518,N_29990,N_29755);
or UO_519 (O_519,N_28947,N_29924);
or UO_520 (O_520,N_29585,N_29728);
or UO_521 (O_521,N_29411,N_29634);
and UO_522 (O_522,N_29026,N_29937);
xor UO_523 (O_523,N_29638,N_29223);
or UO_524 (O_524,N_29240,N_29784);
and UO_525 (O_525,N_29249,N_28903);
nor UO_526 (O_526,N_29710,N_29623);
xnor UO_527 (O_527,N_28892,N_29518);
or UO_528 (O_528,N_29663,N_29968);
nor UO_529 (O_529,N_28941,N_29339);
or UO_530 (O_530,N_29876,N_29274);
and UO_531 (O_531,N_29935,N_29225);
nand UO_532 (O_532,N_29873,N_28834);
xor UO_533 (O_533,N_29181,N_29601);
nand UO_534 (O_534,N_29671,N_28841);
and UO_535 (O_535,N_29160,N_29960);
nand UO_536 (O_536,N_29774,N_29434);
or UO_537 (O_537,N_29546,N_29193);
or UO_538 (O_538,N_29371,N_29146);
and UO_539 (O_539,N_29872,N_29729);
or UO_540 (O_540,N_29934,N_29735);
and UO_541 (O_541,N_29606,N_29130);
xor UO_542 (O_542,N_28924,N_29155);
or UO_543 (O_543,N_28922,N_29708);
nand UO_544 (O_544,N_29541,N_28804);
or UO_545 (O_545,N_29660,N_29123);
and UO_546 (O_546,N_28825,N_29150);
or UO_547 (O_547,N_29456,N_29368);
nor UO_548 (O_548,N_29408,N_29525);
nor UO_549 (O_549,N_29832,N_29743);
and UO_550 (O_550,N_29300,N_28900);
or UO_551 (O_551,N_29305,N_28927);
or UO_552 (O_552,N_29849,N_29242);
nor UO_553 (O_553,N_29337,N_28932);
and UO_554 (O_554,N_28937,N_29172);
nand UO_555 (O_555,N_29447,N_28967);
nand UO_556 (O_556,N_29826,N_29984);
and UO_557 (O_557,N_28835,N_29703);
nand UO_558 (O_558,N_29290,N_29088);
nor UO_559 (O_559,N_29994,N_29097);
nand UO_560 (O_560,N_29046,N_29433);
nand UO_561 (O_561,N_28810,N_29387);
nor UO_562 (O_562,N_29355,N_29672);
xnor UO_563 (O_563,N_29820,N_29711);
nor UO_564 (O_564,N_29284,N_29726);
xor UO_565 (O_565,N_29073,N_29381);
and UO_566 (O_566,N_29008,N_29364);
or UO_567 (O_567,N_29531,N_29426);
and UO_568 (O_568,N_29818,N_29645);
nand UO_569 (O_569,N_29213,N_29714);
nand UO_570 (O_570,N_29569,N_28952);
or UO_571 (O_571,N_29166,N_28807);
or UO_572 (O_572,N_29158,N_29591);
xor UO_573 (O_573,N_29837,N_29018);
xnor UO_574 (O_574,N_29084,N_29835);
xor UO_575 (O_575,N_29537,N_29128);
or UO_576 (O_576,N_29099,N_29271);
or UO_577 (O_577,N_29038,N_29668);
xnor UO_578 (O_578,N_29485,N_29314);
xnor UO_579 (O_579,N_29192,N_29232);
xnor UO_580 (O_580,N_29603,N_29418);
xor UO_581 (O_581,N_29892,N_28853);
nor UO_582 (O_582,N_28989,N_29999);
xnor UO_583 (O_583,N_29329,N_28909);
nand UO_584 (O_584,N_29971,N_29656);
or UO_585 (O_585,N_29862,N_29719);
nand UO_586 (O_586,N_29261,N_29153);
xnor UO_587 (O_587,N_29763,N_29471);
xnor UO_588 (O_588,N_29679,N_29852);
or UO_589 (O_589,N_29561,N_29293);
nand UO_590 (O_590,N_29095,N_29047);
nand UO_591 (O_591,N_29553,N_29785);
or UO_592 (O_592,N_29557,N_29484);
and UO_593 (O_593,N_29615,N_29664);
and UO_594 (O_594,N_28852,N_29020);
nor UO_595 (O_595,N_29724,N_29152);
and UO_596 (O_596,N_29696,N_29713);
nor UO_597 (O_597,N_29469,N_29209);
xor UO_598 (O_598,N_28867,N_29538);
nor UO_599 (O_599,N_29141,N_29795);
nand UO_600 (O_600,N_28992,N_29089);
nand UO_601 (O_601,N_29138,N_29441);
nand UO_602 (O_602,N_29604,N_28803);
nand UO_603 (O_603,N_28873,N_28850);
and UO_604 (O_604,N_29844,N_29362);
nand UO_605 (O_605,N_29827,N_29075);
nor UO_606 (O_606,N_29838,N_29280);
and UO_607 (O_607,N_29556,N_29553);
nor UO_608 (O_608,N_29478,N_29618);
xnor UO_609 (O_609,N_28870,N_29858);
and UO_610 (O_610,N_29493,N_28999);
nand UO_611 (O_611,N_29946,N_29560);
nor UO_612 (O_612,N_29091,N_29377);
or UO_613 (O_613,N_29652,N_29321);
and UO_614 (O_614,N_29377,N_29371);
nor UO_615 (O_615,N_29679,N_29150);
or UO_616 (O_616,N_29185,N_28981);
nand UO_617 (O_617,N_29370,N_29892);
or UO_618 (O_618,N_29585,N_29378);
nand UO_619 (O_619,N_29074,N_29313);
nand UO_620 (O_620,N_29395,N_28979);
and UO_621 (O_621,N_28909,N_29312);
or UO_622 (O_622,N_29669,N_29935);
or UO_623 (O_623,N_28989,N_29390);
xnor UO_624 (O_624,N_29375,N_29224);
nand UO_625 (O_625,N_29609,N_29594);
xnor UO_626 (O_626,N_29960,N_29681);
and UO_627 (O_627,N_29084,N_29320);
xnor UO_628 (O_628,N_29950,N_28951);
nor UO_629 (O_629,N_29944,N_29126);
xor UO_630 (O_630,N_28819,N_29078);
xor UO_631 (O_631,N_29479,N_29884);
or UO_632 (O_632,N_28910,N_29788);
nand UO_633 (O_633,N_29948,N_29490);
xor UO_634 (O_634,N_29406,N_29987);
and UO_635 (O_635,N_29905,N_29168);
or UO_636 (O_636,N_29662,N_28986);
and UO_637 (O_637,N_29657,N_29489);
nand UO_638 (O_638,N_29608,N_29448);
nor UO_639 (O_639,N_29293,N_29709);
nor UO_640 (O_640,N_28816,N_28960);
and UO_641 (O_641,N_29615,N_29972);
nor UO_642 (O_642,N_29498,N_29477);
nor UO_643 (O_643,N_29215,N_28826);
or UO_644 (O_644,N_29644,N_28820);
xnor UO_645 (O_645,N_29236,N_29489);
and UO_646 (O_646,N_29516,N_29726);
and UO_647 (O_647,N_29772,N_29297);
nand UO_648 (O_648,N_29895,N_29425);
nand UO_649 (O_649,N_29164,N_29341);
and UO_650 (O_650,N_29379,N_29342);
nor UO_651 (O_651,N_29794,N_28868);
or UO_652 (O_652,N_29827,N_29500);
xor UO_653 (O_653,N_29575,N_29300);
nor UO_654 (O_654,N_29085,N_29983);
nand UO_655 (O_655,N_28923,N_29337);
nor UO_656 (O_656,N_29194,N_29929);
xor UO_657 (O_657,N_29405,N_29798);
nor UO_658 (O_658,N_29416,N_29689);
or UO_659 (O_659,N_29782,N_29272);
or UO_660 (O_660,N_28908,N_29747);
xnor UO_661 (O_661,N_29754,N_29775);
xnor UO_662 (O_662,N_29081,N_28978);
or UO_663 (O_663,N_29892,N_29886);
nand UO_664 (O_664,N_29307,N_29502);
and UO_665 (O_665,N_28845,N_29607);
or UO_666 (O_666,N_29223,N_29372);
xor UO_667 (O_667,N_29928,N_29043);
or UO_668 (O_668,N_29930,N_29337);
nor UO_669 (O_669,N_29865,N_29901);
or UO_670 (O_670,N_29296,N_29897);
xnor UO_671 (O_671,N_29643,N_29732);
nor UO_672 (O_672,N_29408,N_29445);
nand UO_673 (O_673,N_29048,N_29461);
xor UO_674 (O_674,N_29376,N_29980);
and UO_675 (O_675,N_29409,N_29505);
or UO_676 (O_676,N_28842,N_29551);
or UO_677 (O_677,N_29651,N_29232);
and UO_678 (O_678,N_29150,N_28920);
and UO_679 (O_679,N_29087,N_29036);
or UO_680 (O_680,N_29871,N_29573);
or UO_681 (O_681,N_29787,N_29323);
xnor UO_682 (O_682,N_29846,N_29674);
nand UO_683 (O_683,N_29007,N_29982);
or UO_684 (O_684,N_29864,N_29645);
nand UO_685 (O_685,N_29348,N_29443);
or UO_686 (O_686,N_29058,N_28829);
or UO_687 (O_687,N_29107,N_29720);
and UO_688 (O_688,N_29062,N_29139);
and UO_689 (O_689,N_29154,N_29184);
and UO_690 (O_690,N_29655,N_28809);
nor UO_691 (O_691,N_29132,N_29710);
nor UO_692 (O_692,N_28951,N_29133);
nor UO_693 (O_693,N_29493,N_29771);
xor UO_694 (O_694,N_29483,N_29994);
and UO_695 (O_695,N_29916,N_29800);
xor UO_696 (O_696,N_29668,N_29366);
nor UO_697 (O_697,N_29292,N_28923);
or UO_698 (O_698,N_29317,N_28917);
xor UO_699 (O_699,N_28805,N_29193);
or UO_700 (O_700,N_29614,N_29590);
nor UO_701 (O_701,N_29103,N_29682);
xnor UO_702 (O_702,N_29717,N_29925);
and UO_703 (O_703,N_29695,N_29009);
and UO_704 (O_704,N_29415,N_29551);
nor UO_705 (O_705,N_28921,N_29002);
or UO_706 (O_706,N_29435,N_29050);
xnor UO_707 (O_707,N_29783,N_28819);
nand UO_708 (O_708,N_28911,N_29466);
nand UO_709 (O_709,N_28959,N_29225);
xor UO_710 (O_710,N_29479,N_29405);
and UO_711 (O_711,N_29009,N_28930);
nand UO_712 (O_712,N_29261,N_29502);
and UO_713 (O_713,N_28855,N_28936);
nor UO_714 (O_714,N_29833,N_29236);
xnor UO_715 (O_715,N_29235,N_29158);
and UO_716 (O_716,N_29910,N_28859);
or UO_717 (O_717,N_29245,N_29601);
and UO_718 (O_718,N_28847,N_29390);
nor UO_719 (O_719,N_29098,N_29071);
nor UO_720 (O_720,N_29178,N_29774);
or UO_721 (O_721,N_29312,N_28827);
or UO_722 (O_722,N_28870,N_29476);
or UO_723 (O_723,N_29670,N_28920);
and UO_724 (O_724,N_29354,N_29874);
xnor UO_725 (O_725,N_29368,N_29489);
nand UO_726 (O_726,N_29992,N_29180);
or UO_727 (O_727,N_29406,N_28811);
or UO_728 (O_728,N_29040,N_29722);
nor UO_729 (O_729,N_29566,N_28988);
nor UO_730 (O_730,N_29706,N_29064);
xor UO_731 (O_731,N_28921,N_29906);
or UO_732 (O_732,N_28838,N_29992);
xor UO_733 (O_733,N_29849,N_29431);
nand UO_734 (O_734,N_29288,N_29387);
xor UO_735 (O_735,N_28936,N_29811);
and UO_736 (O_736,N_29753,N_29484);
and UO_737 (O_737,N_28893,N_29123);
nand UO_738 (O_738,N_29973,N_28823);
xor UO_739 (O_739,N_29292,N_28939);
nand UO_740 (O_740,N_29098,N_29474);
xnor UO_741 (O_741,N_29155,N_29165);
nand UO_742 (O_742,N_29755,N_29873);
xor UO_743 (O_743,N_29308,N_29438);
nor UO_744 (O_744,N_29636,N_29101);
or UO_745 (O_745,N_29818,N_29221);
nor UO_746 (O_746,N_29622,N_29178);
and UO_747 (O_747,N_28916,N_29968);
and UO_748 (O_748,N_29489,N_29569);
nor UO_749 (O_749,N_29300,N_29001);
nand UO_750 (O_750,N_29268,N_29829);
or UO_751 (O_751,N_29638,N_29038);
nand UO_752 (O_752,N_29360,N_29225);
nand UO_753 (O_753,N_29338,N_29071);
nor UO_754 (O_754,N_28896,N_29046);
nor UO_755 (O_755,N_28965,N_29069);
nor UO_756 (O_756,N_29013,N_29651);
nor UO_757 (O_757,N_29782,N_29527);
nand UO_758 (O_758,N_29473,N_29667);
xnor UO_759 (O_759,N_28930,N_29960);
nor UO_760 (O_760,N_29752,N_29251);
nand UO_761 (O_761,N_29162,N_29536);
nor UO_762 (O_762,N_29165,N_28822);
nor UO_763 (O_763,N_29913,N_29080);
xor UO_764 (O_764,N_28834,N_29552);
and UO_765 (O_765,N_29014,N_28822);
or UO_766 (O_766,N_29779,N_29396);
and UO_767 (O_767,N_29893,N_29105);
xnor UO_768 (O_768,N_29334,N_28885);
nor UO_769 (O_769,N_28889,N_28878);
xor UO_770 (O_770,N_28827,N_28884);
nor UO_771 (O_771,N_29964,N_29202);
and UO_772 (O_772,N_29572,N_29580);
nor UO_773 (O_773,N_29710,N_29448);
nand UO_774 (O_774,N_29691,N_28888);
nor UO_775 (O_775,N_28918,N_29096);
xor UO_776 (O_776,N_28993,N_29987);
and UO_777 (O_777,N_29289,N_29926);
and UO_778 (O_778,N_29757,N_29529);
xor UO_779 (O_779,N_29007,N_29431);
nand UO_780 (O_780,N_29269,N_29526);
nand UO_781 (O_781,N_29852,N_29496);
xnor UO_782 (O_782,N_28983,N_29976);
nand UO_783 (O_783,N_29855,N_29167);
or UO_784 (O_784,N_29682,N_29395);
and UO_785 (O_785,N_29665,N_28912);
nand UO_786 (O_786,N_29990,N_29646);
or UO_787 (O_787,N_28910,N_28887);
or UO_788 (O_788,N_29934,N_29188);
and UO_789 (O_789,N_28884,N_29462);
xnor UO_790 (O_790,N_29576,N_29681);
xnor UO_791 (O_791,N_29006,N_29882);
nand UO_792 (O_792,N_29239,N_29984);
xnor UO_793 (O_793,N_29880,N_29598);
xor UO_794 (O_794,N_29277,N_29118);
and UO_795 (O_795,N_28936,N_29034);
xnor UO_796 (O_796,N_29696,N_28974);
or UO_797 (O_797,N_29645,N_29450);
xor UO_798 (O_798,N_29721,N_29262);
nor UO_799 (O_799,N_28961,N_29010);
or UO_800 (O_800,N_29143,N_29904);
or UO_801 (O_801,N_29739,N_29023);
or UO_802 (O_802,N_29429,N_29241);
xnor UO_803 (O_803,N_29706,N_29898);
and UO_804 (O_804,N_29167,N_29192);
and UO_805 (O_805,N_29637,N_29926);
nand UO_806 (O_806,N_28804,N_29120);
and UO_807 (O_807,N_29580,N_28938);
nor UO_808 (O_808,N_29373,N_29230);
xnor UO_809 (O_809,N_28945,N_28822);
nand UO_810 (O_810,N_29916,N_29897);
xnor UO_811 (O_811,N_29740,N_28868);
nor UO_812 (O_812,N_29292,N_29737);
xor UO_813 (O_813,N_28882,N_29073);
nand UO_814 (O_814,N_29055,N_29413);
nand UO_815 (O_815,N_29734,N_29711);
nor UO_816 (O_816,N_29741,N_29834);
xnor UO_817 (O_817,N_28920,N_29682);
xor UO_818 (O_818,N_29030,N_29047);
nand UO_819 (O_819,N_28950,N_29893);
nand UO_820 (O_820,N_29291,N_29463);
xor UO_821 (O_821,N_29767,N_29729);
xnor UO_822 (O_822,N_29061,N_29742);
or UO_823 (O_823,N_29124,N_29236);
or UO_824 (O_824,N_29625,N_29757);
nand UO_825 (O_825,N_29772,N_29633);
nor UO_826 (O_826,N_29080,N_28890);
and UO_827 (O_827,N_29637,N_29611);
nand UO_828 (O_828,N_29191,N_29420);
or UO_829 (O_829,N_29340,N_28912);
nand UO_830 (O_830,N_29729,N_28945);
xor UO_831 (O_831,N_29945,N_29669);
and UO_832 (O_832,N_29514,N_28837);
nand UO_833 (O_833,N_29991,N_29796);
nand UO_834 (O_834,N_29414,N_29080);
nor UO_835 (O_835,N_29246,N_29863);
xor UO_836 (O_836,N_29179,N_29365);
nor UO_837 (O_837,N_29200,N_28815);
nor UO_838 (O_838,N_28937,N_29246);
or UO_839 (O_839,N_29553,N_29061);
and UO_840 (O_840,N_29243,N_29576);
or UO_841 (O_841,N_29051,N_29159);
and UO_842 (O_842,N_28856,N_28826);
xnor UO_843 (O_843,N_29326,N_28927);
xnor UO_844 (O_844,N_29598,N_29562);
and UO_845 (O_845,N_29780,N_29797);
or UO_846 (O_846,N_28903,N_29835);
xnor UO_847 (O_847,N_29967,N_29040);
nand UO_848 (O_848,N_29947,N_29410);
nor UO_849 (O_849,N_29061,N_29620);
and UO_850 (O_850,N_28871,N_29995);
nor UO_851 (O_851,N_29454,N_28830);
nor UO_852 (O_852,N_29510,N_28894);
nor UO_853 (O_853,N_29236,N_29354);
nand UO_854 (O_854,N_29876,N_29764);
and UO_855 (O_855,N_29968,N_29038);
and UO_856 (O_856,N_29194,N_29908);
and UO_857 (O_857,N_29188,N_28959);
or UO_858 (O_858,N_29848,N_29274);
nor UO_859 (O_859,N_29441,N_29566);
and UO_860 (O_860,N_29188,N_29099);
nand UO_861 (O_861,N_28818,N_29632);
and UO_862 (O_862,N_29685,N_29256);
nand UO_863 (O_863,N_29762,N_28969);
xnor UO_864 (O_864,N_29336,N_29232);
or UO_865 (O_865,N_29339,N_29201);
and UO_866 (O_866,N_29674,N_29936);
nand UO_867 (O_867,N_29712,N_28875);
and UO_868 (O_868,N_28934,N_28885);
xnor UO_869 (O_869,N_29238,N_29540);
and UO_870 (O_870,N_29419,N_29256);
xnor UO_871 (O_871,N_29992,N_29602);
xor UO_872 (O_872,N_28983,N_29450);
xnor UO_873 (O_873,N_29810,N_29733);
nor UO_874 (O_874,N_29815,N_29032);
nor UO_875 (O_875,N_29221,N_29603);
or UO_876 (O_876,N_29942,N_29712);
xor UO_877 (O_877,N_29299,N_29701);
or UO_878 (O_878,N_29383,N_29276);
and UO_879 (O_879,N_28970,N_29928);
xnor UO_880 (O_880,N_28884,N_29121);
or UO_881 (O_881,N_29847,N_28987);
xor UO_882 (O_882,N_29793,N_29500);
nor UO_883 (O_883,N_29974,N_29490);
xnor UO_884 (O_884,N_29073,N_29454);
xor UO_885 (O_885,N_28936,N_29749);
xor UO_886 (O_886,N_29606,N_28815);
xnor UO_887 (O_887,N_29806,N_29223);
xnor UO_888 (O_888,N_29266,N_29746);
nand UO_889 (O_889,N_28957,N_28982);
or UO_890 (O_890,N_29379,N_29878);
nor UO_891 (O_891,N_29761,N_29552);
nand UO_892 (O_892,N_29556,N_29814);
nand UO_893 (O_893,N_29001,N_29334);
nand UO_894 (O_894,N_28908,N_29382);
nand UO_895 (O_895,N_28840,N_29261);
xor UO_896 (O_896,N_29044,N_29392);
nor UO_897 (O_897,N_29474,N_29207);
xnor UO_898 (O_898,N_28818,N_29680);
nand UO_899 (O_899,N_28919,N_29933);
nor UO_900 (O_900,N_28918,N_29928);
or UO_901 (O_901,N_29969,N_29178);
nand UO_902 (O_902,N_28989,N_29247);
and UO_903 (O_903,N_29309,N_29151);
nand UO_904 (O_904,N_29393,N_29814);
or UO_905 (O_905,N_29000,N_29248);
nand UO_906 (O_906,N_29390,N_28926);
or UO_907 (O_907,N_29593,N_29906);
nand UO_908 (O_908,N_29904,N_29174);
nor UO_909 (O_909,N_29670,N_29535);
nor UO_910 (O_910,N_29723,N_29213);
xor UO_911 (O_911,N_28857,N_29758);
xor UO_912 (O_912,N_29497,N_29086);
and UO_913 (O_913,N_29199,N_29219);
nor UO_914 (O_914,N_28975,N_28961);
or UO_915 (O_915,N_29714,N_29827);
or UO_916 (O_916,N_29491,N_29440);
nor UO_917 (O_917,N_28883,N_28986);
or UO_918 (O_918,N_28946,N_29797);
xnor UO_919 (O_919,N_28943,N_28869);
or UO_920 (O_920,N_29622,N_29641);
nor UO_921 (O_921,N_29316,N_29166);
nand UO_922 (O_922,N_29046,N_29275);
xor UO_923 (O_923,N_29884,N_28961);
and UO_924 (O_924,N_28811,N_29693);
nor UO_925 (O_925,N_28800,N_29271);
nand UO_926 (O_926,N_28960,N_29281);
nand UO_927 (O_927,N_29120,N_29194);
nor UO_928 (O_928,N_29726,N_29958);
nor UO_929 (O_929,N_29462,N_29562);
and UO_930 (O_930,N_28865,N_29545);
nor UO_931 (O_931,N_29745,N_29091);
and UO_932 (O_932,N_29743,N_29746);
or UO_933 (O_933,N_29026,N_29134);
nand UO_934 (O_934,N_29350,N_29933);
nand UO_935 (O_935,N_28843,N_29220);
and UO_936 (O_936,N_29822,N_29357);
and UO_937 (O_937,N_28956,N_28941);
xor UO_938 (O_938,N_29646,N_29149);
and UO_939 (O_939,N_29891,N_29717);
and UO_940 (O_940,N_29080,N_29619);
or UO_941 (O_941,N_29958,N_29823);
or UO_942 (O_942,N_29402,N_29876);
xnor UO_943 (O_943,N_29911,N_29537);
or UO_944 (O_944,N_28945,N_29274);
nand UO_945 (O_945,N_29783,N_28950);
nor UO_946 (O_946,N_29310,N_29388);
or UO_947 (O_947,N_29208,N_29997);
nor UO_948 (O_948,N_29082,N_29411);
and UO_949 (O_949,N_28955,N_29101);
xor UO_950 (O_950,N_28979,N_29021);
or UO_951 (O_951,N_29669,N_29962);
xor UO_952 (O_952,N_29797,N_28876);
and UO_953 (O_953,N_29973,N_29049);
xor UO_954 (O_954,N_28903,N_29487);
nor UO_955 (O_955,N_29544,N_29228);
nor UO_956 (O_956,N_29027,N_29125);
nor UO_957 (O_957,N_29375,N_28911);
or UO_958 (O_958,N_29806,N_29971);
nor UO_959 (O_959,N_29466,N_29832);
nor UO_960 (O_960,N_28913,N_29580);
xor UO_961 (O_961,N_29096,N_28999);
nor UO_962 (O_962,N_29248,N_28936);
and UO_963 (O_963,N_29966,N_29549);
nor UO_964 (O_964,N_28938,N_29819);
nor UO_965 (O_965,N_29963,N_29342);
and UO_966 (O_966,N_28871,N_29799);
nor UO_967 (O_967,N_29308,N_29269);
and UO_968 (O_968,N_29806,N_29642);
or UO_969 (O_969,N_28858,N_29493);
xnor UO_970 (O_970,N_29653,N_29670);
nor UO_971 (O_971,N_29686,N_29865);
nor UO_972 (O_972,N_29833,N_29619);
or UO_973 (O_973,N_29793,N_29944);
and UO_974 (O_974,N_29086,N_29401);
nand UO_975 (O_975,N_29377,N_29651);
xnor UO_976 (O_976,N_28895,N_29965);
xnor UO_977 (O_977,N_29667,N_29923);
or UO_978 (O_978,N_29613,N_29134);
nor UO_979 (O_979,N_29847,N_29239);
and UO_980 (O_980,N_29733,N_29955);
and UO_981 (O_981,N_29706,N_29704);
nand UO_982 (O_982,N_29044,N_28891);
or UO_983 (O_983,N_29494,N_28860);
nor UO_984 (O_984,N_28876,N_29909);
and UO_985 (O_985,N_29202,N_29149);
nand UO_986 (O_986,N_29457,N_28837);
nand UO_987 (O_987,N_29176,N_29475);
nand UO_988 (O_988,N_29246,N_29857);
xor UO_989 (O_989,N_29829,N_29473);
nor UO_990 (O_990,N_29285,N_28853);
nand UO_991 (O_991,N_28912,N_29198);
and UO_992 (O_992,N_29839,N_29411);
or UO_993 (O_993,N_29922,N_29547);
and UO_994 (O_994,N_29949,N_28957);
xnor UO_995 (O_995,N_29224,N_29323);
and UO_996 (O_996,N_29625,N_29318);
or UO_997 (O_997,N_29166,N_29504);
and UO_998 (O_998,N_29190,N_29446);
and UO_999 (O_999,N_29629,N_29905);
nor UO_1000 (O_1000,N_29390,N_29206);
or UO_1001 (O_1001,N_28947,N_29054);
or UO_1002 (O_1002,N_29169,N_29423);
nor UO_1003 (O_1003,N_29581,N_29953);
nand UO_1004 (O_1004,N_29481,N_29618);
and UO_1005 (O_1005,N_29345,N_29851);
or UO_1006 (O_1006,N_29880,N_29017);
xor UO_1007 (O_1007,N_29219,N_29145);
nand UO_1008 (O_1008,N_29043,N_29398);
nor UO_1009 (O_1009,N_28852,N_29605);
nand UO_1010 (O_1010,N_29731,N_29425);
or UO_1011 (O_1011,N_29618,N_29331);
and UO_1012 (O_1012,N_29244,N_29104);
or UO_1013 (O_1013,N_29533,N_29513);
nand UO_1014 (O_1014,N_29624,N_28989);
or UO_1015 (O_1015,N_28802,N_29216);
xor UO_1016 (O_1016,N_28892,N_29256);
nand UO_1017 (O_1017,N_29766,N_29626);
nor UO_1018 (O_1018,N_28970,N_29628);
or UO_1019 (O_1019,N_29387,N_29954);
and UO_1020 (O_1020,N_29880,N_29847);
or UO_1021 (O_1021,N_29177,N_29584);
xnor UO_1022 (O_1022,N_29738,N_28828);
xor UO_1023 (O_1023,N_29853,N_29482);
nor UO_1024 (O_1024,N_29533,N_29232);
nand UO_1025 (O_1025,N_29838,N_29785);
nor UO_1026 (O_1026,N_28897,N_29259);
nand UO_1027 (O_1027,N_29790,N_29854);
xnor UO_1028 (O_1028,N_28868,N_29221);
nand UO_1029 (O_1029,N_29148,N_29535);
xor UO_1030 (O_1030,N_29061,N_29250);
or UO_1031 (O_1031,N_29312,N_29154);
nor UO_1032 (O_1032,N_29308,N_29630);
nand UO_1033 (O_1033,N_28870,N_29263);
or UO_1034 (O_1034,N_29054,N_28940);
xor UO_1035 (O_1035,N_28892,N_28807);
xor UO_1036 (O_1036,N_29675,N_29236);
nand UO_1037 (O_1037,N_29558,N_29618);
xor UO_1038 (O_1038,N_29602,N_28926);
xnor UO_1039 (O_1039,N_29287,N_29925);
and UO_1040 (O_1040,N_29850,N_28903);
or UO_1041 (O_1041,N_29318,N_29376);
or UO_1042 (O_1042,N_29837,N_29221);
and UO_1043 (O_1043,N_29538,N_29947);
nor UO_1044 (O_1044,N_29395,N_29606);
or UO_1045 (O_1045,N_29583,N_28868);
nor UO_1046 (O_1046,N_29760,N_28864);
xnor UO_1047 (O_1047,N_29249,N_29182);
and UO_1048 (O_1048,N_29203,N_29079);
nor UO_1049 (O_1049,N_29500,N_29516);
and UO_1050 (O_1050,N_29691,N_29312);
xor UO_1051 (O_1051,N_29319,N_29693);
xor UO_1052 (O_1052,N_29433,N_29771);
nand UO_1053 (O_1053,N_29006,N_29243);
or UO_1054 (O_1054,N_29993,N_29920);
and UO_1055 (O_1055,N_29637,N_29796);
xnor UO_1056 (O_1056,N_29431,N_29334);
and UO_1057 (O_1057,N_29044,N_29245);
nor UO_1058 (O_1058,N_29678,N_29135);
nor UO_1059 (O_1059,N_29684,N_29548);
or UO_1060 (O_1060,N_29196,N_29222);
nor UO_1061 (O_1061,N_28960,N_29135);
or UO_1062 (O_1062,N_28855,N_29915);
nand UO_1063 (O_1063,N_29928,N_29963);
nand UO_1064 (O_1064,N_29992,N_29879);
xnor UO_1065 (O_1065,N_29787,N_29384);
nor UO_1066 (O_1066,N_28880,N_29606);
xor UO_1067 (O_1067,N_28954,N_29614);
nor UO_1068 (O_1068,N_29660,N_29633);
and UO_1069 (O_1069,N_29868,N_29663);
nand UO_1070 (O_1070,N_29520,N_29177);
and UO_1071 (O_1071,N_29266,N_29921);
and UO_1072 (O_1072,N_29816,N_28859);
or UO_1073 (O_1073,N_29651,N_28876);
or UO_1074 (O_1074,N_28875,N_28808);
or UO_1075 (O_1075,N_29735,N_29663);
nand UO_1076 (O_1076,N_29328,N_29699);
and UO_1077 (O_1077,N_29160,N_29557);
xnor UO_1078 (O_1078,N_29776,N_29505);
and UO_1079 (O_1079,N_29131,N_28968);
nor UO_1080 (O_1080,N_29575,N_29377);
nand UO_1081 (O_1081,N_29667,N_29005);
nor UO_1082 (O_1082,N_29789,N_29715);
and UO_1083 (O_1083,N_28890,N_29379);
xnor UO_1084 (O_1084,N_29120,N_29273);
nand UO_1085 (O_1085,N_29920,N_29625);
xnor UO_1086 (O_1086,N_29015,N_28884);
xor UO_1087 (O_1087,N_29893,N_29442);
xor UO_1088 (O_1088,N_29857,N_28867);
or UO_1089 (O_1089,N_29737,N_28991);
nor UO_1090 (O_1090,N_29520,N_29830);
nand UO_1091 (O_1091,N_29178,N_29498);
or UO_1092 (O_1092,N_28818,N_29384);
and UO_1093 (O_1093,N_29448,N_28967);
nor UO_1094 (O_1094,N_29399,N_29771);
and UO_1095 (O_1095,N_29868,N_29988);
and UO_1096 (O_1096,N_29940,N_29913);
or UO_1097 (O_1097,N_29806,N_29913);
xnor UO_1098 (O_1098,N_29472,N_29429);
xnor UO_1099 (O_1099,N_29357,N_28902);
or UO_1100 (O_1100,N_29775,N_29541);
nand UO_1101 (O_1101,N_29899,N_29835);
or UO_1102 (O_1102,N_29569,N_29598);
nand UO_1103 (O_1103,N_29659,N_28924);
nand UO_1104 (O_1104,N_29107,N_29858);
and UO_1105 (O_1105,N_29584,N_28973);
xnor UO_1106 (O_1106,N_29125,N_29418);
nor UO_1107 (O_1107,N_29456,N_29380);
and UO_1108 (O_1108,N_29509,N_29763);
and UO_1109 (O_1109,N_29269,N_29465);
nor UO_1110 (O_1110,N_29043,N_29507);
nor UO_1111 (O_1111,N_29252,N_29085);
nand UO_1112 (O_1112,N_29399,N_28847);
nand UO_1113 (O_1113,N_29361,N_29172);
xnor UO_1114 (O_1114,N_29829,N_28910);
nand UO_1115 (O_1115,N_29351,N_29910);
xnor UO_1116 (O_1116,N_29932,N_28844);
nor UO_1117 (O_1117,N_29377,N_29200);
and UO_1118 (O_1118,N_29321,N_29750);
and UO_1119 (O_1119,N_29922,N_29777);
or UO_1120 (O_1120,N_29685,N_28845);
nor UO_1121 (O_1121,N_29764,N_29252);
or UO_1122 (O_1122,N_29362,N_28966);
nor UO_1123 (O_1123,N_29625,N_29938);
nor UO_1124 (O_1124,N_28821,N_29689);
or UO_1125 (O_1125,N_29192,N_29004);
and UO_1126 (O_1126,N_28957,N_29600);
nand UO_1127 (O_1127,N_29328,N_29016);
or UO_1128 (O_1128,N_29030,N_29362);
or UO_1129 (O_1129,N_29136,N_29769);
nor UO_1130 (O_1130,N_29987,N_29741);
nand UO_1131 (O_1131,N_28883,N_29879);
nor UO_1132 (O_1132,N_29633,N_29774);
xor UO_1133 (O_1133,N_29479,N_29419);
nand UO_1134 (O_1134,N_29069,N_29792);
and UO_1135 (O_1135,N_29727,N_29457);
xor UO_1136 (O_1136,N_29401,N_29642);
nand UO_1137 (O_1137,N_28881,N_29339);
and UO_1138 (O_1138,N_29189,N_29687);
nand UO_1139 (O_1139,N_28981,N_29931);
or UO_1140 (O_1140,N_28932,N_29769);
or UO_1141 (O_1141,N_29663,N_29936);
nand UO_1142 (O_1142,N_29818,N_29569);
xor UO_1143 (O_1143,N_29169,N_29721);
and UO_1144 (O_1144,N_28839,N_29814);
or UO_1145 (O_1145,N_29667,N_29419);
xnor UO_1146 (O_1146,N_28827,N_29002);
xnor UO_1147 (O_1147,N_29674,N_29546);
and UO_1148 (O_1148,N_29788,N_28824);
nand UO_1149 (O_1149,N_28939,N_29625);
nor UO_1150 (O_1150,N_28823,N_29030);
and UO_1151 (O_1151,N_29802,N_29496);
or UO_1152 (O_1152,N_29707,N_29981);
xnor UO_1153 (O_1153,N_29230,N_29243);
xnor UO_1154 (O_1154,N_29732,N_29469);
and UO_1155 (O_1155,N_29302,N_29671);
or UO_1156 (O_1156,N_29774,N_29703);
xor UO_1157 (O_1157,N_29981,N_29790);
and UO_1158 (O_1158,N_28986,N_29059);
xor UO_1159 (O_1159,N_28836,N_29632);
nand UO_1160 (O_1160,N_29429,N_28861);
nor UO_1161 (O_1161,N_29692,N_28965);
xnor UO_1162 (O_1162,N_29219,N_29938);
nor UO_1163 (O_1163,N_28894,N_29495);
or UO_1164 (O_1164,N_28937,N_29757);
nand UO_1165 (O_1165,N_29539,N_29810);
or UO_1166 (O_1166,N_28915,N_29509);
xnor UO_1167 (O_1167,N_29229,N_29738);
nor UO_1168 (O_1168,N_29422,N_29810);
or UO_1169 (O_1169,N_29111,N_28909);
xor UO_1170 (O_1170,N_29744,N_29804);
and UO_1171 (O_1171,N_29688,N_29303);
xor UO_1172 (O_1172,N_29002,N_29317);
nand UO_1173 (O_1173,N_29963,N_29875);
nor UO_1174 (O_1174,N_29729,N_28917);
nand UO_1175 (O_1175,N_29515,N_29448);
xor UO_1176 (O_1176,N_29711,N_29664);
nor UO_1177 (O_1177,N_29234,N_28858);
nor UO_1178 (O_1178,N_29363,N_28882);
and UO_1179 (O_1179,N_29947,N_29921);
nor UO_1180 (O_1180,N_29158,N_29200);
xor UO_1181 (O_1181,N_29999,N_29095);
xor UO_1182 (O_1182,N_29168,N_29673);
and UO_1183 (O_1183,N_29325,N_29511);
nand UO_1184 (O_1184,N_29771,N_28838);
and UO_1185 (O_1185,N_29150,N_29143);
xor UO_1186 (O_1186,N_28938,N_29843);
and UO_1187 (O_1187,N_28818,N_29610);
and UO_1188 (O_1188,N_28904,N_28906);
nor UO_1189 (O_1189,N_28927,N_29114);
nor UO_1190 (O_1190,N_29059,N_28952);
and UO_1191 (O_1191,N_29108,N_29163);
nand UO_1192 (O_1192,N_29306,N_29749);
nor UO_1193 (O_1193,N_28998,N_29247);
nor UO_1194 (O_1194,N_29819,N_28919);
nor UO_1195 (O_1195,N_28949,N_29216);
xor UO_1196 (O_1196,N_29733,N_29041);
xnor UO_1197 (O_1197,N_29186,N_29773);
nand UO_1198 (O_1198,N_28858,N_29736);
nor UO_1199 (O_1199,N_29106,N_28932);
nand UO_1200 (O_1200,N_29938,N_29952);
nor UO_1201 (O_1201,N_29136,N_29106);
xor UO_1202 (O_1202,N_29971,N_29596);
xor UO_1203 (O_1203,N_29019,N_28986);
xor UO_1204 (O_1204,N_29519,N_28821);
and UO_1205 (O_1205,N_29045,N_29814);
xor UO_1206 (O_1206,N_29129,N_28956);
and UO_1207 (O_1207,N_28863,N_29760);
nor UO_1208 (O_1208,N_29570,N_29025);
nand UO_1209 (O_1209,N_29482,N_29119);
nor UO_1210 (O_1210,N_29344,N_28949);
nand UO_1211 (O_1211,N_28841,N_28966);
and UO_1212 (O_1212,N_29008,N_29371);
xnor UO_1213 (O_1213,N_29869,N_29686);
or UO_1214 (O_1214,N_29537,N_29329);
nor UO_1215 (O_1215,N_29918,N_29828);
and UO_1216 (O_1216,N_29779,N_29335);
xor UO_1217 (O_1217,N_29670,N_29255);
or UO_1218 (O_1218,N_28938,N_29343);
nand UO_1219 (O_1219,N_28916,N_29634);
nor UO_1220 (O_1220,N_29604,N_29709);
xnor UO_1221 (O_1221,N_29308,N_29937);
or UO_1222 (O_1222,N_28894,N_29121);
xor UO_1223 (O_1223,N_29031,N_28895);
nor UO_1224 (O_1224,N_29411,N_28941);
nand UO_1225 (O_1225,N_29660,N_29915);
nor UO_1226 (O_1226,N_29909,N_29249);
xor UO_1227 (O_1227,N_29209,N_29602);
nor UO_1228 (O_1228,N_29770,N_29981);
xnor UO_1229 (O_1229,N_29624,N_29165);
and UO_1230 (O_1230,N_29408,N_29058);
or UO_1231 (O_1231,N_29466,N_29534);
nand UO_1232 (O_1232,N_29598,N_29897);
nor UO_1233 (O_1233,N_29840,N_28939);
nand UO_1234 (O_1234,N_29094,N_29894);
or UO_1235 (O_1235,N_29895,N_28913);
nand UO_1236 (O_1236,N_29210,N_29078);
or UO_1237 (O_1237,N_29481,N_28831);
or UO_1238 (O_1238,N_29505,N_29422);
nor UO_1239 (O_1239,N_29973,N_29495);
xnor UO_1240 (O_1240,N_28929,N_29257);
or UO_1241 (O_1241,N_29931,N_29990);
nor UO_1242 (O_1242,N_29040,N_29036);
nor UO_1243 (O_1243,N_29182,N_29642);
and UO_1244 (O_1244,N_29493,N_29428);
xor UO_1245 (O_1245,N_29620,N_29208);
xor UO_1246 (O_1246,N_29400,N_29061);
or UO_1247 (O_1247,N_29635,N_29187);
xnor UO_1248 (O_1248,N_28924,N_29261);
nor UO_1249 (O_1249,N_28901,N_29772);
or UO_1250 (O_1250,N_29584,N_29593);
nand UO_1251 (O_1251,N_29861,N_29920);
xor UO_1252 (O_1252,N_29655,N_29396);
and UO_1253 (O_1253,N_29450,N_29878);
nor UO_1254 (O_1254,N_29908,N_29993);
xor UO_1255 (O_1255,N_29221,N_29044);
or UO_1256 (O_1256,N_29625,N_29709);
nor UO_1257 (O_1257,N_29827,N_29675);
nor UO_1258 (O_1258,N_29168,N_29011);
nor UO_1259 (O_1259,N_29550,N_29671);
or UO_1260 (O_1260,N_29565,N_28993);
nand UO_1261 (O_1261,N_29104,N_29591);
nand UO_1262 (O_1262,N_29889,N_29246);
xor UO_1263 (O_1263,N_29949,N_29176);
xnor UO_1264 (O_1264,N_29783,N_29681);
and UO_1265 (O_1265,N_29101,N_29753);
or UO_1266 (O_1266,N_28943,N_29135);
nand UO_1267 (O_1267,N_28939,N_29401);
nand UO_1268 (O_1268,N_29076,N_28888);
nor UO_1269 (O_1269,N_29194,N_29365);
or UO_1270 (O_1270,N_29173,N_29433);
or UO_1271 (O_1271,N_29396,N_29837);
nor UO_1272 (O_1272,N_29555,N_29054);
and UO_1273 (O_1273,N_29293,N_29934);
and UO_1274 (O_1274,N_29901,N_29230);
or UO_1275 (O_1275,N_29171,N_29790);
or UO_1276 (O_1276,N_29267,N_28950);
or UO_1277 (O_1277,N_29349,N_29326);
and UO_1278 (O_1278,N_29701,N_29950);
xor UO_1279 (O_1279,N_28884,N_29282);
and UO_1280 (O_1280,N_28913,N_29516);
and UO_1281 (O_1281,N_29887,N_29689);
xor UO_1282 (O_1282,N_29616,N_28942);
and UO_1283 (O_1283,N_29972,N_29212);
xnor UO_1284 (O_1284,N_29261,N_29313);
nand UO_1285 (O_1285,N_29109,N_29564);
and UO_1286 (O_1286,N_29526,N_29682);
nor UO_1287 (O_1287,N_29990,N_29462);
and UO_1288 (O_1288,N_29267,N_29352);
nand UO_1289 (O_1289,N_29815,N_28909);
or UO_1290 (O_1290,N_29121,N_28814);
nor UO_1291 (O_1291,N_29907,N_29762);
nor UO_1292 (O_1292,N_29615,N_29281);
nor UO_1293 (O_1293,N_28996,N_29417);
xor UO_1294 (O_1294,N_29469,N_29460);
or UO_1295 (O_1295,N_29524,N_29797);
xnor UO_1296 (O_1296,N_28959,N_29110);
xor UO_1297 (O_1297,N_29260,N_29931);
or UO_1298 (O_1298,N_29922,N_29362);
and UO_1299 (O_1299,N_28955,N_29124);
xnor UO_1300 (O_1300,N_29918,N_29568);
xnor UO_1301 (O_1301,N_29000,N_29909);
nand UO_1302 (O_1302,N_29223,N_29935);
or UO_1303 (O_1303,N_28815,N_29230);
and UO_1304 (O_1304,N_29614,N_29110);
or UO_1305 (O_1305,N_29285,N_29208);
xnor UO_1306 (O_1306,N_28852,N_29273);
or UO_1307 (O_1307,N_28976,N_29674);
xnor UO_1308 (O_1308,N_29570,N_29736);
and UO_1309 (O_1309,N_29858,N_29855);
and UO_1310 (O_1310,N_29258,N_28892);
or UO_1311 (O_1311,N_28935,N_28828);
nor UO_1312 (O_1312,N_29313,N_29984);
xnor UO_1313 (O_1313,N_29665,N_29170);
nand UO_1314 (O_1314,N_29238,N_29788);
or UO_1315 (O_1315,N_29192,N_29540);
or UO_1316 (O_1316,N_29950,N_29784);
and UO_1317 (O_1317,N_29131,N_29114);
xor UO_1318 (O_1318,N_29091,N_28939);
nor UO_1319 (O_1319,N_29214,N_29304);
xor UO_1320 (O_1320,N_29984,N_29596);
and UO_1321 (O_1321,N_29300,N_29574);
nand UO_1322 (O_1322,N_29913,N_28981);
nand UO_1323 (O_1323,N_29324,N_29184);
or UO_1324 (O_1324,N_29486,N_29573);
nand UO_1325 (O_1325,N_29721,N_29062);
nor UO_1326 (O_1326,N_29158,N_28853);
xnor UO_1327 (O_1327,N_29604,N_29717);
xor UO_1328 (O_1328,N_29722,N_29536);
and UO_1329 (O_1329,N_28898,N_29486);
xnor UO_1330 (O_1330,N_29495,N_29443);
xnor UO_1331 (O_1331,N_29320,N_29706);
nor UO_1332 (O_1332,N_29322,N_29537);
nand UO_1333 (O_1333,N_29387,N_29761);
nor UO_1334 (O_1334,N_29363,N_29762);
or UO_1335 (O_1335,N_29404,N_29499);
nor UO_1336 (O_1336,N_29516,N_28920);
and UO_1337 (O_1337,N_29077,N_29137);
nor UO_1338 (O_1338,N_28882,N_29903);
xor UO_1339 (O_1339,N_29756,N_29231);
or UO_1340 (O_1340,N_28834,N_29709);
xnor UO_1341 (O_1341,N_29237,N_29228);
xnor UO_1342 (O_1342,N_28961,N_29787);
xor UO_1343 (O_1343,N_28829,N_29662);
and UO_1344 (O_1344,N_29284,N_29278);
or UO_1345 (O_1345,N_29767,N_29972);
and UO_1346 (O_1346,N_29392,N_29572);
xnor UO_1347 (O_1347,N_29437,N_29007);
and UO_1348 (O_1348,N_29143,N_29744);
xnor UO_1349 (O_1349,N_29710,N_29102);
and UO_1350 (O_1350,N_29671,N_29133);
and UO_1351 (O_1351,N_29514,N_29763);
and UO_1352 (O_1352,N_29220,N_29962);
or UO_1353 (O_1353,N_28895,N_29564);
or UO_1354 (O_1354,N_29537,N_28943);
xor UO_1355 (O_1355,N_29989,N_29758);
or UO_1356 (O_1356,N_28909,N_28886);
xnor UO_1357 (O_1357,N_29655,N_29650);
xnor UO_1358 (O_1358,N_29372,N_29551);
nor UO_1359 (O_1359,N_29115,N_28815);
or UO_1360 (O_1360,N_29055,N_29253);
or UO_1361 (O_1361,N_29883,N_29692);
or UO_1362 (O_1362,N_29401,N_29648);
nor UO_1363 (O_1363,N_29205,N_29977);
and UO_1364 (O_1364,N_29697,N_29826);
and UO_1365 (O_1365,N_28883,N_29538);
and UO_1366 (O_1366,N_29937,N_29392);
xnor UO_1367 (O_1367,N_29771,N_28969);
or UO_1368 (O_1368,N_29611,N_29869);
and UO_1369 (O_1369,N_29972,N_29589);
or UO_1370 (O_1370,N_29877,N_29732);
or UO_1371 (O_1371,N_29626,N_29107);
xor UO_1372 (O_1372,N_29949,N_28842);
nand UO_1373 (O_1373,N_29230,N_29505);
xor UO_1374 (O_1374,N_29086,N_29534);
xor UO_1375 (O_1375,N_29009,N_29814);
or UO_1376 (O_1376,N_29867,N_29311);
or UO_1377 (O_1377,N_29479,N_29030);
nand UO_1378 (O_1378,N_29189,N_29794);
nand UO_1379 (O_1379,N_29314,N_28990);
xor UO_1380 (O_1380,N_29911,N_28878);
xor UO_1381 (O_1381,N_29926,N_28828);
xnor UO_1382 (O_1382,N_29476,N_28881);
or UO_1383 (O_1383,N_29425,N_29848);
nor UO_1384 (O_1384,N_29546,N_29633);
or UO_1385 (O_1385,N_29259,N_29650);
xor UO_1386 (O_1386,N_29469,N_29548);
nand UO_1387 (O_1387,N_29164,N_29802);
or UO_1388 (O_1388,N_29980,N_29359);
and UO_1389 (O_1389,N_29407,N_29791);
xor UO_1390 (O_1390,N_29542,N_29637);
or UO_1391 (O_1391,N_29025,N_29487);
nand UO_1392 (O_1392,N_29967,N_29061);
nor UO_1393 (O_1393,N_28849,N_29212);
xor UO_1394 (O_1394,N_29111,N_29361);
and UO_1395 (O_1395,N_28982,N_29214);
nand UO_1396 (O_1396,N_28902,N_28986);
nor UO_1397 (O_1397,N_29488,N_29644);
nand UO_1398 (O_1398,N_29694,N_28945);
nor UO_1399 (O_1399,N_29052,N_28853);
nor UO_1400 (O_1400,N_29607,N_29117);
nand UO_1401 (O_1401,N_29881,N_29031);
nor UO_1402 (O_1402,N_29270,N_29950);
and UO_1403 (O_1403,N_29623,N_29534);
nor UO_1404 (O_1404,N_29292,N_29704);
nand UO_1405 (O_1405,N_29335,N_28889);
xor UO_1406 (O_1406,N_29485,N_29289);
and UO_1407 (O_1407,N_28965,N_29374);
xnor UO_1408 (O_1408,N_28964,N_29829);
nor UO_1409 (O_1409,N_29395,N_29853);
xnor UO_1410 (O_1410,N_29317,N_29059);
or UO_1411 (O_1411,N_29715,N_29905);
nand UO_1412 (O_1412,N_29797,N_29995);
and UO_1413 (O_1413,N_29565,N_29254);
nand UO_1414 (O_1414,N_29211,N_29625);
or UO_1415 (O_1415,N_29046,N_29870);
or UO_1416 (O_1416,N_29582,N_29900);
xnor UO_1417 (O_1417,N_28813,N_29125);
xor UO_1418 (O_1418,N_29978,N_28839);
xor UO_1419 (O_1419,N_29999,N_29342);
nor UO_1420 (O_1420,N_29091,N_29239);
nor UO_1421 (O_1421,N_29318,N_28925);
nor UO_1422 (O_1422,N_29870,N_29350);
nand UO_1423 (O_1423,N_29974,N_29070);
or UO_1424 (O_1424,N_29230,N_28884);
or UO_1425 (O_1425,N_29777,N_28927);
nor UO_1426 (O_1426,N_29963,N_29089);
nor UO_1427 (O_1427,N_29284,N_29254);
and UO_1428 (O_1428,N_29896,N_29197);
or UO_1429 (O_1429,N_29848,N_29816);
nor UO_1430 (O_1430,N_28991,N_29669);
or UO_1431 (O_1431,N_29346,N_29983);
xnor UO_1432 (O_1432,N_29042,N_29152);
xnor UO_1433 (O_1433,N_28942,N_29429);
and UO_1434 (O_1434,N_29756,N_29374);
nand UO_1435 (O_1435,N_28820,N_28807);
nand UO_1436 (O_1436,N_29396,N_29148);
and UO_1437 (O_1437,N_29945,N_29722);
nor UO_1438 (O_1438,N_29058,N_29457);
or UO_1439 (O_1439,N_29297,N_29729);
xor UO_1440 (O_1440,N_29871,N_29183);
xor UO_1441 (O_1441,N_29874,N_29520);
xnor UO_1442 (O_1442,N_29973,N_28917);
and UO_1443 (O_1443,N_29790,N_29254);
or UO_1444 (O_1444,N_29481,N_29454);
or UO_1445 (O_1445,N_29551,N_29842);
and UO_1446 (O_1446,N_29855,N_29623);
and UO_1447 (O_1447,N_28810,N_29343);
nand UO_1448 (O_1448,N_29921,N_29141);
nand UO_1449 (O_1449,N_29599,N_29422);
nor UO_1450 (O_1450,N_29921,N_29012);
nand UO_1451 (O_1451,N_29563,N_29205);
nor UO_1452 (O_1452,N_29739,N_29430);
nor UO_1453 (O_1453,N_29809,N_29589);
or UO_1454 (O_1454,N_29108,N_29649);
nor UO_1455 (O_1455,N_29543,N_29082);
nand UO_1456 (O_1456,N_29804,N_28863);
or UO_1457 (O_1457,N_29379,N_29506);
and UO_1458 (O_1458,N_29890,N_29209);
xnor UO_1459 (O_1459,N_29626,N_28966);
xor UO_1460 (O_1460,N_29102,N_29481);
and UO_1461 (O_1461,N_29714,N_29402);
or UO_1462 (O_1462,N_29243,N_29305);
xnor UO_1463 (O_1463,N_29060,N_28901);
or UO_1464 (O_1464,N_29022,N_29797);
xor UO_1465 (O_1465,N_29008,N_29029);
xnor UO_1466 (O_1466,N_28910,N_29071);
nor UO_1467 (O_1467,N_28876,N_29529);
xnor UO_1468 (O_1468,N_29515,N_29059);
nor UO_1469 (O_1469,N_29436,N_28836);
nor UO_1470 (O_1470,N_29778,N_29163);
nor UO_1471 (O_1471,N_29624,N_29136);
xor UO_1472 (O_1472,N_28903,N_29656);
nor UO_1473 (O_1473,N_29961,N_29071);
nor UO_1474 (O_1474,N_29418,N_29492);
xor UO_1475 (O_1475,N_28824,N_29530);
or UO_1476 (O_1476,N_29342,N_29244);
or UO_1477 (O_1477,N_29318,N_29513);
or UO_1478 (O_1478,N_29246,N_29852);
or UO_1479 (O_1479,N_28846,N_28800);
nor UO_1480 (O_1480,N_28810,N_29566);
or UO_1481 (O_1481,N_29324,N_29771);
nand UO_1482 (O_1482,N_29970,N_29705);
nand UO_1483 (O_1483,N_29670,N_28963);
and UO_1484 (O_1484,N_29164,N_29647);
nor UO_1485 (O_1485,N_29830,N_29850);
and UO_1486 (O_1486,N_28905,N_29982);
or UO_1487 (O_1487,N_28923,N_29346);
nand UO_1488 (O_1488,N_29284,N_29512);
nand UO_1489 (O_1489,N_29045,N_29155);
and UO_1490 (O_1490,N_29144,N_29096);
nand UO_1491 (O_1491,N_29364,N_29092);
nor UO_1492 (O_1492,N_29027,N_28998);
nand UO_1493 (O_1493,N_29844,N_29755);
or UO_1494 (O_1494,N_29462,N_29629);
or UO_1495 (O_1495,N_28931,N_28818);
nand UO_1496 (O_1496,N_28929,N_28843);
nand UO_1497 (O_1497,N_29648,N_29546);
and UO_1498 (O_1498,N_29012,N_29497);
nor UO_1499 (O_1499,N_29930,N_29630);
nand UO_1500 (O_1500,N_29952,N_29740);
xnor UO_1501 (O_1501,N_29443,N_29995);
or UO_1502 (O_1502,N_29947,N_28875);
xnor UO_1503 (O_1503,N_29429,N_28884);
nand UO_1504 (O_1504,N_28941,N_28963);
and UO_1505 (O_1505,N_29641,N_29408);
nor UO_1506 (O_1506,N_29050,N_28964);
or UO_1507 (O_1507,N_29165,N_29302);
or UO_1508 (O_1508,N_29744,N_28842);
nor UO_1509 (O_1509,N_29016,N_29633);
and UO_1510 (O_1510,N_29270,N_29161);
and UO_1511 (O_1511,N_29788,N_29303);
nor UO_1512 (O_1512,N_29002,N_29845);
xnor UO_1513 (O_1513,N_29454,N_29587);
xor UO_1514 (O_1514,N_29519,N_29176);
or UO_1515 (O_1515,N_28985,N_29696);
nor UO_1516 (O_1516,N_29849,N_29346);
nand UO_1517 (O_1517,N_29393,N_29461);
nor UO_1518 (O_1518,N_29877,N_29642);
nand UO_1519 (O_1519,N_29983,N_29984);
and UO_1520 (O_1520,N_29683,N_28983);
nand UO_1521 (O_1521,N_28888,N_29580);
nand UO_1522 (O_1522,N_29183,N_29091);
nand UO_1523 (O_1523,N_29925,N_29450);
and UO_1524 (O_1524,N_28978,N_29488);
nand UO_1525 (O_1525,N_28987,N_29816);
xnor UO_1526 (O_1526,N_29137,N_29098);
and UO_1527 (O_1527,N_29698,N_29344);
nor UO_1528 (O_1528,N_29099,N_29142);
nor UO_1529 (O_1529,N_29699,N_29256);
nand UO_1530 (O_1530,N_28908,N_29924);
xor UO_1531 (O_1531,N_29709,N_29137);
nor UO_1532 (O_1532,N_29052,N_28939);
and UO_1533 (O_1533,N_29664,N_29980);
and UO_1534 (O_1534,N_29917,N_29569);
nor UO_1535 (O_1535,N_29478,N_29630);
xnor UO_1536 (O_1536,N_29947,N_29064);
nand UO_1537 (O_1537,N_29569,N_29411);
xor UO_1538 (O_1538,N_29339,N_28897);
and UO_1539 (O_1539,N_29058,N_29146);
or UO_1540 (O_1540,N_28989,N_29420);
xor UO_1541 (O_1541,N_29361,N_29372);
and UO_1542 (O_1542,N_29715,N_29349);
nand UO_1543 (O_1543,N_29000,N_28921);
nor UO_1544 (O_1544,N_28972,N_29347);
nand UO_1545 (O_1545,N_28919,N_29417);
nor UO_1546 (O_1546,N_29801,N_28998);
or UO_1547 (O_1547,N_28936,N_28961);
or UO_1548 (O_1548,N_28928,N_28986);
nor UO_1549 (O_1549,N_29022,N_29789);
or UO_1550 (O_1550,N_29831,N_29982);
xnor UO_1551 (O_1551,N_29737,N_29231);
nand UO_1552 (O_1552,N_29484,N_29518);
nor UO_1553 (O_1553,N_29889,N_29768);
nor UO_1554 (O_1554,N_29468,N_29664);
nand UO_1555 (O_1555,N_28945,N_28883);
nor UO_1556 (O_1556,N_28910,N_29210);
xor UO_1557 (O_1557,N_28865,N_29032);
nand UO_1558 (O_1558,N_29971,N_28841);
nand UO_1559 (O_1559,N_29249,N_29368);
nand UO_1560 (O_1560,N_28865,N_28930);
nor UO_1561 (O_1561,N_29061,N_29849);
and UO_1562 (O_1562,N_29210,N_28961);
nor UO_1563 (O_1563,N_29800,N_29464);
xnor UO_1564 (O_1564,N_29903,N_29305);
xnor UO_1565 (O_1565,N_29186,N_29377);
and UO_1566 (O_1566,N_29935,N_29147);
nand UO_1567 (O_1567,N_28875,N_29886);
and UO_1568 (O_1568,N_29443,N_29359);
nand UO_1569 (O_1569,N_29953,N_29848);
nand UO_1570 (O_1570,N_29221,N_29091);
and UO_1571 (O_1571,N_29513,N_28965);
xor UO_1572 (O_1572,N_29360,N_28939);
and UO_1573 (O_1573,N_29650,N_28920);
and UO_1574 (O_1574,N_29128,N_28914);
nor UO_1575 (O_1575,N_28832,N_29610);
nor UO_1576 (O_1576,N_29317,N_29865);
xnor UO_1577 (O_1577,N_29380,N_29860);
and UO_1578 (O_1578,N_29483,N_29862);
and UO_1579 (O_1579,N_29897,N_29030);
xor UO_1580 (O_1580,N_29461,N_29046);
or UO_1581 (O_1581,N_29803,N_28844);
and UO_1582 (O_1582,N_28893,N_29206);
nor UO_1583 (O_1583,N_29086,N_29357);
or UO_1584 (O_1584,N_29554,N_29480);
and UO_1585 (O_1585,N_29058,N_29874);
or UO_1586 (O_1586,N_29171,N_29438);
nor UO_1587 (O_1587,N_29003,N_29828);
xnor UO_1588 (O_1588,N_29942,N_29025);
nand UO_1589 (O_1589,N_29521,N_29633);
and UO_1590 (O_1590,N_28976,N_29694);
nand UO_1591 (O_1591,N_28970,N_29583);
nand UO_1592 (O_1592,N_29912,N_29443);
and UO_1593 (O_1593,N_29254,N_28847);
or UO_1594 (O_1594,N_28832,N_29203);
nor UO_1595 (O_1595,N_29317,N_28932);
or UO_1596 (O_1596,N_28925,N_29140);
nor UO_1597 (O_1597,N_29801,N_29012);
or UO_1598 (O_1598,N_29671,N_29312);
xor UO_1599 (O_1599,N_29477,N_29562);
and UO_1600 (O_1600,N_29767,N_29428);
nand UO_1601 (O_1601,N_28881,N_29762);
and UO_1602 (O_1602,N_29504,N_29009);
and UO_1603 (O_1603,N_29430,N_29893);
and UO_1604 (O_1604,N_29342,N_29164);
and UO_1605 (O_1605,N_29327,N_29958);
xor UO_1606 (O_1606,N_28828,N_28920);
xnor UO_1607 (O_1607,N_29561,N_29974);
nor UO_1608 (O_1608,N_29989,N_29347);
or UO_1609 (O_1609,N_29933,N_29231);
nor UO_1610 (O_1610,N_29783,N_29326);
xor UO_1611 (O_1611,N_29504,N_29810);
nor UO_1612 (O_1612,N_29407,N_29706);
and UO_1613 (O_1613,N_29595,N_29883);
nor UO_1614 (O_1614,N_28853,N_28905);
nor UO_1615 (O_1615,N_29923,N_29639);
or UO_1616 (O_1616,N_29701,N_29457);
xor UO_1617 (O_1617,N_28985,N_29689);
or UO_1618 (O_1618,N_29096,N_29502);
nand UO_1619 (O_1619,N_28886,N_29817);
nand UO_1620 (O_1620,N_29484,N_29403);
xnor UO_1621 (O_1621,N_29823,N_29627);
nor UO_1622 (O_1622,N_28995,N_29276);
nor UO_1623 (O_1623,N_29215,N_29556);
nand UO_1624 (O_1624,N_29684,N_29498);
nand UO_1625 (O_1625,N_29151,N_28872);
xor UO_1626 (O_1626,N_29904,N_28924);
or UO_1627 (O_1627,N_29142,N_29706);
nor UO_1628 (O_1628,N_29664,N_29709);
nand UO_1629 (O_1629,N_29670,N_29119);
nor UO_1630 (O_1630,N_29185,N_29529);
nand UO_1631 (O_1631,N_29242,N_29150);
or UO_1632 (O_1632,N_29370,N_29731);
and UO_1633 (O_1633,N_29524,N_29157);
nand UO_1634 (O_1634,N_29730,N_29526);
nand UO_1635 (O_1635,N_29006,N_29884);
nand UO_1636 (O_1636,N_28812,N_29349);
nor UO_1637 (O_1637,N_29443,N_28911);
nand UO_1638 (O_1638,N_28998,N_29106);
xnor UO_1639 (O_1639,N_29553,N_28827);
and UO_1640 (O_1640,N_28940,N_29822);
xor UO_1641 (O_1641,N_29508,N_29798);
xor UO_1642 (O_1642,N_29594,N_29059);
or UO_1643 (O_1643,N_29196,N_29329);
nand UO_1644 (O_1644,N_29558,N_29756);
nor UO_1645 (O_1645,N_29730,N_29835);
xnor UO_1646 (O_1646,N_28995,N_28980);
xor UO_1647 (O_1647,N_29664,N_29784);
and UO_1648 (O_1648,N_28982,N_28879);
nor UO_1649 (O_1649,N_28935,N_29064);
xnor UO_1650 (O_1650,N_29017,N_28957);
and UO_1651 (O_1651,N_28866,N_29589);
or UO_1652 (O_1652,N_29691,N_29980);
and UO_1653 (O_1653,N_29236,N_29225);
or UO_1654 (O_1654,N_29666,N_29256);
nand UO_1655 (O_1655,N_28957,N_29063);
xnor UO_1656 (O_1656,N_29698,N_28876);
or UO_1657 (O_1657,N_29550,N_29557);
nand UO_1658 (O_1658,N_29291,N_29909);
nand UO_1659 (O_1659,N_28867,N_29912);
xor UO_1660 (O_1660,N_29896,N_29878);
nor UO_1661 (O_1661,N_29327,N_29340);
nand UO_1662 (O_1662,N_29836,N_29292);
or UO_1663 (O_1663,N_29100,N_29332);
nand UO_1664 (O_1664,N_29884,N_29162);
nor UO_1665 (O_1665,N_29459,N_29750);
xor UO_1666 (O_1666,N_29918,N_29928);
or UO_1667 (O_1667,N_29222,N_29090);
xnor UO_1668 (O_1668,N_29700,N_29081);
xor UO_1669 (O_1669,N_29571,N_29342);
nor UO_1670 (O_1670,N_29798,N_29286);
and UO_1671 (O_1671,N_29302,N_29448);
and UO_1672 (O_1672,N_29452,N_29940);
and UO_1673 (O_1673,N_29930,N_29843);
nand UO_1674 (O_1674,N_29653,N_29765);
nand UO_1675 (O_1675,N_29526,N_29304);
nor UO_1676 (O_1676,N_29244,N_28925);
nand UO_1677 (O_1677,N_29178,N_29937);
or UO_1678 (O_1678,N_29152,N_29542);
and UO_1679 (O_1679,N_29620,N_28916);
nor UO_1680 (O_1680,N_29426,N_28811);
nor UO_1681 (O_1681,N_29588,N_29384);
xnor UO_1682 (O_1682,N_29603,N_28820);
xnor UO_1683 (O_1683,N_29690,N_29873);
nand UO_1684 (O_1684,N_29053,N_29510);
nand UO_1685 (O_1685,N_28803,N_29434);
and UO_1686 (O_1686,N_29281,N_29128);
and UO_1687 (O_1687,N_29826,N_29590);
xnor UO_1688 (O_1688,N_29327,N_29229);
and UO_1689 (O_1689,N_29585,N_29062);
xnor UO_1690 (O_1690,N_28838,N_28930);
nor UO_1691 (O_1691,N_29988,N_29066);
nor UO_1692 (O_1692,N_29698,N_29771);
xor UO_1693 (O_1693,N_29582,N_28871);
nand UO_1694 (O_1694,N_29549,N_29196);
nor UO_1695 (O_1695,N_29619,N_29976);
nor UO_1696 (O_1696,N_29006,N_29183);
xnor UO_1697 (O_1697,N_29788,N_29363);
or UO_1698 (O_1698,N_29289,N_29163);
nor UO_1699 (O_1699,N_28861,N_29127);
or UO_1700 (O_1700,N_29910,N_29045);
xor UO_1701 (O_1701,N_29161,N_29352);
nor UO_1702 (O_1702,N_29101,N_29377);
and UO_1703 (O_1703,N_29747,N_29316);
nand UO_1704 (O_1704,N_29320,N_29068);
and UO_1705 (O_1705,N_29777,N_29096);
and UO_1706 (O_1706,N_29222,N_29414);
and UO_1707 (O_1707,N_29223,N_28953);
nor UO_1708 (O_1708,N_29773,N_29235);
nor UO_1709 (O_1709,N_29066,N_28808);
xor UO_1710 (O_1710,N_29529,N_29315);
or UO_1711 (O_1711,N_29792,N_29705);
and UO_1712 (O_1712,N_28914,N_29517);
nor UO_1713 (O_1713,N_28947,N_29091);
nand UO_1714 (O_1714,N_29785,N_29777);
and UO_1715 (O_1715,N_29296,N_29890);
nor UO_1716 (O_1716,N_29789,N_28897);
and UO_1717 (O_1717,N_29446,N_28866);
and UO_1718 (O_1718,N_28844,N_29352);
nand UO_1719 (O_1719,N_29026,N_29324);
nand UO_1720 (O_1720,N_29530,N_28849);
xor UO_1721 (O_1721,N_28832,N_29962);
nand UO_1722 (O_1722,N_29625,N_29901);
xnor UO_1723 (O_1723,N_29878,N_28819);
xor UO_1724 (O_1724,N_29192,N_29536);
nor UO_1725 (O_1725,N_29402,N_28998);
or UO_1726 (O_1726,N_29813,N_29122);
and UO_1727 (O_1727,N_29536,N_29626);
nor UO_1728 (O_1728,N_28962,N_29061);
and UO_1729 (O_1729,N_29932,N_29542);
and UO_1730 (O_1730,N_29479,N_29271);
and UO_1731 (O_1731,N_29450,N_29669);
nand UO_1732 (O_1732,N_29457,N_28865);
or UO_1733 (O_1733,N_29516,N_29463);
xnor UO_1734 (O_1734,N_29886,N_29569);
xor UO_1735 (O_1735,N_29470,N_29800);
xnor UO_1736 (O_1736,N_29114,N_29123);
nor UO_1737 (O_1737,N_29509,N_29532);
nand UO_1738 (O_1738,N_28895,N_29639);
nor UO_1739 (O_1739,N_29001,N_28986);
xor UO_1740 (O_1740,N_29528,N_28835);
nand UO_1741 (O_1741,N_29642,N_29955);
and UO_1742 (O_1742,N_29481,N_29235);
xor UO_1743 (O_1743,N_29690,N_28953);
nor UO_1744 (O_1744,N_29265,N_29987);
or UO_1745 (O_1745,N_29032,N_29006);
xor UO_1746 (O_1746,N_28947,N_28910);
or UO_1747 (O_1747,N_29595,N_29926);
xnor UO_1748 (O_1748,N_29431,N_29964);
xor UO_1749 (O_1749,N_29067,N_29665);
xor UO_1750 (O_1750,N_29503,N_29725);
nand UO_1751 (O_1751,N_29251,N_28878);
nor UO_1752 (O_1752,N_29120,N_29967);
or UO_1753 (O_1753,N_29021,N_29239);
nand UO_1754 (O_1754,N_29572,N_29459);
nand UO_1755 (O_1755,N_29389,N_29675);
and UO_1756 (O_1756,N_28928,N_29668);
or UO_1757 (O_1757,N_29618,N_29203);
nand UO_1758 (O_1758,N_29130,N_29538);
or UO_1759 (O_1759,N_29944,N_28907);
nor UO_1760 (O_1760,N_29117,N_29553);
nor UO_1761 (O_1761,N_29543,N_29007);
nand UO_1762 (O_1762,N_29380,N_29540);
and UO_1763 (O_1763,N_29574,N_28807);
nand UO_1764 (O_1764,N_29018,N_28804);
xor UO_1765 (O_1765,N_28853,N_29871);
or UO_1766 (O_1766,N_29942,N_28888);
xor UO_1767 (O_1767,N_29852,N_29631);
xor UO_1768 (O_1768,N_29133,N_29588);
nor UO_1769 (O_1769,N_28996,N_29718);
nor UO_1770 (O_1770,N_29821,N_29360);
nor UO_1771 (O_1771,N_29960,N_28814);
or UO_1772 (O_1772,N_29956,N_29812);
xnor UO_1773 (O_1773,N_28985,N_29215);
nand UO_1774 (O_1774,N_29769,N_29915);
nand UO_1775 (O_1775,N_29435,N_29084);
xnor UO_1776 (O_1776,N_29442,N_29933);
or UO_1777 (O_1777,N_29949,N_29442);
and UO_1778 (O_1778,N_29502,N_29245);
xnor UO_1779 (O_1779,N_28858,N_29814);
and UO_1780 (O_1780,N_29730,N_29606);
nor UO_1781 (O_1781,N_29508,N_29560);
and UO_1782 (O_1782,N_28963,N_29411);
and UO_1783 (O_1783,N_29892,N_29603);
nand UO_1784 (O_1784,N_29794,N_29002);
nand UO_1785 (O_1785,N_29217,N_29144);
or UO_1786 (O_1786,N_29466,N_29782);
nand UO_1787 (O_1787,N_29155,N_29550);
or UO_1788 (O_1788,N_29076,N_29308);
xnor UO_1789 (O_1789,N_29705,N_29737);
and UO_1790 (O_1790,N_29956,N_29794);
or UO_1791 (O_1791,N_29100,N_29414);
xor UO_1792 (O_1792,N_29653,N_29172);
or UO_1793 (O_1793,N_29442,N_29415);
nand UO_1794 (O_1794,N_29107,N_29370);
and UO_1795 (O_1795,N_29914,N_29925);
and UO_1796 (O_1796,N_29772,N_29627);
or UO_1797 (O_1797,N_29622,N_28942);
nand UO_1798 (O_1798,N_29434,N_29284);
nand UO_1799 (O_1799,N_29141,N_29932);
and UO_1800 (O_1800,N_29140,N_29014);
or UO_1801 (O_1801,N_29070,N_29292);
xor UO_1802 (O_1802,N_29412,N_29649);
nor UO_1803 (O_1803,N_28974,N_28940);
and UO_1804 (O_1804,N_29375,N_28952);
nand UO_1805 (O_1805,N_28822,N_28950);
or UO_1806 (O_1806,N_29946,N_29799);
xnor UO_1807 (O_1807,N_28900,N_29197);
or UO_1808 (O_1808,N_29210,N_29035);
nor UO_1809 (O_1809,N_28942,N_28946);
or UO_1810 (O_1810,N_29739,N_29014);
nand UO_1811 (O_1811,N_29612,N_29346);
nand UO_1812 (O_1812,N_29613,N_29112);
xor UO_1813 (O_1813,N_29630,N_28963);
or UO_1814 (O_1814,N_29246,N_29977);
and UO_1815 (O_1815,N_29016,N_29511);
xnor UO_1816 (O_1816,N_29453,N_28889);
nand UO_1817 (O_1817,N_28885,N_29402);
nor UO_1818 (O_1818,N_29149,N_29191);
xnor UO_1819 (O_1819,N_28874,N_29343);
nor UO_1820 (O_1820,N_28979,N_29590);
nor UO_1821 (O_1821,N_29754,N_29290);
and UO_1822 (O_1822,N_29843,N_29923);
or UO_1823 (O_1823,N_29809,N_29255);
nand UO_1824 (O_1824,N_29885,N_29054);
and UO_1825 (O_1825,N_29174,N_28934);
and UO_1826 (O_1826,N_29015,N_29203);
nor UO_1827 (O_1827,N_29311,N_29572);
and UO_1828 (O_1828,N_29036,N_28823);
nand UO_1829 (O_1829,N_29078,N_29114);
nand UO_1830 (O_1830,N_28911,N_29986);
xnor UO_1831 (O_1831,N_28951,N_29480);
or UO_1832 (O_1832,N_29294,N_29511);
nor UO_1833 (O_1833,N_28909,N_28907);
xor UO_1834 (O_1834,N_28935,N_29469);
xor UO_1835 (O_1835,N_29017,N_29389);
xnor UO_1836 (O_1836,N_29820,N_29848);
and UO_1837 (O_1837,N_29322,N_29017);
nor UO_1838 (O_1838,N_29198,N_28994);
xnor UO_1839 (O_1839,N_28946,N_28952);
nand UO_1840 (O_1840,N_29923,N_29849);
and UO_1841 (O_1841,N_29285,N_28977);
nor UO_1842 (O_1842,N_29380,N_29836);
and UO_1843 (O_1843,N_29359,N_29795);
xor UO_1844 (O_1844,N_29791,N_29276);
or UO_1845 (O_1845,N_28823,N_29097);
and UO_1846 (O_1846,N_28838,N_29964);
nand UO_1847 (O_1847,N_29991,N_29353);
xnor UO_1848 (O_1848,N_29467,N_29219);
nor UO_1849 (O_1849,N_29614,N_29268);
nand UO_1850 (O_1850,N_29178,N_29308);
or UO_1851 (O_1851,N_29804,N_29099);
xnor UO_1852 (O_1852,N_29641,N_29935);
or UO_1853 (O_1853,N_29809,N_29136);
xor UO_1854 (O_1854,N_28903,N_28992);
and UO_1855 (O_1855,N_29347,N_28905);
nand UO_1856 (O_1856,N_29340,N_29731);
nor UO_1857 (O_1857,N_29663,N_28894);
and UO_1858 (O_1858,N_29550,N_29032);
nor UO_1859 (O_1859,N_29118,N_29611);
or UO_1860 (O_1860,N_29847,N_29649);
nor UO_1861 (O_1861,N_28837,N_29123);
or UO_1862 (O_1862,N_29362,N_29824);
and UO_1863 (O_1863,N_28936,N_29428);
nor UO_1864 (O_1864,N_28963,N_29161);
nand UO_1865 (O_1865,N_29389,N_29678);
xnor UO_1866 (O_1866,N_29303,N_29232);
and UO_1867 (O_1867,N_29274,N_29200);
nand UO_1868 (O_1868,N_29064,N_29192);
nand UO_1869 (O_1869,N_29373,N_29737);
and UO_1870 (O_1870,N_29716,N_28920);
nand UO_1871 (O_1871,N_29570,N_29130);
nand UO_1872 (O_1872,N_29192,N_29116);
or UO_1873 (O_1873,N_29494,N_29845);
nand UO_1874 (O_1874,N_29260,N_29954);
and UO_1875 (O_1875,N_29470,N_29447);
and UO_1876 (O_1876,N_29970,N_29383);
xnor UO_1877 (O_1877,N_28809,N_29525);
xnor UO_1878 (O_1878,N_29403,N_29390);
nand UO_1879 (O_1879,N_28944,N_29578);
nor UO_1880 (O_1880,N_29714,N_29730);
nand UO_1881 (O_1881,N_28840,N_29993);
and UO_1882 (O_1882,N_29303,N_29827);
and UO_1883 (O_1883,N_29136,N_29371);
nor UO_1884 (O_1884,N_29746,N_29831);
nand UO_1885 (O_1885,N_29041,N_29598);
xor UO_1886 (O_1886,N_29016,N_29711);
and UO_1887 (O_1887,N_29413,N_29194);
nand UO_1888 (O_1888,N_29358,N_29821);
xnor UO_1889 (O_1889,N_29249,N_29851);
nor UO_1890 (O_1890,N_29395,N_29935);
nand UO_1891 (O_1891,N_29908,N_29493);
and UO_1892 (O_1892,N_29250,N_29442);
or UO_1893 (O_1893,N_29497,N_29097);
nor UO_1894 (O_1894,N_29591,N_29366);
nor UO_1895 (O_1895,N_28824,N_29525);
and UO_1896 (O_1896,N_29046,N_29710);
and UO_1897 (O_1897,N_28899,N_29433);
and UO_1898 (O_1898,N_29313,N_29435);
nand UO_1899 (O_1899,N_29050,N_28848);
or UO_1900 (O_1900,N_29304,N_29367);
or UO_1901 (O_1901,N_29146,N_29626);
and UO_1902 (O_1902,N_29196,N_29785);
nand UO_1903 (O_1903,N_29983,N_29353);
or UO_1904 (O_1904,N_29282,N_29308);
nor UO_1905 (O_1905,N_29850,N_29932);
nand UO_1906 (O_1906,N_29876,N_29864);
nor UO_1907 (O_1907,N_29712,N_29743);
xor UO_1908 (O_1908,N_28865,N_29714);
and UO_1909 (O_1909,N_28831,N_29316);
nor UO_1910 (O_1910,N_29573,N_29861);
xor UO_1911 (O_1911,N_29488,N_28952);
nor UO_1912 (O_1912,N_29623,N_29915);
nor UO_1913 (O_1913,N_29627,N_28974);
and UO_1914 (O_1914,N_28810,N_29579);
nor UO_1915 (O_1915,N_29702,N_29591);
xor UO_1916 (O_1916,N_29084,N_28848);
xor UO_1917 (O_1917,N_29319,N_29776);
nand UO_1918 (O_1918,N_29454,N_29052);
and UO_1919 (O_1919,N_29025,N_29663);
and UO_1920 (O_1920,N_29344,N_29870);
xnor UO_1921 (O_1921,N_29469,N_29347);
nand UO_1922 (O_1922,N_28855,N_29059);
xor UO_1923 (O_1923,N_28961,N_29866);
or UO_1924 (O_1924,N_29435,N_29966);
nand UO_1925 (O_1925,N_29176,N_29683);
xor UO_1926 (O_1926,N_28842,N_29502);
nor UO_1927 (O_1927,N_29861,N_28961);
xnor UO_1928 (O_1928,N_28851,N_29604);
nand UO_1929 (O_1929,N_29822,N_28847);
xor UO_1930 (O_1930,N_29436,N_29326);
and UO_1931 (O_1931,N_29248,N_28847);
nor UO_1932 (O_1932,N_29292,N_29099);
or UO_1933 (O_1933,N_28885,N_29832);
xnor UO_1934 (O_1934,N_29441,N_29902);
and UO_1935 (O_1935,N_29735,N_29522);
or UO_1936 (O_1936,N_29465,N_29930);
and UO_1937 (O_1937,N_29759,N_28889);
and UO_1938 (O_1938,N_29903,N_29131);
nor UO_1939 (O_1939,N_29176,N_29555);
or UO_1940 (O_1940,N_29626,N_29871);
or UO_1941 (O_1941,N_29660,N_29680);
xor UO_1942 (O_1942,N_29976,N_29931);
and UO_1943 (O_1943,N_29381,N_29241);
and UO_1944 (O_1944,N_29286,N_29190);
nor UO_1945 (O_1945,N_29297,N_29900);
or UO_1946 (O_1946,N_29049,N_29521);
nor UO_1947 (O_1947,N_29282,N_29279);
or UO_1948 (O_1948,N_29954,N_29144);
nor UO_1949 (O_1949,N_29936,N_29259);
or UO_1950 (O_1950,N_29751,N_29957);
xnor UO_1951 (O_1951,N_29542,N_29914);
nand UO_1952 (O_1952,N_29546,N_29520);
or UO_1953 (O_1953,N_29183,N_29524);
or UO_1954 (O_1954,N_29462,N_29099);
and UO_1955 (O_1955,N_29340,N_29687);
xor UO_1956 (O_1956,N_28842,N_29784);
nand UO_1957 (O_1957,N_29525,N_29909);
and UO_1958 (O_1958,N_29630,N_29614);
nand UO_1959 (O_1959,N_29153,N_29635);
xor UO_1960 (O_1960,N_29368,N_29558);
nand UO_1961 (O_1961,N_29731,N_29925);
nor UO_1962 (O_1962,N_28836,N_29004);
nand UO_1963 (O_1963,N_28979,N_29253);
nor UO_1964 (O_1964,N_29431,N_28827);
xor UO_1965 (O_1965,N_29579,N_29967);
nor UO_1966 (O_1966,N_29091,N_29713);
nor UO_1967 (O_1967,N_29977,N_29241);
or UO_1968 (O_1968,N_29416,N_29560);
nor UO_1969 (O_1969,N_29495,N_28810);
and UO_1970 (O_1970,N_29157,N_29319);
nor UO_1971 (O_1971,N_29749,N_29091);
nand UO_1972 (O_1972,N_28924,N_29068);
or UO_1973 (O_1973,N_28917,N_29878);
nand UO_1974 (O_1974,N_29351,N_29202);
nand UO_1975 (O_1975,N_29763,N_29276);
nor UO_1976 (O_1976,N_29290,N_29430);
nor UO_1977 (O_1977,N_28892,N_29739);
nand UO_1978 (O_1978,N_29975,N_28924);
nor UO_1979 (O_1979,N_28992,N_29882);
nor UO_1980 (O_1980,N_29456,N_29450);
nand UO_1981 (O_1981,N_29947,N_28922);
nand UO_1982 (O_1982,N_28927,N_29617);
nand UO_1983 (O_1983,N_29613,N_29128);
and UO_1984 (O_1984,N_29897,N_29108);
nor UO_1985 (O_1985,N_28907,N_29585);
or UO_1986 (O_1986,N_29310,N_29602);
xor UO_1987 (O_1987,N_29083,N_29909);
or UO_1988 (O_1988,N_29367,N_29624);
nor UO_1989 (O_1989,N_29199,N_28977);
nand UO_1990 (O_1990,N_29743,N_28984);
nor UO_1991 (O_1991,N_29889,N_29488);
nor UO_1992 (O_1992,N_29617,N_29910);
and UO_1993 (O_1993,N_29822,N_28885);
nand UO_1994 (O_1994,N_29236,N_29137);
or UO_1995 (O_1995,N_29141,N_29000);
or UO_1996 (O_1996,N_28902,N_29867);
nand UO_1997 (O_1997,N_28841,N_28991);
and UO_1998 (O_1998,N_28805,N_29305);
or UO_1999 (O_1999,N_29010,N_29760);
xor UO_2000 (O_2000,N_29491,N_28992);
and UO_2001 (O_2001,N_29679,N_29592);
xor UO_2002 (O_2002,N_29669,N_29363);
and UO_2003 (O_2003,N_29341,N_28816);
and UO_2004 (O_2004,N_29522,N_28897);
nor UO_2005 (O_2005,N_28861,N_29918);
nand UO_2006 (O_2006,N_29593,N_29695);
or UO_2007 (O_2007,N_29580,N_29425);
nand UO_2008 (O_2008,N_29429,N_29197);
or UO_2009 (O_2009,N_29947,N_29683);
nor UO_2010 (O_2010,N_29179,N_29131);
nor UO_2011 (O_2011,N_29131,N_29180);
or UO_2012 (O_2012,N_29680,N_29278);
nand UO_2013 (O_2013,N_29867,N_29726);
and UO_2014 (O_2014,N_29517,N_29078);
or UO_2015 (O_2015,N_29145,N_28927);
nor UO_2016 (O_2016,N_28974,N_29169);
nor UO_2017 (O_2017,N_29399,N_29854);
nand UO_2018 (O_2018,N_29118,N_29608);
xor UO_2019 (O_2019,N_28881,N_29536);
or UO_2020 (O_2020,N_29333,N_29945);
xor UO_2021 (O_2021,N_28988,N_29132);
nor UO_2022 (O_2022,N_29096,N_29921);
and UO_2023 (O_2023,N_29744,N_29204);
nand UO_2024 (O_2024,N_29332,N_29758);
nand UO_2025 (O_2025,N_29646,N_29692);
nand UO_2026 (O_2026,N_29131,N_29547);
and UO_2027 (O_2027,N_29535,N_29166);
and UO_2028 (O_2028,N_29446,N_29240);
xor UO_2029 (O_2029,N_29068,N_29918);
and UO_2030 (O_2030,N_29937,N_29639);
xor UO_2031 (O_2031,N_29297,N_28957);
nor UO_2032 (O_2032,N_29957,N_29532);
or UO_2033 (O_2033,N_29393,N_29968);
xnor UO_2034 (O_2034,N_29104,N_28889);
or UO_2035 (O_2035,N_29896,N_29544);
nor UO_2036 (O_2036,N_28926,N_29519);
and UO_2037 (O_2037,N_29634,N_29901);
nor UO_2038 (O_2038,N_29864,N_29257);
and UO_2039 (O_2039,N_29346,N_29624);
nor UO_2040 (O_2040,N_29598,N_28896);
nand UO_2041 (O_2041,N_29272,N_29560);
or UO_2042 (O_2042,N_29776,N_28835);
or UO_2043 (O_2043,N_29356,N_28887);
or UO_2044 (O_2044,N_29760,N_29032);
or UO_2045 (O_2045,N_29356,N_29850);
or UO_2046 (O_2046,N_29510,N_29586);
or UO_2047 (O_2047,N_29922,N_29266);
nand UO_2048 (O_2048,N_29356,N_29943);
xnor UO_2049 (O_2049,N_29376,N_29214);
xor UO_2050 (O_2050,N_29203,N_29840);
or UO_2051 (O_2051,N_29710,N_29748);
nand UO_2052 (O_2052,N_29095,N_29802);
nor UO_2053 (O_2053,N_29411,N_29116);
nand UO_2054 (O_2054,N_28868,N_29595);
or UO_2055 (O_2055,N_29340,N_29161);
and UO_2056 (O_2056,N_29482,N_28971);
xor UO_2057 (O_2057,N_29613,N_29101);
and UO_2058 (O_2058,N_29543,N_28851);
or UO_2059 (O_2059,N_29781,N_29960);
xnor UO_2060 (O_2060,N_29753,N_28802);
or UO_2061 (O_2061,N_29599,N_29536);
nand UO_2062 (O_2062,N_29700,N_29095);
nor UO_2063 (O_2063,N_29470,N_29414);
xor UO_2064 (O_2064,N_29460,N_29795);
nor UO_2065 (O_2065,N_29874,N_29682);
or UO_2066 (O_2066,N_29985,N_29344);
xor UO_2067 (O_2067,N_29826,N_29919);
or UO_2068 (O_2068,N_29241,N_28818);
nor UO_2069 (O_2069,N_29661,N_29943);
or UO_2070 (O_2070,N_29574,N_28993);
nand UO_2071 (O_2071,N_29424,N_29853);
nand UO_2072 (O_2072,N_28865,N_29174);
xor UO_2073 (O_2073,N_29951,N_29688);
xor UO_2074 (O_2074,N_29385,N_29188);
and UO_2075 (O_2075,N_29012,N_29593);
and UO_2076 (O_2076,N_29990,N_29236);
nor UO_2077 (O_2077,N_29621,N_29012);
or UO_2078 (O_2078,N_29278,N_29308);
nor UO_2079 (O_2079,N_28962,N_29864);
nand UO_2080 (O_2080,N_28938,N_29304);
nor UO_2081 (O_2081,N_29066,N_29896);
xor UO_2082 (O_2082,N_29580,N_29791);
and UO_2083 (O_2083,N_29433,N_29187);
xor UO_2084 (O_2084,N_28849,N_29546);
xnor UO_2085 (O_2085,N_29629,N_29749);
nor UO_2086 (O_2086,N_28955,N_29146);
or UO_2087 (O_2087,N_29474,N_29638);
nand UO_2088 (O_2088,N_29512,N_29841);
nand UO_2089 (O_2089,N_29021,N_29194);
nor UO_2090 (O_2090,N_29410,N_29875);
nor UO_2091 (O_2091,N_29088,N_29364);
xnor UO_2092 (O_2092,N_28903,N_29705);
nor UO_2093 (O_2093,N_29865,N_29299);
nand UO_2094 (O_2094,N_29876,N_29651);
and UO_2095 (O_2095,N_29833,N_29080);
nor UO_2096 (O_2096,N_29843,N_29295);
and UO_2097 (O_2097,N_29887,N_29705);
nand UO_2098 (O_2098,N_29616,N_29868);
or UO_2099 (O_2099,N_29783,N_28810);
nand UO_2100 (O_2100,N_29619,N_29648);
or UO_2101 (O_2101,N_29024,N_28991);
xor UO_2102 (O_2102,N_29958,N_29503);
and UO_2103 (O_2103,N_29720,N_29131);
nor UO_2104 (O_2104,N_29055,N_29541);
nor UO_2105 (O_2105,N_29003,N_28999);
xor UO_2106 (O_2106,N_28966,N_29563);
nor UO_2107 (O_2107,N_29542,N_29356);
or UO_2108 (O_2108,N_29904,N_29712);
nand UO_2109 (O_2109,N_29869,N_29936);
xor UO_2110 (O_2110,N_29163,N_29735);
and UO_2111 (O_2111,N_29717,N_29017);
xor UO_2112 (O_2112,N_29230,N_29127);
nor UO_2113 (O_2113,N_28947,N_29063);
and UO_2114 (O_2114,N_28801,N_29835);
and UO_2115 (O_2115,N_29813,N_29552);
nor UO_2116 (O_2116,N_29555,N_29145);
nand UO_2117 (O_2117,N_29602,N_29047);
and UO_2118 (O_2118,N_29584,N_29306);
nor UO_2119 (O_2119,N_29685,N_29158);
nor UO_2120 (O_2120,N_29672,N_29934);
or UO_2121 (O_2121,N_29863,N_29184);
xor UO_2122 (O_2122,N_28954,N_29179);
xnor UO_2123 (O_2123,N_29513,N_29354);
or UO_2124 (O_2124,N_29047,N_29134);
xnor UO_2125 (O_2125,N_29995,N_29054);
nand UO_2126 (O_2126,N_29255,N_28927);
nor UO_2127 (O_2127,N_29993,N_29457);
xor UO_2128 (O_2128,N_29269,N_29237);
or UO_2129 (O_2129,N_28946,N_29358);
or UO_2130 (O_2130,N_28820,N_28927);
xnor UO_2131 (O_2131,N_29080,N_28806);
and UO_2132 (O_2132,N_29728,N_28866);
xnor UO_2133 (O_2133,N_29908,N_29249);
xor UO_2134 (O_2134,N_28888,N_28860);
xnor UO_2135 (O_2135,N_28837,N_29024);
and UO_2136 (O_2136,N_28982,N_29854);
or UO_2137 (O_2137,N_29821,N_29717);
nand UO_2138 (O_2138,N_29780,N_28982);
nand UO_2139 (O_2139,N_29502,N_29714);
nand UO_2140 (O_2140,N_28997,N_29590);
nor UO_2141 (O_2141,N_29384,N_29409);
nand UO_2142 (O_2142,N_28803,N_29393);
and UO_2143 (O_2143,N_29391,N_29140);
nor UO_2144 (O_2144,N_29996,N_29855);
and UO_2145 (O_2145,N_29541,N_29567);
nand UO_2146 (O_2146,N_29284,N_29805);
xnor UO_2147 (O_2147,N_29039,N_29215);
or UO_2148 (O_2148,N_29970,N_29980);
and UO_2149 (O_2149,N_29265,N_29136);
nand UO_2150 (O_2150,N_29243,N_29324);
or UO_2151 (O_2151,N_28813,N_28901);
and UO_2152 (O_2152,N_29560,N_29189);
xnor UO_2153 (O_2153,N_29601,N_29970);
and UO_2154 (O_2154,N_29913,N_29116);
or UO_2155 (O_2155,N_29581,N_29469);
nor UO_2156 (O_2156,N_29346,N_29951);
and UO_2157 (O_2157,N_29858,N_29428);
nor UO_2158 (O_2158,N_29424,N_29981);
xor UO_2159 (O_2159,N_29898,N_29762);
xnor UO_2160 (O_2160,N_29890,N_29751);
nand UO_2161 (O_2161,N_29466,N_29813);
xor UO_2162 (O_2162,N_29212,N_28855);
nand UO_2163 (O_2163,N_29433,N_29843);
xnor UO_2164 (O_2164,N_29922,N_29035);
nand UO_2165 (O_2165,N_29442,N_29426);
nor UO_2166 (O_2166,N_29490,N_28949);
xor UO_2167 (O_2167,N_29937,N_29881);
xor UO_2168 (O_2168,N_29663,N_28852);
nor UO_2169 (O_2169,N_28833,N_29650);
and UO_2170 (O_2170,N_29100,N_28857);
or UO_2171 (O_2171,N_29437,N_28989);
nor UO_2172 (O_2172,N_28994,N_29511);
nand UO_2173 (O_2173,N_29342,N_28974);
nand UO_2174 (O_2174,N_29178,N_29023);
or UO_2175 (O_2175,N_28951,N_29157);
xnor UO_2176 (O_2176,N_29293,N_29687);
or UO_2177 (O_2177,N_28930,N_29903);
nand UO_2178 (O_2178,N_29781,N_28888);
nor UO_2179 (O_2179,N_29613,N_29151);
xnor UO_2180 (O_2180,N_29724,N_29342);
nand UO_2181 (O_2181,N_29953,N_29722);
nand UO_2182 (O_2182,N_29021,N_29592);
nor UO_2183 (O_2183,N_29854,N_29058);
nor UO_2184 (O_2184,N_29465,N_29374);
nor UO_2185 (O_2185,N_29495,N_28896);
and UO_2186 (O_2186,N_29140,N_29620);
xor UO_2187 (O_2187,N_29470,N_29051);
xor UO_2188 (O_2188,N_29245,N_28815);
xor UO_2189 (O_2189,N_29263,N_29003);
nor UO_2190 (O_2190,N_29522,N_29482);
or UO_2191 (O_2191,N_29688,N_28881);
nand UO_2192 (O_2192,N_29438,N_29816);
nor UO_2193 (O_2193,N_29983,N_28855);
and UO_2194 (O_2194,N_29895,N_29527);
and UO_2195 (O_2195,N_29874,N_28826);
nand UO_2196 (O_2196,N_28845,N_29332);
nand UO_2197 (O_2197,N_29854,N_28855);
nand UO_2198 (O_2198,N_29510,N_29483);
or UO_2199 (O_2199,N_29578,N_29812);
nand UO_2200 (O_2200,N_29289,N_29726);
or UO_2201 (O_2201,N_29047,N_29912);
xnor UO_2202 (O_2202,N_29214,N_29189);
nand UO_2203 (O_2203,N_29185,N_28950);
nor UO_2204 (O_2204,N_29773,N_29558);
nand UO_2205 (O_2205,N_29342,N_28856);
xnor UO_2206 (O_2206,N_29711,N_29125);
nor UO_2207 (O_2207,N_29148,N_29781);
nor UO_2208 (O_2208,N_29416,N_28845);
or UO_2209 (O_2209,N_29528,N_29533);
nand UO_2210 (O_2210,N_29213,N_28905);
nand UO_2211 (O_2211,N_29653,N_29075);
or UO_2212 (O_2212,N_29543,N_29829);
nand UO_2213 (O_2213,N_29267,N_29393);
or UO_2214 (O_2214,N_29365,N_29056);
xnor UO_2215 (O_2215,N_29838,N_29396);
nor UO_2216 (O_2216,N_29572,N_29780);
xnor UO_2217 (O_2217,N_29126,N_29147);
nor UO_2218 (O_2218,N_29898,N_29254);
or UO_2219 (O_2219,N_29700,N_29652);
or UO_2220 (O_2220,N_29395,N_28802);
or UO_2221 (O_2221,N_28984,N_29256);
nand UO_2222 (O_2222,N_29018,N_29198);
or UO_2223 (O_2223,N_29374,N_29362);
and UO_2224 (O_2224,N_28919,N_29462);
nor UO_2225 (O_2225,N_29995,N_29827);
nand UO_2226 (O_2226,N_29107,N_29676);
xor UO_2227 (O_2227,N_29071,N_29460);
or UO_2228 (O_2228,N_29471,N_29886);
xor UO_2229 (O_2229,N_29574,N_29509);
and UO_2230 (O_2230,N_29607,N_29411);
nor UO_2231 (O_2231,N_29956,N_29177);
xnor UO_2232 (O_2232,N_29954,N_28866);
or UO_2233 (O_2233,N_29092,N_29564);
and UO_2234 (O_2234,N_29108,N_28838);
and UO_2235 (O_2235,N_29630,N_29491);
nand UO_2236 (O_2236,N_29637,N_29270);
and UO_2237 (O_2237,N_29812,N_29888);
nor UO_2238 (O_2238,N_29552,N_29456);
or UO_2239 (O_2239,N_29341,N_28813);
and UO_2240 (O_2240,N_29519,N_29173);
and UO_2241 (O_2241,N_29538,N_28919);
xnor UO_2242 (O_2242,N_29815,N_29921);
nand UO_2243 (O_2243,N_29074,N_29516);
and UO_2244 (O_2244,N_29094,N_28921);
and UO_2245 (O_2245,N_29560,N_29391);
nand UO_2246 (O_2246,N_29083,N_29553);
nor UO_2247 (O_2247,N_29116,N_29191);
nand UO_2248 (O_2248,N_28976,N_29290);
nor UO_2249 (O_2249,N_29615,N_29786);
nor UO_2250 (O_2250,N_29325,N_28872);
xnor UO_2251 (O_2251,N_29956,N_29213);
xor UO_2252 (O_2252,N_29520,N_29154);
and UO_2253 (O_2253,N_29191,N_29016);
and UO_2254 (O_2254,N_29200,N_29195);
nor UO_2255 (O_2255,N_29115,N_29773);
and UO_2256 (O_2256,N_29297,N_29133);
xnor UO_2257 (O_2257,N_28972,N_29809);
xor UO_2258 (O_2258,N_29324,N_29731);
nor UO_2259 (O_2259,N_28998,N_29565);
nand UO_2260 (O_2260,N_29791,N_29698);
nand UO_2261 (O_2261,N_28967,N_29372);
and UO_2262 (O_2262,N_29603,N_29626);
and UO_2263 (O_2263,N_29594,N_29496);
and UO_2264 (O_2264,N_29031,N_28877);
nand UO_2265 (O_2265,N_29387,N_29849);
nand UO_2266 (O_2266,N_29596,N_29689);
nand UO_2267 (O_2267,N_28885,N_28995);
nor UO_2268 (O_2268,N_29327,N_28824);
or UO_2269 (O_2269,N_29609,N_29831);
nand UO_2270 (O_2270,N_29186,N_29666);
or UO_2271 (O_2271,N_29488,N_29951);
xnor UO_2272 (O_2272,N_28934,N_29392);
nand UO_2273 (O_2273,N_29173,N_29452);
nand UO_2274 (O_2274,N_28841,N_28978);
nor UO_2275 (O_2275,N_29268,N_28921);
or UO_2276 (O_2276,N_29890,N_29280);
nand UO_2277 (O_2277,N_29207,N_29342);
nor UO_2278 (O_2278,N_29151,N_29753);
and UO_2279 (O_2279,N_29063,N_29244);
nand UO_2280 (O_2280,N_28864,N_29658);
xnor UO_2281 (O_2281,N_29872,N_29464);
xnor UO_2282 (O_2282,N_29999,N_29755);
and UO_2283 (O_2283,N_28967,N_29718);
or UO_2284 (O_2284,N_29133,N_28916);
nand UO_2285 (O_2285,N_29047,N_29289);
nor UO_2286 (O_2286,N_29499,N_28861);
and UO_2287 (O_2287,N_29943,N_28863);
nand UO_2288 (O_2288,N_28849,N_29578);
or UO_2289 (O_2289,N_29679,N_28869);
or UO_2290 (O_2290,N_29609,N_29481);
xnor UO_2291 (O_2291,N_28946,N_29420);
nor UO_2292 (O_2292,N_28929,N_29889);
nor UO_2293 (O_2293,N_29232,N_29914);
nor UO_2294 (O_2294,N_29583,N_29697);
or UO_2295 (O_2295,N_29917,N_29799);
xnor UO_2296 (O_2296,N_29170,N_28831);
and UO_2297 (O_2297,N_29433,N_29887);
nor UO_2298 (O_2298,N_29210,N_29201);
nor UO_2299 (O_2299,N_28902,N_29812);
nor UO_2300 (O_2300,N_29845,N_29177);
and UO_2301 (O_2301,N_29814,N_29296);
nand UO_2302 (O_2302,N_29647,N_28895);
nand UO_2303 (O_2303,N_29749,N_29360);
nor UO_2304 (O_2304,N_29676,N_29129);
and UO_2305 (O_2305,N_28988,N_29109);
or UO_2306 (O_2306,N_29639,N_29528);
nor UO_2307 (O_2307,N_29571,N_29816);
and UO_2308 (O_2308,N_29108,N_29217);
or UO_2309 (O_2309,N_29659,N_29760);
or UO_2310 (O_2310,N_29098,N_29732);
nor UO_2311 (O_2311,N_29996,N_29086);
or UO_2312 (O_2312,N_28939,N_28957);
or UO_2313 (O_2313,N_29820,N_29774);
and UO_2314 (O_2314,N_29109,N_29952);
or UO_2315 (O_2315,N_29505,N_29424);
and UO_2316 (O_2316,N_29535,N_29248);
nand UO_2317 (O_2317,N_29034,N_29599);
and UO_2318 (O_2318,N_28909,N_29897);
nor UO_2319 (O_2319,N_29816,N_29815);
or UO_2320 (O_2320,N_29595,N_29194);
nand UO_2321 (O_2321,N_29321,N_28803);
nand UO_2322 (O_2322,N_28984,N_29711);
nor UO_2323 (O_2323,N_29860,N_29814);
nor UO_2324 (O_2324,N_29453,N_28988);
or UO_2325 (O_2325,N_28952,N_29819);
nor UO_2326 (O_2326,N_29660,N_28934);
or UO_2327 (O_2327,N_29775,N_29304);
nand UO_2328 (O_2328,N_29294,N_29949);
xor UO_2329 (O_2329,N_29326,N_29208);
xor UO_2330 (O_2330,N_29172,N_29343);
nor UO_2331 (O_2331,N_29799,N_29060);
and UO_2332 (O_2332,N_29061,N_29775);
nor UO_2333 (O_2333,N_29389,N_28808);
or UO_2334 (O_2334,N_29120,N_29696);
nand UO_2335 (O_2335,N_29560,N_29792);
nand UO_2336 (O_2336,N_29976,N_29616);
xor UO_2337 (O_2337,N_29387,N_29523);
or UO_2338 (O_2338,N_29549,N_28962);
xnor UO_2339 (O_2339,N_29797,N_29915);
or UO_2340 (O_2340,N_29816,N_29497);
or UO_2341 (O_2341,N_29577,N_28991);
and UO_2342 (O_2342,N_29173,N_28844);
and UO_2343 (O_2343,N_29655,N_29122);
or UO_2344 (O_2344,N_29960,N_29564);
nor UO_2345 (O_2345,N_28828,N_28886);
xor UO_2346 (O_2346,N_28886,N_29541);
or UO_2347 (O_2347,N_29582,N_29728);
nand UO_2348 (O_2348,N_29398,N_29823);
xnor UO_2349 (O_2349,N_29498,N_29822);
nand UO_2350 (O_2350,N_29586,N_28844);
nand UO_2351 (O_2351,N_29268,N_29310);
nand UO_2352 (O_2352,N_29241,N_29730);
and UO_2353 (O_2353,N_29541,N_29752);
nor UO_2354 (O_2354,N_29298,N_29885);
and UO_2355 (O_2355,N_28989,N_29194);
nor UO_2356 (O_2356,N_29685,N_29662);
and UO_2357 (O_2357,N_29268,N_29421);
nand UO_2358 (O_2358,N_29434,N_29808);
nor UO_2359 (O_2359,N_29273,N_29508);
xnor UO_2360 (O_2360,N_29349,N_29090);
xor UO_2361 (O_2361,N_29029,N_29193);
nand UO_2362 (O_2362,N_28846,N_29176);
nor UO_2363 (O_2363,N_29651,N_29128);
nand UO_2364 (O_2364,N_28973,N_29820);
nor UO_2365 (O_2365,N_29858,N_29775);
nand UO_2366 (O_2366,N_28956,N_29924);
and UO_2367 (O_2367,N_28938,N_29880);
nand UO_2368 (O_2368,N_29239,N_29943);
nand UO_2369 (O_2369,N_29366,N_29015);
xor UO_2370 (O_2370,N_29085,N_29897);
nor UO_2371 (O_2371,N_29257,N_29423);
or UO_2372 (O_2372,N_28888,N_29300);
or UO_2373 (O_2373,N_29355,N_29160);
nand UO_2374 (O_2374,N_29590,N_29855);
nor UO_2375 (O_2375,N_29570,N_29968);
nand UO_2376 (O_2376,N_29303,N_29061);
or UO_2377 (O_2377,N_29957,N_29744);
or UO_2378 (O_2378,N_29967,N_29408);
or UO_2379 (O_2379,N_29019,N_29716);
nand UO_2380 (O_2380,N_29874,N_29186);
nor UO_2381 (O_2381,N_29923,N_28968);
or UO_2382 (O_2382,N_29777,N_29469);
xnor UO_2383 (O_2383,N_28921,N_29413);
nand UO_2384 (O_2384,N_28857,N_28937);
nand UO_2385 (O_2385,N_29131,N_28863);
nor UO_2386 (O_2386,N_29633,N_29610);
nand UO_2387 (O_2387,N_29285,N_29768);
xnor UO_2388 (O_2388,N_29220,N_29955);
or UO_2389 (O_2389,N_29330,N_29539);
nand UO_2390 (O_2390,N_28940,N_29475);
or UO_2391 (O_2391,N_29309,N_29676);
xor UO_2392 (O_2392,N_29905,N_29862);
nor UO_2393 (O_2393,N_29023,N_28814);
or UO_2394 (O_2394,N_29609,N_29284);
xor UO_2395 (O_2395,N_28867,N_29774);
and UO_2396 (O_2396,N_29433,N_29659);
nand UO_2397 (O_2397,N_29431,N_28864);
xor UO_2398 (O_2398,N_29370,N_29077);
or UO_2399 (O_2399,N_29612,N_29698);
nand UO_2400 (O_2400,N_29426,N_28915);
or UO_2401 (O_2401,N_29115,N_29948);
and UO_2402 (O_2402,N_29668,N_29051);
xor UO_2403 (O_2403,N_29820,N_29432);
xnor UO_2404 (O_2404,N_29215,N_29387);
nand UO_2405 (O_2405,N_29438,N_29557);
nor UO_2406 (O_2406,N_29685,N_29364);
and UO_2407 (O_2407,N_29152,N_29490);
xor UO_2408 (O_2408,N_29281,N_28885);
xnor UO_2409 (O_2409,N_28808,N_29251);
nand UO_2410 (O_2410,N_29176,N_29136);
nor UO_2411 (O_2411,N_29421,N_29897);
and UO_2412 (O_2412,N_29863,N_29270);
nand UO_2413 (O_2413,N_29433,N_29024);
xnor UO_2414 (O_2414,N_29595,N_28899);
nand UO_2415 (O_2415,N_29293,N_29143);
and UO_2416 (O_2416,N_29634,N_29620);
and UO_2417 (O_2417,N_29869,N_29095);
and UO_2418 (O_2418,N_29339,N_28940);
nand UO_2419 (O_2419,N_29165,N_29259);
and UO_2420 (O_2420,N_28912,N_29935);
xor UO_2421 (O_2421,N_29315,N_29563);
and UO_2422 (O_2422,N_29836,N_28846);
or UO_2423 (O_2423,N_29464,N_29491);
nor UO_2424 (O_2424,N_29525,N_28819);
and UO_2425 (O_2425,N_29114,N_29744);
nand UO_2426 (O_2426,N_28844,N_29115);
nand UO_2427 (O_2427,N_28947,N_29411);
nor UO_2428 (O_2428,N_29947,N_28803);
nor UO_2429 (O_2429,N_29134,N_29138);
xor UO_2430 (O_2430,N_28916,N_28854);
nor UO_2431 (O_2431,N_29037,N_29366);
nand UO_2432 (O_2432,N_29146,N_28818);
and UO_2433 (O_2433,N_29970,N_29457);
and UO_2434 (O_2434,N_28846,N_29388);
or UO_2435 (O_2435,N_29420,N_29596);
or UO_2436 (O_2436,N_29821,N_29545);
nor UO_2437 (O_2437,N_29523,N_29824);
nor UO_2438 (O_2438,N_29428,N_29918);
xor UO_2439 (O_2439,N_29710,N_28921);
or UO_2440 (O_2440,N_29217,N_29586);
and UO_2441 (O_2441,N_29319,N_29352);
xnor UO_2442 (O_2442,N_29249,N_29473);
or UO_2443 (O_2443,N_29434,N_29239);
nand UO_2444 (O_2444,N_29024,N_28944);
and UO_2445 (O_2445,N_28828,N_29739);
nand UO_2446 (O_2446,N_29696,N_29419);
nand UO_2447 (O_2447,N_29970,N_29325);
nand UO_2448 (O_2448,N_29383,N_29771);
xnor UO_2449 (O_2449,N_29882,N_29314);
and UO_2450 (O_2450,N_29244,N_28996);
nor UO_2451 (O_2451,N_29769,N_28862);
nor UO_2452 (O_2452,N_29030,N_29306);
nand UO_2453 (O_2453,N_29590,N_29625);
and UO_2454 (O_2454,N_28925,N_28939);
and UO_2455 (O_2455,N_29020,N_29440);
and UO_2456 (O_2456,N_29832,N_29900);
nor UO_2457 (O_2457,N_28838,N_29456);
nor UO_2458 (O_2458,N_28805,N_29130);
xnor UO_2459 (O_2459,N_29997,N_29437);
and UO_2460 (O_2460,N_28946,N_29080);
nand UO_2461 (O_2461,N_28923,N_29852);
nand UO_2462 (O_2462,N_29939,N_29227);
nor UO_2463 (O_2463,N_29662,N_29948);
or UO_2464 (O_2464,N_29444,N_29434);
and UO_2465 (O_2465,N_28886,N_29987);
nor UO_2466 (O_2466,N_29264,N_29810);
or UO_2467 (O_2467,N_29053,N_29105);
xor UO_2468 (O_2468,N_29342,N_29121);
or UO_2469 (O_2469,N_29848,N_29934);
or UO_2470 (O_2470,N_29147,N_28838);
and UO_2471 (O_2471,N_29232,N_28945);
or UO_2472 (O_2472,N_29768,N_29132);
nand UO_2473 (O_2473,N_29645,N_29827);
nor UO_2474 (O_2474,N_29493,N_29085);
nand UO_2475 (O_2475,N_29264,N_29200);
xor UO_2476 (O_2476,N_28894,N_29914);
or UO_2477 (O_2477,N_29251,N_29688);
nand UO_2478 (O_2478,N_28887,N_29128);
nor UO_2479 (O_2479,N_29509,N_28969);
xor UO_2480 (O_2480,N_29514,N_29799);
and UO_2481 (O_2481,N_29103,N_29586);
or UO_2482 (O_2482,N_28967,N_29557);
or UO_2483 (O_2483,N_29966,N_29322);
and UO_2484 (O_2484,N_29850,N_29775);
nand UO_2485 (O_2485,N_29030,N_29697);
nand UO_2486 (O_2486,N_29560,N_29617);
or UO_2487 (O_2487,N_29987,N_29039);
nand UO_2488 (O_2488,N_29651,N_29755);
nor UO_2489 (O_2489,N_29382,N_29524);
nor UO_2490 (O_2490,N_29214,N_29756);
xnor UO_2491 (O_2491,N_29639,N_29848);
nand UO_2492 (O_2492,N_28905,N_29086);
xor UO_2493 (O_2493,N_29508,N_29905);
nor UO_2494 (O_2494,N_29423,N_28858);
xor UO_2495 (O_2495,N_29130,N_29246);
or UO_2496 (O_2496,N_29848,N_28952);
nand UO_2497 (O_2497,N_29678,N_29166);
or UO_2498 (O_2498,N_29055,N_29495);
nand UO_2499 (O_2499,N_29184,N_29775);
nor UO_2500 (O_2500,N_29206,N_29675);
nor UO_2501 (O_2501,N_28964,N_29971);
xor UO_2502 (O_2502,N_29965,N_29534);
or UO_2503 (O_2503,N_29941,N_29741);
xnor UO_2504 (O_2504,N_29970,N_29478);
or UO_2505 (O_2505,N_29466,N_28825);
or UO_2506 (O_2506,N_29957,N_29567);
nor UO_2507 (O_2507,N_29680,N_29004);
and UO_2508 (O_2508,N_29139,N_29001);
nand UO_2509 (O_2509,N_29119,N_29169);
or UO_2510 (O_2510,N_28963,N_29702);
xnor UO_2511 (O_2511,N_29103,N_29573);
xor UO_2512 (O_2512,N_29382,N_28963);
xnor UO_2513 (O_2513,N_29183,N_29700);
xnor UO_2514 (O_2514,N_29509,N_29246);
nor UO_2515 (O_2515,N_29054,N_29999);
nor UO_2516 (O_2516,N_29464,N_29447);
nor UO_2517 (O_2517,N_29534,N_29039);
xnor UO_2518 (O_2518,N_29029,N_29280);
xnor UO_2519 (O_2519,N_29627,N_29662);
nand UO_2520 (O_2520,N_29912,N_29893);
and UO_2521 (O_2521,N_28950,N_29982);
xor UO_2522 (O_2522,N_29974,N_28982);
nand UO_2523 (O_2523,N_29794,N_29387);
xnor UO_2524 (O_2524,N_29856,N_29555);
and UO_2525 (O_2525,N_29621,N_29323);
or UO_2526 (O_2526,N_28856,N_29650);
xor UO_2527 (O_2527,N_29197,N_29214);
or UO_2528 (O_2528,N_29451,N_29334);
nor UO_2529 (O_2529,N_29314,N_28934);
nor UO_2530 (O_2530,N_29564,N_29162);
and UO_2531 (O_2531,N_29814,N_29892);
and UO_2532 (O_2532,N_29169,N_29719);
nand UO_2533 (O_2533,N_29802,N_29705);
and UO_2534 (O_2534,N_28885,N_29494);
or UO_2535 (O_2535,N_28908,N_29213);
nor UO_2536 (O_2536,N_29269,N_29593);
or UO_2537 (O_2537,N_29348,N_29662);
or UO_2538 (O_2538,N_29668,N_29703);
xor UO_2539 (O_2539,N_29129,N_29698);
nor UO_2540 (O_2540,N_29874,N_29568);
nand UO_2541 (O_2541,N_29940,N_29052);
xor UO_2542 (O_2542,N_29899,N_29090);
nor UO_2543 (O_2543,N_29619,N_29993);
and UO_2544 (O_2544,N_29270,N_29158);
nor UO_2545 (O_2545,N_29061,N_29109);
xnor UO_2546 (O_2546,N_29476,N_29595);
or UO_2547 (O_2547,N_29764,N_29596);
xnor UO_2548 (O_2548,N_29480,N_28972);
and UO_2549 (O_2549,N_29089,N_29847);
nor UO_2550 (O_2550,N_28879,N_29761);
or UO_2551 (O_2551,N_29839,N_29053);
xor UO_2552 (O_2552,N_29210,N_29047);
or UO_2553 (O_2553,N_29902,N_29525);
or UO_2554 (O_2554,N_29737,N_28851);
nand UO_2555 (O_2555,N_29407,N_29728);
xnor UO_2556 (O_2556,N_29638,N_28819);
and UO_2557 (O_2557,N_28817,N_29200);
nor UO_2558 (O_2558,N_29203,N_28929);
and UO_2559 (O_2559,N_29555,N_29906);
and UO_2560 (O_2560,N_29092,N_29209);
and UO_2561 (O_2561,N_28988,N_29726);
xnor UO_2562 (O_2562,N_28824,N_28842);
nor UO_2563 (O_2563,N_29008,N_29912);
or UO_2564 (O_2564,N_28858,N_29160);
xor UO_2565 (O_2565,N_29537,N_29452);
nor UO_2566 (O_2566,N_29315,N_28852);
xor UO_2567 (O_2567,N_29235,N_29113);
and UO_2568 (O_2568,N_29704,N_28853);
xor UO_2569 (O_2569,N_29871,N_29753);
and UO_2570 (O_2570,N_29753,N_29793);
and UO_2571 (O_2571,N_28997,N_29913);
nand UO_2572 (O_2572,N_29517,N_29438);
or UO_2573 (O_2573,N_29843,N_29810);
xnor UO_2574 (O_2574,N_29681,N_29504);
nand UO_2575 (O_2575,N_29789,N_29754);
nor UO_2576 (O_2576,N_29510,N_29735);
and UO_2577 (O_2577,N_29272,N_29909);
and UO_2578 (O_2578,N_28889,N_29975);
nand UO_2579 (O_2579,N_29068,N_29267);
nor UO_2580 (O_2580,N_29682,N_28839);
xnor UO_2581 (O_2581,N_29195,N_29327);
xnor UO_2582 (O_2582,N_28838,N_28998);
nand UO_2583 (O_2583,N_29437,N_28932);
or UO_2584 (O_2584,N_29545,N_28895);
nor UO_2585 (O_2585,N_29734,N_29180);
nand UO_2586 (O_2586,N_29741,N_29512);
nor UO_2587 (O_2587,N_29852,N_29672);
nand UO_2588 (O_2588,N_29337,N_28940);
nor UO_2589 (O_2589,N_29133,N_29651);
and UO_2590 (O_2590,N_29152,N_28828);
and UO_2591 (O_2591,N_29263,N_29771);
xnor UO_2592 (O_2592,N_29253,N_29310);
nand UO_2593 (O_2593,N_29294,N_29641);
and UO_2594 (O_2594,N_29354,N_29330);
or UO_2595 (O_2595,N_29884,N_28822);
nand UO_2596 (O_2596,N_28971,N_29506);
nand UO_2597 (O_2597,N_29680,N_29628);
xor UO_2598 (O_2598,N_29549,N_29588);
xor UO_2599 (O_2599,N_29985,N_29944);
and UO_2600 (O_2600,N_29868,N_28822);
or UO_2601 (O_2601,N_29696,N_29555);
xnor UO_2602 (O_2602,N_29217,N_28989);
or UO_2603 (O_2603,N_28986,N_29638);
xnor UO_2604 (O_2604,N_28924,N_29644);
or UO_2605 (O_2605,N_29247,N_29864);
and UO_2606 (O_2606,N_29375,N_29403);
or UO_2607 (O_2607,N_29537,N_29798);
nand UO_2608 (O_2608,N_29623,N_29816);
or UO_2609 (O_2609,N_29637,N_28820);
nand UO_2610 (O_2610,N_29872,N_28897);
xnor UO_2611 (O_2611,N_29359,N_28870);
and UO_2612 (O_2612,N_29434,N_29586);
or UO_2613 (O_2613,N_29078,N_29327);
nand UO_2614 (O_2614,N_29825,N_29256);
nand UO_2615 (O_2615,N_29920,N_29997);
nand UO_2616 (O_2616,N_29508,N_29860);
nand UO_2617 (O_2617,N_29111,N_29966);
xor UO_2618 (O_2618,N_29423,N_29565);
and UO_2619 (O_2619,N_28836,N_29225);
xor UO_2620 (O_2620,N_28838,N_29468);
nor UO_2621 (O_2621,N_29041,N_29408);
nor UO_2622 (O_2622,N_29886,N_29950);
nand UO_2623 (O_2623,N_29396,N_29881);
and UO_2624 (O_2624,N_29071,N_29054);
or UO_2625 (O_2625,N_28914,N_29418);
xor UO_2626 (O_2626,N_28808,N_29952);
nand UO_2627 (O_2627,N_29500,N_29049);
nor UO_2628 (O_2628,N_28962,N_29593);
nor UO_2629 (O_2629,N_28897,N_29967);
xnor UO_2630 (O_2630,N_28926,N_29673);
nor UO_2631 (O_2631,N_29273,N_28801);
and UO_2632 (O_2632,N_28998,N_29253);
xor UO_2633 (O_2633,N_29819,N_28935);
and UO_2634 (O_2634,N_29296,N_29359);
nor UO_2635 (O_2635,N_29057,N_29518);
xor UO_2636 (O_2636,N_29414,N_29999);
and UO_2637 (O_2637,N_29613,N_29330);
and UO_2638 (O_2638,N_29715,N_29381);
nor UO_2639 (O_2639,N_29100,N_28825);
nor UO_2640 (O_2640,N_29987,N_28964);
nand UO_2641 (O_2641,N_29773,N_29269);
nand UO_2642 (O_2642,N_29521,N_29345);
nand UO_2643 (O_2643,N_29841,N_29239);
or UO_2644 (O_2644,N_29339,N_29612);
nand UO_2645 (O_2645,N_29765,N_29473);
and UO_2646 (O_2646,N_28850,N_29407);
xor UO_2647 (O_2647,N_29957,N_28958);
nor UO_2648 (O_2648,N_29639,N_29672);
and UO_2649 (O_2649,N_29317,N_29380);
nor UO_2650 (O_2650,N_29387,N_29166);
nor UO_2651 (O_2651,N_29645,N_29455);
nor UO_2652 (O_2652,N_29302,N_29416);
nand UO_2653 (O_2653,N_29280,N_29669);
and UO_2654 (O_2654,N_29306,N_29815);
nor UO_2655 (O_2655,N_29140,N_29539);
or UO_2656 (O_2656,N_29629,N_29236);
or UO_2657 (O_2657,N_29714,N_29178);
and UO_2658 (O_2658,N_29316,N_29549);
or UO_2659 (O_2659,N_29678,N_28811);
nand UO_2660 (O_2660,N_28902,N_28919);
and UO_2661 (O_2661,N_29158,N_29650);
xnor UO_2662 (O_2662,N_29381,N_29552);
xor UO_2663 (O_2663,N_28878,N_28813);
or UO_2664 (O_2664,N_29674,N_29146);
nand UO_2665 (O_2665,N_29493,N_29389);
nor UO_2666 (O_2666,N_29407,N_29361);
nor UO_2667 (O_2667,N_28911,N_29503);
or UO_2668 (O_2668,N_29578,N_29625);
xor UO_2669 (O_2669,N_29251,N_29500);
or UO_2670 (O_2670,N_28801,N_29854);
nand UO_2671 (O_2671,N_29612,N_29354);
and UO_2672 (O_2672,N_29969,N_29359);
xor UO_2673 (O_2673,N_29746,N_29206);
and UO_2674 (O_2674,N_29901,N_29671);
xor UO_2675 (O_2675,N_29109,N_28842);
and UO_2676 (O_2676,N_29679,N_29316);
xor UO_2677 (O_2677,N_28922,N_29715);
or UO_2678 (O_2678,N_29491,N_29978);
xnor UO_2679 (O_2679,N_28961,N_29671);
nor UO_2680 (O_2680,N_28968,N_29952);
nand UO_2681 (O_2681,N_29495,N_29156);
nor UO_2682 (O_2682,N_29307,N_29296);
or UO_2683 (O_2683,N_29478,N_29468);
or UO_2684 (O_2684,N_29372,N_29508);
xor UO_2685 (O_2685,N_29419,N_29425);
and UO_2686 (O_2686,N_29148,N_29594);
or UO_2687 (O_2687,N_29641,N_29894);
and UO_2688 (O_2688,N_29016,N_29770);
nor UO_2689 (O_2689,N_28983,N_29985);
xnor UO_2690 (O_2690,N_29626,N_29412);
or UO_2691 (O_2691,N_29847,N_29863);
xnor UO_2692 (O_2692,N_29577,N_29075);
and UO_2693 (O_2693,N_29029,N_29442);
nand UO_2694 (O_2694,N_29723,N_29386);
and UO_2695 (O_2695,N_29050,N_29171);
xor UO_2696 (O_2696,N_29581,N_29667);
xor UO_2697 (O_2697,N_29705,N_29982);
nor UO_2698 (O_2698,N_29316,N_29006);
or UO_2699 (O_2699,N_29435,N_29224);
xor UO_2700 (O_2700,N_29069,N_29266);
or UO_2701 (O_2701,N_29471,N_28830);
nor UO_2702 (O_2702,N_29964,N_28926);
xnor UO_2703 (O_2703,N_29642,N_29741);
nor UO_2704 (O_2704,N_28880,N_29161);
nand UO_2705 (O_2705,N_29989,N_29838);
nor UO_2706 (O_2706,N_29962,N_28868);
or UO_2707 (O_2707,N_29582,N_29263);
xnor UO_2708 (O_2708,N_28942,N_28844);
or UO_2709 (O_2709,N_29736,N_28835);
and UO_2710 (O_2710,N_29907,N_29320);
and UO_2711 (O_2711,N_29089,N_29676);
xnor UO_2712 (O_2712,N_29844,N_29296);
xor UO_2713 (O_2713,N_29193,N_29686);
and UO_2714 (O_2714,N_29012,N_29007);
and UO_2715 (O_2715,N_29312,N_29448);
nand UO_2716 (O_2716,N_29949,N_29144);
nand UO_2717 (O_2717,N_28877,N_29118);
xor UO_2718 (O_2718,N_29007,N_28874);
and UO_2719 (O_2719,N_29088,N_29094);
xor UO_2720 (O_2720,N_28887,N_29286);
nand UO_2721 (O_2721,N_29425,N_28822);
or UO_2722 (O_2722,N_29492,N_28846);
nand UO_2723 (O_2723,N_29606,N_29566);
nor UO_2724 (O_2724,N_29856,N_28816);
xnor UO_2725 (O_2725,N_29853,N_29767);
xor UO_2726 (O_2726,N_29699,N_29134);
xnor UO_2727 (O_2727,N_29524,N_29572);
nor UO_2728 (O_2728,N_29861,N_29962);
xor UO_2729 (O_2729,N_28893,N_29283);
nor UO_2730 (O_2730,N_29884,N_29510);
nor UO_2731 (O_2731,N_29237,N_28811);
nand UO_2732 (O_2732,N_29567,N_29710);
nand UO_2733 (O_2733,N_29185,N_29785);
nor UO_2734 (O_2734,N_29906,N_29261);
or UO_2735 (O_2735,N_29480,N_29591);
and UO_2736 (O_2736,N_29208,N_29937);
and UO_2737 (O_2737,N_29378,N_29538);
xnor UO_2738 (O_2738,N_28869,N_29655);
xor UO_2739 (O_2739,N_28868,N_28804);
or UO_2740 (O_2740,N_29536,N_29085);
nor UO_2741 (O_2741,N_29137,N_29948);
or UO_2742 (O_2742,N_29700,N_29581);
nand UO_2743 (O_2743,N_29742,N_29530);
nor UO_2744 (O_2744,N_29202,N_29741);
nand UO_2745 (O_2745,N_29160,N_29741);
or UO_2746 (O_2746,N_29855,N_29948);
xnor UO_2747 (O_2747,N_29692,N_29353);
or UO_2748 (O_2748,N_29973,N_29493);
and UO_2749 (O_2749,N_29748,N_28959);
nor UO_2750 (O_2750,N_29106,N_29802);
nor UO_2751 (O_2751,N_29032,N_29690);
nor UO_2752 (O_2752,N_29232,N_29552);
nor UO_2753 (O_2753,N_29570,N_29490);
or UO_2754 (O_2754,N_29395,N_29186);
and UO_2755 (O_2755,N_29415,N_28995);
nand UO_2756 (O_2756,N_28922,N_29535);
or UO_2757 (O_2757,N_29488,N_29131);
and UO_2758 (O_2758,N_29724,N_28965);
nor UO_2759 (O_2759,N_29811,N_29507);
and UO_2760 (O_2760,N_29767,N_29479);
and UO_2761 (O_2761,N_29129,N_29122);
nor UO_2762 (O_2762,N_29236,N_29374);
xnor UO_2763 (O_2763,N_28867,N_29542);
or UO_2764 (O_2764,N_29782,N_29351);
nor UO_2765 (O_2765,N_29428,N_28847);
nor UO_2766 (O_2766,N_29120,N_29607);
nand UO_2767 (O_2767,N_29779,N_29051);
xnor UO_2768 (O_2768,N_29775,N_29438);
xnor UO_2769 (O_2769,N_28934,N_29882);
or UO_2770 (O_2770,N_29681,N_29382);
nand UO_2771 (O_2771,N_28824,N_28833);
nand UO_2772 (O_2772,N_29123,N_29040);
or UO_2773 (O_2773,N_28824,N_29898);
nor UO_2774 (O_2774,N_29469,N_29318);
and UO_2775 (O_2775,N_28991,N_29233);
nor UO_2776 (O_2776,N_28919,N_29568);
xor UO_2777 (O_2777,N_29338,N_29066);
nand UO_2778 (O_2778,N_28945,N_29910);
nand UO_2779 (O_2779,N_29057,N_29916);
and UO_2780 (O_2780,N_29884,N_28859);
or UO_2781 (O_2781,N_29619,N_29800);
nand UO_2782 (O_2782,N_29406,N_28931);
and UO_2783 (O_2783,N_28862,N_29827);
xor UO_2784 (O_2784,N_29739,N_29562);
xor UO_2785 (O_2785,N_29188,N_29528);
xnor UO_2786 (O_2786,N_29889,N_28845);
and UO_2787 (O_2787,N_28979,N_28861);
xnor UO_2788 (O_2788,N_29563,N_29277);
xnor UO_2789 (O_2789,N_29013,N_29010);
xnor UO_2790 (O_2790,N_29621,N_29266);
or UO_2791 (O_2791,N_29364,N_29854);
or UO_2792 (O_2792,N_28837,N_29341);
nor UO_2793 (O_2793,N_29570,N_29955);
xor UO_2794 (O_2794,N_28809,N_29565);
and UO_2795 (O_2795,N_28944,N_28929);
nand UO_2796 (O_2796,N_29591,N_29148);
nand UO_2797 (O_2797,N_29008,N_29016);
nand UO_2798 (O_2798,N_28909,N_29919);
nor UO_2799 (O_2799,N_28984,N_29639);
nor UO_2800 (O_2800,N_29906,N_29448);
xor UO_2801 (O_2801,N_28966,N_29188);
nand UO_2802 (O_2802,N_29369,N_29417);
nor UO_2803 (O_2803,N_29424,N_29388);
or UO_2804 (O_2804,N_29414,N_29493);
xnor UO_2805 (O_2805,N_28917,N_29335);
and UO_2806 (O_2806,N_29144,N_28951);
and UO_2807 (O_2807,N_29739,N_29652);
and UO_2808 (O_2808,N_29682,N_29274);
and UO_2809 (O_2809,N_29041,N_29972);
and UO_2810 (O_2810,N_29453,N_29066);
and UO_2811 (O_2811,N_29042,N_29616);
nor UO_2812 (O_2812,N_29964,N_28868);
and UO_2813 (O_2813,N_29147,N_29685);
nor UO_2814 (O_2814,N_29277,N_29483);
nor UO_2815 (O_2815,N_29404,N_29119);
xnor UO_2816 (O_2816,N_29360,N_29984);
nor UO_2817 (O_2817,N_29008,N_29964);
and UO_2818 (O_2818,N_29217,N_29115);
or UO_2819 (O_2819,N_29568,N_29938);
xor UO_2820 (O_2820,N_29250,N_29111);
nand UO_2821 (O_2821,N_29647,N_29408);
nand UO_2822 (O_2822,N_29393,N_29713);
nand UO_2823 (O_2823,N_29922,N_29220);
or UO_2824 (O_2824,N_29895,N_28900);
and UO_2825 (O_2825,N_29472,N_28859);
xor UO_2826 (O_2826,N_29705,N_29787);
xor UO_2827 (O_2827,N_29310,N_28818);
or UO_2828 (O_2828,N_29865,N_29525);
xnor UO_2829 (O_2829,N_29572,N_29614);
nand UO_2830 (O_2830,N_29370,N_29036);
xnor UO_2831 (O_2831,N_29070,N_29611);
xnor UO_2832 (O_2832,N_29120,N_29326);
and UO_2833 (O_2833,N_28964,N_29139);
and UO_2834 (O_2834,N_29790,N_28844);
and UO_2835 (O_2835,N_29286,N_28815);
or UO_2836 (O_2836,N_29766,N_29750);
nor UO_2837 (O_2837,N_29157,N_29810);
and UO_2838 (O_2838,N_29621,N_28885);
and UO_2839 (O_2839,N_29847,N_28818);
or UO_2840 (O_2840,N_29580,N_28943);
nor UO_2841 (O_2841,N_29351,N_28840);
nand UO_2842 (O_2842,N_29891,N_28899);
xnor UO_2843 (O_2843,N_28801,N_29632);
nor UO_2844 (O_2844,N_29626,N_29613);
xnor UO_2845 (O_2845,N_29974,N_29428);
nand UO_2846 (O_2846,N_29271,N_29637);
xnor UO_2847 (O_2847,N_28944,N_29641);
or UO_2848 (O_2848,N_29562,N_29473);
nor UO_2849 (O_2849,N_28910,N_29480);
nand UO_2850 (O_2850,N_29218,N_28958);
or UO_2851 (O_2851,N_29349,N_29279);
nor UO_2852 (O_2852,N_29787,N_28884);
xnor UO_2853 (O_2853,N_29002,N_28807);
and UO_2854 (O_2854,N_29575,N_29877);
xnor UO_2855 (O_2855,N_29614,N_29463);
nor UO_2856 (O_2856,N_28944,N_29519);
nor UO_2857 (O_2857,N_29860,N_28901);
nor UO_2858 (O_2858,N_29646,N_29988);
xor UO_2859 (O_2859,N_29350,N_28907);
nand UO_2860 (O_2860,N_29221,N_29738);
nor UO_2861 (O_2861,N_29729,N_29208);
or UO_2862 (O_2862,N_28966,N_29560);
nor UO_2863 (O_2863,N_29074,N_29662);
and UO_2864 (O_2864,N_29051,N_29614);
nand UO_2865 (O_2865,N_28815,N_29771);
nand UO_2866 (O_2866,N_29628,N_28824);
or UO_2867 (O_2867,N_29501,N_28896);
or UO_2868 (O_2868,N_29984,N_28827);
and UO_2869 (O_2869,N_29516,N_29442);
nand UO_2870 (O_2870,N_28881,N_29503);
and UO_2871 (O_2871,N_29485,N_29194);
nor UO_2872 (O_2872,N_28919,N_29751);
xor UO_2873 (O_2873,N_28941,N_29949);
nor UO_2874 (O_2874,N_29388,N_29307);
or UO_2875 (O_2875,N_28968,N_29137);
xnor UO_2876 (O_2876,N_29319,N_29375);
or UO_2877 (O_2877,N_29647,N_29243);
nor UO_2878 (O_2878,N_29657,N_29389);
xor UO_2879 (O_2879,N_29847,N_29216);
and UO_2880 (O_2880,N_28863,N_29078);
nor UO_2881 (O_2881,N_29350,N_29067);
and UO_2882 (O_2882,N_29595,N_29726);
nand UO_2883 (O_2883,N_29545,N_29327);
and UO_2884 (O_2884,N_29434,N_29059);
and UO_2885 (O_2885,N_29673,N_29570);
and UO_2886 (O_2886,N_29196,N_29343);
nor UO_2887 (O_2887,N_29327,N_29020);
xnor UO_2888 (O_2888,N_29063,N_29151);
and UO_2889 (O_2889,N_29450,N_29158);
xor UO_2890 (O_2890,N_29162,N_29716);
xor UO_2891 (O_2891,N_29750,N_29384);
nor UO_2892 (O_2892,N_28891,N_28800);
nor UO_2893 (O_2893,N_29667,N_28917);
nor UO_2894 (O_2894,N_29462,N_29275);
nand UO_2895 (O_2895,N_29581,N_29262);
xor UO_2896 (O_2896,N_28838,N_29803);
nor UO_2897 (O_2897,N_29709,N_29125);
or UO_2898 (O_2898,N_28914,N_29817);
xor UO_2899 (O_2899,N_29661,N_28894);
or UO_2900 (O_2900,N_29809,N_29508);
nand UO_2901 (O_2901,N_29559,N_29037);
xnor UO_2902 (O_2902,N_29140,N_29211);
xnor UO_2903 (O_2903,N_29038,N_29190);
xnor UO_2904 (O_2904,N_29270,N_29585);
and UO_2905 (O_2905,N_29275,N_29506);
and UO_2906 (O_2906,N_29129,N_29063);
and UO_2907 (O_2907,N_29705,N_29143);
or UO_2908 (O_2908,N_29872,N_29694);
xnor UO_2909 (O_2909,N_29032,N_29528);
nor UO_2910 (O_2910,N_29374,N_29114);
and UO_2911 (O_2911,N_29106,N_28948);
nand UO_2912 (O_2912,N_28975,N_29043);
nor UO_2913 (O_2913,N_29898,N_29609);
and UO_2914 (O_2914,N_29453,N_29747);
xor UO_2915 (O_2915,N_28942,N_29929);
or UO_2916 (O_2916,N_29898,N_29352);
or UO_2917 (O_2917,N_29370,N_29037);
nand UO_2918 (O_2918,N_29126,N_29605);
nor UO_2919 (O_2919,N_29269,N_29203);
xnor UO_2920 (O_2920,N_29654,N_29939);
or UO_2921 (O_2921,N_28990,N_29607);
xnor UO_2922 (O_2922,N_29261,N_29707);
and UO_2923 (O_2923,N_29582,N_29380);
nor UO_2924 (O_2924,N_28827,N_29691);
or UO_2925 (O_2925,N_29560,N_29326);
or UO_2926 (O_2926,N_29921,N_28966);
nor UO_2927 (O_2927,N_29508,N_29620);
nor UO_2928 (O_2928,N_29678,N_29766);
or UO_2929 (O_2929,N_29709,N_29622);
nor UO_2930 (O_2930,N_29804,N_29655);
xnor UO_2931 (O_2931,N_29715,N_29108);
nand UO_2932 (O_2932,N_29010,N_29094);
xor UO_2933 (O_2933,N_29578,N_29326);
or UO_2934 (O_2934,N_29485,N_28996);
and UO_2935 (O_2935,N_29411,N_29666);
and UO_2936 (O_2936,N_29644,N_29279);
or UO_2937 (O_2937,N_29097,N_29561);
or UO_2938 (O_2938,N_29132,N_29112);
nand UO_2939 (O_2939,N_28896,N_29751);
and UO_2940 (O_2940,N_29862,N_29473);
and UO_2941 (O_2941,N_29295,N_29841);
or UO_2942 (O_2942,N_29690,N_29843);
nor UO_2943 (O_2943,N_29854,N_29120);
or UO_2944 (O_2944,N_29781,N_29166);
nor UO_2945 (O_2945,N_29666,N_29953);
nand UO_2946 (O_2946,N_28972,N_29093);
nand UO_2947 (O_2947,N_29776,N_28992);
and UO_2948 (O_2948,N_29936,N_29828);
nor UO_2949 (O_2949,N_28918,N_29691);
xnor UO_2950 (O_2950,N_29523,N_29567);
nor UO_2951 (O_2951,N_29842,N_29352);
nor UO_2952 (O_2952,N_28975,N_29123);
and UO_2953 (O_2953,N_29027,N_29967);
nor UO_2954 (O_2954,N_29248,N_28885);
and UO_2955 (O_2955,N_28929,N_29726);
or UO_2956 (O_2956,N_28890,N_29922);
and UO_2957 (O_2957,N_28942,N_29861);
xnor UO_2958 (O_2958,N_28920,N_28843);
nand UO_2959 (O_2959,N_29424,N_28870);
or UO_2960 (O_2960,N_29182,N_29635);
or UO_2961 (O_2961,N_29520,N_29936);
xnor UO_2962 (O_2962,N_29296,N_29276);
and UO_2963 (O_2963,N_29394,N_29562);
nand UO_2964 (O_2964,N_29150,N_29882);
nor UO_2965 (O_2965,N_29312,N_29761);
or UO_2966 (O_2966,N_29654,N_29375);
nand UO_2967 (O_2967,N_29706,N_28879);
xnor UO_2968 (O_2968,N_29763,N_28961);
and UO_2969 (O_2969,N_29483,N_29105);
nor UO_2970 (O_2970,N_29189,N_29768);
or UO_2971 (O_2971,N_29538,N_29852);
xor UO_2972 (O_2972,N_29285,N_29229);
nor UO_2973 (O_2973,N_28875,N_28825);
xor UO_2974 (O_2974,N_29456,N_29588);
and UO_2975 (O_2975,N_29719,N_29903);
or UO_2976 (O_2976,N_29334,N_29176);
and UO_2977 (O_2977,N_29668,N_29221);
nor UO_2978 (O_2978,N_29879,N_29636);
or UO_2979 (O_2979,N_29923,N_29437);
xor UO_2980 (O_2980,N_29980,N_29543);
xnor UO_2981 (O_2981,N_29807,N_29713);
xnor UO_2982 (O_2982,N_29389,N_29739);
or UO_2983 (O_2983,N_29466,N_29322);
and UO_2984 (O_2984,N_28912,N_29953);
or UO_2985 (O_2985,N_29975,N_29012);
nor UO_2986 (O_2986,N_29970,N_29829);
xor UO_2987 (O_2987,N_29608,N_29733);
nand UO_2988 (O_2988,N_29498,N_28916);
xor UO_2989 (O_2989,N_29491,N_29133);
nor UO_2990 (O_2990,N_29155,N_29891);
and UO_2991 (O_2991,N_29447,N_29756);
and UO_2992 (O_2992,N_29493,N_29087);
or UO_2993 (O_2993,N_29130,N_29580);
nand UO_2994 (O_2994,N_28975,N_29064);
nor UO_2995 (O_2995,N_29441,N_29350);
or UO_2996 (O_2996,N_29435,N_28918);
nor UO_2997 (O_2997,N_29740,N_28919);
and UO_2998 (O_2998,N_29484,N_28902);
nand UO_2999 (O_2999,N_29484,N_29006);
xnor UO_3000 (O_3000,N_29787,N_29531);
nor UO_3001 (O_3001,N_29783,N_29629);
or UO_3002 (O_3002,N_29723,N_28830);
nor UO_3003 (O_3003,N_29265,N_29221);
and UO_3004 (O_3004,N_29657,N_29471);
or UO_3005 (O_3005,N_29720,N_29175);
or UO_3006 (O_3006,N_29117,N_29988);
xnor UO_3007 (O_3007,N_29150,N_28819);
nor UO_3008 (O_3008,N_29724,N_29003);
and UO_3009 (O_3009,N_29488,N_29948);
or UO_3010 (O_3010,N_28849,N_28946);
and UO_3011 (O_3011,N_28846,N_28816);
nand UO_3012 (O_3012,N_29722,N_28882);
and UO_3013 (O_3013,N_29905,N_29414);
and UO_3014 (O_3014,N_29005,N_29458);
nor UO_3015 (O_3015,N_29220,N_29562);
nor UO_3016 (O_3016,N_28819,N_28963);
xnor UO_3017 (O_3017,N_29476,N_29014);
xor UO_3018 (O_3018,N_29532,N_29452);
or UO_3019 (O_3019,N_28841,N_29110);
and UO_3020 (O_3020,N_29421,N_29942);
nor UO_3021 (O_3021,N_29406,N_28869);
and UO_3022 (O_3022,N_28994,N_29890);
or UO_3023 (O_3023,N_29675,N_29128);
and UO_3024 (O_3024,N_29187,N_29392);
nor UO_3025 (O_3025,N_28806,N_29262);
or UO_3026 (O_3026,N_28961,N_29363);
xnor UO_3027 (O_3027,N_29483,N_29916);
nor UO_3028 (O_3028,N_29138,N_29560);
nand UO_3029 (O_3029,N_29339,N_29535);
xor UO_3030 (O_3030,N_29790,N_29742);
or UO_3031 (O_3031,N_29342,N_29463);
and UO_3032 (O_3032,N_29284,N_29703);
xor UO_3033 (O_3033,N_29031,N_29599);
or UO_3034 (O_3034,N_29045,N_29034);
and UO_3035 (O_3035,N_29650,N_29666);
nand UO_3036 (O_3036,N_28902,N_29791);
xnor UO_3037 (O_3037,N_29007,N_29996);
and UO_3038 (O_3038,N_28813,N_29351);
or UO_3039 (O_3039,N_28939,N_29914);
xor UO_3040 (O_3040,N_29297,N_29535);
or UO_3041 (O_3041,N_29278,N_29660);
or UO_3042 (O_3042,N_29118,N_29628);
xor UO_3043 (O_3043,N_29385,N_29273);
and UO_3044 (O_3044,N_29346,N_28914);
nand UO_3045 (O_3045,N_29284,N_29966);
and UO_3046 (O_3046,N_29646,N_29511);
and UO_3047 (O_3047,N_29260,N_29368);
and UO_3048 (O_3048,N_29053,N_29245);
nor UO_3049 (O_3049,N_28862,N_29165);
nor UO_3050 (O_3050,N_29196,N_29865);
xor UO_3051 (O_3051,N_29751,N_29878);
or UO_3052 (O_3052,N_28970,N_29945);
and UO_3053 (O_3053,N_29511,N_29198);
or UO_3054 (O_3054,N_29552,N_29132);
xnor UO_3055 (O_3055,N_29670,N_29708);
nand UO_3056 (O_3056,N_29353,N_29780);
xnor UO_3057 (O_3057,N_29864,N_29066);
or UO_3058 (O_3058,N_29949,N_29779);
and UO_3059 (O_3059,N_29371,N_29314);
xor UO_3060 (O_3060,N_29562,N_29344);
xnor UO_3061 (O_3061,N_28926,N_29146);
and UO_3062 (O_3062,N_29862,N_29214);
nand UO_3063 (O_3063,N_28903,N_29260);
or UO_3064 (O_3064,N_29528,N_29135);
nand UO_3065 (O_3065,N_29302,N_29677);
and UO_3066 (O_3066,N_28867,N_29011);
and UO_3067 (O_3067,N_29160,N_29726);
xnor UO_3068 (O_3068,N_29210,N_29569);
xnor UO_3069 (O_3069,N_29967,N_29511);
and UO_3070 (O_3070,N_28930,N_29686);
xnor UO_3071 (O_3071,N_29281,N_29186);
nor UO_3072 (O_3072,N_29633,N_28942);
and UO_3073 (O_3073,N_28809,N_29374);
and UO_3074 (O_3074,N_29114,N_29853);
nand UO_3075 (O_3075,N_29899,N_29306);
or UO_3076 (O_3076,N_29443,N_29921);
nor UO_3077 (O_3077,N_28857,N_28898);
xor UO_3078 (O_3078,N_28815,N_29717);
xnor UO_3079 (O_3079,N_29528,N_29138);
nor UO_3080 (O_3080,N_29652,N_29812);
nor UO_3081 (O_3081,N_29192,N_29042);
or UO_3082 (O_3082,N_28952,N_29447);
and UO_3083 (O_3083,N_29206,N_29868);
nor UO_3084 (O_3084,N_29524,N_29314);
nor UO_3085 (O_3085,N_29200,N_29791);
nor UO_3086 (O_3086,N_28886,N_29566);
nand UO_3087 (O_3087,N_28819,N_29107);
nor UO_3088 (O_3088,N_29846,N_29686);
nand UO_3089 (O_3089,N_29397,N_29592);
and UO_3090 (O_3090,N_29176,N_29642);
and UO_3091 (O_3091,N_29641,N_29776);
or UO_3092 (O_3092,N_29522,N_29420);
nand UO_3093 (O_3093,N_29055,N_28888);
nor UO_3094 (O_3094,N_29123,N_29446);
and UO_3095 (O_3095,N_29421,N_29682);
nor UO_3096 (O_3096,N_29214,N_29655);
or UO_3097 (O_3097,N_28826,N_29423);
nor UO_3098 (O_3098,N_29718,N_28822);
nand UO_3099 (O_3099,N_29865,N_29895);
and UO_3100 (O_3100,N_29522,N_29799);
and UO_3101 (O_3101,N_29888,N_29618);
or UO_3102 (O_3102,N_29556,N_29902);
and UO_3103 (O_3103,N_29009,N_29349);
and UO_3104 (O_3104,N_29469,N_29227);
nand UO_3105 (O_3105,N_29139,N_29408);
or UO_3106 (O_3106,N_29184,N_29770);
nor UO_3107 (O_3107,N_29797,N_29964);
or UO_3108 (O_3108,N_29350,N_29490);
and UO_3109 (O_3109,N_29532,N_29553);
nand UO_3110 (O_3110,N_29450,N_28920);
or UO_3111 (O_3111,N_29263,N_29184);
nand UO_3112 (O_3112,N_29747,N_29558);
or UO_3113 (O_3113,N_29551,N_28880);
nor UO_3114 (O_3114,N_28836,N_29825);
xor UO_3115 (O_3115,N_29917,N_29655);
nand UO_3116 (O_3116,N_28911,N_29217);
nand UO_3117 (O_3117,N_29904,N_29602);
xnor UO_3118 (O_3118,N_29308,N_29877);
xor UO_3119 (O_3119,N_28968,N_29318);
and UO_3120 (O_3120,N_29508,N_29412);
or UO_3121 (O_3121,N_29493,N_29373);
and UO_3122 (O_3122,N_29211,N_29440);
nand UO_3123 (O_3123,N_29009,N_29607);
xor UO_3124 (O_3124,N_29797,N_28908);
and UO_3125 (O_3125,N_28823,N_29711);
nand UO_3126 (O_3126,N_29051,N_29277);
nand UO_3127 (O_3127,N_29058,N_29024);
and UO_3128 (O_3128,N_29013,N_29763);
nor UO_3129 (O_3129,N_29027,N_29515);
nor UO_3130 (O_3130,N_28809,N_28867);
nor UO_3131 (O_3131,N_29510,N_28946);
nor UO_3132 (O_3132,N_29627,N_29789);
and UO_3133 (O_3133,N_29836,N_29780);
or UO_3134 (O_3134,N_28863,N_29791);
nor UO_3135 (O_3135,N_28846,N_29046);
nand UO_3136 (O_3136,N_29681,N_29406);
and UO_3137 (O_3137,N_28882,N_29194);
nor UO_3138 (O_3138,N_29864,N_29415);
nand UO_3139 (O_3139,N_29076,N_29640);
and UO_3140 (O_3140,N_29895,N_29430);
nor UO_3141 (O_3141,N_29800,N_29528);
xor UO_3142 (O_3142,N_29454,N_28809);
and UO_3143 (O_3143,N_29397,N_29731);
xnor UO_3144 (O_3144,N_29341,N_29217);
or UO_3145 (O_3145,N_28998,N_29875);
nor UO_3146 (O_3146,N_29192,N_29154);
nor UO_3147 (O_3147,N_29958,N_28966);
or UO_3148 (O_3148,N_29760,N_29387);
nand UO_3149 (O_3149,N_28931,N_29209);
or UO_3150 (O_3150,N_29654,N_29686);
nand UO_3151 (O_3151,N_29081,N_28937);
nor UO_3152 (O_3152,N_29826,N_29227);
nand UO_3153 (O_3153,N_29333,N_29493);
and UO_3154 (O_3154,N_29510,N_29543);
or UO_3155 (O_3155,N_29309,N_29721);
xor UO_3156 (O_3156,N_29612,N_29256);
or UO_3157 (O_3157,N_29058,N_29891);
xor UO_3158 (O_3158,N_29095,N_29778);
and UO_3159 (O_3159,N_28905,N_29658);
nor UO_3160 (O_3160,N_28826,N_29977);
xnor UO_3161 (O_3161,N_29644,N_29692);
nor UO_3162 (O_3162,N_29979,N_29572);
xnor UO_3163 (O_3163,N_29913,N_29878);
or UO_3164 (O_3164,N_29102,N_29614);
and UO_3165 (O_3165,N_29401,N_29679);
nor UO_3166 (O_3166,N_29737,N_29069);
or UO_3167 (O_3167,N_29159,N_29073);
xnor UO_3168 (O_3168,N_28815,N_28911);
or UO_3169 (O_3169,N_29145,N_29221);
nand UO_3170 (O_3170,N_29787,N_29142);
and UO_3171 (O_3171,N_28832,N_29896);
nand UO_3172 (O_3172,N_28944,N_29808);
or UO_3173 (O_3173,N_29540,N_29818);
nor UO_3174 (O_3174,N_29488,N_28838);
xor UO_3175 (O_3175,N_29944,N_29170);
nor UO_3176 (O_3176,N_29294,N_29788);
nand UO_3177 (O_3177,N_29766,N_29427);
or UO_3178 (O_3178,N_29753,N_29279);
xor UO_3179 (O_3179,N_29181,N_29836);
nand UO_3180 (O_3180,N_29880,N_29945);
nand UO_3181 (O_3181,N_29189,N_28983);
nand UO_3182 (O_3182,N_29942,N_29264);
or UO_3183 (O_3183,N_29128,N_29617);
nor UO_3184 (O_3184,N_29541,N_29833);
and UO_3185 (O_3185,N_29280,N_29903);
and UO_3186 (O_3186,N_29653,N_29579);
and UO_3187 (O_3187,N_29201,N_29927);
nor UO_3188 (O_3188,N_28995,N_29033);
or UO_3189 (O_3189,N_29757,N_28839);
xor UO_3190 (O_3190,N_29393,N_29415);
or UO_3191 (O_3191,N_29749,N_29807);
or UO_3192 (O_3192,N_29819,N_29557);
nand UO_3193 (O_3193,N_28944,N_29243);
and UO_3194 (O_3194,N_29178,N_29996);
nand UO_3195 (O_3195,N_28867,N_29141);
and UO_3196 (O_3196,N_29031,N_29783);
xor UO_3197 (O_3197,N_29271,N_29091);
nand UO_3198 (O_3198,N_29248,N_29432);
nor UO_3199 (O_3199,N_28886,N_29506);
or UO_3200 (O_3200,N_29103,N_29512);
and UO_3201 (O_3201,N_29527,N_28942);
xor UO_3202 (O_3202,N_28849,N_28912);
and UO_3203 (O_3203,N_29440,N_29107);
or UO_3204 (O_3204,N_29165,N_29618);
or UO_3205 (O_3205,N_29652,N_28829);
xor UO_3206 (O_3206,N_29186,N_29856);
nor UO_3207 (O_3207,N_29863,N_29695);
nor UO_3208 (O_3208,N_29185,N_29301);
xnor UO_3209 (O_3209,N_29818,N_29250);
xnor UO_3210 (O_3210,N_28848,N_29750);
nor UO_3211 (O_3211,N_29208,N_28885);
xor UO_3212 (O_3212,N_28854,N_29842);
nand UO_3213 (O_3213,N_29404,N_29706);
nand UO_3214 (O_3214,N_29707,N_29429);
or UO_3215 (O_3215,N_29892,N_28816);
xor UO_3216 (O_3216,N_29883,N_29547);
and UO_3217 (O_3217,N_28819,N_29672);
nor UO_3218 (O_3218,N_28871,N_29998);
and UO_3219 (O_3219,N_29779,N_29736);
and UO_3220 (O_3220,N_28909,N_29769);
nor UO_3221 (O_3221,N_28937,N_29278);
and UO_3222 (O_3222,N_29161,N_29608);
nand UO_3223 (O_3223,N_28957,N_29770);
or UO_3224 (O_3224,N_28832,N_29903);
nand UO_3225 (O_3225,N_29833,N_29379);
xnor UO_3226 (O_3226,N_28878,N_29727);
xnor UO_3227 (O_3227,N_29596,N_29849);
xor UO_3228 (O_3228,N_29649,N_29248);
and UO_3229 (O_3229,N_29739,N_29385);
nor UO_3230 (O_3230,N_29235,N_29251);
and UO_3231 (O_3231,N_29293,N_29562);
nor UO_3232 (O_3232,N_28823,N_29929);
or UO_3233 (O_3233,N_29946,N_29487);
xor UO_3234 (O_3234,N_29253,N_29642);
and UO_3235 (O_3235,N_29149,N_28909);
or UO_3236 (O_3236,N_29149,N_29530);
and UO_3237 (O_3237,N_29094,N_29402);
and UO_3238 (O_3238,N_29316,N_29783);
nor UO_3239 (O_3239,N_29935,N_29391);
nor UO_3240 (O_3240,N_29571,N_29454);
and UO_3241 (O_3241,N_29111,N_29969);
and UO_3242 (O_3242,N_29642,N_29568);
xor UO_3243 (O_3243,N_29737,N_28929);
and UO_3244 (O_3244,N_29567,N_29487);
xnor UO_3245 (O_3245,N_29211,N_28900);
xor UO_3246 (O_3246,N_29927,N_29227);
nand UO_3247 (O_3247,N_29846,N_29476);
xnor UO_3248 (O_3248,N_29611,N_29130);
and UO_3249 (O_3249,N_29295,N_29930);
or UO_3250 (O_3250,N_29812,N_29880);
and UO_3251 (O_3251,N_29741,N_28903);
nand UO_3252 (O_3252,N_29970,N_29101);
or UO_3253 (O_3253,N_29798,N_29408);
nor UO_3254 (O_3254,N_28874,N_29733);
xnor UO_3255 (O_3255,N_29085,N_29274);
xnor UO_3256 (O_3256,N_29683,N_29261);
or UO_3257 (O_3257,N_29611,N_29209);
xor UO_3258 (O_3258,N_29548,N_29283);
or UO_3259 (O_3259,N_29946,N_28841);
xnor UO_3260 (O_3260,N_29881,N_28810);
and UO_3261 (O_3261,N_29544,N_29853);
or UO_3262 (O_3262,N_29800,N_29783);
and UO_3263 (O_3263,N_29181,N_29357);
xor UO_3264 (O_3264,N_29672,N_29070);
nor UO_3265 (O_3265,N_28871,N_29925);
and UO_3266 (O_3266,N_29294,N_28946);
nor UO_3267 (O_3267,N_28885,N_29944);
nor UO_3268 (O_3268,N_28949,N_29204);
xnor UO_3269 (O_3269,N_29227,N_29846);
nor UO_3270 (O_3270,N_29925,N_28861);
nor UO_3271 (O_3271,N_29538,N_28901);
or UO_3272 (O_3272,N_29914,N_29868);
or UO_3273 (O_3273,N_29261,N_29600);
nor UO_3274 (O_3274,N_29799,N_28861);
xor UO_3275 (O_3275,N_29648,N_29157);
nand UO_3276 (O_3276,N_29572,N_29361);
xor UO_3277 (O_3277,N_29187,N_29482);
nor UO_3278 (O_3278,N_29431,N_29761);
or UO_3279 (O_3279,N_29155,N_29690);
nor UO_3280 (O_3280,N_29199,N_29838);
or UO_3281 (O_3281,N_28872,N_29858);
or UO_3282 (O_3282,N_29931,N_29628);
or UO_3283 (O_3283,N_29427,N_29644);
or UO_3284 (O_3284,N_29611,N_28836);
xnor UO_3285 (O_3285,N_29246,N_29379);
xor UO_3286 (O_3286,N_28974,N_28981);
xnor UO_3287 (O_3287,N_29741,N_29425);
and UO_3288 (O_3288,N_29917,N_29203);
nor UO_3289 (O_3289,N_29948,N_28979);
nor UO_3290 (O_3290,N_29779,N_29078);
or UO_3291 (O_3291,N_29602,N_29571);
nand UO_3292 (O_3292,N_29385,N_29625);
or UO_3293 (O_3293,N_29102,N_29533);
and UO_3294 (O_3294,N_29824,N_29474);
nand UO_3295 (O_3295,N_29849,N_29915);
nor UO_3296 (O_3296,N_29786,N_29651);
and UO_3297 (O_3297,N_29812,N_29080);
xnor UO_3298 (O_3298,N_29825,N_29683);
xor UO_3299 (O_3299,N_29251,N_28807);
and UO_3300 (O_3300,N_29085,N_29094);
and UO_3301 (O_3301,N_29704,N_29154);
and UO_3302 (O_3302,N_29982,N_29951);
and UO_3303 (O_3303,N_29476,N_29283);
and UO_3304 (O_3304,N_29108,N_29704);
and UO_3305 (O_3305,N_28805,N_28871);
and UO_3306 (O_3306,N_28813,N_29199);
and UO_3307 (O_3307,N_29539,N_29788);
nor UO_3308 (O_3308,N_28880,N_28945);
xor UO_3309 (O_3309,N_29471,N_28901);
nand UO_3310 (O_3310,N_29124,N_29811);
nand UO_3311 (O_3311,N_28919,N_29175);
and UO_3312 (O_3312,N_29284,N_29425);
xnor UO_3313 (O_3313,N_28834,N_29823);
nand UO_3314 (O_3314,N_29703,N_28828);
or UO_3315 (O_3315,N_29770,N_28971);
or UO_3316 (O_3316,N_28952,N_28914);
nand UO_3317 (O_3317,N_29549,N_29431);
nor UO_3318 (O_3318,N_29117,N_29823);
nor UO_3319 (O_3319,N_29082,N_29014);
nand UO_3320 (O_3320,N_29350,N_29546);
xor UO_3321 (O_3321,N_28959,N_29793);
xor UO_3322 (O_3322,N_28824,N_29283);
nor UO_3323 (O_3323,N_29083,N_29897);
nor UO_3324 (O_3324,N_29187,N_28876);
or UO_3325 (O_3325,N_29038,N_29757);
or UO_3326 (O_3326,N_29172,N_29884);
and UO_3327 (O_3327,N_29662,N_29684);
or UO_3328 (O_3328,N_29569,N_29846);
nor UO_3329 (O_3329,N_29098,N_29654);
nand UO_3330 (O_3330,N_29299,N_29678);
nor UO_3331 (O_3331,N_28924,N_28838);
nor UO_3332 (O_3332,N_29411,N_28969);
nor UO_3333 (O_3333,N_29735,N_29813);
and UO_3334 (O_3334,N_29185,N_29833);
and UO_3335 (O_3335,N_29652,N_29533);
nand UO_3336 (O_3336,N_29911,N_29726);
nor UO_3337 (O_3337,N_29999,N_29622);
and UO_3338 (O_3338,N_28874,N_29117);
or UO_3339 (O_3339,N_29172,N_29525);
nand UO_3340 (O_3340,N_28829,N_29425);
and UO_3341 (O_3341,N_29382,N_29609);
or UO_3342 (O_3342,N_29170,N_29084);
xor UO_3343 (O_3343,N_29789,N_29667);
nand UO_3344 (O_3344,N_29585,N_29191);
and UO_3345 (O_3345,N_29787,N_29555);
xnor UO_3346 (O_3346,N_29253,N_29171);
xnor UO_3347 (O_3347,N_29447,N_29065);
nand UO_3348 (O_3348,N_29659,N_28996);
nand UO_3349 (O_3349,N_29636,N_29182);
xor UO_3350 (O_3350,N_29740,N_29122);
nand UO_3351 (O_3351,N_29556,N_28815);
xnor UO_3352 (O_3352,N_29086,N_29523);
nand UO_3353 (O_3353,N_29741,N_28867);
or UO_3354 (O_3354,N_29866,N_29464);
nor UO_3355 (O_3355,N_29910,N_29881);
nand UO_3356 (O_3356,N_29450,N_29056);
and UO_3357 (O_3357,N_29357,N_29703);
nand UO_3358 (O_3358,N_28872,N_29941);
nand UO_3359 (O_3359,N_28920,N_29159);
or UO_3360 (O_3360,N_29512,N_29733);
or UO_3361 (O_3361,N_29680,N_29726);
nor UO_3362 (O_3362,N_29944,N_29342);
nand UO_3363 (O_3363,N_29100,N_29132);
nand UO_3364 (O_3364,N_29567,N_29994);
or UO_3365 (O_3365,N_29929,N_28872);
or UO_3366 (O_3366,N_29210,N_28996);
xor UO_3367 (O_3367,N_29055,N_28812);
and UO_3368 (O_3368,N_29122,N_29728);
or UO_3369 (O_3369,N_29711,N_29203);
and UO_3370 (O_3370,N_29623,N_29463);
xor UO_3371 (O_3371,N_29918,N_29100);
or UO_3372 (O_3372,N_29877,N_28866);
xnor UO_3373 (O_3373,N_29253,N_29507);
nand UO_3374 (O_3374,N_28818,N_29732);
nor UO_3375 (O_3375,N_29400,N_29190);
nand UO_3376 (O_3376,N_29227,N_29011);
xor UO_3377 (O_3377,N_29594,N_29654);
or UO_3378 (O_3378,N_29745,N_29919);
nor UO_3379 (O_3379,N_29578,N_29788);
nand UO_3380 (O_3380,N_29820,N_28828);
and UO_3381 (O_3381,N_29503,N_29462);
xor UO_3382 (O_3382,N_29806,N_29555);
nand UO_3383 (O_3383,N_29333,N_28928);
xor UO_3384 (O_3384,N_29165,N_29327);
xor UO_3385 (O_3385,N_29276,N_29335);
and UO_3386 (O_3386,N_29267,N_28935);
xnor UO_3387 (O_3387,N_29111,N_29746);
xor UO_3388 (O_3388,N_29420,N_29562);
and UO_3389 (O_3389,N_29634,N_29462);
and UO_3390 (O_3390,N_29611,N_29877);
nand UO_3391 (O_3391,N_29903,N_29911);
nor UO_3392 (O_3392,N_29359,N_29454);
or UO_3393 (O_3393,N_29997,N_29202);
and UO_3394 (O_3394,N_29413,N_29548);
or UO_3395 (O_3395,N_29389,N_29223);
nand UO_3396 (O_3396,N_29165,N_29186);
nand UO_3397 (O_3397,N_28839,N_28837);
nand UO_3398 (O_3398,N_29600,N_28896);
or UO_3399 (O_3399,N_29632,N_29596);
and UO_3400 (O_3400,N_29826,N_29572);
and UO_3401 (O_3401,N_29756,N_29215);
xor UO_3402 (O_3402,N_29018,N_28954);
or UO_3403 (O_3403,N_29214,N_29999);
xnor UO_3404 (O_3404,N_29853,N_28974);
xor UO_3405 (O_3405,N_28906,N_29330);
xnor UO_3406 (O_3406,N_29824,N_29983);
nor UO_3407 (O_3407,N_29697,N_29286);
and UO_3408 (O_3408,N_29344,N_29331);
nor UO_3409 (O_3409,N_29329,N_28908);
and UO_3410 (O_3410,N_29288,N_28893);
and UO_3411 (O_3411,N_29624,N_28922);
nand UO_3412 (O_3412,N_29836,N_29765);
nor UO_3413 (O_3413,N_29136,N_29349);
xnor UO_3414 (O_3414,N_29615,N_29688);
xnor UO_3415 (O_3415,N_29635,N_28938);
nand UO_3416 (O_3416,N_29676,N_29539);
and UO_3417 (O_3417,N_29047,N_29252);
xnor UO_3418 (O_3418,N_29939,N_29576);
xnor UO_3419 (O_3419,N_28911,N_29126);
xnor UO_3420 (O_3420,N_29990,N_29492);
or UO_3421 (O_3421,N_29109,N_29415);
xor UO_3422 (O_3422,N_28942,N_29936);
nand UO_3423 (O_3423,N_29933,N_29878);
and UO_3424 (O_3424,N_29418,N_29302);
or UO_3425 (O_3425,N_29774,N_29369);
nand UO_3426 (O_3426,N_29945,N_29589);
nand UO_3427 (O_3427,N_28890,N_28895);
nor UO_3428 (O_3428,N_28877,N_29668);
xnor UO_3429 (O_3429,N_28890,N_29577);
or UO_3430 (O_3430,N_29840,N_29995);
or UO_3431 (O_3431,N_29682,N_28967);
nand UO_3432 (O_3432,N_29887,N_29373);
nand UO_3433 (O_3433,N_29315,N_29880);
or UO_3434 (O_3434,N_29056,N_29198);
nand UO_3435 (O_3435,N_28854,N_29789);
or UO_3436 (O_3436,N_29278,N_29733);
xor UO_3437 (O_3437,N_29479,N_29534);
nand UO_3438 (O_3438,N_29841,N_29025);
nand UO_3439 (O_3439,N_29327,N_29328);
nand UO_3440 (O_3440,N_29843,N_29129);
and UO_3441 (O_3441,N_29782,N_29432);
nor UO_3442 (O_3442,N_29290,N_29390);
and UO_3443 (O_3443,N_29247,N_29602);
nand UO_3444 (O_3444,N_29535,N_29449);
or UO_3445 (O_3445,N_29493,N_29624);
xor UO_3446 (O_3446,N_28823,N_29815);
and UO_3447 (O_3447,N_29529,N_29721);
nand UO_3448 (O_3448,N_29431,N_29038);
nor UO_3449 (O_3449,N_29286,N_29986);
and UO_3450 (O_3450,N_29335,N_28949);
nand UO_3451 (O_3451,N_28953,N_29706);
xnor UO_3452 (O_3452,N_29220,N_29350);
nor UO_3453 (O_3453,N_29153,N_29554);
nand UO_3454 (O_3454,N_29414,N_29186);
nand UO_3455 (O_3455,N_29284,N_29587);
nor UO_3456 (O_3456,N_29320,N_29049);
and UO_3457 (O_3457,N_29092,N_29424);
or UO_3458 (O_3458,N_29672,N_29179);
and UO_3459 (O_3459,N_28829,N_29740);
nor UO_3460 (O_3460,N_29530,N_28893);
xor UO_3461 (O_3461,N_29615,N_29989);
or UO_3462 (O_3462,N_29638,N_29147);
xnor UO_3463 (O_3463,N_29221,N_29727);
nand UO_3464 (O_3464,N_29150,N_28889);
and UO_3465 (O_3465,N_29484,N_29273);
xnor UO_3466 (O_3466,N_29794,N_29750);
or UO_3467 (O_3467,N_29792,N_29724);
nand UO_3468 (O_3468,N_29278,N_29087);
nand UO_3469 (O_3469,N_29920,N_28811);
nand UO_3470 (O_3470,N_28959,N_29538);
nor UO_3471 (O_3471,N_29441,N_29374);
and UO_3472 (O_3472,N_29186,N_29028);
and UO_3473 (O_3473,N_29135,N_29848);
and UO_3474 (O_3474,N_29326,N_28826);
and UO_3475 (O_3475,N_28937,N_28808);
nand UO_3476 (O_3476,N_29071,N_29539);
nor UO_3477 (O_3477,N_29012,N_28803);
nor UO_3478 (O_3478,N_29897,N_29710);
xor UO_3479 (O_3479,N_29150,N_29898);
or UO_3480 (O_3480,N_29602,N_29018);
nand UO_3481 (O_3481,N_29791,N_29001);
and UO_3482 (O_3482,N_29813,N_29915);
xnor UO_3483 (O_3483,N_29583,N_29205);
or UO_3484 (O_3484,N_29682,N_29131);
nand UO_3485 (O_3485,N_29806,N_29617);
or UO_3486 (O_3486,N_29436,N_29787);
and UO_3487 (O_3487,N_29260,N_29834);
xnor UO_3488 (O_3488,N_29714,N_29273);
nor UO_3489 (O_3489,N_29008,N_29576);
xor UO_3490 (O_3490,N_29817,N_29079);
nand UO_3491 (O_3491,N_29202,N_29948);
nor UO_3492 (O_3492,N_29924,N_29134);
xnor UO_3493 (O_3493,N_29874,N_29175);
or UO_3494 (O_3494,N_29727,N_28850);
nand UO_3495 (O_3495,N_29169,N_29551);
xor UO_3496 (O_3496,N_29132,N_29455);
nand UO_3497 (O_3497,N_29504,N_29557);
nor UO_3498 (O_3498,N_29504,N_29923);
nand UO_3499 (O_3499,N_29771,N_29642);
endmodule