module basic_3000_30000_3500_100_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nand U0 (N_0,In_204,In_256);
nor U1 (N_1,In_632,In_875);
nor U2 (N_2,In_1221,In_1840);
xnor U3 (N_3,In_143,In_326);
or U4 (N_4,In_181,In_212);
nor U5 (N_5,In_464,In_766);
nor U6 (N_6,In_2025,In_1694);
nand U7 (N_7,In_835,In_941);
nor U8 (N_8,In_1501,In_2444);
or U9 (N_9,In_1218,In_849);
nor U10 (N_10,In_284,In_365);
or U11 (N_11,In_1096,In_183);
xor U12 (N_12,In_1527,In_211);
and U13 (N_13,In_2091,In_2173);
nand U14 (N_14,In_1627,In_981);
nor U15 (N_15,In_2574,In_2467);
xnor U16 (N_16,In_1749,In_1074);
nor U17 (N_17,In_1412,In_2786);
nor U18 (N_18,In_2503,In_1640);
xor U19 (N_19,In_1498,In_2032);
xor U20 (N_20,In_313,In_1024);
and U21 (N_21,In_568,In_1438);
xor U22 (N_22,In_682,In_1531);
nand U23 (N_23,In_2551,In_1953);
or U24 (N_24,In_1831,In_2047);
nor U25 (N_25,In_778,In_346);
nand U26 (N_26,In_1827,In_2135);
nor U27 (N_27,In_1746,In_1255);
nor U28 (N_28,In_548,In_2908);
and U29 (N_29,In_1951,In_271);
or U30 (N_30,In_2204,In_2322);
nor U31 (N_31,In_1852,In_1509);
nor U32 (N_32,In_536,In_1044);
xnor U33 (N_33,In_2427,In_801);
or U34 (N_34,In_2619,In_208);
or U35 (N_35,In_2363,In_1942);
nand U36 (N_36,In_2562,In_342);
nand U37 (N_37,In_2816,In_2239);
and U38 (N_38,In_852,In_2184);
or U39 (N_39,In_1443,In_1272);
nor U40 (N_40,In_215,In_391);
nor U41 (N_41,In_1916,In_1367);
nor U42 (N_42,In_2585,In_1866);
or U43 (N_43,In_2568,In_531);
or U44 (N_44,In_2354,In_2663);
xor U45 (N_45,In_218,In_2766);
nand U46 (N_46,In_2477,In_2861);
xor U47 (N_47,In_2845,In_279);
or U48 (N_48,In_347,In_2620);
xnor U49 (N_49,In_805,In_914);
nand U50 (N_50,In_2917,In_1517);
nor U51 (N_51,In_1000,In_1493);
nand U52 (N_52,In_2259,In_1086);
nand U53 (N_53,In_1383,In_174);
and U54 (N_54,In_1600,In_483);
nor U55 (N_55,In_2045,In_676);
nand U56 (N_56,In_422,In_1379);
and U57 (N_57,In_1394,In_2633);
nor U58 (N_58,In_657,In_1804);
and U59 (N_59,In_7,In_84);
xnor U60 (N_60,In_2144,In_1664);
nand U61 (N_61,In_675,In_2208);
or U62 (N_62,In_1459,In_2280);
or U63 (N_63,In_1909,In_1109);
nand U64 (N_64,In_268,In_2815);
or U65 (N_65,In_2634,In_2511);
and U66 (N_66,In_1904,In_2145);
nand U67 (N_67,In_1392,In_1043);
xnor U68 (N_68,In_1279,In_1828);
nand U69 (N_69,In_1823,In_1830);
nand U70 (N_70,In_1243,In_1005);
nor U71 (N_71,In_927,In_2580);
xnor U72 (N_72,In_1956,In_468);
and U73 (N_73,In_1097,In_1970);
xor U74 (N_74,In_2946,In_824);
nor U75 (N_75,In_2000,In_586);
nor U76 (N_76,In_2106,In_2901);
and U77 (N_77,In_309,In_2887);
and U78 (N_78,In_2252,In_2903);
nor U79 (N_79,In_2054,In_686);
nand U80 (N_80,In_1886,In_1620);
and U81 (N_81,In_1770,In_104);
and U82 (N_82,In_2851,In_1336);
and U83 (N_83,In_1399,In_721);
and U84 (N_84,In_2140,In_1729);
or U85 (N_85,In_1084,In_2429);
and U86 (N_86,In_2179,In_60);
nand U87 (N_87,In_153,In_519);
nand U88 (N_88,In_2207,In_293);
nand U89 (N_89,In_1666,In_1768);
xnor U90 (N_90,In_2423,In_2066);
or U91 (N_91,In_2577,In_2436);
or U92 (N_92,In_1519,In_2976);
nor U93 (N_93,In_1302,In_125);
nor U94 (N_94,In_1662,In_2027);
xor U95 (N_95,In_2048,In_2369);
and U96 (N_96,In_2166,In_1765);
and U97 (N_97,In_2157,In_564);
or U98 (N_98,In_2463,In_2883);
or U99 (N_99,In_2127,In_785);
xor U100 (N_100,In_2198,In_2717);
and U101 (N_101,In_1069,In_2412);
nand U102 (N_102,In_2142,In_2266);
xnor U103 (N_103,In_1717,In_2933);
or U104 (N_104,In_946,In_2332);
and U105 (N_105,In_168,In_1502);
or U106 (N_106,In_609,In_1688);
nor U107 (N_107,In_2460,In_396);
and U108 (N_108,In_2833,In_2117);
or U109 (N_109,In_1755,In_1888);
and U110 (N_110,In_2616,In_631);
and U111 (N_111,In_2922,In_1016);
xnor U112 (N_112,In_2793,In_1108);
or U113 (N_113,In_2508,In_2549);
nand U114 (N_114,In_2308,In_1982);
xor U115 (N_115,In_1914,In_1801);
and U116 (N_116,In_950,In_407);
nor U117 (N_117,In_1534,In_596);
nor U118 (N_118,In_59,In_2393);
or U119 (N_119,In_2760,In_2488);
nor U120 (N_120,In_2818,In_2489);
nor U121 (N_121,In_1208,In_2645);
xor U122 (N_122,In_2141,In_566);
xor U123 (N_123,In_304,In_255);
xnor U124 (N_124,In_1187,In_1264);
nand U125 (N_125,In_2298,In_2773);
nor U126 (N_126,In_86,In_2124);
nor U127 (N_127,In_1565,In_1997);
and U128 (N_128,In_1633,In_160);
nor U129 (N_129,In_2046,In_1722);
nand U130 (N_130,In_2934,In_1168);
nor U131 (N_131,In_1899,In_508);
nand U132 (N_132,In_791,In_113);
nor U133 (N_133,In_736,In_6);
xnor U134 (N_134,In_2559,In_413);
xnor U135 (N_135,In_2727,In_913);
and U136 (N_136,In_2240,In_1683);
or U137 (N_137,In_1748,In_1071);
xor U138 (N_138,In_307,In_1146);
nor U139 (N_139,In_2176,In_348);
nand U140 (N_140,In_2679,In_565);
or U141 (N_141,In_599,In_1485);
nor U142 (N_142,In_1815,In_1988);
nor U143 (N_143,In_1460,In_2737);
nor U144 (N_144,In_992,In_1891);
and U145 (N_145,In_1607,In_1661);
or U146 (N_146,In_2673,In_2992);
nor U147 (N_147,In_699,In_452);
nand U148 (N_148,In_2509,In_1156);
nor U149 (N_149,In_2019,In_1373);
and U150 (N_150,In_2703,In_1338);
nand U151 (N_151,In_247,In_329);
nand U152 (N_152,In_896,In_1969);
xor U153 (N_153,In_1358,In_2328);
nor U154 (N_154,In_1140,In_597);
or U155 (N_155,In_2235,In_1349);
nor U156 (N_156,In_2878,In_1783);
and U157 (N_157,In_1564,In_196);
or U158 (N_158,In_772,In_2401);
and U159 (N_159,In_2081,In_547);
nand U160 (N_160,In_2797,In_2279);
xor U161 (N_161,In_2012,In_2312);
xor U162 (N_162,In_986,In_2648);
xor U163 (N_163,In_1833,In_2704);
or U164 (N_164,In_1881,In_2109);
and U165 (N_165,In_1781,In_1980);
or U166 (N_166,In_2635,In_2899);
nand U167 (N_167,In_1950,In_487);
xor U168 (N_168,In_1482,In_975);
nor U169 (N_169,In_1769,In_2813);
nor U170 (N_170,In_2195,In_361);
xor U171 (N_171,In_2411,In_67);
and U172 (N_172,In_192,In_2161);
nor U173 (N_173,In_1305,In_915);
or U174 (N_174,In_1491,In_729);
or U175 (N_175,In_2864,In_735);
nand U176 (N_176,In_262,In_2591);
nand U177 (N_177,In_1621,In_1319);
nand U178 (N_178,In_2458,In_2940);
nand U179 (N_179,In_2457,In_1282);
xnor U180 (N_180,In_260,In_2092);
and U181 (N_181,In_1713,In_945);
and U182 (N_182,In_2264,In_2935);
and U183 (N_183,In_1861,In_2691);
and U184 (N_184,In_1719,In_1647);
nor U185 (N_185,In_1613,In_674);
or U186 (N_186,In_512,In_2008);
and U187 (N_187,In_2880,In_867);
xnor U188 (N_188,In_1925,In_2217);
nor U189 (N_189,In_2487,In_206);
and U190 (N_190,In_1316,In_497);
or U191 (N_191,In_1111,In_2267);
and U192 (N_192,In_2599,In_990);
nand U193 (N_193,In_403,In_1428);
nor U194 (N_194,In_795,In_641);
and U195 (N_195,In_1732,In_621);
nor U196 (N_196,In_1691,In_108);
nor U197 (N_197,In_1271,In_924);
xor U198 (N_198,In_1464,In_569);
or U199 (N_199,In_239,In_2228);
nor U200 (N_200,In_745,In_2802);
and U201 (N_201,In_2819,In_1001);
and U202 (N_202,In_576,In_534);
nand U203 (N_203,In_2755,In_2974);
or U204 (N_204,In_2768,In_594);
or U205 (N_205,In_461,In_2534);
xor U206 (N_206,In_1227,In_38);
and U207 (N_207,In_1500,In_722);
or U208 (N_208,In_1018,In_1669);
nand U209 (N_209,In_219,In_2699);
or U210 (N_210,In_2521,In_1064);
or U211 (N_211,In_274,In_1263);
nor U212 (N_212,In_1427,In_1216);
xor U213 (N_213,In_302,In_864);
xor U214 (N_214,In_54,In_213);
nor U215 (N_215,In_291,In_1849);
and U216 (N_216,In_1210,In_861);
or U217 (N_217,In_1308,In_2849);
xnor U218 (N_218,In_2783,In_1289);
xor U219 (N_219,In_886,In_444);
xnor U220 (N_220,In_1575,In_1476);
or U221 (N_221,In_387,In_640);
or U222 (N_222,In_475,In_2447);
and U223 (N_223,In_1526,In_502);
nor U224 (N_224,In_1386,In_433);
and U225 (N_225,In_1674,In_254);
and U226 (N_226,In_2300,In_267);
or U227 (N_227,In_644,In_1405);
or U228 (N_228,In_1961,In_1555);
xnor U229 (N_229,In_770,In_1573);
nand U230 (N_230,In_905,In_767);
nor U231 (N_231,In_393,In_455);
xor U232 (N_232,In_1578,In_250);
and U233 (N_233,In_1177,In_1644);
or U234 (N_234,In_661,In_2218);
nor U235 (N_235,In_1703,In_199);
or U236 (N_236,In_1229,In_121);
nand U237 (N_237,In_2624,In_523);
xor U238 (N_238,In_2398,In_24);
nor U239 (N_239,In_303,In_2594);
nand U240 (N_240,In_2131,In_1400);
xor U241 (N_241,In_1658,In_1230);
and U242 (N_242,In_462,In_101);
and U243 (N_243,In_2897,In_2491);
and U244 (N_244,In_39,In_771);
and U245 (N_245,In_1780,In_2909);
or U246 (N_246,In_2483,In_1137);
and U247 (N_247,In_720,In_740);
xor U248 (N_248,In_639,In_882);
or U249 (N_249,In_360,In_625);
nor U250 (N_250,In_2547,In_1601);
or U251 (N_251,In_1442,In_2099);
and U252 (N_252,In_2852,In_1967);
xor U253 (N_253,In_1039,In_149);
nand U254 (N_254,In_2804,In_294);
xor U255 (N_255,In_718,In_1196);
nand U256 (N_256,In_131,In_2246);
nor U257 (N_257,In_926,In_923);
or U258 (N_258,In_1791,In_2015);
and U259 (N_259,In_763,In_1424);
nor U260 (N_260,In_506,In_976);
xnor U261 (N_261,In_585,In_593);
nand U262 (N_262,In_2567,In_2350);
or U263 (N_263,In_2282,In_636);
and U264 (N_264,In_1013,In_2573);
or U265 (N_265,In_349,In_1774);
nand U266 (N_266,In_1309,In_2998);
nor U267 (N_267,In_2834,In_465);
nor U268 (N_268,In_1634,In_41);
or U269 (N_269,In_622,In_822);
or U270 (N_270,In_1716,In_1790);
or U271 (N_271,In_50,In_1310);
or U272 (N_272,In_1843,In_1);
nor U273 (N_273,In_2021,In_2630);
and U274 (N_274,In_1119,In_2847);
or U275 (N_275,In_2628,In_894);
nand U276 (N_276,In_2516,In_2017);
nor U277 (N_277,In_1511,In_934);
xnor U278 (N_278,In_2010,In_2979);
nor U279 (N_279,In_2656,In_2469);
nand U280 (N_280,In_2471,In_2995);
and U281 (N_281,In_2623,In_1083);
and U282 (N_282,In_1035,In_2096);
or U283 (N_283,In_25,In_844);
or U284 (N_284,In_1902,In_2347);
nor U285 (N_285,In_2669,In_266);
nand U286 (N_286,In_742,In_1080);
nor U287 (N_287,In_994,In_1435);
and U288 (N_288,In_1462,In_2366);
or U289 (N_289,In_774,In_2074);
xor U290 (N_290,In_2103,In_110);
or U291 (N_291,In_1470,In_1418);
and U292 (N_292,In_1085,In_2808);
nand U293 (N_293,In_2806,In_2983);
or U294 (N_294,In_825,In_1265);
xnor U295 (N_295,In_1439,In_330);
and U296 (N_296,In_840,In_1268);
nand U297 (N_297,In_856,In_575);
xnor U298 (N_298,In_1877,In_2285);
and U299 (N_299,In_2653,In_2225);
xnor U300 (N_300,In_51,In_2517);
nand U301 (N_301,In_2771,In_301);
nor U302 (N_302,In_747,In_671);
or U303 (N_303,In_1739,In_2380);
or U304 (N_304,In_2675,In_2924);
xor U305 (N_305,In_901,In_2890);
nor U306 (N_306,In_684,N_261);
nand U307 (N_307,In_1047,N_28);
and U308 (N_308,In_482,In_2943);
and U309 (N_309,In_1672,In_535);
nand U310 (N_310,In_1503,In_1567);
or U311 (N_311,N_210,In_2073);
nand U312 (N_312,In_33,In_1200);
and U313 (N_313,In_1617,In_2877);
xnor U314 (N_314,In_1477,In_2188);
and U315 (N_315,In_873,In_2070);
nor U316 (N_316,In_704,In_1276);
and U317 (N_317,N_152,In_270);
or U318 (N_318,In_749,In_1467);
or U319 (N_319,In_138,In_2676);
or U320 (N_320,In_1454,In_411);
and U321 (N_321,In_618,In_1597);
or U322 (N_322,In_2557,In_490);
nand U323 (N_323,In_2906,In_2809);
or U324 (N_324,In_1700,In_1913);
xnor U325 (N_325,In_1908,In_2371);
nand U326 (N_326,In_1553,In_1247);
xor U327 (N_327,In_1205,In_1903);
or U328 (N_328,In_1262,In_1976);
xor U329 (N_329,N_292,In_1935);
nand U330 (N_330,In_91,In_1639);
nor U331 (N_331,In_2297,In_1298);
and U332 (N_332,In_2111,In_2360);
and U333 (N_333,In_1189,In_2514);
nor U334 (N_334,In_2788,In_787);
xor U335 (N_335,In_1510,In_253);
or U336 (N_336,In_2082,In_2746);
nand U337 (N_337,N_279,In_1887);
xor U338 (N_338,In_2452,In_2478);
and U339 (N_339,In_2595,In_451);
and U340 (N_340,In_1117,In_725);
and U341 (N_341,In_1174,In_2622);
xor U342 (N_342,In_2842,In_2132);
or U343 (N_343,In_1257,In_779);
nor U344 (N_344,In_2529,In_1584);
and U345 (N_345,In_792,N_129);
nand U346 (N_346,In_647,In_762);
nor U347 (N_347,In_2545,In_2378);
xor U348 (N_348,In_2957,In_2163);
nor U349 (N_349,In_2598,In_2868);
xor U350 (N_350,In_2807,In_2453);
xor U351 (N_351,In_16,In_1110);
or U352 (N_352,In_2201,In_0);
xnor U353 (N_353,In_1242,In_1608);
and U354 (N_354,N_40,In_1995);
or U355 (N_355,In_1816,In_1458);
and U356 (N_356,In_904,In_495);
nor U357 (N_357,In_2925,In_258);
nor U358 (N_358,In_532,In_1591);
and U359 (N_359,In_2698,N_240);
xnor U360 (N_360,In_2171,In_2697);
nor U361 (N_361,In_814,In_985);
or U362 (N_362,In_173,N_190);
xnor U363 (N_363,In_760,In_1807);
and U364 (N_364,In_1354,In_1721);
nor U365 (N_365,In_1017,N_110);
xor U366 (N_366,In_2346,In_134);
nor U367 (N_367,In_2642,In_362);
nor U368 (N_368,In_300,In_1619);
xnor U369 (N_369,In_1277,In_1609);
and U370 (N_370,In_764,In_1579);
nand U371 (N_371,In_1051,In_1157);
nor U372 (N_372,In_2647,In_1267);
nor U373 (N_373,In_1274,In_591);
and U374 (N_374,In_344,In_2715);
and U375 (N_375,In_187,In_370);
or U376 (N_376,In_30,In_2168);
nor U377 (N_377,In_2915,In_2859);
or U378 (N_378,In_572,N_258);
or U379 (N_379,In_2997,In_8);
or U380 (N_380,In_1580,In_2058);
and U381 (N_381,In_1735,In_1677);
or U382 (N_382,In_2579,In_1934);
or U383 (N_383,In_751,In_2146);
or U384 (N_384,In_1488,In_2189);
nand U385 (N_385,In_558,In_1102);
and U386 (N_386,N_212,In_99);
nor U387 (N_387,In_1215,In_1931);
and U388 (N_388,In_2299,In_129);
nor U389 (N_389,In_1046,In_1286);
nand U390 (N_390,In_1824,In_405);
nor U391 (N_391,In_2197,In_1994);
or U392 (N_392,In_1602,N_36);
nor U393 (N_393,In_2667,In_898);
xor U394 (N_394,N_270,In_2561);
and U395 (N_395,In_1451,In_2970);
nand U396 (N_396,In_150,In_2353);
and U397 (N_397,In_200,In_1241);
nand U398 (N_398,N_1,In_1468);
xor U399 (N_399,In_2482,In_1456);
or U400 (N_400,In_2973,In_2428);
xor U401 (N_401,In_1876,In_2740);
nand U402 (N_402,In_2836,In_2515);
and U403 (N_403,In_102,In_2442);
nand U404 (N_404,In_1809,In_2410);
nand U405 (N_405,In_2694,In_2982);
nor U406 (N_406,In_2400,In_311);
or U407 (N_407,In_1390,In_865);
nor U408 (N_408,In_1368,N_90);
or U409 (N_409,In_448,In_2250);
nor U410 (N_410,In_2636,In_1297);
or U411 (N_411,In_731,In_1287);
xnor U412 (N_412,In_963,In_887);
xor U413 (N_413,In_1540,In_2650);
xnor U414 (N_414,In_257,In_533);
nand U415 (N_415,In_2067,In_557);
nor U416 (N_416,In_1760,N_65);
or U417 (N_417,In_550,In_191);
and U418 (N_418,In_117,In_1371);
nand U419 (N_419,In_456,In_443);
xor U420 (N_420,In_540,In_697);
xor U421 (N_421,In_1123,In_663);
nor U422 (N_422,In_62,In_1432);
or U423 (N_423,In_571,In_2749);
and U424 (N_424,In_2437,In_188);
and U425 (N_425,In_1325,In_1433);
nor U426 (N_426,In_1372,In_2014);
nor U427 (N_427,In_2537,In_106);
or U428 (N_428,In_2831,In_2961);
nor U429 (N_429,In_1975,In_1183);
and U430 (N_430,In_828,In_2211);
xnor U431 (N_431,In_570,In_1124);
or U432 (N_432,In_310,In_1958);
nor U433 (N_433,In_2719,In_953);
xnor U434 (N_434,In_55,In_2200);
nand U435 (N_435,N_31,In_2661);
nor U436 (N_436,In_2754,N_58);
or U437 (N_437,N_246,In_2958);
xor U438 (N_438,In_1240,In_2147);
nand U439 (N_439,In_1269,In_1740);
and U440 (N_440,In_1714,In_1731);
nor U441 (N_441,In_1965,In_1351);
nand U442 (N_442,In_36,In_2702);
nand U443 (N_443,In_2513,In_1201);
xor U444 (N_444,In_1176,In_2914);
nor U445 (N_445,In_77,In_706);
nand U446 (N_446,N_215,In_1550);
nand U447 (N_447,In_2778,N_264);
and U448 (N_448,In_386,In_1594);
nand U449 (N_449,N_238,In_1948);
nor U450 (N_450,In_2985,In_730);
or U451 (N_451,In_1198,N_177);
nor U452 (N_452,In_1754,In_1733);
nor U453 (N_453,In_2563,In_1614);
nand U454 (N_454,In_1366,In_803);
and U455 (N_455,In_988,In_234);
or U456 (N_456,In_2098,In_2921);
xor U457 (N_457,In_956,N_267);
and U458 (N_458,In_942,In_385);
xnor U459 (N_459,In_820,In_2938);
nor U460 (N_460,In_694,In_551);
nand U461 (N_461,In_2989,In_733);
or U462 (N_462,In_1270,N_281);
nor U463 (N_463,In_440,In_724);
and U464 (N_464,In_2576,In_1258);
or U465 (N_465,In_2586,In_2375);
nand U466 (N_466,In_2911,In_673);
xnor U467 (N_467,In_434,In_135);
and U468 (N_468,In_1589,In_524);
nand U469 (N_469,N_59,In_2451);
or U470 (N_470,In_1989,In_1892);
nor U471 (N_471,In_1962,In_2261);
nor U472 (N_472,In_966,In_574);
xor U473 (N_473,In_665,In_515);
and U474 (N_474,In_2884,In_759);
and U475 (N_475,In_1420,In_2219);
nor U476 (N_476,In_343,In_1068);
nor U477 (N_477,N_27,N_293);
nand U478 (N_478,In_1179,N_234);
and U479 (N_479,In_1549,In_2448);
or U480 (N_480,In_522,N_298);
nand U481 (N_481,In_626,In_637);
nor U482 (N_482,In_2284,In_2062);
or U483 (N_483,In_2381,In_2575);
nand U484 (N_484,In_2268,In_64);
xor U485 (N_485,In_1545,N_184);
and U486 (N_486,In_2782,N_96);
or U487 (N_487,In_1105,In_2986);
and U488 (N_488,N_55,In_2657);
and U489 (N_489,In_1663,In_2449);
nor U490 (N_490,In_431,In_2629);
nor U491 (N_491,In_10,N_68);
nor U492 (N_492,In_2061,In_2687);
nand U493 (N_493,N_260,In_648);
xor U494 (N_494,In_623,In_114);
nor U495 (N_495,In_154,In_2175);
or U496 (N_496,In_94,In_949);
and U497 (N_497,In_120,In_579);
or U498 (N_498,In_1894,In_969);
and U499 (N_499,In_1693,In_2876);
nand U500 (N_500,In_1003,N_14);
nand U501 (N_501,In_2024,In_421);
and U502 (N_502,In_2343,In_1763);
nor U503 (N_503,In_813,In_2714);
or U504 (N_504,In_1859,In_2817);
xnor U505 (N_505,In_1558,In_1655);
nor U506 (N_506,In_2214,In_1330);
nand U507 (N_507,In_2222,In_2869);
xor U508 (N_508,In_220,N_115);
nand U509 (N_509,In_757,N_290);
or U510 (N_510,N_243,In_2572);
nor U511 (N_511,In_406,In_800);
nand U512 (N_512,In_932,In_2858);
and U513 (N_513,In_627,In_2040);
and U514 (N_514,In_1014,In_127);
xor U515 (N_515,In_1727,In_2077);
xnor U516 (N_516,In_1128,N_132);
and U517 (N_517,In_2180,In_2951);
or U518 (N_518,In_20,In_855);
nand U519 (N_519,In_1736,In_1022);
xor U520 (N_520,In_837,N_122);
or U521 (N_521,In_1598,In_1805);
nor U522 (N_522,N_256,In_210);
or U523 (N_523,In_2203,In_1422);
or U524 (N_524,In_1800,In_2383);
or U525 (N_525,In_1237,In_2318);
or U526 (N_526,In_72,In_2368);
nand U527 (N_527,In_646,In_398);
or U528 (N_528,In_1126,N_266);
nand U529 (N_529,In_826,In_1250);
and U530 (N_530,In_859,In_1341);
and U531 (N_531,In_1818,In_1008);
nand U532 (N_532,In_1088,In_235);
nor U533 (N_533,In_264,N_80);
xor U534 (N_534,In_1786,In_1730);
nor U535 (N_535,N_166,In_2611);
nor U536 (N_536,In_2523,In_1955);
or U537 (N_537,In_2525,N_111);
nor U538 (N_538,In_1789,N_153);
xnor U539 (N_539,In_798,In_1963);
or U540 (N_540,In_2659,N_12);
nor U541 (N_541,N_66,In_155);
xor U542 (N_542,In_463,N_183);
nand U543 (N_543,In_1239,In_1949);
nor U544 (N_544,In_1642,In_198);
and U545 (N_545,In_1012,In_2734);
xor U546 (N_546,In_2455,In_2242);
and U547 (N_547,In_2334,In_1184);
xnor U548 (N_548,In_2756,In_2030);
xor U549 (N_549,N_107,In_2932);
nor U550 (N_550,In_1928,In_2419);
xor U551 (N_551,In_653,In_372);
xnor U552 (N_552,In_2926,In_846);
nor U553 (N_553,N_77,In_2565);
nor U554 (N_554,In_1055,N_209);
xor U555 (N_555,In_107,In_358);
nor U556 (N_556,N_167,In_305);
nand U557 (N_557,In_140,In_1518);
nor U558 (N_558,In_1101,In_1673);
nor U559 (N_559,In_2613,In_693);
nand U560 (N_560,In_878,In_1095);
and U561 (N_561,N_57,In_2327);
nand U562 (N_562,In_9,In_545);
and U563 (N_563,In_514,N_164);
xnor U564 (N_564,In_691,In_42);
or U565 (N_565,In_1796,In_769);
and U566 (N_566,N_251,In_1347);
nor U567 (N_567,N_99,In_1798);
or U568 (N_568,In_1724,N_202);
xor U569 (N_569,In_2608,In_978);
nand U570 (N_570,In_1195,In_496);
and U571 (N_571,In_655,In_2801);
xnor U572 (N_572,In_2814,In_1896);
nand U573 (N_573,In_142,In_773);
xor U574 (N_574,In_122,In_1767);
and U575 (N_575,In_292,In_1138);
xnor U576 (N_576,In_1185,In_616);
or U577 (N_577,In_299,In_2528);
nor U578 (N_578,In_402,N_282);
or U579 (N_579,In_388,In_690);
xor U580 (N_580,In_221,In_2507);
nor U581 (N_581,In_1776,In_1259);
nand U582 (N_582,N_193,In_1209);
xor U583 (N_583,In_90,In_2658);
nand U584 (N_584,In_610,In_2763);
xnor U585 (N_585,In_1062,In_1939);
xor U586 (N_586,In_230,N_50);
and U587 (N_587,In_2632,In_2497);
and U588 (N_588,In_871,In_2978);
nor U589 (N_589,N_185,N_29);
nor U590 (N_590,In_2254,In_2721);
and U591 (N_591,In_2238,In_2726);
and U592 (N_592,N_56,N_245);
and U593 (N_593,In_823,In_1037);
or U594 (N_594,In_2470,In_83);
nor U595 (N_595,In_2672,In_885);
or U596 (N_596,In_283,In_893);
or U597 (N_597,N_71,In_1497);
xor U598 (N_598,N_203,In_2745);
nor U599 (N_599,In_2001,In_96);
nand U600 (N_600,In_888,In_701);
and U601 (N_601,N_367,In_1710);
and U602 (N_602,In_2392,In_1979);
and U603 (N_603,In_902,In_838);
or U604 (N_604,In_2258,In_957);
nor U605 (N_605,In_2889,N_436);
or U606 (N_606,In_1636,In_1058);
and U607 (N_607,In_2486,N_583);
and U608 (N_608,N_336,In_935);
xnor U609 (N_609,N_148,In_1260);
and U610 (N_610,N_159,In_1011);
nand U611 (N_611,In_2245,In_592);
xnor U612 (N_612,N_119,In_2069);
nor U613 (N_613,In_1918,In_126);
or U614 (N_614,In_2790,In_1680);
nor U615 (N_615,N_368,In_1369);
and U616 (N_616,In_732,N_491);
nor U617 (N_617,In_649,In_2426);
or U618 (N_618,In_1152,In_2302);
and U619 (N_619,In_931,In_2728);
nor U620 (N_620,In_2005,In_1572);
nand U621 (N_621,In_666,In_1361);
nand U622 (N_622,In_1742,In_2345);
nor U623 (N_623,N_88,In_1076);
nand U624 (N_624,In_2949,N_465);
nand U625 (N_625,In_1235,In_2013);
and U626 (N_626,In_2777,In_63);
nor U627 (N_627,In_1695,In_480);
or U628 (N_628,In_1378,N_410);
xor U629 (N_629,In_761,In_164);
nor U630 (N_630,In_2747,In_1364);
or U631 (N_631,In_286,N_464);
or U632 (N_632,In_1303,In_2454);
nor U633 (N_633,N_562,N_483);
nand U634 (N_634,In_1817,In_1483);
nor U635 (N_635,In_1821,In_1513);
and U636 (N_636,N_230,In_1864);
nand U637 (N_637,In_709,In_689);
nor U638 (N_638,In_921,In_2480);
nand U639 (N_639,In_295,In_48);
xnor U640 (N_640,In_1161,In_681);
nor U641 (N_641,In_1429,N_386);
or U642 (N_642,N_2,N_244);
xor U643 (N_643,N_405,In_2991);
nor U644 (N_644,In_165,In_1167);
or U645 (N_645,In_1697,In_1254);
xnor U646 (N_646,In_2787,In_1616);
nand U647 (N_647,In_781,N_369);
xnor U648 (N_648,In_765,In_2900);
or U649 (N_649,In_209,In_457);
nand U650 (N_650,In_2097,In_510);
xnor U651 (N_651,N_22,In_2683);
nor U652 (N_652,N_235,In_1738);
xor U653 (N_653,In_741,In_601);
nor U654 (N_654,In_2263,In_2306);
or U655 (N_655,In_2137,In_804);
nor U656 (N_656,In_1802,In_2684);
xnor U657 (N_657,In_832,In_2571);
nand U658 (N_658,In_1403,In_76);
and U659 (N_659,In_843,In_817);
or U660 (N_660,In_954,N_427);
xnor U661 (N_661,In_3,In_1920);
nand U662 (N_662,N_195,N_449);
xor U663 (N_663,In_341,In_2036);
xnor U664 (N_664,N_120,N_13);
nor U665 (N_665,In_2186,In_1327);
xor U666 (N_666,In_1495,In_2183);
or U667 (N_667,In_516,In_1253);
and U668 (N_668,In_2272,In_109);
and U669 (N_669,In_1650,In_2307);
or U670 (N_670,In_1339,In_1385);
nor U671 (N_671,In_2155,N_82);
or U672 (N_672,In_543,In_1393);
and U673 (N_673,In_432,In_870);
or U674 (N_674,In_728,In_2413);
or U675 (N_675,In_2649,In_1324);
xnor U676 (N_676,In_2185,N_431);
or U677 (N_677,In_494,In_364);
nor U678 (N_678,N_393,In_2879);
nand U679 (N_679,In_2035,In_2655);
nor U680 (N_680,In_2538,In_351);
nand U681 (N_681,In_2664,In_2006);
or U682 (N_682,In_167,In_325);
nor U683 (N_683,In_1835,In_2765);
nand U684 (N_684,In_1186,In_141);
and U685 (N_685,In_2994,In_2772);
or U686 (N_686,In_2543,N_74);
nor U687 (N_687,In_2693,In_2912);
and U688 (N_688,In_2964,N_274);
and U689 (N_689,In_2828,N_430);
nor U690 (N_690,In_2936,In_1416);
and U691 (N_691,In_650,In_2888);
or U692 (N_692,In_390,In_2257);
nor U693 (N_693,N_182,In_1932);
or U694 (N_694,In_245,N_128);
nor U695 (N_695,In_544,In_1929);
xor U696 (N_696,N_89,In_619);
nor U697 (N_697,In_2643,In_1559);
nor U698 (N_698,In_1957,In_2894);
nor U699 (N_699,In_2316,In_1933);
nor U700 (N_700,In_542,N_586);
nand U701 (N_701,N_42,In_2113);
xor U702 (N_702,In_2827,N_553);
nand U703 (N_703,In_2149,In_252);
nor U704 (N_704,In_1143,In_884);
xnor U705 (N_705,In_426,In_2972);
and U706 (N_706,N_515,N_523);
nand U707 (N_707,In_1065,In_518);
nor U708 (N_708,N_100,N_441);
and U709 (N_709,In_381,In_2680);
nand U710 (N_710,In_2811,In_2210);
nor U711 (N_711,In_2984,In_784);
nand U712 (N_712,In_561,In_2193);
or U713 (N_713,In_872,N_191);
nor U714 (N_714,N_419,In_2277);
nand U715 (N_715,In_2882,In_1759);
xnor U716 (N_716,In_1153,In_1587);
nor U717 (N_717,N_420,In_1678);
and U718 (N_718,In_216,In_1583);
or U719 (N_719,In_57,In_392);
and U720 (N_720,In_2181,In_1514);
xnor U721 (N_721,In_2055,In_1134);
and U722 (N_722,In_2610,In_1027);
or U723 (N_723,N_328,In_1846);
nor U724 (N_724,In_509,In_1512);
nor U725 (N_725,In_2646,N_439);
xor U726 (N_726,In_2089,In_1411);
and U727 (N_727,In_910,In_2438);
nand U728 (N_728,In_214,N_536);
or U729 (N_729,In_1376,In_2233);
nor U730 (N_730,N_49,N_26);
xnor U731 (N_731,In_705,In_2544);
xnor U732 (N_732,N_149,In_58);
xor U733 (N_733,In_2150,N_37);
nor U734 (N_734,In_1340,In_1010);
nand U735 (N_735,N_131,In_484);
or U736 (N_736,In_1417,In_1838);
xor U737 (N_737,In_2533,In_2592);
and U738 (N_738,In_2696,In_2732);
xnor U739 (N_739,In_272,In_797);
nor U740 (N_740,N_301,N_294);
nor U741 (N_741,In_2875,In_1245);
or U742 (N_742,In_982,In_520);
nand U743 (N_743,In_1837,N_444);
and U744 (N_744,In_1726,In_2913);
and U745 (N_745,N_366,In_1959);
nand U746 (N_746,In_1169,N_236);
or U747 (N_747,N_217,In_378);
and U748 (N_748,In_2160,N_335);
xor U749 (N_749,In_1131,In_1414);
xnor U750 (N_750,In_273,In_315);
and U751 (N_751,In_2053,N_319);
and U752 (N_752,In_2051,In_2881);
xor U753 (N_753,In_811,N_118);
nand U754 (N_754,In_1030,In_1938);
or U755 (N_755,In_1409,In_1535);
nor U756 (N_756,N_363,In_1868);
nand U757 (N_757,In_669,In_148);
or U758 (N_758,In_1618,In_1857);
nand U759 (N_759,N_522,N_473);
nor U760 (N_760,In_233,N_349);
nor U761 (N_761,In_1706,In_1548);
nand U762 (N_762,In_2479,In_1292);
or U763 (N_763,In_948,In_4);
or U764 (N_764,In_2108,In_967);
or U765 (N_765,In_1643,N_205);
or U766 (N_766,N_6,In_2920);
nand U767 (N_767,N_332,N_227);
and U768 (N_768,In_974,In_333);
or U769 (N_769,In_1775,In_371);
xor U770 (N_770,In_1983,In_2367);
or U771 (N_771,In_1479,N_138);
nor U772 (N_772,In_1880,In_439);
nor U773 (N_773,In_414,In_409);
and U774 (N_774,In_1944,N_253);
nor U775 (N_775,N_102,In_35);
nand U776 (N_776,In_2301,N_457);
and U777 (N_777,N_355,In_2584);
and U778 (N_778,In_1118,In_755);
nand U779 (N_779,In_2841,In_93);
or U780 (N_780,In_614,In_2558);
and U781 (N_781,N_505,N_141);
or U782 (N_782,In_2873,In_2213);
nor U783 (N_783,In_612,In_229);
nand U784 (N_784,In_2839,N_287);
nor U785 (N_785,In_323,In_1457);
xnor U786 (N_786,N_423,In_1144);
and U787 (N_787,In_559,In_87);
or U788 (N_788,In_602,In_777);
or U789 (N_789,N_275,In_836);
or U790 (N_790,In_707,In_991);
xor U791 (N_791,N_145,In_21);
and U792 (N_792,N_198,In_2609);
and U793 (N_793,In_1050,In_2506);
or U794 (N_794,N_105,In_2358);
and U795 (N_795,In_1547,In_281);
nor U796 (N_796,In_2329,In_1867);
and U797 (N_797,In_1725,N_576);
or U798 (N_798,In_2505,In_1648);
nor U799 (N_799,In_1924,In_306);
nor U800 (N_800,N_378,In_2865);
and U801 (N_801,N_259,N_526);
and U802 (N_802,N_146,In_1212);
and U803 (N_803,In_782,In_2461);
or U804 (N_804,In_1155,In_919);
and U805 (N_805,In_2553,N_316);
and U806 (N_806,In_1622,In_1844);
nand U807 (N_807,N_79,In_2315);
or U808 (N_808,N_547,In_521);
nor U809 (N_809,In_1574,In_1222);
or U810 (N_810,In_1370,N_474);
nor U811 (N_811,In_1132,In_2414);
nor U812 (N_812,In_423,In_2589);
nand U813 (N_813,In_2826,N_162);
and U814 (N_814,In_900,In_2954);
nor U815 (N_815,In_88,In_2910);
or U816 (N_816,In_2652,N_407);
or U817 (N_817,In_1926,In_2402);
and U818 (N_818,In_193,In_1121);
nor U819 (N_819,N_411,N_511);
or U820 (N_820,In_1449,In_1556);
nor U821 (N_821,In_1375,In_298);
xnor U822 (N_822,In_2295,In_1897);
nand U823 (N_823,In_427,N_598);
xnor U824 (N_824,In_353,In_89);
or U825 (N_825,N_399,In_2931);
xnor U826 (N_826,In_2244,In_1473);
xor U827 (N_827,In_2130,N_197);
or U828 (N_828,In_607,N_309);
and U829 (N_829,In_588,In_1797);
nand U830 (N_830,N_454,N_95);
or U831 (N_831,In_1266,In_1288);
or U832 (N_832,In_1328,In_124);
nand U833 (N_833,In_529,In_2191);
nand U834 (N_834,In_399,In_620);
nor U835 (N_835,In_1089,N_75);
nor U836 (N_836,In_1653,In_1981);
nor U837 (N_837,In_1009,N_3);
xnor U838 (N_838,In_1090,In_1684);
nand U839 (N_839,In_1811,In_908);
nor U840 (N_840,In_1782,N_546);
xor U841 (N_841,In_1670,In_1654);
or U842 (N_842,In_1130,N_155);
and U843 (N_843,N_475,In_2527);
nand U844 (N_844,In_1803,N_170);
nor U845 (N_845,In_32,In_1520);
or U846 (N_846,N_460,N_5);
nand U847 (N_847,N_540,In_2421);
nand U848 (N_848,N_337,In_1645);
nor U849 (N_849,In_937,N_161);
and U850 (N_850,In_2009,N_276);
xor U851 (N_851,In_2341,In_61);
and U852 (N_852,In_541,In_2028);
or U853 (N_853,In_889,N_532);
nor U854 (N_854,N_525,In_2087);
or U855 (N_855,In_1440,In_802);
nor U856 (N_856,In_2725,In_2344);
nor U857 (N_857,In_2134,N_516);
and U858 (N_858,In_1494,N_17);
xnor U859 (N_859,N_318,In_2520);
nor U860 (N_860,In_436,N_451);
xor U861 (N_861,In_1941,In_493);
nand U862 (N_862,In_261,In_246);
and U863 (N_863,N_187,In_708);
or U864 (N_864,N_72,N_171);
nand U865 (N_865,In_2496,In_1191);
and U866 (N_866,In_790,In_2321);
xor U867 (N_867,In_577,N_271);
nor U868 (N_868,In_2342,In_442);
xor U869 (N_869,In_660,In_1395);
nor U870 (N_870,In_471,In_507);
and U871 (N_871,In_2433,In_2262);
nand U872 (N_872,N_283,N_497);
and U873 (N_873,N_173,In_395);
or U874 (N_874,In_244,N_537);
or U875 (N_875,In_1345,In_1505);
nand U876 (N_876,N_188,In_2678);
or U877 (N_877,In_680,In_1355);
xor U878 (N_878,In_2465,In_1091);
xnor U879 (N_879,In_1220,In_308);
xor U880 (N_880,In_2542,N_39);
xor U881 (N_881,N_458,In_1871);
or U882 (N_882,In_28,In_2862);
xor U883 (N_883,In_2115,N_500);
xnor U884 (N_884,In_916,In_1704);
and U885 (N_885,In_56,In_1808);
or U886 (N_886,In_752,N_248);
xnor U887 (N_887,N_228,In_1985);
nand U888 (N_888,In_1987,N_356);
nor U889 (N_889,In_1425,In_1326);
nor U890 (N_890,In_973,N_226);
nor U891 (N_891,N_517,In_2850);
nor U892 (N_892,N_16,In_166);
and U893 (N_893,In_1135,In_379);
xor U894 (N_894,N_108,In_2526);
nor U895 (N_895,In_65,In_997);
nand U896 (N_896,In_2153,In_40);
or U897 (N_897,In_2247,In_2919);
nand U898 (N_898,In_2871,In_687);
and U899 (N_899,In_2780,In_1150);
or U900 (N_900,In_567,In_133);
or U901 (N_901,N_385,In_1569);
nand U902 (N_902,N_204,N_813);
nor U903 (N_903,In_382,In_419);
nand U904 (N_904,In_1566,N_704);
xnor U905 (N_905,In_1870,In_478);
xor U906 (N_906,N_296,In_2283);
nor U907 (N_907,N_482,N_640);
and U908 (N_908,In_2956,N_615);
xnor U909 (N_909,N_738,N_467);
nor U910 (N_910,In_1082,In_1915);
nand U911 (N_911,In_186,In_1423);
nand U912 (N_912,In_316,In_2886);
nand U913 (N_913,In_2799,In_881);
nor U914 (N_914,N_117,N_48);
nor U915 (N_915,In_2226,In_679);
or U916 (N_916,N_34,N_842);
or U917 (N_917,In_1628,In_438);
and U918 (N_918,In_2076,N_331);
nand U919 (N_919,In_1581,N_776);
or U920 (N_920,N_852,N_673);
nand U921 (N_921,In_1605,In_205);
and U922 (N_922,N_160,N_792);
and U923 (N_923,In_177,N_521);
xor U924 (N_924,N_163,In_1671);
nor U925 (N_925,In_1890,In_203);
and U926 (N_926,In_481,In_1586);
nor U927 (N_927,N_642,In_2174);
xnor U928 (N_928,N_503,N_299);
or U929 (N_929,In_2789,In_1115);
or U930 (N_930,In_2042,In_377);
or U931 (N_931,N_742,N_866);
nand U932 (N_932,In_2122,In_2038);
and U933 (N_933,N_389,In_2118);
nor U934 (N_934,In_1522,N_8);
nand U935 (N_935,N_424,In_2352);
xor U936 (N_936,In_2626,In_1794);
and U937 (N_937,N_604,In_2810);
nand U938 (N_938,N_780,In_1317);
and U939 (N_939,N_748,In_1825);
or U940 (N_940,N_555,N_343);
nand U941 (N_941,In_2939,N_19);
xnor U942 (N_942,N_179,In_1901);
nor U943 (N_943,In_1334,In_866);
and U944 (N_944,In_184,In_2430);
and U945 (N_945,N_416,In_2158);
nand U946 (N_946,In_1431,In_2466);
or U947 (N_947,In_1492,In_1954);
nor U948 (N_948,In_263,In_2987);
nor U949 (N_949,N_87,N_543);
nand U950 (N_950,In_45,In_2947);
or U951 (N_951,In_863,In_1275);
and U952 (N_952,N_345,In_81);
nand U953 (N_953,In_2969,In_2820);
nor U954 (N_954,In_1359,In_350);
and U955 (N_955,In_750,In_1626);
xor U956 (N_956,In_111,N_443);
nand U957 (N_957,In_466,N_626);
and U958 (N_958,In_2192,N_285);
nor U959 (N_959,N_361,N_797);
nor U960 (N_960,N_800,In_758);
xnor U961 (N_961,In_2965,In_2846);
or U962 (N_962,In_2270,N_189);
xnor U963 (N_963,In_2052,In_1568);
nor U964 (N_964,In_2498,In_1922);
and U965 (N_965,In_2462,In_2151);
or U966 (N_966,N_339,N_853);
nor U967 (N_967,N_874,In_1657);
and U968 (N_968,In_2501,In_1795);
or U969 (N_969,N_708,In_1244);
xnor U970 (N_970,In_2136,In_1993);
or U971 (N_971,N_840,In_416);
and U972 (N_972,N_552,In_1060);
or U973 (N_973,In_366,In_2356);
nor U974 (N_974,In_1067,N_735);
xnor U975 (N_975,In_2570,In_1335);
nand U976 (N_976,In_2475,N_395);
nor U977 (N_977,N_781,In_922);
xnor U978 (N_978,In_1059,In_400);
xnor U979 (N_979,N_607,N_476);
or U980 (N_980,N_254,N_354);
nor U981 (N_981,In_1213,In_2681);
and U982 (N_982,In_340,In_2101);
or U983 (N_983,In_2490,In_918);
or U984 (N_984,In_1280,In_959);
nand U985 (N_985,N_861,N_502);
nor U986 (N_986,In_331,N_855);
nor U987 (N_987,In_2331,In_2840);
xor U988 (N_988,In_1075,N_712);
xor U989 (N_989,In_259,In_2377);
and U990 (N_990,N_825,In_2739);
nor U991 (N_991,N_684,In_1623);
nand U992 (N_992,In_276,In_115);
or U993 (N_993,In_2003,In_1974);
or U994 (N_994,In_1940,In_1872);
xnor U995 (N_995,In_1772,In_2769);
xnor U996 (N_996,In_473,In_652);
xor U997 (N_997,In_1745,In_2317);
or U998 (N_998,In_995,In_1487);
nor U999 (N_999,In_1723,N_851);
nor U1000 (N_1000,N_756,In_2116);
nor U1001 (N_1001,In_1996,In_2123);
nand U1002 (N_1002,In_1604,In_1638);
nor U1003 (N_1003,In_2403,In_1851);
and U1004 (N_1004,N_843,In_907);
nor U1005 (N_1005,In_2405,In_1606);
nor U1006 (N_1006,N_849,In_1019);
xor U1007 (N_1007,In_1562,In_2339);
nor U1008 (N_1008,In_2615,N_584);
and U1009 (N_1009,In_2742,In_1972);
xor U1010 (N_1010,In_389,N_252);
and U1011 (N_1011,In_2337,In_1927);
xor U1012 (N_1012,In_321,In_27);
xor U1013 (N_1013,In_1635,In_2260);
nand U1014 (N_1014,In_1397,N_667);
nand U1015 (N_1015,N_893,In_839);
or U1016 (N_1016,In_1410,N_556);
and U1017 (N_1017,N_382,In_2148);
xor U1018 (N_1018,N_365,In_1389);
nor U1019 (N_1019,In_290,N_638);
and U1020 (N_1020,In_1148,In_2971);
xnor U1021 (N_1021,N_388,N_750);
and U1022 (N_1022,N_621,In_2338);
xnor U1023 (N_1023,In_1163,In_630);
nor U1024 (N_1024,N_359,N_670);
or U1025 (N_1025,In_1842,In_2229);
nor U1026 (N_1026,In_930,N_600);
nor U1027 (N_1027,N_716,N_741);
nand U1028 (N_1028,In_1448,In_1348);
and U1029 (N_1029,In_2063,In_2605);
or U1030 (N_1030,In_525,In_2408);
and U1031 (N_1031,In_1391,N_213);
nor U1032 (N_1032,In_672,N_728);
and U1033 (N_1033,N_494,In_667);
nor U1034 (N_1034,In_1715,N_323);
and U1035 (N_1035,N_325,N_406);
or U1036 (N_1036,In_716,In_1173);
and U1037 (N_1037,In_2441,N_577);
nor U1038 (N_1038,N_211,In_477);
nor U1039 (N_1039,In_1530,In_269);
xor U1040 (N_1040,In_1708,In_780);
xnor U1041 (N_1041,In_746,In_2395);
or U1042 (N_1042,In_1125,In_2929);
xor U1043 (N_1043,In_1002,In_1525);
nand U1044 (N_1044,In_1792,N_709);
nor U1045 (N_1045,In_2689,In_172);
nand U1046 (N_1046,N_625,In_1858);
nand U1047 (N_1047,In_82,In_1402);
and U1048 (N_1048,In_603,In_2710);
or U1049 (N_1049,In_853,In_1300);
or U1050 (N_1050,N_46,N_718);
nor U1051 (N_1051,N_223,In_1181);
and U1052 (N_1052,In_664,In_2654);
xor U1053 (N_1053,In_22,In_2324);
or U1054 (N_1054,In_925,In_850);
nor U1055 (N_1055,In_1675,In_1711);
nor U1056 (N_1056,In_2443,In_2167);
and U1057 (N_1057,N_663,In_2293);
nand U1058 (N_1058,N_890,In_1078);
xnor U1059 (N_1059,In_2977,In_2178);
nor U1060 (N_1060,In_123,In_2056);
xnor U1061 (N_1061,In_613,In_2370);
nor U1062 (N_1062,In_2065,In_334);
nor U1063 (N_1063,In_34,N_400);
xnor U1064 (N_1064,N_769,In_1499);
or U1065 (N_1065,In_1952,N_9);
or U1066 (N_1066,In_2446,In_2154);
nor U1067 (N_1067,N_429,In_2937);
nor U1068 (N_1068,N_317,In_1905);
nand U1069 (N_1069,In_726,In_2835);
or U1070 (N_1070,In_2843,In_1434);
nand U1071 (N_1071,N_533,N_493);
xnor U1072 (N_1072,N_143,N_448);
nand U1073 (N_1073,In_130,In_834);
nand U1074 (N_1074,In_2493,In_562);
nor U1075 (N_1075,In_2289,In_938);
nor U1076 (N_1076,N_498,N_779);
xor U1077 (N_1077,In_2682,In_1194);
or U1078 (N_1078,In_2172,N_97);
or U1079 (N_1079,In_1398,In_600);
nor U1080 (N_1080,In_1087,In_1436);
nand U1081 (N_1081,N_480,In_2671);
xor U1082 (N_1082,In_1986,N_326);
nand U1083 (N_1083,N_619,In_2274);
nor U1084 (N_1084,In_2752,N_81);
nor U1085 (N_1085,N_194,In_723);
nor U1086 (N_1086,N_578,In_2415);
and U1087 (N_1087,In_1158,N_624);
xnor U1088 (N_1088,In_2304,In_1192);
nand U1089 (N_1089,In_2407,In_799);
nor U1090 (N_1090,In_2215,In_2644);
nand U1091 (N_1091,In_899,In_285);
or U1092 (N_1092,In_275,In_136);
nand U1093 (N_1093,In_1889,In_2785);
nand U1094 (N_1094,In_1136,N_798);
nor U1095 (N_1095,N_788,N_821);
and U1096 (N_1096,N_320,N_871);
nand U1097 (N_1097,In_194,N_846);
nand U1098 (N_1098,In_1133,In_1261);
xnor U1099 (N_1099,N_696,N_807);
xnor U1100 (N_1100,In_1329,In_2399);
and U1101 (N_1101,In_2720,In_2376);
nor U1102 (N_1102,N_127,In_1063);
xnor U1103 (N_1103,N_743,N_381);
nand U1104 (N_1104,N_752,N_746);
and U1105 (N_1105,N_495,In_2271);
and U1106 (N_1106,N_338,In_2596);
xnor U1107 (N_1107,In_1374,N_815);
and U1108 (N_1108,N_487,In_892);
or U1109 (N_1109,In_1667,In_1836);
nor U1110 (N_1110,In_1188,N_803);
and U1111 (N_1111,In_430,N_315);
or U1112 (N_1112,In_1490,In_2668);
nor U1113 (N_1113,N_805,In_776);
nand U1114 (N_1114,N_308,In_1656);
xor U1115 (N_1115,In_2107,In_685);
nor U1116 (N_1116,N_658,In_1696);
nor U1117 (N_1117,In_2662,In_2665);
and U1118 (N_1118,N_342,In_1362);
nand U1119 (N_1119,In_1474,In_1689);
nor U1120 (N_1120,In_2741,In_2102);
xor U1121 (N_1121,In_1552,In_1528);
or U1122 (N_1122,In_670,In_1461);
and U1123 (N_1123,In_2431,N_892);
and U1124 (N_1124,N_875,N_297);
or U1125 (N_1125,N_885,N_809);
and U1126 (N_1126,N_422,N_888);
nor U1127 (N_1127,N_11,N_758);
xor U1128 (N_1128,In_642,In_1992);
nand U1129 (N_1129,In_1966,In_2079);
nand U1130 (N_1130,N_588,In_971);
nor U1131 (N_1131,In_1363,In_1228);
xor U1132 (N_1132,In_527,In_538);
and U1133 (N_1133,N_876,In_1506);
or U1134 (N_1134,In_345,In_1869);
and U1135 (N_1135,In_2753,In_1353);
and U1136 (N_1136,In_1751,N_836);
and U1137 (N_1137,N_585,In_2796);
or U1138 (N_1138,In_556,In_2853);
nor U1139 (N_1139,In_876,N_341);
nand U1140 (N_1140,In_2128,N_262);
and U1141 (N_1141,N_304,N_174);
xnor U1142 (N_1142,In_2230,In_983);
nand U1143 (N_1143,N_679,In_412);
nor U1144 (N_1144,In_1214,In_1480);
and U1145 (N_1145,N_864,In_1311);
and U1146 (N_1146,In_2382,In_1652);
nor U1147 (N_1147,In_472,In_2907);
nand U1148 (N_1148,N_513,In_1103);
nor U1149 (N_1149,N_707,In_1346);
or U1150 (N_1150,In_984,N_740);
nand U1151 (N_1151,In_2265,In_2510);
nor U1152 (N_1152,In_2844,N_496);
and U1153 (N_1153,N_333,In_998);
or U1154 (N_1154,N_862,In_2824);
nor U1155 (N_1155,In_105,In_1649);
or U1156 (N_1156,In_1450,In_2588);
nor U1157 (N_1157,In_2129,In_2026);
xor U1158 (N_1158,N_353,In_2364);
nand U1159 (N_1159,In_1945,In_2313);
or U1160 (N_1160,N_644,In_1331);
and U1161 (N_1161,In_207,N_514);
nand U1162 (N_1162,In_1624,In_955);
and U1163 (N_1163,In_2417,N_33);
nor U1164 (N_1164,In_615,N_247);
nor U1165 (N_1165,In_2695,N_877);
and U1166 (N_1166,N_883,In_2731);
or U1167 (N_1167,In_977,N_639);
nand U1168 (N_1168,N_897,N_590);
nand U1169 (N_1169,In_605,In_2237);
nand U1170 (N_1170,N_18,In_2495);
or U1171 (N_1171,N_249,In_1352);
and U1172 (N_1172,In_1283,In_2690);
xnor U1173 (N_1173,In_714,N_828);
and U1174 (N_1174,In_2722,In_338);
xor U1175 (N_1175,In_862,N_373);
or U1176 (N_1176,In_1052,In_972);
nor U1177 (N_1177,In_2248,N_848);
nand U1178 (N_1178,N_782,In_2359);
and U1179 (N_1179,In_712,In_492);
or U1180 (N_1180,N_668,N_802);
nand U1181 (N_1181,In_2121,In_474);
or U1182 (N_1182,N_518,N_647);
xor U1183 (N_1183,N_865,In_1551);
nand U1184 (N_1184,In_424,In_240);
and U1185 (N_1185,N_603,In_936);
or U1186 (N_1186,In_236,In_2800);
xor U1187 (N_1187,In_2182,N_857);
nand U1188 (N_1188,In_1219,In_920);
or U1189 (N_1189,In_14,In_12);
or U1190 (N_1190,N_41,In_1819);
nand U1191 (N_1191,N_806,In_2548);
or U1192 (N_1192,In_1576,In_546);
or U1193 (N_1193,In_2418,N_477);
xor U1194 (N_1194,N_589,N_814);
xor U1195 (N_1195,N_440,In_2404);
xor U1196 (N_1196,In_1380,In_2767);
or U1197 (N_1197,In_152,In_1127);
nand U1198 (N_1198,In_46,In_526);
or U1199 (N_1199,N_452,N_112);
nor U1200 (N_1200,N_535,In_753);
xnor U1201 (N_1201,N_824,N_947);
and U1202 (N_1202,N_545,N_433);
or U1203 (N_1203,In_52,In_231);
xor U1204 (N_1204,In_2004,In_1977);
xnor U1205 (N_1205,In_314,N_269);
or U1206 (N_1206,In_2104,In_1304);
or U1207 (N_1207,N_456,N_1128);
nand U1208 (N_1208,N_450,In_2774);
or U1209 (N_1209,N_1166,In_2587);
nor U1210 (N_1210,N_425,In_1541);
and U1211 (N_1211,N_1009,N_933);
nor U1212 (N_1212,In_2860,N_488);
or U1213 (N_1213,In_369,In_789);
or U1214 (N_1214,In_2023,In_2792);
nor U1215 (N_1215,In_1515,In_2968);
and U1216 (N_1216,In_162,In_2251);
nor U1217 (N_1217,N_478,In_2473);
nor U1218 (N_1218,N_201,In_1165);
xor U1219 (N_1219,In_965,N_506);
nor U1220 (N_1220,In_2711,N_371);
nand U1221 (N_1221,In_2385,In_929);
and U1222 (N_1222,N_157,In_2757);
nor U1223 (N_1223,N_554,In_2224);
xnor U1224 (N_1224,N_551,N_786);
nor U1225 (N_1225,N_565,In_2743);
xor U1226 (N_1226,In_2556,In_2333);
nor U1227 (N_1227,In_1546,N_1030);
and U1228 (N_1228,N_765,In_598);
or U1229 (N_1229,N_688,N_1151);
nor U1230 (N_1230,In_1295,N_899);
and U1231 (N_1231,In_2078,N_1055);
nand U1232 (N_1232,N_1104,N_956);
nand U1233 (N_1233,In_2564,In_2942);
and U1234 (N_1234,N_692,In_2855);
and U1235 (N_1235,In_2159,In_1860);
nand U1236 (N_1236,In_1045,In_19);
nand U1237 (N_1237,In_810,In_1033);
nand U1238 (N_1238,In_2365,N_1065);
xor U1239 (N_1239,In_2518,N_109);
nor U1240 (N_1240,N_992,In_2708);
nor U1241 (N_1241,N_946,N_1035);
nor U1242 (N_1242,In_2143,N_1011);
nor U1243 (N_1243,In_2569,In_112);
nor U1244 (N_1244,In_909,N_437);
and U1245 (N_1245,In_808,In_1320);
nor U1246 (N_1246,In_2805,In_441);
or U1247 (N_1247,In_1092,In_2232);
nand U1248 (N_1248,N_1187,In_831);
nor U1249 (N_1249,N_116,N_438);
and U1250 (N_1250,In_1968,In_2072);
xnor U1251 (N_1251,In_1122,In_1875);
and U1252 (N_1252,In_1233,In_1641);
nor U1253 (N_1253,N_620,N_988);
or U1254 (N_1254,In_1036,N_1186);
or U1255 (N_1255,N_384,N_678);
nor U1256 (N_1256,N_937,In_1307);
nor U1257 (N_1257,N_605,In_1895);
nand U1258 (N_1258,In_2241,N_1080);
nor U1259 (N_1259,In_2759,In_2593);
nor U1260 (N_1260,In_404,N_730);
nand U1261 (N_1261,N_306,N_531);
nor U1262 (N_1262,In_513,In_2440);
and U1263 (N_1263,In_1430,N_945);
and U1264 (N_1264,N_1013,N_61);
and U1265 (N_1265,In_116,In_2614);
or U1266 (N_1266,N_1044,In_2276);
nand U1267 (N_1267,In_1028,N_169);
or U1268 (N_1268,N_878,N_510);
and U1269 (N_1269,In_324,N_622);
xnor U1270 (N_1270,In_2057,In_958);
xor U1271 (N_1271,In_2373,In_1223);
or U1272 (N_1272,In_2677,N_950);
xnor U1273 (N_1273,In_1469,In_1031);
and U1274 (N_1274,In_960,In_2083);
nor U1275 (N_1275,In_312,N_442);
nor U1276 (N_1276,In_857,In_2194);
nor U1277 (N_1277,N_557,In_289);
nor U1278 (N_1278,N_997,N_392);
nand U1279 (N_1279,N_426,In_2029);
and U1280 (N_1280,In_2590,N_62);
and U1281 (N_1281,In_1061,N_1109);
or U1282 (N_1282,N_402,N_869);
xnor U1283 (N_1283,In_2941,In_2416);
nand U1284 (N_1284,N_1163,In_2716);
nor U1285 (N_1285,In_2583,N_953);
nor U1286 (N_1286,N_760,In_1203);
nand U1287 (N_1287,In_2114,N_766);
nand U1288 (N_1288,In_1632,N_186);
xor U1289 (N_1289,N_327,N_759);
nand U1290 (N_1290,N_1198,N_770);
nand U1291 (N_1291,In_74,In_1741);
or U1292 (N_1292,In_2988,In_890);
nand U1293 (N_1293,N_726,In_2256);
nand U1294 (N_1294,N_137,N_689);
and U1295 (N_1295,N_1034,N_15);
nor U1296 (N_1296,In_2960,N_1020);
xnor U1297 (N_1297,In_1784,In_1593);
xor U1298 (N_1298,In_85,In_897);
nand U1299 (N_1299,In_2918,N_686);
and U1300 (N_1300,In_1225,In_793);
nor U1301 (N_1301,In_95,N_35);
nand U1302 (N_1302,N_935,In_1936);
or U1303 (N_1303,N_1130,In_277);
nor U1304 (N_1304,N_73,N_199);
or U1305 (N_1305,N_1063,In_1306);
or U1306 (N_1306,In_979,In_1863);
or U1307 (N_1307,In_128,N_314);
nand U1308 (N_1308,In_97,In_2362);
nand U1309 (N_1309,N_913,In_408);
nor U1310 (N_1310,N_550,N_1098);
nor U1311 (N_1311,In_1707,In_1862);
xnor U1312 (N_1312,N_541,In_1747);
and U1313 (N_1313,In_1029,In_903);
nor U1314 (N_1314,In_1533,In_2504);
and U1315 (N_1315,N_1108,In_158);
nor U1316 (N_1316,N_206,N_867);
nor U1317 (N_1317,In_190,N_1038);
xnor U1318 (N_1318,N_1070,N_713);
nor U1319 (N_1319,In_2406,N_1018);
nand U1320 (N_1320,In_354,N_1091);
nand U1321 (N_1321,N_573,In_628);
nor U1322 (N_1322,N_508,N_970);
xnor U1323 (N_1323,In_1452,In_851);
or U1324 (N_1324,N_396,In_2896);
or U1325 (N_1325,N_858,N_1092);
nor U1326 (N_1326,N_459,In_2340);
xor U1327 (N_1327,In_1557,In_2112);
nor U1328 (N_1328,In_2733,In_2798);
and U1329 (N_1329,N_542,In_437);
xor U1330 (N_1330,N_596,N_91);
and U1331 (N_1331,N_1115,N_86);
nor U1332 (N_1332,In_176,N_1062);
nand U1333 (N_1333,N_1014,In_1094);
and U1334 (N_1334,In_2560,N_894);
nand U1335 (N_1335,N_1029,In_288);
nand U1336 (N_1336,In_1172,In_238);
and U1337 (N_1337,N_221,N_499);
and U1338 (N_1338,N_1160,In_748);
nand U1339 (N_1339,In_1793,N_654);
xor U1340 (N_1340,N_10,N_978);
nor U1341 (N_1341,N_492,In_2822);
nor U1342 (N_1342,In_1839,N_106);
and U1343 (N_1343,N_446,In_2764);
nor U1344 (N_1344,N_957,In_1570);
nor U1345 (N_1345,N_614,In_2205);
xnor U1346 (N_1346,N_969,N_561);
nor U1347 (N_1347,In_2165,In_842);
or U1348 (N_1348,In_222,N_761);
nor U1349 (N_1349,N_606,N_613);
xor U1350 (N_1350,N_808,In_1070);
and U1351 (N_1351,N_826,N_548);
or U1352 (N_1352,N_466,In_980);
or U1353 (N_1353,N_697,N_699);
or U1354 (N_1354,In_1679,N_237);
or U1355 (N_1355,In_1407,In_1919);
or U1356 (N_1356,N_1019,In_1856);
nor U1357 (N_1357,N_1016,In_638);
nor U1358 (N_1358,In_1773,In_49);
and U1359 (N_1359,N_911,In_363);
nand U1360 (N_1360,In_2923,N_773);
and U1361 (N_1361,In_944,N_616);
nor U1362 (N_1362,N_1061,N_471);
nand U1363 (N_1363,In_2892,N_463);
nor U1364 (N_1364,In_2539,In_11);
xnor U1365 (N_1365,N_1140,In_1799);
or U1366 (N_1366,In_2955,In_359);
nand U1367 (N_1367,N_787,N_632);
nor U1368 (N_1368,N_51,In_2948);
xor U1369 (N_1369,In_1879,In_2779);
and U1370 (N_1370,N_819,N_421);
and U1371 (N_1371,N_717,N_582);
xnor U1372 (N_1372,In_587,N_990);
nand U1373 (N_1373,N_351,N_949);
nor U1374 (N_1374,In_2895,In_2566);
xnor U1375 (N_1375,In_2930,In_2094);
nand U1376 (N_1376,N_330,In_611);
and U1377 (N_1377,N_731,N_1004);
nand U1378 (N_1378,In_397,N_1001);
and U1379 (N_1379,In_768,In_703);
or U1380 (N_1380,N_963,N_268);
xnor U1381 (N_1381,In_227,In_1960);
and U1382 (N_1382,In_2950,In_912);
nand U1383 (N_1383,N_468,In_987);
and U1384 (N_1384,N_307,N_241);
xor U1385 (N_1385,In_29,In_1343);
or U1386 (N_1386,In_1106,N_922);
nand U1387 (N_1387,In_147,In_968);
nand U1388 (N_1388,N_900,N_1076);
nand U1389 (N_1389,In_1874,In_100);
and U1390 (N_1390,In_1224,In_1883);
nand U1391 (N_1391,In_2660,In_2374);
xnor U1392 (N_1392,In_2275,N_774);
and U1393 (N_1393,N_114,In_2602);
xnor U1394 (N_1394,In_578,N_455);
or U1395 (N_1395,N_739,In_617);
xnor U1396 (N_1396,N_733,In_2499);
nand U1397 (N_1397,In_1093,In_1204);
xor U1398 (N_1398,N_841,N_856);
and U1399 (N_1399,In_2016,N_794);
or U1400 (N_1400,In_157,N_981);
or U1401 (N_1401,In_2597,In_2435);
nor U1402 (N_1402,In_70,In_833);
and U1403 (N_1403,In_447,N_418);
nor U1404 (N_1404,In_182,In_2607);
xnor U1405 (N_1405,N_698,N_727);
and U1406 (N_1406,In_906,In_2651);
or U1407 (N_1407,In_1032,In_879);
xnor U1408 (N_1408,In_1637,N_567);
nor U1409 (N_1409,In_1406,In_2825);
or U1410 (N_1410,In_2086,In_2857);
nand U1411 (N_1411,N_1075,N_895);
nor U1412 (N_1412,In_401,N_1129);
xnor U1413 (N_1413,In_604,In_2893);
and U1414 (N_1414,N_987,In_2775);
nor U1415 (N_1415,N_835,N_334);
and U1416 (N_1416,In_1668,In_2612);
xnor U1417 (N_1417,N_1133,N_1025);
xor U1418 (N_1418,In_2033,In_1381);
nand U1419 (N_1419,In_1178,N_302);
nand U1420 (N_1420,In_734,In_2532);
or U1421 (N_1421,In_144,N_32);
xor U1422 (N_1422,In_1426,In_1764);
and U1423 (N_1423,In_2829,In_2854);
and U1424 (N_1424,In_2724,In_1342);
nand U1425 (N_1425,N_85,In_2618);
nand U1426 (N_1426,In_169,N_837);
nand U1427 (N_1427,In_2795,N_801);
nand U1428 (N_1428,In_2320,In_2169);
nand U1429 (N_1429,In_1463,In_1984);
or U1430 (N_1430,N_272,In_2536);
xor U1431 (N_1431,N_690,N_1094);
or U1432 (N_1432,In_132,In_2044);
nor U1433 (N_1433,In_939,N_1093);
nand U1434 (N_1434,N_397,N_350);
xnor U1435 (N_1435,In_1766,In_1193);
xor U1436 (N_1436,N_1107,In_2959);
or U1437 (N_1437,In_993,In_217);
and U1438 (N_1438,N_134,In_47);
or U1439 (N_1439,In_2902,N_665);
or U1440 (N_1440,In_719,N_139);
nand U1441 (N_1441,In_337,N_1138);
nand U1442 (N_1442,In_2110,In_2761);
xor U1443 (N_1443,N_358,N_597);
or U1444 (N_1444,N_693,N_156);
or U1445 (N_1445,N_995,N_1181);
or U1446 (N_1446,In_2705,N_559);
nand U1447 (N_1447,In_582,In_2870);
or U1448 (N_1448,In_659,In_695);
nor U1449 (N_1449,N_1069,N_136);
and U1450 (N_1450,In_1756,N_154);
nand U1451 (N_1451,N_1105,N_387);
nor U1452 (N_1452,In_1964,N_563);
or U1453 (N_1453,N_657,N_133);
or U1454 (N_1454,In_1523,In_1357);
nor U1455 (N_1455,In_2812,N_732);
nand U1456 (N_1456,N_67,In_336);
and U1457 (N_1457,In_1596,In_2425);
xor U1458 (N_1458,In_297,In_2601);
or U1459 (N_1459,In_1990,In_1529);
and U1460 (N_1460,N_778,N_408);
nor U1461 (N_1461,N_1189,N_312);
nor U1462 (N_1462,In_2856,In_2162);
and U1463 (N_1463,In_1686,N_172);
nor U1464 (N_1464,N_1000,In_2361);
xnor U1465 (N_1465,N_1136,N_925);
xor U1466 (N_1466,In_454,In_1114);
nand U1467 (N_1467,In_1175,N_509);
nor U1468 (N_1468,In_2712,In_1472);
xor U1469 (N_1469,In_962,In_573);
nor U1470 (N_1470,N_1089,N_687);
or U1471 (N_1471,N_231,In_2512);
nand U1472 (N_1472,In_940,In_794);
xnor U1473 (N_1473,In_1910,In_2355);
nand U1474 (N_1474,N_207,In_1595);
or U1475 (N_1475,N_882,N_347);
or U1476 (N_1476,In_1481,In_1007);
xnor U1477 (N_1477,In_786,In_2541);
xor U1478 (N_1478,N_176,In_700);
or U1479 (N_1479,N_1142,N_219);
nor U1480 (N_1480,In_1832,In_1850);
nor U1481 (N_1481,N_1100,N_1161);
or U1482 (N_1482,In_1207,N_1168);
nand U1483 (N_1483,In_1682,N_340);
nor U1484 (N_1484,N_811,In_500);
nand U1485 (N_1485,N_560,N_472);
nand U1486 (N_1486,N_352,N_705);
or U1487 (N_1487,In_1893,In_1532);
or U1488 (N_1488,N_544,In_1350);
or U1489 (N_1489,In_530,In_1753);
xnor U1490 (N_1490,N_121,N_489);
and U1491 (N_1491,N_1005,In_1521);
nor U1492 (N_1492,N_1046,In_374);
or U1493 (N_1493,In_161,N_661);
xor U1494 (N_1494,In_1778,N_1157);
nand U1495 (N_1495,In_2031,In_1356);
or U1496 (N_1496,In_2474,N_793);
xor U1497 (N_1497,In_698,N_409);
or U1498 (N_1498,In_645,N_754);
or U1499 (N_1499,In_1999,N_1068);
and U1500 (N_1500,N_901,N_831);
nor U1501 (N_1501,In_2303,In_2090);
or U1502 (N_1502,N_1274,N_646);
xor U1503 (N_1503,In_658,In_505);
and U1504 (N_1504,N_1477,In_1625);
nand U1505 (N_1505,In_917,In_606);
or U1506 (N_1506,In_367,In_511);
nand U1507 (N_1507,N_123,N_486);
and U1508 (N_1508,In_662,In_1810);
xor U1509 (N_1509,In_1419,In_2744);
xor U1510 (N_1510,N_1365,N_966);
nand U1511 (N_1511,N_1334,In_1447);
nand U1512 (N_1512,N_682,N_795);
nand U1513 (N_1513,In_883,N_1357);
nand U1514 (N_1514,N_1413,In_1592);
nand U1515 (N_1515,In_1937,In_1542);
xor U1516 (N_1516,In_2996,In_249);
nor U1517 (N_1517,N_1284,In_1651);
and U1518 (N_1518,N_1026,N_1267);
and U1519 (N_1519,N_1444,N_1301);
xor U1520 (N_1520,In_1273,N_914);
or U1521 (N_1521,N_372,N_1196);
nand U1522 (N_1522,In_1947,N_677);
or U1523 (N_1523,N_1373,N_1305);
xnor U1524 (N_1524,N_1437,N_609);
nor U1525 (N_1525,N_1340,N_1333);
and U1526 (N_1526,N_4,In_2450);
or U1527 (N_1527,N_98,N_1318);
and U1528 (N_1528,In_1073,N_144);
or U1529 (N_1529,N_1303,N_1280);
and U1530 (N_1530,N_1294,N_1469);
and U1531 (N_1531,N_1411,In_453);
or U1532 (N_1532,In_1226,N_1182);
xor U1533 (N_1533,In_1077,N_965);
or U1534 (N_1534,In_2093,In_1788);
or U1535 (N_1535,N_1229,In_23);
nor U1536 (N_1536,In_629,In_185);
nand U1537 (N_1537,N_7,N_790);
xnor U1538 (N_1538,In_1814,In_1702);
nand U1539 (N_1539,N_1310,In_2018);
or U1540 (N_1540,N_1353,In_1829);
nand U1541 (N_1541,N_1470,In_2718);
xnor U1542 (N_1542,In_69,N_374);
xnor U1543 (N_1543,N_1453,In_1100);
and U1544 (N_1544,In_1806,N_1165);
nand U1545 (N_1545,In_1120,In_2685);
nor U1546 (N_1546,N_655,N_1306);
nand U1547 (N_1547,In_1611,In_1246);
nor U1548 (N_1548,N_1430,In_228);
or U1549 (N_1549,N_1400,In_2550);
nor U1550 (N_1550,N_192,In_265);
xor U1551 (N_1551,In_445,N_1224);
nand U1552 (N_1552,In_232,N_1380);
or U1553 (N_1553,In_429,In_2309);
xnor U1554 (N_1554,N_1364,In_2898);
and U1555 (N_1555,N_1090,N_1427);
nor U1556 (N_1556,In_2323,N_1204);
nand U1557 (N_1557,In_26,In_827);
nand U1558 (N_1558,N_1499,In_66);
nor U1559 (N_1559,N_1296,N_1483);
xnor U1560 (N_1560,N_823,In_1571);
xor U1561 (N_1561,N_664,In_1705);
or U1562 (N_1562,N_1304,In_1079);
nor U1563 (N_1563,In_2434,In_415);
or U1564 (N_1564,N_1436,N_1227);
nor U1565 (N_1565,In_2823,In_2071);
nor U1566 (N_1566,N_1338,N_1386);
nand U1567 (N_1567,N_1325,In_420);
and U1568 (N_1568,N_1327,In_180);
nor U1569 (N_1569,N_744,In_1291);
and U1570 (N_1570,N_1007,In_2980);
xor U1571 (N_1571,N_324,N_972);
xnor U1572 (N_1572,In_2386,N_612);
or U1573 (N_1573,In_479,In_17);
and U1574 (N_1574,N_1111,N_1145);
or U1575 (N_1575,N_1010,N_376);
nor U1576 (N_1576,N_1118,N_681);
or U1577 (N_1577,N_940,N_1258);
or U1578 (N_1578,N_200,N_1257);
nand U1579 (N_1579,In_503,In_1021);
nor U1580 (N_1580,N_23,In_2928);
and U1581 (N_1581,N_1336,N_968);
or U1582 (N_1582,N_1067,In_1779);
nand U1583 (N_1583,In_1322,In_1845);
or U1584 (N_1584,In_2738,In_2227);
nand U1585 (N_1585,N_783,N_608);
and U1586 (N_1586,N_630,In_1057);
nand U1587 (N_1587,In_1973,In_296);
nor U1588 (N_1588,In_868,N_539);
nor U1589 (N_1589,N_1322,N_1113);
xnor U1590 (N_1590,N_1086,N_311);
nand U1591 (N_1591,In_1038,In_678);
nor U1592 (N_1592,In_197,N_364);
nor U1593 (N_1593,N_1099,In_2750);
nor U1594 (N_1594,In_2472,N_971);
xor U1595 (N_1595,N_1399,In_241);
xnor U1596 (N_1596,N_1329,N_1147);
nand U1597 (N_1597,N_273,N_928);
or U1598 (N_1598,N_636,N_910);
or U1599 (N_1599,In_1615,In_368);
nand U1600 (N_1600,N_377,In_2020);
xnor U1601 (N_1601,N_838,N_1081);
and U1602 (N_1602,N_659,In_1197);
or U1603 (N_1603,N_1362,N_1275);
xnor U1604 (N_1604,In_947,N_936);
and U1605 (N_1605,In_1171,N_887);
nand U1606 (N_1606,N_208,N_912);
and U1607 (N_1607,In_1041,N_1320);
or U1608 (N_1608,N_1321,N_434);
nand U1609 (N_1609,N_1423,In_1712);
nor U1610 (N_1610,In_2866,N_962);
nor U1611 (N_1611,N_1169,N_764);
xnor U1612 (N_1612,N_719,N_1201);
nand U1613 (N_1613,In_727,In_2387);
nor U1614 (N_1614,N_618,In_1560);
or U1615 (N_1615,N_810,N_1176);
xnor U1616 (N_1616,In_841,N_595);
nor U1617 (N_1617,N_1170,N_1192);
nand U1618 (N_1618,N_1475,N_1146);
nor U1619 (N_1619,N_1324,N_685);
nand U1620 (N_1620,In_2292,In_1299);
and U1621 (N_1621,N_1226,In_2791);
nand U1622 (N_1622,N_993,In_2848);
xor U1623 (N_1623,N_1456,In_1421);
or U1624 (N_1624,N_1418,N_1292);
or U1625 (N_1625,In_2707,In_608);
or U1626 (N_1626,In_1107,N_1234);
and U1627 (N_1627,N_958,N_0);
nor U1628 (N_1628,N_404,In_139);
nand U1629 (N_1629,In_2011,In_251);
nand U1630 (N_1630,In_2674,N_751);
and U1631 (N_1631,N_21,In_668);
nor U1632 (N_1632,N_1359,In_2639);
nor U1633 (N_1633,In_355,N_30);
and U1634 (N_1634,In_1762,N_706);
and U1635 (N_1635,N_1419,N_635);
nand U1636 (N_1636,In_1337,In_2120);
xor U1637 (N_1637,In_1912,In_1853);
xor U1638 (N_1638,N_453,In_53);
or U1639 (N_1639,In_854,N_1323);
or U1640 (N_1640,N_512,In_2540);
xnor U1641 (N_1641,In_2075,N_979);
nor U1642 (N_1642,In_2209,N_1127);
nand U1643 (N_1643,In_78,In_159);
and U1644 (N_1644,In_2311,N_581);
and U1645 (N_1645,In_2838,In_2291);
nor U1646 (N_1646,In_179,In_1865);
xor U1647 (N_1647,N_902,In_1042);
nand U1648 (N_1648,N_975,In_2420);
xor U1649 (N_1649,N_479,In_1699);
nand U1650 (N_1650,In_1486,N_627);
nand U1651 (N_1651,In_1020,N_1241);
xnor U1652 (N_1652,In_2519,N_1197);
or U1653 (N_1653,N_558,N_1200);
or U1654 (N_1654,N_579,In_2578);
nor U1655 (N_1655,N_1458,N_1159);
nor U1656 (N_1656,N_611,N_934);
xnor U1657 (N_1657,In_1445,In_634);
nand U1658 (N_1658,In_970,N_1208);
or U1659 (N_1659,In_2335,N_69);
xor U1660 (N_1660,N_1066,In_2554);
or U1661 (N_1661,In_1690,N_481);
nor U1662 (N_1662,In_1415,N_1497);
nor U1663 (N_1663,N_1466,N_1367);
nand U1664 (N_1664,In_1991,N_1332);
xor U1665 (N_1665,In_539,N_529);
or U1666 (N_1666,N_960,In_2390);
nand U1667 (N_1667,N_1215,N_672);
nand U1668 (N_1668,In_2336,In_2781);
nand U1669 (N_1669,N_1144,N_1405);
xor U1670 (N_1670,N_1179,N_757);
nor U1671 (N_1671,In_2253,In_1199);
or U1672 (N_1672,In_2485,In_1524);
and U1673 (N_1673,N_1431,In_2700);
nor U1674 (N_1674,In_2640,In_830);
nor U1675 (N_1675,In_1408,N_1374);
nand U1676 (N_1676,N_873,N_1027);
nor U1677 (N_1677,N_1045,N_724);
and U1678 (N_1678,N_1207,N_1440);
and U1679 (N_1679,N_284,N_1228);
or U1680 (N_1680,N_126,N_1236);
nor U1681 (N_1681,N_691,In_383);
nor U1682 (N_1682,In_2885,In_1318);
nor U1683 (N_1683,N_710,N_1043);
nor U1684 (N_1684,N_310,In_1516);
nor U1685 (N_1685,In_1660,In_320);
xnor U1686 (N_1686,N_322,In_1160);
xnor U1687 (N_1687,In_2310,In_1025);
nand U1688 (N_1688,N_1297,In_1743);
and U1689 (N_1689,N_1432,N_1391);
nor U1690 (N_1690,N_920,In_1612);
xor U1691 (N_1691,In_710,In_2126);
nor U1692 (N_1692,In_2445,In_1978);
nand U1693 (N_1693,N_1370,N_844);
and U1694 (N_1694,In_2231,In_1687);
xnor U1695 (N_1695,In_469,In_2459);
nand U1696 (N_1696,N_996,N_747);
xor U1697 (N_1697,N_998,N_1002);
and U1698 (N_1698,N_165,In_1081);
or U1699 (N_1699,In_1465,N_660);
xnor U1700 (N_1700,N_370,In_1911);
and U1701 (N_1701,N_1124,N_1287);
xor U1702 (N_1702,N_1202,In_1847);
xnor U1703 (N_1703,N_889,N_924);
and U1704 (N_1704,In_2287,N_926);
nand U1705 (N_1705,N_1078,In_2686);
xor U1706 (N_1706,N_1331,In_1822);
and U1707 (N_1707,N_1206,In_356);
xor U1708 (N_1708,In_1906,N_1481);
nand U1709 (N_1709,In_1180,In_2278);
xor U1710 (N_1710,In_1113,N_1376);
nor U1711 (N_1711,In_2494,N_1446);
nand U1712 (N_1712,N_1377,N_683);
nand U1713 (N_1713,In_2059,In_2637);
or U1714 (N_1714,In_485,N_379);
nand U1715 (N_1715,N_1442,N_904);
nand U1716 (N_1716,N_125,N_1358);
or U1717 (N_1717,N_891,In_2397);
and U1718 (N_1718,N_1148,N_669);
nor U1719 (N_1719,N_1238,N_1302);
xor U1720 (N_1720,In_553,In_486);
and U1721 (N_1721,In_1659,In_1147);
nand U1722 (N_1722,In_394,N_63);
and U1723 (N_1723,N_881,N_1412);
nand U1724 (N_1724,In_2891,N_1343);
nand U1725 (N_1725,N_789,In_322);
nand U1726 (N_1726,N_929,N_1397);
nand U1727 (N_1727,N_1282,In_2952);
nor U1728 (N_1728,N_906,N_1194);
xor U1729 (N_1729,In_1718,In_417);
and U1730 (N_1730,In_425,N_1433);
xor U1731 (N_1731,N_1269,In_171);
or U1732 (N_1732,N_1450,N_1474);
nor U1733 (N_1733,In_1446,In_317);
xnor U1734 (N_1734,N_1220,N_1385);
nand U1735 (N_1735,In_590,In_2170);
or U1736 (N_1736,In_847,N_1314);
or U1737 (N_1737,In_952,In_2319);
xnor U1738 (N_1738,In_891,N_92);
and U1739 (N_1739,In_1537,N_43);
nand U1740 (N_1740,In_2325,N_220);
nand U1741 (N_1741,N_1149,N_1461);
xnor U1742 (N_1742,In_1112,In_2713);
and U1743 (N_1743,N_1225,In_2993);
nor U1744 (N_1744,In_15,N_580);
or U1745 (N_1745,In_2216,N_1486);
xnor U1746 (N_1746,In_2037,N_1495);
and U1747 (N_1747,N_1394,In_818);
and U1748 (N_1748,In_1752,In_2357);
nand U1749 (N_1749,N_1487,N_959);
nand U1750 (N_1750,N_834,N_1361);
or U1751 (N_1751,In_1820,In_2830);
nand U1752 (N_1752,In_999,N_1451);
and U1753 (N_1753,N_1485,N_564);
and U1754 (N_1754,In_1471,In_1049);
and U1755 (N_1755,In_1834,N_1337);
xor U1756 (N_1756,N_1221,N_923);
nor U1757 (N_1757,N_850,N_1480);
nand U1758 (N_1758,N_1134,N_948);
nor U1759 (N_1759,In_2631,In_2388);
and U1760 (N_1760,In_1293,N_938);
xor U1761 (N_1761,In_943,N_216);
or U1762 (N_1762,In_2701,In_895);
nor U1763 (N_1763,In_2837,In_319);
xnor U1764 (N_1764,In_1504,In_1630);
xnor U1765 (N_1765,N_225,N_674);
and U1766 (N_1766,N_1188,In_1496);
nor U1767 (N_1767,In_2621,N_403);
or U1768 (N_1768,N_1268,In_2627);
or U1769 (N_1769,N_1183,N_263);
nor U1770 (N_1770,In_201,In_2872);
or U1771 (N_1771,N_1288,N_822);
or U1772 (N_1772,N_507,N_357);
and U1773 (N_1773,N_952,N_151);
and U1774 (N_1774,In_2088,N_1132);
nor U1775 (N_1775,N_1003,In_711);
nand U1776 (N_1776,In_737,N_1356);
or U1777 (N_1777,In_43,N_818);
and U1778 (N_1778,N_1434,In_2492);
nand U1779 (N_1779,In_1141,In_1681);
and U1780 (N_1780,N_860,In_1554);
nor U1781 (N_1781,In_237,N_1349);
and U1782 (N_1782,In_584,N_1378);
and U1783 (N_1783,In_1631,In_2953);
nor U1784 (N_1784,N_1355,N_1116);
or U1785 (N_1785,N_1193,In_1056);
or U1786 (N_1786,In_2945,N_1414);
xor U1787 (N_1787,N_380,In_467);
xor U1788 (N_1788,In_2084,In_2269);
or U1789 (N_1789,N_1033,N_767);
nor U1790 (N_1790,N_1317,N_1449);
and U1791 (N_1791,In_18,N_939);
nor U1792 (N_1792,In_1248,N_1463);
nand U1793 (N_1793,In_2723,N_524);
nor U1794 (N_1794,In_1234,N_1389);
and U1795 (N_1795,N_64,In_717);
and U1796 (N_1796,N_313,N_587);
and U1797 (N_1797,N_1464,In_1900);
xnor U1798 (N_1798,N_390,In_278);
nor U1799 (N_1799,N_1254,N_999);
nor U1800 (N_1800,N_1256,N_1235);
nand U1801 (N_1801,N_1199,N_833);
xnor U1802 (N_1802,N_1162,N_1088);
and U1803 (N_1803,N_1260,N_1614);
nand U1804 (N_1804,In_2002,In_1285);
xnor U1805 (N_1805,In_1026,N_1758);
nor U1806 (N_1806,N_1543,N_1574);
nor U1807 (N_1807,N_214,N_415);
nand U1808 (N_1808,In_754,N_1683);
nor U1809 (N_1809,N_1760,N_534);
nor U1810 (N_1810,N_1335,N_1692);
nor U1811 (N_1811,N_977,N_1577);
nor U1812 (N_1812,N_520,N_1096);
nor U1813 (N_1813,N_1372,In_435);
xor U1814 (N_1814,N_1222,N_1773);
or U1815 (N_1815,N_1715,In_2348);
nand U1816 (N_1816,N_1668,N_1375);
nand U1817 (N_1817,N_1625,N_1508);
nand U1818 (N_1818,In_318,N_1748);
nand U1819 (N_1819,N_1278,N_1388);
or U1820 (N_1820,In_1170,N_1780);
nor U1821 (N_1821,N_1053,N_1384);
or U1822 (N_1822,N_1523,In_1841);
nor U1823 (N_1823,N_1718,N_1520);
nor U1824 (N_1824,N_1547,N_1734);
nand U1825 (N_1825,N_470,N_1060);
and U1826 (N_1826,In_563,N_1195);
or U1827 (N_1827,N_649,N_484);
nor U1828 (N_1828,N_1549,In_119);
nor U1829 (N_1829,N_714,In_2190);
nand U1830 (N_1830,N_951,N_1048);
nor U1831 (N_1831,N_702,N_417);
or U1832 (N_1832,N_113,N_447);
nand U1833 (N_1833,N_1447,N_1587);
or U1834 (N_1834,In_287,In_2432);
xnor U1835 (N_1835,In_2604,N_1750);
or U1836 (N_1836,N_1071,N_1119);
and U1837 (N_1837,N_1650,N_1512);
and U1838 (N_1838,In_2666,N_222);
nand U1839 (N_1839,N_1219,N_1694);
and U1840 (N_1840,N_1530,N_1686);
xnor U1841 (N_1841,In_282,N_1240);
or U1842 (N_1842,N_1040,In_1129);
nor U1843 (N_1843,N_1590,In_549);
xnor U1844 (N_1844,In_739,In_352);
xor U1845 (N_1845,N_599,N_1612);
nor U1846 (N_1846,N_1106,In_2439);
or U1847 (N_1847,N_1698,In_71);
nor U1848 (N_1848,N_1368,N_346);
and U1849 (N_1849,N_1513,N_1319);
and U1850 (N_1850,N_804,In_1344);
nor U1851 (N_1851,N_1723,N_1299);
or U1852 (N_1852,N_1554,N_1568);
xor U1853 (N_1853,In_1588,N_1050);
and U1854 (N_1854,N_1796,N_1671);
nor U1855 (N_1855,N_24,In_2552);
xor U1856 (N_1856,N_1232,N_1687);
nor U1857 (N_1857,N_1261,In_145);
nor U1858 (N_1858,N_1742,In_103);
nand U1859 (N_1859,In_2095,In_1466);
xor U1860 (N_1860,N_1714,N_1585);
and U1861 (N_1861,N_44,N_1315);
xor U1862 (N_1862,N_1737,N_1379);
xnor U1863 (N_1863,N_1592,N_898);
or U1864 (N_1864,N_1732,N_1231);
xor U1865 (N_1865,N_985,N_1602);
nand U1866 (N_1866,In_1676,N_428);
nor U1867 (N_1867,N_1604,N_964);
and U1868 (N_1868,N_575,N_1768);
nor U1869 (N_1869,N_676,In_1162);
nand U1870 (N_1870,N_1628,In_1489);
nand U1871 (N_1871,N_771,N_413);
or U1872 (N_1872,N_1503,N_1247);
nor U1873 (N_1873,N_1669,In_2281);
or U1874 (N_1874,In_1758,N_1793);
and U1875 (N_1875,In_2372,N_1350);
nand U1876 (N_1876,N_461,N_1680);
nand U1877 (N_1877,In_1278,N_233);
or U1878 (N_1878,In_858,N_1639);
nand U1879 (N_1879,In_118,N_1605);
xor U1880 (N_1880,N_490,N_1710);
and U1881 (N_1881,In_1139,N_1713);
nor U1882 (N_1882,N_1699,In_1217);
nor U1883 (N_1883,In_2581,In_2794);
and U1884 (N_1884,N_721,N_1542);
or U1885 (N_1885,N_1597,N_1652);
xnor U1886 (N_1886,In_1190,N_181);
nand U1887 (N_1887,N_1289,In_2916);
and U1888 (N_1888,In_989,In_2234);
nor U1889 (N_1889,In_1054,N_1363);
and U1890 (N_1890,N_1428,N_1759);
nand U1891 (N_1891,N_1276,N_1312);
nor U1892 (N_1892,N_623,In_589);
nand U1893 (N_1893,N_1681,In_2422);
nand U1894 (N_1894,N_816,N_1672);
xor U1895 (N_1895,N_1012,In_458);
or U1896 (N_1896,N_1755,N_1563);
and U1897 (N_1897,N_1556,In_2296);
or U1898 (N_1898,In_581,N_1735);
xor U1899 (N_1899,N_1239,N_462);
or U1900 (N_1900,In_328,N_1569);
and U1901 (N_1901,N_435,N_1150);
nor U1902 (N_1902,N_530,N_398);
nand U1903 (N_1903,N_1178,N_1797);
nor U1904 (N_1904,In_1750,N_38);
nand U1905 (N_1905,N_135,N_1515);
nand U1906 (N_1906,N_1415,N_394);
xor U1907 (N_1907,N_289,In_476);
nand U1908 (N_1908,N_1462,In_1701);
xnor U1909 (N_1909,In_815,N_955);
xnor U1910 (N_1910,N_1248,N_1778);
and U1911 (N_1911,N_982,N_1242);
nor U1912 (N_1912,N_1533,In_2314);
xor U1913 (N_1913,N_1212,In_1484);
nand U1914 (N_1914,N_1703,N_1244);
and U1915 (N_1915,In_2464,N_1711);
xnor U1916 (N_1916,N_694,N_645);
nor U1917 (N_1917,N_1311,N_943);
or U1918 (N_1918,N_918,In_1396);
or U1919 (N_1919,In_1301,In_517);
nand U1920 (N_1920,In_92,N_1135);
nor U1921 (N_1921,N_1398,N_1402);
or U1922 (N_1922,N_1445,N_594);
xor U1923 (N_1923,N_1716,N_1342);
or U1924 (N_1924,N_755,N_360);
and U1925 (N_1925,In_335,N_1164);
xor U1926 (N_1926,In_2243,N_602);
xor U1927 (N_1927,N_662,N_1056);
nor U1928 (N_1928,N_1216,In_2085);
xor U1929 (N_1929,N_980,N_648);
nand U1930 (N_1930,N_984,In_501);
and U1931 (N_1931,N_1684,In_2709);
nand U1932 (N_1932,In_537,N_916);
xor U1933 (N_1933,In_1314,In_80);
nand U1934 (N_1934,In_635,N_917);
nand U1935 (N_1935,N_391,N_591);
or U1936 (N_1936,N_1561,In_1692);
xor U1937 (N_1937,In_2867,N_432);
xnor U1938 (N_1938,N_1214,N_1610);
nand U1939 (N_1939,In_2706,In_692);
xor U1940 (N_1940,In_2603,N_1460);
nor U1941 (N_1941,In_1066,N_1740);
xnor U1942 (N_1942,In_2530,N_1730);
nor U1943 (N_1943,N_1706,N_1032);
nor U1944 (N_1944,N_1217,N_1017);
xor U1945 (N_1945,N_1117,N_1522);
nor U1946 (N_1946,N_799,N_1184);
and U1947 (N_1947,In_2187,In_552);
xnor U1948 (N_1948,N_1223,N_736);
xor U1949 (N_1949,N_1660,N_47);
xnor U1950 (N_1950,In_175,In_2821);
or U1951 (N_1951,N_70,N_1576);
nor U1952 (N_1952,N_1251,N_1283);
or U1953 (N_1953,In_783,In_1365);
xnor U1954 (N_1954,In_633,N_1298);
or U1955 (N_1955,N_362,N_1422);
nor U1956 (N_1956,N_1396,N_908);
nor U1957 (N_1957,N_1191,N_414);
nor U1958 (N_1958,N_300,N_1608);
and U1959 (N_1959,In_1508,N_232);
or U1960 (N_1960,In_1728,In_860);
and U1961 (N_1961,N_1072,In_1116);
nor U1962 (N_1962,N_93,N_1122);
nor U1963 (N_1963,In_1404,N_1521);
xor U1964 (N_1964,N_1541,In_2966);
and U1965 (N_1965,In_643,In_2638);
nand U1966 (N_1966,N_1689,N_886);
and U1967 (N_1967,N_1443,In_2119);
nand U1968 (N_1968,N_1213,N_1790);
or U1969 (N_1969,In_1151,In_2481);
nand U1970 (N_1970,N_1787,N_1525);
nand U1971 (N_1971,N_1125,N_879);
or U1972 (N_1972,In_1166,N_1496);
xor U1973 (N_1973,N_1659,N_839);
nand U1974 (N_1974,N_1727,In_13);
xor U1975 (N_1975,In_2199,In_1154);
nand U1976 (N_1976,N_1491,N_1006);
or U1977 (N_1977,N_1152,N_1273);
and U1978 (N_1978,In_928,N_845);
xnor U1979 (N_1979,N_1262,In_1563);
nor U1980 (N_1980,N_1473,In_1313);
xor U1981 (N_1981,N_1721,N_1588);
or U1982 (N_1982,In_1159,N_1403);
and U1983 (N_1983,In_1053,N_286);
nand U1984 (N_1984,N_175,N_1555);
nor U1985 (N_1985,N_257,N_305);
xor U1986 (N_1986,N_986,N_1783);
xnor U1987 (N_1987,In_1582,N_784);
and U1988 (N_1988,In_583,N_1682);
nand U1989 (N_1989,In_654,N_976);
and U1990 (N_1990,N_1657,In_1885);
nand U1991 (N_1991,N_1630,N_1120);
xor U1992 (N_1992,N_504,N_880);
xor U1993 (N_1993,In_1777,N_1448);
xor U1994 (N_1994,N_571,N_868);
and U1995 (N_1995,N_1272,N_1454);
and U1996 (N_1996,N_1277,N_1532);
nand U1997 (N_1997,N_1285,N_633);
nand U1998 (N_1998,In_2125,N_1772);
and U1999 (N_1999,N_528,In_1142);
nor U2000 (N_2000,N_178,N_1326);
or U2001 (N_2001,In_743,In_1685);
nand U2002 (N_2002,N_1596,In_504);
or U2003 (N_2003,N_651,N_631);
or U2004 (N_2004,In_2273,In_1478);
and U2005 (N_2005,N_1233,N_1155);
nor U2006 (N_2006,N_469,N_1205);
xor U2007 (N_2007,N_1631,N_1103);
xnor U2008 (N_2008,In_2770,N_1354);
nor U2009 (N_2009,N_1154,In_459);
nand U2010 (N_2010,N_1559,N_1180);
nand U2011 (N_2011,N_1290,N_1566);
and U2012 (N_2012,N_265,In_1971);
nor U2013 (N_2013,N_1564,N_1765);
or U2014 (N_2014,In_1720,In_2863);
xor U2015 (N_2015,N_1479,N_1616);
nor U2016 (N_2016,N_1051,N_944);
and U2017 (N_2017,N_1210,N_1572);
xnor U2018 (N_2018,In_812,N_1465);
nand U2019 (N_2019,In_1917,In_1543);
xor U2020 (N_2020,In_2905,N_1546);
nand U2021 (N_2021,In_1315,N_903);
xnor U2022 (N_2022,N_53,In_1238);
or U2023 (N_2023,N_1634,N_1506);
or U2024 (N_2024,In_2305,In_2100);
nor U2025 (N_2025,N_280,In_788);
nand U2026 (N_2026,In_848,N_1316);
or U2027 (N_2027,N_1185,N_703);
xnor U2028 (N_2028,N_1558,In_195);
and U2029 (N_2029,N_1557,In_2990);
xor U2030 (N_2030,In_1884,In_1734);
xor U2031 (N_2031,N_1230,N_1494);
and U2032 (N_2032,In_2999,N_1670);
nor U2033 (N_2033,In_31,N_1203);
nand U2034 (N_2034,In_1249,N_60);
xnor U2035 (N_2035,In_1453,In_151);
or U2036 (N_2036,In_595,In_499);
nor U2037 (N_2037,N_1074,N_1545);
nand U2038 (N_2038,In_1930,N_1279);
and U2039 (N_2039,N_1728,N_1606);
nor U2040 (N_2040,N_224,In_2156);
and U2041 (N_2041,N_1253,In_1855);
xor U2042 (N_2042,In_1206,N_76);
nor U2043 (N_2043,In_2904,In_2500);
nand U2044 (N_2044,In_816,N_1617);
nor U2045 (N_2045,N_288,N_1504);
nand U2046 (N_2046,In_683,N_927);
nor U2047 (N_2047,N_1595,In_877);
nor U2048 (N_2048,N_1517,In_375);
or U2049 (N_2049,N_785,N_666);
xor U2050 (N_2050,In_2468,N_1249);
xnor U2051 (N_2051,N_1008,N_1536);
or U2052 (N_2052,N_218,In_226);
nand U2053 (N_2053,N_196,In_2349);
or U2054 (N_2054,N_1764,N_1255);
nor U2055 (N_2055,N_896,N_25);
and U2056 (N_2056,N_641,N_617);
and U2057 (N_2057,In_224,N_1770);
or U2058 (N_2058,In_2039,N_629);
nand U2059 (N_2059,N_242,In_384);
nand U2060 (N_2060,In_2476,N_1591);
and U2061 (N_2061,N_1167,N_54);
nand U2062 (N_2062,N_1393,In_2139);
xor U2063 (N_2063,N_643,N_1761);
nor U2064 (N_2064,In_373,N_375);
xnor U2065 (N_2065,N_1382,In_1599);
nand U2066 (N_2066,N_1156,N_1560);
xnor U2067 (N_2067,N_1636,N_1675);
and U2068 (N_2068,N_1528,In_75);
nand U2069 (N_2069,N_104,In_2582);
nand U2070 (N_2070,In_2389,In_163);
nand U2071 (N_2071,N_1571,In_964);
and U2072 (N_2072,N_1584,N_1691);
or U2073 (N_2073,N_961,N_1052);
nand U2074 (N_2074,In_2975,N_445);
and U2075 (N_2075,In_2927,N_1724);
or U2076 (N_2076,N_401,N_1293);
nor U2077 (N_2077,N_796,In_829);
or U2078 (N_2078,N_1745,N_1792);
nand U2079 (N_2079,N_1348,In_1812);
xnor U2080 (N_2080,In_2007,In_656);
or U2081 (N_2081,N_1705,In_225);
or U2082 (N_2082,In_380,N_905);
nor U2083 (N_2083,In_37,N_870);
or U2084 (N_2084,N_1578,N_150);
or U2085 (N_2085,In_339,N_1381);
nor U2086 (N_2086,In_809,N_775);
nor U2087 (N_2087,N_1776,In_744);
nand U2088 (N_2088,N_930,In_248);
or U2089 (N_2089,In_2424,N_1615);
xnor U2090 (N_2090,In_2223,N_1779);
nor U2091 (N_2091,N_830,N_1387);
nor U2092 (N_2092,In_1744,In_2064);
or U2093 (N_2093,N_1190,In_2484);
and U2094 (N_2094,N_45,N_1529);
and U2095 (N_2095,In_1698,N_1095);
nor U2096 (N_2096,In_2294,In_450);
nand U2097 (N_2097,N_1583,N_1039);
nor U2098 (N_2098,In_2409,In_1787);
xor U2099 (N_2099,N_1439,N_763);
xnor U2100 (N_2100,N_1678,N_1539);
nand U2101 (N_2101,N_124,N_1757);
and U2102 (N_2102,N_1410,In_1296);
nor U2103 (N_2103,N_1101,N_1979);
nand U2104 (N_2104,N_723,N_921);
or U2105 (N_2105,N_1077,N_1492);
and U2106 (N_2106,N_1822,N_1264);
or U2107 (N_2107,In_1444,N_1909);
nand U2108 (N_2108,N_1548,N_1218);
xnor U2109 (N_2109,N_2078,N_277);
and U2110 (N_2110,N_1704,In_156);
nor U2111 (N_2111,N_1871,In_1281);
nor U2112 (N_2112,N_2079,N_1902);
or U2113 (N_2113,N_1897,In_2080);
or U2114 (N_2114,N_1884,N_1579);
or U2115 (N_2115,N_1806,N_1752);
nand U2116 (N_2116,N_1960,N_1534);
nor U2117 (N_2117,N_680,N_1812);
nand U2118 (N_2118,N_1696,N_2083);
nand U2119 (N_2119,N_1637,N_2085);
xor U2120 (N_2120,In_189,N_1843);
nand U2121 (N_2121,N_2009,N_1295);
or U2122 (N_2122,N_989,In_1771);
and U2123 (N_2123,N_1781,N_610);
and U2124 (N_2124,N_1417,In_2874);
xnor U2125 (N_2125,N_1237,N_2090);
and U2126 (N_2126,N_1927,N_1345);
xnor U2127 (N_2127,N_1749,N_1824);
nand U2128 (N_2128,N_2070,N_1172);
and U2129 (N_2129,N_1263,N_1177);
xor U2130 (N_2130,N_2003,N_915);
or U2131 (N_2131,N_2080,N_2054);
nor U2132 (N_2132,In_1104,N_2007);
nand U2133 (N_2133,N_1919,N_348);
and U2134 (N_2134,N_2052,N_1695);
xor U2135 (N_2135,In_178,In_2152);
nand U2136 (N_2136,In_560,In_819);
xor U2137 (N_2137,N_1985,N_1751);
nor U2138 (N_2138,N_907,In_806);
nor U2139 (N_2139,N_1421,N_1490);
or U2140 (N_2140,N_1153,N_1907);
nand U2141 (N_2141,N_954,N_527);
and U2142 (N_2142,N_1863,N_239);
or U2143 (N_2143,In_332,N_1435);
nand U2144 (N_2144,N_1839,N_1501);
nand U2145 (N_2145,N_2065,N_1505);
nand U2146 (N_2146,N_1883,In_2606);
nand U2147 (N_2147,N_1246,In_1252);
xnor U2148 (N_2148,N_2071,N_729);
xor U2149 (N_2149,In_1665,N_1920);
and U2150 (N_2150,N_1409,N_2077);
and U2151 (N_2151,N_1846,N_1805);
or U2152 (N_2152,N_1609,In_449);
or U2153 (N_2153,N_1137,N_2064);
and U2154 (N_2154,In_1998,N_2063);
or U2155 (N_2155,N_1531,N_1601);
and U2156 (N_2156,In_580,In_446);
nand U2157 (N_2157,N_1841,N_2084);
nand U2158 (N_2158,N_1931,N_1064);
xor U2159 (N_2159,N_1990,N_909);
and U2160 (N_2160,In_688,N_2046);
xor U2161 (N_2161,N_1425,N_1873);
nor U2162 (N_2162,In_2043,N_1586);
xor U2163 (N_2163,N_1633,In_2177);
nor U2164 (N_2164,N_737,N_1955);
nor U2165 (N_2165,N_1344,N_1281);
nor U2166 (N_2166,N_1967,N_1874);
or U2167 (N_2167,N_1567,In_775);
nand U2168 (N_2168,N_1848,N_1383);
xor U2169 (N_2169,N_1946,In_2133);
and U2170 (N_2170,N_1934,N_2072);
nand U2171 (N_2171,N_2022,N_1767);
nor U2172 (N_2172,N_2069,N_1995);
nand U2173 (N_2173,N_1114,N_863);
xor U2174 (N_2174,N_142,In_2290);
nor U2175 (N_2175,N_519,N_78);
or U2176 (N_2176,N_762,N_2067);
and U2177 (N_2177,N_1832,N_1756);
xnor U2178 (N_2178,N_1408,In_1544);
and U2179 (N_2179,In_1737,N_1493);
xor U2180 (N_2180,N_1058,N_1954);
nor U2181 (N_2181,N_1036,N_1598);
or U2182 (N_2182,N_1112,N_1476);
nor U2183 (N_2183,N_501,N_1847);
nand U2184 (N_2184,In_68,N_1994);
xnor U2185 (N_2185,N_2015,In_1882);
and U2186 (N_2186,N_1987,N_1860);
nor U2187 (N_2187,N_1693,N_1509);
nand U2188 (N_2188,N_2012,N_1785);
and U2189 (N_2189,In_491,In_2981);
nand U2190 (N_2190,In_1034,N_967);
nand U2191 (N_2191,N_1526,N_2036);
xor U2192 (N_2192,N_1827,N_1392);
and U2193 (N_2193,In_2391,In_489);
nor U2194 (N_2194,N_1964,N_250);
and U2195 (N_2195,In_470,N_637);
nor U2196 (N_2196,In_1294,N_1245);
and U2197 (N_2197,N_1544,N_1655);
nand U2198 (N_2198,N_1986,N_1800);
xor U2199 (N_2199,In_1921,N_1950);
xnor U2200 (N_2200,N_2000,N_1788);
or U2201 (N_2201,N_1878,N_1643);
nor U2202 (N_2202,N_2028,N_383);
or U2203 (N_2203,N_1880,N_1801);
or U2204 (N_2204,N_2089,N_1339);
nor U2205 (N_2205,N_1830,In_327);
nand U2206 (N_2206,N_872,N_1959);
nand U2207 (N_2207,N_2074,N_1881);
nand U2208 (N_2208,In_807,N_1972);
nand U2209 (N_2209,N_2040,In_2034);
nor U2210 (N_2210,N_1939,N_1498);
xor U2211 (N_2211,N_1965,N_1457);
or U2212 (N_2212,N_1867,N_1097);
nand U2213 (N_2213,N_1849,N_1665);
or U2214 (N_2214,N_1707,N_1736);
xnor U2215 (N_2215,In_1236,N_817);
and U2216 (N_2216,N_1777,N_2021);
and U2217 (N_2217,In_1202,In_1377);
nor U2218 (N_2218,N_180,N_329);
xnor U2219 (N_2219,N_2066,N_1426);
or U2220 (N_2220,N_1762,N_1524);
or U2221 (N_2221,N_1904,In_418);
nor U2222 (N_2222,N_1865,N_1673);
or U2223 (N_2223,N_1838,N_1581);
nand U2224 (N_2224,N_1250,N_1618);
nand U2225 (N_2225,N_2027,In_1577);
nand U2226 (N_2226,N_574,N_1935);
and U2227 (N_2227,N_2039,N_1708);
and U2228 (N_2228,N_1110,N_1252);
xor U2229 (N_2229,N_1818,N_1925);
nand U2230 (N_2230,N_2050,N_1891);
and U2231 (N_2231,N_1983,N_2011);
or U2232 (N_2232,N_1401,N_140);
nor U2233 (N_2233,N_2048,N_1700);
nor U2234 (N_2234,N_2008,N_1690);
nand U2235 (N_2235,In_2326,N_2060);
nand U2236 (N_2236,N_1915,N_1943);
or U2237 (N_2237,N_1998,N_1901);
xnor U2238 (N_2238,N_1514,N_1390);
or U2239 (N_2239,N_1763,N_1869);
and U2240 (N_2240,N_1593,N_1916);
or U2241 (N_2241,N_2062,In_1898);
and U2242 (N_2242,N_1791,In_1585);
nor U2243 (N_2243,In_1387,N_1307);
nand U2244 (N_2244,N_1733,N_2016);
or U2245 (N_2245,N_1823,N_1968);
or U2246 (N_2246,N_1313,In_2138);
xnor U2247 (N_2247,In_2330,In_2748);
and U2248 (N_2248,N_1037,In_554);
or U2249 (N_2249,N_1429,N_1482);
nor U2250 (N_2250,N_1666,N_1804);
nand U2251 (N_2251,N_1837,N_1688);
nand U2252 (N_2252,N_1817,N_2019);
nand U2253 (N_2253,N_1057,N_1271);
and U2254 (N_2254,N_1936,In_2060);
nor U2255 (N_2255,N_1623,N_1887);
or U2256 (N_2256,In_2196,In_869);
xor U2257 (N_2257,N_255,N_593);
xnor U2258 (N_2258,N_1538,N_1484);
or U2259 (N_2259,N_2094,N_1810);
and U2260 (N_2260,In_428,N_1816);
and U2261 (N_2261,N_1406,In_2762);
nand U2262 (N_2262,In_1072,N_1857);
or U2263 (N_2263,N_772,In_2531);
xnor U2264 (N_2264,In_1099,N_1021);
nor U2265 (N_2265,N_1653,In_1785);
nand U2266 (N_2266,N_1798,N_1500);
xnor U2267 (N_2267,N_2051,In_1164);
nor U2268 (N_2268,N_1913,In_911);
xnor U2269 (N_2269,N_1489,In_756);
nor U2270 (N_2270,N_569,N_1259);
and U2271 (N_2271,N_1855,N_1243);
nand U2272 (N_2272,N_1352,N_1638);
xnor U2273 (N_2273,N_1938,In_1040);
and U2274 (N_2274,N_1175,N_1641);
xnor U2275 (N_2275,N_1459,In_1323);
or U2276 (N_2276,In_2049,In_2220);
or U2277 (N_2277,N_1291,N_1371);
nand U2278 (N_2278,N_695,In_2379);
and U2279 (N_2279,N_1347,In_98);
and U2280 (N_2280,N_1807,N_1888);
or U2281 (N_2281,N_1047,N_1042);
xnor U2282 (N_2282,N_566,N_1024);
nor U2283 (N_2283,In_1290,In_796);
and U2284 (N_2284,In_1757,N_1015);
xnor U2285 (N_2285,N_1308,N_1082);
xor U2286 (N_2286,N_1488,N_1121);
xnor U2287 (N_2287,N_1784,N_832);
xnor U2288 (N_2288,In_488,N_1958);
nor U2289 (N_2289,In_2068,N_1662);
and U2290 (N_2290,N_1717,N_1741);
nor U2291 (N_2291,In_651,N_1813);
nor U2292 (N_2292,In_1441,N_1859);
nor U2293 (N_2293,In_2729,N_1341);
or U2294 (N_2294,In_170,N_2005);
nand U2295 (N_2295,In_1384,N_1795);
or U2296 (N_2296,N_1821,In_528);
nand U2297 (N_2297,N_1864,N_991);
and U2298 (N_2298,N_1991,N_2026);
or U2299 (N_2299,N_1856,N_1719);
and U2300 (N_2300,N_1853,In_2963);
xor U2301 (N_2301,N_1369,N_1754);
nor U2302 (N_2302,In_624,N_2033);
and U2303 (N_2303,In_1943,In_821);
xnor U2304 (N_2304,N_1831,N_1731);
or U2305 (N_2305,N_1085,N_2087);
nor U2306 (N_2306,N_1535,N_1646);
nor U2307 (N_2307,N_1942,In_410);
xor U2308 (N_2308,In_2212,N_1102);
nor U2309 (N_2309,In_223,N_1825);
nor U2310 (N_2310,N_1265,N_1782);
and U2311 (N_2311,N_1651,In_1455);
or U2312 (N_2312,N_1656,N_1918);
or U2313 (N_2313,N_1041,In_202);
nand U2314 (N_2314,N_1933,N_1766);
nor U2315 (N_2315,N_2023,In_1437);
nand U2316 (N_2316,N_1562,In_874);
and U2317 (N_2317,N_1980,N_1420);
and U2318 (N_2318,N_1516,In_1413);
xor U2319 (N_2319,N_1158,N_650);
nor U2320 (N_2320,N_1550,N_1141);
or U2321 (N_2321,N_1895,N_942);
and U2322 (N_2322,N_2076,N_1603);
xnor U2323 (N_2323,N_1738,N_1573);
xnor U2324 (N_2324,N_1890,N_2025);
and U2325 (N_2325,N_568,N_291);
or U2326 (N_2326,N_1803,N_1613);
nand U2327 (N_2327,N_1580,In_2050);
nand U2328 (N_2328,N_2018,N_1973);
and U2329 (N_2329,N_1808,In_1561);
xor U2330 (N_2330,In_242,N_653);
xor U2331 (N_2331,N_1629,N_1877);
and U2332 (N_2332,N_1607,N_1876);
and U2333 (N_2333,N_1974,N_2086);
and U2334 (N_2334,N_601,N_2045);
nand U2335 (N_2335,N_1870,N_791);
xor U2336 (N_2336,N_83,N_2056);
and U2337 (N_2337,N_1858,In_1231);
nor U2338 (N_2338,N_1844,N_671);
xnor U2339 (N_2339,In_2456,N_1330);
or U2340 (N_2340,N_1552,N_1518);
nand U2341 (N_2341,In_555,In_1854);
nor U2342 (N_2342,N_1502,N_2098);
or U2343 (N_2343,In_1149,In_1536);
xor U2344 (N_2344,N_1962,N_1565);
nand U2345 (N_2345,N_1209,N_1885);
nor U2346 (N_2346,N_1911,In_2670);
and U2347 (N_2347,N_974,In_1475);
nor U2348 (N_2348,In_1004,N_2099);
nor U2349 (N_2349,N_1645,N_2073);
xor U2350 (N_2350,In_1251,N_1908);
or U2351 (N_2351,N_1944,N_745);
or U2352 (N_2352,N_1969,N_2001);
or U2353 (N_2353,N_2010,N_2006);
xor U2354 (N_2354,N_1677,In_1332);
and U2355 (N_2355,N_1720,N_549);
nand U2356 (N_2356,N_711,N_2059);
or U2357 (N_2357,N_1739,N_1211);
or U2358 (N_2358,N_1945,N_1407);
or U2359 (N_2359,N_1900,N_1360);
or U2360 (N_2360,N_2096,N_1854);
and U2361 (N_2361,N_1589,N_1632);
and U2362 (N_2362,N_1982,N_1988);
and U2363 (N_2363,N_1851,N_101);
or U2364 (N_2364,N_1952,N_919);
nor U2365 (N_2365,N_1351,N_827);
or U2366 (N_2366,N_1087,N_1441);
xor U2367 (N_2367,N_1828,N_1941);
xnor U2368 (N_2368,N_1903,N_1932);
or U2369 (N_2369,N_1619,In_2202);
or U2370 (N_2370,N_1647,N_1875);
nand U2371 (N_2371,N_1886,N_592);
nor U2372 (N_2372,N_2081,N_2047);
nand U2373 (N_2373,N_2014,In_1603);
nand U2374 (N_2374,In_1006,N_1951);
nor U2375 (N_2375,In_2736,N_2029);
xor U2376 (N_2376,N_2095,N_130);
and U2377 (N_2377,In_1182,N_1624);
or U2378 (N_2378,N_1771,In_996);
and U2379 (N_2379,N_1395,N_859);
or U2380 (N_2380,N_1917,N_652);
xor U2381 (N_2381,In_2221,N_1309);
xor U2382 (N_2382,In_1610,In_1232);
nor U2383 (N_2383,In_1507,N_2031);
and U2384 (N_2384,N_1799,In_2688);
xor U2385 (N_2385,N_777,N_2037);
nor U2386 (N_2386,N_1366,N_344);
nor U2387 (N_2387,N_1031,In_2384);
or U2388 (N_2388,N_829,N_1510);
and U2389 (N_2389,N_1809,N_1600);
nor U2390 (N_2390,In_2962,N_1977);
nand U2391 (N_2391,In_1878,N_572);
and U2392 (N_2392,In_696,N_1892);
and U2393 (N_2393,N_1712,In_738);
or U2394 (N_2394,N_715,N_1644);
and U2395 (N_2395,In_715,In_2944);
and U2396 (N_2396,N_1519,N_1923);
nor U2397 (N_2397,In_1360,In_2394);
xnor U2398 (N_2398,N_303,N_1914);
nand U2399 (N_2399,In_1284,N_1992);
nor U2400 (N_2400,N_1836,N_2300);
nand U2401 (N_2401,N_2365,N_1511);
and U2402 (N_2402,N_2210,N_2188);
xor U2403 (N_2403,In_1709,N_1621);
xnor U2404 (N_2404,N_2255,N_2311);
and U2405 (N_2405,In_880,N_2305);
nor U2406 (N_2406,N_1852,N_2262);
nand U2407 (N_2407,N_1139,N_2284);
or U2408 (N_2408,N_2348,In_2);
or U2409 (N_2409,N_820,In_2625);
nor U2410 (N_2410,N_1814,N_2091);
and U2411 (N_2411,In_1048,N_1746);
xor U2412 (N_2412,N_1676,N_2041);
nand U2413 (N_2413,N_2307,In_1321);
xnor U2414 (N_2414,In_1145,N_2251);
and U2415 (N_2415,In_1826,N_2245);
xor U2416 (N_2416,N_2119,N_2239);
or U2417 (N_2417,N_2265,N_2211);
and U2418 (N_2418,N_2334,N_1769);
and U2419 (N_2419,N_2189,N_2299);
and U2420 (N_2420,N_1981,N_1654);
xnor U2421 (N_2421,In_1333,N_2227);
and U2422 (N_2422,N_2234,N_1084);
nand U2423 (N_2423,N_634,N_2075);
nor U2424 (N_2424,N_2017,N_2323);
xor U2425 (N_2425,In_2396,N_2143);
nand U2426 (N_2426,N_2331,N_2329);
xor U2427 (N_2427,N_1940,N_628);
or U2428 (N_2428,N_2145,N_2061);
or U2429 (N_2429,N_1906,N_2164);
xnor U2430 (N_2430,N_2285,N_1661);
xor U2431 (N_2431,N_2277,N_2319);
xnor U2432 (N_2432,N_2185,In_2255);
xor U2433 (N_2433,N_2364,In_498);
or U2434 (N_2434,N_1834,N_2173);
or U2435 (N_2435,N_2375,N_1131);
or U2436 (N_2436,N_941,N_2356);
xnor U2437 (N_2437,In_1907,N_2387);
and U2438 (N_2438,N_1905,N_2366);
nand U2439 (N_2439,N_1924,N_1956);
or U2440 (N_2440,In_961,N_2159);
nand U2441 (N_2441,N_1582,N_2004);
and U2442 (N_2442,In_1923,N_2035);
xnor U2443 (N_2443,N_2124,In_44);
nor U2444 (N_2444,N_2309,N_2147);
nand U2445 (N_2445,In_2555,N_2157);
xnor U2446 (N_2446,N_2398,N_1073);
or U2447 (N_2447,N_2377,N_2088);
and U2448 (N_2448,N_2032,N_1649);
nor U2449 (N_2449,N_2136,N_2043);
nand U2450 (N_2450,N_2146,N_2391);
and U2451 (N_2451,In_1256,N_2370);
and U2452 (N_2452,N_2114,N_2340);
nand U2453 (N_2453,N_2182,N_1953);
or U2454 (N_2454,N_2002,N_2161);
or U2455 (N_2455,In_2535,N_2024);
and U2456 (N_2456,N_2163,N_1286);
and U2457 (N_2457,In_2692,N_2058);
and U2458 (N_2458,N_2332,N_1611);
and U2459 (N_2459,N_1123,N_295);
nor U2460 (N_2460,N_2252,N_2168);
nand U2461 (N_2461,In_2288,N_2106);
and U2462 (N_2462,N_2256,N_1594);
nor U2463 (N_2463,N_2201,N_1143);
and U2464 (N_2464,N_2140,N_2053);
xor U2465 (N_2465,N_2363,N_2344);
and U2466 (N_2466,N_2178,N_2294);
or U2467 (N_2467,In_1646,In_2249);
nand U2468 (N_2468,N_2233,In_2236);
nand U2469 (N_2469,N_2381,N_1346);
nand U2470 (N_2470,N_2303,N_2194);
or U2471 (N_2471,N_103,N_1894);
xnor U2472 (N_2472,N_1023,N_2330);
or U2473 (N_2473,N_2133,N_2186);
or U2474 (N_2474,N_2295,N_994);
nand U2475 (N_2475,N_2144,N_1626);
or U2476 (N_2476,N_768,N_1815);
or U2477 (N_2477,N_538,N_2200);
nor U2478 (N_2478,N_2121,N_1811);
and U2479 (N_2479,N_2343,N_1472);
and U2480 (N_2480,N_2281,N_2111);
nand U2481 (N_2481,N_1553,N_2279);
or U2482 (N_2482,N_2212,N_2013);
or U2483 (N_2483,N_2341,N_2373);
xnor U2484 (N_2484,In_1382,N_2278);
xor U2485 (N_2485,N_2165,N_1862);
or U2486 (N_2486,N_2167,N_52);
nor U2487 (N_2487,N_2280,N_158);
nor U2488 (N_2488,N_749,N_1664);
xnor U2489 (N_2489,N_2350,N_2263);
and U2490 (N_2490,N_2202,N_1083);
xor U2491 (N_2491,N_2132,N_2175);
xor U2492 (N_2492,In_1098,N_1835);
nand U2493 (N_2493,N_1889,N_1126);
xnor U2494 (N_2494,N_2390,N_2354);
or U2495 (N_2495,N_973,N_2395);
nand U2496 (N_2496,N_1786,N_2257);
nand U2497 (N_2497,N_1455,N_1658);
and U2498 (N_2498,N_2226,N_983);
and U2499 (N_2499,N_2374,N_2170);
or U2500 (N_2500,N_2214,N_2247);
or U2501 (N_2501,N_1266,N_2399);
nand U2502 (N_2502,N_2191,N_229);
nor U2503 (N_2503,N_2162,In_2286);
nand U2504 (N_2504,In_2041,N_2034);
or U2505 (N_2505,N_1622,N_1059);
nor U2506 (N_2506,N_2180,N_1993);
nor U2507 (N_2507,N_2313,In_1211);
and U2508 (N_2508,N_2044,In_951);
or U2509 (N_2509,In_1813,N_2135);
nand U2510 (N_2510,N_1948,N_2179);
nand U2511 (N_2511,N_2123,N_2266);
xor U2512 (N_2512,N_2393,N_1079);
or U2513 (N_2513,In_137,In_1401);
xnor U2514 (N_2514,N_2215,N_1997);
and U2515 (N_2515,N_1478,N_1912);
and U2516 (N_2516,N_1725,N_2203);
and U2517 (N_2517,N_2122,N_2310);
nor U2518 (N_2518,N_2240,In_677);
and U2519 (N_2519,N_1540,N_2108);
or U2520 (N_2520,N_1467,In_79);
or U2521 (N_2521,N_2338,N_2297);
xor U2522 (N_2522,N_2103,N_2093);
and U2523 (N_2523,N_1049,N_753);
nand U2524 (N_2524,N_321,N_1471);
and U2525 (N_2525,In_1761,N_2296);
nor U2526 (N_2526,N_2317,N_2358);
nand U2527 (N_2527,N_2092,N_2142);
xor U2528 (N_2528,N_2198,N_2286);
or U2529 (N_2529,N_1899,N_2130);
nand U2530 (N_2530,N_2288,N_2392);
nand U2531 (N_2531,N_1537,N_2207);
nand U2532 (N_2532,N_2246,N_2290);
xnor U2533 (N_2533,N_2128,N_2148);
nand U2534 (N_2534,N_2160,In_2803);
xnor U2535 (N_2535,N_2264,N_2361);
and U2536 (N_2536,N_2020,N_1744);
and U2537 (N_2537,N_2154,N_1424);
and U2538 (N_2538,N_2183,N_2291);
nor U2539 (N_2539,N_2321,N_2376);
and U2540 (N_2540,N_2176,N_2057);
nand U2541 (N_2541,N_1774,N_2378);
and U2542 (N_2542,In_845,N_2222);
or U2543 (N_2543,In_280,In_702);
and U2544 (N_2544,N_2232,N_2342);
nand U2545 (N_2545,N_1054,N_2253);
nor U2546 (N_2546,N_2213,N_2353);
nor U2547 (N_2547,In_73,N_2208);
nand U2548 (N_2548,N_2055,N_1709);
and U2549 (N_2549,N_2243,N_2388);
or U2550 (N_2550,N_94,N_2269);
and U2551 (N_2551,In_2502,In_1015);
nor U2552 (N_2552,In_2617,N_2038);
or U2553 (N_2553,N_1910,N_2324);
and U2554 (N_2554,N_1743,N_2367);
nand U2555 (N_2555,N_2315,N_1842);
or U2556 (N_2556,N_20,In_5);
nor U2557 (N_2557,In_2546,N_701);
and U2558 (N_2558,N_2349,N_1702);
or U2559 (N_2559,N_720,N_2267);
or U2560 (N_2560,N_1527,N_2220);
nor U2561 (N_2561,In_2206,N_1575);
nand U2562 (N_2562,N_2125,N_884);
xnor U2563 (N_2563,N_2328,N_1978);
xnor U2564 (N_2564,In_2751,N_734);
nand U2565 (N_2565,N_2134,In_2164);
nand U2566 (N_2566,N_2141,N_1984);
and U2567 (N_2567,N_1947,N_2357);
xnor U2568 (N_2568,N_1949,N_2152);
nor U2569 (N_2569,N_2270,N_2261);
or U2570 (N_2570,N_2386,N_412);
nand U2571 (N_2571,N_1679,N_1551);
or U2572 (N_2572,N_2150,N_1879);
and U2573 (N_2573,N_1642,N_1922);
nand U2574 (N_2574,N_675,N_1627);
nand U2575 (N_2575,N_1966,N_1416);
xnor U2576 (N_2576,N_1685,In_2967);
xnor U2577 (N_2577,N_2101,In_2022);
or U2578 (N_2578,N_2137,N_2120);
xor U2579 (N_2579,N_1452,N_2371);
nand U2580 (N_2580,N_1882,N_1970);
nand U2581 (N_2581,N_1404,N_1845);
or U2582 (N_2582,N_2217,N_2314);
nor U2583 (N_2583,N_2221,N_2231);
nand U2584 (N_2584,In_2105,N_1328);
nand U2585 (N_2585,N_1930,N_2337);
or U2586 (N_2586,N_1270,N_2308);
nor U2587 (N_2587,N_2254,N_2320);
or U2588 (N_2588,N_168,N_2129);
nand U2589 (N_2589,N_2118,N_2115);
nand U2590 (N_2590,N_2117,N_1989);
nor U2591 (N_2591,N_2197,N_1507);
or U2592 (N_2592,N_2322,N_1640);
nor U2593 (N_2593,In_1538,N_1937);
nor U2594 (N_2594,N_2241,In_1590);
and U2595 (N_2595,N_725,N_1850);
and U2596 (N_2596,N_278,N_2394);
xnor U2597 (N_2597,N_2192,In_1312);
xnor U2598 (N_2598,N_2351,N_1726);
nor U2599 (N_2599,In_2641,N_2369);
or U2600 (N_2600,N_2384,N_2382);
nor U2601 (N_2601,N_2352,In_243);
or U2602 (N_2602,N_1674,N_1775);
and U2603 (N_2603,N_2204,N_2346);
and U2604 (N_2604,N_2171,N_2287);
and U2605 (N_2605,N_2228,N_2223);
nand U2606 (N_2606,N_2318,N_2237);
nand U2607 (N_2607,N_1861,In_713);
or U2608 (N_2608,N_1820,In_1539);
xnor U2609 (N_2609,In_1848,N_2049);
nor U2610 (N_2610,N_1976,N_1926);
and U2611 (N_2611,N_2260,N_2383);
xor U2612 (N_2612,N_2190,In_2735);
or U2613 (N_2613,N_2302,N_2181);
nor U2614 (N_2614,N_2271,N_2199);
or U2615 (N_2615,N_1570,N_2206);
nand U2616 (N_2616,N_1921,N_2249);
or U2617 (N_2617,N_2274,N_1893);
nand U2618 (N_2618,N_84,N_854);
nand U2619 (N_2619,N_2301,N_1794);
nand U2620 (N_2620,N_2100,N_2276);
nand U2621 (N_2621,N_1928,In_1629);
nor U2622 (N_2622,N_1999,N_1957);
or U2623 (N_2623,N_2282,N_847);
xor U2624 (N_2624,N_2312,N_1620);
nand U2625 (N_2625,N_2250,N_2304);
nand U2626 (N_2626,N_2333,N_2139);
and U2627 (N_2627,N_2316,N_2177);
nand U2628 (N_2628,N_2104,N_2397);
xor U2629 (N_2629,N_2244,N_2109);
or U2630 (N_2630,N_1174,N_2292);
nor U2631 (N_2631,N_2097,N_2380);
nor U2632 (N_2632,In_2758,N_1028);
nand U2633 (N_2633,N_2258,N_2345);
nand U2634 (N_2634,N_1996,N_722);
nand U2635 (N_2635,N_1468,N_2230);
nand U2636 (N_2636,N_2110,N_1022);
or U2637 (N_2637,N_1701,N_1929);
nand U2638 (N_2638,N_2379,N_2275);
nand U2639 (N_2639,N_1826,N_1171);
or U2640 (N_2640,N_2158,N_2396);
or U2641 (N_2641,N_2116,N_2238);
nand U2642 (N_2642,N_2209,N_2298);
and U2643 (N_2643,N_2112,N_1789);
and U2644 (N_2644,N_2360,N_2131);
nor U2645 (N_2645,N_2336,N_2107);
nand U2646 (N_2646,N_2105,N_1829);
or U2647 (N_2647,N_2156,N_2347);
xnor U2648 (N_2648,In_2522,N_2218);
and U2649 (N_2649,N_2068,In_357);
or U2650 (N_2650,N_1173,N_1667);
xnor U2651 (N_2651,In_2784,N_2195);
or U2652 (N_2652,N_1961,N_1872);
xnor U2653 (N_2653,N_1840,N_1753);
nand U2654 (N_2654,N_2326,N_2283);
or U2655 (N_2655,N_2042,N_1866);
xor U2656 (N_2656,N_570,N_1300);
and U2657 (N_2657,N_2184,N_932);
xor U2658 (N_2658,N_1635,N_2225);
xor U2659 (N_2659,N_2293,N_2166);
nand U2660 (N_2660,N_485,In_2351);
or U2661 (N_2661,In_2730,N_2385);
nand U2662 (N_2662,N_2193,N_1802);
nor U2663 (N_2663,N_2355,N_2248);
nand U2664 (N_2664,In_2832,N_2259);
nor U2665 (N_2665,N_1722,N_2372);
or U2666 (N_2666,N_2151,N_2339);
and U2667 (N_2667,N_2368,In_1023);
xnor U2668 (N_2668,N_931,N_2289);
and U2669 (N_2669,N_2229,In_2600);
or U2670 (N_2670,N_2030,N_1819);
xnor U2671 (N_2671,N_2174,In_460);
xor U2672 (N_2672,N_2216,N_2219);
or U2673 (N_2673,N_1648,N_1438);
and U2674 (N_2674,N_700,N_2155);
nand U2675 (N_2675,N_1971,In_376);
xor U2676 (N_2676,N_1729,N_1898);
xor U2677 (N_2677,N_1697,In_1873);
or U2678 (N_2678,N_656,N_147);
xnor U2679 (N_2679,In_1388,N_1747);
nand U2680 (N_2680,N_2196,In_1946);
and U2681 (N_2681,N_2335,N_2082);
or U2682 (N_2682,N_2113,N_2268);
nor U2683 (N_2683,N_2102,N_1963);
nand U2684 (N_2684,N_1896,N_2138);
nand U2685 (N_2685,N_2327,In_933);
nor U2686 (N_2686,N_2362,In_2524);
and U2687 (N_2687,N_2127,N_2205);
nor U2688 (N_2688,N_2126,N_2153);
nor U2689 (N_2689,N_2149,N_2273);
or U2690 (N_2690,N_2236,N_1663);
and U2691 (N_2691,N_812,N_2325);
nor U2692 (N_2692,N_2359,N_2187);
nand U2693 (N_2693,In_146,N_2169);
xor U2694 (N_2694,In_2776,N_2306);
or U2695 (N_2695,N_1975,N_2235);
or U2696 (N_2696,N_1599,N_2172);
nor U2697 (N_2697,N_2242,N_1833);
xor U2698 (N_2698,N_2389,N_2272);
or U2699 (N_2699,N_1868,N_2224);
nor U2700 (N_2700,N_2535,N_2655);
xor U2701 (N_2701,N_2558,N_2493);
and U2702 (N_2702,N_2433,N_2657);
and U2703 (N_2703,N_2568,N_2596);
or U2704 (N_2704,N_2446,N_2414);
or U2705 (N_2705,N_2450,N_2503);
xor U2706 (N_2706,N_2653,N_2511);
nand U2707 (N_2707,N_2483,N_2530);
nand U2708 (N_2708,N_2420,N_2679);
xor U2709 (N_2709,N_2622,N_2667);
nand U2710 (N_2710,N_2510,N_2630);
nand U2711 (N_2711,N_2699,N_2520);
nor U2712 (N_2712,N_2545,N_2532);
xnor U2713 (N_2713,N_2424,N_2557);
nor U2714 (N_2714,N_2439,N_2482);
or U2715 (N_2715,N_2475,N_2467);
nor U2716 (N_2716,N_2489,N_2683);
nor U2717 (N_2717,N_2636,N_2539);
nand U2718 (N_2718,N_2518,N_2624);
and U2719 (N_2719,N_2650,N_2675);
nand U2720 (N_2720,N_2544,N_2674);
or U2721 (N_2721,N_2517,N_2639);
xor U2722 (N_2722,N_2481,N_2434);
and U2723 (N_2723,N_2419,N_2500);
and U2724 (N_2724,N_2522,N_2519);
and U2725 (N_2725,N_2549,N_2660);
or U2726 (N_2726,N_2637,N_2688);
or U2727 (N_2727,N_2432,N_2437);
and U2728 (N_2728,N_2413,N_2560);
or U2729 (N_2729,N_2659,N_2646);
or U2730 (N_2730,N_2598,N_2571);
nor U2731 (N_2731,N_2572,N_2612);
or U2732 (N_2732,N_2595,N_2526);
nand U2733 (N_2733,N_2480,N_2603);
nor U2734 (N_2734,N_2471,N_2602);
nor U2735 (N_2735,N_2425,N_2628);
or U2736 (N_2736,N_2634,N_2491);
and U2737 (N_2737,N_2690,N_2554);
or U2738 (N_2738,N_2421,N_2502);
nand U2739 (N_2739,N_2696,N_2469);
nor U2740 (N_2740,N_2626,N_2508);
nor U2741 (N_2741,N_2618,N_2490);
nor U2742 (N_2742,N_2548,N_2627);
xnor U2743 (N_2743,N_2487,N_2542);
nor U2744 (N_2744,N_2666,N_2463);
nand U2745 (N_2745,N_2400,N_2547);
nor U2746 (N_2746,N_2577,N_2476);
xor U2747 (N_2747,N_2609,N_2497);
xnor U2748 (N_2748,N_2524,N_2582);
nand U2749 (N_2749,N_2606,N_2431);
and U2750 (N_2750,N_2691,N_2640);
or U2751 (N_2751,N_2623,N_2440);
nor U2752 (N_2752,N_2682,N_2485);
and U2753 (N_2753,N_2589,N_2460);
nor U2754 (N_2754,N_2405,N_2677);
nand U2755 (N_2755,N_2513,N_2562);
or U2756 (N_2756,N_2470,N_2583);
nand U2757 (N_2757,N_2496,N_2629);
nand U2758 (N_2758,N_2694,N_2506);
or U2759 (N_2759,N_2617,N_2473);
xnor U2760 (N_2760,N_2417,N_2680);
xor U2761 (N_2761,N_2403,N_2587);
or U2762 (N_2762,N_2592,N_2649);
or U2763 (N_2763,N_2527,N_2507);
nor U2764 (N_2764,N_2418,N_2515);
nor U2765 (N_2765,N_2559,N_2692);
xor U2766 (N_2766,N_2436,N_2590);
nor U2767 (N_2767,N_2455,N_2474);
nand U2768 (N_2768,N_2406,N_2564);
nand U2769 (N_2769,N_2631,N_2468);
nor U2770 (N_2770,N_2614,N_2448);
xor U2771 (N_2771,N_2563,N_2625);
nand U2772 (N_2772,N_2600,N_2556);
xnor U2773 (N_2773,N_2408,N_2578);
and U2774 (N_2774,N_2427,N_2575);
nand U2775 (N_2775,N_2642,N_2525);
and U2776 (N_2776,N_2415,N_2494);
nand U2777 (N_2777,N_2528,N_2457);
nand U2778 (N_2778,N_2697,N_2435);
nor U2779 (N_2779,N_2607,N_2635);
and U2780 (N_2780,N_2536,N_2576);
or U2781 (N_2781,N_2512,N_2404);
nor U2782 (N_2782,N_2426,N_2488);
or U2783 (N_2783,N_2671,N_2505);
nand U2784 (N_2784,N_2477,N_2462);
xor U2785 (N_2785,N_2654,N_2591);
nor U2786 (N_2786,N_2501,N_2584);
nand U2787 (N_2787,N_2401,N_2565);
nor U2788 (N_2788,N_2521,N_2566);
nor U2789 (N_2789,N_2423,N_2543);
nor U2790 (N_2790,N_2541,N_2581);
and U2791 (N_2791,N_2676,N_2416);
nor U2792 (N_2792,N_2597,N_2540);
xnor U2793 (N_2793,N_2686,N_2593);
and U2794 (N_2794,N_2644,N_2689);
or U2795 (N_2795,N_2656,N_2523);
or U2796 (N_2796,N_2454,N_2537);
and U2797 (N_2797,N_2601,N_2464);
nand U2798 (N_2798,N_2407,N_2531);
and U2799 (N_2799,N_2453,N_2402);
nand U2800 (N_2800,N_2621,N_2638);
nor U2801 (N_2801,N_2615,N_2410);
nand U2802 (N_2802,N_2461,N_2573);
xor U2803 (N_2803,N_2668,N_2672);
and U2804 (N_2804,N_2599,N_2498);
or U2805 (N_2805,N_2611,N_2447);
xnor U2806 (N_2806,N_2579,N_2588);
nand U2807 (N_2807,N_2445,N_2553);
xnor U2808 (N_2808,N_2438,N_2459);
nand U2809 (N_2809,N_2516,N_2685);
or U2810 (N_2810,N_2669,N_2484);
nor U2811 (N_2811,N_2651,N_2452);
nor U2812 (N_2812,N_2570,N_2665);
and U2813 (N_2813,N_2604,N_2580);
and U2814 (N_2814,N_2687,N_2495);
xnor U2815 (N_2815,N_2693,N_2546);
and U2816 (N_2816,N_2661,N_2529);
xnor U2817 (N_2817,N_2514,N_2633);
and U2818 (N_2818,N_2613,N_2662);
or U2819 (N_2819,N_2632,N_2533);
nor U2820 (N_2820,N_2586,N_2479);
and U2821 (N_2821,N_2443,N_2678);
and U2822 (N_2822,N_2673,N_2670);
nor U2823 (N_2823,N_2616,N_2648);
nor U2824 (N_2824,N_2534,N_2422);
and U2825 (N_2825,N_2429,N_2478);
and U2826 (N_2826,N_2663,N_2647);
and U2827 (N_2827,N_2574,N_2610);
nand U2828 (N_2828,N_2451,N_2698);
nor U2829 (N_2829,N_2550,N_2695);
nor U2830 (N_2830,N_2641,N_2585);
nor U2831 (N_2831,N_2552,N_2412);
nand U2832 (N_2832,N_2684,N_2486);
or U2833 (N_2833,N_2608,N_2472);
or U2834 (N_2834,N_2409,N_2444);
xor U2835 (N_2835,N_2652,N_2428);
or U2836 (N_2836,N_2465,N_2411);
nor U2837 (N_2837,N_2555,N_2551);
and U2838 (N_2838,N_2645,N_2538);
and U2839 (N_2839,N_2620,N_2449);
xnor U2840 (N_2840,N_2504,N_2681);
xor U2841 (N_2841,N_2658,N_2561);
xor U2842 (N_2842,N_2466,N_2619);
xnor U2843 (N_2843,N_2594,N_2605);
and U2844 (N_2844,N_2442,N_2441);
xnor U2845 (N_2845,N_2458,N_2569);
xnor U2846 (N_2846,N_2567,N_2509);
nor U2847 (N_2847,N_2499,N_2492);
xor U2848 (N_2848,N_2456,N_2664);
and U2849 (N_2849,N_2643,N_2430);
nand U2850 (N_2850,N_2530,N_2531);
nand U2851 (N_2851,N_2400,N_2409);
xor U2852 (N_2852,N_2518,N_2446);
and U2853 (N_2853,N_2651,N_2699);
and U2854 (N_2854,N_2460,N_2521);
xnor U2855 (N_2855,N_2515,N_2613);
and U2856 (N_2856,N_2505,N_2410);
nand U2857 (N_2857,N_2476,N_2613);
nor U2858 (N_2858,N_2560,N_2563);
xor U2859 (N_2859,N_2584,N_2559);
nand U2860 (N_2860,N_2610,N_2453);
or U2861 (N_2861,N_2675,N_2694);
nand U2862 (N_2862,N_2573,N_2681);
or U2863 (N_2863,N_2591,N_2430);
or U2864 (N_2864,N_2518,N_2586);
nand U2865 (N_2865,N_2570,N_2603);
or U2866 (N_2866,N_2490,N_2474);
nand U2867 (N_2867,N_2631,N_2523);
and U2868 (N_2868,N_2502,N_2563);
xor U2869 (N_2869,N_2410,N_2495);
nand U2870 (N_2870,N_2448,N_2431);
nand U2871 (N_2871,N_2564,N_2412);
or U2872 (N_2872,N_2610,N_2612);
nor U2873 (N_2873,N_2522,N_2548);
xnor U2874 (N_2874,N_2406,N_2560);
and U2875 (N_2875,N_2572,N_2635);
and U2876 (N_2876,N_2669,N_2464);
and U2877 (N_2877,N_2578,N_2672);
and U2878 (N_2878,N_2418,N_2513);
and U2879 (N_2879,N_2574,N_2536);
or U2880 (N_2880,N_2650,N_2521);
or U2881 (N_2881,N_2463,N_2542);
and U2882 (N_2882,N_2423,N_2501);
nor U2883 (N_2883,N_2606,N_2598);
nor U2884 (N_2884,N_2464,N_2470);
and U2885 (N_2885,N_2506,N_2586);
nand U2886 (N_2886,N_2573,N_2472);
nand U2887 (N_2887,N_2598,N_2484);
nand U2888 (N_2888,N_2546,N_2423);
and U2889 (N_2889,N_2542,N_2530);
xnor U2890 (N_2890,N_2501,N_2434);
nand U2891 (N_2891,N_2497,N_2671);
and U2892 (N_2892,N_2552,N_2676);
xor U2893 (N_2893,N_2601,N_2660);
nor U2894 (N_2894,N_2471,N_2447);
nor U2895 (N_2895,N_2487,N_2602);
xnor U2896 (N_2896,N_2596,N_2539);
nor U2897 (N_2897,N_2592,N_2601);
xor U2898 (N_2898,N_2698,N_2682);
and U2899 (N_2899,N_2693,N_2427);
nand U2900 (N_2900,N_2509,N_2611);
and U2901 (N_2901,N_2621,N_2520);
or U2902 (N_2902,N_2492,N_2618);
xor U2903 (N_2903,N_2513,N_2659);
nand U2904 (N_2904,N_2582,N_2591);
nand U2905 (N_2905,N_2507,N_2488);
xnor U2906 (N_2906,N_2419,N_2631);
and U2907 (N_2907,N_2476,N_2650);
xnor U2908 (N_2908,N_2594,N_2568);
or U2909 (N_2909,N_2677,N_2637);
and U2910 (N_2910,N_2621,N_2676);
nor U2911 (N_2911,N_2609,N_2450);
nand U2912 (N_2912,N_2658,N_2534);
nand U2913 (N_2913,N_2480,N_2658);
xnor U2914 (N_2914,N_2561,N_2582);
nand U2915 (N_2915,N_2674,N_2635);
nand U2916 (N_2916,N_2625,N_2461);
or U2917 (N_2917,N_2406,N_2670);
nor U2918 (N_2918,N_2514,N_2676);
and U2919 (N_2919,N_2517,N_2498);
or U2920 (N_2920,N_2623,N_2683);
or U2921 (N_2921,N_2517,N_2464);
nor U2922 (N_2922,N_2574,N_2510);
nand U2923 (N_2923,N_2594,N_2514);
nor U2924 (N_2924,N_2404,N_2504);
nand U2925 (N_2925,N_2542,N_2492);
and U2926 (N_2926,N_2437,N_2583);
nand U2927 (N_2927,N_2635,N_2411);
nand U2928 (N_2928,N_2569,N_2555);
xnor U2929 (N_2929,N_2444,N_2572);
nand U2930 (N_2930,N_2600,N_2448);
xnor U2931 (N_2931,N_2651,N_2694);
nor U2932 (N_2932,N_2518,N_2409);
nor U2933 (N_2933,N_2541,N_2511);
nor U2934 (N_2934,N_2458,N_2692);
and U2935 (N_2935,N_2632,N_2430);
nand U2936 (N_2936,N_2441,N_2557);
or U2937 (N_2937,N_2534,N_2476);
or U2938 (N_2938,N_2629,N_2405);
nand U2939 (N_2939,N_2636,N_2557);
or U2940 (N_2940,N_2582,N_2450);
and U2941 (N_2941,N_2541,N_2478);
and U2942 (N_2942,N_2597,N_2579);
nand U2943 (N_2943,N_2531,N_2454);
and U2944 (N_2944,N_2683,N_2667);
xnor U2945 (N_2945,N_2513,N_2572);
nand U2946 (N_2946,N_2500,N_2606);
xnor U2947 (N_2947,N_2492,N_2573);
or U2948 (N_2948,N_2684,N_2539);
xnor U2949 (N_2949,N_2402,N_2452);
nor U2950 (N_2950,N_2525,N_2416);
xor U2951 (N_2951,N_2438,N_2421);
xnor U2952 (N_2952,N_2671,N_2429);
xnor U2953 (N_2953,N_2647,N_2449);
xnor U2954 (N_2954,N_2436,N_2415);
or U2955 (N_2955,N_2486,N_2532);
nand U2956 (N_2956,N_2547,N_2417);
nor U2957 (N_2957,N_2554,N_2613);
or U2958 (N_2958,N_2504,N_2486);
and U2959 (N_2959,N_2619,N_2523);
nor U2960 (N_2960,N_2661,N_2554);
or U2961 (N_2961,N_2507,N_2693);
nand U2962 (N_2962,N_2438,N_2629);
and U2963 (N_2963,N_2500,N_2502);
nor U2964 (N_2964,N_2474,N_2572);
xor U2965 (N_2965,N_2450,N_2694);
nand U2966 (N_2966,N_2582,N_2447);
nand U2967 (N_2967,N_2565,N_2622);
nor U2968 (N_2968,N_2561,N_2412);
nor U2969 (N_2969,N_2567,N_2462);
or U2970 (N_2970,N_2442,N_2516);
nand U2971 (N_2971,N_2500,N_2686);
nand U2972 (N_2972,N_2695,N_2611);
and U2973 (N_2973,N_2575,N_2482);
nand U2974 (N_2974,N_2446,N_2589);
nand U2975 (N_2975,N_2404,N_2446);
and U2976 (N_2976,N_2484,N_2594);
nand U2977 (N_2977,N_2418,N_2540);
nor U2978 (N_2978,N_2561,N_2521);
and U2979 (N_2979,N_2611,N_2437);
nor U2980 (N_2980,N_2442,N_2679);
or U2981 (N_2981,N_2478,N_2525);
or U2982 (N_2982,N_2485,N_2622);
nand U2983 (N_2983,N_2558,N_2415);
nor U2984 (N_2984,N_2419,N_2437);
or U2985 (N_2985,N_2607,N_2667);
and U2986 (N_2986,N_2636,N_2637);
nand U2987 (N_2987,N_2643,N_2512);
and U2988 (N_2988,N_2671,N_2442);
and U2989 (N_2989,N_2517,N_2574);
or U2990 (N_2990,N_2628,N_2525);
xor U2991 (N_2991,N_2697,N_2671);
xnor U2992 (N_2992,N_2444,N_2690);
nor U2993 (N_2993,N_2530,N_2676);
or U2994 (N_2994,N_2693,N_2535);
and U2995 (N_2995,N_2446,N_2645);
nand U2996 (N_2996,N_2662,N_2661);
nor U2997 (N_2997,N_2596,N_2613);
nand U2998 (N_2998,N_2697,N_2592);
or U2999 (N_2999,N_2627,N_2637);
xnor U3000 (N_3000,N_2879,N_2811);
nand U3001 (N_3001,N_2702,N_2808);
and U3002 (N_3002,N_2777,N_2883);
and U3003 (N_3003,N_2706,N_2867);
or U3004 (N_3004,N_2926,N_2701);
nand U3005 (N_3005,N_2875,N_2866);
xor U3006 (N_3006,N_2742,N_2954);
xor U3007 (N_3007,N_2748,N_2959);
or U3008 (N_3008,N_2878,N_2714);
nor U3009 (N_3009,N_2924,N_2919);
and U3010 (N_3010,N_2884,N_2915);
or U3011 (N_3011,N_2792,N_2759);
nor U3012 (N_3012,N_2882,N_2910);
nand U3013 (N_3013,N_2781,N_2987);
xor U3014 (N_3014,N_2881,N_2846);
nand U3015 (N_3015,N_2942,N_2906);
nand U3016 (N_3016,N_2946,N_2757);
and U3017 (N_3017,N_2817,N_2780);
nand U3018 (N_3018,N_2952,N_2752);
nand U3019 (N_3019,N_2833,N_2857);
or U3020 (N_3020,N_2912,N_2718);
or U3021 (N_3021,N_2859,N_2813);
xor U3022 (N_3022,N_2704,N_2730);
xor U3023 (N_3023,N_2711,N_2843);
nor U3024 (N_3024,N_2838,N_2986);
nor U3025 (N_3025,N_2799,N_2904);
xnor U3026 (N_3026,N_2767,N_2963);
and U3027 (N_3027,N_2880,N_2970);
and U3028 (N_3028,N_2864,N_2721);
or U3029 (N_3029,N_2788,N_2708);
xor U3030 (N_3030,N_2796,N_2933);
xnor U3031 (N_3031,N_2950,N_2802);
and U3032 (N_3032,N_2705,N_2839);
or U3033 (N_3033,N_2732,N_2888);
and U3034 (N_3034,N_2819,N_2871);
or U3035 (N_3035,N_2897,N_2984);
and U3036 (N_3036,N_2981,N_2887);
xnor U3037 (N_3037,N_2971,N_2991);
xor U3038 (N_3038,N_2768,N_2929);
or U3039 (N_3039,N_2840,N_2961);
nand U3040 (N_3040,N_2725,N_2921);
and U3041 (N_3041,N_2820,N_2724);
nand U3042 (N_3042,N_2974,N_2823);
nand U3043 (N_3043,N_2927,N_2824);
xnor U3044 (N_3044,N_2737,N_2918);
nor U3045 (N_3045,N_2898,N_2922);
and U3046 (N_3046,N_2789,N_2966);
and U3047 (N_3047,N_2791,N_2993);
or U3048 (N_3048,N_2896,N_2903);
or U3049 (N_3049,N_2814,N_2821);
xor U3050 (N_3050,N_2745,N_2995);
and U3051 (N_3051,N_2837,N_2766);
nor U3052 (N_3052,N_2805,N_2720);
nand U3053 (N_3053,N_2928,N_2723);
or U3054 (N_3054,N_2938,N_2743);
and U3055 (N_3055,N_2769,N_2907);
xnor U3056 (N_3056,N_2877,N_2944);
nand U3057 (N_3057,N_2914,N_2947);
nor U3058 (N_3058,N_2822,N_2795);
nand U3059 (N_3059,N_2889,N_2832);
and U3060 (N_3060,N_2847,N_2932);
or U3061 (N_3061,N_2960,N_2800);
nor U3062 (N_3062,N_2784,N_2749);
or U3063 (N_3063,N_2983,N_2809);
nand U3064 (N_3064,N_2873,N_2764);
and U3065 (N_3065,N_2774,N_2707);
or U3066 (N_3066,N_2958,N_2943);
xor U3067 (N_3067,N_2850,N_2801);
and U3068 (N_3068,N_2710,N_2747);
nor U3069 (N_3069,N_2951,N_2853);
nor U3070 (N_3070,N_2890,N_2876);
nand U3071 (N_3071,N_2856,N_2962);
nand U3072 (N_3072,N_2729,N_2739);
nand U3073 (N_3073,N_2715,N_2977);
xor U3074 (N_3074,N_2980,N_2936);
nand U3075 (N_3075,N_2787,N_2865);
and U3076 (N_3076,N_2999,N_2778);
xnor U3077 (N_3077,N_2783,N_2753);
or U3078 (N_3078,N_2874,N_2863);
xor U3079 (N_3079,N_2978,N_2967);
nand U3080 (N_3080,N_2803,N_2841);
xor U3081 (N_3081,N_2899,N_2770);
nand U3082 (N_3082,N_2937,N_2949);
nor U3083 (N_3083,N_2858,N_2891);
nand U3084 (N_3084,N_2860,N_2964);
or U3085 (N_3085,N_2760,N_2996);
nor U3086 (N_3086,N_2852,N_2893);
or U3087 (N_3087,N_2908,N_2969);
nor U3088 (N_3088,N_2761,N_2975);
or U3089 (N_3089,N_2754,N_2731);
and U3090 (N_3090,N_2741,N_2826);
nor U3091 (N_3091,N_2793,N_2712);
xnor U3092 (N_3092,N_2744,N_2807);
nor U3093 (N_3093,N_2968,N_2930);
or U3094 (N_3094,N_2940,N_2998);
and U3095 (N_3095,N_2939,N_2709);
xor U3096 (N_3096,N_2935,N_2872);
xor U3097 (N_3097,N_2772,N_2941);
and U3098 (N_3098,N_2869,N_2804);
nand U3099 (N_3099,N_2909,N_2786);
and U3100 (N_3100,N_2797,N_2756);
or U3101 (N_3101,N_2886,N_2994);
nor U3102 (N_3102,N_2901,N_2776);
and U3103 (N_3103,N_2955,N_2989);
and U3104 (N_3104,N_2845,N_2844);
and U3105 (N_3105,N_2785,N_2920);
xor U3106 (N_3106,N_2990,N_2746);
or U3107 (N_3107,N_2816,N_2700);
or U3108 (N_3108,N_2957,N_2894);
or U3109 (N_3109,N_2735,N_2728);
or U3110 (N_3110,N_2762,N_2733);
or U3111 (N_3111,N_2719,N_2885);
xor U3112 (N_3112,N_2985,N_2758);
nor U3113 (N_3113,N_2988,N_2842);
and U3114 (N_3114,N_2854,N_2848);
nor U3115 (N_3115,N_2790,N_2779);
xnor U3116 (N_3116,N_2972,N_2925);
xor U3117 (N_3117,N_2782,N_2818);
xnor U3118 (N_3118,N_2827,N_2763);
and U3119 (N_3119,N_2750,N_2849);
and U3120 (N_3120,N_2836,N_2895);
xnor U3121 (N_3121,N_2851,N_2870);
nor U3122 (N_3122,N_2734,N_2953);
nand U3123 (N_3123,N_2911,N_2855);
xnor U3124 (N_3124,N_2794,N_2726);
xnor U3125 (N_3125,N_2830,N_2703);
or U3126 (N_3126,N_2965,N_2979);
nor U3127 (N_3127,N_2765,N_2755);
and U3128 (N_3128,N_2976,N_2740);
nand U3129 (N_3129,N_2900,N_2917);
xnor U3130 (N_3130,N_2923,N_2831);
nand U3131 (N_3131,N_2773,N_2861);
nor U3132 (N_3132,N_2913,N_2997);
or U3133 (N_3133,N_2956,N_2931);
nor U3134 (N_3134,N_2982,N_2713);
nor U3135 (N_3135,N_2973,N_2916);
or U3136 (N_3136,N_2812,N_2892);
nand U3137 (N_3137,N_2810,N_2945);
and U3138 (N_3138,N_2738,N_2862);
nand U3139 (N_3139,N_2868,N_2751);
and U3140 (N_3140,N_2902,N_2825);
nor U3141 (N_3141,N_2727,N_2736);
nand U3142 (N_3142,N_2829,N_2722);
xnor U3143 (N_3143,N_2828,N_2934);
and U3144 (N_3144,N_2815,N_2948);
nor U3145 (N_3145,N_2716,N_2835);
or U3146 (N_3146,N_2798,N_2992);
or U3147 (N_3147,N_2834,N_2905);
and U3148 (N_3148,N_2775,N_2717);
and U3149 (N_3149,N_2806,N_2771);
and U3150 (N_3150,N_2764,N_2872);
or U3151 (N_3151,N_2772,N_2768);
nor U3152 (N_3152,N_2724,N_2843);
or U3153 (N_3153,N_2838,N_2895);
nor U3154 (N_3154,N_2758,N_2936);
nor U3155 (N_3155,N_2712,N_2987);
nand U3156 (N_3156,N_2869,N_2844);
or U3157 (N_3157,N_2994,N_2950);
and U3158 (N_3158,N_2833,N_2723);
or U3159 (N_3159,N_2811,N_2888);
and U3160 (N_3160,N_2896,N_2757);
nor U3161 (N_3161,N_2876,N_2830);
nor U3162 (N_3162,N_2753,N_2917);
and U3163 (N_3163,N_2766,N_2956);
nand U3164 (N_3164,N_2756,N_2818);
and U3165 (N_3165,N_2971,N_2868);
and U3166 (N_3166,N_2935,N_2722);
nor U3167 (N_3167,N_2913,N_2701);
nand U3168 (N_3168,N_2867,N_2942);
nand U3169 (N_3169,N_2891,N_2702);
or U3170 (N_3170,N_2956,N_2923);
or U3171 (N_3171,N_2941,N_2770);
or U3172 (N_3172,N_2711,N_2752);
nand U3173 (N_3173,N_2933,N_2883);
nor U3174 (N_3174,N_2731,N_2948);
and U3175 (N_3175,N_2782,N_2866);
xnor U3176 (N_3176,N_2997,N_2742);
or U3177 (N_3177,N_2738,N_2835);
xnor U3178 (N_3178,N_2853,N_2919);
nand U3179 (N_3179,N_2966,N_2711);
nand U3180 (N_3180,N_2915,N_2847);
or U3181 (N_3181,N_2906,N_2853);
and U3182 (N_3182,N_2858,N_2925);
and U3183 (N_3183,N_2905,N_2913);
and U3184 (N_3184,N_2740,N_2973);
nand U3185 (N_3185,N_2900,N_2845);
or U3186 (N_3186,N_2842,N_2875);
xor U3187 (N_3187,N_2971,N_2853);
xor U3188 (N_3188,N_2924,N_2889);
or U3189 (N_3189,N_2977,N_2951);
or U3190 (N_3190,N_2722,N_2922);
nor U3191 (N_3191,N_2937,N_2980);
nand U3192 (N_3192,N_2932,N_2969);
nand U3193 (N_3193,N_2871,N_2824);
or U3194 (N_3194,N_2888,N_2912);
nor U3195 (N_3195,N_2787,N_2842);
nor U3196 (N_3196,N_2902,N_2731);
or U3197 (N_3197,N_2723,N_2885);
and U3198 (N_3198,N_2855,N_2894);
nand U3199 (N_3199,N_2985,N_2744);
and U3200 (N_3200,N_2788,N_2973);
or U3201 (N_3201,N_2970,N_2810);
or U3202 (N_3202,N_2819,N_2944);
or U3203 (N_3203,N_2993,N_2737);
or U3204 (N_3204,N_2736,N_2992);
and U3205 (N_3205,N_2709,N_2774);
and U3206 (N_3206,N_2962,N_2963);
xor U3207 (N_3207,N_2877,N_2703);
xor U3208 (N_3208,N_2884,N_2787);
nand U3209 (N_3209,N_2879,N_2744);
nor U3210 (N_3210,N_2962,N_2871);
and U3211 (N_3211,N_2849,N_2888);
and U3212 (N_3212,N_2729,N_2791);
nand U3213 (N_3213,N_2923,N_2919);
and U3214 (N_3214,N_2798,N_2789);
nand U3215 (N_3215,N_2811,N_2980);
nand U3216 (N_3216,N_2736,N_2833);
or U3217 (N_3217,N_2747,N_2740);
and U3218 (N_3218,N_2926,N_2934);
nor U3219 (N_3219,N_2816,N_2825);
or U3220 (N_3220,N_2929,N_2773);
nor U3221 (N_3221,N_2897,N_2835);
nand U3222 (N_3222,N_2961,N_2754);
or U3223 (N_3223,N_2916,N_2733);
xor U3224 (N_3224,N_2803,N_2773);
nand U3225 (N_3225,N_2918,N_2793);
nor U3226 (N_3226,N_2758,N_2760);
xor U3227 (N_3227,N_2990,N_2925);
xor U3228 (N_3228,N_2738,N_2859);
xor U3229 (N_3229,N_2846,N_2847);
xor U3230 (N_3230,N_2859,N_2714);
nand U3231 (N_3231,N_2717,N_2796);
xor U3232 (N_3232,N_2926,N_2788);
xnor U3233 (N_3233,N_2914,N_2987);
xnor U3234 (N_3234,N_2888,N_2893);
or U3235 (N_3235,N_2928,N_2890);
and U3236 (N_3236,N_2913,N_2741);
or U3237 (N_3237,N_2952,N_2889);
and U3238 (N_3238,N_2711,N_2900);
and U3239 (N_3239,N_2801,N_2819);
and U3240 (N_3240,N_2701,N_2795);
xnor U3241 (N_3241,N_2960,N_2766);
nor U3242 (N_3242,N_2963,N_2794);
nand U3243 (N_3243,N_2834,N_2790);
xor U3244 (N_3244,N_2840,N_2764);
nand U3245 (N_3245,N_2903,N_2715);
and U3246 (N_3246,N_2711,N_2862);
nor U3247 (N_3247,N_2731,N_2932);
or U3248 (N_3248,N_2937,N_2759);
nand U3249 (N_3249,N_2938,N_2913);
and U3250 (N_3250,N_2828,N_2855);
xor U3251 (N_3251,N_2831,N_2943);
nand U3252 (N_3252,N_2812,N_2744);
xor U3253 (N_3253,N_2743,N_2795);
nand U3254 (N_3254,N_2790,N_2945);
xnor U3255 (N_3255,N_2979,N_2828);
and U3256 (N_3256,N_2933,N_2781);
and U3257 (N_3257,N_2837,N_2971);
nand U3258 (N_3258,N_2939,N_2702);
nand U3259 (N_3259,N_2920,N_2991);
nor U3260 (N_3260,N_2943,N_2769);
or U3261 (N_3261,N_2911,N_2790);
or U3262 (N_3262,N_2962,N_2850);
nor U3263 (N_3263,N_2872,N_2949);
xnor U3264 (N_3264,N_2774,N_2916);
nand U3265 (N_3265,N_2825,N_2968);
nand U3266 (N_3266,N_2877,N_2875);
and U3267 (N_3267,N_2948,N_2712);
nand U3268 (N_3268,N_2935,N_2869);
or U3269 (N_3269,N_2958,N_2977);
and U3270 (N_3270,N_2966,N_2797);
nor U3271 (N_3271,N_2984,N_2817);
or U3272 (N_3272,N_2799,N_2930);
xor U3273 (N_3273,N_2785,N_2759);
nand U3274 (N_3274,N_2876,N_2715);
xnor U3275 (N_3275,N_2930,N_2868);
or U3276 (N_3276,N_2954,N_2996);
xnor U3277 (N_3277,N_2808,N_2858);
nor U3278 (N_3278,N_2772,N_2851);
and U3279 (N_3279,N_2989,N_2879);
nand U3280 (N_3280,N_2736,N_2762);
and U3281 (N_3281,N_2853,N_2832);
nand U3282 (N_3282,N_2790,N_2891);
nand U3283 (N_3283,N_2976,N_2991);
xnor U3284 (N_3284,N_2819,N_2767);
xor U3285 (N_3285,N_2842,N_2978);
nand U3286 (N_3286,N_2776,N_2958);
xor U3287 (N_3287,N_2837,N_2954);
nand U3288 (N_3288,N_2875,N_2814);
nor U3289 (N_3289,N_2705,N_2983);
nand U3290 (N_3290,N_2966,N_2977);
xnor U3291 (N_3291,N_2941,N_2721);
xor U3292 (N_3292,N_2727,N_2747);
nand U3293 (N_3293,N_2800,N_2994);
and U3294 (N_3294,N_2785,N_2889);
and U3295 (N_3295,N_2856,N_2996);
or U3296 (N_3296,N_2989,N_2914);
xnor U3297 (N_3297,N_2832,N_2850);
nor U3298 (N_3298,N_2984,N_2838);
or U3299 (N_3299,N_2846,N_2792);
xor U3300 (N_3300,N_3012,N_3108);
nand U3301 (N_3301,N_3250,N_3002);
and U3302 (N_3302,N_3280,N_3230);
or U3303 (N_3303,N_3198,N_3253);
or U3304 (N_3304,N_3089,N_3096);
or U3305 (N_3305,N_3080,N_3019);
nor U3306 (N_3306,N_3142,N_3136);
and U3307 (N_3307,N_3183,N_3097);
xor U3308 (N_3308,N_3286,N_3231);
nor U3309 (N_3309,N_3232,N_3299);
xnor U3310 (N_3310,N_3221,N_3157);
or U3311 (N_3311,N_3148,N_3155);
xor U3312 (N_3312,N_3113,N_3005);
xnor U3313 (N_3313,N_3125,N_3256);
or U3314 (N_3314,N_3193,N_3276);
nand U3315 (N_3315,N_3179,N_3237);
nand U3316 (N_3316,N_3199,N_3001);
and U3317 (N_3317,N_3251,N_3226);
and U3318 (N_3318,N_3249,N_3123);
nor U3319 (N_3319,N_3266,N_3078);
or U3320 (N_3320,N_3139,N_3034);
or U3321 (N_3321,N_3172,N_3118);
and U3322 (N_3322,N_3244,N_3067);
or U3323 (N_3323,N_3160,N_3072);
nor U3324 (N_3324,N_3233,N_3141);
xor U3325 (N_3325,N_3043,N_3240);
or U3326 (N_3326,N_3059,N_3079);
or U3327 (N_3327,N_3047,N_3115);
or U3328 (N_3328,N_3050,N_3098);
and U3329 (N_3329,N_3282,N_3196);
nor U3330 (N_3330,N_3051,N_3081);
or U3331 (N_3331,N_3158,N_3101);
nand U3332 (N_3332,N_3065,N_3154);
nand U3333 (N_3333,N_3246,N_3235);
or U3334 (N_3334,N_3187,N_3126);
nor U3335 (N_3335,N_3053,N_3285);
nor U3336 (N_3336,N_3049,N_3117);
nor U3337 (N_3337,N_3087,N_3074);
nand U3338 (N_3338,N_3234,N_3213);
xnor U3339 (N_3339,N_3110,N_3046);
nor U3340 (N_3340,N_3175,N_3063);
nor U3341 (N_3341,N_3182,N_3228);
or U3342 (N_3342,N_3248,N_3144);
or U3343 (N_3343,N_3243,N_3219);
xor U3344 (N_3344,N_3057,N_3014);
xor U3345 (N_3345,N_3007,N_3104);
and U3346 (N_3346,N_3298,N_3162);
nor U3347 (N_3347,N_3236,N_3190);
and U3348 (N_3348,N_3058,N_3178);
nand U3349 (N_3349,N_3060,N_3261);
xor U3350 (N_3350,N_3177,N_3024);
nand U3351 (N_3351,N_3093,N_3003);
and U3352 (N_3352,N_3090,N_3056);
and U3353 (N_3353,N_3135,N_3086);
and U3354 (N_3354,N_3044,N_3011);
nor U3355 (N_3355,N_3171,N_3062);
and U3356 (N_3356,N_3241,N_3023);
or U3357 (N_3357,N_3255,N_3119);
xnor U3358 (N_3358,N_3273,N_3132);
xnor U3359 (N_3359,N_3114,N_3208);
xor U3360 (N_3360,N_3022,N_3120);
nand U3361 (N_3361,N_3009,N_3103);
or U3362 (N_3362,N_3209,N_3018);
xor U3363 (N_3363,N_3128,N_3068);
nor U3364 (N_3364,N_3224,N_3216);
and U3365 (N_3365,N_3167,N_3165);
and U3366 (N_3366,N_3033,N_3263);
or U3367 (N_3367,N_3291,N_3279);
or U3368 (N_3368,N_3035,N_3295);
nand U3369 (N_3369,N_3166,N_3211);
nand U3370 (N_3370,N_3085,N_3017);
or U3371 (N_3371,N_3077,N_3127);
xor U3372 (N_3372,N_3073,N_3170);
xor U3373 (N_3373,N_3239,N_3100);
nand U3374 (N_3374,N_3200,N_3048);
and U3375 (N_3375,N_3297,N_3066);
and U3376 (N_3376,N_3289,N_3185);
xnor U3377 (N_3377,N_3222,N_3070);
or U3378 (N_3378,N_3025,N_3265);
xor U3379 (N_3379,N_3124,N_3064);
and U3380 (N_3380,N_3242,N_3094);
and U3381 (N_3381,N_3036,N_3076);
and U3382 (N_3382,N_3267,N_3102);
xor U3383 (N_3383,N_3122,N_3288);
and U3384 (N_3384,N_3069,N_3164);
nand U3385 (N_3385,N_3210,N_3278);
nand U3386 (N_3386,N_3109,N_3111);
xor U3387 (N_3387,N_3082,N_3192);
xnor U3388 (N_3388,N_3238,N_3262);
nor U3389 (N_3389,N_3021,N_3268);
nor U3390 (N_3390,N_3191,N_3257);
nand U3391 (N_3391,N_3112,N_3030);
nand U3392 (N_3392,N_3130,N_3099);
or U3393 (N_3393,N_3189,N_3287);
or U3394 (N_3394,N_3004,N_3174);
or U3395 (N_3395,N_3169,N_3106);
nand U3396 (N_3396,N_3054,N_3000);
or U3397 (N_3397,N_3258,N_3296);
xnor U3398 (N_3398,N_3156,N_3163);
and U3399 (N_3399,N_3283,N_3161);
or U3400 (N_3400,N_3041,N_3186);
xnor U3401 (N_3401,N_3245,N_3173);
and U3402 (N_3402,N_3181,N_3028);
and U3403 (N_3403,N_3040,N_3091);
nand U3404 (N_3404,N_3042,N_3247);
nor U3405 (N_3405,N_3252,N_3061);
or U3406 (N_3406,N_3205,N_3176);
and U3407 (N_3407,N_3052,N_3008);
xor U3408 (N_3408,N_3134,N_3277);
or U3409 (N_3409,N_3088,N_3194);
xnor U3410 (N_3410,N_3201,N_3140);
or U3411 (N_3411,N_3055,N_3197);
and U3412 (N_3412,N_3206,N_3149);
xnor U3413 (N_3413,N_3188,N_3184);
and U3414 (N_3414,N_3202,N_3281);
xnor U3415 (N_3415,N_3284,N_3152);
nand U3416 (N_3416,N_3227,N_3015);
xor U3417 (N_3417,N_3029,N_3092);
and U3418 (N_3418,N_3269,N_3032);
nor U3419 (N_3419,N_3138,N_3150);
xnor U3420 (N_3420,N_3151,N_3294);
nand U3421 (N_3421,N_3214,N_3006);
and U3422 (N_3422,N_3037,N_3027);
nor U3423 (N_3423,N_3010,N_3146);
nor U3424 (N_3424,N_3039,N_3204);
or U3425 (N_3425,N_3145,N_3168);
or U3426 (N_3426,N_3212,N_3223);
nand U3427 (N_3427,N_3045,N_3083);
or U3428 (N_3428,N_3292,N_3260);
and U3429 (N_3429,N_3272,N_3038);
nor U3430 (N_3430,N_3095,N_3116);
nand U3431 (N_3431,N_3031,N_3264);
or U3432 (N_3432,N_3105,N_3215);
nand U3433 (N_3433,N_3071,N_3075);
nand U3434 (N_3434,N_3225,N_3217);
nor U3435 (N_3435,N_3153,N_3195);
xnor U3436 (N_3436,N_3218,N_3275);
or U3437 (N_3437,N_3137,N_3229);
or U3438 (N_3438,N_3016,N_3274);
nor U3439 (N_3439,N_3254,N_3020);
nand U3440 (N_3440,N_3133,N_3203);
or U3441 (N_3441,N_3026,N_3220);
xnor U3442 (N_3442,N_3129,N_3013);
xor U3443 (N_3443,N_3271,N_3259);
or U3444 (N_3444,N_3180,N_3107);
or U3445 (N_3445,N_3084,N_3207);
and U3446 (N_3446,N_3121,N_3159);
nand U3447 (N_3447,N_3147,N_3270);
nand U3448 (N_3448,N_3290,N_3131);
nand U3449 (N_3449,N_3293,N_3143);
and U3450 (N_3450,N_3197,N_3105);
nor U3451 (N_3451,N_3198,N_3055);
or U3452 (N_3452,N_3086,N_3156);
or U3453 (N_3453,N_3032,N_3074);
and U3454 (N_3454,N_3290,N_3019);
nor U3455 (N_3455,N_3237,N_3111);
xnor U3456 (N_3456,N_3017,N_3077);
nor U3457 (N_3457,N_3128,N_3151);
nor U3458 (N_3458,N_3188,N_3225);
or U3459 (N_3459,N_3206,N_3199);
xnor U3460 (N_3460,N_3072,N_3281);
xor U3461 (N_3461,N_3172,N_3155);
and U3462 (N_3462,N_3040,N_3144);
and U3463 (N_3463,N_3183,N_3275);
nand U3464 (N_3464,N_3152,N_3006);
nor U3465 (N_3465,N_3136,N_3046);
or U3466 (N_3466,N_3008,N_3225);
xor U3467 (N_3467,N_3281,N_3060);
and U3468 (N_3468,N_3105,N_3036);
or U3469 (N_3469,N_3066,N_3071);
nand U3470 (N_3470,N_3241,N_3171);
nand U3471 (N_3471,N_3276,N_3087);
nor U3472 (N_3472,N_3252,N_3064);
xnor U3473 (N_3473,N_3227,N_3112);
nor U3474 (N_3474,N_3206,N_3147);
and U3475 (N_3475,N_3203,N_3135);
and U3476 (N_3476,N_3004,N_3023);
nor U3477 (N_3477,N_3221,N_3129);
xnor U3478 (N_3478,N_3248,N_3038);
nand U3479 (N_3479,N_3048,N_3169);
nand U3480 (N_3480,N_3156,N_3137);
nor U3481 (N_3481,N_3150,N_3075);
xor U3482 (N_3482,N_3037,N_3028);
xnor U3483 (N_3483,N_3171,N_3214);
or U3484 (N_3484,N_3202,N_3071);
xnor U3485 (N_3485,N_3274,N_3108);
and U3486 (N_3486,N_3015,N_3163);
nor U3487 (N_3487,N_3089,N_3002);
or U3488 (N_3488,N_3276,N_3095);
nor U3489 (N_3489,N_3131,N_3293);
xor U3490 (N_3490,N_3194,N_3249);
and U3491 (N_3491,N_3000,N_3268);
nand U3492 (N_3492,N_3028,N_3001);
nand U3493 (N_3493,N_3104,N_3288);
nand U3494 (N_3494,N_3132,N_3248);
nand U3495 (N_3495,N_3217,N_3188);
and U3496 (N_3496,N_3150,N_3011);
xor U3497 (N_3497,N_3100,N_3214);
nor U3498 (N_3498,N_3143,N_3248);
nor U3499 (N_3499,N_3191,N_3265);
and U3500 (N_3500,N_3172,N_3024);
or U3501 (N_3501,N_3242,N_3013);
nand U3502 (N_3502,N_3010,N_3212);
nor U3503 (N_3503,N_3071,N_3088);
nor U3504 (N_3504,N_3245,N_3267);
nor U3505 (N_3505,N_3223,N_3195);
nor U3506 (N_3506,N_3286,N_3077);
and U3507 (N_3507,N_3150,N_3096);
nor U3508 (N_3508,N_3039,N_3173);
nand U3509 (N_3509,N_3207,N_3166);
nand U3510 (N_3510,N_3284,N_3104);
nand U3511 (N_3511,N_3166,N_3236);
nand U3512 (N_3512,N_3227,N_3192);
xnor U3513 (N_3513,N_3054,N_3013);
nor U3514 (N_3514,N_3008,N_3246);
and U3515 (N_3515,N_3220,N_3017);
nor U3516 (N_3516,N_3223,N_3090);
nand U3517 (N_3517,N_3190,N_3158);
nand U3518 (N_3518,N_3050,N_3223);
and U3519 (N_3519,N_3187,N_3267);
nand U3520 (N_3520,N_3091,N_3220);
xor U3521 (N_3521,N_3054,N_3213);
nor U3522 (N_3522,N_3246,N_3147);
nor U3523 (N_3523,N_3022,N_3200);
xor U3524 (N_3524,N_3138,N_3297);
nor U3525 (N_3525,N_3195,N_3094);
and U3526 (N_3526,N_3088,N_3083);
or U3527 (N_3527,N_3263,N_3231);
nand U3528 (N_3528,N_3186,N_3182);
nand U3529 (N_3529,N_3020,N_3246);
or U3530 (N_3530,N_3225,N_3048);
nand U3531 (N_3531,N_3277,N_3059);
nor U3532 (N_3532,N_3040,N_3003);
or U3533 (N_3533,N_3029,N_3272);
nand U3534 (N_3534,N_3291,N_3263);
nor U3535 (N_3535,N_3080,N_3201);
nand U3536 (N_3536,N_3108,N_3293);
and U3537 (N_3537,N_3074,N_3153);
xnor U3538 (N_3538,N_3229,N_3258);
nor U3539 (N_3539,N_3061,N_3294);
or U3540 (N_3540,N_3119,N_3275);
and U3541 (N_3541,N_3247,N_3015);
or U3542 (N_3542,N_3090,N_3128);
and U3543 (N_3543,N_3207,N_3295);
or U3544 (N_3544,N_3256,N_3247);
or U3545 (N_3545,N_3169,N_3049);
nand U3546 (N_3546,N_3072,N_3133);
and U3547 (N_3547,N_3129,N_3089);
xnor U3548 (N_3548,N_3245,N_3282);
nand U3549 (N_3549,N_3063,N_3147);
nand U3550 (N_3550,N_3274,N_3121);
xnor U3551 (N_3551,N_3147,N_3009);
nand U3552 (N_3552,N_3152,N_3175);
and U3553 (N_3553,N_3179,N_3195);
or U3554 (N_3554,N_3204,N_3231);
and U3555 (N_3555,N_3151,N_3115);
and U3556 (N_3556,N_3290,N_3003);
xnor U3557 (N_3557,N_3019,N_3152);
or U3558 (N_3558,N_3081,N_3060);
and U3559 (N_3559,N_3223,N_3152);
or U3560 (N_3560,N_3185,N_3154);
or U3561 (N_3561,N_3202,N_3146);
xnor U3562 (N_3562,N_3263,N_3003);
nand U3563 (N_3563,N_3022,N_3184);
nand U3564 (N_3564,N_3199,N_3095);
and U3565 (N_3565,N_3127,N_3220);
or U3566 (N_3566,N_3242,N_3243);
and U3567 (N_3567,N_3193,N_3287);
nand U3568 (N_3568,N_3066,N_3184);
nand U3569 (N_3569,N_3177,N_3015);
nor U3570 (N_3570,N_3280,N_3294);
and U3571 (N_3571,N_3037,N_3048);
nand U3572 (N_3572,N_3014,N_3019);
nor U3573 (N_3573,N_3068,N_3110);
and U3574 (N_3574,N_3267,N_3080);
nand U3575 (N_3575,N_3266,N_3252);
xor U3576 (N_3576,N_3192,N_3122);
or U3577 (N_3577,N_3226,N_3050);
nor U3578 (N_3578,N_3061,N_3280);
and U3579 (N_3579,N_3275,N_3179);
or U3580 (N_3580,N_3194,N_3055);
nand U3581 (N_3581,N_3213,N_3267);
nand U3582 (N_3582,N_3182,N_3180);
or U3583 (N_3583,N_3233,N_3227);
xnor U3584 (N_3584,N_3111,N_3110);
nor U3585 (N_3585,N_3179,N_3076);
or U3586 (N_3586,N_3217,N_3219);
xnor U3587 (N_3587,N_3090,N_3166);
nand U3588 (N_3588,N_3102,N_3298);
and U3589 (N_3589,N_3250,N_3281);
nor U3590 (N_3590,N_3127,N_3115);
and U3591 (N_3591,N_3045,N_3115);
nor U3592 (N_3592,N_3050,N_3218);
xor U3593 (N_3593,N_3131,N_3126);
or U3594 (N_3594,N_3257,N_3023);
nand U3595 (N_3595,N_3217,N_3012);
nor U3596 (N_3596,N_3030,N_3235);
xor U3597 (N_3597,N_3090,N_3229);
nor U3598 (N_3598,N_3133,N_3181);
and U3599 (N_3599,N_3205,N_3237);
or U3600 (N_3600,N_3323,N_3310);
or U3601 (N_3601,N_3529,N_3425);
xor U3602 (N_3602,N_3391,N_3538);
xor U3603 (N_3603,N_3513,N_3500);
and U3604 (N_3604,N_3351,N_3535);
xor U3605 (N_3605,N_3522,N_3347);
or U3606 (N_3606,N_3461,N_3301);
xor U3607 (N_3607,N_3587,N_3599);
and U3608 (N_3608,N_3597,N_3525);
or U3609 (N_3609,N_3305,N_3490);
xor U3610 (N_3610,N_3455,N_3492);
or U3611 (N_3611,N_3449,N_3337);
xor U3612 (N_3612,N_3592,N_3434);
or U3613 (N_3613,N_3575,N_3381);
and U3614 (N_3614,N_3586,N_3325);
or U3615 (N_3615,N_3510,N_3591);
and U3616 (N_3616,N_3559,N_3590);
nand U3617 (N_3617,N_3536,N_3481);
and U3618 (N_3618,N_3317,N_3565);
nor U3619 (N_3619,N_3556,N_3541);
nand U3620 (N_3620,N_3560,N_3393);
and U3621 (N_3621,N_3331,N_3533);
or U3622 (N_3622,N_3466,N_3563);
or U3623 (N_3623,N_3454,N_3552);
nand U3624 (N_3624,N_3468,N_3499);
xor U3625 (N_3625,N_3319,N_3375);
xor U3626 (N_3626,N_3444,N_3428);
and U3627 (N_3627,N_3568,N_3507);
or U3628 (N_3628,N_3504,N_3459);
nand U3629 (N_3629,N_3399,N_3390);
or U3630 (N_3630,N_3540,N_3387);
nand U3631 (N_3631,N_3572,N_3350);
or U3632 (N_3632,N_3363,N_3379);
or U3633 (N_3633,N_3372,N_3557);
and U3634 (N_3634,N_3440,N_3416);
nand U3635 (N_3635,N_3402,N_3366);
nor U3636 (N_3636,N_3333,N_3546);
xnor U3637 (N_3637,N_3594,N_3340);
and U3638 (N_3638,N_3589,N_3571);
nand U3639 (N_3639,N_3397,N_3324);
or U3640 (N_3640,N_3561,N_3421);
xnor U3641 (N_3641,N_3514,N_3473);
nor U3642 (N_3642,N_3370,N_3503);
and U3643 (N_3643,N_3361,N_3443);
nand U3644 (N_3644,N_3482,N_3479);
or U3645 (N_3645,N_3422,N_3532);
nand U3646 (N_3646,N_3498,N_3329);
or U3647 (N_3647,N_3530,N_3446);
xor U3648 (N_3648,N_3314,N_3388);
and U3649 (N_3649,N_3554,N_3356);
nand U3650 (N_3650,N_3573,N_3398);
nand U3651 (N_3651,N_3445,N_3489);
or U3652 (N_3652,N_3374,N_3593);
xor U3653 (N_3653,N_3389,N_3496);
or U3654 (N_3654,N_3400,N_3584);
or U3655 (N_3655,N_3544,N_3477);
or U3656 (N_3656,N_3417,N_3537);
nand U3657 (N_3657,N_3569,N_3352);
and U3658 (N_3658,N_3467,N_3553);
or U3659 (N_3659,N_3579,N_3437);
nand U3660 (N_3660,N_3419,N_3339);
nand U3661 (N_3661,N_3558,N_3345);
or U3662 (N_3662,N_3453,N_3436);
xor U3663 (N_3663,N_3516,N_3312);
nor U3664 (N_3664,N_3472,N_3377);
nor U3665 (N_3665,N_3539,N_3346);
nand U3666 (N_3666,N_3395,N_3386);
nor U3667 (N_3667,N_3450,N_3457);
and U3668 (N_3668,N_3509,N_3595);
xnor U3669 (N_3669,N_3458,N_3407);
xor U3670 (N_3670,N_3564,N_3439);
xor U3671 (N_3671,N_3543,N_3475);
or U3672 (N_3672,N_3414,N_3574);
and U3673 (N_3673,N_3410,N_3527);
nand U3674 (N_3674,N_3369,N_3313);
nor U3675 (N_3675,N_3442,N_3567);
xor U3676 (N_3676,N_3409,N_3338);
nand U3677 (N_3677,N_3460,N_3365);
or U3678 (N_3678,N_3511,N_3570);
and U3679 (N_3679,N_3478,N_3315);
nor U3680 (N_3680,N_3451,N_3506);
nand U3681 (N_3681,N_3578,N_3348);
xor U3682 (N_3682,N_3581,N_3431);
nor U3683 (N_3683,N_3429,N_3380);
nand U3684 (N_3684,N_3502,N_3524);
nor U3685 (N_3685,N_3336,N_3357);
or U3686 (N_3686,N_3394,N_3342);
or U3687 (N_3687,N_3588,N_3542);
and U3688 (N_3688,N_3367,N_3550);
xnor U3689 (N_3689,N_3327,N_3435);
or U3690 (N_3690,N_3353,N_3330);
or U3691 (N_3691,N_3476,N_3344);
nor U3692 (N_3692,N_3562,N_3358);
or U3693 (N_3693,N_3545,N_3306);
nor U3694 (N_3694,N_3470,N_3354);
nand U3695 (N_3695,N_3335,N_3448);
and U3696 (N_3696,N_3474,N_3549);
nand U3697 (N_3697,N_3528,N_3308);
nand U3698 (N_3698,N_3401,N_3495);
xnor U3699 (N_3699,N_3364,N_3403);
nor U3700 (N_3700,N_3368,N_3480);
and U3701 (N_3701,N_3512,N_3566);
nand U3702 (N_3702,N_3383,N_3580);
xor U3703 (N_3703,N_3547,N_3508);
or U3704 (N_3704,N_3487,N_3378);
nor U3705 (N_3705,N_3463,N_3302);
nor U3706 (N_3706,N_3328,N_3355);
or U3707 (N_3707,N_3430,N_3334);
and U3708 (N_3708,N_3362,N_3307);
nand U3709 (N_3709,N_3465,N_3382);
xor U3710 (N_3710,N_3485,N_3464);
or U3711 (N_3711,N_3418,N_3491);
nor U3712 (N_3712,N_3520,N_3517);
xor U3713 (N_3713,N_3384,N_3322);
nand U3714 (N_3714,N_3548,N_3577);
or U3715 (N_3715,N_3483,N_3304);
and U3716 (N_3716,N_3427,N_3341);
and U3717 (N_3717,N_3598,N_3462);
and U3718 (N_3718,N_3413,N_3484);
and U3719 (N_3719,N_3396,N_3371);
and U3720 (N_3720,N_3526,N_3488);
and U3721 (N_3721,N_3300,N_3497);
and U3722 (N_3722,N_3349,N_3424);
and U3723 (N_3723,N_3471,N_3452);
xnor U3724 (N_3724,N_3555,N_3332);
nor U3725 (N_3725,N_3469,N_3385);
nor U3726 (N_3726,N_3456,N_3518);
and U3727 (N_3727,N_3534,N_3309);
nand U3728 (N_3728,N_3486,N_3505);
and U3729 (N_3729,N_3432,N_3423);
and U3730 (N_3730,N_3596,N_3438);
xor U3731 (N_3731,N_3320,N_3415);
nand U3732 (N_3732,N_3420,N_3585);
or U3733 (N_3733,N_3426,N_3316);
nor U3734 (N_3734,N_3493,N_3447);
xnor U3735 (N_3735,N_3501,N_3343);
xnor U3736 (N_3736,N_3318,N_3411);
or U3737 (N_3737,N_3412,N_3441);
xnor U3738 (N_3738,N_3373,N_3408);
nand U3739 (N_3739,N_3359,N_3376);
nand U3740 (N_3740,N_3582,N_3521);
xnor U3741 (N_3741,N_3303,N_3523);
nand U3742 (N_3742,N_3551,N_3531);
nand U3743 (N_3743,N_3404,N_3406);
nand U3744 (N_3744,N_3392,N_3583);
and U3745 (N_3745,N_3360,N_3494);
nand U3746 (N_3746,N_3405,N_3311);
nor U3747 (N_3747,N_3515,N_3519);
nor U3748 (N_3748,N_3326,N_3576);
nor U3749 (N_3749,N_3433,N_3321);
xor U3750 (N_3750,N_3584,N_3345);
or U3751 (N_3751,N_3503,N_3516);
and U3752 (N_3752,N_3345,N_3314);
and U3753 (N_3753,N_3411,N_3324);
or U3754 (N_3754,N_3592,N_3430);
nor U3755 (N_3755,N_3556,N_3534);
nor U3756 (N_3756,N_3331,N_3314);
nand U3757 (N_3757,N_3457,N_3339);
xnor U3758 (N_3758,N_3458,N_3493);
nor U3759 (N_3759,N_3570,N_3479);
or U3760 (N_3760,N_3423,N_3388);
xor U3761 (N_3761,N_3545,N_3522);
xor U3762 (N_3762,N_3496,N_3327);
nand U3763 (N_3763,N_3555,N_3392);
nor U3764 (N_3764,N_3385,N_3529);
xor U3765 (N_3765,N_3430,N_3444);
nand U3766 (N_3766,N_3326,N_3507);
nand U3767 (N_3767,N_3458,N_3422);
nand U3768 (N_3768,N_3370,N_3563);
xor U3769 (N_3769,N_3329,N_3578);
or U3770 (N_3770,N_3358,N_3382);
nand U3771 (N_3771,N_3436,N_3501);
xnor U3772 (N_3772,N_3454,N_3514);
and U3773 (N_3773,N_3533,N_3535);
nor U3774 (N_3774,N_3380,N_3529);
xor U3775 (N_3775,N_3527,N_3491);
and U3776 (N_3776,N_3553,N_3515);
nor U3777 (N_3777,N_3495,N_3376);
and U3778 (N_3778,N_3577,N_3440);
or U3779 (N_3779,N_3480,N_3471);
xnor U3780 (N_3780,N_3354,N_3467);
and U3781 (N_3781,N_3473,N_3572);
and U3782 (N_3782,N_3493,N_3466);
xnor U3783 (N_3783,N_3327,N_3480);
and U3784 (N_3784,N_3476,N_3433);
or U3785 (N_3785,N_3409,N_3493);
or U3786 (N_3786,N_3488,N_3405);
or U3787 (N_3787,N_3385,N_3520);
and U3788 (N_3788,N_3468,N_3534);
nand U3789 (N_3789,N_3511,N_3521);
and U3790 (N_3790,N_3569,N_3475);
nand U3791 (N_3791,N_3383,N_3407);
xnor U3792 (N_3792,N_3526,N_3318);
nor U3793 (N_3793,N_3551,N_3321);
nor U3794 (N_3794,N_3471,N_3361);
nand U3795 (N_3795,N_3347,N_3465);
and U3796 (N_3796,N_3512,N_3481);
nand U3797 (N_3797,N_3377,N_3318);
xor U3798 (N_3798,N_3381,N_3587);
or U3799 (N_3799,N_3370,N_3596);
nand U3800 (N_3800,N_3566,N_3534);
and U3801 (N_3801,N_3368,N_3329);
nand U3802 (N_3802,N_3542,N_3517);
nand U3803 (N_3803,N_3429,N_3500);
or U3804 (N_3804,N_3583,N_3321);
xor U3805 (N_3805,N_3598,N_3549);
and U3806 (N_3806,N_3568,N_3377);
xor U3807 (N_3807,N_3415,N_3414);
and U3808 (N_3808,N_3463,N_3439);
or U3809 (N_3809,N_3357,N_3472);
or U3810 (N_3810,N_3499,N_3398);
nand U3811 (N_3811,N_3548,N_3441);
nand U3812 (N_3812,N_3505,N_3348);
nor U3813 (N_3813,N_3457,N_3546);
or U3814 (N_3814,N_3486,N_3509);
nor U3815 (N_3815,N_3538,N_3465);
nand U3816 (N_3816,N_3539,N_3492);
nand U3817 (N_3817,N_3329,N_3395);
or U3818 (N_3818,N_3353,N_3359);
and U3819 (N_3819,N_3554,N_3493);
and U3820 (N_3820,N_3329,N_3373);
nor U3821 (N_3821,N_3564,N_3453);
and U3822 (N_3822,N_3421,N_3480);
xor U3823 (N_3823,N_3383,N_3314);
and U3824 (N_3824,N_3510,N_3411);
xor U3825 (N_3825,N_3397,N_3536);
nor U3826 (N_3826,N_3467,N_3430);
nand U3827 (N_3827,N_3395,N_3571);
nand U3828 (N_3828,N_3434,N_3536);
xnor U3829 (N_3829,N_3489,N_3407);
nor U3830 (N_3830,N_3534,N_3463);
xnor U3831 (N_3831,N_3517,N_3359);
and U3832 (N_3832,N_3377,N_3309);
or U3833 (N_3833,N_3350,N_3481);
and U3834 (N_3834,N_3448,N_3490);
or U3835 (N_3835,N_3449,N_3522);
or U3836 (N_3836,N_3353,N_3515);
xnor U3837 (N_3837,N_3480,N_3469);
and U3838 (N_3838,N_3468,N_3445);
nand U3839 (N_3839,N_3347,N_3313);
and U3840 (N_3840,N_3336,N_3328);
nor U3841 (N_3841,N_3365,N_3359);
nor U3842 (N_3842,N_3527,N_3393);
nand U3843 (N_3843,N_3567,N_3517);
or U3844 (N_3844,N_3587,N_3434);
nand U3845 (N_3845,N_3354,N_3403);
nand U3846 (N_3846,N_3491,N_3443);
and U3847 (N_3847,N_3341,N_3368);
nand U3848 (N_3848,N_3339,N_3475);
nand U3849 (N_3849,N_3375,N_3500);
xor U3850 (N_3850,N_3511,N_3546);
xnor U3851 (N_3851,N_3367,N_3472);
or U3852 (N_3852,N_3374,N_3427);
nand U3853 (N_3853,N_3531,N_3586);
nor U3854 (N_3854,N_3305,N_3377);
or U3855 (N_3855,N_3544,N_3377);
nor U3856 (N_3856,N_3508,N_3561);
nor U3857 (N_3857,N_3494,N_3340);
nor U3858 (N_3858,N_3538,N_3590);
or U3859 (N_3859,N_3460,N_3459);
and U3860 (N_3860,N_3509,N_3482);
xnor U3861 (N_3861,N_3401,N_3456);
or U3862 (N_3862,N_3336,N_3564);
xnor U3863 (N_3863,N_3482,N_3440);
xnor U3864 (N_3864,N_3456,N_3533);
xor U3865 (N_3865,N_3356,N_3405);
nand U3866 (N_3866,N_3363,N_3431);
nand U3867 (N_3867,N_3546,N_3527);
nor U3868 (N_3868,N_3588,N_3476);
nor U3869 (N_3869,N_3589,N_3544);
xor U3870 (N_3870,N_3536,N_3516);
xnor U3871 (N_3871,N_3459,N_3395);
or U3872 (N_3872,N_3523,N_3411);
xor U3873 (N_3873,N_3433,N_3322);
xnor U3874 (N_3874,N_3384,N_3477);
nand U3875 (N_3875,N_3353,N_3564);
nand U3876 (N_3876,N_3534,N_3316);
or U3877 (N_3877,N_3446,N_3481);
nand U3878 (N_3878,N_3428,N_3356);
xnor U3879 (N_3879,N_3364,N_3394);
nand U3880 (N_3880,N_3350,N_3305);
nand U3881 (N_3881,N_3447,N_3546);
xnor U3882 (N_3882,N_3430,N_3362);
xnor U3883 (N_3883,N_3486,N_3469);
or U3884 (N_3884,N_3344,N_3546);
and U3885 (N_3885,N_3484,N_3483);
nand U3886 (N_3886,N_3441,N_3545);
or U3887 (N_3887,N_3372,N_3334);
nor U3888 (N_3888,N_3363,N_3464);
and U3889 (N_3889,N_3545,N_3406);
and U3890 (N_3890,N_3381,N_3551);
nor U3891 (N_3891,N_3587,N_3516);
nor U3892 (N_3892,N_3458,N_3447);
xnor U3893 (N_3893,N_3565,N_3483);
nor U3894 (N_3894,N_3420,N_3483);
or U3895 (N_3895,N_3539,N_3597);
xor U3896 (N_3896,N_3447,N_3545);
nor U3897 (N_3897,N_3470,N_3554);
nor U3898 (N_3898,N_3418,N_3388);
and U3899 (N_3899,N_3353,N_3369);
nand U3900 (N_3900,N_3718,N_3762);
nand U3901 (N_3901,N_3677,N_3625);
or U3902 (N_3902,N_3651,N_3787);
or U3903 (N_3903,N_3786,N_3867);
or U3904 (N_3904,N_3745,N_3803);
nand U3905 (N_3905,N_3874,N_3802);
nand U3906 (N_3906,N_3796,N_3737);
nor U3907 (N_3907,N_3878,N_3889);
and U3908 (N_3908,N_3828,N_3845);
xor U3909 (N_3909,N_3750,N_3612);
nand U3910 (N_3910,N_3731,N_3735);
nor U3911 (N_3911,N_3881,N_3720);
xor U3912 (N_3912,N_3780,N_3690);
xor U3913 (N_3913,N_3623,N_3713);
and U3914 (N_3914,N_3806,N_3835);
xnor U3915 (N_3915,N_3888,N_3733);
xnor U3916 (N_3916,N_3817,N_3675);
and U3917 (N_3917,N_3716,N_3781);
nand U3918 (N_3918,N_3822,N_3634);
nor U3919 (N_3919,N_3691,N_3616);
nand U3920 (N_3920,N_3665,N_3614);
and U3921 (N_3921,N_3622,N_3722);
or U3922 (N_3922,N_3818,N_3648);
nand U3923 (N_3923,N_3746,N_3724);
and U3924 (N_3924,N_3788,N_3608);
xor U3925 (N_3925,N_3683,N_3668);
or U3926 (N_3926,N_3671,N_3710);
xnor U3927 (N_3927,N_3784,N_3891);
xor U3928 (N_3928,N_3744,N_3755);
or U3929 (N_3929,N_3662,N_3840);
or U3930 (N_3930,N_3858,N_3851);
or U3931 (N_3931,N_3830,N_3853);
and U3932 (N_3932,N_3761,N_3846);
nor U3933 (N_3933,N_3844,N_3615);
xnor U3934 (N_3934,N_3887,N_3613);
nand U3935 (N_3935,N_3639,N_3813);
xor U3936 (N_3936,N_3816,N_3884);
or U3937 (N_3937,N_3848,N_3606);
nand U3938 (N_3938,N_3740,N_3669);
nand U3939 (N_3939,N_3605,N_3836);
xor U3940 (N_3940,N_3689,N_3892);
or U3941 (N_3941,N_3667,N_3661);
or U3942 (N_3942,N_3857,N_3795);
nor U3943 (N_3943,N_3783,N_3793);
xor U3944 (N_3944,N_3820,N_3753);
nor U3945 (N_3945,N_3772,N_3704);
xor U3946 (N_3946,N_3672,N_3798);
nor U3947 (N_3947,N_3859,N_3712);
and U3948 (N_3948,N_3785,N_3607);
xnor U3949 (N_3949,N_3684,N_3601);
xnor U3950 (N_3950,N_3760,N_3764);
xnor U3951 (N_3951,N_3626,N_3794);
nor U3952 (N_3952,N_3657,N_3666);
and U3953 (N_3953,N_3637,N_3656);
nand U3954 (N_3954,N_3842,N_3875);
nor U3955 (N_3955,N_3638,N_3885);
xnor U3956 (N_3956,N_3777,N_3664);
xnor U3957 (N_3957,N_3653,N_3826);
xnor U3958 (N_3958,N_3629,N_3654);
xnor U3959 (N_3959,N_3870,N_3834);
and U3960 (N_3960,N_3749,N_3847);
nand U3961 (N_3961,N_3701,N_3670);
or U3962 (N_3962,N_3682,N_3633);
and U3963 (N_3963,N_3739,N_3636);
or U3964 (N_3964,N_3610,N_3824);
nor U3965 (N_3965,N_3688,N_3645);
nand U3966 (N_3966,N_3797,N_3642);
or U3967 (N_3967,N_3838,N_3694);
nand U3968 (N_3968,N_3640,N_3896);
nor U3969 (N_3969,N_3877,N_3717);
nor U3970 (N_3970,N_3759,N_3897);
nand U3971 (N_3971,N_3650,N_3821);
nand U3972 (N_3972,N_3705,N_3685);
nand U3973 (N_3973,N_3829,N_3679);
or U3974 (N_3974,N_3841,N_3680);
and U3975 (N_3975,N_3758,N_3766);
nor U3976 (N_3976,N_3812,N_3603);
xor U3977 (N_3977,N_3831,N_3873);
or U3978 (N_3978,N_3769,N_3620);
and U3979 (N_3979,N_3678,N_3736);
and U3980 (N_3980,N_3658,N_3602);
nand U3981 (N_3981,N_3839,N_3808);
nor U3982 (N_3982,N_3600,N_3631);
nand U3983 (N_3983,N_3827,N_3630);
nor U3984 (N_3984,N_3673,N_3728);
nand U3985 (N_3985,N_3810,N_3837);
or U3986 (N_3986,N_3635,N_3864);
xor U3987 (N_3987,N_3632,N_3660);
xor U3988 (N_3988,N_3641,N_3687);
and U3989 (N_3989,N_3833,N_3729);
nand U3990 (N_3990,N_3702,N_3895);
and U3991 (N_3991,N_3799,N_3748);
and U3992 (N_3992,N_3770,N_3757);
or U3993 (N_3993,N_3789,N_3681);
nor U3994 (N_3994,N_3696,N_3815);
nor U3995 (N_3995,N_3611,N_3819);
nor U3996 (N_3996,N_3862,N_3856);
and U3997 (N_3997,N_3801,N_3843);
or U3998 (N_3998,N_3619,N_3778);
nor U3999 (N_3999,N_3709,N_3768);
xor U4000 (N_4000,N_3741,N_3898);
and U4001 (N_4001,N_3861,N_3699);
nor U4002 (N_4002,N_3686,N_3860);
and U4003 (N_4003,N_3866,N_3617);
or U4004 (N_4004,N_3854,N_3697);
and U4005 (N_4005,N_3730,N_3621);
nor U4006 (N_4006,N_3751,N_3775);
nand U4007 (N_4007,N_3782,N_3644);
nand U4008 (N_4008,N_3707,N_3773);
xnor U4009 (N_4009,N_3894,N_3804);
or U4010 (N_4010,N_3871,N_3872);
xnor U4011 (N_4011,N_3890,N_3734);
and U4012 (N_4012,N_3809,N_3883);
nand U4013 (N_4013,N_3850,N_3792);
nand U4014 (N_4014,N_3832,N_3695);
and U4015 (N_4015,N_3880,N_3719);
nor U4016 (N_4016,N_3643,N_3742);
and U4017 (N_4017,N_3869,N_3727);
nand U4018 (N_4018,N_3714,N_3693);
nor U4019 (N_4019,N_3790,N_3868);
nand U4020 (N_4020,N_3700,N_3765);
and U4021 (N_4021,N_3655,N_3852);
or U4022 (N_4022,N_3715,N_3706);
xor U4023 (N_4023,N_3646,N_3723);
nor U4024 (N_4024,N_3774,N_3747);
or U4025 (N_4025,N_3879,N_3767);
or U4026 (N_4026,N_3849,N_3618);
xor U4027 (N_4027,N_3676,N_3604);
and U4028 (N_4028,N_3823,N_3624);
xor U4029 (N_4029,N_3863,N_3721);
xnor U4030 (N_4030,N_3752,N_3791);
and U4031 (N_4031,N_3814,N_3865);
nor U4032 (N_4032,N_3652,N_3698);
nand U4033 (N_4033,N_3855,N_3609);
xnor U4034 (N_4034,N_3732,N_3763);
xor U4035 (N_4035,N_3692,N_3627);
or U4036 (N_4036,N_3779,N_3756);
and U4037 (N_4037,N_3886,N_3805);
nor U4038 (N_4038,N_3899,N_3659);
and U4039 (N_4039,N_3726,N_3725);
or U4040 (N_4040,N_3649,N_3754);
nor U4041 (N_4041,N_3893,N_3771);
xnor U4042 (N_4042,N_3674,N_3876);
nand U4043 (N_4043,N_3743,N_3663);
or U4044 (N_4044,N_3807,N_3825);
or U4045 (N_4045,N_3776,N_3628);
or U4046 (N_4046,N_3811,N_3708);
and U4047 (N_4047,N_3647,N_3711);
and U4048 (N_4048,N_3703,N_3800);
nor U4049 (N_4049,N_3738,N_3882);
nor U4050 (N_4050,N_3633,N_3893);
nor U4051 (N_4051,N_3731,N_3709);
or U4052 (N_4052,N_3775,N_3894);
nor U4053 (N_4053,N_3607,N_3637);
nand U4054 (N_4054,N_3787,N_3652);
nor U4055 (N_4055,N_3731,N_3897);
nor U4056 (N_4056,N_3797,N_3863);
or U4057 (N_4057,N_3670,N_3671);
and U4058 (N_4058,N_3834,N_3767);
nor U4059 (N_4059,N_3860,N_3763);
or U4060 (N_4060,N_3684,N_3686);
and U4061 (N_4061,N_3852,N_3636);
nand U4062 (N_4062,N_3765,N_3627);
or U4063 (N_4063,N_3627,N_3760);
or U4064 (N_4064,N_3893,N_3691);
nor U4065 (N_4065,N_3613,N_3700);
nor U4066 (N_4066,N_3821,N_3793);
nand U4067 (N_4067,N_3643,N_3826);
nand U4068 (N_4068,N_3620,N_3810);
xnor U4069 (N_4069,N_3617,N_3668);
nor U4070 (N_4070,N_3822,N_3759);
nor U4071 (N_4071,N_3772,N_3738);
nand U4072 (N_4072,N_3770,N_3740);
nor U4073 (N_4073,N_3704,N_3702);
nor U4074 (N_4074,N_3868,N_3883);
and U4075 (N_4075,N_3866,N_3792);
xor U4076 (N_4076,N_3752,N_3765);
nor U4077 (N_4077,N_3604,N_3714);
nor U4078 (N_4078,N_3649,N_3732);
nand U4079 (N_4079,N_3786,N_3750);
or U4080 (N_4080,N_3887,N_3642);
nor U4081 (N_4081,N_3636,N_3897);
xor U4082 (N_4082,N_3735,N_3823);
nor U4083 (N_4083,N_3823,N_3730);
and U4084 (N_4084,N_3853,N_3778);
nor U4085 (N_4085,N_3825,N_3683);
xnor U4086 (N_4086,N_3769,N_3845);
xnor U4087 (N_4087,N_3794,N_3779);
or U4088 (N_4088,N_3795,N_3665);
or U4089 (N_4089,N_3786,N_3601);
and U4090 (N_4090,N_3612,N_3614);
nor U4091 (N_4091,N_3637,N_3892);
and U4092 (N_4092,N_3687,N_3703);
or U4093 (N_4093,N_3855,N_3851);
and U4094 (N_4094,N_3614,N_3723);
nand U4095 (N_4095,N_3677,N_3733);
xor U4096 (N_4096,N_3697,N_3868);
nor U4097 (N_4097,N_3815,N_3716);
or U4098 (N_4098,N_3888,N_3860);
and U4099 (N_4099,N_3843,N_3874);
or U4100 (N_4100,N_3884,N_3638);
or U4101 (N_4101,N_3676,N_3645);
or U4102 (N_4102,N_3832,N_3603);
or U4103 (N_4103,N_3890,N_3761);
nand U4104 (N_4104,N_3859,N_3766);
nand U4105 (N_4105,N_3742,N_3744);
nand U4106 (N_4106,N_3683,N_3727);
nor U4107 (N_4107,N_3798,N_3680);
xor U4108 (N_4108,N_3881,N_3618);
or U4109 (N_4109,N_3859,N_3836);
and U4110 (N_4110,N_3686,N_3728);
nor U4111 (N_4111,N_3686,N_3861);
xnor U4112 (N_4112,N_3682,N_3676);
or U4113 (N_4113,N_3847,N_3848);
or U4114 (N_4114,N_3643,N_3664);
nand U4115 (N_4115,N_3654,N_3665);
nand U4116 (N_4116,N_3656,N_3742);
nand U4117 (N_4117,N_3601,N_3788);
or U4118 (N_4118,N_3777,N_3660);
and U4119 (N_4119,N_3674,N_3646);
xnor U4120 (N_4120,N_3755,N_3801);
xnor U4121 (N_4121,N_3795,N_3704);
xor U4122 (N_4122,N_3751,N_3815);
nand U4123 (N_4123,N_3602,N_3616);
nor U4124 (N_4124,N_3759,N_3695);
nor U4125 (N_4125,N_3610,N_3646);
and U4126 (N_4126,N_3835,N_3712);
nor U4127 (N_4127,N_3695,N_3692);
nor U4128 (N_4128,N_3766,N_3662);
nor U4129 (N_4129,N_3754,N_3705);
nor U4130 (N_4130,N_3888,N_3671);
or U4131 (N_4131,N_3606,N_3662);
xor U4132 (N_4132,N_3695,N_3617);
or U4133 (N_4133,N_3834,N_3893);
and U4134 (N_4134,N_3628,N_3679);
and U4135 (N_4135,N_3888,N_3730);
xor U4136 (N_4136,N_3604,N_3765);
or U4137 (N_4137,N_3676,N_3784);
xnor U4138 (N_4138,N_3784,N_3680);
or U4139 (N_4139,N_3754,N_3825);
xor U4140 (N_4140,N_3827,N_3808);
xnor U4141 (N_4141,N_3853,N_3684);
nor U4142 (N_4142,N_3809,N_3774);
or U4143 (N_4143,N_3747,N_3777);
xnor U4144 (N_4144,N_3896,N_3843);
and U4145 (N_4145,N_3694,N_3776);
xor U4146 (N_4146,N_3706,N_3615);
and U4147 (N_4147,N_3607,N_3852);
xnor U4148 (N_4148,N_3689,N_3786);
xor U4149 (N_4149,N_3691,N_3839);
nand U4150 (N_4150,N_3767,N_3796);
xnor U4151 (N_4151,N_3687,N_3662);
and U4152 (N_4152,N_3629,N_3678);
and U4153 (N_4153,N_3744,N_3890);
and U4154 (N_4154,N_3895,N_3843);
or U4155 (N_4155,N_3721,N_3738);
or U4156 (N_4156,N_3725,N_3758);
nand U4157 (N_4157,N_3861,N_3874);
nor U4158 (N_4158,N_3886,N_3870);
nor U4159 (N_4159,N_3800,N_3738);
and U4160 (N_4160,N_3778,N_3650);
nand U4161 (N_4161,N_3799,N_3876);
xnor U4162 (N_4162,N_3634,N_3772);
nor U4163 (N_4163,N_3774,N_3780);
or U4164 (N_4164,N_3737,N_3800);
and U4165 (N_4165,N_3745,N_3887);
nand U4166 (N_4166,N_3785,N_3893);
xor U4167 (N_4167,N_3707,N_3887);
nand U4168 (N_4168,N_3649,N_3676);
nand U4169 (N_4169,N_3864,N_3825);
xor U4170 (N_4170,N_3849,N_3642);
nand U4171 (N_4171,N_3729,N_3634);
or U4172 (N_4172,N_3685,N_3720);
or U4173 (N_4173,N_3622,N_3632);
nor U4174 (N_4174,N_3704,N_3898);
xnor U4175 (N_4175,N_3810,N_3862);
or U4176 (N_4176,N_3614,N_3666);
nor U4177 (N_4177,N_3802,N_3865);
and U4178 (N_4178,N_3767,N_3623);
and U4179 (N_4179,N_3889,N_3861);
xor U4180 (N_4180,N_3602,N_3719);
xnor U4181 (N_4181,N_3614,N_3852);
nor U4182 (N_4182,N_3771,N_3637);
nor U4183 (N_4183,N_3898,N_3639);
or U4184 (N_4184,N_3726,N_3636);
nand U4185 (N_4185,N_3642,N_3622);
xor U4186 (N_4186,N_3698,N_3741);
xnor U4187 (N_4187,N_3818,N_3839);
or U4188 (N_4188,N_3885,N_3663);
nor U4189 (N_4189,N_3821,N_3836);
xnor U4190 (N_4190,N_3620,N_3899);
nor U4191 (N_4191,N_3688,N_3722);
xnor U4192 (N_4192,N_3896,N_3624);
nand U4193 (N_4193,N_3745,N_3808);
or U4194 (N_4194,N_3842,N_3713);
xnor U4195 (N_4195,N_3833,N_3605);
nor U4196 (N_4196,N_3730,N_3802);
and U4197 (N_4197,N_3819,N_3820);
nor U4198 (N_4198,N_3638,N_3883);
nor U4199 (N_4199,N_3613,N_3605);
nand U4200 (N_4200,N_3949,N_3959);
and U4201 (N_4201,N_4139,N_4076);
nor U4202 (N_4202,N_4052,N_4071);
xor U4203 (N_4203,N_4006,N_4027);
and U4204 (N_4204,N_3929,N_3928);
nand U4205 (N_4205,N_4144,N_4099);
or U4206 (N_4206,N_3901,N_4054);
or U4207 (N_4207,N_4080,N_3990);
nand U4208 (N_4208,N_4060,N_3907);
nand U4209 (N_4209,N_4170,N_4079);
nor U4210 (N_4210,N_3988,N_4048);
nor U4211 (N_4211,N_3913,N_4164);
or U4212 (N_4212,N_3960,N_3912);
xnor U4213 (N_4213,N_4166,N_3980);
or U4214 (N_4214,N_3934,N_4065);
nand U4215 (N_4215,N_4188,N_4009);
and U4216 (N_4216,N_4125,N_4094);
or U4217 (N_4217,N_4191,N_4105);
nor U4218 (N_4218,N_3968,N_4152);
xor U4219 (N_4219,N_4167,N_4151);
nor U4220 (N_4220,N_4121,N_4040);
nor U4221 (N_4221,N_4103,N_4180);
and U4222 (N_4222,N_3975,N_3918);
and U4223 (N_4223,N_4174,N_3950);
nor U4224 (N_4224,N_4134,N_4148);
xor U4225 (N_4225,N_4022,N_3937);
nand U4226 (N_4226,N_3941,N_4101);
or U4227 (N_4227,N_3974,N_4136);
xnor U4228 (N_4228,N_3940,N_3970);
nor U4229 (N_4229,N_4003,N_4111);
nand U4230 (N_4230,N_4176,N_4190);
xnor U4231 (N_4231,N_4091,N_3945);
or U4232 (N_4232,N_4020,N_4186);
nor U4233 (N_4233,N_4074,N_3948);
xor U4234 (N_4234,N_3911,N_4118);
and U4235 (N_4235,N_4171,N_4175);
nor U4236 (N_4236,N_3909,N_4081);
and U4237 (N_4237,N_4072,N_3919);
nand U4238 (N_4238,N_4024,N_3964);
and U4239 (N_4239,N_3967,N_3930);
xnor U4240 (N_4240,N_4128,N_4078);
xor U4241 (N_4241,N_4117,N_4042);
and U4242 (N_4242,N_3927,N_3916);
nor U4243 (N_4243,N_4077,N_3935);
nand U4244 (N_4244,N_3951,N_4088);
or U4245 (N_4245,N_4033,N_4126);
xnor U4246 (N_4246,N_4001,N_4084);
or U4247 (N_4247,N_4199,N_4122);
xor U4248 (N_4248,N_4127,N_3996);
nor U4249 (N_4249,N_4098,N_4132);
xnor U4250 (N_4250,N_4093,N_4012);
xnor U4251 (N_4251,N_4133,N_3963);
nand U4252 (N_4252,N_3947,N_3903);
nand U4253 (N_4253,N_4029,N_4181);
xnor U4254 (N_4254,N_4082,N_3946);
xor U4255 (N_4255,N_3914,N_4124);
nor U4256 (N_4256,N_4142,N_4067);
nor U4257 (N_4257,N_4141,N_4197);
nand U4258 (N_4258,N_3938,N_4109);
nand U4259 (N_4259,N_4000,N_4187);
nand U4260 (N_4260,N_4092,N_4032);
or U4261 (N_4261,N_4043,N_3915);
xor U4262 (N_4262,N_4157,N_4189);
nor U4263 (N_4263,N_4096,N_3943);
or U4264 (N_4264,N_4041,N_4162);
xor U4265 (N_4265,N_3979,N_4194);
and U4266 (N_4266,N_3992,N_4120);
xor U4267 (N_4267,N_4063,N_3993);
nor U4268 (N_4268,N_4031,N_3976);
nand U4269 (N_4269,N_3983,N_4073);
xor U4270 (N_4270,N_4049,N_4149);
and U4271 (N_4271,N_4070,N_4016);
nand U4272 (N_4272,N_4097,N_4156);
or U4273 (N_4273,N_4123,N_4058);
nand U4274 (N_4274,N_3921,N_3944);
nor U4275 (N_4275,N_4178,N_4193);
and U4276 (N_4276,N_4083,N_3999);
and U4277 (N_4277,N_4037,N_4100);
nor U4278 (N_4278,N_4116,N_3982);
nand U4279 (N_4279,N_4147,N_4046);
nand U4280 (N_4280,N_3920,N_4008);
nor U4281 (N_4281,N_4115,N_4165);
xor U4282 (N_4282,N_3966,N_4026);
nand U4283 (N_4283,N_4168,N_3923);
xnor U4284 (N_4284,N_4062,N_4055);
xnor U4285 (N_4285,N_3962,N_4159);
or U4286 (N_4286,N_4085,N_4137);
xnor U4287 (N_4287,N_4028,N_3936);
nand U4288 (N_4288,N_4007,N_4179);
or U4289 (N_4289,N_3987,N_3926);
nor U4290 (N_4290,N_4021,N_4034);
and U4291 (N_4291,N_4114,N_3986);
nand U4292 (N_4292,N_4195,N_4064);
and U4293 (N_4293,N_3942,N_4131);
xnor U4294 (N_4294,N_4038,N_3917);
nor U4295 (N_4295,N_4086,N_4013);
nor U4296 (N_4296,N_4010,N_4095);
and U4297 (N_4297,N_4112,N_4153);
or U4298 (N_4298,N_4035,N_3953);
nor U4299 (N_4299,N_4160,N_3922);
nand U4300 (N_4300,N_3902,N_4158);
xnor U4301 (N_4301,N_4161,N_3985);
or U4302 (N_4302,N_4196,N_4089);
or U4303 (N_4303,N_4107,N_4075);
or U4304 (N_4304,N_4025,N_3954);
nor U4305 (N_4305,N_4106,N_4011);
nor U4306 (N_4306,N_3904,N_3955);
nor U4307 (N_4307,N_4023,N_4039);
nor U4308 (N_4308,N_4017,N_4154);
nand U4309 (N_4309,N_4155,N_4177);
or U4310 (N_4310,N_4184,N_3910);
nor U4311 (N_4311,N_3924,N_4019);
and U4312 (N_4312,N_3965,N_3977);
xor U4313 (N_4313,N_3939,N_4018);
nor U4314 (N_4314,N_4135,N_4146);
nor U4315 (N_4315,N_3957,N_4004);
nand U4316 (N_4316,N_3932,N_4172);
or U4317 (N_4317,N_4061,N_3933);
and U4318 (N_4318,N_3905,N_3971);
nor U4319 (N_4319,N_4104,N_3906);
or U4320 (N_4320,N_4045,N_4087);
nand U4321 (N_4321,N_3958,N_4108);
or U4322 (N_4322,N_4183,N_3961);
and U4323 (N_4323,N_4014,N_4044);
nand U4324 (N_4324,N_4102,N_3972);
nand U4325 (N_4325,N_4090,N_4015);
nor U4326 (N_4326,N_4002,N_3973);
nor U4327 (N_4327,N_3991,N_3981);
nand U4328 (N_4328,N_3908,N_4138);
nand U4329 (N_4329,N_4185,N_4066);
or U4330 (N_4330,N_4050,N_3978);
xor U4331 (N_4331,N_4047,N_4140);
or U4332 (N_4332,N_3997,N_3998);
nor U4333 (N_4333,N_4150,N_4030);
nand U4334 (N_4334,N_4129,N_4113);
nor U4335 (N_4335,N_4051,N_4192);
nor U4336 (N_4336,N_3952,N_4182);
nor U4337 (N_4337,N_4053,N_4059);
nor U4338 (N_4338,N_4173,N_3969);
nor U4339 (N_4339,N_4068,N_3989);
nor U4340 (N_4340,N_3931,N_4163);
and U4341 (N_4341,N_3995,N_3984);
and U4342 (N_4342,N_4130,N_4198);
nand U4343 (N_4343,N_4169,N_4110);
nand U4344 (N_4344,N_3956,N_4036);
nor U4345 (N_4345,N_4143,N_3994);
and U4346 (N_4346,N_4145,N_3925);
xnor U4347 (N_4347,N_4005,N_3900);
xor U4348 (N_4348,N_4056,N_4057);
or U4349 (N_4349,N_4069,N_4119);
or U4350 (N_4350,N_4141,N_4195);
nor U4351 (N_4351,N_4188,N_4117);
or U4352 (N_4352,N_4165,N_3917);
nand U4353 (N_4353,N_4189,N_4138);
and U4354 (N_4354,N_4030,N_4080);
and U4355 (N_4355,N_4148,N_4120);
or U4356 (N_4356,N_4198,N_4184);
xnor U4357 (N_4357,N_3970,N_4168);
nor U4358 (N_4358,N_4180,N_4008);
nand U4359 (N_4359,N_4001,N_4172);
nand U4360 (N_4360,N_4029,N_4022);
and U4361 (N_4361,N_3942,N_3944);
nor U4362 (N_4362,N_4056,N_3970);
or U4363 (N_4363,N_3953,N_3931);
nor U4364 (N_4364,N_4164,N_3914);
nor U4365 (N_4365,N_4190,N_3909);
or U4366 (N_4366,N_4178,N_4145);
nor U4367 (N_4367,N_4162,N_3929);
xor U4368 (N_4368,N_4079,N_4073);
or U4369 (N_4369,N_3947,N_4002);
nor U4370 (N_4370,N_4038,N_3968);
or U4371 (N_4371,N_4089,N_4029);
and U4372 (N_4372,N_4009,N_4128);
and U4373 (N_4373,N_4087,N_4005);
or U4374 (N_4374,N_4097,N_3966);
nand U4375 (N_4375,N_3992,N_4003);
or U4376 (N_4376,N_3934,N_4035);
nand U4377 (N_4377,N_3954,N_4118);
or U4378 (N_4378,N_4147,N_3958);
nand U4379 (N_4379,N_3934,N_3975);
xnor U4380 (N_4380,N_3976,N_4028);
xnor U4381 (N_4381,N_3971,N_4192);
and U4382 (N_4382,N_4197,N_4049);
xor U4383 (N_4383,N_3947,N_3930);
nand U4384 (N_4384,N_4055,N_4064);
or U4385 (N_4385,N_4041,N_4028);
or U4386 (N_4386,N_3956,N_4050);
xnor U4387 (N_4387,N_4144,N_3932);
xnor U4388 (N_4388,N_3996,N_3926);
nor U4389 (N_4389,N_4023,N_3922);
nand U4390 (N_4390,N_4099,N_4100);
nand U4391 (N_4391,N_4165,N_4024);
xor U4392 (N_4392,N_3982,N_3925);
and U4393 (N_4393,N_4129,N_4122);
nor U4394 (N_4394,N_4107,N_4147);
or U4395 (N_4395,N_3964,N_3987);
and U4396 (N_4396,N_3979,N_4182);
xor U4397 (N_4397,N_4060,N_3982);
nor U4398 (N_4398,N_3975,N_4085);
or U4399 (N_4399,N_4025,N_4010);
and U4400 (N_4400,N_4166,N_4061);
or U4401 (N_4401,N_4142,N_4136);
or U4402 (N_4402,N_4103,N_4072);
xor U4403 (N_4403,N_3967,N_4196);
and U4404 (N_4404,N_4099,N_4154);
nand U4405 (N_4405,N_4052,N_3926);
nand U4406 (N_4406,N_4045,N_4081);
nor U4407 (N_4407,N_4028,N_3916);
nand U4408 (N_4408,N_4073,N_4007);
and U4409 (N_4409,N_3914,N_4088);
nor U4410 (N_4410,N_3945,N_3926);
xor U4411 (N_4411,N_4083,N_3944);
and U4412 (N_4412,N_4168,N_3977);
xnor U4413 (N_4413,N_4077,N_4141);
nor U4414 (N_4414,N_4187,N_4177);
xor U4415 (N_4415,N_4096,N_3966);
or U4416 (N_4416,N_3917,N_3903);
xnor U4417 (N_4417,N_4117,N_4101);
or U4418 (N_4418,N_4183,N_3992);
nand U4419 (N_4419,N_4072,N_4107);
or U4420 (N_4420,N_3982,N_4069);
and U4421 (N_4421,N_4067,N_3940);
and U4422 (N_4422,N_4153,N_3953);
and U4423 (N_4423,N_4121,N_3996);
or U4424 (N_4424,N_4046,N_3938);
and U4425 (N_4425,N_3938,N_4033);
nor U4426 (N_4426,N_3937,N_4006);
nand U4427 (N_4427,N_4169,N_3902);
nor U4428 (N_4428,N_3900,N_4170);
xor U4429 (N_4429,N_3940,N_4165);
and U4430 (N_4430,N_4198,N_4106);
or U4431 (N_4431,N_4101,N_4194);
nand U4432 (N_4432,N_4140,N_4013);
and U4433 (N_4433,N_3978,N_4184);
nand U4434 (N_4434,N_4039,N_3904);
nand U4435 (N_4435,N_4181,N_4089);
xnor U4436 (N_4436,N_4008,N_4015);
nand U4437 (N_4437,N_4095,N_4140);
xor U4438 (N_4438,N_4026,N_3900);
nand U4439 (N_4439,N_3949,N_3920);
or U4440 (N_4440,N_4054,N_3911);
nand U4441 (N_4441,N_3918,N_4044);
and U4442 (N_4442,N_3962,N_4183);
or U4443 (N_4443,N_3955,N_3993);
nand U4444 (N_4444,N_3926,N_4188);
and U4445 (N_4445,N_3960,N_4071);
nor U4446 (N_4446,N_3990,N_3908);
nor U4447 (N_4447,N_4057,N_4011);
nand U4448 (N_4448,N_4064,N_4090);
or U4449 (N_4449,N_4179,N_3957);
or U4450 (N_4450,N_3936,N_3940);
nand U4451 (N_4451,N_3926,N_4029);
xor U4452 (N_4452,N_3943,N_3990);
nand U4453 (N_4453,N_4160,N_3944);
or U4454 (N_4454,N_4192,N_3994);
nand U4455 (N_4455,N_3901,N_3965);
or U4456 (N_4456,N_4171,N_3959);
or U4457 (N_4457,N_4076,N_3939);
nand U4458 (N_4458,N_3942,N_3929);
xnor U4459 (N_4459,N_4106,N_3998);
nand U4460 (N_4460,N_3998,N_3982);
xor U4461 (N_4461,N_4021,N_3906);
nand U4462 (N_4462,N_4123,N_3965);
xnor U4463 (N_4463,N_3933,N_3935);
nor U4464 (N_4464,N_4056,N_3916);
or U4465 (N_4465,N_3903,N_4075);
and U4466 (N_4466,N_4114,N_3998);
or U4467 (N_4467,N_3989,N_4056);
xor U4468 (N_4468,N_4036,N_4007);
or U4469 (N_4469,N_4185,N_4148);
nor U4470 (N_4470,N_4174,N_4054);
or U4471 (N_4471,N_4068,N_4039);
nor U4472 (N_4472,N_4111,N_4151);
xor U4473 (N_4473,N_3989,N_4030);
and U4474 (N_4474,N_3911,N_4170);
nor U4475 (N_4475,N_4111,N_4138);
xnor U4476 (N_4476,N_3955,N_3938);
xor U4477 (N_4477,N_4148,N_4147);
xor U4478 (N_4478,N_3903,N_3960);
and U4479 (N_4479,N_4147,N_4170);
or U4480 (N_4480,N_4094,N_4025);
or U4481 (N_4481,N_4091,N_4066);
or U4482 (N_4482,N_4178,N_4043);
xnor U4483 (N_4483,N_4095,N_4176);
nand U4484 (N_4484,N_4058,N_4173);
nor U4485 (N_4485,N_3946,N_4084);
nor U4486 (N_4486,N_4186,N_3938);
and U4487 (N_4487,N_4073,N_3933);
nand U4488 (N_4488,N_3900,N_4199);
nor U4489 (N_4489,N_4099,N_4112);
or U4490 (N_4490,N_4006,N_3996);
nor U4491 (N_4491,N_3984,N_4006);
and U4492 (N_4492,N_4061,N_3964);
nor U4493 (N_4493,N_3960,N_4198);
or U4494 (N_4494,N_4191,N_4014);
xor U4495 (N_4495,N_4128,N_4074);
or U4496 (N_4496,N_3909,N_3932);
nand U4497 (N_4497,N_4164,N_4048);
or U4498 (N_4498,N_4158,N_4108);
or U4499 (N_4499,N_4039,N_4128);
nand U4500 (N_4500,N_4209,N_4319);
and U4501 (N_4501,N_4301,N_4421);
and U4502 (N_4502,N_4461,N_4413);
xnor U4503 (N_4503,N_4239,N_4351);
nor U4504 (N_4504,N_4419,N_4369);
nor U4505 (N_4505,N_4485,N_4360);
nor U4506 (N_4506,N_4221,N_4252);
xor U4507 (N_4507,N_4352,N_4288);
or U4508 (N_4508,N_4247,N_4225);
xnor U4509 (N_4509,N_4498,N_4346);
xnor U4510 (N_4510,N_4431,N_4425);
nand U4511 (N_4511,N_4276,N_4202);
xor U4512 (N_4512,N_4244,N_4359);
nor U4513 (N_4513,N_4255,N_4416);
xor U4514 (N_4514,N_4430,N_4483);
or U4515 (N_4515,N_4312,N_4365);
xnor U4516 (N_4516,N_4337,N_4249);
nand U4517 (N_4517,N_4242,N_4408);
or U4518 (N_4518,N_4227,N_4281);
xor U4519 (N_4519,N_4257,N_4208);
xor U4520 (N_4520,N_4477,N_4395);
xnor U4521 (N_4521,N_4275,N_4349);
nand U4522 (N_4522,N_4488,N_4348);
nor U4523 (N_4523,N_4353,N_4471);
or U4524 (N_4524,N_4380,N_4424);
xor U4525 (N_4525,N_4320,N_4458);
nand U4526 (N_4526,N_4334,N_4279);
or U4527 (N_4527,N_4292,N_4377);
or U4528 (N_4528,N_4266,N_4315);
nor U4529 (N_4529,N_4495,N_4381);
or U4530 (N_4530,N_4434,N_4466);
xor U4531 (N_4531,N_4364,N_4305);
xnor U4532 (N_4532,N_4476,N_4340);
nand U4533 (N_4533,N_4243,N_4287);
nor U4534 (N_4534,N_4286,N_4330);
or U4535 (N_4535,N_4267,N_4251);
nor U4536 (N_4536,N_4248,N_4354);
and U4537 (N_4537,N_4259,N_4426);
or U4538 (N_4538,N_4390,N_4326);
and U4539 (N_4539,N_4236,N_4270);
nor U4540 (N_4540,N_4378,N_4428);
and U4541 (N_4541,N_4423,N_4448);
and U4542 (N_4542,N_4432,N_4379);
nand U4543 (N_4543,N_4333,N_4284);
xor U4544 (N_4544,N_4226,N_4499);
or U4545 (N_4545,N_4382,N_4258);
and U4546 (N_4546,N_4289,N_4433);
xnor U4547 (N_4547,N_4232,N_4366);
nand U4548 (N_4548,N_4456,N_4472);
xor U4549 (N_4549,N_4293,N_4399);
nor U4550 (N_4550,N_4435,N_4216);
xor U4551 (N_4551,N_4262,N_4487);
or U4552 (N_4552,N_4411,N_4321);
or U4553 (N_4553,N_4250,N_4205);
and U4554 (N_4554,N_4338,N_4478);
and U4555 (N_4555,N_4318,N_4441);
and U4556 (N_4556,N_4278,N_4297);
and U4557 (N_4557,N_4410,N_4260);
xnor U4558 (N_4558,N_4218,N_4264);
and U4559 (N_4559,N_4482,N_4357);
nor U4560 (N_4560,N_4223,N_4463);
and U4561 (N_4561,N_4265,N_4462);
xnor U4562 (N_4562,N_4316,N_4392);
nor U4563 (N_4563,N_4263,N_4491);
and U4564 (N_4564,N_4389,N_4234);
xor U4565 (N_4565,N_4212,N_4460);
or U4566 (N_4566,N_4210,N_4347);
nand U4567 (N_4567,N_4299,N_4361);
and U4568 (N_4568,N_4325,N_4474);
nand U4569 (N_4569,N_4317,N_4256);
xnor U4570 (N_4570,N_4277,N_4261);
xor U4571 (N_4571,N_4231,N_4489);
nand U4572 (N_4572,N_4345,N_4385);
or U4573 (N_4573,N_4343,N_4412);
and U4574 (N_4574,N_4497,N_4233);
nor U4575 (N_4575,N_4417,N_4329);
and U4576 (N_4576,N_4291,N_4418);
xnor U4577 (N_4577,N_4407,N_4387);
xnor U4578 (N_4578,N_4254,N_4207);
xor U4579 (N_4579,N_4335,N_4304);
xnor U4580 (N_4580,N_4375,N_4484);
xnor U4581 (N_4581,N_4269,N_4447);
xnor U4582 (N_4582,N_4341,N_4427);
nor U4583 (N_4583,N_4420,N_4450);
or U4584 (N_4584,N_4213,N_4440);
xor U4585 (N_4585,N_4444,N_4229);
and U4586 (N_4586,N_4309,N_4394);
xor U4587 (N_4587,N_4453,N_4300);
nand U4588 (N_4588,N_4451,N_4356);
and U4589 (N_4589,N_4211,N_4268);
nor U4590 (N_4590,N_4469,N_4457);
nor U4591 (N_4591,N_4459,N_4400);
nand U4592 (N_4592,N_4238,N_4245);
nor U4593 (N_4593,N_4342,N_4465);
xor U4594 (N_4594,N_4401,N_4355);
or U4595 (N_4595,N_4443,N_4396);
or U4596 (N_4596,N_4405,N_4228);
or U4597 (N_4597,N_4295,N_4328);
nor U4598 (N_4598,N_4336,N_4403);
nor U4599 (N_4599,N_4473,N_4429);
or U4600 (N_4600,N_4445,N_4310);
nand U4601 (N_4601,N_4294,N_4449);
nor U4602 (N_4602,N_4303,N_4439);
or U4603 (N_4603,N_4271,N_4383);
nand U4604 (N_4604,N_4308,N_4496);
or U4605 (N_4605,N_4367,N_4393);
or U4606 (N_4606,N_4398,N_4214);
xnor U4607 (N_4607,N_4282,N_4368);
nand U4608 (N_4608,N_4493,N_4344);
nand U4609 (N_4609,N_4220,N_4215);
nand U4610 (N_4610,N_4224,N_4492);
nor U4611 (N_4611,N_4467,N_4422);
or U4612 (N_4612,N_4388,N_4332);
or U4613 (N_4613,N_4339,N_4376);
or U4614 (N_4614,N_4241,N_4217);
xor U4615 (N_4615,N_4222,N_4290);
nand U4616 (N_4616,N_4322,N_4363);
and U4617 (N_4617,N_4273,N_4454);
xnor U4618 (N_4618,N_4311,N_4203);
or U4619 (N_4619,N_4285,N_4442);
or U4620 (N_4620,N_4272,N_4253);
and U4621 (N_4621,N_4404,N_4206);
or U4622 (N_4622,N_4490,N_4494);
nor U4623 (N_4623,N_4362,N_4437);
or U4624 (N_4624,N_4237,N_4280);
and U4625 (N_4625,N_4470,N_4274);
or U4626 (N_4626,N_4386,N_4371);
nor U4627 (N_4627,N_4464,N_4452);
nor U4628 (N_4628,N_4415,N_4324);
and U4629 (N_4629,N_4372,N_4327);
nand U4630 (N_4630,N_4246,N_4350);
or U4631 (N_4631,N_4374,N_4313);
or U4632 (N_4632,N_4200,N_4323);
nor U4633 (N_4633,N_4201,N_4283);
or U4634 (N_4634,N_4302,N_4240);
nand U4635 (N_4635,N_4235,N_4314);
or U4636 (N_4636,N_4397,N_4406);
nand U4637 (N_4637,N_4414,N_4391);
nand U4638 (N_4638,N_4446,N_4455);
nand U4639 (N_4639,N_4409,N_4298);
xor U4640 (N_4640,N_4296,N_4307);
or U4641 (N_4641,N_4384,N_4480);
nor U4642 (N_4642,N_4230,N_4436);
and U4643 (N_4643,N_4219,N_4331);
and U4644 (N_4644,N_4204,N_4373);
xnor U4645 (N_4645,N_4370,N_4402);
or U4646 (N_4646,N_4486,N_4438);
and U4647 (N_4647,N_4481,N_4306);
nand U4648 (N_4648,N_4479,N_4468);
nor U4649 (N_4649,N_4358,N_4475);
nand U4650 (N_4650,N_4418,N_4448);
nor U4651 (N_4651,N_4309,N_4289);
nand U4652 (N_4652,N_4364,N_4259);
nand U4653 (N_4653,N_4404,N_4289);
nor U4654 (N_4654,N_4324,N_4318);
nor U4655 (N_4655,N_4263,N_4360);
and U4656 (N_4656,N_4468,N_4351);
nand U4657 (N_4657,N_4444,N_4326);
or U4658 (N_4658,N_4412,N_4241);
xor U4659 (N_4659,N_4253,N_4216);
and U4660 (N_4660,N_4314,N_4477);
nand U4661 (N_4661,N_4361,N_4480);
nand U4662 (N_4662,N_4389,N_4358);
or U4663 (N_4663,N_4330,N_4432);
and U4664 (N_4664,N_4496,N_4383);
nor U4665 (N_4665,N_4470,N_4391);
xor U4666 (N_4666,N_4324,N_4329);
and U4667 (N_4667,N_4297,N_4391);
and U4668 (N_4668,N_4314,N_4356);
and U4669 (N_4669,N_4382,N_4491);
or U4670 (N_4670,N_4467,N_4203);
xor U4671 (N_4671,N_4383,N_4297);
xnor U4672 (N_4672,N_4312,N_4317);
nand U4673 (N_4673,N_4402,N_4321);
and U4674 (N_4674,N_4311,N_4231);
xor U4675 (N_4675,N_4366,N_4242);
or U4676 (N_4676,N_4234,N_4418);
or U4677 (N_4677,N_4255,N_4231);
nor U4678 (N_4678,N_4400,N_4366);
xor U4679 (N_4679,N_4373,N_4464);
and U4680 (N_4680,N_4437,N_4340);
nor U4681 (N_4681,N_4401,N_4379);
nand U4682 (N_4682,N_4273,N_4226);
and U4683 (N_4683,N_4214,N_4244);
nand U4684 (N_4684,N_4229,N_4411);
and U4685 (N_4685,N_4238,N_4435);
nor U4686 (N_4686,N_4475,N_4472);
or U4687 (N_4687,N_4456,N_4387);
or U4688 (N_4688,N_4451,N_4478);
nor U4689 (N_4689,N_4254,N_4397);
and U4690 (N_4690,N_4313,N_4309);
nand U4691 (N_4691,N_4360,N_4232);
nor U4692 (N_4692,N_4260,N_4378);
nor U4693 (N_4693,N_4469,N_4249);
xor U4694 (N_4694,N_4415,N_4335);
or U4695 (N_4695,N_4393,N_4362);
or U4696 (N_4696,N_4496,N_4317);
and U4697 (N_4697,N_4264,N_4293);
and U4698 (N_4698,N_4482,N_4346);
nand U4699 (N_4699,N_4268,N_4462);
and U4700 (N_4700,N_4411,N_4268);
or U4701 (N_4701,N_4297,N_4416);
or U4702 (N_4702,N_4438,N_4404);
nand U4703 (N_4703,N_4397,N_4342);
nor U4704 (N_4704,N_4461,N_4425);
nor U4705 (N_4705,N_4492,N_4403);
or U4706 (N_4706,N_4413,N_4203);
and U4707 (N_4707,N_4393,N_4285);
or U4708 (N_4708,N_4338,N_4212);
and U4709 (N_4709,N_4381,N_4451);
nor U4710 (N_4710,N_4429,N_4484);
xnor U4711 (N_4711,N_4314,N_4439);
xor U4712 (N_4712,N_4403,N_4431);
nand U4713 (N_4713,N_4273,N_4258);
xnor U4714 (N_4714,N_4201,N_4342);
or U4715 (N_4715,N_4219,N_4469);
xnor U4716 (N_4716,N_4243,N_4416);
or U4717 (N_4717,N_4292,N_4243);
xnor U4718 (N_4718,N_4380,N_4301);
or U4719 (N_4719,N_4446,N_4200);
nor U4720 (N_4720,N_4414,N_4260);
xor U4721 (N_4721,N_4488,N_4491);
nor U4722 (N_4722,N_4363,N_4494);
nor U4723 (N_4723,N_4476,N_4380);
xnor U4724 (N_4724,N_4432,N_4282);
xor U4725 (N_4725,N_4380,N_4256);
xnor U4726 (N_4726,N_4260,N_4352);
nand U4727 (N_4727,N_4464,N_4363);
nand U4728 (N_4728,N_4407,N_4442);
xor U4729 (N_4729,N_4284,N_4467);
nand U4730 (N_4730,N_4250,N_4319);
and U4731 (N_4731,N_4497,N_4381);
or U4732 (N_4732,N_4369,N_4246);
nor U4733 (N_4733,N_4400,N_4206);
nor U4734 (N_4734,N_4463,N_4317);
nand U4735 (N_4735,N_4317,N_4388);
nand U4736 (N_4736,N_4411,N_4261);
nand U4737 (N_4737,N_4444,N_4376);
xor U4738 (N_4738,N_4400,N_4214);
nand U4739 (N_4739,N_4430,N_4426);
nand U4740 (N_4740,N_4398,N_4303);
nor U4741 (N_4741,N_4477,N_4244);
xor U4742 (N_4742,N_4252,N_4255);
xnor U4743 (N_4743,N_4372,N_4437);
and U4744 (N_4744,N_4411,N_4224);
nor U4745 (N_4745,N_4336,N_4445);
nor U4746 (N_4746,N_4485,N_4441);
nor U4747 (N_4747,N_4316,N_4375);
and U4748 (N_4748,N_4343,N_4229);
nor U4749 (N_4749,N_4432,N_4492);
nor U4750 (N_4750,N_4215,N_4428);
nand U4751 (N_4751,N_4438,N_4223);
nor U4752 (N_4752,N_4265,N_4491);
or U4753 (N_4753,N_4445,N_4295);
nor U4754 (N_4754,N_4420,N_4269);
xor U4755 (N_4755,N_4369,N_4248);
nor U4756 (N_4756,N_4302,N_4443);
or U4757 (N_4757,N_4253,N_4262);
nand U4758 (N_4758,N_4454,N_4296);
and U4759 (N_4759,N_4217,N_4301);
xnor U4760 (N_4760,N_4276,N_4398);
or U4761 (N_4761,N_4354,N_4477);
nand U4762 (N_4762,N_4230,N_4327);
nand U4763 (N_4763,N_4205,N_4396);
nand U4764 (N_4764,N_4280,N_4404);
or U4765 (N_4765,N_4246,N_4490);
nor U4766 (N_4766,N_4465,N_4221);
or U4767 (N_4767,N_4487,N_4473);
or U4768 (N_4768,N_4282,N_4443);
and U4769 (N_4769,N_4364,N_4311);
nand U4770 (N_4770,N_4329,N_4436);
or U4771 (N_4771,N_4354,N_4266);
nor U4772 (N_4772,N_4205,N_4323);
nand U4773 (N_4773,N_4413,N_4404);
nand U4774 (N_4774,N_4251,N_4226);
and U4775 (N_4775,N_4304,N_4391);
and U4776 (N_4776,N_4468,N_4373);
nor U4777 (N_4777,N_4484,N_4225);
or U4778 (N_4778,N_4259,N_4249);
or U4779 (N_4779,N_4383,N_4402);
and U4780 (N_4780,N_4412,N_4335);
nor U4781 (N_4781,N_4231,N_4461);
or U4782 (N_4782,N_4409,N_4312);
or U4783 (N_4783,N_4419,N_4203);
nor U4784 (N_4784,N_4219,N_4307);
or U4785 (N_4785,N_4432,N_4320);
xor U4786 (N_4786,N_4302,N_4259);
nand U4787 (N_4787,N_4206,N_4208);
nor U4788 (N_4788,N_4349,N_4497);
xnor U4789 (N_4789,N_4203,N_4245);
nand U4790 (N_4790,N_4353,N_4394);
xor U4791 (N_4791,N_4256,N_4226);
nand U4792 (N_4792,N_4494,N_4472);
and U4793 (N_4793,N_4380,N_4223);
xor U4794 (N_4794,N_4462,N_4391);
nand U4795 (N_4795,N_4347,N_4325);
xnor U4796 (N_4796,N_4352,N_4462);
xor U4797 (N_4797,N_4232,N_4458);
nand U4798 (N_4798,N_4289,N_4429);
nor U4799 (N_4799,N_4312,N_4465);
xor U4800 (N_4800,N_4536,N_4684);
nor U4801 (N_4801,N_4560,N_4688);
or U4802 (N_4802,N_4517,N_4769);
xnor U4803 (N_4803,N_4544,N_4683);
nor U4804 (N_4804,N_4547,N_4647);
nand U4805 (N_4805,N_4537,N_4749);
nor U4806 (N_4806,N_4739,N_4648);
nand U4807 (N_4807,N_4759,N_4670);
nor U4808 (N_4808,N_4755,N_4539);
xor U4809 (N_4809,N_4658,N_4766);
xor U4810 (N_4810,N_4611,N_4543);
and U4811 (N_4811,N_4607,N_4520);
or U4812 (N_4812,N_4643,N_4770);
xor U4813 (N_4813,N_4518,N_4660);
xnor U4814 (N_4814,N_4720,N_4525);
nor U4815 (N_4815,N_4619,N_4712);
nor U4816 (N_4816,N_4602,N_4693);
and U4817 (N_4817,N_4592,N_4620);
nand U4818 (N_4818,N_4733,N_4638);
and U4819 (N_4819,N_4600,N_4776);
nand U4820 (N_4820,N_4781,N_4758);
nand U4821 (N_4821,N_4663,N_4651);
xnor U4822 (N_4822,N_4687,N_4504);
nor U4823 (N_4823,N_4669,N_4700);
and U4824 (N_4824,N_4737,N_4787);
nand U4825 (N_4825,N_4696,N_4586);
nand U4826 (N_4826,N_4774,N_4747);
or U4827 (N_4827,N_4532,N_4514);
nand U4828 (N_4828,N_4513,N_4574);
and U4829 (N_4829,N_4576,N_4634);
nor U4830 (N_4830,N_4557,N_4545);
or U4831 (N_4831,N_4605,N_4784);
or U4832 (N_4832,N_4778,N_4569);
xor U4833 (N_4833,N_4640,N_4649);
or U4834 (N_4834,N_4705,N_4673);
or U4835 (N_4835,N_4555,N_4780);
and U4836 (N_4836,N_4568,N_4501);
and U4837 (N_4837,N_4637,N_4527);
and U4838 (N_4838,N_4727,N_4535);
or U4839 (N_4839,N_4507,N_4762);
and U4840 (N_4840,N_4551,N_4612);
or U4841 (N_4841,N_4718,N_4521);
and U4842 (N_4842,N_4799,N_4742);
and U4843 (N_4843,N_4571,N_4548);
and U4844 (N_4844,N_4515,N_4645);
xor U4845 (N_4845,N_4666,N_4579);
xnor U4846 (N_4846,N_4782,N_4785);
nor U4847 (N_4847,N_4661,N_4724);
and U4848 (N_4848,N_4655,N_4790);
xor U4849 (N_4849,N_4764,N_4662);
or U4850 (N_4850,N_4546,N_4624);
nand U4851 (N_4851,N_4697,N_4756);
and U4852 (N_4852,N_4563,N_4786);
nand U4853 (N_4853,N_4503,N_4511);
nand U4854 (N_4854,N_4795,N_4614);
and U4855 (N_4855,N_4589,N_4702);
and U4856 (N_4856,N_4601,N_4797);
nor U4857 (N_4857,N_4652,N_4584);
xnor U4858 (N_4858,N_4644,N_4646);
nand U4859 (N_4859,N_4711,N_4523);
or U4860 (N_4860,N_4744,N_4665);
nand U4861 (N_4861,N_4567,N_4676);
or U4862 (N_4862,N_4509,N_4659);
nor U4863 (N_4863,N_4768,N_4668);
nand U4864 (N_4864,N_4765,N_4510);
nor U4865 (N_4865,N_4623,N_4533);
and U4866 (N_4866,N_4577,N_4740);
nand U4867 (N_4867,N_4783,N_4512);
or U4868 (N_4868,N_4708,N_4570);
nor U4869 (N_4869,N_4717,N_4671);
xor U4870 (N_4870,N_4657,N_4745);
or U4871 (N_4871,N_4541,N_4595);
or U4872 (N_4872,N_4604,N_4751);
or U4873 (N_4873,N_4788,N_4679);
and U4874 (N_4874,N_4641,N_4771);
nand U4875 (N_4875,N_4729,N_4752);
or U4876 (N_4876,N_4738,N_4534);
nand U4877 (N_4877,N_4538,N_4627);
nor U4878 (N_4878,N_4722,N_4698);
nand U4879 (N_4879,N_4672,N_4713);
nor U4880 (N_4880,N_4508,N_4691);
xor U4881 (N_4881,N_4714,N_4581);
xnor U4882 (N_4882,N_4734,N_4767);
xor U4883 (N_4883,N_4599,N_4617);
nor U4884 (N_4884,N_4726,N_4591);
nand U4885 (N_4885,N_4542,N_4593);
and U4886 (N_4886,N_4685,N_4789);
nor U4887 (N_4887,N_4753,N_4674);
and U4888 (N_4888,N_4585,N_4716);
or U4889 (N_4889,N_4632,N_4594);
nand U4890 (N_4890,N_4692,N_4530);
nor U4891 (N_4891,N_4572,N_4522);
or U4892 (N_4892,N_4610,N_4709);
or U4893 (N_4893,N_4606,N_4682);
nor U4894 (N_4894,N_4629,N_4502);
or U4895 (N_4895,N_4754,N_4675);
xor U4896 (N_4896,N_4553,N_4615);
nand U4897 (N_4897,N_4621,N_4562);
xnor U4898 (N_4898,N_4519,N_4796);
or U4899 (N_4899,N_4772,N_4625);
and U4900 (N_4900,N_4635,N_4680);
nand U4901 (N_4901,N_4773,N_4793);
or U4902 (N_4902,N_4681,N_4794);
xor U4903 (N_4903,N_4609,N_4721);
or U4904 (N_4904,N_4703,N_4580);
or U4905 (N_4905,N_4775,N_4531);
xnor U4906 (N_4906,N_4642,N_4598);
and U4907 (N_4907,N_4761,N_4719);
and U4908 (N_4908,N_4706,N_4707);
xnor U4909 (N_4909,N_4516,N_4656);
and U4910 (N_4910,N_4779,N_4667);
and U4911 (N_4911,N_4686,N_4735);
nor U4912 (N_4912,N_4528,N_4622);
and U4913 (N_4913,N_4626,N_4583);
and U4914 (N_4914,N_4540,N_4777);
or U4915 (N_4915,N_4550,N_4728);
or U4916 (N_4916,N_4603,N_4613);
nand U4917 (N_4917,N_4588,N_4798);
xor U4918 (N_4918,N_4500,N_4616);
and U4919 (N_4919,N_4561,N_4582);
xnor U4920 (N_4920,N_4549,N_4630);
xor U4921 (N_4921,N_4763,N_4618);
or U4922 (N_4922,N_4732,N_4701);
nor U4923 (N_4923,N_4566,N_4608);
nand U4924 (N_4924,N_4636,N_4597);
or U4925 (N_4925,N_4596,N_4699);
nor U4926 (N_4926,N_4748,N_4746);
or U4927 (N_4927,N_4524,N_4715);
nand U4928 (N_4928,N_4639,N_4505);
or U4929 (N_4929,N_4578,N_4730);
and U4930 (N_4930,N_4565,N_4633);
nor U4931 (N_4931,N_4506,N_4760);
nor U4932 (N_4932,N_4757,N_4694);
nand U4933 (N_4933,N_4587,N_4654);
nand U4934 (N_4934,N_4791,N_4723);
or U4935 (N_4935,N_4690,N_4559);
nor U4936 (N_4936,N_4556,N_4689);
nor U4937 (N_4937,N_4573,N_4575);
nor U4938 (N_4938,N_4558,N_4750);
xor U4939 (N_4939,N_4710,N_4695);
xnor U4940 (N_4940,N_4529,N_4631);
nor U4941 (N_4941,N_4731,N_4792);
xnor U4942 (N_4942,N_4650,N_4743);
nand U4943 (N_4943,N_4677,N_4526);
and U4944 (N_4944,N_4704,N_4628);
and U4945 (N_4945,N_4736,N_4554);
nor U4946 (N_4946,N_4741,N_4678);
xor U4947 (N_4947,N_4664,N_4564);
nor U4948 (N_4948,N_4590,N_4725);
nand U4949 (N_4949,N_4653,N_4552);
nand U4950 (N_4950,N_4651,N_4619);
and U4951 (N_4951,N_4552,N_4615);
xor U4952 (N_4952,N_4632,N_4780);
xnor U4953 (N_4953,N_4544,N_4643);
and U4954 (N_4954,N_4715,N_4784);
nor U4955 (N_4955,N_4546,N_4562);
nand U4956 (N_4956,N_4635,N_4647);
nand U4957 (N_4957,N_4727,N_4642);
nor U4958 (N_4958,N_4725,N_4782);
and U4959 (N_4959,N_4639,N_4574);
nor U4960 (N_4960,N_4653,N_4521);
xor U4961 (N_4961,N_4626,N_4744);
and U4962 (N_4962,N_4581,N_4626);
or U4963 (N_4963,N_4761,N_4581);
and U4964 (N_4964,N_4772,N_4767);
xor U4965 (N_4965,N_4731,N_4700);
nor U4966 (N_4966,N_4726,N_4577);
nand U4967 (N_4967,N_4653,N_4775);
and U4968 (N_4968,N_4620,N_4644);
and U4969 (N_4969,N_4744,N_4696);
or U4970 (N_4970,N_4663,N_4737);
or U4971 (N_4971,N_4523,N_4736);
and U4972 (N_4972,N_4547,N_4797);
and U4973 (N_4973,N_4546,N_4740);
nand U4974 (N_4974,N_4732,N_4611);
xnor U4975 (N_4975,N_4715,N_4723);
xnor U4976 (N_4976,N_4586,N_4625);
nor U4977 (N_4977,N_4697,N_4644);
nor U4978 (N_4978,N_4729,N_4777);
and U4979 (N_4979,N_4791,N_4522);
or U4980 (N_4980,N_4610,N_4769);
nor U4981 (N_4981,N_4708,N_4761);
xnor U4982 (N_4982,N_4693,N_4671);
nand U4983 (N_4983,N_4622,N_4731);
or U4984 (N_4984,N_4524,N_4686);
nand U4985 (N_4985,N_4796,N_4556);
xor U4986 (N_4986,N_4668,N_4587);
or U4987 (N_4987,N_4639,N_4625);
and U4988 (N_4988,N_4678,N_4639);
or U4989 (N_4989,N_4677,N_4603);
nor U4990 (N_4990,N_4784,N_4535);
and U4991 (N_4991,N_4623,N_4571);
or U4992 (N_4992,N_4658,N_4566);
xor U4993 (N_4993,N_4646,N_4555);
or U4994 (N_4994,N_4659,N_4721);
nand U4995 (N_4995,N_4666,N_4525);
nor U4996 (N_4996,N_4704,N_4667);
xnor U4997 (N_4997,N_4585,N_4534);
xor U4998 (N_4998,N_4588,N_4632);
or U4999 (N_4999,N_4696,N_4689);
nor U5000 (N_5000,N_4682,N_4623);
nor U5001 (N_5001,N_4750,N_4771);
and U5002 (N_5002,N_4714,N_4569);
nand U5003 (N_5003,N_4736,N_4752);
or U5004 (N_5004,N_4536,N_4798);
and U5005 (N_5005,N_4555,N_4503);
xor U5006 (N_5006,N_4628,N_4748);
nand U5007 (N_5007,N_4611,N_4521);
xnor U5008 (N_5008,N_4668,N_4730);
nand U5009 (N_5009,N_4734,N_4729);
and U5010 (N_5010,N_4781,N_4667);
or U5011 (N_5011,N_4599,N_4589);
nor U5012 (N_5012,N_4627,N_4672);
and U5013 (N_5013,N_4526,N_4734);
nand U5014 (N_5014,N_4517,N_4504);
and U5015 (N_5015,N_4795,N_4562);
nand U5016 (N_5016,N_4546,N_4650);
or U5017 (N_5017,N_4637,N_4592);
nor U5018 (N_5018,N_4557,N_4585);
nand U5019 (N_5019,N_4777,N_4618);
and U5020 (N_5020,N_4761,N_4676);
or U5021 (N_5021,N_4512,N_4680);
xnor U5022 (N_5022,N_4665,N_4758);
nor U5023 (N_5023,N_4723,N_4579);
xor U5024 (N_5024,N_4762,N_4654);
or U5025 (N_5025,N_4707,N_4642);
or U5026 (N_5026,N_4646,N_4527);
nor U5027 (N_5027,N_4758,N_4776);
and U5028 (N_5028,N_4706,N_4682);
nor U5029 (N_5029,N_4762,N_4566);
xor U5030 (N_5030,N_4616,N_4672);
nor U5031 (N_5031,N_4663,N_4669);
xnor U5032 (N_5032,N_4666,N_4518);
or U5033 (N_5033,N_4502,N_4624);
and U5034 (N_5034,N_4790,N_4695);
xnor U5035 (N_5035,N_4695,N_4573);
nor U5036 (N_5036,N_4643,N_4525);
xor U5037 (N_5037,N_4557,N_4796);
nor U5038 (N_5038,N_4792,N_4544);
nand U5039 (N_5039,N_4738,N_4630);
nor U5040 (N_5040,N_4559,N_4740);
nand U5041 (N_5041,N_4554,N_4584);
and U5042 (N_5042,N_4574,N_4528);
xor U5043 (N_5043,N_4678,N_4709);
nand U5044 (N_5044,N_4799,N_4696);
or U5045 (N_5045,N_4519,N_4625);
or U5046 (N_5046,N_4681,N_4727);
xor U5047 (N_5047,N_4707,N_4725);
xor U5048 (N_5048,N_4687,N_4556);
and U5049 (N_5049,N_4752,N_4669);
or U5050 (N_5050,N_4763,N_4743);
nand U5051 (N_5051,N_4603,N_4621);
xor U5052 (N_5052,N_4552,N_4721);
nor U5053 (N_5053,N_4629,N_4727);
nor U5054 (N_5054,N_4574,N_4669);
and U5055 (N_5055,N_4752,N_4758);
and U5056 (N_5056,N_4700,N_4595);
and U5057 (N_5057,N_4791,N_4521);
xnor U5058 (N_5058,N_4556,N_4502);
nor U5059 (N_5059,N_4742,N_4559);
and U5060 (N_5060,N_4764,N_4610);
xnor U5061 (N_5061,N_4668,N_4763);
and U5062 (N_5062,N_4502,N_4788);
nand U5063 (N_5063,N_4517,N_4605);
xor U5064 (N_5064,N_4529,N_4758);
xnor U5065 (N_5065,N_4544,N_4634);
nor U5066 (N_5066,N_4659,N_4573);
and U5067 (N_5067,N_4701,N_4503);
and U5068 (N_5068,N_4650,N_4672);
or U5069 (N_5069,N_4746,N_4500);
or U5070 (N_5070,N_4604,N_4734);
nand U5071 (N_5071,N_4759,N_4673);
nor U5072 (N_5072,N_4527,N_4763);
xor U5073 (N_5073,N_4658,N_4651);
and U5074 (N_5074,N_4504,N_4787);
nor U5075 (N_5075,N_4556,N_4626);
nand U5076 (N_5076,N_4748,N_4505);
nand U5077 (N_5077,N_4717,N_4573);
and U5078 (N_5078,N_4564,N_4524);
xnor U5079 (N_5079,N_4684,N_4667);
or U5080 (N_5080,N_4620,N_4654);
nand U5081 (N_5081,N_4516,N_4720);
xor U5082 (N_5082,N_4660,N_4639);
xnor U5083 (N_5083,N_4512,N_4572);
or U5084 (N_5084,N_4657,N_4689);
xor U5085 (N_5085,N_4636,N_4701);
xnor U5086 (N_5086,N_4664,N_4686);
and U5087 (N_5087,N_4783,N_4774);
xnor U5088 (N_5088,N_4541,N_4528);
and U5089 (N_5089,N_4556,N_4654);
nor U5090 (N_5090,N_4612,N_4555);
nand U5091 (N_5091,N_4669,N_4711);
or U5092 (N_5092,N_4727,N_4785);
or U5093 (N_5093,N_4687,N_4564);
or U5094 (N_5094,N_4784,N_4729);
or U5095 (N_5095,N_4689,N_4511);
or U5096 (N_5096,N_4539,N_4579);
xnor U5097 (N_5097,N_4771,N_4788);
xnor U5098 (N_5098,N_4785,N_4647);
nand U5099 (N_5099,N_4657,N_4607);
nand U5100 (N_5100,N_4834,N_4922);
nor U5101 (N_5101,N_4883,N_5061);
and U5102 (N_5102,N_4837,N_4844);
nand U5103 (N_5103,N_5076,N_5043);
nor U5104 (N_5104,N_4979,N_4890);
or U5105 (N_5105,N_4963,N_4929);
nand U5106 (N_5106,N_5028,N_4868);
xnor U5107 (N_5107,N_5044,N_4820);
nor U5108 (N_5108,N_5010,N_4931);
xnor U5109 (N_5109,N_4977,N_4826);
xnor U5110 (N_5110,N_5016,N_4809);
and U5111 (N_5111,N_4892,N_5069);
nand U5112 (N_5112,N_4864,N_4806);
and U5113 (N_5113,N_5032,N_5045);
xnor U5114 (N_5114,N_4999,N_5097);
nor U5115 (N_5115,N_4872,N_4901);
and U5116 (N_5116,N_5006,N_5053);
and U5117 (N_5117,N_5077,N_4807);
and U5118 (N_5118,N_4866,N_4930);
and U5119 (N_5119,N_4902,N_4849);
xor U5120 (N_5120,N_4874,N_4813);
or U5121 (N_5121,N_4989,N_5040);
or U5122 (N_5122,N_4921,N_5056);
nor U5123 (N_5123,N_4869,N_5064);
xnor U5124 (N_5124,N_4815,N_4986);
or U5125 (N_5125,N_4919,N_4926);
xnor U5126 (N_5126,N_5093,N_4908);
xnor U5127 (N_5127,N_4937,N_5081);
nor U5128 (N_5128,N_5018,N_5058);
and U5129 (N_5129,N_5059,N_4958);
and U5130 (N_5130,N_4915,N_4992);
nor U5131 (N_5131,N_4973,N_4862);
nor U5132 (N_5132,N_4842,N_4821);
or U5133 (N_5133,N_4932,N_5037);
xor U5134 (N_5134,N_5000,N_4832);
nand U5135 (N_5135,N_4917,N_4845);
xor U5136 (N_5136,N_4838,N_4893);
nand U5137 (N_5137,N_5070,N_5096);
nand U5138 (N_5138,N_4889,N_4853);
nor U5139 (N_5139,N_4810,N_5078);
xnor U5140 (N_5140,N_4985,N_4880);
nand U5141 (N_5141,N_4833,N_5080);
or U5142 (N_5142,N_5021,N_4903);
nand U5143 (N_5143,N_4897,N_5051);
nand U5144 (N_5144,N_5029,N_5013);
xor U5145 (N_5145,N_5079,N_5035);
nor U5146 (N_5146,N_4996,N_4942);
xnor U5147 (N_5147,N_4854,N_4819);
nor U5148 (N_5148,N_4995,N_4952);
or U5149 (N_5149,N_4863,N_4953);
xnor U5150 (N_5150,N_4873,N_4882);
nor U5151 (N_5151,N_4935,N_4961);
and U5152 (N_5152,N_4914,N_5022);
and U5153 (N_5153,N_4936,N_4877);
or U5154 (N_5154,N_5025,N_4885);
and U5155 (N_5155,N_5048,N_5020);
nor U5156 (N_5156,N_4924,N_4934);
nand U5157 (N_5157,N_4894,N_4907);
nor U5158 (N_5158,N_5039,N_4899);
xnor U5159 (N_5159,N_5094,N_4971);
nand U5160 (N_5160,N_5031,N_4804);
nand U5161 (N_5161,N_4841,N_4951);
or U5162 (N_5162,N_4997,N_5068);
or U5163 (N_5163,N_4801,N_4956);
and U5164 (N_5164,N_4895,N_5073);
and U5165 (N_5165,N_4876,N_4857);
xnor U5166 (N_5166,N_4925,N_4896);
and U5167 (N_5167,N_4949,N_4911);
and U5168 (N_5168,N_5015,N_4990);
nor U5169 (N_5169,N_4858,N_5047);
and U5170 (N_5170,N_4966,N_4982);
nor U5171 (N_5171,N_4984,N_5042);
or U5172 (N_5172,N_4861,N_5086);
xnor U5173 (N_5173,N_4847,N_4825);
xnor U5174 (N_5174,N_4927,N_5034);
or U5175 (N_5175,N_4916,N_4887);
nand U5176 (N_5176,N_5027,N_4960);
or U5177 (N_5177,N_4939,N_4957);
xnor U5178 (N_5178,N_5063,N_4822);
nor U5179 (N_5179,N_5055,N_4848);
nand U5180 (N_5180,N_4944,N_5007);
xnor U5181 (N_5181,N_4840,N_5092);
xor U5182 (N_5182,N_4867,N_4830);
xnor U5183 (N_5183,N_4886,N_4967);
xnor U5184 (N_5184,N_4905,N_4988);
or U5185 (N_5185,N_4817,N_4964);
nand U5186 (N_5186,N_4884,N_5074);
xor U5187 (N_5187,N_4969,N_4870);
or U5188 (N_5188,N_5099,N_5041);
nand U5189 (N_5189,N_4912,N_4846);
xor U5190 (N_5190,N_5002,N_5009);
and U5191 (N_5191,N_5030,N_4972);
and U5192 (N_5192,N_4976,N_4947);
and U5193 (N_5193,N_4965,N_4933);
nor U5194 (N_5194,N_4802,N_4943);
and U5195 (N_5195,N_4814,N_4856);
and U5196 (N_5196,N_4811,N_4835);
nor U5197 (N_5197,N_4998,N_5090);
or U5198 (N_5198,N_4987,N_5049);
and U5199 (N_5199,N_5017,N_4888);
nand U5200 (N_5200,N_4974,N_5089);
nand U5201 (N_5201,N_4991,N_5098);
xor U5202 (N_5202,N_5033,N_5065);
nand U5203 (N_5203,N_5024,N_4891);
and U5204 (N_5204,N_5008,N_4871);
or U5205 (N_5205,N_5003,N_4923);
nor U5206 (N_5206,N_5057,N_4975);
and U5207 (N_5207,N_5075,N_4818);
nor U5208 (N_5208,N_5062,N_4909);
or U5209 (N_5209,N_5087,N_5011);
nand U5210 (N_5210,N_4993,N_4968);
nand U5211 (N_5211,N_4962,N_5084);
nor U5212 (N_5212,N_4855,N_4828);
nand U5213 (N_5213,N_4865,N_4827);
and U5214 (N_5214,N_4829,N_4878);
nor U5215 (N_5215,N_4970,N_5072);
or U5216 (N_5216,N_4824,N_5060);
nor U5217 (N_5217,N_4839,N_5038);
xnor U5218 (N_5218,N_4803,N_5014);
or U5219 (N_5219,N_4852,N_4831);
nor U5220 (N_5220,N_4823,N_5001);
nor U5221 (N_5221,N_4859,N_5004);
and U5222 (N_5222,N_4941,N_5066);
and U5223 (N_5223,N_5026,N_4910);
or U5224 (N_5224,N_4816,N_4881);
nor U5225 (N_5225,N_4938,N_4805);
and U5226 (N_5226,N_4978,N_4950);
nand U5227 (N_5227,N_5012,N_5082);
nor U5228 (N_5228,N_4904,N_4980);
nand U5229 (N_5229,N_4808,N_4955);
xor U5230 (N_5230,N_4954,N_4812);
and U5231 (N_5231,N_5019,N_5083);
nor U5232 (N_5232,N_5088,N_4875);
nand U5233 (N_5233,N_4983,N_5067);
nand U5234 (N_5234,N_4994,N_5095);
nor U5235 (N_5235,N_5046,N_4913);
nor U5236 (N_5236,N_4948,N_4900);
nor U5237 (N_5237,N_4928,N_4800);
nor U5238 (N_5238,N_4920,N_5085);
xnor U5239 (N_5239,N_5050,N_4945);
nand U5240 (N_5240,N_5052,N_5071);
nand U5241 (N_5241,N_4860,N_4851);
or U5242 (N_5242,N_4879,N_5005);
nand U5243 (N_5243,N_5023,N_4843);
or U5244 (N_5244,N_4940,N_4959);
and U5245 (N_5245,N_4981,N_4946);
xnor U5246 (N_5246,N_5091,N_4850);
nor U5247 (N_5247,N_5054,N_4918);
and U5248 (N_5248,N_4898,N_5036);
nand U5249 (N_5249,N_4906,N_4836);
nor U5250 (N_5250,N_4976,N_4983);
and U5251 (N_5251,N_5002,N_4809);
nor U5252 (N_5252,N_4843,N_4862);
or U5253 (N_5253,N_4896,N_5029);
nor U5254 (N_5254,N_4963,N_4872);
or U5255 (N_5255,N_4836,N_4846);
nand U5256 (N_5256,N_4876,N_5053);
and U5257 (N_5257,N_5087,N_5001);
nor U5258 (N_5258,N_4912,N_4851);
nor U5259 (N_5259,N_4910,N_4848);
or U5260 (N_5260,N_4813,N_4982);
nor U5261 (N_5261,N_4898,N_4975);
nand U5262 (N_5262,N_5055,N_4967);
and U5263 (N_5263,N_4938,N_4833);
nand U5264 (N_5264,N_4862,N_5084);
or U5265 (N_5265,N_4976,N_5039);
and U5266 (N_5266,N_4882,N_5077);
or U5267 (N_5267,N_4956,N_5016);
and U5268 (N_5268,N_5021,N_5054);
or U5269 (N_5269,N_5046,N_4824);
xor U5270 (N_5270,N_4819,N_4977);
and U5271 (N_5271,N_5035,N_4948);
xnor U5272 (N_5272,N_4843,N_4959);
xor U5273 (N_5273,N_4870,N_4973);
xnor U5274 (N_5274,N_4885,N_5036);
xnor U5275 (N_5275,N_4989,N_4986);
xnor U5276 (N_5276,N_5016,N_5046);
or U5277 (N_5277,N_5081,N_5070);
and U5278 (N_5278,N_4928,N_4963);
or U5279 (N_5279,N_4822,N_4987);
nand U5280 (N_5280,N_5015,N_4856);
xnor U5281 (N_5281,N_5013,N_4887);
nand U5282 (N_5282,N_4938,N_4936);
or U5283 (N_5283,N_4915,N_4857);
xnor U5284 (N_5284,N_4826,N_4808);
nand U5285 (N_5285,N_4867,N_4910);
or U5286 (N_5286,N_4923,N_4846);
and U5287 (N_5287,N_4831,N_4833);
nor U5288 (N_5288,N_5022,N_4931);
and U5289 (N_5289,N_4945,N_4847);
nand U5290 (N_5290,N_4914,N_4905);
or U5291 (N_5291,N_5029,N_4884);
and U5292 (N_5292,N_5048,N_4890);
and U5293 (N_5293,N_5079,N_4855);
xor U5294 (N_5294,N_4852,N_4992);
nor U5295 (N_5295,N_4822,N_5024);
and U5296 (N_5296,N_5083,N_4915);
or U5297 (N_5297,N_4925,N_5065);
xnor U5298 (N_5298,N_4910,N_4801);
nand U5299 (N_5299,N_4875,N_4929);
nor U5300 (N_5300,N_5026,N_4842);
or U5301 (N_5301,N_5060,N_4946);
or U5302 (N_5302,N_4993,N_4875);
or U5303 (N_5303,N_5038,N_4864);
and U5304 (N_5304,N_4886,N_4828);
nand U5305 (N_5305,N_4838,N_4883);
and U5306 (N_5306,N_5045,N_4998);
or U5307 (N_5307,N_5010,N_4972);
nand U5308 (N_5308,N_5099,N_5055);
nand U5309 (N_5309,N_4940,N_4994);
nand U5310 (N_5310,N_4888,N_5006);
and U5311 (N_5311,N_4969,N_4952);
or U5312 (N_5312,N_4853,N_5017);
nor U5313 (N_5313,N_4929,N_5077);
nand U5314 (N_5314,N_4861,N_4808);
and U5315 (N_5315,N_5084,N_5057);
or U5316 (N_5316,N_4822,N_4932);
nand U5317 (N_5317,N_4889,N_4958);
nor U5318 (N_5318,N_4876,N_4880);
or U5319 (N_5319,N_4978,N_4915);
and U5320 (N_5320,N_4855,N_5020);
and U5321 (N_5321,N_4848,N_4964);
nor U5322 (N_5322,N_4960,N_5033);
and U5323 (N_5323,N_5043,N_5003);
nand U5324 (N_5324,N_4990,N_4987);
xnor U5325 (N_5325,N_4871,N_4885);
or U5326 (N_5326,N_5067,N_4811);
nor U5327 (N_5327,N_5081,N_5094);
and U5328 (N_5328,N_5048,N_5039);
nor U5329 (N_5329,N_4947,N_4827);
or U5330 (N_5330,N_5072,N_5018);
nor U5331 (N_5331,N_4885,N_4858);
nand U5332 (N_5332,N_4906,N_5087);
nor U5333 (N_5333,N_4908,N_5089);
or U5334 (N_5334,N_4996,N_4884);
xnor U5335 (N_5335,N_4999,N_4897);
and U5336 (N_5336,N_4842,N_4831);
or U5337 (N_5337,N_4849,N_5026);
and U5338 (N_5338,N_4826,N_4830);
nor U5339 (N_5339,N_5024,N_5036);
xor U5340 (N_5340,N_4921,N_5061);
nand U5341 (N_5341,N_4820,N_5054);
and U5342 (N_5342,N_4895,N_4961);
or U5343 (N_5343,N_4990,N_4881);
or U5344 (N_5344,N_5097,N_4985);
nor U5345 (N_5345,N_5062,N_4868);
nor U5346 (N_5346,N_4920,N_4897);
nor U5347 (N_5347,N_5073,N_5046);
nor U5348 (N_5348,N_5053,N_5092);
nor U5349 (N_5349,N_4803,N_5045);
xor U5350 (N_5350,N_5071,N_5051);
and U5351 (N_5351,N_4963,N_4972);
or U5352 (N_5352,N_4970,N_5087);
nor U5353 (N_5353,N_5085,N_4803);
nor U5354 (N_5354,N_5063,N_4845);
nor U5355 (N_5355,N_5083,N_5006);
or U5356 (N_5356,N_5078,N_4803);
nand U5357 (N_5357,N_5096,N_4854);
and U5358 (N_5358,N_5059,N_4957);
xnor U5359 (N_5359,N_5098,N_4806);
xnor U5360 (N_5360,N_4926,N_4884);
or U5361 (N_5361,N_5014,N_5034);
nor U5362 (N_5362,N_4826,N_4835);
and U5363 (N_5363,N_4869,N_4976);
xnor U5364 (N_5364,N_4886,N_4907);
xnor U5365 (N_5365,N_5007,N_5047);
or U5366 (N_5366,N_4943,N_4944);
xnor U5367 (N_5367,N_4859,N_5040);
xnor U5368 (N_5368,N_5084,N_4956);
or U5369 (N_5369,N_4824,N_4844);
nand U5370 (N_5370,N_5046,N_5047);
or U5371 (N_5371,N_4995,N_4861);
nand U5372 (N_5372,N_5002,N_4880);
nor U5373 (N_5373,N_5010,N_4938);
or U5374 (N_5374,N_5094,N_4898);
or U5375 (N_5375,N_4941,N_4814);
nor U5376 (N_5376,N_5010,N_5000);
nand U5377 (N_5377,N_5070,N_4956);
nor U5378 (N_5378,N_4898,N_5006);
and U5379 (N_5379,N_4916,N_4918);
or U5380 (N_5380,N_4842,N_4805);
or U5381 (N_5381,N_4986,N_5093);
and U5382 (N_5382,N_5085,N_4967);
or U5383 (N_5383,N_4818,N_4910);
or U5384 (N_5384,N_4887,N_4996);
or U5385 (N_5385,N_5021,N_4888);
nor U5386 (N_5386,N_5027,N_5047);
xnor U5387 (N_5387,N_4875,N_4994);
nor U5388 (N_5388,N_5059,N_5074);
nor U5389 (N_5389,N_4925,N_5019);
xnor U5390 (N_5390,N_5054,N_5088);
and U5391 (N_5391,N_4920,N_4831);
nand U5392 (N_5392,N_5065,N_4988);
nor U5393 (N_5393,N_4990,N_5066);
or U5394 (N_5394,N_4997,N_4998);
and U5395 (N_5395,N_5007,N_5094);
and U5396 (N_5396,N_5060,N_4934);
xor U5397 (N_5397,N_4983,N_5098);
nor U5398 (N_5398,N_5082,N_5068);
nor U5399 (N_5399,N_4946,N_4841);
or U5400 (N_5400,N_5103,N_5102);
nor U5401 (N_5401,N_5119,N_5105);
or U5402 (N_5402,N_5158,N_5265);
nor U5403 (N_5403,N_5214,N_5222);
or U5404 (N_5404,N_5246,N_5306);
xnor U5405 (N_5405,N_5388,N_5113);
xor U5406 (N_5406,N_5123,N_5327);
and U5407 (N_5407,N_5284,N_5258);
xnor U5408 (N_5408,N_5263,N_5337);
and U5409 (N_5409,N_5131,N_5330);
or U5410 (N_5410,N_5107,N_5278);
nand U5411 (N_5411,N_5377,N_5348);
or U5412 (N_5412,N_5269,N_5101);
nand U5413 (N_5413,N_5199,N_5262);
and U5414 (N_5414,N_5231,N_5351);
nand U5415 (N_5415,N_5106,N_5271);
and U5416 (N_5416,N_5386,N_5396);
nand U5417 (N_5417,N_5184,N_5310);
nand U5418 (N_5418,N_5373,N_5216);
nand U5419 (N_5419,N_5175,N_5364);
and U5420 (N_5420,N_5145,N_5155);
and U5421 (N_5421,N_5266,N_5339);
xnor U5422 (N_5422,N_5198,N_5352);
and U5423 (N_5423,N_5303,N_5305);
nor U5424 (N_5424,N_5148,N_5341);
nor U5425 (N_5425,N_5354,N_5210);
nand U5426 (N_5426,N_5363,N_5253);
nand U5427 (N_5427,N_5161,N_5191);
and U5428 (N_5428,N_5178,N_5116);
or U5429 (N_5429,N_5343,N_5204);
or U5430 (N_5430,N_5293,N_5152);
nor U5431 (N_5431,N_5108,N_5261);
and U5432 (N_5432,N_5164,N_5301);
xor U5433 (N_5433,N_5180,N_5366);
nand U5434 (N_5434,N_5112,N_5125);
nand U5435 (N_5435,N_5357,N_5296);
nand U5436 (N_5436,N_5273,N_5250);
xnor U5437 (N_5437,N_5147,N_5317);
nand U5438 (N_5438,N_5136,N_5240);
and U5439 (N_5439,N_5227,N_5398);
and U5440 (N_5440,N_5194,N_5212);
or U5441 (N_5441,N_5137,N_5270);
nor U5442 (N_5442,N_5228,N_5361);
or U5443 (N_5443,N_5344,N_5104);
and U5444 (N_5444,N_5213,N_5384);
nor U5445 (N_5445,N_5189,N_5200);
and U5446 (N_5446,N_5132,N_5259);
nand U5447 (N_5447,N_5291,N_5346);
and U5448 (N_5448,N_5391,N_5368);
and U5449 (N_5449,N_5252,N_5362);
nor U5450 (N_5450,N_5138,N_5181);
nand U5451 (N_5451,N_5129,N_5130);
or U5452 (N_5452,N_5335,N_5334);
xnor U5453 (N_5453,N_5294,N_5358);
nand U5454 (N_5454,N_5122,N_5295);
nand U5455 (N_5455,N_5172,N_5292);
and U5456 (N_5456,N_5353,N_5190);
nor U5457 (N_5457,N_5382,N_5326);
and U5458 (N_5458,N_5387,N_5196);
nand U5459 (N_5459,N_5340,N_5342);
nor U5460 (N_5460,N_5168,N_5128);
nor U5461 (N_5461,N_5383,N_5218);
nand U5462 (N_5462,N_5365,N_5345);
and U5463 (N_5463,N_5311,N_5225);
or U5464 (N_5464,N_5338,N_5211);
nand U5465 (N_5465,N_5224,N_5126);
nor U5466 (N_5466,N_5230,N_5399);
or U5467 (N_5467,N_5118,N_5234);
nor U5468 (N_5468,N_5195,N_5146);
nand U5469 (N_5469,N_5205,N_5376);
xor U5470 (N_5470,N_5217,N_5251);
xor U5471 (N_5471,N_5202,N_5397);
nand U5472 (N_5472,N_5187,N_5329);
nand U5473 (N_5473,N_5374,N_5332);
or U5474 (N_5474,N_5223,N_5283);
xor U5475 (N_5475,N_5257,N_5312);
or U5476 (N_5476,N_5307,N_5390);
or U5477 (N_5477,N_5157,N_5394);
xor U5478 (N_5478,N_5179,N_5149);
and U5479 (N_5479,N_5153,N_5115);
nand U5480 (N_5480,N_5208,N_5282);
or U5481 (N_5481,N_5281,N_5162);
or U5482 (N_5482,N_5197,N_5323);
xnor U5483 (N_5483,N_5276,N_5372);
nand U5484 (N_5484,N_5272,N_5275);
nor U5485 (N_5485,N_5209,N_5371);
or U5486 (N_5486,N_5241,N_5226);
xnor U5487 (N_5487,N_5308,N_5177);
xnor U5488 (N_5488,N_5267,N_5159);
or U5489 (N_5489,N_5170,N_5313);
or U5490 (N_5490,N_5300,N_5121);
or U5491 (N_5491,N_5206,N_5381);
nor U5492 (N_5492,N_5120,N_5183);
nor U5493 (N_5493,N_5264,N_5299);
nor U5494 (N_5494,N_5268,N_5165);
or U5495 (N_5495,N_5277,N_5304);
or U5496 (N_5496,N_5156,N_5385);
and U5497 (N_5497,N_5150,N_5221);
nand U5498 (N_5498,N_5135,N_5359);
nand U5499 (N_5499,N_5247,N_5349);
and U5500 (N_5500,N_5256,N_5314);
nor U5501 (N_5501,N_5239,N_5287);
nand U5502 (N_5502,N_5370,N_5243);
and U5503 (N_5503,N_5176,N_5143);
or U5504 (N_5504,N_5237,N_5144);
xor U5505 (N_5505,N_5254,N_5114);
nor U5506 (N_5506,N_5169,N_5193);
or U5507 (N_5507,N_5201,N_5203);
xor U5508 (N_5508,N_5229,N_5333);
xor U5509 (N_5509,N_5356,N_5297);
nor U5510 (N_5510,N_5100,N_5290);
xor U5511 (N_5511,N_5235,N_5173);
nor U5512 (N_5512,N_5302,N_5380);
xor U5513 (N_5513,N_5124,N_5244);
nor U5514 (N_5514,N_5166,N_5260);
xor U5515 (N_5515,N_5133,N_5255);
and U5516 (N_5516,N_5319,N_5318);
or U5517 (N_5517,N_5274,N_5298);
or U5518 (N_5518,N_5315,N_5378);
and U5519 (N_5519,N_5288,N_5154);
nand U5520 (N_5520,N_5233,N_5188);
nand U5521 (N_5521,N_5309,N_5395);
nor U5522 (N_5522,N_5220,N_5171);
xnor U5523 (N_5523,N_5232,N_5110);
nand U5524 (N_5524,N_5393,N_5127);
and U5525 (N_5525,N_5360,N_5167);
nor U5526 (N_5526,N_5139,N_5207);
xnor U5527 (N_5527,N_5289,N_5236);
xor U5528 (N_5528,N_5392,N_5248);
and U5529 (N_5529,N_5321,N_5367);
xor U5530 (N_5530,N_5185,N_5219);
nor U5531 (N_5531,N_5331,N_5186);
xor U5532 (N_5532,N_5322,N_5324);
or U5533 (N_5533,N_5141,N_5336);
nand U5534 (N_5534,N_5245,N_5182);
nand U5535 (N_5535,N_5347,N_5369);
and U5536 (N_5536,N_5350,N_5238);
xnor U5537 (N_5537,N_5174,N_5215);
xor U5538 (N_5538,N_5109,N_5242);
or U5539 (N_5539,N_5285,N_5325);
xor U5540 (N_5540,N_5280,N_5140);
nor U5541 (N_5541,N_5379,N_5249);
nor U5542 (N_5542,N_5160,N_5375);
xnor U5543 (N_5543,N_5111,N_5117);
nand U5544 (N_5544,N_5286,N_5389);
and U5545 (N_5545,N_5316,N_5320);
and U5546 (N_5546,N_5328,N_5151);
nand U5547 (N_5547,N_5142,N_5192);
nor U5548 (N_5548,N_5279,N_5163);
or U5549 (N_5549,N_5134,N_5355);
nor U5550 (N_5550,N_5114,N_5228);
nand U5551 (N_5551,N_5254,N_5295);
or U5552 (N_5552,N_5117,N_5184);
nor U5553 (N_5553,N_5174,N_5354);
xnor U5554 (N_5554,N_5103,N_5281);
or U5555 (N_5555,N_5149,N_5246);
and U5556 (N_5556,N_5383,N_5324);
nor U5557 (N_5557,N_5172,N_5345);
nand U5558 (N_5558,N_5391,N_5218);
and U5559 (N_5559,N_5243,N_5141);
nor U5560 (N_5560,N_5221,N_5229);
and U5561 (N_5561,N_5311,N_5367);
xor U5562 (N_5562,N_5123,N_5294);
nand U5563 (N_5563,N_5308,N_5370);
or U5564 (N_5564,N_5393,N_5263);
or U5565 (N_5565,N_5116,N_5282);
nor U5566 (N_5566,N_5231,N_5381);
and U5567 (N_5567,N_5208,N_5111);
nor U5568 (N_5568,N_5360,N_5279);
xnor U5569 (N_5569,N_5370,N_5221);
nand U5570 (N_5570,N_5394,N_5308);
nand U5571 (N_5571,N_5308,N_5269);
nand U5572 (N_5572,N_5154,N_5171);
nor U5573 (N_5573,N_5161,N_5224);
or U5574 (N_5574,N_5231,N_5207);
nor U5575 (N_5575,N_5100,N_5161);
nand U5576 (N_5576,N_5308,N_5315);
or U5577 (N_5577,N_5254,N_5116);
xor U5578 (N_5578,N_5344,N_5371);
nand U5579 (N_5579,N_5175,N_5120);
and U5580 (N_5580,N_5213,N_5252);
nor U5581 (N_5581,N_5204,N_5163);
nor U5582 (N_5582,N_5158,N_5367);
nor U5583 (N_5583,N_5362,N_5391);
xnor U5584 (N_5584,N_5167,N_5201);
xnor U5585 (N_5585,N_5366,N_5168);
nor U5586 (N_5586,N_5275,N_5266);
and U5587 (N_5587,N_5154,N_5313);
xor U5588 (N_5588,N_5119,N_5258);
nor U5589 (N_5589,N_5191,N_5324);
nor U5590 (N_5590,N_5367,N_5308);
and U5591 (N_5591,N_5208,N_5299);
and U5592 (N_5592,N_5385,N_5315);
or U5593 (N_5593,N_5388,N_5212);
nand U5594 (N_5594,N_5340,N_5104);
and U5595 (N_5595,N_5307,N_5147);
nor U5596 (N_5596,N_5131,N_5382);
and U5597 (N_5597,N_5399,N_5372);
nor U5598 (N_5598,N_5177,N_5389);
or U5599 (N_5599,N_5198,N_5222);
nor U5600 (N_5600,N_5209,N_5173);
nand U5601 (N_5601,N_5346,N_5189);
nand U5602 (N_5602,N_5256,N_5346);
nor U5603 (N_5603,N_5273,N_5368);
nand U5604 (N_5604,N_5373,N_5195);
xnor U5605 (N_5605,N_5175,N_5114);
xor U5606 (N_5606,N_5394,N_5377);
xnor U5607 (N_5607,N_5277,N_5241);
and U5608 (N_5608,N_5302,N_5140);
xnor U5609 (N_5609,N_5239,N_5241);
nor U5610 (N_5610,N_5274,N_5364);
nand U5611 (N_5611,N_5323,N_5327);
and U5612 (N_5612,N_5364,N_5231);
nor U5613 (N_5613,N_5206,N_5289);
or U5614 (N_5614,N_5217,N_5283);
nand U5615 (N_5615,N_5357,N_5160);
and U5616 (N_5616,N_5330,N_5267);
nor U5617 (N_5617,N_5314,N_5174);
or U5618 (N_5618,N_5315,N_5307);
or U5619 (N_5619,N_5139,N_5254);
nor U5620 (N_5620,N_5315,N_5341);
nor U5621 (N_5621,N_5325,N_5116);
nand U5622 (N_5622,N_5163,N_5331);
nand U5623 (N_5623,N_5114,N_5205);
and U5624 (N_5624,N_5195,N_5150);
xor U5625 (N_5625,N_5221,N_5216);
nand U5626 (N_5626,N_5395,N_5388);
nand U5627 (N_5627,N_5237,N_5319);
nand U5628 (N_5628,N_5123,N_5255);
nor U5629 (N_5629,N_5370,N_5232);
and U5630 (N_5630,N_5359,N_5292);
xnor U5631 (N_5631,N_5360,N_5286);
nand U5632 (N_5632,N_5352,N_5371);
or U5633 (N_5633,N_5262,N_5360);
or U5634 (N_5634,N_5174,N_5344);
and U5635 (N_5635,N_5208,N_5281);
nand U5636 (N_5636,N_5286,N_5156);
and U5637 (N_5637,N_5131,N_5264);
nor U5638 (N_5638,N_5127,N_5380);
nand U5639 (N_5639,N_5250,N_5198);
or U5640 (N_5640,N_5152,N_5221);
and U5641 (N_5641,N_5332,N_5161);
nor U5642 (N_5642,N_5197,N_5108);
or U5643 (N_5643,N_5183,N_5235);
nor U5644 (N_5644,N_5325,N_5328);
nor U5645 (N_5645,N_5392,N_5217);
and U5646 (N_5646,N_5210,N_5242);
nor U5647 (N_5647,N_5392,N_5243);
and U5648 (N_5648,N_5199,N_5180);
nor U5649 (N_5649,N_5260,N_5230);
xnor U5650 (N_5650,N_5166,N_5333);
nand U5651 (N_5651,N_5234,N_5179);
or U5652 (N_5652,N_5354,N_5318);
or U5653 (N_5653,N_5354,N_5238);
or U5654 (N_5654,N_5123,N_5168);
and U5655 (N_5655,N_5210,N_5262);
and U5656 (N_5656,N_5186,N_5330);
and U5657 (N_5657,N_5369,N_5261);
nor U5658 (N_5658,N_5332,N_5111);
nand U5659 (N_5659,N_5386,N_5129);
or U5660 (N_5660,N_5128,N_5214);
nand U5661 (N_5661,N_5137,N_5382);
nand U5662 (N_5662,N_5126,N_5337);
or U5663 (N_5663,N_5160,N_5198);
and U5664 (N_5664,N_5380,N_5258);
nand U5665 (N_5665,N_5119,N_5154);
nor U5666 (N_5666,N_5102,N_5310);
nand U5667 (N_5667,N_5396,N_5174);
nor U5668 (N_5668,N_5301,N_5231);
nor U5669 (N_5669,N_5268,N_5199);
and U5670 (N_5670,N_5333,N_5126);
nand U5671 (N_5671,N_5228,N_5168);
nor U5672 (N_5672,N_5152,N_5163);
xnor U5673 (N_5673,N_5152,N_5389);
and U5674 (N_5674,N_5118,N_5182);
or U5675 (N_5675,N_5351,N_5244);
nand U5676 (N_5676,N_5309,N_5225);
or U5677 (N_5677,N_5149,N_5209);
xor U5678 (N_5678,N_5196,N_5242);
xor U5679 (N_5679,N_5346,N_5216);
nand U5680 (N_5680,N_5164,N_5290);
nor U5681 (N_5681,N_5356,N_5386);
nand U5682 (N_5682,N_5239,N_5171);
and U5683 (N_5683,N_5391,N_5238);
nand U5684 (N_5684,N_5352,N_5353);
xor U5685 (N_5685,N_5115,N_5181);
nor U5686 (N_5686,N_5245,N_5311);
and U5687 (N_5687,N_5293,N_5200);
nor U5688 (N_5688,N_5322,N_5160);
or U5689 (N_5689,N_5233,N_5179);
or U5690 (N_5690,N_5244,N_5163);
nand U5691 (N_5691,N_5234,N_5373);
nor U5692 (N_5692,N_5116,N_5377);
and U5693 (N_5693,N_5118,N_5326);
nor U5694 (N_5694,N_5261,N_5237);
nand U5695 (N_5695,N_5167,N_5292);
nor U5696 (N_5696,N_5205,N_5239);
or U5697 (N_5697,N_5119,N_5178);
nand U5698 (N_5698,N_5324,N_5163);
nor U5699 (N_5699,N_5299,N_5125);
or U5700 (N_5700,N_5410,N_5405);
nand U5701 (N_5701,N_5422,N_5430);
or U5702 (N_5702,N_5468,N_5624);
xor U5703 (N_5703,N_5485,N_5686);
or U5704 (N_5704,N_5527,N_5577);
or U5705 (N_5705,N_5623,N_5497);
and U5706 (N_5706,N_5655,N_5532);
and U5707 (N_5707,N_5506,N_5505);
xor U5708 (N_5708,N_5564,N_5523);
or U5709 (N_5709,N_5669,N_5674);
nor U5710 (N_5710,N_5607,N_5442);
xnor U5711 (N_5711,N_5647,N_5608);
nand U5712 (N_5712,N_5519,N_5446);
or U5713 (N_5713,N_5551,N_5401);
and U5714 (N_5714,N_5511,N_5616);
and U5715 (N_5715,N_5627,N_5416);
nand U5716 (N_5716,N_5621,N_5681);
nor U5717 (N_5717,N_5515,N_5633);
or U5718 (N_5718,N_5455,N_5646);
xnor U5719 (N_5719,N_5672,N_5571);
and U5720 (N_5720,N_5593,N_5481);
and U5721 (N_5721,N_5406,N_5563);
nand U5722 (N_5722,N_5685,N_5544);
xnor U5723 (N_5723,N_5676,N_5413);
nor U5724 (N_5724,N_5661,N_5484);
xnor U5725 (N_5725,N_5635,N_5565);
nand U5726 (N_5726,N_5463,N_5494);
nand U5727 (N_5727,N_5696,N_5656);
or U5728 (N_5728,N_5659,N_5456);
and U5729 (N_5729,N_5566,N_5574);
xnor U5730 (N_5730,N_5412,N_5586);
xnor U5731 (N_5731,N_5678,N_5622);
nor U5732 (N_5732,N_5640,N_5517);
nor U5733 (N_5733,N_5503,N_5490);
and U5734 (N_5734,N_5618,N_5437);
and U5735 (N_5735,N_5535,N_5510);
nand U5736 (N_5736,N_5499,N_5459);
xor U5737 (N_5737,N_5454,N_5534);
nand U5738 (N_5738,N_5617,N_5429);
xor U5739 (N_5739,N_5435,N_5426);
or U5740 (N_5740,N_5525,N_5407);
and U5741 (N_5741,N_5480,N_5495);
and U5742 (N_5742,N_5698,N_5414);
nor U5743 (N_5743,N_5561,N_5651);
xor U5744 (N_5744,N_5440,N_5599);
and U5745 (N_5745,N_5626,N_5460);
nor U5746 (N_5746,N_5541,N_5464);
and U5747 (N_5747,N_5552,N_5689);
nor U5748 (N_5748,N_5664,N_5634);
or U5749 (N_5749,N_5555,N_5628);
xnor U5750 (N_5750,N_5516,N_5501);
or U5751 (N_5751,N_5478,N_5691);
nand U5752 (N_5752,N_5467,N_5508);
xnor U5753 (N_5753,N_5677,N_5504);
xnor U5754 (N_5754,N_5680,N_5600);
nor U5755 (N_5755,N_5648,N_5584);
xnor U5756 (N_5756,N_5500,N_5598);
nand U5757 (N_5757,N_5668,N_5663);
nand U5758 (N_5758,N_5424,N_5575);
xor U5759 (N_5759,N_5556,N_5675);
and U5760 (N_5760,N_5447,N_5486);
nand U5761 (N_5761,N_5404,N_5502);
xnor U5762 (N_5762,N_5548,N_5694);
or U5763 (N_5763,N_5639,N_5521);
nand U5764 (N_5764,N_5580,N_5493);
nand U5765 (N_5765,N_5550,N_5400);
xnor U5766 (N_5766,N_5590,N_5539);
or U5767 (N_5767,N_5529,N_5449);
nand U5768 (N_5768,N_5409,N_5625);
and U5769 (N_5769,N_5475,N_5636);
nor U5770 (N_5770,N_5549,N_5473);
and U5771 (N_5771,N_5643,N_5433);
nand U5772 (N_5772,N_5432,N_5649);
and U5773 (N_5773,N_5419,N_5583);
xor U5774 (N_5774,N_5644,N_5434);
nor U5775 (N_5775,N_5684,N_5582);
nand U5776 (N_5776,N_5595,N_5425);
or U5777 (N_5777,N_5488,N_5579);
or U5778 (N_5778,N_5472,N_5458);
nor U5779 (N_5779,N_5572,N_5526);
xnor U5780 (N_5780,N_5568,N_5557);
nand U5781 (N_5781,N_5692,N_5452);
xor U5782 (N_5782,N_5610,N_5697);
xnor U5783 (N_5783,N_5606,N_5487);
nand U5784 (N_5784,N_5642,N_5597);
nand U5785 (N_5785,N_5469,N_5638);
and U5786 (N_5786,N_5542,N_5604);
nor U5787 (N_5787,N_5524,N_5522);
and U5788 (N_5788,N_5512,N_5547);
xnor U5789 (N_5789,N_5443,N_5531);
and U5790 (N_5790,N_5543,N_5602);
nor U5791 (N_5791,N_5431,N_5613);
or U5792 (N_5792,N_5630,N_5546);
and U5793 (N_5793,N_5496,N_5665);
nand U5794 (N_5794,N_5587,N_5662);
and U5795 (N_5795,N_5650,N_5417);
nand U5796 (N_5796,N_5415,N_5423);
nand U5797 (N_5797,N_5679,N_5601);
nand U5798 (N_5798,N_5445,N_5660);
nor U5799 (N_5799,N_5457,N_5513);
or U5800 (N_5800,N_5554,N_5611);
nor U5801 (N_5801,N_5652,N_5418);
or U5802 (N_5802,N_5609,N_5666);
nor U5803 (N_5803,N_5687,N_5581);
nor U5804 (N_5804,N_5466,N_5538);
and U5805 (N_5805,N_5537,N_5629);
nand U5806 (N_5806,N_5567,N_5540);
nor U5807 (N_5807,N_5612,N_5578);
and U5808 (N_5808,N_5667,N_5569);
or U5809 (N_5809,N_5637,N_5470);
and U5810 (N_5810,N_5570,N_5444);
nor U5811 (N_5811,N_5465,N_5619);
and U5812 (N_5812,N_5530,N_5682);
and U5813 (N_5813,N_5411,N_5670);
nand U5814 (N_5814,N_5479,N_5483);
nor U5815 (N_5815,N_5588,N_5509);
and U5816 (N_5816,N_5427,N_5631);
nor U5817 (N_5817,N_5438,N_5491);
xor U5818 (N_5818,N_5690,N_5498);
xor U5819 (N_5819,N_5695,N_5441);
nor U5820 (N_5820,N_5592,N_5573);
and U5821 (N_5821,N_5576,N_5461);
nand U5822 (N_5822,N_5699,N_5632);
nand U5823 (N_5823,N_5589,N_5673);
nor U5824 (N_5824,N_5536,N_5520);
or U5825 (N_5825,N_5428,N_5671);
or U5826 (N_5826,N_5474,N_5507);
nor U5827 (N_5827,N_5558,N_5492);
nor U5828 (N_5828,N_5591,N_5645);
or U5829 (N_5829,N_5653,N_5658);
nand U5830 (N_5830,N_5453,N_5436);
xnor U5831 (N_5831,N_5562,N_5482);
xor U5832 (N_5832,N_5641,N_5514);
and U5833 (N_5833,N_5471,N_5605);
nand U5834 (N_5834,N_5657,N_5585);
nand U5835 (N_5835,N_5439,N_5545);
or U5836 (N_5836,N_5594,N_5693);
and U5837 (N_5837,N_5553,N_5559);
and U5838 (N_5838,N_5489,N_5654);
and U5839 (N_5839,N_5450,N_5615);
nand U5840 (N_5840,N_5528,N_5560);
xor U5841 (N_5841,N_5683,N_5688);
and U5842 (N_5842,N_5476,N_5462);
nand U5843 (N_5843,N_5408,N_5596);
nand U5844 (N_5844,N_5451,N_5420);
or U5845 (N_5845,N_5533,N_5603);
nand U5846 (N_5846,N_5421,N_5620);
nor U5847 (N_5847,N_5448,N_5518);
nand U5848 (N_5848,N_5477,N_5402);
or U5849 (N_5849,N_5614,N_5403);
xnor U5850 (N_5850,N_5403,N_5423);
nor U5851 (N_5851,N_5413,N_5412);
xnor U5852 (N_5852,N_5460,N_5483);
or U5853 (N_5853,N_5611,N_5476);
and U5854 (N_5854,N_5508,N_5577);
and U5855 (N_5855,N_5654,N_5487);
nand U5856 (N_5856,N_5597,N_5625);
nand U5857 (N_5857,N_5428,N_5406);
or U5858 (N_5858,N_5604,N_5669);
and U5859 (N_5859,N_5583,N_5480);
nor U5860 (N_5860,N_5474,N_5555);
nand U5861 (N_5861,N_5405,N_5661);
xor U5862 (N_5862,N_5544,N_5450);
or U5863 (N_5863,N_5411,N_5485);
nor U5864 (N_5864,N_5639,N_5426);
or U5865 (N_5865,N_5546,N_5559);
xor U5866 (N_5866,N_5695,N_5474);
or U5867 (N_5867,N_5638,N_5501);
or U5868 (N_5868,N_5473,N_5665);
nor U5869 (N_5869,N_5539,N_5421);
or U5870 (N_5870,N_5587,N_5448);
nor U5871 (N_5871,N_5486,N_5571);
nor U5872 (N_5872,N_5490,N_5401);
nand U5873 (N_5873,N_5540,N_5661);
nor U5874 (N_5874,N_5584,N_5668);
or U5875 (N_5875,N_5512,N_5523);
or U5876 (N_5876,N_5521,N_5579);
xnor U5877 (N_5877,N_5476,N_5675);
and U5878 (N_5878,N_5509,N_5685);
nand U5879 (N_5879,N_5599,N_5557);
nor U5880 (N_5880,N_5538,N_5436);
nor U5881 (N_5881,N_5479,N_5539);
nand U5882 (N_5882,N_5684,N_5598);
and U5883 (N_5883,N_5552,N_5594);
and U5884 (N_5884,N_5471,N_5519);
xor U5885 (N_5885,N_5424,N_5688);
xnor U5886 (N_5886,N_5551,N_5601);
xor U5887 (N_5887,N_5431,N_5589);
and U5888 (N_5888,N_5418,N_5426);
nor U5889 (N_5889,N_5462,N_5513);
xor U5890 (N_5890,N_5459,N_5576);
xnor U5891 (N_5891,N_5427,N_5693);
nor U5892 (N_5892,N_5623,N_5697);
or U5893 (N_5893,N_5609,N_5691);
nand U5894 (N_5894,N_5564,N_5479);
nand U5895 (N_5895,N_5400,N_5588);
or U5896 (N_5896,N_5670,N_5525);
xnor U5897 (N_5897,N_5525,N_5579);
or U5898 (N_5898,N_5688,N_5685);
and U5899 (N_5899,N_5546,N_5594);
nand U5900 (N_5900,N_5620,N_5636);
and U5901 (N_5901,N_5555,N_5697);
and U5902 (N_5902,N_5406,N_5522);
and U5903 (N_5903,N_5578,N_5601);
xor U5904 (N_5904,N_5632,N_5698);
nand U5905 (N_5905,N_5546,N_5576);
and U5906 (N_5906,N_5696,N_5655);
nor U5907 (N_5907,N_5659,N_5553);
nand U5908 (N_5908,N_5455,N_5426);
xor U5909 (N_5909,N_5514,N_5419);
nor U5910 (N_5910,N_5548,N_5606);
nand U5911 (N_5911,N_5617,N_5667);
nor U5912 (N_5912,N_5510,N_5461);
nor U5913 (N_5913,N_5682,N_5447);
xor U5914 (N_5914,N_5435,N_5522);
xnor U5915 (N_5915,N_5431,N_5420);
and U5916 (N_5916,N_5666,N_5635);
xnor U5917 (N_5917,N_5465,N_5512);
or U5918 (N_5918,N_5519,N_5452);
nand U5919 (N_5919,N_5626,N_5561);
and U5920 (N_5920,N_5436,N_5430);
or U5921 (N_5921,N_5410,N_5637);
or U5922 (N_5922,N_5506,N_5655);
nor U5923 (N_5923,N_5649,N_5528);
and U5924 (N_5924,N_5465,N_5679);
nand U5925 (N_5925,N_5428,N_5404);
or U5926 (N_5926,N_5699,N_5643);
nor U5927 (N_5927,N_5595,N_5466);
xnor U5928 (N_5928,N_5605,N_5449);
and U5929 (N_5929,N_5623,N_5500);
nand U5930 (N_5930,N_5529,N_5508);
xor U5931 (N_5931,N_5539,N_5696);
xnor U5932 (N_5932,N_5545,N_5498);
nor U5933 (N_5933,N_5499,N_5678);
nand U5934 (N_5934,N_5523,N_5577);
or U5935 (N_5935,N_5578,N_5490);
nor U5936 (N_5936,N_5473,N_5529);
xnor U5937 (N_5937,N_5416,N_5545);
or U5938 (N_5938,N_5588,N_5650);
and U5939 (N_5939,N_5474,N_5536);
and U5940 (N_5940,N_5517,N_5510);
and U5941 (N_5941,N_5495,N_5659);
nor U5942 (N_5942,N_5428,N_5418);
nor U5943 (N_5943,N_5674,N_5466);
or U5944 (N_5944,N_5689,N_5599);
nor U5945 (N_5945,N_5424,N_5613);
nand U5946 (N_5946,N_5482,N_5536);
nand U5947 (N_5947,N_5693,N_5407);
nor U5948 (N_5948,N_5660,N_5413);
or U5949 (N_5949,N_5431,N_5558);
nand U5950 (N_5950,N_5697,N_5542);
and U5951 (N_5951,N_5444,N_5646);
xor U5952 (N_5952,N_5495,N_5400);
or U5953 (N_5953,N_5545,N_5450);
and U5954 (N_5954,N_5601,N_5631);
or U5955 (N_5955,N_5522,N_5514);
nand U5956 (N_5956,N_5666,N_5651);
or U5957 (N_5957,N_5523,N_5529);
or U5958 (N_5958,N_5691,N_5545);
nand U5959 (N_5959,N_5588,N_5487);
xnor U5960 (N_5960,N_5633,N_5454);
and U5961 (N_5961,N_5457,N_5585);
nand U5962 (N_5962,N_5500,N_5618);
nor U5963 (N_5963,N_5555,N_5463);
or U5964 (N_5964,N_5403,N_5484);
xor U5965 (N_5965,N_5493,N_5522);
nand U5966 (N_5966,N_5584,N_5441);
nand U5967 (N_5967,N_5533,N_5562);
nand U5968 (N_5968,N_5446,N_5421);
xor U5969 (N_5969,N_5414,N_5574);
nor U5970 (N_5970,N_5508,N_5569);
and U5971 (N_5971,N_5482,N_5644);
nand U5972 (N_5972,N_5431,N_5495);
and U5973 (N_5973,N_5449,N_5665);
nor U5974 (N_5974,N_5533,N_5430);
xnor U5975 (N_5975,N_5670,N_5553);
nor U5976 (N_5976,N_5493,N_5471);
nor U5977 (N_5977,N_5595,N_5558);
xor U5978 (N_5978,N_5603,N_5434);
nor U5979 (N_5979,N_5527,N_5675);
xnor U5980 (N_5980,N_5504,N_5641);
or U5981 (N_5981,N_5425,N_5612);
nand U5982 (N_5982,N_5519,N_5630);
nand U5983 (N_5983,N_5568,N_5513);
nand U5984 (N_5984,N_5486,N_5539);
nand U5985 (N_5985,N_5620,N_5469);
or U5986 (N_5986,N_5532,N_5459);
or U5987 (N_5987,N_5535,N_5561);
and U5988 (N_5988,N_5522,N_5598);
nor U5989 (N_5989,N_5651,N_5436);
nand U5990 (N_5990,N_5480,N_5599);
or U5991 (N_5991,N_5506,N_5448);
or U5992 (N_5992,N_5568,N_5426);
xnor U5993 (N_5993,N_5645,N_5601);
nor U5994 (N_5994,N_5577,N_5504);
xor U5995 (N_5995,N_5459,N_5614);
or U5996 (N_5996,N_5566,N_5653);
and U5997 (N_5997,N_5554,N_5560);
or U5998 (N_5998,N_5569,N_5500);
and U5999 (N_5999,N_5471,N_5488);
and U6000 (N_6000,N_5947,N_5816);
and U6001 (N_6001,N_5932,N_5759);
or U6002 (N_6002,N_5858,N_5910);
nor U6003 (N_6003,N_5953,N_5722);
nor U6004 (N_6004,N_5749,N_5831);
nand U6005 (N_6005,N_5824,N_5745);
xnor U6006 (N_6006,N_5769,N_5944);
or U6007 (N_6007,N_5950,N_5987);
and U6008 (N_6008,N_5941,N_5841);
xnor U6009 (N_6009,N_5978,N_5893);
and U6010 (N_6010,N_5871,N_5717);
xor U6011 (N_6011,N_5888,N_5994);
and U6012 (N_6012,N_5988,N_5891);
nand U6013 (N_6013,N_5815,N_5892);
and U6014 (N_6014,N_5995,N_5836);
and U6015 (N_6015,N_5737,N_5964);
xnor U6016 (N_6016,N_5889,N_5743);
xor U6017 (N_6017,N_5733,N_5999);
or U6018 (N_6018,N_5726,N_5900);
nor U6019 (N_6019,N_5912,N_5904);
and U6020 (N_6020,N_5913,N_5935);
or U6021 (N_6021,N_5742,N_5794);
xor U6022 (N_6022,N_5847,N_5886);
or U6023 (N_6023,N_5774,N_5908);
xor U6024 (N_6024,N_5830,N_5919);
nor U6025 (N_6025,N_5977,N_5755);
nor U6026 (N_6026,N_5704,N_5760);
nor U6027 (N_6027,N_5712,N_5776);
and U6028 (N_6028,N_5739,N_5738);
xor U6029 (N_6029,N_5865,N_5821);
and U6030 (N_6030,N_5915,N_5960);
or U6031 (N_6031,N_5967,N_5877);
nor U6032 (N_6032,N_5906,N_5780);
and U6033 (N_6033,N_5867,N_5850);
xor U6034 (N_6034,N_5724,N_5720);
nand U6035 (N_6035,N_5806,N_5853);
or U6036 (N_6036,N_5903,N_5949);
nor U6037 (N_6037,N_5800,N_5946);
xnor U6038 (N_6038,N_5939,N_5719);
nor U6039 (N_6039,N_5775,N_5822);
or U6040 (N_6040,N_5835,N_5894);
and U6041 (N_6041,N_5721,N_5789);
nand U6042 (N_6042,N_5880,N_5917);
xnor U6043 (N_6043,N_5864,N_5765);
xor U6044 (N_6044,N_5884,N_5703);
and U6045 (N_6045,N_5741,N_5996);
xnor U6046 (N_6046,N_5753,N_5873);
or U6047 (N_6047,N_5730,N_5861);
nand U6048 (N_6048,N_5907,N_5971);
and U6049 (N_6049,N_5786,N_5767);
and U6050 (N_6050,N_5825,N_5808);
or U6051 (N_6051,N_5832,N_5940);
and U6052 (N_6052,N_5772,N_5827);
and U6053 (N_6053,N_5833,N_5708);
nand U6054 (N_6054,N_5933,N_5883);
or U6055 (N_6055,N_5968,N_5844);
or U6056 (N_6056,N_5998,N_5709);
and U6057 (N_6057,N_5705,N_5823);
nor U6058 (N_6058,N_5779,N_5793);
nand U6059 (N_6059,N_5807,N_5909);
or U6060 (N_6060,N_5798,N_5862);
nor U6061 (N_6061,N_5879,N_5711);
nor U6062 (N_6062,N_5736,N_5973);
or U6063 (N_6063,N_5819,N_5734);
nand U6064 (N_6064,N_5896,N_5937);
xnor U6065 (N_6065,N_5875,N_5934);
nand U6066 (N_6066,N_5963,N_5868);
or U6067 (N_6067,N_5961,N_5898);
nor U6068 (N_6068,N_5989,N_5969);
nor U6069 (N_6069,N_5936,N_5802);
nor U6070 (N_6070,N_5837,N_5810);
or U6071 (N_6071,N_5731,N_5895);
xnor U6072 (N_6072,N_5990,N_5899);
and U6073 (N_6073,N_5809,N_5838);
and U6074 (N_6074,N_5992,N_5956);
nand U6075 (N_6075,N_5812,N_5966);
xor U6076 (N_6076,N_5938,N_5795);
nor U6077 (N_6077,N_5984,N_5855);
or U6078 (N_6078,N_5757,N_5834);
and U6079 (N_6079,N_5714,N_5878);
nand U6080 (N_6080,N_5788,N_5754);
xnor U6081 (N_6081,N_5848,N_5783);
xnor U6082 (N_6082,N_5785,N_5986);
or U6083 (N_6083,N_5744,N_5974);
and U6084 (N_6084,N_5991,N_5732);
and U6085 (N_6085,N_5751,N_5980);
or U6086 (N_6086,N_5700,N_5931);
xnor U6087 (N_6087,N_5778,N_5747);
or U6088 (N_6088,N_5828,N_5911);
or U6089 (N_6089,N_5857,N_5920);
nor U6090 (N_6090,N_5791,N_5870);
and U6091 (N_6091,N_5887,N_5852);
nand U6092 (N_6092,N_5860,N_5885);
and U6093 (N_6093,N_5985,N_5943);
and U6094 (N_6094,N_5829,N_5972);
xor U6095 (N_6095,N_5797,N_5901);
xor U6096 (N_6096,N_5840,N_5763);
and U6097 (N_6097,N_5856,N_5817);
and U6098 (N_6098,N_5805,N_5761);
nand U6099 (N_6099,N_5997,N_5784);
nor U6100 (N_6100,N_5758,N_5770);
xnor U6101 (N_6101,N_5928,N_5727);
or U6102 (N_6102,N_5849,N_5923);
nor U6103 (N_6103,N_5787,N_5890);
xnor U6104 (N_6104,N_5914,N_5916);
nor U6105 (N_6105,N_5970,N_5811);
or U6106 (N_6106,N_5866,N_5948);
nand U6107 (N_6107,N_5799,N_5728);
or U6108 (N_6108,N_5843,N_5740);
nand U6109 (N_6109,N_5748,N_5975);
or U6110 (N_6110,N_5801,N_5976);
and U6111 (N_6111,N_5902,N_5777);
or U6112 (N_6112,N_5876,N_5762);
xor U6113 (N_6113,N_5842,N_5905);
or U6114 (N_6114,N_5897,N_5735);
nand U6115 (N_6115,N_5818,N_5983);
and U6116 (N_6116,N_5803,N_5945);
or U6117 (N_6117,N_5782,N_5796);
or U6118 (N_6118,N_5882,N_5746);
or U6119 (N_6119,N_5716,N_5925);
and U6120 (N_6120,N_5965,N_5962);
or U6121 (N_6121,N_5713,N_5826);
nand U6122 (N_6122,N_5959,N_5957);
or U6123 (N_6123,N_5872,N_5942);
or U6124 (N_6124,N_5874,N_5924);
nor U6125 (N_6125,N_5955,N_5710);
and U6126 (N_6126,N_5839,N_5952);
or U6127 (N_6127,N_5814,N_5951);
nand U6128 (N_6128,N_5725,N_5851);
nor U6129 (N_6129,N_5706,N_5718);
nor U6130 (N_6130,N_5922,N_5771);
nor U6131 (N_6131,N_5881,N_5790);
and U6132 (N_6132,N_5927,N_5854);
xnor U6133 (N_6133,N_5804,N_5979);
nor U6134 (N_6134,N_5859,N_5921);
nor U6135 (N_6135,N_5756,N_5813);
xnor U6136 (N_6136,N_5766,N_5845);
xor U6137 (N_6137,N_5701,N_5869);
and U6138 (N_6138,N_5773,N_5954);
xnor U6139 (N_6139,N_5715,N_5930);
and U6140 (N_6140,N_5729,N_5918);
xnor U6141 (N_6141,N_5982,N_5993);
or U6142 (N_6142,N_5846,N_5820);
and U6143 (N_6143,N_5929,N_5764);
or U6144 (N_6144,N_5863,N_5981);
nor U6145 (N_6145,N_5958,N_5723);
nor U6146 (N_6146,N_5707,N_5926);
nand U6147 (N_6147,N_5752,N_5781);
nand U6148 (N_6148,N_5750,N_5702);
nand U6149 (N_6149,N_5792,N_5768);
xor U6150 (N_6150,N_5886,N_5829);
or U6151 (N_6151,N_5730,N_5834);
xnor U6152 (N_6152,N_5722,N_5834);
or U6153 (N_6153,N_5948,N_5747);
or U6154 (N_6154,N_5834,N_5839);
or U6155 (N_6155,N_5761,N_5999);
nand U6156 (N_6156,N_5977,N_5716);
and U6157 (N_6157,N_5948,N_5933);
and U6158 (N_6158,N_5832,N_5925);
nand U6159 (N_6159,N_5995,N_5867);
nand U6160 (N_6160,N_5873,N_5805);
xnor U6161 (N_6161,N_5928,N_5993);
or U6162 (N_6162,N_5843,N_5808);
and U6163 (N_6163,N_5989,N_5850);
nand U6164 (N_6164,N_5731,N_5763);
or U6165 (N_6165,N_5833,N_5752);
nand U6166 (N_6166,N_5965,N_5836);
and U6167 (N_6167,N_5982,N_5750);
nand U6168 (N_6168,N_5966,N_5732);
nor U6169 (N_6169,N_5879,N_5906);
xor U6170 (N_6170,N_5983,N_5900);
nand U6171 (N_6171,N_5889,N_5985);
xnor U6172 (N_6172,N_5710,N_5724);
xor U6173 (N_6173,N_5809,N_5954);
or U6174 (N_6174,N_5936,N_5990);
nand U6175 (N_6175,N_5936,N_5773);
or U6176 (N_6176,N_5961,N_5822);
nor U6177 (N_6177,N_5743,N_5838);
or U6178 (N_6178,N_5976,N_5710);
nand U6179 (N_6179,N_5869,N_5870);
or U6180 (N_6180,N_5965,N_5951);
nand U6181 (N_6181,N_5803,N_5965);
xnor U6182 (N_6182,N_5789,N_5712);
xnor U6183 (N_6183,N_5787,N_5858);
nand U6184 (N_6184,N_5750,N_5840);
xor U6185 (N_6185,N_5740,N_5790);
nor U6186 (N_6186,N_5793,N_5814);
or U6187 (N_6187,N_5853,N_5875);
xor U6188 (N_6188,N_5756,N_5763);
nor U6189 (N_6189,N_5962,N_5784);
xor U6190 (N_6190,N_5850,N_5780);
and U6191 (N_6191,N_5915,N_5781);
nand U6192 (N_6192,N_5980,N_5735);
xor U6193 (N_6193,N_5868,N_5827);
and U6194 (N_6194,N_5819,N_5712);
and U6195 (N_6195,N_5981,N_5917);
or U6196 (N_6196,N_5872,N_5877);
nor U6197 (N_6197,N_5768,N_5957);
or U6198 (N_6198,N_5752,N_5846);
nor U6199 (N_6199,N_5801,N_5836);
nand U6200 (N_6200,N_5958,N_5790);
xnor U6201 (N_6201,N_5744,N_5768);
xor U6202 (N_6202,N_5862,N_5820);
nor U6203 (N_6203,N_5701,N_5745);
nor U6204 (N_6204,N_5884,N_5810);
nand U6205 (N_6205,N_5849,N_5703);
or U6206 (N_6206,N_5827,N_5995);
nand U6207 (N_6207,N_5784,N_5858);
nor U6208 (N_6208,N_5731,N_5882);
xor U6209 (N_6209,N_5746,N_5716);
nand U6210 (N_6210,N_5721,N_5886);
nand U6211 (N_6211,N_5789,N_5982);
and U6212 (N_6212,N_5905,N_5843);
xor U6213 (N_6213,N_5982,N_5742);
nor U6214 (N_6214,N_5890,N_5705);
nor U6215 (N_6215,N_5730,N_5999);
and U6216 (N_6216,N_5967,N_5868);
or U6217 (N_6217,N_5932,N_5800);
and U6218 (N_6218,N_5989,N_5973);
nor U6219 (N_6219,N_5717,N_5711);
and U6220 (N_6220,N_5945,N_5781);
nand U6221 (N_6221,N_5750,N_5947);
nor U6222 (N_6222,N_5831,N_5931);
nand U6223 (N_6223,N_5963,N_5708);
and U6224 (N_6224,N_5897,N_5847);
or U6225 (N_6225,N_5812,N_5915);
and U6226 (N_6226,N_5898,N_5704);
or U6227 (N_6227,N_5743,N_5957);
nor U6228 (N_6228,N_5927,N_5809);
xnor U6229 (N_6229,N_5721,N_5733);
or U6230 (N_6230,N_5910,N_5991);
or U6231 (N_6231,N_5959,N_5723);
nor U6232 (N_6232,N_5763,N_5745);
nand U6233 (N_6233,N_5730,N_5758);
and U6234 (N_6234,N_5966,N_5765);
and U6235 (N_6235,N_5770,N_5792);
and U6236 (N_6236,N_5803,N_5859);
nor U6237 (N_6237,N_5984,N_5974);
or U6238 (N_6238,N_5975,N_5903);
nand U6239 (N_6239,N_5772,N_5862);
and U6240 (N_6240,N_5957,N_5715);
and U6241 (N_6241,N_5982,N_5903);
nor U6242 (N_6242,N_5707,N_5715);
nand U6243 (N_6243,N_5737,N_5858);
xnor U6244 (N_6244,N_5752,N_5842);
and U6245 (N_6245,N_5918,N_5979);
or U6246 (N_6246,N_5881,N_5729);
xor U6247 (N_6247,N_5960,N_5961);
xnor U6248 (N_6248,N_5762,N_5709);
or U6249 (N_6249,N_5984,N_5751);
xnor U6250 (N_6250,N_5769,N_5800);
nor U6251 (N_6251,N_5747,N_5996);
and U6252 (N_6252,N_5746,N_5872);
nor U6253 (N_6253,N_5895,N_5952);
nand U6254 (N_6254,N_5932,N_5861);
xnor U6255 (N_6255,N_5905,N_5980);
or U6256 (N_6256,N_5892,N_5712);
nor U6257 (N_6257,N_5837,N_5997);
nand U6258 (N_6258,N_5795,N_5826);
or U6259 (N_6259,N_5956,N_5952);
or U6260 (N_6260,N_5884,N_5804);
nand U6261 (N_6261,N_5895,N_5925);
or U6262 (N_6262,N_5888,N_5772);
and U6263 (N_6263,N_5827,N_5933);
nor U6264 (N_6264,N_5765,N_5795);
and U6265 (N_6265,N_5962,N_5746);
or U6266 (N_6266,N_5798,N_5750);
or U6267 (N_6267,N_5790,N_5854);
nor U6268 (N_6268,N_5802,N_5755);
and U6269 (N_6269,N_5910,N_5909);
nor U6270 (N_6270,N_5814,N_5864);
xnor U6271 (N_6271,N_5877,N_5837);
and U6272 (N_6272,N_5917,N_5924);
or U6273 (N_6273,N_5831,N_5872);
xnor U6274 (N_6274,N_5984,N_5979);
xor U6275 (N_6275,N_5997,N_5711);
nor U6276 (N_6276,N_5858,N_5935);
nand U6277 (N_6277,N_5827,N_5852);
xnor U6278 (N_6278,N_5954,N_5713);
xor U6279 (N_6279,N_5779,N_5899);
nand U6280 (N_6280,N_5723,N_5956);
nand U6281 (N_6281,N_5756,N_5947);
nand U6282 (N_6282,N_5990,N_5725);
and U6283 (N_6283,N_5902,N_5732);
and U6284 (N_6284,N_5820,N_5849);
xor U6285 (N_6285,N_5723,N_5847);
nand U6286 (N_6286,N_5767,N_5922);
nand U6287 (N_6287,N_5783,N_5987);
xor U6288 (N_6288,N_5837,N_5922);
xnor U6289 (N_6289,N_5935,N_5780);
nand U6290 (N_6290,N_5769,N_5896);
or U6291 (N_6291,N_5996,N_5760);
or U6292 (N_6292,N_5825,N_5970);
nor U6293 (N_6293,N_5724,N_5796);
nand U6294 (N_6294,N_5892,N_5998);
and U6295 (N_6295,N_5760,N_5701);
or U6296 (N_6296,N_5948,N_5915);
nand U6297 (N_6297,N_5853,N_5851);
xnor U6298 (N_6298,N_5709,N_5852);
xor U6299 (N_6299,N_5926,N_5807);
or U6300 (N_6300,N_6265,N_6091);
and U6301 (N_6301,N_6213,N_6177);
and U6302 (N_6302,N_6049,N_6042);
xnor U6303 (N_6303,N_6250,N_6240);
xor U6304 (N_6304,N_6053,N_6127);
and U6305 (N_6305,N_6179,N_6243);
nand U6306 (N_6306,N_6267,N_6224);
and U6307 (N_6307,N_6124,N_6286);
xnor U6308 (N_6308,N_6114,N_6222);
xnor U6309 (N_6309,N_6132,N_6058);
nor U6310 (N_6310,N_6256,N_6219);
nor U6311 (N_6311,N_6043,N_6259);
xnor U6312 (N_6312,N_6068,N_6212);
nand U6313 (N_6313,N_6063,N_6125);
nand U6314 (N_6314,N_6210,N_6131);
nor U6315 (N_6315,N_6294,N_6065);
nand U6316 (N_6316,N_6180,N_6153);
and U6317 (N_6317,N_6106,N_6077);
or U6318 (N_6318,N_6261,N_6118);
nor U6319 (N_6319,N_6099,N_6148);
xor U6320 (N_6320,N_6023,N_6150);
xnor U6321 (N_6321,N_6012,N_6297);
or U6322 (N_6322,N_6191,N_6158);
nor U6323 (N_6323,N_6190,N_6088);
nand U6324 (N_6324,N_6016,N_6045);
or U6325 (N_6325,N_6144,N_6229);
nor U6326 (N_6326,N_6247,N_6037);
nand U6327 (N_6327,N_6123,N_6139);
or U6328 (N_6328,N_6014,N_6225);
nor U6329 (N_6329,N_6112,N_6075);
nor U6330 (N_6330,N_6015,N_6121);
and U6331 (N_6331,N_6167,N_6164);
and U6332 (N_6332,N_6149,N_6097);
xnor U6333 (N_6333,N_6020,N_6241);
nor U6334 (N_6334,N_6017,N_6258);
nand U6335 (N_6335,N_6296,N_6071);
or U6336 (N_6336,N_6155,N_6072);
nand U6337 (N_6337,N_6070,N_6129);
xnor U6338 (N_6338,N_6178,N_6052);
nand U6339 (N_6339,N_6204,N_6059);
nor U6340 (N_6340,N_6223,N_6298);
nand U6341 (N_6341,N_6232,N_6018);
nand U6342 (N_6342,N_6001,N_6218);
or U6343 (N_6343,N_6110,N_6120);
or U6344 (N_6344,N_6086,N_6207);
or U6345 (N_6345,N_6184,N_6214);
nand U6346 (N_6346,N_6032,N_6255);
nor U6347 (N_6347,N_6274,N_6287);
nand U6348 (N_6348,N_6289,N_6067);
xnor U6349 (N_6349,N_6084,N_6085);
and U6350 (N_6350,N_6281,N_6299);
nand U6351 (N_6351,N_6290,N_6193);
xor U6352 (N_6352,N_6007,N_6248);
xnor U6353 (N_6353,N_6116,N_6113);
or U6354 (N_6354,N_6292,N_6126);
nand U6355 (N_6355,N_6137,N_6119);
nor U6356 (N_6356,N_6117,N_6040);
or U6357 (N_6357,N_6244,N_6048);
xnor U6358 (N_6358,N_6203,N_6216);
and U6359 (N_6359,N_6080,N_6231);
xnor U6360 (N_6360,N_6188,N_6268);
nor U6361 (N_6361,N_6108,N_6079);
xnor U6362 (N_6362,N_6227,N_6090);
or U6363 (N_6363,N_6027,N_6073);
and U6364 (N_6364,N_6181,N_6235);
nor U6365 (N_6365,N_6279,N_6169);
or U6366 (N_6366,N_6271,N_6262);
and U6367 (N_6367,N_6096,N_6002);
nand U6368 (N_6368,N_6173,N_6208);
nand U6369 (N_6369,N_6233,N_6172);
nor U6370 (N_6370,N_6009,N_6295);
xor U6371 (N_6371,N_6003,N_6192);
or U6372 (N_6372,N_6034,N_6162);
nor U6373 (N_6373,N_6130,N_6076);
xor U6374 (N_6374,N_6205,N_6157);
or U6375 (N_6375,N_6128,N_6101);
or U6376 (N_6376,N_6095,N_6238);
and U6377 (N_6377,N_6166,N_6004);
and U6378 (N_6378,N_6031,N_6064);
or U6379 (N_6379,N_6107,N_6239);
nand U6380 (N_6380,N_6154,N_6082);
and U6381 (N_6381,N_6156,N_6038);
nor U6382 (N_6382,N_6275,N_6060);
nand U6383 (N_6383,N_6291,N_6028);
and U6384 (N_6384,N_6021,N_6211);
and U6385 (N_6385,N_6026,N_6109);
and U6386 (N_6386,N_6094,N_6252);
and U6387 (N_6387,N_6196,N_6103);
xnor U6388 (N_6388,N_6189,N_6257);
nand U6389 (N_6389,N_6185,N_6264);
or U6390 (N_6390,N_6285,N_6140);
or U6391 (N_6391,N_6022,N_6010);
nor U6392 (N_6392,N_6242,N_6276);
nand U6393 (N_6393,N_6019,N_6260);
or U6394 (N_6394,N_6175,N_6174);
and U6395 (N_6395,N_6221,N_6011);
nor U6396 (N_6396,N_6236,N_6098);
nand U6397 (N_6397,N_6036,N_6284);
nor U6398 (N_6398,N_6066,N_6230);
nand U6399 (N_6399,N_6138,N_6074);
xnor U6400 (N_6400,N_6089,N_6092);
xor U6401 (N_6401,N_6163,N_6033);
and U6402 (N_6402,N_6263,N_6159);
nor U6403 (N_6403,N_6000,N_6194);
and U6404 (N_6404,N_6087,N_6245);
or U6405 (N_6405,N_6270,N_6135);
or U6406 (N_6406,N_6186,N_6100);
nand U6407 (N_6407,N_6145,N_6209);
or U6408 (N_6408,N_6187,N_6199);
nand U6409 (N_6409,N_6057,N_6115);
and U6410 (N_6410,N_6134,N_6136);
or U6411 (N_6411,N_6217,N_6030);
or U6412 (N_6412,N_6054,N_6168);
or U6413 (N_6413,N_6201,N_6046);
and U6414 (N_6414,N_6039,N_6215);
xnor U6415 (N_6415,N_6234,N_6249);
nor U6416 (N_6416,N_6288,N_6269);
or U6417 (N_6417,N_6282,N_6226);
nor U6418 (N_6418,N_6151,N_6293);
or U6419 (N_6419,N_6202,N_6013);
nand U6420 (N_6420,N_6147,N_6228);
and U6421 (N_6421,N_6025,N_6006);
or U6422 (N_6422,N_6143,N_6195);
or U6423 (N_6423,N_6104,N_6220);
xnor U6424 (N_6424,N_6083,N_6253);
xor U6425 (N_6425,N_6206,N_6024);
xor U6426 (N_6426,N_6005,N_6122);
or U6427 (N_6427,N_6246,N_6283);
xor U6428 (N_6428,N_6272,N_6176);
nand U6429 (N_6429,N_6183,N_6062);
and U6430 (N_6430,N_6160,N_6041);
and U6431 (N_6431,N_6266,N_6047);
nor U6432 (N_6432,N_6198,N_6251);
xor U6433 (N_6433,N_6141,N_6161);
xor U6434 (N_6434,N_6278,N_6200);
xor U6435 (N_6435,N_6069,N_6170);
xor U6436 (N_6436,N_6093,N_6197);
xnor U6437 (N_6437,N_6105,N_6044);
or U6438 (N_6438,N_6050,N_6171);
nor U6439 (N_6439,N_6152,N_6182);
nand U6440 (N_6440,N_6111,N_6056);
or U6441 (N_6441,N_6078,N_6061);
and U6442 (N_6442,N_6280,N_6008);
nor U6443 (N_6443,N_6237,N_6142);
nand U6444 (N_6444,N_6254,N_6273);
nor U6445 (N_6445,N_6146,N_6051);
or U6446 (N_6446,N_6133,N_6102);
xnor U6447 (N_6447,N_6029,N_6035);
xor U6448 (N_6448,N_6081,N_6165);
xor U6449 (N_6449,N_6277,N_6055);
and U6450 (N_6450,N_6249,N_6051);
nor U6451 (N_6451,N_6032,N_6052);
nand U6452 (N_6452,N_6170,N_6078);
nor U6453 (N_6453,N_6157,N_6124);
and U6454 (N_6454,N_6084,N_6168);
or U6455 (N_6455,N_6033,N_6201);
and U6456 (N_6456,N_6065,N_6175);
nand U6457 (N_6457,N_6253,N_6118);
nand U6458 (N_6458,N_6052,N_6187);
nand U6459 (N_6459,N_6266,N_6042);
xor U6460 (N_6460,N_6244,N_6030);
xor U6461 (N_6461,N_6112,N_6259);
nor U6462 (N_6462,N_6158,N_6200);
nand U6463 (N_6463,N_6131,N_6231);
nand U6464 (N_6464,N_6150,N_6042);
nand U6465 (N_6465,N_6232,N_6254);
nor U6466 (N_6466,N_6155,N_6119);
or U6467 (N_6467,N_6001,N_6237);
or U6468 (N_6468,N_6099,N_6089);
or U6469 (N_6469,N_6030,N_6122);
and U6470 (N_6470,N_6116,N_6182);
nor U6471 (N_6471,N_6231,N_6060);
nand U6472 (N_6472,N_6198,N_6013);
and U6473 (N_6473,N_6048,N_6158);
and U6474 (N_6474,N_6219,N_6162);
and U6475 (N_6475,N_6011,N_6116);
or U6476 (N_6476,N_6218,N_6145);
xnor U6477 (N_6477,N_6044,N_6001);
xnor U6478 (N_6478,N_6088,N_6133);
nand U6479 (N_6479,N_6286,N_6208);
xor U6480 (N_6480,N_6110,N_6209);
nand U6481 (N_6481,N_6163,N_6070);
or U6482 (N_6482,N_6297,N_6141);
nand U6483 (N_6483,N_6200,N_6228);
xor U6484 (N_6484,N_6082,N_6008);
nand U6485 (N_6485,N_6154,N_6242);
nor U6486 (N_6486,N_6248,N_6179);
or U6487 (N_6487,N_6248,N_6187);
xor U6488 (N_6488,N_6012,N_6094);
and U6489 (N_6489,N_6227,N_6118);
nor U6490 (N_6490,N_6145,N_6210);
nor U6491 (N_6491,N_6295,N_6282);
nand U6492 (N_6492,N_6262,N_6017);
or U6493 (N_6493,N_6217,N_6008);
nand U6494 (N_6494,N_6180,N_6192);
and U6495 (N_6495,N_6165,N_6045);
or U6496 (N_6496,N_6299,N_6170);
nand U6497 (N_6497,N_6102,N_6065);
xnor U6498 (N_6498,N_6193,N_6214);
or U6499 (N_6499,N_6296,N_6026);
and U6500 (N_6500,N_6041,N_6044);
nand U6501 (N_6501,N_6060,N_6033);
or U6502 (N_6502,N_6178,N_6263);
or U6503 (N_6503,N_6031,N_6081);
nor U6504 (N_6504,N_6150,N_6154);
xnor U6505 (N_6505,N_6238,N_6142);
and U6506 (N_6506,N_6110,N_6155);
and U6507 (N_6507,N_6049,N_6115);
or U6508 (N_6508,N_6175,N_6153);
nor U6509 (N_6509,N_6042,N_6106);
nand U6510 (N_6510,N_6065,N_6159);
and U6511 (N_6511,N_6293,N_6298);
and U6512 (N_6512,N_6139,N_6269);
xor U6513 (N_6513,N_6297,N_6191);
and U6514 (N_6514,N_6283,N_6256);
and U6515 (N_6515,N_6165,N_6102);
nor U6516 (N_6516,N_6057,N_6203);
nor U6517 (N_6517,N_6044,N_6012);
or U6518 (N_6518,N_6259,N_6287);
and U6519 (N_6519,N_6123,N_6228);
nor U6520 (N_6520,N_6065,N_6248);
nor U6521 (N_6521,N_6281,N_6024);
and U6522 (N_6522,N_6024,N_6299);
nand U6523 (N_6523,N_6233,N_6109);
nand U6524 (N_6524,N_6290,N_6036);
nor U6525 (N_6525,N_6006,N_6120);
xnor U6526 (N_6526,N_6272,N_6213);
nor U6527 (N_6527,N_6115,N_6172);
nand U6528 (N_6528,N_6193,N_6172);
or U6529 (N_6529,N_6071,N_6215);
and U6530 (N_6530,N_6123,N_6012);
nand U6531 (N_6531,N_6048,N_6259);
and U6532 (N_6532,N_6179,N_6220);
nor U6533 (N_6533,N_6294,N_6129);
nand U6534 (N_6534,N_6085,N_6267);
xnor U6535 (N_6535,N_6177,N_6197);
or U6536 (N_6536,N_6251,N_6159);
or U6537 (N_6537,N_6092,N_6035);
nand U6538 (N_6538,N_6216,N_6215);
nor U6539 (N_6539,N_6139,N_6287);
xnor U6540 (N_6540,N_6202,N_6170);
nor U6541 (N_6541,N_6020,N_6140);
or U6542 (N_6542,N_6174,N_6029);
nor U6543 (N_6543,N_6148,N_6064);
xor U6544 (N_6544,N_6194,N_6083);
xnor U6545 (N_6545,N_6002,N_6054);
xnor U6546 (N_6546,N_6010,N_6248);
or U6547 (N_6547,N_6122,N_6265);
xor U6548 (N_6548,N_6282,N_6025);
nand U6549 (N_6549,N_6173,N_6110);
nor U6550 (N_6550,N_6194,N_6283);
and U6551 (N_6551,N_6292,N_6253);
and U6552 (N_6552,N_6177,N_6210);
nor U6553 (N_6553,N_6038,N_6238);
nor U6554 (N_6554,N_6021,N_6287);
nor U6555 (N_6555,N_6079,N_6158);
or U6556 (N_6556,N_6269,N_6110);
xnor U6557 (N_6557,N_6128,N_6213);
nor U6558 (N_6558,N_6278,N_6055);
nand U6559 (N_6559,N_6075,N_6215);
nand U6560 (N_6560,N_6141,N_6025);
nand U6561 (N_6561,N_6212,N_6168);
nand U6562 (N_6562,N_6075,N_6046);
xnor U6563 (N_6563,N_6149,N_6197);
or U6564 (N_6564,N_6262,N_6221);
nand U6565 (N_6565,N_6156,N_6081);
and U6566 (N_6566,N_6188,N_6194);
xor U6567 (N_6567,N_6095,N_6015);
nor U6568 (N_6568,N_6279,N_6007);
or U6569 (N_6569,N_6027,N_6100);
xor U6570 (N_6570,N_6060,N_6041);
xor U6571 (N_6571,N_6211,N_6193);
or U6572 (N_6572,N_6022,N_6209);
nand U6573 (N_6573,N_6161,N_6204);
xnor U6574 (N_6574,N_6017,N_6214);
xnor U6575 (N_6575,N_6195,N_6276);
and U6576 (N_6576,N_6271,N_6108);
nor U6577 (N_6577,N_6153,N_6215);
or U6578 (N_6578,N_6049,N_6279);
xnor U6579 (N_6579,N_6188,N_6233);
nor U6580 (N_6580,N_6299,N_6217);
and U6581 (N_6581,N_6000,N_6060);
or U6582 (N_6582,N_6178,N_6240);
nor U6583 (N_6583,N_6094,N_6255);
xor U6584 (N_6584,N_6162,N_6039);
xnor U6585 (N_6585,N_6196,N_6027);
xor U6586 (N_6586,N_6229,N_6250);
and U6587 (N_6587,N_6295,N_6093);
nor U6588 (N_6588,N_6249,N_6199);
and U6589 (N_6589,N_6213,N_6079);
xnor U6590 (N_6590,N_6164,N_6181);
and U6591 (N_6591,N_6060,N_6028);
nor U6592 (N_6592,N_6083,N_6042);
xor U6593 (N_6593,N_6195,N_6002);
or U6594 (N_6594,N_6255,N_6050);
and U6595 (N_6595,N_6058,N_6279);
and U6596 (N_6596,N_6095,N_6056);
nor U6597 (N_6597,N_6147,N_6208);
and U6598 (N_6598,N_6232,N_6069);
xnor U6599 (N_6599,N_6070,N_6031);
nor U6600 (N_6600,N_6353,N_6418);
nor U6601 (N_6601,N_6582,N_6317);
xor U6602 (N_6602,N_6384,N_6374);
nand U6603 (N_6603,N_6562,N_6462);
nand U6604 (N_6604,N_6400,N_6505);
or U6605 (N_6605,N_6307,N_6591);
nor U6606 (N_6606,N_6388,N_6576);
nor U6607 (N_6607,N_6381,N_6389);
or U6608 (N_6608,N_6395,N_6529);
and U6609 (N_6609,N_6548,N_6579);
nand U6610 (N_6610,N_6348,N_6513);
or U6611 (N_6611,N_6435,N_6446);
and U6612 (N_6612,N_6492,N_6525);
nand U6613 (N_6613,N_6451,N_6373);
nor U6614 (N_6614,N_6394,N_6443);
nand U6615 (N_6615,N_6523,N_6588);
nand U6616 (N_6616,N_6575,N_6584);
xnor U6617 (N_6617,N_6300,N_6427);
xnor U6618 (N_6618,N_6482,N_6517);
and U6619 (N_6619,N_6314,N_6372);
or U6620 (N_6620,N_6359,N_6557);
nor U6621 (N_6621,N_6397,N_6454);
nand U6622 (N_6622,N_6542,N_6409);
or U6623 (N_6623,N_6500,N_6568);
xor U6624 (N_6624,N_6577,N_6375);
nand U6625 (N_6625,N_6530,N_6464);
nor U6626 (N_6626,N_6326,N_6340);
and U6627 (N_6627,N_6324,N_6322);
and U6628 (N_6628,N_6356,N_6350);
or U6629 (N_6629,N_6567,N_6479);
xnor U6630 (N_6630,N_6485,N_6414);
and U6631 (N_6631,N_6571,N_6332);
and U6632 (N_6632,N_6501,N_6558);
nand U6633 (N_6633,N_6364,N_6316);
nand U6634 (N_6634,N_6449,N_6452);
nor U6635 (N_6635,N_6483,N_6425);
xor U6636 (N_6636,N_6396,N_6367);
nor U6637 (N_6637,N_6407,N_6382);
nor U6638 (N_6638,N_6355,N_6599);
nor U6639 (N_6639,N_6570,N_6403);
nand U6640 (N_6640,N_6554,N_6478);
or U6641 (N_6641,N_6553,N_6448);
xor U6642 (N_6642,N_6499,N_6420);
nand U6643 (N_6643,N_6543,N_6487);
nand U6644 (N_6644,N_6460,N_6555);
and U6645 (N_6645,N_6365,N_6496);
or U6646 (N_6646,N_6419,N_6323);
and U6647 (N_6647,N_6561,N_6327);
or U6648 (N_6648,N_6595,N_6472);
nor U6649 (N_6649,N_6301,N_6598);
nand U6650 (N_6650,N_6559,N_6309);
nor U6651 (N_6651,N_6578,N_6489);
xor U6652 (N_6652,N_6539,N_6563);
and U6653 (N_6653,N_6380,N_6476);
nor U6654 (N_6654,N_6336,N_6346);
and U6655 (N_6655,N_6508,N_6383);
and U6656 (N_6656,N_6502,N_6564);
nand U6657 (N_6657,N_6371,N_6465);
and U6658 (N_6658,N_6376,N_6402);
nor U6659 (N_6659,N_6410,N_6440);
nand U6660 (N_6660,N_6593,N_6498);
nor U6661 (N_6661,N_6484,N_6493);
nor U6662 (N_6662,N_6426,N_6412);
nand U6663 (N_6663,N_6488,N_6325);
nand U6664 (N_6664,N_6428,N_6431);
xor U6665 (N_6665,N_6461,N_6321);
xor U6666 (N_6666,N_6315,N_6494);
xnor U6667 (N_6667,N_6444,N_6587);
xor U6668 (N_6668,N_6515,N_6308);
xnor U6669 (N_6669,N_6415,N_6351);
or U6670 (N_6670,N_6343,N_6437);
nor U6671 (N_6671,N_6497,N_6596);
xnor U6672 (N_6672,N_6399,N_6469);
xnor U6673 (N_6673,N_6463,N_6474);
or U6674 (N_6674,N_6586,N_6337);
xnor U6675 (N_6675,N_6320,N_6349);
nand U6676 (N_6676,N_6572,N_6527);
or U6677 (N_6677,N_6522,N_6470);
xor U6678 (N_6678,N_6339,N_6416);
and U6679 (N_6679,N_6441,N_6556);
or U6680 (N_6680,N_6512,N_6581);
and U6681 (N_6681,N_6473,N_6592);
nor U6682 (N_6682,N_6541,N_6358);
xor U6683 (N_6683,N_6370,N_6342);
nor U6684 (N_6684,N_6516,N_6504);
xor U6685 (N_6685,N_6503,N_6331);
xnor U6686 (N_6686,N_6589,N_6368);
nand U6687 (N_6687,N_6413,N_6514);
nor U6688 (N_6688,N_6405,N_6585);
xor U6689 (N_6689,N_6490,N_6534);
nand U6690 (N_6690,N_6573,N_6310);
nand U6691 (N_6691,N_6574,N_6481);
and U6692 (N_6692,N_6477,N_6361);
or U6693 (N_6693,N_6552,N_6445);
or U6694 (N_6694,N_6520,N_6486);
and U6695 (N_6695,N_6432,N_6304);
or U6696 (N_6696,N_6433,N_6495);
or U6697 (N_6697,N_6545,N_6392);
xnor U6698 (N_6698,N_6305,N_6533);
nand U6699 (N_6699,N_6546,N_6347);
nand U6700 (N_6700,N_6569,N_6471);
nand U6701 (N_6701,N_6518,N_6436);
nor U6702 (N_6702,N_6306,N_6366);
xor U6703 (N_6703,N_6531,N_6565);
or U6704 (N_6704,N_6458,N_6362);
nand U6705 (N_6705,N_6333,N_6434);
xnor U6706 (N_6706,N_6302,N_6447);
nand U6707 (N_6707,N_6597,N_6429);
or U6708 (N_6708,N_6453,N_6424);
nor U6709 (N_6709,N_6551,N_6345);
and U6710 (N_6710,N_6590,N_6526);
xnor U6711 (N_6711,N_6338,N_6456);
and U6712 (N_6712,N_6430,N_6311);
and U6713 (N_6713,N_6450,N_6401);
xor U6714 (N_6714,N_6580,N_6510);
or U6715 (N_6715,N_6385,N_6538);
nor U6716 (N_6716,N_6344,N_6594);
or U6717 (N_6717,N_6330,N_6536);
nand U6718 (N_6718,N_6411,N_6377);
nor U6719 (N_6719,N_6352,N_6519);
xor U6720 (N_6720,N_6303,N_6480);
or U6721 (N_6721,N_6438,N_6335);
or U6722 (N_6722,N_6406,N_6532);
nor U6723 (N_6723,N_6421,N_6360);
or U6724 (N_6724,N_6475,N_6491);
nand U6725 (N_6725,N_6468,N_6540);
nand U6726 (N_6726,N_6398,N_6455);
nor U6727 (N_6727,N_6408,N_6369);
nand U6728 (N_6728,N_6459,N_6312);
nor U6729 (N_6729,N_6391,N_6319);
and U6730 (N_6730,N_6549,N_6457);
xnor U6731 (N_6731,N_6387,N_6439);
nor U6732 (N_6732,N_6357,N_6524);
xor U6733 (N_6733,N_6404,N_6442);
or U6734 (N_6734,N_6417,N_6544);
nand U6735 (N_6735,N_6509,N_6537);
and U6736 (N_6736,N_6560,N_6378);
or U6737 (N_6737,N_6528,N_6390);
or U6738 (N_6738,N_6393,N_6422);
nor U6739 (N_6739,N_6328,N_6511);
or U6740 (N_6740,N_6379,N_6341);
nor U6741 (N_6741,N_6466,N_6318);
or U6742 (N_6742,N_6583,N_6386);
and U6743 (N_6743,N_6566,N_6507);
or U6744 (N_6744,N_6506,N_6550);
xnor U6745 (N_6745,N_6521,N_6329);
nand U6746 (N_6746,N_6535,N_6334);
and U6747 (N_6747,N_6547,N_6354);
nand U6748 (N_6748,N_6423,N_6363);
or U6749 (N_6749,N_6313,N_6467);
or U6750 (N_6750,N_6559,N_6358);
and U6751 (N_6751,N_6392,N_6425);
nor U6752 (N_6752,N_6475,N_6324);
xnor U6753 (N_6753,N_6589,N_6315);
nand U6754 (N_6754,N_6509,N_6373);
and U6755 (N_6755,N_6564,N_6438);
nand U6756 (N_6756,N_6313,N_6407);
nand U6757 (N_6757,N_6398,N_6495);
nand U6758 (N_6758,N_6516,N_6541);
nand U6759 (N_6759,N_6354,N_6361);
xor U6760 (N_6760,N_6532,N_6593);
nor U6761 (N_6761,N_6404,N_6406);
nor U6762 (N_6762,N_6317,N_6319);
nand U6763 (N_6763,N_6442,N_6389);
nor U6764 (N_6764,N_6594,N_6316);
xor U6765 (N_6765,N_6417,N_6580);
or U6766 (N_6766,N_6395,N_6330);
nand U6767 (N_6767,N_6520,N_6316);
or U6768 (N_6768,N_6539,N_6491);
xor U6769 (N_6769,N_6441,N_6564);
nor U6770 (N_6770,N_6397,N_6573);
nand U6771 (N_6771,N_6407,N_6584);
nand U6772 (N_6772,N_6363,N_6325);
xor U6773 (N_6773,N_6343,N_6344);
and U6774 (N_6774,N_6559,N_6534);
or U6775 (N_6775,N_6364,N_6306);
and U6776 (N_6776,N_6396,N_6479);
and U6777 (N_6777,N_6577,N_6479);
and U6778 (N_6778,N_6444,N_6354);
xnor U6779 (N_6779,N_6393,N_6562);
nor U6780 (N_6780,N_6483,N_6442);
and U6781 (N_6781,N_6365,N_6420);
nand U6782 (N_6782,N_6448,N_6403);
nor U6783 (N_6783,N_6497,N_6494);
nor U6784 (N_6784,N_6576,N_6425);
or U6785 (N_6785,N_6482,N_6564);
nand U6786 (N_6786,N_6392,N_6447);
and U6787 (N_6787,N_6438,N_6484);
xnor U6788 (N_6788,N_6503,N_6535);
or U6789 (N_6789,N_6413,N_6406);
or U6790 (N_6790,N_6301,N_6431);
and U6791 (N_6791,N_6310,N_6517);
nand U6792 (N_6792,N_6398,N_6347);
and U6793 (N_6793,N_6595,N_6441);
and U6794 (N_6794,N_6497,N_6307);
and U6795 (N_6795,N_6547,N_6398);
xnor U6796 (N_6796,N_6362,N_6596);
xnor U6797 (N_6797,N_6442,N_6481);
xnor U6798 (N_6798,N_6395,N_6389);
and U6799 (N_6799,N_6426,N_6445);
xnor U6800 (N_6800,N_6560,N_6359);
nor U6801 (N_6801,N_6368,N_6574);
xor U6802 (N_6802,N_6555,N_6386);
nor U6803 (N_6803,N_6404,N_6545);
and U6804 (N_6804,N_6318,N_6453);
xor U6805 (N_6805,N_6595,N_6473);
or U6806 (N_6806,N_6354,N_6380);
xor U6807 (N_6807,N_6419,N_6315);
or U6808 (N_6808,N_6395,N_6525);
or U6809 (N_6809,N_6316,N_6428);
or U6810 (N_6810,N_6415,N_6383);
nor U6811 (N_6811,N_6425,N_6528);
nand U6812 (N_6812,N_6424,N_6313);
or U6813 (N_6813,N_6510,N_6362);
xor U6814 (N_6814,N_6457,N_6330);
nor U6815 (N_6815,N_6568,N_6442);
and U6816 (N_6816,N_6314,N_6461);
and U6817 (N_6817,N_6573,N_6384);
nor U6818 (N_6818,N_6325,N_6569);
nand U6819 (N_6819,N_6440,N_6422);
xnor U6820 (N_6820,N_6415,N_6426);
nor U6821 (N_6821,N_6489,N_6400);
nand U6822 (N_6822,N_6489,N_6478);
and U6823 (N_6823,N_6356,N_6599);
and U6824 (N_6824,N_6336,N_6530);
xor U6825 (N_6825,N_6538,N_6311);
xnor U6826 (N_6826,N_6320,N_6548);
or U6827 (N_6827,N_6570,N_6596);
nand U6828 (N_6828,N_6459,N_6585);
xnor U6829 (N_6829,N_6371,N_6479);
xnor U6830 (N_6830,N_6596,N_6496);
xor U6831 (N_6831,N_6316,N_6383);
nand U6832 (N_6832,N_6525,N_6305);
nor U6833 (N_6833,N_6387,N_6338);
xnor U6834 (N_6834,N_6321,N_6585);
or U6835 (N_6835,N_6314,N_6591);
nand U6836 (N_6836,N_6513,N_6571);
nor U6837 (N_6837,N_6336,N_6516);
or U6838 (N_6838,N_6308,N_6506);
xnor U6839 (N_6839,N_6416,N_6526);
and U6840 (N_6840,N_6412,N_6569);
xnor U6841 (N_6841,N_6446,N_6413);
and U6842 (N_6842,N_6429,N_6446);
or U6843 (N_6843,N_6435,N_6443);
xnor U6844 (N_6844,N_6356,N_6503);
nand U6845 (N_6845,N_6467,N_6428);
or U6846 (N_6846,N_6563,N_6598);
or U6847 (N_6847,N_6552,N_6554);
nor U6848 (N_6848,N_6365,N_6446);
nor U6849 (N_6849,N_6446,N_6375);
nor U6850 (N_6850,N_6352,N_6313);
nor U6851 (N_6851,N_6304,N_6496);
xor U6852 (N_6852,N_6303,N_6313);
xor U6853 (N_6853,N_6571,N_6595);
and U6854 (N_6854,N_6337,N_6307);
or U6855 (N_6855,N_6569,N_6375);
and U6856 (N_6856,N_6437,N_6380);
xnor U6857 (N_6857,N_6495,N_6598);
nand U6858 (N_6858,N_6524,N_6495);
nand U6859 (N_6859,N_6390,N_6431);
xnor U6860 (N_6860,N_6432,N_6341);
nand U6861 (N_6861,N_6408,N_6481);
nand U6862 (N_6862,N_6370,N_6514);
nand U6863 (N_6863,N_6470,N_6546);
and U6864 (N_6864,N_6515,N_6582);
or U6865 (N_6865,N_6399,N_6470);
and U6866 (N_6866,N_6300,N_6404);
xor U6867 (N_6867,N_6314,N_6385);
or U6868 (N_6868,N_6415,N_6473);
nor U6869 (N_6869,N_6363,N_6368);
nor U6870 (N_6870,N_6463,N_6444);
nand U6871 (N_6871,N_6532,N_6334);
or U6872 (N_6872,N_6336,N_6356);
xor U6873 (N_6873,N_6314,N_6406);
nor U6874 (N_6874,N_6498,N_6457);
nor U6875 (N_6875,N_6325,N_6476);
nor U6876 (N_6876,N_6396,N_6459);
or U6877 (N_6877,N_6362,N_6599);
or U6878 (N_6878,N_6597,N_6352);
xor U6879 (N_6879,N_6380,N_6556);
and U6880 (N_6880,N_6501,N_6517);
xnor U6881 (N_6881,N_6371,N_6363);
and U6882 (N_6882,N_6559,N_6466);
or U6883 (N_6883,N_6324,N_6561);
or U6884 (N_6884,N_6494,N_6448);
nand U6885 (N_6885,N_6372,N_6433);
and U6886 (N_6886,N_6448,N_6487);
nor U6887 (N_6887,N_6373,N_6576);
xor U6888 (N_6888,N_6518,N_6530);
or U6889 (N_6889,N_6363,N_6352);
or U6890 (N_6890,N_6420,N_6437);
nor U6891 (N_6891,N_6554,N_6527);
and U6892 (N_6892,N_6553,N_6514);
nand U6893 (N_6893,N_6342,N_6358);
or U6894 (N_6894,N_6563,N_6463);
nor U6895 (N_6895,N_6488,N_6412);
nor U6896 (N_6896,N_6591,N_6337);
nor U6897 (N_6897,N_6533,N_6407);
and U6898 (N_6898,N_6551,N_6390);
nand U6899 (N_6899,N_6371,N_6345);
xor U6900 (N_6900,N_6696,N_6871);
xor U6901 (N_6901,N_6748,N_6688);
xnor U6902 (N_6902,N_6681,N_6726);
and U6903 (N_6903,N_6812,N_6623);
and U6904 (N_6904,N_6723,N_6889);
or U6905 (N_6905,N_6783,N_6790);
nor U6906 (N_6906,N_6635,N_6788);
xnor U6907 (N_6907,N_6618,N_6606);
and U6908 (N_6908,N_6874,N_6837);
and U6909 (N_6909,N_6785,N_6757);
nand U6910 (N_6910,N_6625,N_6722);
nand U6911 (N_6911,N_6829,N_6714);
or U6912 (N_6912,N_6744,N_6616);
or U6913 (N_6913,N_6642,N_6737);
nand U6914 (N_6914,N_6674,N_6730);
nand U6915 (N_6915,N_6878,N_6686);
or U6916 (N_6916,N_6643,N_6716);
or U6917 (N_6917,N_6665,N_6848);
and U6918 (N_6918,N_6819,N_6866);
xor U6919 (N_6919,N_6739,N_6808);
and U6920 (N_6920,N_6891,N_6633);
and U6921 (N_6921,N_6738,N_6707);
or U6922 (N_6922,N_6851,N_6823);
xor U6923 (N_6923,N_6613,N_6895);
nor U6924 (N_6924,N_6845,N_6651);
or U6925 (N_6925,N_6787,N_6774);
and U6926 (N_6926,N_6600,N_6629);
nor U6927 (N_6927,N_6666,N_6610);
or U6928 (N_6928,N_6863,N_6644);
or U6929 (N_6929,N_6695,N_6641);
or U6930 (N_6930,N_6862,N_6800);
nor U6931 (N_6931,N_6830,N_6620);
nor U6932 (N_6932,N_6802,N_6685);
nand U6933 (N_6933,N_6835,N_6637);
xor U6934 (N_6934,N_6877,N_6694);
nor U6935 (N_6935,N_6728,N_6631);
and U6936 (N_6936,N_6893,N_6670);
or U6937 (N_6937,N_6806,N_6619);
nor U6938 (N_6938,N_6671,N_6669);
xnor U6939 (N_6939,N_6883,N_6717);
nand U6940 (N_6940,N_6655,N_6745);
xor U6941 (N_6941,N_6645,N_6750);
xor U6942 (N_6942,N_6746,N_6693);
or U6943 (N_6943,N_6658,N_6634);
nand U6944 (N_6944,N_6626,N_6821);
nor U6945 (N_6945,N_6804,N_6697);
nor U6946 (N_6946,N_6815,N_6660);
or U6947 (N_6947,N_6715,N_6628);
xor U6948 (N_6948,N_6896,N_6703);
xnor U6949 (N_6949,N_6838,N_6736);
nor U6950 (N_6950,N_6711,N_6720);
nand U6951 (N_6951,N_6710,N_6854);
xnor U6952 (N_6952,N_6604,N_6791);
or U6953 (N_6953,N_6731,N_6872);
xor U6954 (N_6954,N_6782,N_6667);
nand U6955 (N_6955,N_6621,N_6640);
nor U6956 (N_6956,N_6760,N_6721);
nor U6957 (N_6957,N_6868,N_6807);
nor U6958 (N_6958,N_6701,N_6841);
and U6959 (N_6959,N_6647,N_6803);
and U6960 (N_6960,N_6649,N_6733);
xor U6961 (N_6961,N_6654,N_6755);
nand U6962 (N_6962,N_6776,N_6741);
nand U6963 (N_6963,N_6699,N_6826);
and U6964 (N_6964,N_6814,N_6622);
xnor U6965 (N_6965,N_6691,N_6801);
or U6966 (N_6966,N_6844,N_6885);
nand U6967 (N_6967,N_6832,N_6767);
nor U6968 (N_6968,N_6831,N_6648);
xnor U6969 (N_6969,N_6705,N_6784);
nor U6970 (N_6970,N_6611,N_6735);
or U6971 (N_6971,N_6601,N_6873);
and U6972 (N_6972,N_6798,N_6754);
and U6973 (N_6973,N_6780,N_6732);
and U6974 (N_6974,N_6657,N_6865);
xnor U6975 (N_6975,N_6608,N_6759);
or U6976 (N_6976,N_6603,N_6857);
nand U6977 (N_6977,N_6663,N_6743);
nand U6978 (N_6978,N_6624,N_6605);
or U6979 (N_6979,N_6880,N_6734);
nand U6980 (N_6980,N_6638,N_6824);
nand U6981 (N_6981,N_6779,N_6692);
nor U6982 (N_6982,N_6842,N_6795);
nand U6983 (N_6983,N_6833,N_6789);
or U6984 (N_6984,N_6849,N_6724);
and U6985 (N_6985,N_6810,N_6747);
xnor U6986 (N_6986,N_6664,N_6709);
and U6987 (N_6987,N_6888,N_6775);
xor U6988 (N_6988,N_6773,N_6673);
or U6989 (N_6989,N_6828,N_6676);
nand U6990 (N_6990,N_6811,N_6727);
nor U6991 (N_6991,N_6753,N_6713);
and U6992 (N_6992,N_6698,N_6839);
nand U6993 (N_6993,N_6627,N_6708);
xnor U6994 (N_6994,N_6702,N_6672);
xnor U6995 (N_6995,N_6617,N_6781);
or U6996 (N_6996,N_6884,N_6678);
or U6997 (N_6997,N_6867,N_6840);
and U6998 (N_6998,N_6770,N_6882);
nor U6999 (N_6999,N_6856,N_6719);
nand U7000 (N_7000,N_6765,N_6805);
nor U7001 (N_7001,N_6843,N_6763);
xor U7002 (N_7002,N_6766,N_6656);
nor U7003 (N_7003,N_6677,N_6899);
and U7004 (N_7004,N_6890,N_6725);
xor U7005 (N_7005,N_6768,N_6659);
or U7006 (N_7006,N_6809,N_6836);
nand U7007 (N_7007,N_6636,N_6858);
xor U7008 (N_7008,N_6652,N_6853);
nor U7009 (N_7009,N_6751,N_6879);
and U7010 (N_7010,N_6630,N_6876);
nor U7011 (N_7011,N_6825,N_6761);
and U7012 (N_7012,N_6817,N_6861);
nor U7013 (N_7013,N_6749,N_6680);
xor U7014 (N_7014,N_6886,N_6850);
nor U7015 (N_7015,N_6778,N_6609);
nand U7016 (N_7016,N_6846,N_6793);
or U7017 (N_7017,N_6662,N_6771);
and U7018 (N_7018,N_6892,N_6847);
xnor U7019 (N_7019,N_6614,N_6772);
and U7020 (N_7020,N_6786,N_6792);
and U7021 (N_7021,N_6700,N_6799);
nor U7022 (N_7022,N_6816,N_6852);
nand U7023 (N_7023,N_6650,N_6875);
and U7024 (N_7024,N_6668,N_6687);
nand U7025 (N_7025,N_6762,N_6712);
or U7026 (N_7026,N_6887,N_6881);
nand U7027 (N_7027,N_6639,N_6704);
xor U7028 (N_7028,N_6769,N_6706);
and U7029 (N_7029,N_6615,N_6718);
xnor U7030 (N_7030,N_6756,N_6646);
or U7031 (N_7031,N_6834,N_6607);
xor U7032 (N_7032,N_6679,N_6860);
and U7033 (N_7033,N_6740,N_6752);
nand U7034 (N_7034,N_6827,N_6894);
or U7035 (N_7035,N_6683,N_6897);
xor U7036 (N_7036,N_6602,N_6684);
nand U7037 (N_7037,N_6764,N_6758);
or U7038 (N_7038,N_6632,N_6661);
nor U7039 (N_7039,N_6682,N_6742);
and U7040 (N_7040,N_6820,N_6777);
nand U7041 (N_7041,N_6864,N_6653);
xor U7042 (N_7042,N_6822,N_6870);
xnor U7043 (N_7043,N_6797,N_6689);
nor U7044 (N_7044,N_6869,N_6859);
xnor U7045 (N_7045,N_6898,N_6794);
xnor U7046 (N_7046,N_6813,N_6796);
and U7047 (N_7047,N_6675,N_6612);
nor U7048 (N_7048,N_6855,N_6729);
xor U7049 (N_7049,N_6818,N_6690);
xor U7050 (N_7050,N_6733,N_6874);
xnor U7051 (N_7051,N_6600,N_6714);
and U7052 (N_7052,N_6609,N_6890);
or U7053 (N_7053,N_6646,N_6741);
xor U7054 (N_7054,N_6720,N_6821);
nand U7055 (N_7055,N_6742,N_6828);
xor U7056 (N_7056,N_6700,N_6712);
or U7057 (N_7057,N_6750,N_6795);
or U7058 (N_7058,N_6647,N_6804);
or U7059 (N_7059,N_6848,N_6819);
nand U7060 (N_7060,N_6896,N_6893);
and U7061 (N_7061,N_6819,N_6611);
nor U7062 (N_7062,N_6793,N_6666);
and U7063 (N_7063,N_6692,N_6620);
xor U7064 (N_7064,N_6619,N_6832);
nor U7065 (N_7065,N_6624,N_6686);
and U7066 (N_7066,N_6614,N_6663);
nor U7067 (N_7067,N_6680,N_6872);
and U7068 (N_7068,N_6747,N_6863);
xor U7069 (N_7069,N_6889,N_6601);
xor U7070 (N_7070,N_6718,N_6866);
nand U7071 (N_7071,N_6701,N_6676);
or U7072 (N_7072,N_6853,N_6725);
or U7073 (N_7073,N_6762,N_6857);
or U7074 (N_7074,N_6643,N_6750);
nor U7075 (N_7075,N_6822,N_6707);
nor U7076 (N_7076,N_6640,N_6658);
and U7077 (N_7077,N_6805,N_6778);
and U7078 (N_7078,N_6633,N_6817);
nand U7079 (N_7079,N_6829,N_6633);
or U7080 (N_7080,N_6646,N_6879);
or U7081 (N_7081,N_6806,N_6648);
and U7082 (N_7082,N_6782,N_6734);
xnor U7083 (N_7083,N_6739,N_6666);
and U7084 (N_7084,N_6752,N_6697);
nand U7085 (N_7085,N_6638,N_6887);
and U7086 (N_7086,N_6830,N_6765);
or U7087 (N_7087,N_6880,N_6624);
xor U7088 (N_7088,N_6887,N_6842);
nand U7089 (N_7089,N_6693,N_6738);
xor U7090 (N_7090,N_6635,N_6608);
nand U7091 (N_7091,N_6668,N_6665);
xor U7092 (N_7092,N_6812,N_6772);
and U7093 (N_7093,N_6815,N_6622);
nand U7094 (N_7094,N_6785,N_6664);
or U7095 (N_7095,N_6601,N_6631);
xnor U7096 (N_7096,N_6826,N_6837);
nand U7097 (N_7097,N_6876,N_6632);
or U7098 (N_7098,N_6837,N_6891);
xnor U7099 (N_7099,N_6887,N_6773);
and U7100 (N_7100,N_6660,N_6790);
nand U7101 (N_7101,N_6789,N_6693);
nand U7102 (N_7102,N_6698,N_6648);
nand U7103 (N_7103,N_6775,N_6748);
nand U7104 (N_7104,N_6625,N_6624);
or U7105 (N_7105,N_6820,N_6656);
and U7106 (N_7106,N_6697,N_6772);
xor U7107 (N_7107,N_6839,N_6699);
and U7108 (N_7108,N_6873,N_6798);
nand U7109 (N_7109,N_6827,N_6617);
and U7110 (N_7110,N_6606,N_6806);
or U7111 (N_7111,N_6788,N_6851);
xor U7112 (N_7112,N_6888,N_6682);
nand U7113 (N_7113,N_6699,N_6861);
xnor U7114 (N_7114,N_6671,N_6611);
nand U7115 (N_7115,N_6815,N_6776);
nor U7116 (N_7116,N_6865,N_6674);
nor U7117 (N_7117,N_6862,N_6885);
and U7118 (N_7118,N_6612,N_6695);
and U7119 (N_7119,N_6699,N_6850);
xor U7120 (N_7120,N_6680,N_6825);
and U7121 (N_7121,N_6663,N_6811);
nand U7122 (N_7122,N_6793,N_6765);
xor U7123 (N_7123,N_6610,N_6797);
or U7124 (N_7124,N_6685,N_6759);
nor U7125 (N_7125,N_6725,N_6603);
and U7126 (N_7126,N_6823,N_6815);
nor U7127 (N_7127,N_6702,N_6668);
or U7128 (N_7128,N_6617,N_6751);
and U7129 (N_7129,N_6794,N_6695);
nor U7130 (N_7130,N_6688,N_6757);
and U7131 (N_7131,N_6731,N_6759);
or U7132 (N_7132,N_6621,N_6747);
xor U7133 (N_7133,N_6612,N_6829);
and U7134 (N_7134,N_6610,N_6697);
and U7135 (N_7135,N_6646,N_6847);
xnor U7136 (N_7136,N_6852,N_6857);
and U7137 (N_7137,N_6739,N_6750);
nand U7138 (N_7138,N_6707,N_6680);
or U7139 (N_7139,N_6777,N_6794);
nor U7140 (N_7140,N_6732,N_6734);
or U7141 (N_7141,N_6625,N_6700);
or U7142 (N_7142,N_6894,N_6871);
and U7143 (N_7143,N_6802,N_6897);
nor U7144 (N_7144,N_6637,N_6772);
nand U7145 (N_7145,N_6620,N_6707);
or U7146 (N_7146,N_6671,N_6810);
or U7147 (N_7147,N_6818,N_6810);
xor U7148 (N_7148,N_6725,N_6897);
nor U7149 (N_7149,N_6675,N_6621);
nand U7150 (N_7150,N_6839,N_6791);
nor U7151 (N_7151,N_6757,N_6712);
or U7152 (N_7152,N_6879,N_6644);
nor U7153 (N_7153,N_6758,N_6835);
or U7154 (N_7154,N_6899,N_6762);
and U7155 (N_7155,N_6781,N_6702);
nand U7156 (N_7156,N_6729,N_6666);
or U7157 (N_7157,N_6802,N_6668);
nor U7158 (N_7158,N_6856,N_6724);
or U7159 (N_7159,N_6865,N_6718);
and U7160 (N_7160,N_6820,N_6795);
xor U7161 (N_7161,N_6782,N_6880);
or U7162 (N_7162,N_6707,N_6865);
nand U7163 (N_7163,N_6690,N_6657);
or U7164 (N_7164,N_6691,N_6854);
or U7165 (N_7165,N_6674,N_6758);
xor U7166 (N_7166,N_6787,N_6884);
or U7167 (N_7167,N_6793,N_6678);
or U7168 (N_7168,N_6635,N_6835);
nand U7169 (N_7169,N_6603,N_6820);
or U7170 (N_7170,N_6790,N_6641);
nor U7171 (N_7171,N_6840,N_6645);
nor U7172 (N_7172,N_6749,N_6773);
and U7173 (N_7173,N_6787,N_6603);
or U7174 (N_7174,N_6826,N_6705);
nor U7175 (N_7175,N_6821,N_6802);
nand U7176 (N_7176,N_6745,N_6812);
or U7177 (N_7177,N_6844,N_6803);
nor U7178 (N_7178,N_6859,N_6834);
or U7179 (N_7179,N_6720,N_6616);
nor U7180 (N_7180,N_6782,N_6638);
nand U7181 (N_7181,N_6732,N_6847);
xnor U7182 (N_7182,N_6884,N_6710);
and U7183 (N_7183,N_6809,N_6705);
or U7184 (N_7184,N_6785,N_6678);
or U7185 (N_7185,N_6633,N_6707);
nor U7186 (N_7186,N_6873,N_6653);
nand U7187 (N_7187,N_6831,N_6688);
xor U7188 (N_7188,N_6686,N_6681);
xor U7189 (N_7189,N_6741,N_6875);
xnor U7190 (N_7190,N_6846,N_6715);
nand U7191 (N_7191,N_6638,N_6758);
nand U7192 (N_7192,N_6725,N_6623);
xor U7193 (N_7193,N_6662,N_6757);
and U7194 (N_7194,N_6722,N_6841);
nor U7195 (N_7195,N_6741,N_6638);
nand U7196 (N_7196,N_6778,N_6710);
and U7197 (N_7197,N_6889,N_6606);
nor U7198 (N_7198,N_6620,N_6651);
and U7199 (N_7199,N_6791,N_6730);
nand U7200 (N_7200,N_6992,N_6910);
and U7201 (N_7201,N_7106,N_7196);
or U7202 (N_7202,N_6974,N_7095);
or U7203 (N_7203,N_7148,N_7161);
nand U7204 (N_7204,N_6917,N_7039);
nor U7205 (N_7205,N_7042,N_7064);
xnor U7206 (N_7206,N_6970,N_7025);
and U7207 (N_7207,N_7047,N_6997);
nand U7208 (N_7208,N_7040,N_6998);
and U7209 (N_7209,N_6919,N_7140);
nor U7210 (N_7210,N_7084,N_6980);
nor U7211 (N_7211,N_6906,N_7092);
xor U7212 (N_7212,N_6944,N_7043);
xnor U7213 (N_7213,N_7108,N_6966);
and U7214 (N_7214,N_7125,N_7197);
or U7215 (N_7215,N_7158,N_7101);
nand U7216 (N_7216,N_7018,N_7166);
or U7217 (N_7217,N_7147,N_6907);
nor U7218 (N_7218,N_6968,N_7036);
xnor U7219 (N_7219,N_6905,N_7071);
or U7220 (N_7220,N_7055,N_7009);
nand U7221 (N_7221,N_7053,N_7031);
or U7222 (N_7222,N_7184,N_6949);
xnor U7223 (N_7223,N_6911,N_7020);
or U7224 (N_7224,N_7153,N_7017);
xnor U7225 (N_7225,N_7026,N_7127);
and U7226 (N_7226,N_7014,N_6908);
or U7227 (N_7227,N_7165,N_6912);
xor U7228 (N_7228,N_6999,N_6946);
nor U7229 (N_7229,N_7123,N_7183);
and U7230 (N_7230,N_7162,N_6929);
nor U7231 (N_7231,N_7006,N_7087);
and U7232 (N_7232,N_7152,N_6941);
nor U7233 (N_7233,N_7103,N_6916);
nor U7234 (N_7234,N_6952,N_6902);
and U7235 (N_7235,N_7016,N_7062);
nand U7236 (N_7236,N_7021,N_7195);
xnor U7237 (N_7237,N_7027,N_6918);
or U7238 (N_7238,N_6933,N_7137);
nand U7239 (N_7239,N_6950,N_7054);
or U7240 (N_7240,N_6947,N_7120);
nand U7241 (N_7241,N_7116,N_6951);
and U7242 (N_7242,N_7181,N_6954);
nand U7243 (N_7243,N_7034,N_7169);
xor U7244 (N_7244,N_7046,N_7049);
nand U7245 (N_7245,N_7198,N_6971);
nor U7246 (N_7246,N_6931,N_7154);
or U7247 (N_7247,N_7004,N_7105);
and U7248 (N_7248,N_7001,N_7131);
nand U7249 (N_7249,N_7175,N_7012);
nand U7250 (N_7250,N_7061,N_7068);
and U7251 (N_7251,N_7121,N_7080);
xor U7252 (N_7252,N_7044,N_6948);
xnor U7253 (N_7253,N_7079,N_6994);
and U7254 (N_7254,N_7019,N_7011);
nand U7255 (N_7255,N_7122,N_6965);
nand U7256 (N_7256,N_7075,N_7150);
nor U7257 (N_7257,N_6995,N_6961);
nor U7258 (N_7258,N_6983,N_7104);
or U7259 (N_7259,N_7010,N_7167);
and U7260 (N_7260,N_6930,N_7090);
xnor U7261 (N_7261,N_7124,N_7088);
nor U7262 (N_7262,N_7135,N_7155);
nand U7263 (N_7263,N_6923,N_6936);
or U7264 (N_7264,N_7118,N_6981);
nand U7265 (N_7265,N_7005,N_7115);
xor U7266 (N_7266,N_7048,N_6996);
or U7267 (N_7267,N_7179,N_7182);
and U7268 (N_7268,N_6925,N_7096);
and U7269 (N_7269,N_7111,N_7093);
xnor U7270 (N_7270,N_7045,N_7149);
xnor U7271 (N_7271,N_7141,N_7022);
nor U7272 (N_7272,N_7091,N_7156);
nand U7273 (N_7273,N_7003,N_7085);
xor U7274 (N_7274,N_6921,N_7015);
nand U7275 (N_7275,N_6987,N_7109);
and U7276 (N_7276,N_7157,N_6937);
and U7277 (N_7277,N_7177,N_7063);
xnor U7278 (N_7278,N_7142,N_7083);
nor U7279 (N_7279,N_6920,N_7190);
or U7280 (N_7280,N_7024,N_7082);
nand U7281 (N_7281,N_7151,N_6964);
nor U7282 (N_7282,N_7180,N_7078);
or U7283 (N_7283,N_7089,N_7112);
xnor U7284 (N_7284,N_7186,N_7066);
nor U7285 (N_7285,N_7086,N_6935);
nor U7286 (N_7286,N_7037,N_7099);
nor U7287 (N_7287,N_6953,N_7173);
and U7288 (N_7288,N_7192,N_7008);
or U7289 (N_7289,N_6962,N_7132);
nor U7290 (N_7290,N_6969,N_7065);
nor U7291 (N_7291,N_6928,N_7168);
nand U7292 (N_7292,N_7129,N_7038);
or U7293 (N_7293,N_7117,N_7160);
xor U7294 (N_7294,N_6956,N_6982);
nand U7295 (N_7295,N_7189,N_6955);
or U7296 (N_7296,N_7143,N_7050);
and U7297 (N_7297,N_6901,N_7171);
nor U7298 (N_7298,N_7035,N_7072);
xor U7299 (N_7299,N_7114,N_7119);
xor U7300 (N_7300,N_7130,N_6963);
or U7301 (N_7301,N_6915,N_6986);
and U7302 (N_7302,N_7029,N_6957);
xor U7303 (N_7303,N_7194,N_7128);
xor U7304 (N_7304,N_6940,N_7159);
or U7305 (N_7305,N_6993,N_7199);
xnor U7306 (N_7306,N_7052,N_7172);
or U7307 (N_7307,N_6958,N_7176);
and U7308 (N_7308,N_7033,N_6914);
or U7309 (N_7309,N_7013,N_6984);
and U7310 (N_7310,N_7056,N_7163);
or U7311 (N_7311,N_6990,N_6991);
nor U7312 (N_7312,N_6959,N_7170);
and U7313 (N_7313,N_7102,N_7144);
and U7314 (N_7314,N_7188,N_7145);
nor U7315 (N_7315,N_6939,N_6900);
nor U7316 (N_7316,N_6960,N_6967);
or U7317 (N_7317,N_7059,N_7094);
xor U7318 (N_7318,N_7193,N_6978);
xnor U7319 (N_7319,N_7076,N_6985);
and U7320 (N_7320,N_6973,N_7070);
xor U7321 (N_7321,N_7057,N_7133);
xor U7322 (N_7322,N_7178,N_7074);
nand U7323 (N_7323,N_6988,N_6932);
and U7324 (N_7324,N_7051,N_7028);
xnor U7325 (N_7325,N_6989,N_7041);
nor U7326 (N_7326,N_7107,N_6924);
nand U7327 (N_7327,N_7073,N_6904);
nand U7328 (N_7328,N_6927,N_6903);
and U7329 (N_7329,N_7134,N_6942);
or U7330 (N_7330,N_7058,N_7138);
xnor U7331 (N_7331,N_7023,N_7185);
or U7332 (N_7332,N_6979,N_7126);
or U7333 (N_7333,N_6926,N_6945);
and U7334 (N_7334,N_6934,N_7007);
nor U7335 (N_7335,N_7069,N_6977);
nand U7336 (N_7336,N_7187,N_6976);
nand U7337 (N_7337,N_7000,N_7164);
and U7338 (N_7338,N_7146,N_7191);
nand U7339 (N_7339,N_7030,N_7081);
xnor U7340 (N_7340,N_7097,N_6913);
nand U7341 (N_7341,N_6922,N_6972);
or U7342 (N_7342,N_7098,N_7110);
or U7343 (N_7343,N_7032,N_7060);
xor U7344 (N_7344,N_7077,N_6943);
xor U7345 (N_7345,N_7100,N_7113);
xnor U7346 (N_7346,N_7002,N_6938);
or U7347 (N_7347,N_7136,N_7174);
or U7348 (N_7348,N_6975,N_7067);
xnor U7349 (N_7349,N_7139,N_6909);
and U7350 (N_7350,N_7193,N_7094);
nor U7351 (N_7351,N_7165,N_7020);
nand U7352 (N_7352,N_7037,N_6922);
nor U7353 (N_7353,N_6970,N_6977);
nand U7354 (N_7354,N_6957,N_6960);
or U7355 (N_7355,N_7122,N_7096);
and U7356 (N_7356,N_6984,N_7083);
and U7357 (N_7357,N_7065,N_6924);
nor U7358 (N_7358,N_7055,N_7038);
nor U7359 (N_7359,N_6979,N_7055);
xor U7360 (N_7360,N_7146,N_7108);
xor U7361 (N_7361,N_7036,N_7127);
or U7362 (N_7362,N_6960,N_7149);
nor U7363 (N_7363,N_7145,N_7063);
or U7364 (N_7364,N_6913,N_7079);
and U7365 (N_7365,N_7015,N_6904);
xnor U7366 (N_7366,N_6975,N_7048);
or U7367 (N_7367,N_7038,N_7067);
xor U7368 (N_7368,N_7018,N_7007);
and U7369 (N_7369,N_6951,N_6969);
nand U7370 (N_7370,N_6916,N_7004);
nand U7371 (N_7371,N_6979,N_7074);
nor U7372 (N_7372,N_7094,N_7196);
nand U7373 (N_7373,N_7079,N_7022);
nand U7374 (N_7374,N_7017,N_7092);
or U7375 (N_7375,N_6950,N_7185);
nand U7376 (N_7376,N_7166,N_6959);
and U7377 (N_7377,N_6920,N_7106);
nand U7378 (N_7378,N_6906,N_7002);
nand U7379 (N_7379,N_6994,N_6986);
xor U7380 (N_7380,N_7071,N_7051);
nand U7381 (N_7381,N_6908,N_7133);
and U7382 (N_7382,N_6965,N_6985);
nor U7383 (N_7383,N_7055,N_7137);
and U7384 (N_7384,N_7126,N_6913);
nand U7385 (N_7385,N_7093,N_6966);
and U7386 (N_7386,N_7180,N_6937);
or U7387 (N_7387,N_7117,N_7170);
nand U7388 (N_7388,N_7198,N_7172);
and U7389 (N_7389,N_7120,N_6933);
nand U7390 (N_7390,N_7018,N_6915);
or U7391 (N_7391,N_7044,N_7164);
xor U7392 (N_7392,N_7067,N_7195);
and U7393 (N_7393,N_6950,N_7041);
nand U7394 (N_7394,N_7199,N_7014);
nor U7395 (N_7395,N_6991,N_7137);
nor U7396 (N_7396,N_6918,N_7118);
or U7397 (N_7397,N_7120,N_6916);
xor U7398 (N_7398,N_7176,N_7108);
nor U7399 (N_7399,N_7097,N_6935);
xor U7400 (N_7400,N_6900,N_6948);
or U7401 (N_7401,N_7069,N_7027);
or U7402 (N_7402,N_7051,N_7099);
or U7403 (N_7403,N_6984,N_6949);
nor U7404 (N_7404,N_7129,N_7099);
or U7405 (N_7405,N_7109,N_6909);
and U7406 (N_7406,N_6959,N_7123);
nand U7407 (N_7407,N_7195,N_7199);
and U7408 (N_7408,N_6983,N_7130);
nand U7409 (N_7409,N_6912,N_6971);
and U7410 (N_7410,N_7071,N_6956);
xnor U7411 (N_7411,N_6931,N_7125);
and U7412 (N_7412,N_6991,N_7159);
nor U7413 (N_7413,N_7144,N_6947);
and U7414 (N_7414,N_6916,N_7171);
or U7415 (N_7415,N_6904,N_6969);
nor U7416 (N_7416,N_7196,N_7046);
and U7417 (N_7417,N_7136,N_7105);
and U7418 (N_7418,N_7155,N_6983);
xnor U7419 (N_7419,N_6958,N_6980);
xnor U7420 (N_7420,N_7012,N_7070);
xnor U7421 (N_7421,N_7055,N_6971);
nor U7422 (N_7422,N_7106,N_7131);
nand U7423 (N_7423,N_6988,N_7010);
and U7424 (N_7424,N_7051,N_7112);
and U7425 (N_7425,N_6982,N_7142);
and U7426 (N_7426,N_7096,N_6913);
nor U7427 (N_7427,N_6959,N_6971);
or U7428 (N_7428,N_7007,N_7072);
nand U7429 (N_7429,N_6937,N_7044);
xnor U7430 (N_7430,N_7062,N_7075);
nor U7431 (N_7431,N_6924,N_7159);
and U7432 (N_7432,N_7136,N_7069);
or U7433 (N_7433,N_7015,N_7026);
xnor U7434 (N_7434,N_7065,N_7035);
nand U7435 (N_7435,N_7052,N_7016);
nand U7436 (N_7436,N_7027,N_7116);
nand U7437 (N_7437,N_7029,N_7036);
xnor U7438 (N_7438,N_7075,N_7035);
nor U7439 (N_7439,N_7111,N_6964);
nand U7440 (N_7440,N_6917,N_7006);
xor U7441 (N_7441,N_7187,N_6955);
xor U7442 (N_7442,N_7177,N_7010);
nand U7443 (N_7443,N_7014,N_7119);
xnor U7444 (N_7444,N_6906,N_7147);
and U7445 (N_7445,N_7128,N_7146);
and U7446 (N_7446,N_6940,N_7116);
nand U7447 (N_7447,N_6952,N_6997);
xor U7448 (N_7448,N_7196,N_7034);
nand U7449 (N_7449,N_6949,N_7132);
nand U7450 (N_7450,N_7034,N_7195);
and U7451 (N_7451,N_6905,N_7163);
and U7452 (N_7452,N_7121,N_6968);
nand U7453 (N_7453,N_7059,N_7010);
or U7454 (N_7454,N_6944,N_7057);
xnor U7455 (N_7455,N_6969,N_7097);
and U7456 (N_7456,N_7052,N_7198);
nand U7457 (N_7457,N_7020,N_7088);
nand U7458 (N_7458,N_6914,N_7010);
or U7459 (N_7459,N_7126,N_6968);
xnor U7460 (N_7460,N_7000,N_6953);
nor U7461 (N_7461,N_7159,N_6919);
xnor U7462 (N_7462,N_6910,N_7028);
nor U7463 (N_7463,N_7002,N_6979);
xnor U7464 (N_7464,N_7125,N_7053);
nor U7465 (N_7465,N_7176,N_6926);
or U7466 (N_7466,N_6930,N_6934);
or U7467 (N_7467,N_6922,N_7005);
xnor U7468 (N_7468,N_7168,N_6958);
and U7469 (N_7469,N_7008,N_7058);
and U7470 (N_7470,N_7198,N_6952);
or U7471 (N_7471,N_7111,N_6943);
xor U7472 (N_7472,N_6901,N_6983);
or U7473 (N_7473,N_6975,N_7183);
nand U7474 (N_7474,N_7109,N_7137);
and U7475 (N_7475,N_6956,N_6950);
and U7476 (N_7476,N_6934,N_7119);
nand U7477 (N_7477,N_7005,N_7116);
nor U7478 (N_7478,N_7082,N_7121);
and U7479 (N_7479,N_7110,N_7152);
nor U7480 (N_7480,N_7127,N_7142);
nand U7481 (N_7481,N_6901,N_7030);
xor U7482 (N_7482,N_7043,N_7180);
nand U7483 (N_7483,N_7142,N_7113);
xnor U7484 (N_7484,N_7083,N_6964);
nor U7485 (N_7485,N_6928,N_6946);
nand U7486 (N_7486,N_7191,N_7000);
nor U7487 (N_7487,N_7034,N_7191);
nor U7488 (N_7488,N_7115,N_7086);
or U7489 (N_7489,N_6975,N_7063);
nand U7490 (N_7490,N_7102,N_7046);
nand U7491 (N_7491,N_7199,N_7186);
and U7492 (N_7492,N_7052,N_7183);
and U7493 (N_7493,N_7079,N_7047);
or U7494 (N_7494,N_7013,N_7149);
nand U7495 (N_7495,N_7044,N_6970);
or U7496 (N_7496,N_7061,N_7144);
nand U7497 (N_7497,N_7193,N_6977);
nor U7498 (N_7498,N_7001,N_7063);
xnor U7499 (N_7499,N_7113,N_7009);
xor U7500 (N_7500,N_7332,N_7406);
nor U7501 (N_7501,N_7261,N_7490);
xor U7502 (N_7502,N_7316,N_7343);
xor U7503 (N_7503,N_7437,N_7205);
nor U7504 (N_7504,N_7268,N_7452);
nor U7505 (N_7505,N_7424,N_7213);
and U7506 (N_7506,N_7459,N_7248);
and U7507 (N_7507,N_7445,N_7203);
nand U7508 (N_7508,N_7410,N_7481);
and U7509 (N_7509,N_7357,N_7280);
nor U7510 (N_7510,N_7216,N_7446);
xnor U7511 (N_7511,N_7463,N_7394);
xor U7512 (N_7512,N_7389,N_7412);
xnor U7513 (N_7513,N_7351,N_7432);
or U7514 (N_7514,N_7498,N_7326);
or U7515 (N_7515,N_7226,N_7384);
nand U7516 (N_7516,N_7461,N_7386);
nor U7517 (N_7517,N_7322,N_7349);
nor U7518 (N_7518,N_7355,N_7473);
or U7519 (N_7519,N_7240,N_7257);
nand U7520 (N_7520,N_7364,N_7373);
or U7521 (N_7521,N_7362,N_7426);
nand U7522 (N_7522,N_7247,N_7238);
nor U7523 (N_7523,N_7487,N_7414);
xor U7524 (N_7524,N_7296,N_7360);
nand U7525 (N_7525,N_7344,N_7251);
nor U7526 (N_7526,N_7223,N_7417);
nand U7527 (N_7527,N_7407,N_7214);
nand U7528 (N_7528,N_7273,N_7259);
nand U7529 (N_7529,N_7413,N_7207);
nor U7530 (N_7530,N_7376,N_7474);
xor U7531 (N_7531,N_7350,N_7381);
or U7532 (N_7532,N_7225,N_7365);
nor U7533 (N_7533,N_7244,N_7329);
or U7534 (N_7534,N_7428,N_7265);
or U7535 (N_7535,N_7366,N_7287);
nand U7536 (N_7536,N_7380,N_7224);
nand U7537 (N_7537,N_7334,N_7438);
or U7538 (N_7538,N_7267,N_7399);
xor U7539 (N_7539,N_7484,N_7402);
and U7540 (N_7540,N_7263,N_7305);
or U7541 (N_7541,N_7297,N_7489);
or U7542 (N_7542,N_7482,N_7204);
or U7543 (N_7543,N_7272,N_7450);
or U7544 (N_7544,N_7290,N_7411);
nand U7545 (N_7545,N_7444,N_7246);
and U7546 (N_7546,N_7234,N_7488);
nand U7547 (N_7547,N_7243,N_7395);
and U7548 (N_7548,N_7393,N_7369);
and U7549 (N_7549,N_7420,N_7492);
xnor U7550 (N_7550,N_7325,N_7338);
or U7551 (N_7551,N_7404,N_7464);
nor U7552 (N_7552,N_7242,N_7200);
nor U7553 (N_7553,N_7422,N_7477);
nor U7554 (N_7554,N_7397,N_7258);
xnor U7555 (N_7555,N_7491,N_7310);
nor U7556 (N_7556,N_7237,N_7390);
xnor U7557 (N_7557,N_7330,N_7283);
and U7558 (N_7558,N_7289,N_7228);
nor U7559 (N_7559,N_7494,N_7304);
xnor U7560 (N_7560,N_7496,N_7254);
nand U7561 (N_7561,N_7210,N_7448);
and U7562 (N_7562,N_7279,N_7443);
or U7563 (N_7563,N_7308,N_7398);
xor U7564 (N_7564,N_7486,N_7231);
nand U7565 (N_7565,N_7229,N_7485);
and U7566 (N_7566,N_7453,N_7433);
or U7567 (N_7567,N_7460,N_7337);
and U7568 (N_7568,N_7206,N_7359);
nand U7569 (N_7569,N_7233,N_7209);
or U7570 (N_7570,N_7201,N_7430);
nand U7571 (N_7571,N_7408,N_7314);
nor U7572 (N_7572,N_7429,N_7219);
nand U7573 (N_7573,N_7375,N_7468);
xnor U7574 (N_7574,N_7348,N_7286);
and U7575 (N_7575,N_7275,N_7483);
or U7576 (N_7576,N_7327,N_7335);
or U7577 (N_7577,N_7409,N_7449);
and U7578 (N_7578,N_7467,N_7479);
nand U7579 (N_7579,N_7253,N_7227);
and U7580 (N_7580,N_7379,N_7340);
xnor U7581 (N_7581,N_7300,N_7385);
nor U7582 (N_7582,N_7454,N_7425);
nor U7583 (N_7583,N_7271,N_7215);
xnor U7584 (N_7584,N_7220,N_7469);
nor U7585 (N_7585,N_7298,N_7260);
xor U7586 (N_7586,N_7321,N_7456);
or U7587 (N_7587,N_7388,N_7442);
nor U7588 (N_7588,N_7371,N_7288);
nor U7589 (N_7589,N_7396,N_7281);
or U7590 (N_7590,N_7249,N_7478);
nor U7591 (N_7591,N_7235,N_7358);
and U7592 (N_7592,N_7370,N_7236);
and U7593 (N_7593,N_7341,N_7306);
nor U7594 (N_7594,N_7339,N_7311);
xor U7595 (N_7595,N_7317,N_7245);
nand U7596 (N_7596,N_7319,N_7202);
xnor U7597 (N_7597,N_7400,N_7284);
nor U7598 (N_7598,N_7212,N_7301);
and U7599 (N_7599,N_7367,N_7434);
nor U7600 (N_7600,N_7354,N_7217);
and U7601 (N_7601,N_7345,N_7392);
xnor U7602 (N_7602,N_7313,N_7466);
nand U7603 (N_7603,N_7269,N_7277);
xnor U7604 (N_7604,N_7493,N_7285);
nor U7605 (N_7605,N_7328,N_7232);
and U7606 (N_7606,N_7480,N_7346);
and U7607 (N_7607,N_7457,N_7256);
and U7608 (N_7608,N_7415,N_7418);
and U7609 (N_7609,N_7472,N_7447);
and U7610 (N_7610,N_7250,N_7318);
xnor U7611 (N_7611,N_7405,N_7382);
and U7612 (N_7612,N_7458,N_7419);
and U7613 (N_7613,N_7372,N_7374);
nand U7614 (N_7614,N_7208,N_7470);
xor U7615 (N_7615,N_7387,N_7497);
or U7616 (N_7616,N_7293,N_7211);
and U7617 (N_7617,N_7423,N_7476);
xor U7618 (N_7618,N_7307,N_7391);
xor U7619 (N_7619,N_7299,N_7241);
and U7620 (N_7620,N_7222,N_7383);
nor U7621 (N_7621,N_7309,N_7302);
and U7622 (N_7622,N_7427,N_7441);
xnor U7623 (N_7623,N_7295,N_7439);
xor U7624 (N_7624,N_7462,N_7218);
or U7625 (N_7625,N_7471,N_7352);
nor U7626 (N_7626,N_7377,N_7292);
or U7627 (N_7627,N_7331,N_7303);
nor U7628 (N_7628,N_7368,N_7270);
or U7629 (N_7629,N_7440,N_7431);
nand U7630 (N_7630,N_7255,N_7221);
and U7631 (N_7631,N_7291,N_7323);
nor U7632 (N_7632,N_7276,N_7436);
xnor U7633 (N_7633,N_7347,N_7336);
and U7634 (N_7634,N_7239,N_7451);
nor U7635 (N_7635,N_7499,N_7421);
and U7636 (N_7636,N_7294,N_7361);
nand U7637 (N_7637,N_7435,N_7356);
xor U7638 (N_7638,N_7252,N_7353);
or U7639 (N_7639,N_7320,N_7278);
xor U7640 (N_7640,N_7315,N_7324);
nor U7641 (N_7641,N_7378,N_7465);
nand U7642 (N_7642,N_7495,N_7262);
nor U7643 (N_7643,N_7403,N_7312);
xor U7644 (N_7644,N_7230,N_7274);
nand U7645 (N_7645,N_7333,N_7401);
and U7646 (N_7646,N_7475,N_7264);
xnor U7647 (N_7647,N_7416,N_7266);
or U7648 (N_7648,N_7455,N_7282);
xor U7649 (N_7649,N_7342,N_7363);
or U7650 (N_7650,N_7218,N_7251);
xnor U7651 (N_7651,N_7395,N_7203);
nor U7652 (N_7652,N_7485,N_7407);
or U7653 (N_7653,N_7361,N_7453);
xor U7654 (N_7654,N_7488,N_7428);
xor U7655 (N_7655,N_7472,N_7334);
nor U7656 (N_7656,N_7488,N_7281);
or U7657 (N_7657,N_7440,N_7379);
nand U7658 (N_7658,N_7369,N_7487);
nor U7659 (N_7659,N_7476,N_7292);
nor U7660 (N_7660,N_7314,N_7252);
and U7661 (N_7661,N_7313,N_7328);
and U7662 (N_7662,N_7291,N_7454);
xor U7663 (N_7663,N_7215,N_7281);
nor U7664 (N_7664,N_7258,N_7242);
and U7665 (N_7665,N_7345,N_7325);
xnor U7666 (N_7666,N_7460,N_7255);
and U7667 (N_7667,N_7333,N_7279);
xnor U7668 (N_7668,N_7356,N_7261);
nor U7669 (N_7669,N_7407,N_7433);
nor U7670 (N_7670,N_7452,N_7305);
nor U7671 (N_7671,N_7476,N_7429);
nor U7672 (N_7672,N_7207,N_7480);
or U7673 (N_7673,N_7233,N_7495);
nand U7674 (N_7674,N_7266,N_7337);
and U7675 (N_7675,N_7446,N_7480);
or U7676 (N_7676,N_7431,N_7353);
or U7677 (N_7677,N_7290,N_7472);
xnor U7678 (N_7678,N_7440,N_7302);
nor U7679 (N_7679,N_7263,N_7439);
xor U7680 (N_7680,N_7275,N_7496);
or U7681 (N_7681,N_7451,N_7395);
nor U7682 (N_7682,N_7368,N_7328);
or U7683 (N_7683,N_7453,N_7490);
nor U7684 (N_7684,N_7238,N_7405);
nand U7685 (N_7685,N_7327,N_7390);
xor U7686 (N_7686,N_7499,N_7410);
xor U7687 (N_7687,N_7355,N_7361);
nor U7688 (N_7688,N_7358,N_7280);
nor U7689 (N_7689,N_7274,N_7353);
nor U7690 (N_7690,N_7221,N_7274);
xor U7691 (N_7691,N_7259,N_7209);
nand U7692 (N_7692,N_7392,N_7486);
xor U7693 (N_7693,N_7284,N_7331);
xor U7694 (N_7694,N_7478,N_7364);
xor U7695 (N_7695,N_7492,N_7237);
nor U7696 (N_7696,N_7414,N_7488);
and U7697 (N_7697,N_7338,N_7244);
and U7698 (N_7698,N_7377,N_7432);
xor U7699 (N_7699,N_7254,N_7473);
and U7700 (N_7700,N_7420,N_7391);
xnor U7701 (N_7701,N_7413,N_7296);
nand U7702 (N_7702,N_7233,N_7299);
or U7703 (N_7703,N_7248,N_7220);
nand U7704 (N_7704,N_7333,N_7395);
or U7705 (N_7705,N_7468,N_7382);
xnor U7706 (N_7706,N_7207,N_7237);
and U7707 (N_7707,N_7355,N_7488);
xor U7708 (N_7708,N_7424,N_7267);
nor U7709 (N_7709,N_7299,N_7335);
nand U7710 (N_7710,N_7352,N_7351);
xnor U7711 (N_7711,N_7363,N_7241);
and U7712 (N_7712,N_7293,N_7495);
and U7713 (N_7713,N_7443,N_7442);
and U7714 (N_7714,N_7399,N_7438);
xor U7715 (N_7715,N_7218,N_7222);
or U7716 (N_7716,N_7216,N_7204);
and U7717 (N_7717,N_7200,N_7492);
xnor U7718 (N_7718,N_7287,N_7437);
and U7719 (N_7719,N_7498,N_7258);
xor U7720 (N_7720,N_7223,N_7443);
and U7721 (N_7721,N_7219,N_7303);
nand U7722 (N_7722,N_7262,N_7486);
and U7723 (N_7723,N_7313,N_7298);
xor U7724 (N_7724,N_7258,N_7225);
nand U7725 (N_7725,N_7390,N_7213);
xnor U7726 (N_7726,N_7443,N_7419);
nand U7727 (N_7727,N_7488,N_7339);
nor U7728 (N_7728,N_7350,N_7420);
xnor U7729 (N_7729,N_7478,N_7243);
and U7730 (N_7730,N_7289,N_7247);
nor U7731 (N_7731,N_7212,N_7281);
nor U7732 (N_7732,N_7267,N_7367);
nor U7733 (N_7733,N_7435,N_7480);
xor U7734 (N_7734,N_7415,N_7392);
nor U7735 (N_7735,N_7400,N_7406);
or U7736 (N_7736,N_7234,N_7260);
nor U7737 (N_7737,N_7227,N_7327);
xnor U7738 (N_7738,N_7452,N_7351);
nand U7739 (N_7739,N_7453,N_7471);
nand U7740 (N_7740,N_7287,N_7466);
xor U7741 (N_7741,N_7437,N_7485);
or U7742 (N_7742,N_7476,N_7303);
or U7743 (N_7743,N_7316,N_7390);
and U7744 (N_7744,N_7430,N_7420);
or U7745 (N_7745,N_7221,N_7389);
nor U7746 (N_7746,N_7379,N_7427);
nand U7747 (N_7747,N_7384,N_7283);
or U7748 (N_7748,N_7267,N_7249);
or U7749 (N_7749,N_7260,N_7327);
xnor U7750 (N_7750,N_7351,N_7202);
and U7751 (N_7751,N_7373,N_7421);
nor U7752 (N_7752,N_7365,N_7209);
xor U7753 (N_7753,N_7264,N_7344);
nand U7754 (N_7754,N_7362,N_7301);
nand U7755 (N_7755,N_7379,N_7473);
or U7756 (N_7756,N_7453,N_7301);
or U7757 (N_7757,N_7327,N_7429);
and U7758 (N_7758,N_7337,N_7226);
nor U7759 (N_7759,N_7327,N_7463);
or U7760 (N_7760,N_7399,N_7306);
nand U7761 (N_7761,N_7408,N_7343);
and U7762 (N_7762,N_7417,N_7255);
and U7763 (N_7763,N_7313,N_7327);
nand U7764 (N_7764,N_7218,N_7472);
nor U7765 (N_7765,N_7454,N_7241);
nor U7766 (N_7766,N_7443,N_7434);
nand U7767 (N_7767,N_7360,N_7319);
xor U7768 (N_7768,N_7270,N_7249);
and U7769 (N_7769,N_7290,N_7237);
and U7770 (N_7770,N_7357,N_7375);
xnor U7771 (N_7771,N_7361,N_7482);
and U7772 (N_7772,N_7223,N_7268);
or U7773 (N_7773,N_7286,N_7260);
nand U7774 (N_7774,N_7428,N_7381);
nor U7775 (N_7775,N_7318,N_7372);
or U7776 (N_7776,N_7366,N_7479);
nand U7777 (N_7777,N_7406,N_7386);
or U7778 (N_7778,N_7481,N_7325);
nand U7779 (N_7779,N_7313,N_7465);
nand U7780 (N_7780,N_7448,N_7364);
nor U7781 (N_7781,N_7475,N_7447);
or U7782 (N_7782,N_7219,N_7263);
nor U7783 (N_7783,N_7429,N_7399);
nand U7784 (N_7784,N_7454,N_7224);
nand U7785 (N_7785,N_7388,N_7308);
xnor U7786 (N_7786,N_7370,N_7460);
or U7787 (N_7787,N_7477,N_7269);
nand U7788 (N_7788,N_7368,N_7263);
and U7789 (N_7789,N_7372,N_7379);
and U7790 (N_7790,N_7446,N_7351);
nor U7791 (N_7791,N_7370,N_7485);
or U7792 (N_7792,N_7305,N_7310);
or U7793 (N_7793,N_7231,N_7446);
or U7794 (N_7794,N_7320,N_7349);
or U7795 (N_7795,N_7295,N_7319);
nand U7796 (N_7796,N_7270,N_7473);
nor U7797 (N_7797,N_7257,N_7398);
and U7798 (N_7798,N_7312,N_7330);
nand U7799 (N_7799,N_7428,N_7390);
nand U7800 (N_7800,N_7642,N_7557);
and U7801 (N_7801,N_7524,N_7713);
xnor U7802 (N_7802,N_7781,N_7652);
nor U7803 (N_7803,N_7640,N_7653);
nand U7804 (N_7804,N_7687,N_7747);
nand U7805 (N_7805,N_7596,N_7796);
nand U7806 (N_7806,N_7750,N_7778);
and U7807 (N_7807,N_7589,N_7725);
nor U7808 (N_7808,N_7583,N_7741);
xor U7809 (N_7809,N_7537,N_7768);
nor U7810 (N_7810,N_7686,N_7798);
nand U7811 (N_7811,N_7777,N_7516);
nand U7812 (N_7812,N_7716,N_7606);
or U7813 (N_7813,N_7502,N_7654);
and U7814 (N_7814,N_7613,N_7793);
and U7815 (N_7815,N_7564,N_7795);
or U7816 (N_7816,N_7761,N_7568);
or U7817 (N_7817,N_7505,N_7539);
and U7818 (N_7818,N_7544,N_7678);
nor U7819 (N_7819,N_7555,N_7666);
xor U7820 (N_7820,N_7649,N_7522);
xnor U7821 (N_7821,N_7710,N_7753);
or U7822 (N_7822,N_7657,N_7594);
nand U7823 (N_7823,N_7540,N_7500);
xnor U7824 (N_7824,N_7785,N_7592);
xnor U7825 (N_7825,N_7569,N_7791);
xnor U7826 (N_7826,N_7633,N_7685);
xor U7827 (N_7827,N_7681,N_7530);
xor U7828 (N_7828,N_7717,N_7617);
and U7829 (N_7829,N_7578,N_7663);
or U7830 (N_7830,N_7698,N_7584);
nand U7831 (N_7831,N_7621,N_7514);
or U7832 (N_7832,N_7748,N_7743);
nor U7833 (N_7833,N_7734,N_7581);
or U7834 (N_7834,N_7675,N_7655);
xnor U7835 (N_7835,N_7535,N_7672);
xnor U7836 (N_7836,N_7566,N_7570);
or U7837 (N_7837,N_7546,N_7545);
xor U7838 (N_7838,N_7595,N_7727);
xnor U7839 (N_7839,N_7776,N_7782);
and U7840 (N_7840,N_7549,N_7771);
xor U7841 (N_7841,N_7508,N_7627);
nor U7842 (N_7842,N_7588,N_7562);
or U7843 (N_7843,N_7533,N_7561);
nand U7844 (N_7844,N_7553,N_7680);
nand U7845 (N_7845,N_7651,N_7630);
nand U7846 (N_7846,N_7575,N_7550);
or U7847 (N_7847,N_7611,N_7673);
and U7848 (N_7848,N_7792,N_7664);
or U7849 (N_7849,N_7737,N_7740);
nand U7850 (N_7850,N_7629,N_7697);
nand U7851 (N_7851,N_7523,N_7679);
and U7852 (N_7852,N_7758,N_7705);
and U7853 (N_7853,N_7756,N_7631);
xor U7854 (N_7854,N_7577,N_7552);
and U7855 (N_7855,N_7724,N_7751);
nor U7856 (N_7856,N_7789,N_7572);
nand U7857 (N_7857,N_7775,N_7706);
and U7858 (N_7858,N_7536,N_7610);
nand U7859 (N_7859,N_7718,N_7542);
xor U7860 (N_7860,N_7684,N_7723);
nor U7861 (N_7861,N_7767,N_7504);
xor U7862 (N_7862,N_7731,N_7515);
and U7863 (N_7863,N_7677,N_7576);
and U7864 (N_7864,N_7556,N_7721);
nand U7865 (N_7865,N_7625,N_7607);
nor U7866 (N_7866,N_7587,N_7511);
nor U7867 (N_7867,N_7643,N_7788);
nor U7868 (N_7868,N_7551,N_7567);
or U7869 (N_7869,N_7730,N_7670);
or U7870 (N_7870,N_7528,N_7790);
nand U7871 (N_7871,N_7695,N_7582);
nand U7872 (N_7872,N_7779,N_7512);
or U7873 (N_7873,N_7614,N_7650);
nand U7874 (N_7874,N_7591,N_7676);
and U7875 (N_7875,N_7637,N_7531);
or U7876 (N_7876,N_7719,N_7736);
xor U7877 (N_7877,N_7527,N_7770);
nand U7878 (N_7878,N_7593,N_7605);
or U7879 (N_7879,N_7780,N_7704);
nand U7880 (N_7880,N_7692,N_7754);
nand U7881 (N_7881,N_7688,N_7709);
xnor U7882 (N_7882,N_7707,N_7525);
or U7883 (N_7883,N_7714,N_7752);
nand U7884 (N_7884,N_7547,N_7619);
xnor U7885 (N_7885,N_7674,N_7520);
or U7886 (N_7886,N_7759,N_7700);
xnor U7887 (N_7887,N_7501,N_7656);
xnor U7888 (N_7888,N_7636,N_7609);
xnor U7889 (N_7889,N_7558,N_7660);
and U7890 (N_7890,N_7510,N_7765);
and U7891 (N_7891,N_7634,N_7598);
or U7892 (N_7892,N_7784,N_7521);
xor U7893 (N_7893,N_7541,N_7799);
or U7894 (N_7894,N_7526,N_7711);
nand U7895 (N_7895,N_7623,N_7665);
or U7896 (N_7896,N_7755,N_7513);
nand U7897 (N_7897,N_7559,N_7735);
xor U7898 (N_7898,N_7694,N_7565);
or U7899 (N_7899,N_7738,N_7733);
or U7900 (N_7900,N_7794,N_7662);
nand U7901 (N_7901,N_7646,N_7715);
and U7902 (N_7902,N_7626,N_7543);
nand U7903 (N_7903,N_7638,N_7766);
nand U7904 (N_7904,N_7615,N_7658);
or U7905 (N_7905,N_7762,N_7519);
or U7906 (N_7906,N_7554,N_7722);
nand U7907 (N_7907,N_7534,N_7529);
xnor U7908 (N_7908,N_7693,N_7600);
nor U7909 (N_7909,N_7708,N_7571);
and U7910 (N_7910,N_7538,N_7602);
nor U7911 (N_7911,N_7639,N_7760);
nand U7912 (N_7912,N_7671,N_7742);
nor U7913 (N_7913,N_7732,N_7597);
nor U7914 (N_7914,N_7560,N_7509);
nor U7915 (N_7915,N_7635,N_7618);
nor U7916 (N_7916,N_7548,N_7746);
and U7917 (N_7917,N_7659,N_7506);
nand U7918 (N_7918,N_7667,N_7763);
xnor U7919 (N_7919,N_7644,N_7616);
xor U7920 (N_7920,N_7749,N_7797);
nor U7921 (N_7921,N_7507,N_7601);
and U7922 (N_7922,N_7787,N_7590);
and U7923 (N_7923,N_7699,N_7712);
nand U7924 (N_7924,N_7608,N_7628);
xor U7925 (N_7925,N_7757,N_7691);
nand U7926 (N_7926,N_7586,N_7774);
nor U7927 (N_7927,N_7585,N_7701);
xor U7928 (N_7928,N_7517,N_7683);
xor U7929 (N_7929,N_7620,N_7703);
xor U7930 (N_7930,N_7745,N_7573);
or U7931 (N_7931,N_7744,N_7668);
nor U7932 (N_7932,N_7624,N_7574);
xnor U7933 (N_7933,N_7690,N_7612);
xor U7934 (N_7934,N_7632,N_7689);
nor U7935 (N_7935,N_7518,N_7503);
xnor U7936 (N_7936,N_7661,N_7702);
and U7937 (N_7937,N_7764,N_7603);
xnor U7938 (N_7938,N_7647,N_7648);
and U7939 (N_7939,N_7739,N_7696);
or U7940 (N_7940,N_7783,N_7579);
and U7941 (N_7941,N_7786,N_7773);
xnor U7942 (N_7942,N_7599,N_7720);
and U7943 (N_7943,N_7729,N_7728);
and U7944 (N_7944,N_7772,N_7563);
xor U7945 (N_7945,N_7726,N_7604);
nand U7946 (N_7946,N_7580,N_7532);
nand U7947 (N_7947,N_7682,N_7669);
or U7948 (N_7948,N_7622,N_7645);
xor U7949 (N_7949,N_7641,N_7769);
nand U7950 (N_7950,N_7758,N_7685);
and U7951 (N_7951,N_7644,N_7578);
nor U7952 (N_7952,N_7589,N_7665);
nand U7953 (N_7953,N_7726,N_7518);
and U7954 (N_7954,N_7689,N_7681);
nand U7955 (N_7955,N_7579,N_7591);
and U7956 (N_7956,N_7783,N_7709);
nand U7957 (N_7957,N_7671,N_7607);
nor U7958 (N_7958,N_7669,N_7652);
or U7959 (N_7959,N_7746,N_7544);
or U7960 (N_7960,N_7601,N_7518);
nor U7961 (N_7961,N_7534,N_7704);
nand U7962 (N_7962,N_7787,N_7694);
or U7963 (N_7963,N_7675,N_7587);
nor U7964 (N_7964,N_7749,N_7541);
and U7965 (N_7965,N_7758,N_7595);
or U7966 (N_7966,N_7516,N_7797);
nand U7967 (N_7967,N_7785,N_7534);
xor U7968 (N_7968,N_7581,N_7727);
or U7969 (N_7969,N_7752,N_7656);
xor U7970 (N_7970,N_7631,N_7768);
and U7971 (N_7971,N_7727,N_7569);
or U7972 (N_7972,N_7773,N_7745);
and U7973 (N_7973,N_7705,N_7780);
nor U7974 (N_7974,N_7522,N_7650);
xor U7975 (N_7975,N_7760,N_7764);
nand U7976 (N_7976,N_7730,N_7544);
and U7977 (N_7977,N_7731,N_7615);
and U7978 (N_7978,N_7786,N_7614);
and U7979 (N_7979,N_7690,N_7775);
nand U7980 (N_7980,N_7625,N_7694);
and U7981 (N_7981,N_7553,N_7640);
nor U7982 (N_7982,N_7595,N_7753);
or U7983 (N_7983,N_7564,N_7798);
and U7984 (N_7984,N_7513,N_7749);
xor U7985 (N_7985,N_7521,N_7789);
or U7986 (N_7986,N_7757,N_7603);
xnor U7987 (N_7987,N_7687,N_7567);
nor U7988 (N_7988,N_7628,N_7501);
xor U7989 (N_7989,N_7581,N_7606);
nor U7990 (N_7990,N_7723,N_7512);
or U7991 (N_7991,N_7719,N_7673);
nor U7992 (N_7992,N_7710,N_7589);
and U7993 (N_7993,N_7637,N_7731);
nand U7994 (N_7994,N_7717,N_7770);
nand U7995 (N_7995,N_7776,N_7733);
xor U7996 (N_7996,N_7633,N_7699);
and U7997 (N_7997,N_7672,N_7729);
and U7998 (N_7998,N_7538,N_7606);
nand U7999 (N_7999,N_7602,N_7506);
nand U8000 (N_8000,N_7697,N_7606);
and U8001 (N_8001,N_7738,N_7730);
xnor U8002 (N_8002,N_7741,N_7664);
nand U8003 (N_8003,N_7719,N_7510);
and U8004 (N_8004,N_7732,N_7634);
nor U8005 (N_8005,N_7628,N_7742);
xor U8006 (N_8006,N_7662,N_7753);
and U8007 (N_8007,N_7570,N_7597);
or U8008 (N_8008,N_7635,N_7523);
or U8009 (N_8009,N_7502,N_7770);
or U8010 (N_8010,N_7547,N_7777);
or U8011 (N_8011,N_7679,N_7668);
and U8012 (N_8012,N_7692,N_7563);
or U8013 (N_8013,N_7782,N_7671);
nand U8014 (N_8014,N_7619,N_7684);
and U8015 (N_8015,N_7572,N_7613);
xnor U8016 (N_8016,N_7661,N_7562);
or U8017 (N_8017,N_7566,N_7500);
nor U8018 (N_8018,N_7606,N_7710);
nand U8019 (N_8019,N_7780,N_7553);
nor U8020 (N_8020,N_7718,N_7752);
or U8021 (N_8021,N_7767,N_7662);
nor U8022 (N_8022,N_7768,N_7774);
and U8023 (N_8023,N_7659,N_7571);
nand U8024 (N_8024,N_7681,N_7632);
and U8025 (N_8025,N_7533,N_7781);
nor U8026 (N_8026,N_7603,N_7765);
nor U8027 (N_8027,N_7667,N_7698);
and U8028 (N_8028,N_7645,N_7715);
and U8029 (N_8029,N_7585,N_7627);
xnor U8030 (N_8030,N_7635,N_7605);
nand U8031 (N_8031,N_7719,N_7592);
or U8032 (N_8032,N_7755,N_7621);
nor U8033 (N_8033,N_7764,N_7509);
or U8034 (N_8034,N_7562,N_7645);
and U8035 (N_8035,N_7620,N_7693);
or U8036 (N_8036,N_7711,N_7567);
nand U8037 (N_8037,N_7529,N_7639);
nand U8038 (N_8038,N_7793,N_7536);
nor U8039 (N_8039,N_7523,N_7623);
nand U8040 (N_8040,N_7573,N_7501);
or U8041 (N_8041,N_7546,N_7681);
and U8042 (N_8042,N_7564,N_7659);
or U8043 (N_8043,N_7739,N_7536);
xor U8044 (N_8044,N_7746,N_7669);
nor U8045 (N_8045,N_7732,N_7613);
xnor U8046 (N_8046,N_7745,N_7608);
xor U8047 (N_8047,N_7672,N_7725);
nand U8048 (N_8048,N_7639,N_7553);
and U8049 (N_8049,N_7572,N_7693);
xnor U8050 (N_8050,N_7700,N_7641);
or U8051 (N_8051,N_7577,N_7621);
nand U8052 (N_8052,N_7768,N_7565);
and U8053 (N_8053,N_7674,N_7712);
or U8054 (N_8054,N_7734,N_7567);
and U8055 (N_8055,N_7734,N_7524);
and U8056 (N_8056,N_7693,N_7617);
xnor U8057 (N_8057,N_7516,N_7628);
or U8058 (N_8058,N_7699,N_7548);
and U8059 (N_8059,N_7747,N_7619);
and U8060 (N_8060,N_7702,N_7504);
and U8061 (N_8061,N_7667,N_7774);
and U8062 (N_8062,N_7601,N_7707);
or U8063 (N_8063,N_7710,N_7537);
xnor U8064 (N_8064,N_7720,N_7562);
nor U8065 (N_8065,N_7754,N_7501);
or U8066 (N_8066,N_7730,N_7520);
or U8067 (N_8067,N_7506,N_7666);
xnor U8068 (N_8068,N_7759,N_7507);
nand U8069 (N_8069,N_7712,N_7758);
and U8070 (N_8070,N_7798,N_7553);
and U8071 (N_8071,N_7569,N_7682);
nor U8072 (N_8072,N_7609,N_7665);
and U8073 (N_8073,N_7749,N_7596);
and U8074 (N_8074,N_7657,N_7761);
or U8075 (N_8075,N_7760,N_7734);
xnor U8076 (N_8076,N_7523,N_7556);
or U8077 (N_8077,N_7644,N_7793);
xor U8078 (N_8078,N_7710,N_7619);
xnor U8079 (N_8079,N_7580,N_7681);
nand U8080 (N_8080,N_7635,N_7514);
nor U8081 (N_8081,N_7736,N_7629);
xor U8082 (N_8082,N_7790,N_7742);
or U8083 (N_8083,N_7607,N_7567);
or U8084 (N_8084,N_7705,N_7755);
xor U8085 (N_8085,N_7658,N_7611);
or U8086 (N_8086,N_7580,N_7731);
nor U8087 (N_8087,N_7549,N_7628);
nor U8088 (N_8088,N_7542,N_7674);
nor U8089 (N_8089,N_7638,N_7765);
xnor U8090 (N_8090,N_7775,N_7666);
or U8091 (N_8091,N_7794,N_7711);
xor U8092 (N_8092,N_7779,N_7651);
nand U8093 (N_8093,N_7600,N_7514);
nor U8094 (N_8094,N_7675,N_7752);
xnor U8095 (N_8095,N_7647,N_7502);
nor U8096 (N_8096,N_7751,N_7587);
xnor U8097 (N_8097,N_7605,N_7546);
xor U8098 (N_8098,N_7611,N_7601);
or U8099 (N_8099,N_7743,N_7772);
xnor U8100 (N_8100,N_8093,N_7912);
and U8101 (N_8101,N_7980,N_8074);
nor U8102 (N_8102,N_7897,N_7917);
nor U8103 (N_8103,N_7857,N_7900);
xor U8104 (N_8104,N_7875,N_7825);
or U8105 (N_8105,N_7847,N_7932);
or U8106 (N_8106,N_7883,N_7863);
or U8107 (N_8107,N_7866,N_8010);
nor U8108 (N_8108,N_7987,N_7864);
nor U8109 (N_8109,N_7972,N_8024);
xor U8110 (N_8110,N_8003,N_8091);
or U8111 (N_8111,N_7975,N_8078);
or U8112 (N_8112,N_8057,N_8069);
xnor U8113 (N_8113,N_7874,N_8046);
or U8114 (N_8114,N_7877,N_7999);
nand U8115 (N_8115,N_7843,N_7837);
nor U8116 (N_8116,N_7887,N_7815);
nor U8117 (N_8117,N_8020,N_7803);
and U8118 (N_8118,N_8041,N_7898);
xnor U8119 (N_8119,N_8067,N_7964);
nor U8120 (N_8120,N_7858,N_7902);
or U8121 (N_8121,N_7833,N_7878);
or U8122 (N_8122,N_7926,N_7855);
nand U8123 (N_8123,N_8099,N_7827);
and U8124 (N_8124,N_8030,N_7846);
nand U8125 (N_8125,N_7981,N_7823);
and U8126 (N_8126,N_8080,N_7945);
or U8127 (N_8127,N_7831,N_8051);
nor U8128 (N_8128,N_7891,N_7916);
or U8129 (N_8129,N_7807,N_7920);
xnor U8130 (N_8130,N_8098,N_7885);
or U8131 (N_8131,N_8092,N_7995);
xor U8132 (N_8132,N_7871,N_7923);
or U8133 (N_8133,N_8026,N_7809);
nor U8134 (N_8134,N_8090,N_7997);
xor U8135 (N_8135,N_7895,N_7973);
nand U8136 (N_8136,N_7860,N_8081);
and U8137 (N_8137,N_7880,N_7838);
or U8138 (N_8138,N_7948,N_7955);
and U8139 (N_8139,N_7947,N_7940);
nor U8140 (N_8140,N_8094,N_8083);
or U8141 (N_8141,N_7852,N_7942);
and U8142 (N_8142,N_7805,N_7960);
xor U8143 (N_8143,N_7918,N_8012);
or U8144 (N_8144,N_7950,N_7908);
nand U8145 (N_8145,N_7856,N_7894);
nand U8146 (N_8146,N_7817,N_8004);
nand U8147 (N_8147,N_7931,N_8054);
xor U8148 (N_8148,N_8071,N_8015);
nand U8149 (N_8149,N_7909,N_7978);
and U8150 (N_8150,N_8076,N_7892);
nor U8151 (N_8151,N_7806,N_7849);
nor U8152 (N_8152,N_7826,N_7914);
or U8153 (N_8153,N_8043,N_7937);
nand U8154 (N_8154,N_7934,N_7861);
nand U8155 (N_8155,N_8022,N_7802);
nor U8156 (N_8156,N_7876,N_7842);
and U8157 (N_8157,N_8055,N_8047);
and U8158 (N_8158,N_7910,N_8050);
or U8159 (N_8159,N_7813,N_8096);
or U8160 (N_8160,N_8001,N_7824);
and U8161 (N_8161,N_8000,N_7906);
and U8162 (N_8162,N_7896,N_7800);
xnor U8163 (N_8163,N_7822,N_8097);
and U8164 (N_8164,N_7921,N_8082);
xnor U8165 (N_8165,N_7996,N_7966);
xor U8166 (N_8166,N_7974,N_7929);
and U8167 (N_8167,N_8014,N_7927);
nor U8168 (N_8168,N_7977,N_7954);
xnor U8169 (N_8169,N_8007,N_8018);
and U8170 (N_8170,N_7834,N_8029);
xor U8171 (N_8171,N_8059,N_8056);
nor U8172 (N_8172,N_7911,N_8009);
nor U8173 (N_8173,N_7936,N_8019);
or U8174 (N_8174,N_7935,N_7904);
or U8175 (N_8175,N_7924,N_7991);
and U8176 (N_8176,N_7844,N_7839);
or U8177 (N_8177,N_8036,N_7941);
or U8178 (N_8178,N_7946,N_8023);
nor U8179 (N_8179,N_8049,N_7998);
or U8180 (N_8180,N_7841,N_8085);
nor U8181 (N_8181,N_8031,N_7938);
xnor U8182 (N_8182,N_7867,N_7939);
or U8183 (N_8183,N_7928,N_7890);
and U8184 (N_8184,N_7899,N_7814);
or U8185 (N_8185,N_7956,N_7969);
nor U8186 (N_8186,N_7949,N_8033);
nand U8187 (N_8187,N_8064,N_8035);
or U8188 (N_8188,N_7905,N_7865);
nor U8189 (N_8189,N_7882,N_8028);
xor U8190 (N_8190,N_7970,N_8002);
xnor U8191 (N_8191,N_7993,N_8040);
xor U8192 (N_8192,N_7903,N_7990);
nor U8193 (N_8193,N_8070,N_7836);
xnor U8194 (N_8194,N_8073,N_7840);
nor U8195 (N_8195,N_7830,N_7951);
nand U8196 (N_8196,N_7992,N_7888);
or U8197 (N_8197,N_8008,N_8013);
nand U8198 (N_8198,N_8011,N_7957);
nand U8199 (N_8199,N_7832,N_8044);
nand U8200 (N_8200,N_7944,N_7961);
xor U8201 (N_8201,N_8025,N_7901);
xor U8202 (N_8202,N_7982,N_8065);
and U8203 (N_8203,N_8060,N_8042);
nor U8204 (N_8204,N_7952,N_7873);
nand U8205 (N_8205,N_8045,N_8048);
and U8206 (N_8206,N_7854,N_7818);
nor U8207 (N_8207,N_8079,N_7859);
and U8208 (N_8208,N_8005,N_7853);
or U8209 (N_8209,N_8017,N_7919);
nand U8210 (N_8210,N_8088,N_8021);
nor U8211 (N_8211,N_7862,N_7835);
and U8212 (N_8212,N_8038,N_7821);
nand U8213 (N_8213,N_8032,N_7979);
and U8214 (N_8214,N_8075,N_7870);
xnor U8215 (N_8215,N_7913,N_8027);
nand U8216 (N_8216,N_8016,N_7804);
nor U8217 (N_8217,N_7983,N_8084);
and U8218 (N_8218,N_7933,N_8095);
xnor U8219 (N_8219,N_8039,N_7968);
nand U8220 (N_8220,N_7881,N_7850);
and U8221 (N_8221,N_8052,N_8086);
nand U8222 (N_8222,N_8068,N_7958);
or U8223 (N_8223,N_7963,N_8006);
xnor U8224 (N_8224,N_7925,N_7848);
nand U8225 (N_8225,N_8063,N_7922);
xor U8226 (N_8226,N_7810,N_8072);
or U8227 (N_8227,N_7959,N_7893);
and U8228 (N_8228,N_7965,N_8077);
nor U8229 (N_8229,N_7884,N_8062);
nor U8230 (N_8230,N_7851,N_7953);
or U8231 (N_8231,N_7801,N_8087);
nand U8232 (N_8232,N_8089,N_8061);
nand U8233 (N_8233,N_7889,N_7820);
nor U8234 (N_8234,N_7869,N_7879);
xor U8235 (N_8235,N_7816,N_7985);
xor U8236 (N_8236,N_7986,N_8066);
or U8237 (N_8237,N_7845,N_7886);
nand U8238 (N_8238,N_8058,N_7962);
nor U8239 (N_8239,N_7989,N_7808);
nand U8240 (N_8240,N_8037,N_7943);
nor U8241 (N_8241,N_8053,N_7994);
xnor U8242 (N_8242,N_7971,N_7984);
xnor U8243 (N_8243,N_8034,N_7819);
or U8244 (N_8244,N_7872,N_7868);
nor U8245 (N_8245,N_7988,N_7976);
and U8246 (N_8246,N_7811,N_7828);
nor U8247 (N_8247,N_7829,N_7930);
nand U8248 (N_8248,N_7967,N_7907);
or U8249 (N_8249,N_7915,N_7812);
nor U8250 (N_8250,N_7912,N_7944);
and U8251 (N_8251,N_7803,N_7888);
nor U8252 (N_8252,N_8070,N_8093);
xor U8253 (N_8253,N_7831,N_7894);
nor U8254 (N_8254,N_7892,N_7938);
or U8255 (N_8255,N_7834,N_7929);
or U8256 (N_8256,N_7809,N_8008);
or U8257 (N_8257,N_8012,N_8072);
or U8258 (N_8258,N_7875,N_8083);
or U8259 (N_8259,N_7988,N_8042);
nand U8260 (N_8260,N_7844,N_7819);
or U8261 (N_8261,N_7808,N_8036);
or U8262 (N_8262,N_7848,N_8045);
and U8263 (N_8263,N_7800,N_7838);
xor U8264 (N_8264,N_8079,N_7955);
xor U8265 (N_8265,N_8058,N_7844);
nor U8266 (N_8266,N_8025,N_8028);
nand U8267 (N_8267,N_7943,N_7873);
or U8268 (N_8268,N_7916,N_7944);
nor U8269 (N_8269,N_7909,N_7853);
nor U8270 (N_8270,N_8092,N_8073);
nor U8271 (N_8271,N_7954,N_8013);
and U8272 (N_8272,N_8051,N_7847);
xnor U8273 (N_8273,N_7831,N_8006);
nand U8274 (N_8274,N_7923,N_7836);
and U8275 (N_8275,N_8056,N_8003);
and U8276 (N_8276,N_7808,N_7822);
nand U8277 (N_8277,N_8065,N_8080);
nand U8278 (N_8278,N_7990,N_8022);
nor U8279 (N_8279,N_7849,N_8040);
xnor U8280 (N_8280,N_7921,N_8006);
or U8281 (N_8281,N_8056,N_8029);
nor U8282 (N_8282,N_8099,N_8045);
or U8283 (N_8283,N_8008,N_8030);
xor U8284 (N_8284,N_7805,N_8099);
nor U8285 (N_8285,N_7943,N_7911);
nand U8286 (N_8286,N_7877,N_7809);
or U8287 (N_8287,N_8003,N_8027);
nor U8288 (N_8288,N_7867,N_8045);
and U8289 (N_8289,N_7828,N_7886);
and U8290 (N_8290,N_8083,N_7950);
nor U8291 (N_8291,N_7898,N_8007);
and U8292 (N_8292,N_8050,N_7843);
or U8293 (N_8293,N_8046,N_7823);
xor U8294 (N_8294,N_7883,N_8038);
nor U8295 (N_8295,N_7828,N_7993);
nor U8296 (N_8296,N_7953,N_7934);
or U8297 (N_8297,N_7909,N_7852);
or U8298 (N_8298,N_7882,N_7803);
xnor U8299 (N_8299,N_7824,N_8069);
nand U8300 (N_8300,N_7979,N_7952);
or U8301 (N_8301,N_7994,N_8039);
xnor U8302 (N_8302,N_7827,N_8053);
nor U8303 (N_8303,N_8050,N_7917);
xor U8304 (N_8304,N_8077,N_7855);
and U8305 (N_8305,N_8003,N_7993);
and U8306 (N_8306,N_7933,N_7925);
nor U8307 (N_8307,N_7918,N_7857);
nor U8308 (N_8308,N_8084,N_7887);
or U8309 (N_8309,N_8095,N_8043);
nor U8310 (N_8310,N_7855,N_8026);
nand U8311 (N_8311,N_8046,N_7849);
and U8312 (N_8312,N_7834,N_8056);
and U8313 (N_8313,N_7949,N_7930);
nor U8314 (N_8314,N_7859,N_7821);
nand U8315 (N_8315,N_7863,N_8011);
nor U8316 (N_8316,N_7964,N_7940);
xor U8317 (N_8317,N_7910,N_8051);
nor U8318 (N_8318,N_7904,N_8047);
xnor U8319 (N_8319,N_8079,N_8075);
nand U8320 (N_8320,N_7804,N_7912);
nor U8321 (N_8321,N_8067,N_7923);
or U8322 (N_8322,N_7874,N_7973);
xor U8323 (N_8323,N_8034,N_7927);
and U8324 (N_8324,N_7918,N_7887);
or U8325 (N_8325,N_8076,N_7900);
or U8326 (N_8326,N_7923,N_8044);
nor U8327 (N_8327,N_8024,N_7898);
nor U8328 (N_8328,N_7923,N_7848);
xnor U8329 (N_8329,N_8006,N_7968);
xnor U8330 (N_8330,N_8055,N_7996);
nand U8331 (N_8331,N_8097,N_7840);
and U8332 (N_8332,N_8091,N_7973);
nand U8333 (N_8333,N_7878,N_7992);
nand U8334 (N_8334,N_8044,N_7899);
xnor U8335 (N_8335,N_7957,N_8044);
nand U8336 (N_8336,N_8027,N_8079);
and U8337 (N_8337,N_8059,N_7956);
nand U8338 (N_8338,N_8073,N_8036);
or U8339 (N_8339,N_8038,N_7896);
and U8340 (N_8340,N_8028,N_7984);
or U8341 (N_8341,N_7893,N_8076);
xnor U8342 (N_8342,N_7983,N_7986);
and U8343 (N_8343,N_8029,N_8024);
or U8344 (N_8344,N_8038,N_8013);
nor U8345 (N_8345,N_7958,N_7841);
and U8346 (N_8346,N_7900,N_8061);
or U8347 (N_8347,N_8087,N_8069);
xnor U8348 (N_8348,N_8007,N_7974);
and U8349 (N_8349,N_8027,N_8086);
and U8350 (N_8350,N_7836,N_7838);
nor U8351 (N_8351,N_7982,N_7811);
or U8352 (N_8352,N_8094,N_7889);
or U8353 (N_8353,N_7939,N_8032);
xor U8354 (N_8354,N_7901,N_8073);
and U8355 (N_8355,N_7958,N_7859);
nand U8356 (N_8356,N_7943,N_7905);
and U8357 (N_8357,N_7894,N_7918);
nor U8358 (N_8358,N_7887,N_7951);
nor U8359 (N_8359,N_7802,N_7974);
nand U8360 (N_8360,N_7972,N_8032);
xnor U8361 (N_8361,N_7806,N_7883);
or U8362 (N_8362,N_7972,N_8016);
nand U8363 (N_8363,N_7844,N_7936);
nor U8364 (N_8364,N_7811,N_7824);
nor U8365 (N_8365,N_7904,N_7826);
xor U8366 (N_8366,N_7915,N_8015);
nand U8367 (N_8367,N_7830,N_7929);
xor U8368 (N_8368,N_7968,N_7919);
or U8369 (N_8369,N_8034,N_7899);
nand U8370 (N_8370,N_8020,N_7882);
nand U8371 (N_8371,N_8074,N_7897);
xor U8372 (N_8372,N_8047,N_7944);
nor U8373 (N_8373,N_7953,N_8034);
and U8374 (N_8374,N_7918,N_7868);
nand U8375 (N_8375,N_7882,N_7853);
or U8376 (N_8376,N_7865,N_8013);
and U8377 (N_8377,N_8069,N_7941);
and U8378 (N_8378,N_8021,N_7907);
nand U8379 (N_8379,N_7952,N_7971);
nand U8380 (N_8380,N_8011,N_8079);
nor U8381 (N_8381,N_7911,N_7910);
nand U8382 (N_8382,N_7872,N_7989);
nor U8383 (N_8383,N_7949,N_7811);
xnor U8384 (N_8384,N_7970,N_7885);
nor U8385 (N_8385,N_7931,N_8071);
nor U8386 (N_8386,N_8073,N_7859);
nor U8387 (N_8387,N_7811,N_8054);
nor U8388 (N_8388,N_8078,N_8088);
nor U8389 (N_8389,N_7947,N_8010);
nand U8390 (N_8390,N_7962,N_7997);
nand U8391 (N_8391,N_8057,N_8058);
or U8392 (N_8392,N_8046,N_7992);
xnor U8393 (N_8393,N_8021,N_7962);
nor U8394 (N_8394,N_8091,N_7993);
nor U8395 (N_8395,N_8062,N_7941);
or U8396 (N_8396,N_7919,N_8090);
nor U8397 (N_8397,N_7846,N_7993);
or U8398 (N_8398,N_7896,N_8063);
xnor U8399 (N_8399,N_8073,N_7975);
nand U8400 (N_8400,N_8318,N_8243);
nand U8401 (N_8401,N_8224,N_8305);
and U8402 (N_8402,N_8369,N_8126);
xor U8403 (N_8403,N_8306,N_8356);
nor U8404 (N_8404,N_8276,N_8112);
nand U8405 (N_8405,N_8185,N_8107);
nor U8406 (N_8406,N_8157,N_8178);
and U8407 (N_8407,N_8390,N_8182);
or U8408 (N_8408,N_8140,N_8314);
xnor U8409 (N_8409,N_8193,N_8268);
or U8410 (N_8410,N_8387,N_8102);
or U8411 (N_8411,N_8395,N_8329);
xnor U8412 (N_8412,N_8325,N_8374);
nor U8413 (N_8413,N_8304,N_8239);
nor U8414 (N_8414,N_8352,N_8308);
xor U8415 (N_8415,N_8150,N_8353);
and U8416 (N_8416,N_8364,N_8257);
and U8417 (N_8417,N_8132,N_8171);
nor U8418 (N_8418,N_8203,N_8251);
or U8419 (N_8419,N_8265,N_8238);
nand U8420 (N_8420,N_8322,N_8146);
xor U8421 (N_8421,N_8263,N_8255);
nor U8422 (N_8422,N_8281,N_8247);
nand U8423 (N_8423,N_8365,N_8259);
xnor U8424 (N_8424,N_8350,N_8335);
nand U8425 (N_8425,N_8381,N_8375);
or U8426 (N_8426,N_8346,N_8175);
nor U8427 (N_8427,N_8160,N_8371);
xor U8428 (N_8428,N_8168,N_8159);
nand U8429 (N_8429,N_8229,N_8167);
nor U8430 (N_8430,N_8279,N_8372);
xor U8431 (N_8431,N_8202,N_8319);
nor U8432 (N_8432,N_8170,N_8331);
nor U8433 (N_8433,N_8339,N_8392);
xnor U8434 (N_8434,N_8122,N_8378);
nand U8435 (N_8435,N_8271,N_8248);
or U8436 (N_8436,N_8256,N_8245);
nand U8437 (N_8437,N_8343,N_8184);
nor U8438 (N_8438,N_8153,N_8137);
xor U8439 (N_8439,N_8336,N_8138);
or U8440 (N_8440,N_8292,N_8133);
nand U8441 (N_8441,N_8234,N_8384);
xor U8442 (N_8442,N_8382,N_8301);
nor U8443 (N_8443,N_8135,N_8192);
nand U8444 (N_8444,N_8164,N_8210);
or U8445 (N_8445,N_8345,N_8307);
and U8446 (N_8446,N_8337,N_8377);
nor U8447 (N_8447,N_8199,N_8187);
xnor U8448 (N_8448,N_8396,N_8101);
and U8449 (N_8449,N_8373,N_8209);
xnor U8450 (N_8450,N_8389,N_8129);
or U8451 (N_8451,N_8127,N_8363);
xnor U8452 (N_8452,N_8147,N_8399);
nand U8453 (N_8453,N_8262,N_8113);
nand U8454 (N_8454,N_8286,N_8354);
xnor U8455 (N_8455,N_8278,N_8130);
nand U8456 (N_8456,N_8148,N_8252);
nand U8457 (N_8457,N_8172,N_8144);
nand U8458 (N_8458,N_8273,N_8212);
xor U8459 (N_8459,N_8360,N_8228);
or U8460 (N_8460,N_8161,N_8289);
and U8461 (N_8461,N_8211,N_8358);
nor U8462 (N_8462,N_8200,N_8328);
nor U8463 (N_8463,N_8244,N_8183);
xnor U8464 (N_8464,N_8264,N_8297);
and U8465 (N_8465,N_8205,N_8317);
xnor U8466 (N_8466,N_8320,N_8221);
or U8467 (N_8467,N_8355,N_8338);
nor U8468 (N_8468,N_8176,N_8272);
or U8469 (N_8469,N_8299,N_8333);
nand U8470 (N_8470,N_8115,N_8136);
xor U8471 (N_8471,N_8283,N_8284);
xor U8472 (N_8472,N_8206,N_8368);
xor U8473 (N_8473,N_8311,N_8195);
nor U8474 (N_8474,N_8242,N_8323);
nor U8475 (N_8475,N_8121,N_8258);
xor U8476 (N_8476,N_8109,N_8204);
nor U8477 (N_8477,N_8312,N_8142);
xor U8478 (N_8478,N_8391,N_8223);
nand U8479 (N_8479,N_8222,N_8191);
nor U8480 (N_8480,N_8327,N_8118);
nor U8481 (N_8481,N_8145,N_8134);
xor U8482 (N_8482,N_8119,N_8326);
nor U8483 (N_8483,N_8198,N_8298);
or U8484 (N_8484,N_8232,N_8341);
xor U8485 (N_8485,N_8186,N_8174);
xor U8486 (N_8486,N_8190,N_8347);
nand U8487 (N_8487,N_8310,N_8131);
xnor U8488 (N_8488,N_8141,N_8287);
or U8489 (N_8489,N_8106,N_8367);
xor U8490 (N_8490,N_8386,N_8351);
and U8491 (N_8491,N_8316,N_8117);
nand U8492 (N_8492,N_8240,N_8154);
and U8493 (N_8493,N_8366,N_8296);
and U8494 (N_8494,N_8197,N_8393);
or U8495 (N_8495,N_8397,N_8380);
and U8496 (N_8496,N_8215,N_8213);
nor U8497 (N_8497,N_8293,N_8230);
nor U8498 (N_8498,N_8165,N_8383);
or U8499 (N_8499,N_8250,N_8340);
nand U8500 (N_8500,N_8321,N_8196);
nand U8501 (N_8501,N_8158,N_8156);
or U8502 (N_8502,N_8181,N_8249);
nor U8503 (N_8503,N_8235,N_8225);
xor U8504 (N_8504,N_8166,N_8285);
nor U8505 (N_8505,N_8385,N_8108);
nor U8506 (N_8506,N_8388,N_8324);
nand U8507 (N_8507,N_8237,N_8163);
xnor U8508 (N_8508,N_8344,N_8100);
nor U8509 (N_8509,N_8103,N_8313);
and U8510 (N_8510,N_8280,N_8201);
nor U8511 (N_8511,N_8120,N_8295);
nand U8512 (N_8512,N_8116,N_8180);
xor U8513 (N_8513,N_8216,N_8291);
and U8514 (N_8514,N_8348,N_8110);
xor U8515 (N_8515,N_8309,N_8398);
and U8516 (N_8516,N_8188,N_8143);
nand U8517 (N_8517,N_8357,N_8227);
nor U8518 (N_8518,N_8236,N_8139);
nand U8519 (N_8519,N_8288,N_8123);
xnor U8520 (N_8520,N_8349,N_8274);
xnor U8521 (N_8521,N_8394,N_8155);
and U8522 (N_8522,N_8246,N_8342);
or U8523 (N_8523,N_8253,N_8151);
nor U8524 (N_8524,N_8125,N_8359);
or U8525 (N_8525,N_8332,N_8294);
nor U8526 (N_8526,N_8208,N_8105);
and U8527 (N_8527,N_8303,N_8162);
nand U8528 (N_8528,N_8315,N_8362);
nor U8529 (N_8529,N_8330,N_8282);
and U8530 (N_8530,N_8214,N_8173);
xnor U8531 (N_8531,N_8370,N_8220);
or U8532 (N_8532,N_8169,N_8300);
nand U8533 (N_8533,N_8241,N_8217);
nand U8534 (N_8534,N_8334,N_8218);
nand U8535 (N_8535,N_8104,N_8260);
nor U8536 (N_8536,N_8207,N_8267);
xor U8537 (N_8537,N_8226,N_8379);
nand U8538 (N_8538,N_8277,N_8290);
nor U8539 (N_8539,N_8266,N_8128);
nor U8540 (N_8540,N_8361,N_8219);
nand U8541 (N_8541,N_8152,N_8302);
nand U8542 (N_8542,N_8275,N_8189);
and U8543 (N_8543,N_8179,N_8270);
nand U8544 (N_8544,N_8261,N_8149);
nor U8545 (N_8545,N_8114,N_8194);
and U8546 (N_8546,N_8231,N_8269);
and U8547 (N_8547,N_8233,N_8124);
and U8548 (N_8548,N_8177,N_8111);
nand U8549 (N_8549,N_8376,N_8254);
xnor U8550 (N_8550,N_8319,N_8184);
or U8551 (N_8551,N_8321,N_8223);
nor U8552 (N_8552,N_8341,N_8321);
nand U8553 (N_8553,N_8236,N_8334);
xor U8554 (N_8554,N_8341,N_8205);
or U8555 (N_8555,N_8356,N_8273);
and U8556 (N_8556,N_8105,N_8229);
nand U8557 (N_8557,N_8304,N_8386);
nand U8558 (N_8558,N_8181,N_8118);
and U8559 (N_8559,N_8242,N_8113);
and U8560 (N_8560,N_8131,N_8196);
xor U8561 (N_8561,N_8386,N_8211);
and U8562 (N_8562,N_8287,N_8239);
xor U8563 (N_8563,N_8391,N_8353);
nand U8564 (N_8564,N_8318,N_8398);
and U8565 (N_8565,N_8236,N_8158);
or U8566 (N_8566,N_8141,N_8255);
nor U8567 (N_8567,N_8242,N_8216);
nand U8568 (N_8568,N_8169,N_8132);
nor U8569 (N_8569,N_8237,N_8267);
and U8570 (N_8570,N_8376,N_8314);
and U8571 (N_8571,N_8110,N_8345);
nand U8572 (N_8572,N_8391,N_8202);
nand U8573 (N_8573,N_8231,N_8220);
nand U8574 (N_8574,N_8280,N_8374);
and U8575 (N_8575,N_8172,N_8387);
and U8576 (N_8576,N_8144,N_8213);
and U8577 (N_8577,N_8166,N_8102);
nand U8578 (N_8578,N_8164,N_8147);
and U8579 (N_8579,N_8119,N_8396);
nand U8580 (N_8580,N_8193,N_8106);
xnor U8581 (N_8581,N_8368,N_8258);
nor U8582 (N_8582,N_8163,N_8188);
nor U8583 (N_8583,N_8259,N_8244);
and U8584 (N_8584,N_8103,N_8220);
nor U8585 (N_8585,N_8290,N_8236);
nor U8586 (N_8586,N_8374,N_8289);
and U8587 (N_8587,N_8359,N_8342);
and U8588 (N_8588,N_8164,N_8391);
xor U8589 (N_8589,N_8325,N_8289);
and U8590 (N_8590,N_8101,N_8208);
xor U8591 (N_8591,N_8175,N_8232);
and U8592 (N_8592,N_8351,N_8303);
nor U8593 (N_8593,N_8397,N_8231);
and U8594 (N_8594,N_8148,N_8154);
nor U8595 (N_8595,N_8228,N_8342);
or U8596 (N_8596,N_8316,N_8241);
and U8597 (N_8597,N_8364,N_8328);
or U8598 (N_8598,N_8191,N_8335);
xor U8599 (N_8599,N_8314,N_8393);
nor U8600 (N_8600,N_8126,N_8159);
nand U8601 (N_8601,N_8255,N_8146);
xor U8602 (N_8602,N_8398,N_8259);
nor U8603 (N_8603,N_8193,N_8131);
and U8604 (N_8604,N_8326,N_8324);
and U8605 (N_8605,N_8179,N_8183);
or U8606 (N_8606,N_8358,N_8326);
nand U8607 (N_8607,N_8246,N_8245);
or U8608 (N_8608,N_8130,N_8299);
or U8609 (N_8609,N_8357,N_8249);
and U8610 (N_8610,N_8126,N_8144);
or U8611 (N_8611,N_8397,N_8272);
nor U8612 (N_8612,N_8297,N_8188);
and U8613 (N_8613,N_8139,N_8193);
xor U8614 (N_8614,N_8130,N_8158);
nand U8615 (N_8615,N_8128,N_8212);
or U8616 (N_8616,N_8318,N_8372);
nand U8617 (N_8617,N_8331,N_8184);
and U8618 (N_8618,N_8137,N_8343);
nor U8619 (N_8619,N_8283,N_8301);
and U8620 (N_8620,N_8182,N_8142);
or U8621 (N_8621,N_8133,N_8280);
nand U8622 (N_8622,N_8281,N_8321);
nor U8623 (N_8623,N_8321,N_8110);
and U8624 (N_8624,N_8390,N_8292);
and U8625 (N_8625,N_8356,N_8376);
nand U8626 (N_8626,N_8310,N_8136);
and U8627 (N_8627,N_8251,N_8103);
nand U8628 (N_8628,N_8385,N_8247);
nand U8629 (N_8629,N_8333,N_8286);
nand U8630 (N_8630,N_8174,N_8102);
and U8631 (N_8631,N_8314,N_8275);
and U8632 (N_8632,N_8392,N_8320);
nor U8633 (N_8633,N_8116,N_8364);
xnor U8634 (N_8634,N_8374,N_8270);
or U8635 (N_8635,N_8343,N_8247);
nor U8636 (N_8636,N_8106,N_8130);
nand U8637 (N_8637,N_8240,N_8244);
and U8638 (N_8638,N_8178,N_8330);
and U8639 (N_8639,N_8385,N_8196);
and U8640 (N_8640,N_8247,N_8357);
nand U8641 (N_8641,N_8268,N_8281);
and U8642 (N_8642,N_8178,N_8149);
or U8643 (N_8643,N_8314,N_8247);
nor U8644 (N_8644,N_8225,N_8333);
or U8645 (N_8645,N_8269,N_8309);
or U8646 (N_8646,N_8111,N_8290);
or U8647 (N_8647,N_8344,N_8174);
nor U8648 (N_8648,N_8378,N_8359);
nand U8649 (N_8649,N_8228,N_8199);
and U8650 (N_8650,N_8244,N_8342);
xor U8651 (N_8651,N_8220,N_8192);
or U8652 (N_8652,N_8296,N_8113);
nand U8653 (N_8653,N_8270,N_8241);
nand U8654 (N_8654,N_8302,N_8173);
and U8655 (N_8655,N_8310,N_8388);
nor U8656 (N_8656,N_8304,N_8278);
or U8657 (N_8657,N_8323,N_8163);
and U8658 (N_8658,N_8149,N_8145);
or U8659 (N_8659,N_8185,N_8326);
nand U8660 (N_8660,N_8252,N_8194);
and U8661 (N_8661,N_8103,N_8211);
xor U8662 (N_8662,N_8138,N_8184);
or U8663 (N_8663,N_8271,N_8261);
and U8664 (N_8664,N_8137,N_8373);
nor U8665 (N_8665,N_8230,N_8366);
nor U8666 (N_8666,N_8335,N_8332);
or U8667 (N_8667,N_8190,N_8140);
or U8668 (N_8668,N_8381,N_8258);
xnor U8669 (N_8669,N_8306,N_8150);
and U8670 (N_8670,N_8133,N_8283);
or U8671 (N_8671,N_8348,N_8237);
nor U8672 (N_8672,N_8213,N_8111);
nand U8673 (N_8673,N_8274,N_8398);
and U8674 (N_8674,N_8265,N_8183);
or U8675 (N_8675,N_8316,N_8332);
nor U8676 (N_8676,N_8152,N_8150);
xor U8677 (N_8677,N_8213,N_8137);
xnor U8678 (N_8678,N_8188,N_8158);
xor U8679 (N_8679,N_8330,N_8115);
and U8680 (N_8680,N_8198,N_8361);
xor U8681 (N_8681,N_8274,N_8262);
and U8682 (N_8682,N_8168,N_8267);
or U8683 (N_8683,N_8241,N_8214);
nand U8684 (N_8684,N_8383,N_8222);
xor U8685 (N_8685,N_8319,N_8299);
xnor U8686 (N_8686,N_8174,N_8356);
xor U8687 (N_8687,N_8106,N_8354);
nor U8688 (N_8688,N_8155,N_8287);
nand U8689 (N_8689,N_8351,N_8396);
or U8690 (N_8690,N_8207,N_8191);
nor U8691 (N_8691,N_8143,N_8112);
xnor U8692 (N_8692,N_8263,N_8231);
and U8693 (N_8693,N_8384,N_8115);
nor U8694 (N_8694,N_8109,N_8231);
and U8695 (N_8695,N_8246,N_8102);
or U8696 (N_8696,N_8109,N_8100);
nand U8697 (N_8697,N_8208,N_8319);
nand U8698 (N_8698,N_8171,N_8203);
or U8699 (N_8699,N_8398,N_8170);
nand U8700 (N_8700,N_8423,N_8613);
xnor U8701 (N_8701,N_8517,N_8579);
and U8702 (N_8702,N_8584,N_8467);
xnor U8703 (N_8703,N_8448,N_8561);
nand U8704 (N_8704,N_8475,N_8491);
nand U8705 (N_8705,N_8618,N_8424);
or U8706 (N_8706,N_8521,N_8673);
nand U8707 (N_8707,N_8648,N_8470);
or U8708 (N_8708,N_8615,N_8401);
nor U8709 (N_8709,N_8505,N_8434);
xnor U8710 (N_8710,N_8578,N_8688);
or U8711 (N_8711,N_8426,N_8440);
and U8712 (N_8712,N_8554,N_8576);
nor U8713 (N_8713,N_8632,N_8452);
and U8714 (N_8714,N_8485,N_8597);
and U8715 (N_8715,N_8680,N_8450);
xnor U8716 (N_8716,N_8410,N_8690);
xnor U8717 (N_8717,N_8626,N_8533);
nand U8718 (N_8718,N_8596,N_8464);
nand U8719 (N_8719,N_8620,N_8551);
and U8720 (N_8720,N_8590,N_8635);
xor U8721 (N_8721,N_8670,N_8520);
and U8722 (N_8722,N_8624,N_8549);
nand U8723 (N_8723,N_8543,N_8659);
nand U8724 (N_8724,N_8519,N_8693);
xor U8725 (N_8725,N_8556,N_8604);
or U8726 (N_8726,N_8478,N_8495);
xnor U8727 (N_8727,N_8665,N_8600);
and U8728 (N_8728,N_8555,N_8611);
nor U8729 (N_8729,N_8638,N_8487);
nor U8730 (N_8730,N_8686,N_8658);
xnor U8731 (N_8731,N_8559,N_8443);
and U8732 (N_8732,N_8647,N_8449);
xnor U8733 (N_8733,N_8523,N_8537);
and U8734 (N_8734,N_8593,N_8545);
xnor U8735 (N_8735,N_8570,N_8546);
nand U8736 (N_8736,N_8544,N_8674);
and U8737 (N_8737,N_8627,N_8640);
nand U8738 (N_8738,N_8431,N_8493);
and U8739 (N_8739,N_8438,N_8528);
or U8740 (N_8740,N_8535,N_8451);
and U8741 (N_8741,N_8583,N_8502);
nand U8742 (N_8742,N_8433,N_8422);
nand U8743 (N_8743,N_8661,N_8617);
nand U8744 (N_8744,N_8653,N_8650);
xnor U8745 (N_8745,N_8633,N_8514);
nor U8746 (N_8746,N_8466,N_8622);
and U8747 (N_8747,N_8513,N_8542);
and U8748 (N_8748,N_8420,N_8530);
nand U8749 (N_8749,N_8529,N_8527);
nor U8750 (N_8750,N_8492,N_8508);
or U8751 (N_8751,N_8403,N_8500);
xnor U8752 (N_8752,N_8415,N_8419);
or U8753 (N_8753,N_8531,N_8616);
xnor U8754 (N_8754,N_8473,N_8516);
nor U8755 (N_8755,N_8557,N_8462);
or U8756 (N_8756,N_8538,N_8453);
xor U8757 (N_8757,N_8581,N_8414);
nand U8758 (N_8758,N_8479,N_8636);
nand U8759 (N_8759,N_8628,N_8501);
xor U8760 (N_8760,N_8458,N_8660);
nor U8761 (N_8761,N_8646,N_8698);
xor U8762 (N_8762,N_8631,N_8413);
xor U8763 (N_8763,N_8696,N_8418);
xnor U8764 (N_8764,N_8656,N_8643);
xor U8765 (N_8765,N_8577,N_8678);
nor U8766 (N_8766,N_8573,N_8614);
nor U8767 (N_8767,N_8663,N_8691);
or U8768 (N_8768,N_8540,N_8507);
or U8769 (N_8769,N_8655,N_8598);
nor U8770 (N_8770,N_8454,N_8547);
or U8771 (N_8771,N_8474,N_8667);
nand U8772 (N_8772,N_8601,N_8687);
xor U8773 (N_8773,N_8496,N_8476);
or U8774 (N_8774,N_8605,N_8683);
xor U8775 (N_8775,N_8697,N_8651);
nor U8776 (N_8776,N_8400,N_8587);
nor U8777 (N_8777,N_8506,N_8518);
nand U8778 (N_8778,N_8405,N_8439);
nand U8779 (N_8779,N_8417,N_8565);
xor U8780 (N_8780,N_8681,N_8652);
and U8781 (N_8781,N_8568,N_8599);
nor U8782 (N_8782,N_8629,N_8482);
xnor U8783 (N_8783,N_8428,N_8526);
xor U8784 (N_8784,N_8436,N_8645);
nor U8785 (N_8785,N_8657,N_8689);
xnor U8786 (N_8786,N_8582,N_8494);
xnor U8787 (N_8787,N_8532,N_8457);
or U8788 (N_8788,N_8606,N_8447);
xnor U8789 (N_8789,N_8490,N_8484);
nand U8790 (N_8790,N_8682,N_8563);
xnor U8791 (N_8791,N_8404,N_8621);
nand U8792 (N_8792,N_8463,N_8639);
or U8793 (N_8793,N_8664,N_8602);
or U8794 (N_8794,N_8619,N_8625);
and U8795 (N_8795,N_8432,N_8416);
and U8796 (N_8796,N_8679,N_8407);
and U8797 (N_8797,N_8497,N_8566);
or U8798 (N_8798,N_8504,N_8649);
and U8799 (N_8799,N_8610,N_8692);
xnor U8800 (N_8800,N_8553,N_8435);
xor U8801 (N_8801,N_8609,N_8522);
nand U8802 (N_8802,N_8575,N_8552);
nor U8803 (N_8803,N_8525,N_8548);
xor U8804 (N_8804,N_8562,N_8511);
xnor U8805 (N_8805,N_8580,N_8489);
xnor U8806 (N_8806,N_8498,N_8699);
xor U8807 (N_8807,N_8477,N_8441);
xnor U8808 (N_8808,N_8595,N_8574);
nor U8809 (N_8809,N_8586,N_8402);
xor U8810 (N_8810,N_8445,N_8503);
nor U8811 (N_8811,N_8499,N_8571);
nor U8812 (N_8812,N_8666,N_8472);
xor U8813 (N_8813,N_8671,N_8483);
xnor U8814 (N_8814,N_8471,N_8572);
nor U8815 (N_8815,N_8588,N_8408);
nor U8816 (N_8816,N_8409,N_8406);
xor U8817 (N_8817,N_8642,N_8594);
nand U8818 (N_8818,N_8567,N_8480);
xor U8819 (N_8819,N_8607,N_8486);
nor U8820 (N_8820,N_8672,N_8677);
nor U8821 (N_8821,N_8564,N_8539);
nor U8822 (N_8822,N_8468,N_8534);
nor U8823 (N_8823,N_8469,N_8481);
nor U8824 (N_8824,N_8459,N_8460);
and U8825 (N_8825,N_8591,N_8644);
and U8826 (N_8826,N_8694,N_8411);
or U8827 (N_8827,N_8592,N_8429);
or U8828 (N_8828,N_8536,N_8560);
nand U8829 (N_8829,N_8662,N_8510);
or U8830 (N_8830,N_8675,N_8465);
nand U8831 (N_8831,N_8676,N_8455);
xor U8832 (N_8832,N_8603,N_8585);
nand U8833 (N_8833,N_8437,N_8442);
nand U8834 (N_8834,N_8488,N_8654);
nor U8835 (N_8835,N_8608,N_8637);
xnor U8836 (N_8836,N_8412,N_8541);
or U8837 (N_8837,N_8524,N_8550);
nor U8838 (N_8838,N_8684,N_8612);
xnor U8839 (N_8839,N_8512,N_8669);
and U8840 (N_8840,N_8668,N_8634);
and U8841 (N_8841,N_8558,N_8427);
and U8842 (N_8842,N_8461,N_8695);
nor U8843 (N_8843,N_8444,N_8589);
nor U8844 (N_8844,N_8430,N_8509);
or U8845 (N_8845,N_8425,N_8569);
or U8846 (N_8846,N_8630,N_8623);
xnor U8847 (N_8847,N_8421,N_8685);
xor U8848 (N_8848,N_8641,N_8515);
or U8849 (N_8849,N_8456,N_8446);
nor U8850 (N_8850,N_8683,N_8606);
or U8851 (N_8851,N_8669,N_8530);
and U8852 (N_8852,N_8451,N_8561);
and U8853 (N_8853,N_8449,N_8600);
nand U8854 (N_8854,N_8642,N_8511);
nand U8855 (N_8855,N_8656,N_8507);
xor U8856 (N_8856,N_8657,N_8654);
and U8857 (N_8857,N_8467,N_8689);
or U8858 (N_8858,N_8462,N_8486);
nand U8859 (N_8859,N_8667,N_8485);
nand U8860 (N_8860,N_8523,N_8647);
nor U8861 (N_8861,N_8412,N_8492);
nand U8862 (N_8862,N_8642,N_8540);
or U8863 (N_8863,N_8468,N_8476);
or U8864 (N_8864,N_8556,N_8690);
nand U8865 (N_8865,N_8626,N_8527);
and U8866 (N_8866,N_8600,N_8661);
nand U8867 (N_8867,N_8655,N_8677);
nand U8868 (N_8868,N_8501,N_8513);
nor U8869 (N_8869,N_8527,N_8407);
or U8870 (N_8870,N_8513,N_8578);
and U8871 (N_8871,N_8575,N_8421);
xnor U8872 (N_8872,N_8451,N_8526);
and U8873 (N_8873,N_8579,N_8450);
xor U8874 (N_8874,N_8465,N_8571);
or U8875 (N_8875,N_8594,N_8431);
or U8876 (N_8876,N_8617,N_8534);
and U8877 (N_8877,N_8470,N_8577);
nor U8878 (N_8878,N_8508,N_8407);
xnor U8879 (N_8879,N_8696,N_8552);
xnor U8880 (N_8880,N_8581,N_8401);
nor U8881 (N_8881,N_8519,N_8603);
xor U8882 (N_8882,N_8513,N_8685);
and U8883 (N_8883,N_8572,N_8501);
nand U8884 (N_8884,N_8546,N_8588);
or U8885 (N_8885,N_8637,N_8402);
and U8886 (N_8886,N_8557,N_8527);
and U8887 (N_8887,N_8421,N_8500);
nor U8888 (N_8888,N_8491,N_8402);
xnor U8889 (N_8889,N_8598,N_8517);
nand U8890 (N_8890,N_8607,N_8595);
xnor U8891 (N_8891,N_8582,N_8410);
and U8892 (N_8892,N_8636,N_8464);
or U8893 (N_8893,N_8507,N_8685);
nor U8894 (N_8894,N_8449,N_8481);
and U8895 (N_8895,N_8558,N_8698);
or U8896 (N_8896,N_8586,N_8614);
xor U8897 (N_8897,N_8537,N_8429);
or U8898 (N_8898,N_8502,N_8493);
xnor U8899 (N_8899,N_8429,N_8473);
nand U8900 (N_8900,N_8525,N_8630);
nor U8901 (N_8901,N_8458,N_8691);
and U8902 (N_8902,N_8493,N_8533);
nor U8903 (N_8903,N_8499,N_8426);
and U8904 (N_8904,N_8441,N_8485);
nor U8905 (N_8905,N_8528,N_8550);
xnor U8906 (N_8906,N_8606,N_8442);
and U8907 (N_8907,N_8601,N_8437);
and U8908 (N_8908,N_8484,N_8640);
xor U8909 (N_8909,N_8639,N_8429);
and U8910 (N_8910,N_8508,N_8571);
xor U8911 (N_8911,N_8666,N_8553);
or U8912 (N_8912,N_8455,N_8614);
or U8913 (N_8913,N_8456,N_8414);
or U8914 (N_8914,N_8626,N_8496);
nor U8915 (N_8915,N_8561,N_8471);
and U8916 (N_8916,N_8688,N_8446);
nor U8917 (N_8917,N_8630,N_8543);
nor U8918 (N_8918,N_8408,N_8611);
nor U8919 (N_8919,N_8634,N_8442);
or U8920 (N_8920,N_8470,N_8483);
nand U8921 (N_8921,N_8498,N_8672);
or U8922 (N_8922,N_8611,N_8423);
and U8923 (N_8923,N_8435,N_8630);
or U8924 (N_8924,N_8458,N_8672);
xnor U8925 (N_8925,N_8617,N_8468);
xor U8926 (N_8926,N_8586,N_8620);
nand U8927 (N_8927,N_8421,N_8529);
or U8928 (N_8928,N_8450,N_8476);
nor U8929 (N_8929,N_8540,N_8667);
nand U8930 (N_8930,N_8520,N_8505);
or U8931 (N_8931,N_8669,N_8471);
xor U8932 (N_8932,N_8668,N_8447);
xnor U8933 (N_8933,N_8462,N_8480);
and U8934 (N_8934,N_8488,N_8587);
or U8935 (N_8935,N_8448,N_8696);
nor U8936 (N_8936,N_8520,N_8548);
and U8937 (N_8937,N_8597,N_8401);
nor U8938 (N_8938,N_8574,N_8522);
and U8939 (N_8939,N_8418,N_8480);
nand U8940 (N_8940,N_8411,N_8480);
nand U8941 (N_8941,N_8473,N_8582);
or U8942 (N_8942,N_8427,N_8540);
or U8943 (N_8943,N_8583,N_8639);
and U8944 (N_8944,N_8408,N_8570);
nand U8945 (N_8945,N_8589,N_8605);
xnor U8946 (N_8946,N_8584,N_8480);
xor U8947 (N_8947,N_8436,N_8676);
and U8948 (N_8948,N_8528,N_8552);
nor U8949 (N_8949,N_8610,N_8582);
or U8950 (N_8950,N_8500,N_8431);
and U8951 (N_8951,N_8565,N_8567);
and U8952 (N_8952,N_8480,N_8624);
or U8953 (N_8953,N_8590,N_8562);
and U8954 (N_8954,N_8570,N_8633);
nor U8955 (N_8955,N_8476,N_8523);
xor U8956 (N_8956,N_8582,N_8499);
nand U8957 (N_8957,N_8508,N_8598);
xnor U8958 (N_8958,N_8606,N_8685);
or U8959 (N_8959,N_8511,N_8430);
nor U8960 (N_8960,N_8617,N_8487);
nor U8961 (N_8961,N_8650,N_8439);
nor U8962 (N_8962,N_8554,N_8650);
nor U8963 (N_8963,N_8653,N_8473);
nand U8964 (N_8964,N_8682,N_8483);
nor U8965 (N_8965,N_8581,N_8471);
or U8966 (N_8966,N_8474,N_8611);
or U8967 (N_8967,N_8469,N_8555);
nor U8968 (N_8968,N_8480,N_8558);
and U8969 (N_8969,N_8529,N_8462);
or U8970 (N_8970,N_8668,N_8692);
nor U8971 (N_8971,N_8689,N_8496);
or U8972 (N_8972,N_8472,N_8618);
nor U8973 (N_8973,N_8547,N_8657);
and U8974 (N_8974,N_8488,N_8465);
or U8975 (N_8975,N_8496,N_8627);
and U8976 (N_8976,N_8498,N_8441);
and U8977 (N_8977,N_8684,N_8445);
xnor U8978 (N_8978,N_8658,N_8678);
and U8979 (N_8979,N_8636,N_8502);
nor U8980 (N_8980,N_8423,N_8625);
or U8981 (N_8981,N_8545,N_8651);
xor U8982 (N_8982,N_8630,N_8653);
nand U8983 (N_8983,N_8448,N_8429);
and U8984 (N_8984,N_8600,N_8506);
or U8985 (N_8985,N_8478,N_8567);
and U8986 (N_8986,N_8680,N_8560);
xnor U8987 (N_8987,N_8402,N_8411);
nand U8988 (N_8988,N_8580,N_8418);
nor U8989 (N_8989,N_8402,N_8636);
nor U8990 (N_8990,N_8699,N_8563);
or U8991 (N_8991,N_8481,N_8685);
or U8992 (N_8992,N_8695,N_8648);
xnor U8993 (N_8993,N_8526,N_8669);
and U8994 (N_8994,N_8446,N_8641);
nor U8995 (N_8995,N_8610,N_8438);
or U8996 (N_8996,N_8508,N_8594);
nor U8997 (N_8997,N_8596,N_8663);
nor U8998 (N_8998,N_8639,N_8484);
and U8999 (N_8999,N_8508,N_8590);
nand U9000 (N_9000,N_8736,N_8705);
nor U9001 (N_9001,N_8886,N_8795);
nand U9002 (N_9002,N_8717,N_8992);
xnor U9003 (N_9003,N_8939,N_8990);
and U9004 (N_9004,N_8991,N_8942);
and U9005 (N_9005,N_8719,N_8732);
or U9006 (N_9006,N_8853,N_8781);
nand U9007 (N_9007,N_8811,N_8891);
or U9008 (N_9008,N_8801,N_8815);
and U9009 (N_9009,N_8807,N_8957);
or U9010 (N_9010,N_8924,N_8912);
and U9011 (N_9011,N_8978,N_8998);
nor U9012 (N_9012,N_8723,N_8704);
nand U9013 (N_9013,N_8779,N_8786);
xnor U9014 (N_9014,N_8973,N_8843);
nand U9015 (N_9015,N_8730,N_8819);
and U9016 (N_9016,N_8768,N_8989);
nand U9017 (N_9017,N_8933,N_8858);
nor U9018 (N_9018,N_8837,N_8767);
or U9019 (N_9019,N_8985,N_8970);
nor U9020 (N_9020,N_8983,N_8936);
or U9021 (N_9021,N_8851,N_8904);
nand U9022 (N_9022,N_8722,N_8804);
or U9023 (N_9023,N_8935,N_8889);
nor U9024 (N_9024,N_8824,N_8972);
nand U9025 (N_9025,N_8900,N_8757);
nand U9026 (N_9026,N_8981,N_8871);
or U9027 (N_9027,N_8910,N_8783);
or U9028 (N_9028,N_8741,N_8731);
or U9029 (N_9029,N_8729,N_8774);
xor U9030 (N_9030,N_8833,N_8735);
nor U9031 (N_9031,N_8840,N_8812);
and U9032 (N_9032,N_8802,N_8911);
and U9033 (N_9033,N_8790,N_8818);
and U9034 (N_9034,N_8969,N_8711);
and U9035 (N_9035,N_8895,N_8993);
nor U9036 (N_9036,N_8700,N_8964);
xnor U9037 (N_9037,N_8893,N_8852);
nand U9038 (N_9038,N_8808,N_8874);
or U9039 (N_9039,N_8763,N_8728);
or U9040 (N_9040,N_8997,N_8845);
and U9041 (N_9041,N_8965,N_8762);
or U9042 (N_9042,N_8913,N_8870);
and U9043 (N_9043,N_8953,N_8876);
nor U9044 (N_9044,N_8968,N_8785);
xor U9045 (N_9045,N_8944,N_8820);
and U9046 (N_9046,N_8756,N_8882);
nor U9047 (N_9047,N_8869,N_8842);
xnor U9048 (N_9048,N_8943,N_8707);
xnor U9049 (N_9049,N_8841,N_8794);
nor U9050 (N_9050,N_8923,N_8834);
nand U9051 (N_9051,N_8823,N_8960);
xnor U9052 (N_9052,N_8987,N_8919);
nor U9053 (N_9053,N_8878,N_8701);
and U9054 (N_9054,N_8772,N_8715);
and U9055 (N_9055,N_8927,N_8793);
and U9056 (N_9056,N_8879,N_8934);
nor U9057 (N_9057,N_8962,N_8784);
nor U9058 (N_9058,N_8721,N_8737);
xor U9059 (N_9059,N_8856,N_8855);
nand U9060 (N_9060,N_8996,N_8980);
and U9061 (N_9061,N_8847,N_8798);
nor U9062 (N_9062,N_8775,N_8850);
or U9063 (N_9063,N_8747,N_8930);
and U9064 (N_9064,N_8838,N_8931);
nand U9065 (N_9065,N_8748,N_8733);
nor U9066 (N_9066,N_8734,N_8988);
nand U9067 (N_9067,N_8865,N_8956);
or U9068 (N_9068,N_8765,N_8742);
xor U9069 (N_9069,N_8799,N_8776);
xnor U9070 (N_9070,N_8901,N_8976);
and U9071 (N_9071,N_8846,N_8894);
nand U9072 (N_9072,N_8849,N_8769);
or U9073 (N_9073,N_8884,N_8710);
and U9074 (N_9074,N_8803,N_8750);
xor U9075 (N_9075,N_8825,N_8921);
nand U9076 (N_9076,N_8753,N_8726);
and U9077 (N_9077,N_8863,N_8963);
xor U9078 (N_9078,N_8917,N_8961);
xor U9079 (N_9079,N_8826,N_8702);
and U9080 (N_9080,N_8787,N_8938);
nand U9081 (N_9081,N_8848,N_8809);
xnor U9082 (N_9082,N_8906,N_8760);
nand U9083 (N_9083,N_8885,N_8830);
and U9084 (N_9084,N_8745,N_8868);
or U9085 (N_9085,N_8971,N_8788);
and U9086 (N_9086,N_8982,N_8725);
xor U9087 (N_9087,N_8955,N_8881);
nand U9088 (N_9088,N_8718,N_8800);
or U9089 (N_9089,N_8810,N_8709);
nand U9090 (N_9090,N_8909,N_8951);
or U9091 (N_9091,N_8859,N_8797);
xnor U9092 (N_9092,N_8791,N_8892);
xnor U9093 (N_9093,N_8937,N_8862);
xor U9094 (N_9094,N_8975,N_8984);
and U9095 (N_9095,N_8905,N_8860);
nor U9096 (N_9096,N_8764,N_8727);
nand U9097 (N_9097,N_8780,N_8922);
nor U9098 (N_9098,N_8835,N_8925);
and U9099 (N_9099,N_8898,N_8873);
or U9100 (N_9100,N_8744,N_8857);
nand U9101 (N_9101,N_8806,N_8714);
or U9102 (N_9102,N_8887,N_8782);
or U9103 (N_9103,N_8954,N_8703);
and U9104 (N_9104,N_8754,N_8817);
or U9105 (N_9105,N_8949,N_8777);
nand U9106 (N_9106,N_8899,N_8914);
or U9107 (N_9107,N_8945,N_8896);
nor U9108 (N_9108,N_8720,N_8813);
nor U9109 (N_9109,N_8792,N_8883);
nand U9110 (N_9110,N_8816,N_8831);
or U9111 (N_9111,N_8920,N_8854);
nor U9112 (N_9112,N_8827,N_8716);
and U9113 (N_9113,N_8929,N_8867);
nand U9114 (N_9114,N_8759,N_8928);
or U9115 (N_9115,N_8789,N_8959);
and U9116 (N_9116,N_8941,N_8713);
xnor U9117 (N_9117,N_8844,N_8986);
xnor U9118 (N_9118,N_8828,N_8805);
and U9119 (N_9119,N_8712,N_8839);
and U9120 (N_9120,N_8773,N_8977);
xnor U9121 (N_9121,N_8740,N_8796);
nand U9122 (N_9122,N_8888,N_8761);
xor U9123 (N_9123,N_8708,N_8994);
and U9124 (N_9124,N_8932,N_8766);
nor U9125 (N_9125,N_8822,N_8755);
xor U9126 (N_9126,N_8967,N_8814);
and U9127 (N_9127,N_8770,N_8752);
or U9128 (N_9128,N_8903,N_8999);
and U9129 (N_9129,N_8958,N_8907);
or U9130 (N_9130,N_8771,N_8866);
and U9131 (N_9131,N_8880,N_8947);
and U9132 (N_9132,N_8821,N_8738);
nand U9133 (N_9133,N_8749,N_8974);
nand U9134 (N_9134,N_8940,N_8890);
nor U9135 (N_9135,N_8724,N_8778);
nand U9136 (N_9136,N_8872,N_8897);
nor U9137 (N_9137,N_8832,N_8916);
or U9138 (N_9138,N_8946,N_8751);
nor U9139 (N_9139,N_8915,N_8758);
and U9140 (N_9140,N_8902,N_8950);
nor U9141 (N_9141,N_8829,N_8864);
nand U9142 (N_9142,N_8861,N_8743);
and U9143 (N_9143,N_8908,N_8952);
or U9144 (N_9144,N_8918,N_8948);
or U9145 (N_9145,N_8746,N_8995);
nor U9146 (N_9146,N_8966,N_8979);
nand U9147 (N_9147,N_8706,N_8836);
or U9148 (N_9148,N_8875,N_8926);
and U9149 (N_9149,N_8877,N_8739);
or U9150 (N_9150,N_8880,N_8734);
nor U9151 (N_9151,N_8751,N_8810);
xnor U9152 (N_9152,N_8929,N_8794);
nand U9153 (N_9153,N_8864,N_8708);
nor U9154 (N_9154,N_8775,N_8829);
nand U9155 (N_9155,N_8925,N_8751);
nand U9156 (N_9156,N_8909,N_8786);
or U9157 (N_9157,N_8727,N_8817);
and U9158 (N_9158,N_8850,N_8804);
nor U9159 (N_9159,N_8962,N_8707);
and U9160 (N_9160,N_8786,N_8714);
nor U9161 (N_9161,N_8834,N_8933);
and U9162 (N_9162,N_8965,N_8905);
nand U9163 (N_9163,N_8823,N_8894);
xor U9164 (N_9164,N_8973,N_8757);
xnor U9165 (N_9165,N_8729,N_8823);
and U9166 (N_9166,N_8886,N_8726);
or U9167 (N_9167,N_8754,N_8910);
and U9168 (N_9168,N_8920,N_8771);
and U9169 (N_9169,N_8853,N_8901);
nor U9170 (N_9170,N_8983,N_8854);
or U9171 (N_9171,N_8866,N_8917);
nand U9172 (N_9172,N_8791,N_8811);
xnor U9173 (N_9173,N_8768,N_8934);
or U9174 (N_9174,N_8915,N_8764);
xnor U9175 (N_9175,N_8949,N_8962);
nor U9176 (N_9176,N_8954,N_8791);
xor U9177 (N_9177,N_8780,N_8738);
or U9178 (N_9178,N_8788,N_8933);
xnor U9179 (N_9179,N_8798,N_8852);
nand U9180 (N_9180,N_8943,N_8706);
nor U9181 (N_9181,N_8802,N_8813);
xnor U9182 (N_9182,N_8986,N_8738);
and U9183 (N_9183,N_8774,N_8757);
nor U9184 (N_9184,N_8927,N_8945);
or U9185 (N_9185,N_8741,N_8785);
and U9186 (N_9186,N_8862,N_8882);
or U9187 (N_9187,N_8771,N_8994);
xor U9188 (N_9188,N_8813,N_8778);
or U9189 (N_9189,N_8943,N_8894);
nand U9190 (N_9190,N_8867,N_8781);
nor U9191 (N_9191,N_8875,N_8824);
nor U9192 (N_9192,N_8732,N_8794);
nand U9193 (N_9193,N_8893,N_8912);
nand U9194 (N_9194,N_8743,N_8947);
or U9195 (N_9195,N_8714,N_8861);
or U9196 (N_9196,N_8710,N_8913);
or U9197 (N_9197,N_8751,N_8750);
nand U9198 (N_9198,N_8946,N_8983);
or U9199 (N_9199,N_8955,N_8958);
nand U9200 (N_9200,N_8925,N_8705);
nand U9201 (N_9201,N_8702,N_8812);
nor U9202 (N_9202,N_8906,N_8721);
nor U9203 (N_9203,N_8770,N_8822);
nor U9204 (N_9204,N_8771,N_8912);
or U9205 (N_9205,N_8772,N_8976);
nand U9206 (N_9206,N_8990,N_8947);
nand U9207 (N_9207,N_8724,N_8954);
or U9208 (N_9208,N_8940,N_8804);
nor U9209 (N_9209,N_8741,N_8943);
xnor U9210 (N_9210,N_8752,N_8798);
or U9211 (N_9211,N_8749,N_8938);
xor U9212 (N_9212,N_8773,N_8847);
or U9213 (N_9213,N_8843,N_8808);
xor U9214 (N_9214,N_8778,N_8894);
nor U9215 (N_9215,N_8795,N_8970);
nor U9216 (N_9216,N_8715,N_8738);
or U9217 (N_9217,N_8858,N_8709);
and U9218 (N_9218,N_8865,N_8922);
and U9219 (N_9219,N_8859,N_8798);
nor U9220 (N_9220,N_8702,N_8755);
and U9221 (N_9221,N_8852,N_8950);
and U9222 (N_9222,N_8971,N_8945);
nand U9223 (N_9223,N_8785,N_8978);
nor U9224 (N_9224,N_8898,N_8890);
and U9225 (N_9225,N_8778,N_8815);
nand U9226 (N_9226,N_8905,N_8777);
and U9227 (N_9227,N_8810,N_8717);
xor U9228 (N_9228,N_8949,N_8999);
nand U9229 (N_9229,N_8739,N_8988);
and U9230 (N_9230,N_8735,N_8988);
nand U9231 (N_9231,N_8995,N_8903);
nand U9232 (N_9232,N_8894,N_8910);
xnor U9233 (N_9233,N_8989,N_8723);
xnor U9234 (N_9234,N_8754,N_8947);
or U9235 (N_9235,N_8980,N_8840);
nor U9236 (N_9236,N_8822,N_8707);
or U9237 (N_9237,N_8722,N_8898);
and U9238 (N_9238,N_8865,N_8974);
or U9239 (N_9239,N_8948,N_8786);
or U9240 (N_9240,N_8910,N_8908);
nand U9241 (N_9241,N_8822,N_8915);
nand U9242 (N_9242,N_8900,N_8869);
and U9243 (N_9243,N_8974,N_8883);
xnor U9244 (N_9244,N_8976,N_8739);
xnor U9245 (N_9245,N_8788,N_8791);
and U9246 (N_9246,N_8704,N_8843);
or U9247 (N_9247,N_8721,N_8883);
nor U9248 (N_9248,N_8871,N_8735);
nand U9249 (N_9249,N_8953,N_8823);
and U9250 (N_9250,N_8794,N_8909);
or U9251 (N_9251,N_8789,N_8734);
and U9252 (N_9252,N_8869,N_8734);
or U9253 (N_9253,N_8790,N_8983);
nor U9254 (N_9254,N_8887,N_8839);
nor U9255 (N_9255,N_8716,N_8760);
and U9256 (N_9256,N_8971,N_8934);
nand U9257 (N_9257,N_8815,N_8822);
nor U9258 (N_9258,N_8809,N_8976);
xor U9259 (N_9259,N_8721,N_8846);
and U9260 (N_9260,N_8760,N_8819);
and U9261 (N_9261,N_8860,N_8994);
or U9262 (N_9262,N_8845,N_8946);
or U9263 (N_9263,N_8782,N_8810);
and U9264 (N_9264,N_8943,N_8788);
nand U9265 (N_9265,N_8896,N_8844);
or U9266 (N_9266,N_8714,N_8796);
and U9267 (N_9267,N_8765,N_8841);
nor U9268 (N_9268,N_8966,N_8760);
xnor U9269 (N_9269,N_8727,N_8771);
nand U9270 (N_9270,N_8855,N_8793);
nor U9271 (N_9271,N_8987,N_8973);
xor U9272 (N_9272,N_8887,N_8905);
nor U9273 (N_9273,N_8797,N_8831);
xor U9274 (N_9274,N_8942,N_8950);
nor U9275 (N_9275,N_8720,N_8984);
and U9276 (N_9276,N_8908,N_8773);
xor U9277 (N_9277,N_8916,N_8895);
or U9278 (N_9278,N_8804,N_8835);
or U9279 (N_9279,N_8984,N_8957);
nand U9280 (N_9280,N_8801,N_8769);
nand U9281 (N_9281,N_8898,N_8715);
nand U9282 (N_9282,N_8818,N_8841);
or U9283 (N_9283,N_8981,N_8844);
xor U9284 (N_9284,N_8703,N_8702);
nor U9285 (N_9285,N_8827,N_8977);
nand U9286 (N_9286,N_8719,N_8912);
and U9287 (N_9287,N_8884,N_8740);
or U9288 (N_9288,N_8837,N_8858);
and U9289 (N_9289,N_8753,N_8854);
nor U9290 (N_9290,N_8869,N_8875);
nand U9291 (N_9291,N_8974,N_8700);
and U9292 (N_9292,N_8931,N_8719);
nand U9293 (N_9293,N_8986,N_8975);
xnor U9294 (N_9294,N_8867,N_8764);
nor U9295 (N_9295,N_8957,N_8994);
and U9296 (N_9296,N_8713,N_8912);
nand U9297 (N_9297,N_8882,N_8884);
nor U9298 (N_9298,N_8919,N_8959);
nor U9299 (N_9299,N_8924,N_8734);
nand U9300 (N_9300,N_9238,N_9001);
xor U9301 (N_9301,N_9081,N_9107);
nor U9302 (N_9302,N_9009,N_9070);
xnor U9303 (N_9303,N_9297,N_9188);
or U9304 (N_9304,N_9292,N_9236);
nor U9305 (N_9305,N_9082,N_9088);
and U9306 (N_9306,N_9258,N_9167);
and U9307 (N_9307,N_9166,N_9117);
or U9308 (N_9308,N_9128,N_9155);
or U9309 (N_9309,N_9169,N_9220);
xnor U9310 (N_9310,N_9203,N_9273);
nand U9311 (N_9311,N_9071,N_9060);
and U9312 (N_9312,N_9296,N_9079);
nand U9313 (N_9313,N_9113,N_9294);
xor U9314 (N_9314,N_9014,N_9245);
nor U9315 (N_9315,N_9241,N_9231);
or U9316 (N_9316,N_9176,N_9265);
or U9317 (N_9317,N_9186,N_9073);
nor U9318 (N_9318,N_9227,N_9084);
and U9319 (N_9319,N_9183,N_9062);
nor U9320 (N_9320,N_9123,N_9051);
xor U9321 (N_9321,N_9067,N_9233);
nand U9322 (N_9322,N_9112,N_9223);
nor U9323 (N_9323,N_9216,N_9008);
nor U9324 (N_9324,N_9201,N_9029);
or U9325 (N_9325,N_9196,N_9246);
or U9326 (N_9326,N_9004,N_9281);
or U9327 (N_9327,N_9111,N_9106);
nor U9328 (N_9328,N_9030,N_9219);
and U9329 (N_9329,N_9198,N_9025);
nor U9330 (N_9330,N_9044,N_9141);
nor U9331 (N_9331,N_9157,N_9228);
nand U9332 (N_9332,N_9164,N_9287);
xnor U9333 (N_9333,N_9200,N_9115);
and U9334 (N_9334,N_9146,N_9269);
nor U9335 (N_9335,N_9126,N_9142);
nor U9336 (N_9336,N_9075,N_9197);
nor U9337 (N_9337,N_9251,N_9013);
nor U9338 (N_9338,N_9211,N_9256);
or U9339 (N_9339,N_9179,N_9119);
and U9340 (N_9340,N_9168,N_9077);
or U9341 (N_9341,N_9005,N_9208);
xnor U9342 (N_9342,N_9006,N_9063);
nand U9343 (N_9343,N_9074,N_9270);
nand U9344 (N_9344,N_9289,N_9272);
xor U9345 (N_9345,N_9140,N_9124);
or U9346 (N_9346,N_9138,N_9175);
xor U9347 (N_9347,N_9174,N_9259);
nand U9348 (N_9348,N_9143,N_9016);
nand U9349 (N_9349,N_9205,N_9047);
and U9350 (N_9350,N_9056,N_9280);
or U9351 (N_9351,N_9114,N_9226);
nand U9352 (N_9352,N_9087,N_9058);
or U9353 (N_9353,N_9007,N_9125);
nor U9354 (N_9354,N_9103,N_9210);
nor U9355 (N_9355,N_9178,N_9089);
nor U9356 (N_9356,N_9024,N_9012);
xnor U9357 (N_9357,N_9232,N_9086);
and U9358 (N_9358,N_9285,N_9261);
and U9359 (N_9359,N_9017,N_9116);
and U9360 (N_9360,N_9131,N_9181);
nand U9361 (N_9361,N_9028,N_9290);
xor U9362 (N_9362,N_9102,N_9221);
and U9363 (N_9363,N_9054,N_9298);
or U9364 (N_9364,N_9249,N_9096);
xnor U9365 (N_9365,N_9148,N_9254);
nor U9366 (N_9366,N_9121,N_9133);
xnor U9367 (N_9367,N_9078,N_9235);
nand U9368 (N_9368,N_9244,N_9043);
and U9369 (N_9369,N_9109,N_9118);
xnor U9370 (N_9370,N_9206,N_9120);
and U9371 (N_9371,N_9253,N_9020);
nand U9372 (N_9372,N_9100,N_9263);
nor U9373 (N_9373,N_9032,N_9215);
and U9374 (N_9374,N_9202,N_9291);
nand U9375 (N_9375,N_9271,N_9127);
xnor U9376 (N_9376,N_9094,N_9190);
or U9377 (N_9377,N_9003,N_9156);
nand U9378 (N_9378,N_9212,N_9098);
nor U9379 (N_9379,N_9171,N_9053);
and U9380 (N_9380,N_9042,N_9153);
nand U9381 (N_9381,N_9031,N_9173);
xor U9382 (N_9382,N_9237,N_9194);
and U9383 (N_9383,N_9260,N_9110);
and U9384 (N_9384,N_9192,N_9204);
nand U9385 (N_9385,N_9019,N_9209);
or U9386 (N_9386,N_9234,N_9161);
nor U9387 (N_9387,N_9274,N_9189);
nor U9388 (N_9388,N_9162,N_9105);
and U9389 (N_9389,N_9072,N_9275);
nand U9390 (N_9390,N_9160,N_9247);
nand U9391 (N_9391,N_9158,N_9187);
or U9392 (N_9392,N_9010,N_9000);
nand U9393 (N_9393,N_9191,N_9037);
xnor U9394 (N_9394,N_9276,N_9252);
or U9395 (N_9395,N_9027,N_9299);
nand U9396 (N_9396,N_9177,N_9182);
nand U9397 (N_9397,N_9093,N_9057);
nand U9398 (N_9398,N_9050,N_9250);
xor U9399 (N_9399,N_9277,N_9264);
or U9400 (N_9400,N_9243,N_9195);
and U9401 (N_9401,N_9268,N_9033);
and U9402 (N_9402,N_9257,N_9026);
xnor U9403 (N_9403,N_9217,N_9130);
or U9404 (N_9404,N_9122,N_9021);
nor U9405 (N_9405,N_9242,N_9076);
and U9406 (N_9406,N_9011,N_9065);
and U9407 (N_9407,N_9092,N_9214);
or U9408 (N_9408,N_9136,N_9288);
nor U9409 (N_9409,N_9267,N_9036);
or U9410 (N_9410,N_9180,N_9097);
nand U9411 (N_9411,N_9279,N_9207);
xor U9412 (N_9412,N_9066,N_9080);
nand U9413 (N_9413,N_9163,N_9150);
nor U9414 (N_9414,N_9152,N_9135);
and U9415 (N_9415,N_9040,N_9023);
or U9416 (N_9416,N_9048,N_9049);
nor U9417 (N_9417,N_9295,N_9230);
nor U9418 (N_9418,N_9283,N_9213);
nand U9419 (N_9419,N_9059,N_9278);
or U9420 (N_9420,N_9159,N_9018);
or U9421 (N_9421,N_9284,N_9239);
nor U9422 (N_9422,N_9108,N_9095);
nor U9423 (N_9423,N_9022,N_9090);
and U9424 (N_9424,N_9240,N_9035);
nand U9425 (N_9425,N_9085,N_9099);
and U9426 (N_9426,N_9229,N_9132);
xor U9427 (N_9427,N_9282,N_9045);
xor U9428 (N_9428,N_9069,N_9055);
or U9429 (N_9429,N_9149,N_9137);
and U9430 (N_9430,N_9129,N_9052);
and U9431 (N_9431,N_9061,N_9224);
or U9432 (N_9432,N_9139,N_9151);
nand U9433 (N_9433,N_9064,N_9145);
or U9434 (N_9434,N_9068,N_9104);
xor U9435 (N_9435,N_9193,N_9199);
nor U9436 (N_9436,N_9248,N_9218);
or U9437 (N_9437,N_9165,N_9185);
xor U9438 (N_9438,N_9034,N_9091);
or U9439 (N_9439,N_9154,N_9170);
xor U9440 (N_9440,N_9039,N_9184);
and U9441 (N_9441,N_9083,N_9002);
nor U9442 (N_9442,N_9038,N_9293);
nor U9443 (N_9443,N_9101,N_9222);
nor U9444 (N_9444,N_9172,N_9147);
and U9445 (N_9445,N_9046,N_9266);
or U9446 (N_9446,N_9041,N_9262);
xor U9447 (N_9447,N_9286,N_9225);
nor U9448 (N_9448,N_9015,N_9134);
xor U9449 (N_9449,N_9255,N_9144);
nand U9450 (N_9450,N_9126,N_9282);
xnor U9451 (N_9451,N_9029,N_9123);
nand U9452 (N_9452,N_9104,N_9285);
or U9453 (N_9453,N_9002,N_9224);
xnor U9454 (N_9454,N_9207,N_9070);
or U9455 (N_9455,N_9189,N_9058);
or U9456 (N_9456,N_9025,N_9055);
or U9457 (N_9457,N_9258,N_9294);
nand U9458 (N_9458,N_9144,N_9106);
xor U9459 (N_9459,N_9112,N_9206);
nand U9460 (N_9460,N_9005,N_9022);
nor U9461 (N_9461,N_9109,N_9024);
nor U9462 (N_9462,N_9248,N_9266);
nor U9463 (N_9463,N_9270,N_9102);
or U9464 (N_9464,N_9056,N_9209);
or U9465 (N_9465,N_9232,N_9284);
nor U9466 (N_9466,N_9073,N_9065);
nor U9467 (N_9467,N_9152,N_9134);
or U9468 (N_9468,N_9232,N_9157);
and U9469 (N_9469,N_9213,N_9078);
nand U9470 (N_9470,N_9288,N_9153);
or U9471 (N_9471,N_9150,N_9279);
nand U9472 (N_9472,N_9054,N_9270);
nand U9473 (N_9473,N_9003,N_9015);
xor U9474 (N_9474,N_9133,N_9256);
nor U9475 (N_9475,N_9020,N_9097);
or U9476 (N_9476,N_9200,N_9295);
and U9477 (N_9477,N_9122,N_9267);
and U9478 (N_9478,N_9023,N_9078);
and U9479 (N_9479,N_9165,N_9057);
and U9480 (N_9480,N_9130,N_9292);
or U9481 (N_9481,N_9238,N_9011);
and U9482 (N_9482,N_9247,N_9290);
nand U9483 (N_9483,N_9162,N_9159);
nor U9484 (N_9484,N_9038,N_9122);
and U9485 (N_9485,N_9076,N_9074);
xor U9486 (N_9486,N_9105,N_9118);
nor U9487 (N_9487,N_9046,N_9179);
and U9488 (N_9488,N_9295,N_9097);
nor U9489 (N_9489,N_9270,N_9243);
and U9490 (N_9490,N_9071,N_9295);
xor U9491 (N_9491,N_9045,N_9245);
xor U9492 (N_9492,N_9244,N_9221);
xor U9493 (N_9493,N_9131,N_9045);
or U9494 (N_9494,N_9188,N_9141);
nand U9495 (N_9495,N_9224,N_9291);
nand U9496 (N_9496,N_9090,N_9298);
nand U9497 (N_9497,N_9172,N_9195);
or U9498 (N_9498,N_9065,N_9041);
and U9499 (N_9499,N_9273,N_9276);
and U9500 (N_9500,N_9288,N_9066);
or U9501 (N_9501,N_9041,N_9261);
nand U9502 (N_9502,N_9166,N_9032);
nor U9503 (N_9503,N_9080,N_9221);
xnor U9504 (N_9504,N_9104,N_9034);
and U9505 (N_9505,N_9199,N_9239);
nand U9506 (N_9506,N_9178,N_9064);
or U9507 (N_9507,N_9058,N_9298);
nand U9508 (N_9508,N_9282,N_9285);
xor U9509 (N_9509,N_9048,N_9160);
and U9510 (N_9510,N_9247,N_9282);
or U9511 (N_9511,N_9015,N_9235);
and U9512 (N_9512,N_9091,N_9127);
and U9513 (N_9513,N_9066,N_9282);
nand U9514 (N_9514,N_9223,N_9269);
nand U9515 (N_9515,N_9027,N_9063);
and U9516 (N_9516,N_9007,N_9068);
nand U9517 (N_9517,N_9119,N_9283);
nand U9518 (N_9518,N_9105,N_9095);
xor U9519 (N_9519,N_9227,N_9297);
xnor U9520 (N_9520,N_9216,N_9298);
or U9521 (N_9521,N_9248,N_9017);
nor U9522 (N_9522,N_9164,N_9288);
xnor U9523 (N_9523,N_9007,N_9071);
nor U9524 (N_9524,N_9004,N_9192);
xnor U9525 (N_9525,N_9284,N_9032);
and U9526 (N_9526,N_9290,N_9156);
or U9527 (N_9527,N_9159,N_9163);
or U9528 (N_9528,N_9059,N_9219);
nand U9529 (N_9529,N_9287,N_9040);
nor U9530 (N_9530,N_9026,N_9282);
nor U9531 (N_9531,N_9067,N_9169);
nor U9532 (N_9532,N_9170,N_9178);
nor U9533 (N_9533,N_9093,N_9130);
or U9534 (N_9534,N_9168,N_9115);
nand U9535 (N_9535,N_9212,N_9059);
or U9536 (N_9536,N_9089,N_9275);
nor U9537 (N_9537,N_9085,N_9002);
xnor U9538 (N_9538,N_9154,N_9000);
nand U9539 (N_9539,N_9029,N_9152);
nor U9540 (N_9540,N_9108,N_9079);
nand U9541 (N_9541,N_9198,N_9045);
xor U9542 (N_9542,N_9242,N_9140);
or U9543 (N_9543,N_9244,N_9023);
nor U9544 (N_9544,N_9229,N_9278);
nor U9545 (N_9545,N_9244,N_9179);
nand U9546 (N_9546,N_9166,N_9077);
nor U9547 (N_9547,N_9137,N_9036);
nor U9548 (N_9548,N_9183,N_9012);
nand U9549 (N_9549,N_9103,N_9170);
nor U9550 (N_9550,N_9142,N_9160);
xor U9551 (N_9551,N_9061,N_9059);
nor U9552 (N_9552,N_9072,N_9053);
or U9553 (N_9553,N_9046,N_9290);
or U9554 (N_9554,N_9116,N_9296);
or U9555 (N_9555,N_9069,N_9060);
and U9556 (N_9556,N_9143,N_9230);
or U9557 (N_9557,N_9106,N_9158);
or U9558 (N_9558,N_9092,N_9116);
xnor U9559 (N_9559,N_9190,N_9131);
xor U9560 (N_9560,N_9107,N_9090);
or U9561 (N_9561,N_9081,N_9187);
or U9562 (N_9562,N_9279,N_9199);
and U9563 (N_9563,N_9211,N_9089);
nor U9564 (N_9564,N_9128,N_9188);
nor U9565 (N_9565,N_9224,N_9179);
nor U9566 (N_9566,N_9233,N_9109);
nand U9567 (N_9567,N_9099,N_9168);
xor U9568 (N_9568,N_9176,N_9187);
xnor U9569 (N_9569,N_9265,N_9056);
or U9570 (N_9570,N_9074,N_9183);
xor U9571 (N_9571,N_9235,N_9198);
nand U9572 (N_9572,N_9137,N_9197);
and U9573 (N_9573,N_9271,N_9249);
or U9574 (N_9574,N_9010,N_9223);
and U9575 (N_9575,N_9048,N_9011);
nand U9576 (N_9576,N_9289,N_9155);
xor U9577 (N_9577,N_9191,N_9035);
nand U9578 (N_9578,N_9186,N_9232);
and U9579 (N_9579,N_9063,N_9013);
xor U9580 (N_9580,N_9196,N_9102);
and U9581 (N_9581,N_9065,N_9172);
xor U9582 (N_9582,N_9270,N_9002);
nor U9583 (N_9583,N_9073,N_9213);
nand U9584 (N_9584,N_9057,N_9198);
nor U9585 (N_9585,N_9268,N_9058);
and U9586 (N_9586,N_9176,N_9101);
and U9587 (N_9587,N_9075,N_9142);
nand U9588 (N_9588,N_9165,N_9174);
xnor U9589 (N_9589,N_9188,N_9172);
nand U9590 (N_9590,N_9043,N_9232);
or U9591 (N_9591,N_9069,N_9052);
or U9592 (N_9592,N_9022,N_9271);
nor U9593 (N_9593,N_9118,N_9266);
nand U9594 (N_9594,N_9163,N_9289);
nand U9595 (N_9595,N_9155,N_9284);
xor U9596 (N_9596,N_9017,N_9104);
nand U9597 (N_9597,N_9238,N_9236);
nand U9598 (N_9598,N_9188,N_9222);
and U9599 (N_9599,N_9043,N_9075);
and U9600 (N_9600,N_9579,N_9576);
xnor U9601 (N_9601,N_9459,N_9553);
nand U9602 (N_9602,N_9414,N_9425);
and U9603 (N_9603,N_9389,N_9448);
xnor U9604 (N_9604,N_9497,N_9421);
xor U9605 (N_9605,N_9572,N_9442);
nor U9606 (N_9606,N_9557,N_9368);
nor U9607 (N_9607,N_9565,N_9312);
and U9608 (N_9608,N_9470,N_9570);
and U9609 (N_9609,N_9371,N_9452);
xor U9610 (N_9610,N_9357,N_9303);
or U9611 (N_9611,N_9339,N_9592);
nor U9612 (N_9612,N_9411,N_9590);
and U9613 (N_9613,N_9443,N_9372);
or U9614 (N_9614,N_9410,N_9597);
and U9615 (N_9615,N_9507,N_9511);
nor U9616 (N_9616,N_9323,N_9340);
and U9617 (N_9617,N_9502,N_9439);
xnor U9618 (N_9618,N_9310,N_9516);
or U9619 (N_9619,N_9462,N_9466);
xnor U9620 (N_9620,N_9324,N_9517);
or U9621 (N_9621,N_9495,N_9307);
and U9622 (N_9622,N_9444,N_9388);
nor U9623 (N_9623,N_9467,N_9407);
and U9624 (N_9624,N_9583,N_9377);
nand U9625 (N_9625,N_9413,N_9376);
nor U9626 (N_9626,N_9496,N_9363);
or U9627 (N_9627,N_9447,N_9539);
or U9628 (N_9628,N_9374,N_9334);
or U9629 (N_9629,N_9544,N_9332);
xor U9630 (N_9630,N_9586,N_9370);
nand U9631 (N_9631,N_9355,N_9529);
nor U9632 (N_9632,N_9518,N_9533);
nor U9633 (N_9633,N_9338,N_9432);
nor U9634 (N_9634,N_9541,N_9362);
xnor U9635 (N_9635,N_9306,N_9395);
nor U9636 (N_9636,N_9598,N_9406);
and U9637 (N_9637,N_9397,N_9361);
nand U9638 (N_9638,N_9385,N_9418);
nor U9639 (N_9639,N_9559,N_9500);
xnor U9640 (N_9640,N_9348,N_9480);
and U9641 (N_9641,N_9350,N_9580);
xor U9642 (N_9642,N_9409,N_9364);
and U9643 (N_9643,N_9524,N_9486);
xor U9644 (N_9644,N_9562,N_9584);
or U9645 (N_9645,N_9322,N_9531);
nand U9646 (N_9646,N_9532,N_9551);
xnor U9647 (N_9647,N_9594,N_9352);
and U9648 (N_9648,N_9316,N_9542);
and U9649 (N_9649,N_9429,N_9346);
and U9650 (N_9650,N_9521,N_9547);
and U9651 (N_9651,N_9564,N_9506);
nor U9652 (N_9652,N_9420,N_9481);
or U9653 (N_9653,N_9373,N_9479);
and U9654 (N_9654,N_9314,N_9461);
and U9655 (N_9655,N_9484,N_9379);
xor U9656 (N_9656,N_9560,N_9319);
xnor U9657 (N_9657,N_9440,N_9555);
or U9658 (N_9658,N_9499,N_9434);
and U9659 (N_9659,N_9399,N_9475);
xnor U9660 (N_9660,N_9549,N_9454);
nor U9661 (N_9661,N_9522,N_9577);
nand U9662 (N_9662,N_9417,N_9477);
or U9663 (N_9663,N_9330,N_9599);
xor U9664 (N_9664,N_9453,N_9327);
nand U9665 (N_9665,N_9311,N_9302);
and U9666 (N_9666,N_9498,N_9589);
nand U9667 (N_9667,N_9527,N_9463);
and U9668 (N_9668,N_9438,N_9483);
nor U9669 (N_9669,N_9501,N_9424);
and U9670 (N_9670,N_9416,N_9456);
nor U9671 (N_9671,N_9471,N_9445);
and U9672 (N_9672,N_9404,N_9573);
nor U9673 (N_9673,N_9490,N_9568);
and U9674 (N_9674,N_9489,N_9578);
nand U9675 (N_9675,N_9386,N_9505);
or U9676 (N_9676,N_9315,N_9582);
xnor U9677 (N_9677,N_9367,N_9353);
nand U9678 (N_9678,N_9396,N_9530);
nor U9679 (N_9679,N_9535,N_9394);
nor U9680 (N_9680,N_9405,N_9308);
nand U9681 (N_9681,N_9476,N_9423);
or U9682 (N_9682,N_9342,N_9528);
nor U9683 (N_9683,N_9400,N_9335);
and U9684 (N_9684,N_9366,N_9493);
or U9685 (N_9685,N_9369,N_9333);
nor U9686 (N_9686,N_9548,N_9300);
nor U9687 (N_9687,N_9356,N_9343);
nor U9688 (N_9688,N_9510,N_9581);
nor U9689 (N_9689,N_9523,N_9391);
nor U9690 (N_9690,N_9354,N_9545);
nand U9691 (N_9691,N_9422,N_9464);
and U9692 (N_9692,N_9537,N_9474);
nor U9693 (N_9693,N_9450,N_9345);
nand U9694 (N_9694,N_9383,N_9328);
nor U9695 (N_9695,N_9550,N_9558);
nand U9696 (N_9696,N_9384,N_9381);
or U9697 (N_9697,N_9556,N_9344);
xor U9698 (N_9698,N_9575,N_9401);
or U9699 (N_9699,N_9419,N_9596);
nor U9700 (N_9700,N_9441,N_9359);
or U9701 (N_9701,N_9321,N_9593);
nor U9702 (N_9702,N_9472,N_9437);
and U9703 (N_9703,N_9378,N_9552);
and U9704 (N_9704,N_9478,N_9318);
and U9705 (N_9705,N_9554,N_9536);
xnor U9706 (N_9706,N_9341,N_9387);
nand U9707 (N_9707,N_9426,N_9504);
nor U9708 (N_9708,N_9513,N_9431);
nor U9709 (N_9709,N_9512,N_9412);
xnor U9710 (N_9710,N_9543,N_9465);
nand U9711 (N_9711,N_9309,N_9473);
xor U9712 (N_9712,N_9313,N_9569);
xor U9713 (N_9713,N_9514,N_9337);
xor U9714 (N_9714,N_9415,N_9520);
or U9715 (N_9715,N_9561,N_9455);
nand U9716 (N_9716,N_9390,N_9403);
or U9717 (N_9717,N_9430,N_9492);
nand U9718 (N_9718,N_9317,N_9457);
nor U9719 (N_9719,N_9358,N_9408);
nand U9720 (N_9720,N_9538,N_9347);
nand U9721 (N_9721,N_9451,N_9574);
and U9722 (N_9722,N_9380,N_9460);
nor U9723 (N_9723,N_9587,N_9546);
nor U9724 (N_9724,N_9508,N_9349);
and U9725 (N_9725,N_9382,N_9433);
or U9726 (N_9726,N_9436,N_9428);
xnor U9727 (N_9727,N_9304,N_9360);
nand U9728 (N_9728,N_9365,N_9458);
nand U9729 (N_9729,N_9427,N_9301);
and U9730 (N_9730,N_9540,N_9595);
xor U9731 (N_9731,N_9534,N_9487);
nand U9732 (N_9732,N_9329,N_9526);
nand U9733 (N_9733,N_9326,N_9567);
and U9734 (N_9734,N_9402,N_9336);
or U9735 (N_9735,N_9585,N_9525);
or U9736 (N_9736,N_9488,N_9588);
xnor U9737 (N_9737,N_9566,N_9325);
nand U9738 (N_9738,N_9398,N_9591);
nand U9739 (N_9739,N_9519,N_9393);
or U9740 (N_9740,N_9331,N_9509);
and U9741 (N_9741,N_9468,N_9392);
or U9742 (N_9742,N_9503,N_9491);
and U9743 (N_9743,N_9482,N_9320);
or U9744 (N_9744,N_9515,N_9446);
nor U9745 (N_9745,N_9494,N_9375);
nand U9746 (N_9746,N_9435,N_9571);
xor U9747 (N_9747,N_9485,N_9351);
nand U9748 (N_9748,N_9469,N_9449);
nand U9749 (N_9749,N_9305,N_9563);
and U9750 (N_9750,N_9464,N_9321);
xor U9751 (N_9751,N_9397,N_9313);
nand U9752 (N_9752,N_9421,N_9357);
nor U9753 (N_9753,N_9372,N_9571);
nand U9754 (N_9754,N_9447,N_9367);
or U9755 (N_9755,N_9332,N_9307);
nor U9756 (N_9756,N_9426,N_9525);
or U9757 (N_9757,N_9345,N_9406);
or U9758 (N_9758,N_9301,N_9409);
xnor U9759 (N_9759,N_9447,N_9488);
nor U9760 (N_9760,N_9577,N_9386);
nand U9761 (N_9761,N_9531,N_9352);
nand U9762 (N_9762,N_9340,N_9544);
nor U9763 (N_9763,N_9535,N_9505);
xnor U9764 (N_9764,N_9469,N_9360);
and U9765 (N_9765,N_9567,N_9438);
and U9766 (N_9766,N_9311,N_9423);
and U9767 (N_9767,N_9406,N_9344);
and U9768 (N_9768,N_9343,N_9425);
nand U9769 (N_9769,N_9462,N_9473);
and U9770 (N_9770,N_9443,N_9470);
xor U9771 (N_9771,N_9453,N_9526);
and U9772 (N_9772,N_9576,N_9564);
nand U9773 (N_9773,N_9364,N_9441);
or U9774 (N_9774,N_9390,N_9324);
and U9775 (N_9775,N_9388,N_9518);
and U9776 (N_9776,N_9560,N_9433);
nor U9777 (N_9777,N_9350,N_9324);
nor U9778 (N_9778,N_9359,N_9513);
xnor U9779 (N_9779,N_9450,N_9312);
xnor U9780 (N_9780,N_9445,N_9389);
nand U9781 (N_9781,N_9480,N_9546);
xnor U9782 (N_9782,N_9335,N_9446);
or U9783 (N_9783,N_9323,N_9438);
or U9784 (N_9784,N_9494,N_9432);
nor U9785 (N_9785,N_9407,N_9390);
xor U9786 (N_9786,N_9426,N_9486);
xnor U9787 (N_9787,N_9579,N_9435);
nor U9788 (N_9788,N_9380,N_9382);
xnor U9789 (N_9789,N_9435,N_9364);
nand U9790 (N_9790,N_9595,N_9583);
xor U9791 (N_9791,N_9473,N_9496);
xor U9792 (N_9792,N_9560,N_9527);
xnor U9793 (N_9793,N_9415,N_9331);
nor U9794 (N_9794,N_9491,N_9481);
nand U9795 (N_9795,N_9410,N_9536);
xor U9796 (N_9796,N_9523,N_9587);
xor U9797 (N_9797,N_9374,N_9337);
nand U9798 (N_9798,N_9547,N_9442);
or U9799 (N_9799,N_9487,N_9372);
nor U9800 (N_9800,N_9390,N_9469);
nor U9801 (N_9801,N_9495,N_9587);
and U9802 (N_9802,N_9323,N_9328);
xor U9803 (N_9803,N_9494,N_9455);
xor U9804 (N_9804,N_9389,N_9324);
and U9805 (N_9805,N_9422,N_9507);
xnor U9806 (N_9806,N_9377,N_9523);
nand U9807 (N_9807,N_9306,N_9457);
or U9808 (N_9808,N_9578,N_9539);
nor U9809 (N_9809,N_9340,N_9596);
nand U9810 (N_9810,N_9391,N_9520);
xor U9811 (N_9811,N_9484,N_9560);
nor U9812 (N_9812,N_9474,N_9448);
and U9813 (N_9813,N_9454,N_9555);
or U9814 (N_9814,N_9533,N_9361);
or U9815 (N_9815,N_9488,N_9326);
xnor U9816 (N_9816,N_9364,N_9389);
and U9817 (N_9817,N_9454,N_9325);
nand U9818 (N_9818,N_9436,N_9442);
and U9819 (N_9819,N_9370,N_9561);
and U9820 (N_9820,N_9384,N_9567);
xor U9821 (N_9821,N_9498,N_9431);
nand U9822 (N_9822,N_9538,N_9582);
nand U9823 (N_9823,N_9586,N_9478);
or U9824 (N_9824,N_9524,N_9342);
and U9825 (N_9825,N_9586,N_9333);
or U9826 (N_9826,N_9376,N_9434);
and U9827 (N_9827,N_9365,N_9576);
or U9828 (N_9828,N_9503,N_9368);
and U9829 (N_9829,N_9491,N_9432);
and U9830 (N_9830,N_9310,N_9443);
nor U9831 (N_9831,N_9369,N_9512);
nand U9832 (N_9832,N_9357,N_9317);
nor U9833 (N_9833,N_9451,N_9584);
nor U9834 (N_9834,N_9462,N_9434);
nand U9835 (N_9835,N_9403,N_9357);
xor U9836 (N_9836,N_9558,N_9577);
nor U9837 (N_9837,N_9483,N_9348);
or U9838 (N_9838,N_9579,N_9527);
xor U9839 (N_9839,N_9358,N_9444);
and U9840 (N_9840,N_9327,N_9410);
nand U9841 (N_9841,N_9381,N_9583);
and U9842 (N_9842,N_9425,N_9550);
nor U9843 (N_9843,N_9401,N_9583);
nand U9844 (N_9844,N_9325,N_9414);
or U9845 (N_9845,N_9340,N_9322);
or U9846 (N_9846,N_9361,N_9589);
nor U9847 (N_9847,N_9477,N_9469);
xor U9848 (N_9848,N_9442,N_9404);
or U9849 (N_9849,N_9576,N_9364);
and U9850 (N_9850,N_9576,N_9397);
and U9851 (N_9851,N_9502,N_9305);
nor U9852 (N_9852,N_9489,N_9586);
xor U9853 (N_9853,N_9300,N_9499);
xnor U9854 (N_9854,N_9457,N_9300);
and U9855 (N_9855,N_9583,N_9403);
and U9856 (N_9856,N_9442,N_9599);
nand U9857 (N_9857,N_9553,N_9597);
xnor U9858 (N_9858,N_9430,N_9330);
nand U9859 (N_9859,N_9349,N_9412);
and U9860 (N_9860,N_9315,N_9360);
or U9861 (N_9861,N_9407,N_9417);
nand U9862 (N_9862,N_9500,N_9522);
xor U9863 (N_9863,N_9467,N_9400);
nand U9864 (N_9864,N_9379,N_9359);
and U9865 (N_9865,N_9543,N_9365);
nor U9866 (N_9866,N_9596,N_9530);
nor U9867 (N_9867,N_9407,N_9496);
nand U9868 (N_9868,N_9526,N_9534);
nor U9869 (N_9869,N_9569,N_9474);
or U9870 (N_9870,N_9553,N_9526);
or U9871 (N_9871,N_9469,N_9321);
nand U9872 (N_9872,N_9369,N_9487);
xor U9873 (N_9873,N_9404,N_9422);
nand U9874 (N_9874,N_9305,N_9595);
or U9875 (N_9875,N_9477,N_9563);
nor U9876 (N_9876,N_9458,N_9596);
nor U9877 (N_9877,N_9355,N_9316);
or U9878 (N_9878,N_9397,N_9587);
nor U9879 (N_9879,N_9403,N_9479);
xor U9880 (N_9880,N_9446,N_9440);
nor U9881 (N_9881,N_9543,N_9482);
or U9882 (N_9882,N_9348,N_9326);
nand U9883 (N_9883,N_9472,N_9511);
or U9884 (N_9884,N_9556,N_9345);
xnor U9885 (N_9885,N_9537,N_9373);
nor U9886 (N_9886,N_9482,N_9578);
nand U9887 (N_9887,N_9429,N_9472);
xor U9888 (N_9888,N_9503,N_9385);
nor U9889 (N_9889,N_9411,N_9594);
and U9890 (N_9890,N_9420,N_9463);
nor U9891 (N_9891,N_9463,N_9345);
xor U9892 (N_9892,N_9415,N_9445);
or U9893 (N_9893,N_9324,N_9379);
nor U9894 (N_9894,N_9591,N_9353);
or U9895 (N_9895,N_9541,N_9396);
nor U9896 (N_9896,N_9581,N_9477);
nand U9897 (N_9897,N_9346,N_9479);
nor U9898 (N_9898,N_9581,N_9414);
xnor U9899 (N_9899,N_9388,N_9436);
nand U9900 (N_9900,N_9639,N_9830);
and U9901 (N_9901,N_9844,N_9877);
nand U9902 (N_9902,N_9689,N_9737);
nor U9903 (N_9903,N_9703,N_9768);
xor U9904 (N_9904,N_9808,N_9848);
nor U9905 (N_9905,N_9731,N_9748);
or U9906 (N_9906,N_9684,N_9774);
and U9907 (N_9907,N_9632,N_9734);
nor U9908 (N_9908,N_9652,N_9716);
or U9909 (N_9909,N_9681,N_9875);
xor U9910 (N_9910,N_9701,N_9710);
nand U9911 (N_9911,N_9854,N_9725);
or U9912 (N_9912,N_9658,N_9866);
nand U9913 (N_9913,N_9800,N_9787);
nand U9914 (N_9914,N_9894,N_9745);
or U9915 (N_9915,N_9782,N_9872);
nand U9916 (N_9916,N_9620,N_9727);
nand U9917 (N_9917,N_9677,N_9751);
nor U9918 (N_9918,N_9646,N_9899);
nor U9919 (N_9919,N_9694,N_9799);
or U9920 (N_9920,N_9649,N_9680);
and U9921 (N_9921,N_9753,N_9766);
xor U9922 (N_9922,N_9641,N_9744);
xnor U9923 (N_9923,N_9823,N_9874);
xnor U9924 (N_9924,N_9780,N_9818);
nor U9925 (N_9925,N_9837,N_9869);
or U9926 (N_9926,N_9765,N_9759);
and U9927 (N_9927,N_9806,N_9674);
nor U9928 (N_9928,N_9855,N_9643);
or U9929 (N_9929,N_9749,N_9743);
or U9930 (N_9930,N_9802,N_9856);
and U9931 (N_9931,N_9746,N_9878);
xnor U9932 (N_9932,N_9757,N_9690);
nor U9933 (N_9933,N_9608,N_9688);
nand U9934 (N_9934,N_9756,N_9871);
nand U9935 (N_9935,N_9668,N_9648);
nand U9936 (N_9936,N_9772,N_9807);
xor U9937 (N_9937,N_9687,N_9650);
nor U9938 (N_9938,N_9676,N_9885);
nand U9939 (N_9939,N_9637,N_9662);
nor U9940 (N_9940,N_9600,N_9669);
xnor U9941 (N_9941,N_9794,N_9859);
nor U9942 (N_9942,N_9758,N_9798);
or U9943 (N_9943,N_9776,N_9860);
or U9944 (N_9944,N_9773,N_9699);
xor U9945 (N_9945,N_9867,N_9720);
or U9946 (N_9946,N_9602,N_9609);
nand U9947 (N_9947,N_9863,N_9730);
xnor U9948 (N_9948,N_9616,N_9812);
and U9949 (N_9949,N_9835,N_9685);
nor U9950 (N_9950,N_9660,N_9884);
or U9951 (N_9951,N_9709,N_9706);
nand U9952 (N_9952,N_9811,N_9849);
or U9953 (N_9953,N_9656,N_9777);
and U9954 (N_9954,N_9850,N_9796);
or U9955 (N_9955,N_9740,N_9624);
or U9956 (N_9956,N_9612,N_9779);
and U9957 (N_9957,N_9852,N_9733);
and U9958 (N_9958,N_9864,N_9630);
xor U9959 (N_9959,N_9892,N_9728);
and U9960 (N_9960,N_9771,N_9718);
or U9961 (N_9961,N_9761,N_9770);
nor U9962 (N_9962,N_9722,N_9832);
and U9963 (N_9963,N_9791,N_9789);
and U9964 (N_9964,N_9805,N_9784);
nor U9965 (N_9965,N_9762,N_9895);
nor U9966 (N_9966,N_9673,N_9755);
nand U9967 (N_9967,N_9611,N_9619);
nand U9968 (N_9968,N_9801,N_9723);
and U9969 (N_9969,N_9814,N_9605);
nand U9970 (N_9970,N_9691,N_9678);
nand U9971 (N_9971,N_9767,N_9741);
or U9972 (N_9972,N_9781,N_9702);
nor U9973 (N_9973,N_9713,N_9626);
and U9974 (N_9974,N_9833,N_9888);
or U9975 (N_9975,N_9868,N_9786);
and U9976 (N_9976,N_9829,N_9627);
and U9977 (N_9977,N_9613,N_9695);
nand U9978 (N_9978,N_9655,N_9657);
xor U9979 (N_9979,N_9838,N_9622);
xnor U9980 (N_9980,N_9826,N_9634);
and U9981 (N_9981,N_9631,N_9845);
nor U9982 (N_9982,N_9846,N_9865);
and U9983 (N_9983,N_9760,N_9642);
or U9984 (N_9984,N_9831,N_9752);
and U9985 (N_9985,N_9711,N_9819);
and U9986 (N_9986,N_9862,N_9610);
nor U9987 (N_9987,N_9636,N_9738);
nor U9988 (N_9988,N_9742,N_9842);
xnor U9989 (N_9989,N_9825,N_9769);
or U9990 (N_9990,N_9783,N_9893);
nand U9991 (N_9991,N_9654,N_9890);
nand U9992 (N_9992,N_9778,N_9601);
and U9993 (N_9993,N_9763,N_9841);
xnor U9994 (N_9994,N_9827,N_9675);
or U9995 (N_9995,N_9793,N_9615);
and U9996 (N_9996,N_9853,N_9617);
xnor U9997 (N_9997,N_9698,N_9614);
nand U9998 (N_9998,N_9635,N_9876);
or U9999 (N_9999,N_9822,N_9809);
nor U10000 (N_10000,N_9700,N_9795);
nor U10001 (N_10001,N_9788,N_9647);
and U10002 (N_10002,N_9664,N_9847);
nand U10003 (N_10003,N_9651,N_9873);
nor U10004 (N_10004,N_9804,N_9666);
or U10005 (N_10005,N_9712,N_9817);
xnor U10006 (N_10006,N_9882,N_9686);
nor U10007 (N_10007,N_9603,N_9886);
nand U10008 (N_10008,N_9625,N_9663);
nor U10009 (N_10009,N_9840,N_9638);
nor U10010 (N_10010,N_9633,N_9790);
nor U10011 (N_10011,N_9623,N_9618);
nand U10012 (N_10012,N_9764,N_9870);
or U10013 (N_10013,N_9607,N_9661);
and U10014 (N_10014,N_9682,N_9824);
xnor U10015 (N_10015,N_9815,N_9851);
and U10016 (N_10016,N_9621,N_9785);
nor U10017 (N_10017,N_9821,N_9653);
nand U10018 (N_10018,N_9732,N_9735);
or U10019 (N_10019,N_9628,N_9820);
nand U10020 (N_10020,N_9750,N_9747);
nand U10021 (N_10021,N_9705,N_9896);
and U10022 (N_10022,N_9816,N_9670);
nand U10023 (N_10023,N_9891,N_9729);
nor U10024 (N_10024,N_9714,N_9887);
xor U10025 (N_10025,N_9667,N_9828);
or U10026 (N_10026,N_9679,N_9645);
or U10027 (N_10027,N_9861,N_9803);
xnor U10028 (N_10028,N_9629,N_9834);
nor U10029 (N_10029,N_9898,N_9897);
and U10030 (N_10030,N_9683,N_9693);
nor U10031 (N_10031,N_9775,N_9792);
nand U10032 (N_10032,N_9715,N_9836);
xor U10033 (N_10033,N_9797,N_9721);
or U10034 (N_10034,N_9881,N_9813);
xnor U10035 (N_10035,N_9665,N_9697);
or U10036 (N_10036,N_9606,N_9754);
xnor U10037 (N_10037,N_9707,N_9640);
xor U10038 (N_10038,N_9810,N_9839);
or U10039 (N_10039,N_9724,N_9672);
and U10040 (N_10040,N_9843,N_9644);
and U10041 (N_10041,N_9879,N_9883);
or U10042 (N_10042,N_9659,N_9857);
xnor U10043 (N_10043,N_9726,N_9739);
or U10044 (N_10044,N_9696,N_9889);
and U10045 (N_10045,N_9604,N_9736);
and U10046 (N_10046,N_9719,N_9717);
and U10047 (N_10047,N_9692,N_9671);
and U10048 (N_10048,N_9880,N_9858);
nand U10049 (N_10049,N_9708,N_9704);
or U10050 (N_10050,N_9703,N_9637);
and U10051 (N_10051,N_9716,N_9886);
nand U10052 (N_10052,N_9812,N_9776);
nand U10053 (N_10053,N_9603,N_9817);
nand U10054 (N_10054,N_9687,N_9696);
and U10055 (N_10055,N_9685,N_9640);
and U10056 (N_10056,N_9633,N_9878);
nand U10057 (N_10057,N_9844,N_9767);
and U10058 (N_10058,N_9769,N_9844);
or U10059 (N_10059,N_9748,N_9813);
and U10060 (N_10060,N_9780,N_9690);
and U10061 (N_10061,N_9858,N_9770);
nor U10062 (N_10062,N_9879,N_9760);
nand U10063 (N_10063,N_9784,N_9800);
nand U10064 (N_10064,N_9793,N_9647);
xnor U10065 (N_10065,N_9880,N_9666);
or U10066 (N_10066,N_9848,N_9674);
or U10067 (N_10067,N_9850,N_9872);
and U10068 (N_10068,N_9644,N_9896);
nand U10069 (N_10069,N_9888,N_9803);
nand U10070 (N_10070,N_9696,N_9748);
nor U10071 (N_10071,N_9748,N_9752);
nand U10072 (N_10072,N_9729,N_9601);
or U10073 (N_10073,N_9869,N_9642);
nor U10074 (N_10074,N_9778,N_9838);
or U10075 (N_10075,N_9759,N_9772);
xor U10076 (N_10076,N_9783,N_9690);
or U10077 (N_10077,N_9623,N_9681);
nor U10078 (N_10078,N_9894,N_9867);
xor U10079 (N_10079,N_9888,N_9699);
nand U10080 (N_10080,N_9797,N_9717);
nor U10081 (N_10081,N_9601,N_9834);
nand U10082 (N_10082,N_9810,N_9643);
xnor U10083 (N_10083,N_9620,N_9762);
or U10084 (N_10084,N_9791,N_9878);
and U10085 (N_10085,N_9655,N_9793);
nand U10086 (N_10086,N_9735,N_9757);
nor U10087 (N_10087,N_9858,N_9888);
or U10088 (N_10088,N_9706,N_9778);
or U10089 (N_10089,N_9675,N_9649);
nand U10090 (N_10090,N_9841,N_9787);
xor U10091 (N_10091,N_9863,N_9767);
and U10092 (N_10092,N_9752,N_9838);
and U10093 (N_10093,N_9858,N_9819);
xor U10094 (N_10094,N_9785,N_9859);
nand U10095 (N_10095,N_9824,N_9774);
or U10096 (N_10096,N_9643,N_9889);
or U10097 (N_10097,N_9816,N_9728);
and U10098 (N_10098,N_9776,N_9766);
or U10099 (N_10099,N_9641,N_9720);
nand U10100 (N_10100,N_9868,N_9707);
nor U10101 (N_10101,N_9849,N_9709);
nor U10102 (N_10102,N_9712,N_9679);
nor U10103 (N_10103,N_9803,N_9766);
xor U10104 (N_10104,N_9820,N_9698);
nor U10105 (N_10105,N_9894,N_9790);
nor U10106 (N_10106,N_9675,N_9876);
or U10107 (N_10107,N_9607,N_9732);
nand U10108 (N_10108,N_9720,N_9863);
xor U10109 (N_10109,N_9742,N_9651);
nand U10110 (N_10110,N_9849,N_9860);
or U10111 (N_10111,N_9609,N_9672);
nor U10112 (N_10112,N_9627,N_9649);
nand U10113 (N_10113,N_9793,N_9763);
nor U10114 (N_10114,N_9712,N_9684);
nor U10115 (N_10115,N_9872,N_9835);
nor U10116 (N_10116,N_9780,N_9754);
and U10117 (N_10117,N_9840,N_9660);
xor U10118 (N_10118,N_9742,N_9737);
nor U10119 (N_10119,N_9743,N_9847);
nor U10120 (N_10120,N_9894,N_9672);
nor U10121 (N_10121,N_9670,N_9734);
xor U10122 (N_10122,N_9734,N_9857);
nand U10123 (N_10123,N_9718,N_9660);
or U10124 (N_10124,N_9704,N_9742);
nor U10125 (N_10125,N_9750,N_9611);
nor U10126 (N_10126,N_9846,N_9764);
or U10127 (N_10127,N_9732,N_9862);
or U10128 (N_10128,N_9630,N_9708);
and U10129 (N_10129,N_9873,N_9864);
nor U10130 (N_10130,N_9865,N_9821);
nand U10131 (N_10131,N_9789,N_9620);
or U10132 (N_10132,N_9867,N_9850);
nand U10133 (N_10133,N_9833,N_9625);
or U10134 (N_10134,N_9664,N_9827);
or U10135 (N_10135,N_9719,N_9616);
xor U10136 (N_10136,N_9643,N_9715);
xnor U10137 (N_10137,N_9714,N_9615);
nor U10138 (N_10138,N_9715,N_9873);
or U10139 (N_10139,N_9838,N_9755);
xnor U10140 (N_10140,N_9643,N_9672);
xnor U10141 (N_10141,N_9748,N_9794);
xnor U10142 (N_10142,N_9778,N_9801);
or U10143 (N_10143,N_9690,N_9654);
nand U10144 (N_10144,N_9737,N_9702);
and U10145 (N_10145,N_9876,N_9783);
nor U10146 (N_10146,N_9883,N_9626);
or U10147 (N_10147,N_9804,N_9884);
nand U10148 (N_10148,N_9873,N_9899);
nand U10149 (N_10149,N_9710,N_9692);
nor U10150 (N_10150,N_9885,N_9757);
and U10151 (N_10151,N_9754,N_9719);
nand U10152 (N_10152,N_9789,N_9859);
nor U10153 (N_10153,N_9678,N_9844);
or U10154 (N_10154,N_9716,N_9613);
and U10155 (N_10155,N_9794,N_9650);
nand U10156 (N_10156,N_9781,N_9824);
xnor U10157 (N_10157,N_9667,N_9888);
nor U10158 (N_10158,N_9815,N_9789);
nor U10159 (N_10159,N_9859,N_9880);
or U10160 (N_10160,N_9870,N_9620);
or U10161 (N_10161,N_9767,N_9609);
nand U10162 (N_10162,N_9768,N_9781);
nor U10163 (N_10163,N_9836,N_9675);
xor U10164 (N_10164,N_9835,N_9799);
and U10165 (N_10165,N_9692,N_9737);
nand U10166 (N_10166,N_9768,N_9647);
or U10167 (N_10167,N_9622,N_9688);
and U10168 (N_10168,N_9802,N_9788);
or U10169 (N_10169,N_9772,N_9627);
and U10170 (N_10170,N_9663,N_9814);
nand U10171 (N_10171,N_9709,N_9691);
xor U10172 (N_10172,N_9680,N_9804);
nor U10173 (N_10173,N_9770,N_9890);
or U10174 (N_10174,N_9884,N_9814);
nand U10175 (N_10175,N_9753,N_9687);
xnor U10176 (N_10176,N_9712,N_9625);
and U10177 (N_10177,N_9896,N_9669);
nand U10178 (N_10178,N_9750,N_9881);
or U10179 (N_10179,N_9747,N_9878);
nor U10180 (N_10180,N_9798,N_9613);
nand U10181 (N_10181,N_9828,N_9807);
xnor U10182 (N_10182,N_9783,N_9822);
and U10183 (N_10183,N_9655,N_9896);
or U10184 (N_10184,N_9686,N_9886);
or U10185 (N_10185,N_9750,N_9851);
nand U10186 (N_10186,N_9606,N_9616);
xnor U10187 (N_10187,N_9827,N_9899);
xor U10188 (N_10188,N_9619,N_9869);
xnor U10189 (N_10189,N_9796,N_9692);
and U10190 (N_10190,N_9785,N_9716);
nand U10191 (N_10191,N_9841,N_9884);
nand U10192 (N_10192,N_9888,N_9634);
xnor U10193 (N_10193,N_9867,N_9864);
and U10194 (N_10194,N_9881,N_9820);
and U10195 (N_10195,N_9673,N_9613);
nor U10196 (N_10196,N_9890,N_9849);
or U10197 (N_10197,N_9665,N_9810);
or U10198 (N_10198,N_9676,N_9615);
or U10199 (N_10199,N_9701,N_9779);
and U10200 (N_10200,N_9955,N_10041);
nor U10201 (N_10201,N_10018,N_9918);
nand U10202 (N_10202,N_9946,N_9959);
nor U10203 (N_10203,N_9969,N_9984);
xnor U10204 (N_10204,N_10145,N_10023);
or U10205 (N_10205,N_9906,N_10102);
nor U10206 (N_10206,N_9975,N_10127);
xor U10207 (N_10207,N_10110,N_10176);
and U10208 (N_10208,N_9968,N_10155);
xnor U10209 (N_10209,N_10188,N_9915);
or U10210 (N_10210,N_10111,N_9910);
or U10211 (N_10211,N_10129,N_9940);
nor U10212 (N_10212,N_9972,N_10099);
xnor U10213 (N_10213,N_9988,N_10170);
or U10214 (N_10214,N_10094,N_10156);
or U10215 (N_10215,N_10043,N_10124);
or U10216 (N_10216,N_10029,N_9919);
nand U10217 (N_10217,N_10052,N_10025);
and U10218 (N_10218,N_10087,N_10195);
and U10219 (N_10219,N_10016,N_9938);
nor U10220 (N_10220,N_10134,N_10001);
nor U10221 (N_10221,N_10101,N_9914);
nand U10222 (N_10222,N_9996,N_10165);
nand U10223 (N_10223,N_9930,N_10148);
nor U10224 (N_10224,N_10081,N_9971);
nand U10225 (N_10225,N_9932,N_10046);
xnor U10226 (N_10226,N_9987,N_10003);
or U10227 (N_10227,N_10075,N_10189);
nor U10228 (N_10228,N_10019,N_9980);
xor U10229 (N_10229,N_9937,N_10096);
xor U10230 (N_10230,N_10097,N_9907);
xor U10231 (N_10231,N_9999,N_10157);
xor U10232 (N_10232,N_10083,N_10106);
nor U10233 (N_10233,N_9982,N_9953);
xor U10234 (N_10234,N_9952,N_10153);
or U10235 (N_10235,N_10090,N_10143);
nor U10236 (N_10236,N_10053,N_9989);
nand U10237 (N_10237,N_10071,N_10063);
and U10238 (N_10238,N_10120,N_10002);
and U10239 (N_10239,N_10047,N_9998);
xnor U10240 (N_10240,N_10114,N_9961);
xor U10241 (N_10241,N_10118,N_10100);
and U10242 (N_10242,N_10072,N_10054);
xnor U10243 (N_10243,N_9990,N_10040);
xor U10244 (N_10244,N_10051,N_10123);
nor U10245 (N_10245,N_10020,N_10125);
and U10246 (N_10246,N_10098,N_9993);
xnor U10247 (N_10247,N_10042,N_10180);
or U10248 (N_10248,N_9921,N_10192);
xnor U10249 (N_10249,N_10166,N_10130);
nand U10250 (N_10250,N_9957,N_9905);
or U10251 (N_10251,N_10161,N_10035);
or U10252 (N_10252,N_10034,N_10048);
nor U10253 (N_10253,N_10158,N_9978);
nor U10254 (N_10254,N_10162,N_9974);
nor U10255 (N_10255,N_10128,N_10109);
nor U10256 (N_10256,N_9979,N_10138);
or U10257 (N_10257,N_10191,N_10171);
and U10258 (N_10258,N_10131,N_9950);
nor U10259 (N_10259,N_9970,N_10050);
or U10260 (N_10260,N_10070,N_10066);
xor U10261 (N_10261,N_9908,N_10177);
or U10262 (N_10262,N_9903,N_9928);
and U10263 (N_10263,N_9941,N_10108);
nand U10264 (N_10264,N_10168,N_10039);
nor U10265 (N_10265,N_10086,N_10167);
nor U10266 (N_10266,N_9934,N_10062);
xnor U10267 (N_10267,N_9922,N_9951);
nor U10268 (N_10268,N_10154,N_9913);
or U10269 (N_10269,N_10007,N_10080);
nor U10270 (N_10270,N_10144,N_9949);
nand U10271 (N_10271,N_10017,N_10008);
nand U10272 (N_10272,N_10164,N_10027);
nand U10273 (N_10273,N_9991,N_10181);
or U10274 (N_10274,N_9945,N_9962);
nor U10275 (N_10275,N_10067,N_10059);
and U10276 (N_10276,N_10178,N_10163);
nor U10277 (N_10277,N_10079,N_9977);
xor U10278 (N_10278,N_10150,N_10006);
or U10279 (N_10279,N_10000,N_9995);
and U10280 (N_10280,N_9933,N_10116);
and U10281 (N_10281,N_10172,N_9965);
or U10282 (N_10282,N_10031,N_10038);
and U10283 (N_10283,N_10026,N_10073);
xor U10284 (N_10284,N_10015,N_10119);
xor U10285 (N_10285,N_10175,N_9997);
or U10286 (N_10286,N_10121,N_10126);
xnor U10287 (N_10287,N_10169,N_10179);
and U10288 (N_10288,N_9911,N_10021);
nor U10289 (N_10289,N_9931,N_10193);
xor U10290 (N_10290,N_9939,N_9904);
xor U10291 (N_10291,N_10077,N_10057);
xor U10292 (N_10292,N_10122,N_9900);
nand U10293 (N_10293,N_9917,N_10136);
nand U10294 (N_10294,N_9901,N_9964);
nand U10295 (N_10295,N_10095,N_9994);
nor U10296 (N_10296,N_10084,N_10159);
or U10297 (N_10297,N_9935,N_10183);
and U10298 (N_10298,N_9916,N_10012);
and U10299 (N_10299,N_10078,N_10089);
or U10300 (N_10300,N_9954,N_10187);
xnor U10301 (N_10301,N_10194,N_9967);
nor U10302 (N_10302,N_9960,N_10068);
xor U10303 (N_10303,N_10152,N_9942);
and U10304 (N_10304,N_10049,N_10088);
nand U10305 (N_10305,N_10104,N_10190);
nand U10306 (N_10306,N_9912,N_9920);
nand U10307 (N_10307,N_10082,N_10032);
nand U10308 (N_10308,N_10140,N_9926);
and U10309 (N_10309,N_9927,N_10037);
and U10310 (N_10310,N_10009,N_10093);
or U10311 (N_10311,N_10044,N_10036);
nand U10312 (N_10312,N_10107,N_9976);
or U10313 (N_10313,N_10182,N_10173);
nand U10314 (N_10314,N_10139,N_10135);
nand U10315 (N_10315,N_9963,N_10147);
and U10316 (N_10316,N_10004,N_10091);
nor U10317 (N_10317,N_10058,N_10103);
nor U10318 (N_10318,N_10185,N_10069);
and U10319 (N_10319,N_9944,N_9948);
or U10320 (N_10320,N_10151,N_10092);
and U10321 (N_10321,N_9985,N_10011);
and U10322 (N_10322,N_9992,N_9958);
nand U10323 (N_10323,N_10186,N_9943);
nor U10324 (N_10324,N_10014,N_10022);
xnor U10325 (N_10325,N_10056,N_10184);
nor U10326 (N_10326,N_9983,N_10141);
nor U10327 (N_10327,N_10065,N_9902);
nor U10328 (N_10328,N_10085,N_10113);
nor U10329 (N_10329,N_10028,N_9909);
or U10330 (N_10330,N_9923,N_10076);
nor U10331 (N_10331,N_10174,N_10117);
and U10332 (N_10332,N_9924,N_10060);
nand U10333 (N_10333,N_9966,N_10055);
or U10334 (N_10334,N_10074,N_9981);
nand U10335 (N_10335,N_10137,N_10045);
nand U10336 (N_10336,N_10112,N_10030);
xnor U10337 (N_10337,N_10160,N_10199);
and U10338 (N_10338,N_10061,N_10149);
nand U10339 (N_10339,N_10196,N_10198);
nand U10340 (N_10340,N_10105,N_9956);
nand U10341 (N_10341,N_10010,N_10115);
or U10342 (N_10342,N_10132,N_10197);
nand U10343 (N_10343,N_9936,N_9947);
nand U10344 (N_10344,N_10064,N_9929);
xor U10345 (N_10345,N_10133,N_10146);
and U10346 (N_10346,N_10013,N_10005);
xor U10347 (N_10347,N_9986,N_10142);
or U10348 (N_10348,N_9925,N_10024);
or U10349 (N_10349,N_10033,N_9973);
nand U10350 (N_10350,N_10159,N_10054);
nand U10351 (N_10351,N_10152,N_9928);
and U10352 (N_10352,N_10175,N_10109);
or U10353 (N_10353,N_10067,N_10179);
nor U10354 (N_10354,N_10038,N_10153);
nor U10355 (N_10355,N_10010,N_10158);
or U10356 (N_10356,N_9951,N_10072);
xor U10357 (N_10357,N_9984,N_9975);
nor U10358 (N_10358,N_10038,N_10155);
or U10359 (N_10359,N_10040,N_10038);
nor U10360 (N_10360,N_10064,N_9956);
and U10361 (N_10361,N_10010,N_9997);
nor U10362 (N_10362,N_10002,N_9978);
xnor U10363 (N_10363,N_10110,N_9934);
nand U10364 (N_10364,N_10146,N_9933);
nand U10365 (N_10365,N_10085,N_10077);
or U10366 (N_10366,N_9991,N_9945);
or U10367 (N_10367,N_9945,N_10017);
xnor U10368 (N_10368,N_10176,N_10106);
and U10369 (N_10369,N_9938,N_10103);
xor U10370 (N_10370,N_9905,N_10151);
xor U10371 (N_10371,N_10146,N_9996);
nand U10372 (N_10372,N_9927,N_10103);
or U10373 (N_10373,N_10074,N_10026);
or U10374 (N_10374,N_10108,N_10051);
and U10375 (N_10375,N_9905,N_9931);
or U10376 (N_10376,N_10033,N_10148);
nand U10377 (N_10377,N_10146,N_10188);
xnor U10378 (N_10378,N_10071,N_9941);
or U10379 (N_10379,N_9957,N_10171);
nand U10380 (N_10380,N_10012,N_9908);
or U10381 (N_10381,N_10134,N_9917);
nor U10382 (N_10382,N_9985,N_10133);
nor U10383 (N_10383,N_10130,N_10093);
or U10384 (N_10384,N_10130,N_9929);
or U10385 (N_10385,N_9973,N_10169);
or U10386 (N_10386,N_10001,N_10095);
or U10387 (N_10387,N_10046,N_10090);
nand U10388 (N_10388,N_9932,N_10132);
nand U10389 (N_10389,N_9975,N_10159);
or U10390 (N_10390,N_10178,N_10031);
nor U10391 (N_10391,N_10079,N_10051);
nand U10392 (N_10392,N_9963,N_10125);
nand U10393 (N_10393,N_10158,N_10001);
xor U10394 (N_10394,N_9976,N_10141);
nand U10395 (N_10395,N_10063,N_10097);
nor U10396 (N_10396,N_10003,N_10130);
nand U10397 (N_10397,N_9931,N_9932);
nand U10398 (N_10398,N_10055,N_10072);
and U10399 (N_10399,N_10078,N_10080);
nor U10400 (N_10400,N_10181,N_9904);
or U10401 (N_10401,N_10167,N_10125);
xor U10402 (N_10402,N_9990,N_9949);
and U10403 (N_10403,N_10036,N_9926);
xnor U10404 (N_10404,N_10098,N_10184);
and U10405 (N_10405,N_10006,N_10052);
and U10406 (N_10406,N_9999,N_10102);
or U10407 (N_10407,N_9908,N_10157);
or U10408 (N_10408,N_10019,N_10004);
xor U10409 (N_10409,N_9925,N_9903);
and U10410 (N_10410,N_10159,N_9922);
and U10411 (N_10411,N_10015,N_10111);
nor U10412 (N_10412,N_10073,N_10118);
xnor U10413 (N_10413,N_10184,N_9939);
nor U10414 (N_10414,N_9955,N_10150);
nor U10415 (N_10415,N_9986,N_10170);
or U10416 (N_10416,N_9911,N_9973);
nor U10417 (N_10417,N_9906,N_10031);
nor U10418 (N_10418,N_9930,N_9954);
and U10419 (N_10419,N_10024,N_10085);
nand U10420 (N_10420,N_10055,N_9978);
and U10421 (N_10421,N_10036,N_9954);
and U10422 (N_10422,N_10104,N_10068);
nor U10423 (N_10423,N_10004,N_10024);
and U10424 (N_10424,N_9999,N_9915);
nor U10425 (N_10425,N_10139,N_9902);
nand U10426 (N_10426,N_9946,N_10133);
or U10427 (N_10427,N_10197,N_10187);
and U10428 (N_10428,N_9909,N_10048);
nor U10429 (N_10429,N_10019,N_10142);
and U10430 (N_10430,N_10058,N_10070);
or U10431 (N_10431,N_10060,N_10129);
xnor U10432 (N_10432,N_10148,N_10174);
nor U10433 (N_10433,N_10105,N_9950);
xor U10434 (N_10434,N_10121,N_9951);
nor U10435 (N_10435,N_10028,N_10071);
nor U10436 (N_10436,N_9963,N_9916);
nor U10437 (N_10437,N_9990,N_10066);
xor U10438 (N_10438,N_9903,N_10193);
or U10439 (N_10439,N_10181,N_10003);
nor U10440 (N_10440,N_10074,N_9923);
and U10441 (N_10441,N_10028,N_9945);
or U10442 (N_10442,N_9972,N_10011);
xor U10443 (N_10443,N_10171,N_10176);
xnor U10444 (N_10444,N_10153,N_10184);
xnor U10445 (N_10445,N_10118,N_10008);
and U10446 (N_10446,N_9997,N_9945);
nor U10447 (N_10447,N_10084,N_10101);
xor U10448 (N_10448,N_9905,N_10043);
nand U10449 (N_10449,N_10115,N_10179);
nor U10450 (N_10450,N_9925,N_9921);
nor U10451 (N_10451,N_10099,N_10015);
xnor U10452 (N_10452,N_10003,N_10099);
nor U10453 (N_10453,N_10132,N_10122);
nor U10454 (N_10454,N_9949,N_9935);
or U10455 (N_10455,N_9920,N_9969);
and U10456 (N_10456,N_9970,N_9928);
and U10457 (N_10457,N_10112,N_10174);
or U10458 (N_10458,N_10147,N_10056);
or U10459 (N_10459,N_9980,N_10053);
or U10460 (N_10460,N_10019,N_9912);
xor U10461 (N_10461,N_10188,N_10039);
nand U10462 (N_10462,N_9923,N_10161);
or U10463 (N_10463,N_10181,N_9956);
or U10464 (N_10464,N_10038,N_10008);
xor U10465 (N_10465,N_10190,N_10162);
nand U10466 (N_10466,N_9971,N_9960);
or U10467 (N_10467,N_10174,N_9988);
nand U10468 (N_10468,N_10072,N_10050);
and U10469 (N_10469,N_9965,N_10154);
and U10470 (N_10470,N_10124,N_9998);
or U10471 (N_10471,N_10007,N_9933);
or U10472 (N_10472,N_10093,N_9960);
and U10473 (N_10473,N_9955,N_10026);
and U10474 (N_10474,N_10152,N_10177);
and U10475 (N_10475,N_9957,N_9996);
xor U10476 (N_10476,N_10126,N_10008);
or U10477 (N_10477,N_9907,N_10091);
or U10478 (N_10478,N_9930,N_10078);
nand U10479 (N_10479,N_9929,N_9983);
xnor U10480 (N_10480,N_10118,N_10064);
nor U10481 (N_10481,N_10156,N_10160);
xnor U10482 (N_10482,N_10110,N_10084);
nor U10483 (N_10483,N_10199,N_10174);
xnor U10484 (N_10484,N_10137,N_9917);
and U10485 (N_10485,N_9994,N_10173);
nand U10486 (N_10486,N_10123,N_9994);
nor U10487 (N_10487,N_10024,N_10090);
xnor U10488 (N_10488,N_10163,N_10037);
and U10489 (N_10489,N_10159,N_9952);
or U10490 (N_10490,N_10046,N_9933);
nor U10491 (N_10491,N_10070,N_9932);
nor U10492 (N_10492,N_10171,N_10100);
nor U10493 (N_10493,N_9921,N_9916);
nor U10494 (N_10494,N_10108,N_10113);
or U10495 (N_10495,N_9935,N_10129);
and U10496 (N_10496,N_10139,N_10006);
and U10497 (N_10497,N_10018,N_10039);
or U10498 (N_10498,N_9917,N_9932);
and U10499 (N_10499,N_10190,N_10021);
nor U10500 (N_10500,N_10366,N_10325);
xor U10501 (N_10501,N_10293,N_10439);
nor U10502 (N_10502,N_10255,N_10280);
and U10503 (N_10503,N_10324,N_10215);
nand U10504 (N_10504,N_10236,N_10436);
and U10505 (N_10505,N_10284,N_10239);
xor U10506 (N_10506,N_10445,N_10268);
or U10507 (N_10507,N_10313,N_10406);
nor U10508 (N_10508,N_10435,N_10283);
and U10509 (N_10509,N_10465,N_10491);
xnor U10510 (N_10510,N_10235,N_10487);
xnor U10511 (N_10511,N_10404,N_10291);
and U10512 (N_10512,N_10372,N_10222);
or U10513 (N_10513,N_10490,N_10365);
nor U10514 (N_10514,N_10401,N_10202);
and U10515 (N_10515,N_10356,N_10444);
nor U10516 (N_10516,N_10303,N_10273);
nand U10517 (N_10517,N_10389,N_10361);
or U10518 (N_10518,N_10319,N_10346);
xnor U10519 (N_10519,N_10269,N_10305);
xor U10520 (N_10520,N_10419,N_10320);
nor U10521 (N_10521,N_10249,N_10351);
or U10522 (N_10522,N_10224,N_10450);
or U10523 (N_10523,N_10331,N_10229);
or U10524 (N_10524,N_10262,N_10385);
nor U10525 (N_10525,N_10295,N_10272);
nor U10526 (N_10526,N_10399,N_10230);
and U10527 (N_10527,N_10397,N_10413);
or U10528 (N_10528,N_10422,N_10207);
and U10529 (N_10529,N_10471,N_10321);
or U10530 (N_10530,N_10288,N_10352);
nand U10531 (N_10531,N_10474,N_10381);
and U10532 (N_10532,N_10271,N_10452);
nand U10533 (N_10533,N_10355,N_10276);
nand U10534 (N_10534,N_10393,N_10316);
nor U10535 (N_10535,N_10424,N_10226);
nand U10536 (N_10536,N_10300,N_10387);
and U10537 (N_10537,N_10277,N_10213);
or U10538 (N_10538,N_10473,N_10302);
and U10539 (N_10539,N_10468,N_10250);
nor U10540 (N_10540,N_10309,N_10344);
or U10541 (N_10541,N_10247,N_10314);
and U10542 (N_10542,N_10498,N_10263);
nand U10543 (N_10543,N_10231,N_10223);
and U10544 (N_10544,N_10257,N_10426);
xor U10545 (N_10545,N_10376,N_10217);
nand U10546 (N_10546,N_10308,N_10335);
nor U10547 (N_10547,N_10488,N_10287);
nor U10548 (N_10548,N_10336,N_10294);
nand U10549 (N_10549,N_10265,N_10279);
and U10550 (N_10550,N_10274,N_10216);
xnor U10551 (N_10551,N_10275,N_10353);
nor U10552 (N_10552,N_10359,N_10464);
nor U10553 (N_10553,N_10453,N_10375);
nor U10554 (N_10554,N_10296,N_10469);
and U10555 (N_10555,N_10396,N_10438);
and U10556 (N_10556,N_10330,N_10432);
nor U10557 (N_10557,N_10204,N_10493);
xor U10558 (N_10558,N_10433,N_10259);
and U10559 (N_10559,N_10443,N_10323);
nand U10560 (N_10560,N_10383,N_10253);
xnor U10561 (N_10561,N_10244,N_10270);
and U10562 (N_10562,N_10329,N_10341);
or U10563 (N_10563,N_10460,N_10251);
or U10564 (N_10564,N_10298,N_10260);
or U10565 (N_10565,N_10338,N_10348);
or U10566 (N_10566,N_10201,N_10340);
and U10567 (N_10567,N_10403,N_10417);
and U10568 (N_10568,N_10237,N_10499);
nor U10569 (N_10569,N_10437,N_10379);
and U10570 (N_10570,N_10392,N_10412);
and U10571 (N_10571,N_10382,N_10306);
and U10572 (N_10572,N_10241,N_10307);
nor U10573 (N_10573,N_10484,N_10343);
nor U10574 (N_10574,N_10354,N_10221);
or U10575 (N_10575,N_10481,N_10496);
nor U10576 (N_10576,N_10391,N_10282);
xnor U10577 (N_10577,N_10357,N_10225);
xnor U10578 (N_10578,N_10281,N_10394);
xnor U10579 (N_10579,N_10209,N_10371);
and U10580 (N_10580,N_10358,N_10342);
or U10581 (N_10581,N_10486,N_10203);
or U10582 (N_10582,N_10364,N_10467);
xnor U10583 (N_10583,N_10256,N_10278);
and U10584 (N_10584,N_10388,N_10440);
nor U10585 (N_10585,N_10373,N_10483);
nand U10586 (N_10586,N_10326,N_10350);
and U10587 (N_10587,N_10240,N_10299);
and U10588 (N_10588,N_10434,N_10214);
nor U10589 (N_10589,N_10349,N_10328);
xnor U10590 (N_10590,N_10233,N_10398);
nand U10591 (N_10591,N_10384,N_10420);
xor U10592 (N_10592,N_10347,N_10470);
and U10593 (N_10593,N_10285,N_10458);
xor U10594 (N_10594,N_10267,N_10414);
xnor U10595 (N_10595,N_10489,N_10334);
or U10596 (N_10596,N_10457,N_10451);
xnor U10597 (N_10597,N_10418,N_10243);
or U10598 (N_10598,N_10246,N_10345);
nor U10599 (N_10599,N_10461,N_10315);
nand U10600 (N_10600,N_10421,N_10415);
or U10601 (N_10601,N_10258,N_10339);
nand U10602 (N_10602,N_10475,N_10322);
nor U10603 (N_10603,N_10264,N_10368);
nor U10604 (N_10604,N_10261,N_10416);
or U10605 (N_10605,N_10390,N_10304);
nor U10606 (N_10606,N_10459,N_10477);
or U10607 (N_10607,N_10362,N_10200);
xor U10608 (N_10608,N_10482,N_10462);
or U10609 (N_10609,N_10378,N_10312);
xor U10610 (N_10610,N_10428,N_10289);
nor U10611 (N_10611,N_10286,N_10219);
nand U10612 (N_10612,N_10211,N_10408);
or U10613 (N_10613,N_10363,N_10380);
nor U10614 (N_10614,N_10292,N_10218);
nand U10615 (N_10615,N_10429,N_10370);
xnor U10616 (N_10616,N_10455,N_10497);
or U10617 (N_10617,N_10310,N_10234);
or U10618 (N_10618,N_10411,N_10409);
nor U10619 (N_10619,N_10400,N_10386);
or U10620 (N_10620,N_10248,N_10242);
and U10621 (N_10621,N_10447,N_10466);
nand U10622 (N_10622,N_10377,N_10205);
or U10623 (N_10623,N_10252,N_10301);
or U10624 (N_10624,N_10318,N_10448);
nand U10625 (N_10625,N_10430,N_10232);
nand U10626 (N_10626,N_10478,N_10427);
nor U10627 (N_10627,N_10446,N_10492);
xor U10628 (N_10628,N_10212,N_10206);
xnor U10629 (N_10629,N_10208,N_10311);
and U10630 (N_10630,N_10449,N_10266);
nor U10631 (N_10631,N_10442,N_10463);
xor U10632 (N_10632,N_10407,N_10494);
or U10633 (N_10633,N_10425,N_10431);
nor U10634 (N_10634,N_10297,N_10228);
nand U10635 (N_10635,N_10410,N_10290);
xor U10636 (N_10636,N_10327,N_10480);
or U10637 (N_10637,N_10472,N_10441);
and U10638 (N_10638,N_10227,N_10454);
nand U10639 (N_10639,N_10254,N_10360);
nor U10640 (N_10640,N_10374,N_10220);
or U10641 (N_10641,N_10238,N_10495);
and U10642 (N_10642,N_10317,N_10485);
nand U10643 (N_10643,N_10210,N_10479);
nor U10644 (N_10644,N_10456,N_10337);
xnor U10645 (N_10645,N_10245,N_10476);
nor U10646 (N_10646,N_10405,N_10367);
nor U10647 (N_10647,N_10423,N_10333);
nor U10648 (N_10648,N_10402,N_10369);
xnor U10649 (N_10649,N_10395,N_10332);
nor U10650 (N_10650,N_10332,N_10250);
or U10651 (N_10651,N_10492,N_10437);
nor U10652 (N_10652,N_10486,N_10340);
or U10653 (N_10653,N_10203,N_10263);
and U10654 (N_10654,N_10236,N_10306);
nand U10655 (N_10655,N_10267,N_10429);
or U10656 (N_10656,N_10394,N_10392);
xor U10657 (N_10657,N_10283,N_10212);
and U10658 (N_10658,N_10354,N_10236);
nand U10659 (N_10659,N_10438,N_10486);
nand U10660 (N_10660,N_10221,N_10388);
nor U10661 (N_10661,N_10493,N_10414);
nor U10662 (N_10662,N_10272,N_10328);
or U10663 (N_10663,N_10214,N_10291);
nor U10664 (N_10664,N_10306,N_10273);
nor U10665 (N_10665,N_10272,N_10317);
and U10666 (N_10666,N_10437,N_10461);
nand U10667 (N_10667,N_10370,N_10357);
xor U10668 (N_10668,N_10441,N_10353);
or U10669 (N_10669,N_10430,N_10237);
nor U10670 (N_10670,N_10302,N_10439);
or U10671 (N_10671,N_10418,N_10415);
and U10672 (N_10672,N_10491,N_10475);
and U10673 (N_10673,N_10228,N_10390);
xor U10674 (N_10674,N_10362,N_10213);
nand U10675 (N_10675,N_10219,N_10440);
or U10676 (N_10676,N_10489,N_10448);
nand U10677 (N_10677,N_10426,N_10259);
nand U10678 (N_10678,N_10459,N_10251);
xnor U10679 (N_10679,N_10408,N_10260);
or U10680 (N_10680,N_10280,N_10396);
nor U10681 (N_10681,N_10265,N_10427);
nand U10682 (N_10682,N_10314,N_10223);
or U10683 (N_10683,N_10269,N_10452);
xor U10684 (N_10684,N_10265,N_10482);
nor U10685 (N_10685,N_10229,N_10392);
or U10686 (N_10686,N_10349,N_10407);
or U10687 (N_10687,N_10219,N_10224);
nor U10688 (N_10688,N_10240,N_10447);
or U10689 (N_10689,N_10474,N_10444);
nand U10690 (N_10690,N_10413,N_10355);
xor U10691 (N_10691,N_10294,N_10390);
xor U10692 (N_10692,N_10437,N_10456);
nand U10693 (N_10693,N_10386,N_10268);
nand U10694 (N_10694,N_10369,N_10378);
nand U10695 (N_10695,N_10386,N_10215);
xnor U10696 (N_10696,N_10413,N_10352);
nand U10697 (N_10697,N_10273,N_10323);
nand U10698 (N_10698,N_10455,N_10424);
or U10699 (N_10699,N_10432,N_10243);
nand U10700 (N_10700,N_10353,N_10352);
or U10701 (N_10701,N_10290,N_10270);
nand U10702 (N_10702,N_10462,N_10269);
or U10703 (N_10703,N_10375,N_10300);
and U10704 (N_10704,N_10450,N_10401);
nand U10705 (N_10705,N_10377,N_10341);
or U10706 (N_10706,N_10322,N_10262);
and U10707 (N_10707,N_10320,N_10277);
nor U10708 (N_10708,N_10355,N_10473);
nor U10709 (N_10709,N_10422,N_10455);
xnor U10710 (N_10710,N_10410,N_10462);
or U10711 (N_10711,N_10245,N_10422);
xnor U10712 (N_10712,N_10265,N_10308);
xor U10713 (N_10713,N_10327,N_10209);
xor U10714 (N_10714,N_10215,N_10333);
xnor U10715 (N_10715,N_10492,N_10422);
or U10716 (N_10716,N_10287,N_10452);
and U10717 (N_10717,N_10241,N_10377);
nand U10718 (N_10718,N_10455,N_10209);
or U10719 (N_10719,N_10324,N_10201);
nor U10720 (N_10720,N_10247,N_10406);
and U10721 (N_10721,N_10435,N_10221);
nand U10722 (N_10722,N_10357,N_10243);
or U10723 (N_10723,N_10347,N_10219);
or U10724 (N_10724,N_10409,N_10254);
nand U10725 (N_10725,N_10359,N_10474);
nand U10726 (N_10726,N_10369,N_10313);
nand U10727 (N_10727,N_10409,N_10230);
xnor U10728 (N_10728,N_10476,N_10475);
nor U10729 (N_10729,N_10425,N_10405);
nand U10730 (N_10730,N_10324,N_10413);
nand U10731 (N_10731,N_10441,N_10358);
or U10732 (N_10732,N_10427,N_10210);
and U10733 (N_10733,N_10459,N_10264);
xnor U10734 (N_10734,N_10429,N_10230);
and U10735 (N_10735,N_10379,N_10206);
xor U10736 (N_10736,N_10419,N_10213);
nor U10737 (N_10737,N_10426,N_10271);
xor U10738 (N_10738,N_10388,N_10267);
nand U10739 (N_10739,N_10263,N_10335);
and U10740 (N_10740,N_10206,N_10492);
nand U10741 (N_10741,N_10290,N_10327);
or U10742 (N_10742,N_10338,N_10290);
nand U10743 (N_10743,N_10472,N_10409);
nand U10744 (N_10744,N_10491,N_10383);
and U10745 (N_10745,N_10488,N_10284);
xor U10746 (N_10746,N_10414,N_10341);
or U10747 (N_10747,N_10389,N_10473);
or U10748 (N_10748,N_10320,N_10404);
and U10749 (N_10749,N_10314,N_10308);
nand U10750 (N_10750,N_10393,N_10349);
xnor U10751 (N_10751,N_10386,N_10249);
nor U10752 (N_10752,N_10263,N_10212);
nor U10753 (N_10753,N_10374,N_10266);
or U10754 (N_10754,N_10293,N_10277);
xnor U10755 (N_10755,N_10492,N_10298);
nor U10756 (N_10756,N_10420,N_10490);
xnor U10757 (N_10757,N_10296,N_10271);
and U10758 (N_10758,N_10423,N_10247);
and U10759 (N_10759,N_10394,N_10457);
xnor U10760 (N_10760,N_10286,N_10227);
nor U10761 (N_10761,N_10422,N_10234);
nor U10762 (N_10762,N_10347,N_10479);
xor U10763 (N_10763,N_10210,N_10482);
or U10764 (N_10764,N_10419,N_10219);
or U10765 (N_10765,N_10262,N_10241);
and U10766 (N_10766,N_10307,N_10319);
nand U10767 (N_10767,N_10407,N_10489);
or U10768 (N_10768,N_10457,N_10264);
or U10769 (N_10769,N_10364,N_10395);
or U10770 (N_10770,N_10318,N_10389);
and U10771 (N_10771,N_10239,N_10419);
and U10772 (N_10772,N_10225,N_10213);
nor U10773 (N_10773,N_10399,N_10261);
and U10774 (N_10774,N_10241,N_10267);
nand U10775 (N_10775,N_10386,N_10402);
nor U10776 (N_10776,N_10425,N_10368);
or U10777 (N_10777,N_10269,N_10273);
nor U10778 (N_10778,N_10374,N_10413);
xnor U10779 (N_10779,N_10463,N_10384);
nand U10780 (N_10780,N_10276,N_10333);
nand U10781 (N_10781,N_10206,N_10387);
xnor U10782 (N_10782,N_10306,N_10419);
nand U10783 (N_10783,N_10214,N_10323);
xnor U10784 (N_10784,N_10288,N_10279);
nor U10785 (N_10785,N_10216,N_10326);
nor U10786 (N_10786,N_10418,N_10222);
xnor U10787 (N_10787,N_10487,N_10413);
and U10788 (N_10788,N_10446,N_10447);
nor U10789 (N_10789,N_10331,N_10232);
or U10790 (N_10790,N_10376,N_10363);
nand U10791 (N_10791,N_10343,N_10446);
or U10792 (N_10792,N_10334,N_10254);
and U10793 (N_10793,N_10446,N_10211);
xnor U10794 (N_10794,N_10229,N_10376);
nor U10795 (N_10795,N_10298,N_10249);
and U10796 (N_10796,N_10258,N_10439);
nand U10797 (N_10797,N_10251,N_10392);
and U10798 (N_10798,N_10368,N_10232);
and U10799 (N_10799,N_10497,N_10415);
nand U10800 (N_10800,N_10568,N_10573);
nor U10801 (N_10801,N_10588,N_10669);
nor U10802 (N_10802,N_10641,N_10512);
nand U10803 (N_10803,N_10535,N_10635);
nand U10804 (N_10804,N_10707,N_10737);
or U10805 (N_10805,N_10628,N_10760);
or U10806 (N_10806,N_10636,N_10735);
nand U10807 (N_10807,N_10786,N_10689);
nor U10808 (N_10808,N_10711,N_10534);
nor U10809 (N_10809,N_10649,N_10703);
nor U10810 (N_10810,N_10759,N_10688);
and U10811 (N_10811,N_10666,N_10548);
nor U10812 (N_10812,N_10640,N_10506);
and U10813 (N_10813,N_10772,N_10712);
nand U10814 (N_10814,N_10673,N_10753);
and U10815 (N_10815,N_10721,N_10773);
nor U10816 (N_10816,N_10608,N_10555);
and U10817 (N_10817,N_10579,N_10587);
xor U10818 (N_10818,N_10768,N_10706);
or U10819 (N_10819,N_10668,N_10532);
and U10820 (N_10820,N_10651,N_10634);
and U10821 (N_10821,N_10739,N_10769);
and U10822 (N_10822,N_10544,N_10530);
or U10823 (N_10823,N_10740,N_10536);
nand U10824 (N_10824,N_10732,N_10552);
xnor U10825 (N_10825,N_10779,N_10572);
and U10826 (N_10826,N_10744,N_10676);
nand U10827 (N_10827,N_10545,N_10715);
xor U10828 (N_10828,N_10664,N_10694);
nand U10829 (N_10829,N_10750,N_10583);
nand U10830 (N_10830,N_10595,N_10723);
nand U10831 (N_10831,N_10550,N_10604);
xnor U10832 (N_10832,N_10585,N_10594);
nand U10833 (N_10833,N_10660,N_10639);
nand U10834 (N_10834,N_10708,N_10751);
nand U10835 (N_10835,N_10613,N_10597);
nor U10836 (N_10836,N_10790,N_10500);
nand U10837 (N_10837,N_10637,N_10659);
xor U10838 (N_10838,N_10575,N_10531);
or U10839 (N_10839,N_10704,N_10513);
nor U10840 (N_10840,N_10690,N_10701);
xnor U10841 (N_10841,N_10736,N_10782);
xnor U10842 (N_10842,N_10565,N_10799);
nor U10843 (N_10843,N_10798,N_10691);
and U10844 (N_10844,N_10619,N_10655);
or U10845 (N_10845,N_10741,N_10516);
nor U10846 (N_10846,N_10503,N_10792);
xor U10847 (N_10847,N_10593,N_10724);
xor U10848 (N_10848,N_10557,N_10770);
and U10849 (N_10849,N_10700,N_10617);
nand U10850 (N_10850,N_10648,N_10783);
nor U10851 (N_10851,N_10778,N_10598);
nand U10852 (N_10852,N_10729,N_10791);
and U10853 (N_10853,N_10519,N_10510);
nor U10854 (N_10854,N_10713,N_10757);
and U10855 (N_10855,N_10775,N_10638);
or U10856 (N_10856,N_10733,N_10776);
nor U10857 (N_10857,N_10787,N_10797);
nor U10858 (N_10858,N_10501,N_10549);
nor U10859 (N_10859,N_10680,N_10656);
or U10860 (N_10860,N_10607,N_10710);
nor U10861 (N_10861,N_10631,N_10674);
nor U10862 (N_10862,N_10521,N_10654);
nand U10863 (N_10863,N_10561,N_10794);
nor U10864 (N_10864,N_10747,N_10749);
nor U10865 (N_10865,N_10616,N_10709);
nor U10866 (N_10866,N_10560,N_10785);
nand U10867 (N_10867,N_10681,N_10745);
and U10868 (N_10868,N_10695,N_10586);
or U10869 (N_10869,N_10767,N_10652);
or U10870 (N_10870,N_10558,N_10539);
xnor U10871 (N_10871,N_10542,N_10731);
or U10872 (N_10872,N_10756,N_10599);
nor U10873 (N_10873,N_10528,N_10761);
xnor U10874 (N_10874,N_10625,N_10765);
and U10875 (N_10875,N_10702,N_10717);
nor U10876 (N_10876,N_10738,N_10553);
nor U10877 (N_10877,N_10611,N_10533);
or U10878 (N_10878,N_10784,N_10564);
or U10879 (N_10879,N_10662,N_10679);
and U10880 (N_10880,N_10657,N_10621);
or U10881 (N_10881,N_10562,N_10686);
or U10882 (N_10882,N_10600,N_10626);
or U10883 (N_10883,N_10527,N_10623);
xnor U10884 (N_10884,N_10620,N_10559);
xnor U10885 (N_10885,N_10726,N_10793);
nor U10886 (N_10886,N_10722,N_10644);
and U10887 (N_10887,N_10788,N_10622);
or U10888 (N_10888,N_10685,N_10509);
or U10889 (N_10889,N_10571,N_10692);
xor U10890 (N_10890,N_10525,N_10720);
or U10891 (N_10891,N_10678,N_10672);
xnor U10892 (N_10892,N_10671,N_10524);
xnor U10893 (N_10893,N_10755,N_10538);
nor U10894 (N_10894,N_10719,N_10526);
xnor U10895 (N_10895,N_10610,N_10502);
xnor U10896 (N_10896,N_10795,N_10667);
nand U10897 (N_10897,N_10504,N_10606);
nor U10898 (N_10898,N_10627,N_10609);
nor U10899 (N_10899,N_10796,N_10596);
or U10900 (N_10900,N_10716,N_10658);
or U10901 (N_10901,N_10577,N_10675);
xor U10902 (N_10902,N_10683,N_10718);
nand U10903 (N_10903,N_10781,N_10647);
or U10904 (N_10904,N_10643,N_10762);
xor U10905 (N_10905,N_10777,N_10546);
or U10906 (N_10906,N_10734,N_10727);
or U10907 (N_10907,N_10684,N_10508);
and U10908 (N_10908,N_10511,N_10601);
and U10909 (N_10909,N_10780,N_10774);
nand U10910 (N_10910,N_10551,N_10578);
nor U10911 (N_10911,N_10584,N_10730);
and U10912 (N_10912,N_10646,N_10752);
nand U10913 (N_10913,N_10515,N_10696);
and U10914 (N_10914,N_10592,N_10624);
nor U10915 (N_10915,N_10563,N_10520);
xor U10916 (N_10916,N_10580,N_10582);
and U10917 (N_10917,N_10540,N_10505);
nand U10918 (N_10918,N_10605,N_10556);
and U10919 (N_10919,N_10693,N_10661);
or U10920 (N_10920,N_10554,N_10523);
and U10921 (N_10921,N_10642,N_10514);
nor U10922 (N_10922,N_10529,N_10748);
nand U10923 (N_10923,N_10618,N_10746);
and U10924 (N_10924,N_10771,N_10650);
xnor U10925 (N_10925,N_10633,N_10522);
and U10926 (N_10926,N_10602,N_10518);
or U10927 (N_10927,N_10589,N_10645);
or U10928 (N_10928,N_10728,N_10543);
nand U10929 (N_10929,N_10742,N_10614);
xor U10930 (N_10930,N_10590,N_10570);
and U10931 (N_10931,N_10663,N_10537);
or U10932 (N_10932,N_10758,N_10567);
xnor U10933 (N_10933,N_10687,N_10603);
xnor U10934 (N_10934,N_10698,N_10591);
xor U10935 (N_10935,N_10612,N_10517);
or U10936 (N_10936,N_10697,N_10653);
or U10937 (N_10937,N_10789,N_10566);
or U10938 (N_10938,N_10743,N_10541);
or U10939 (N_10939,N_10576,N_10670);
xor U10940 (N_10940,N_10581,N_10677);
xor U10941 (N_10941,N_10574,N_10705);
nor U10942 (N_10942,N_10547,N_10766);
xor U10943 (N_10943,N_10615,N_10665);
or U10944 (N_10944,N_10725,N_10569);
or U10945 (N_10945,N_10714,N_10764);
nand U10946 (N_10946,N_10507,N_10629);
or U10947 (N_10947,N_10754,N_10699);
xor U10948 (N_10948,N_10632,N_10630);
nand U10949 (N_10949,N_10763,N_10682);
nand U10950 (N_10950,N_10592,N_10729);
xor U10951 (N_10951,N_10547,N_10654);
or U10952 (N_10952,N_10678,N_10639);
xnor U10953 (N_10953,N_10679,N_10643);
nand U10954 (N_10954,N_10661,N_10586);
nand U10955 (N_10955,N_10678,N_10571);
xnor U10956 (N_10956,N_10745,N_10744);
and U10957 (N_10957,N_10545,N_10617);
nand U10958 (N_10958,N_10676,N_10582);
xnor U10959 (N_10959,N_10771,N_10705);
nor U10960 (N_10960,N_10532,N_10520);
or U10961 (N_10961,N_10668,N_10764);
nand U10962 (N_10962,N_10614,N_10616);
nor U10963 (N_10963,N_10576,N_10565);
xnor U10964 (N_10964,N_10739,N_10642);
or U10965 (N_10965,N_10535,N_10618);
nand U10966 (N_10966,N_10784,N_10591);
and U10967 (N_10967,N_10608,N_10732);
or U10968 (N_10968,N_10721,N_10716);
or U10969 (N_10969,N_10527,N_10710);
nor U10970 (N_10970,N_10666,N_10699);
nand U10971 (N_10971,N_10795,N_10766);
xnor U10972 (N_10972,N_10659,N_10695);
nor U10973 (N_10973,N_10635,N_10545);
and U10974 (N_10974,N_10696,N_10577);
nand U10975 (N_10975,N_10524,N_10783);
nor U10976 (N_10976,N_10705,N_10525);
xnor U10977 (N_10977,N_10679,N_10676);
and U10978 (N_10978,N_10500,N_10540);
nor U10979 (N_10979,N_10747,N_10657);
nor U10980 (N_10980,N_10679,N_10657);
nand U10981 (N_10981,N_10793,N_10691);
nand U10982 (N_10982,N_10542,N_10787);
and U10983 (N_10983,N_10693,N_10719);
nand U10984 (N_10984,N_10602,N_10502);
xnor U10985 (N_10985,N_10767,N_10657);
and U10986 (N_10986,N_10691,N_10777);
or U10987 (N_10987,N_10619,N_10580);
or U10988 (N_10988,N_10625,N_10732);
and U10989 (N_10989,N_10652,N_10502);
nor U10990 (N_10990,N_10758,N_10682);
or U10991 (N_10991,N_10727,N_10654);
nand U10992 (N_10992,N_10600,N_10574);
nand U10993 (N_10993,N_10549,N_10541);
and U10994 (N_10994,N_10596,N_10548);
and U10995 (N_10995,N_10721,N_10751);
and U10996 (N_10996,N_10649,N_10599);
nand U10997 (N_10997,N_10710,N_10523);
or U10998 (N_10998,N_10513,N_10517);
or U10999 (N_10999,N_10705,N_10557);
nand U11000 (N_11000,N_10718,N_10648);
xor U11001 (N_11001,N_10616,N_10593);
xnor U11002 (N_11002,N_10759,N_10507);
and U11003 (N_11003,N_10591,N_10789);
and U11004 (N_11004,N_10695,N_10758);
nor U11005 (N_11005,N_10637,N_10626);
nor U11006 (N_11006,N_10531,N_10628);
xor U11007 (N_11007,N_10687,N_10728);
nor U11008 (N_11008,N_10724,N_10577);
nand U11009 (N_11009,N_10706,N_10789);
nand U11010 (N_11010,N_10777,N_10796);
nand U11011 (N_11011,N_10550,N_10674);
nor U11012 (N_11012,N_10659,N_10720);
or U11013 (N_11013,N_10766,N_10588);
or U11014 (N_11014,N_10707,N_10641);
and U11015 (N_11015,N_10616,N_10503);
nand U11016 (N_11016,N_10516,N_10740);
nand U11017 (N_11017,N_10507,N_10649);
nor U11018 (N_11018,N_10726,N_10760);
xnor U11019 (N_11019,N_10707,N_10751);
nor U11020 (N_11020,N_10591,N_10734);
nand U11021 (N_11021,N_10500,N_10508);
xor U11022 (N_11022,N_10647,N_10765);
nand U11023 (N_11023,N_10601,N_10675);
nand U11024 (N_11024,N_10676,N_10725);
nor U11025 (N_11025,N_10777,N_10635);
nand U11026 (N_11026,N_10585,N_10763);
and U11027 (N_11027,N_10577,N_10533);
nor U11028 (N_11028,N_10786,N_10623);
and U11029 (N_11029,N_10673,N_10574);
xor U11030 (N_11030,N_10503,N_10738);
xor U11031 (N_11031,N_10506,N_10532);
nand U11032 (N_11032,N_10749,N_10717);
nor U11033 (N_11033,N_10582,N_10650);
nor U11034 (N_11034,N_10587,N_10755);
nor U11035 (N_11035,N_10750,N_10765);
nand U11036 (N_11036,N_10595,N_10799);
xnor U11037 (N_11037,N_10770,N_10680);
nor U11038 (N_11038,N_10739,N_10732);
and U11039 (N_11039,N_10750,N_10565);
nor U11040 (N_11040,N_10609,N_10635);
nand U11041 (N_11041,N_10764,N_10566);
or U11042 (N_11042,N_10604,N_10627);
nor U11043 (N_11043,N_10557,N_10738);
and U11044 (N_11044,N_10724,N_10694);
or U11045 (N_11045,N_10614,N_10546);
and U11046 (N_11046,N_10560,N_10789);
and U11047 (N_11047,N_10736,N_10506);
nand U11048 (N_11048,N_10616,N_10781);
nor U11049 (N_11049,N_10626,N_10741);
or U11050 (N_11050,N_10584,N_10551);
xnor U11051 (N_11051,N_10653,N_10717);
nand U11052 (N_11052,N_10777,N_10740);
and U11053 (N_11053,N_10568,N_10556);
nor U11054 (N_11054,N_10616,N_10702);
nand U11055 (N_11055,N_10742,N_10766);
nor U11056 (N_11056,N_10796,N_10568);
or U11057 (N_11057,N_10728,N_10573);
nor U11058 (N_11058,N_10595,N_10714);
or U11059 (N_11059,N_10639,N_10521);
nand U11060 (N_11060,N_10577,N_10641);
xor U11061 (N_11061,N_10656,N_10704);
nor U11062 (N_11062,N_10537,N_10787);
xor U11063 (N_11063,N_10787,N_10535);
or U11064 (N_11064,N_10697,N_10535);
and U11065 (N_11065,N_10535,N_10657);
and U11066 (N_11066,N_10532,N_10708);
nand U11067 (N_11067,N_10541,N_10576);
nand U11068 (N_11068,N_10693,N_10506);
xor U11069 (N_11069,N_10687,N_10723);
nor U11070 (N_11070,N_10537,N_10699);
or U11071 (N_11071,N_10543,N_10777);
and U11072 (N_11072,N_10575,N_10526);
or U11073 (N_11073,N_10610,N_10569);
nor U11074 (N_11074,N_10500,N_10672);
and U11075 (N_11075,N_10509,N_10664);
or U11076 (N_11076,N_10733,N_10608);
or U11077 (N_11077,N_10781,N_10669);
nor U11078 (N_11078,N_10621,N_10552);
nand U11079 (N_11079,N_10761,N_10537);
xnor U11080 (N_11080,N_10538,N_10503);
and U11081 (N_11081,N_10518,N_10524);
and U11082 (N_11082,N_10520,N_10547);
or U11083 (N_11083,N_10723,N_10525);
or U11084 (N_11084,N_10654,N_10742);
and U11085 (N_11085,N_10533,N_10723);
and U11086 (N_11086,N_10522,N_10779);
nand U11087 (N_11087,N_10553,N_10613);
nor U11088 (N_11088,N_10776,N_10771);
nor U11089 (N_11089,N_10623,N_10628);
or U11090 (N_11090,N_10553,N_10579);
or U11091 (N_11091,N_10609,N_10679);
and U11092 (N_11092,N_10545,N_10619);
xnor U11093 (N_11093,N_10566,N_10755);
and U11094 (N_11094,N_10574,N_10767);
and U11095 (N_11095,N_10741,N_10728);
nand U11096 (N_11096,N_10648,N_10510);
and U11097 (N_11097,N_10543,N_10699);
nand U11098 (N_11098,N_10507,N_10593);
nand U11099 (N_11099,N_10571,N_10658);
and U11100 (N_11100,N_11086,N_10802);
and U11101 (N_11101,N_10971,N_10958);
and U11102 (N_11102,N_10817,N_10933);
nand U11103 (N_11103,N_10917,N_10912);
or U11104 (N_11104,N_11098,N_10808);
xnor U11105 (N_11105,N_11078,N_10834);
and U11106 (N_11106,N_11048,N_10998);
or U11107 (N_11107,N_10982,N_11032);
or U11108 (N_11108,N_10919,N_10824);
nor U11109 (N_11109,N_11093,N_10907);
xnor U11110 (N_11110,N_10818,N_11064);
xor U11111 (N_11111,N_11017,N_10828);
nor U11112 (N_11112,N_10858,N_10811);
nand U11113 (N_11113,N_11010,N_11031);
nand U11114 (N_11114,N_10804,N_11035);
xnor U11115 (N_11115,N_10955,N_11057);
and U11116 (N_11116,N_10904,N_10974);
nand U11117 (N_11117,N_10987,N_10978);
nand U11118 (N_11118,N_10908,N_11020);
or U11119 (N_11119,N_10941,N_10999);
xor U11120 (N_11120,N_10867,N_10859);
and U11121 (N_11121,N_10868,N_10961);
nand U11122 (N_11122,N_11019,N_10841);
and U11123 (N_11123,N_10898,N_11099);
nor U11124 (N_11124,N_10969,N_10889);
nor U11125 (N_11125,N_10922,N_10989);
and U11126 (N_11126,N_11083,N_10803);
or U11127 (N_11127,N_11040,N_10927);
nor U11128 (N_11128,N_10945,N_10923);
or U11129 (N_11129,N_10988,N_10994);
or U11130 (N_11130,N_11054,N_10921);
or U11131 (N_11131,N_10997,N_10925);
nor U11132 (N_11132,N_10870,N_11074);
xor U11133 (N_11133,N_11015,N_10881);
nor U11134 (N_11134,N_11034,N_11059);
nand U11135 (N_11135,N_11061,N_10831);
or U11136 (N_11136,N_11039,N_11067);
or U11137 (N_11137,N_11030,N_11055);
or U11138 (N_11138,N_11065,N_10821);
and U11139 (N_11139,N_10950,N_10833);
nand U11140 (N_11140,N_11066,N_10916);
nor U11141 (N_11141,N_11043,N_10822);
and U11142 (N_11142,N_10810,N_11089);
nor U11143 (N_11143,N_11044,N_10943);
or U11144 (N_11144,N_10948,N_10836);
xor U11145 (N_11145,N_10886,N_11016);
or U11146 (N_11146,N_10965,N_10814);
nand U11147 (N_11147,N_11033,N_10806);
and U11148 (N_11148,N_10954,N_10995);
nand U11149 (N_11149,N_10911,N_10844);
nand U11150 (N_11150,N_10897,N_10928);
nand U11151 (N_11151,N_10830,N_10996);
and U11152 (N_11152,N_11041,N_10891);
and U11153 (N_11153,N_10825,N_10873);
nand U11154 (N_11154,N_10871,N_10863);
or U11155 (N_11155,N_10930,N_10918);
nor U11156 (N_11156,N_10937,N_11029);
nor U11157 (N_11157,N_10846,N_10849);
and U11158 (N_11158,N_10915,N_10966);
or U11159 (N_11159,N_11052,N_11011);
or U11160 (N_11160,N_11087,N_10905);
or U11161 (N_11161,N_10843,N_11008);
and U11162 (N_11162,N_10942,N_11051);
and U11163 (N_11163,N_11042,N_10901);
and U11164 (N_11164,N_11005,N_10936);
nand U11165 (N_11165,N_11025,N_10957);
nor U11166 (N_11166,N_10924,N_11081);
or U11167 (N_11167,N_11028,N_11076);
nor U11168 (N_11168,N_10883,N_10894);
xor U11169 (N_11169,N_10862,N_11094);
xnor U11170 (N_11170,N_10837,N_11056);
nor U11171 (N_11171,N_10852,N_10827);
nor U11172 (N_11172,N_10953,N_11072);
and U11173 (N_11173,N_11069,N_11013);
and U11174 (N_11174,N_10812,N_10877);
xnor U11175 (N_11175,N_11018,N_10845);
and U11176 (N_11176,N_10882,N_10880);
and U11177 (N_11177,N_10931,N_10972);
nand U11178 (N_11178,N_10983,N_10888);
nand U11179 (N_11179,N_11082,N_10902);
and U11180 (N_11180,N_10975,N_10885);
xnor U11181 (N_11181,N_11077,N_11026);
or U11182 (N_11182,N_10920,N_10913);
and U11183 (N_11183,N_11000,N_11009);
xnor U11184 (N_11184,N_11097,N_10842);
nand U11185 (N_11185,N_11095,N_11027);
or U11186 (N_11186,N_10856,N_11004);
nand U11187 (N_11187,N_11024,N_11012);
or U11188 (N_11188,N_10850,N_10979);
or U11189 (N_11189,N_10990,N_10986);
or U11190 (N_11190,N_10939,N_10840);
xnor U11191 (N_11191,N_10815,N_10860);
and U11192 (N_11192,N_11038,N_10906);
nor U11193 (N_11193,N_10855,N_10964);
xor U11194 (N_11194,N_11096,N_10847);
and U11195 (N_11195,N_10884,N_11070);
and U11196 (N_11196,N_11002,N_10993);
or U11197 (N_11197,N_10940,N_11080);
nand U11198 (N_11198,N_11058,N_10853);
nand U11199 (N_11199,N_10960,N_10929);
and U11200 (N_11200,N_11014,N_10946);
or U11201 (N_11201,N_10962,N_10878);
nand U11202 (N_11202,N_10984,N_10848);
xnor U11203 (N_11203,N_10952,N_10816);
nor U11204 (N_11204,N_10887,N_10977);
or U11205 (N_11205,N_10820,N_10899);
or U11206 (N_11206,N_10864,N_11036);
or U11207 (N_11207,N_10890,N_10926);
or U11208 (N_11208,N_10963,N_10896);
nor U11209 (N_11209,N_10985,N_11037);
or U11210 (N_11210,N_10823,N_10970);
nor U11211 (N_11211,N_10934,N_11050);
nand U11212 (N_11212,N_11068,N_11046);
and U11213 (N_11213,N_10968,N_10892);
nor U11214 (N_11214,N_10947,N_10809);
nand U11215 (N_11215,N_11085,N_10819);
and U11216 (N_11216,N_10959,N_10938);
nor U11217 (N_11217,N_10976,N_10967);
xor U11218 (N_11218,N_10865,N_10944);
nand U11219 (N_11219,N_11090,N_10932);
nor U11220 (N_11220,N_10876,N_11023);
or U11221 (N_11221,N_10813,N_11063);
nand U11222 (N_11222,N_10903,N_11075);
nor U11223 (N_11223,N_10951,N_10861);
nor U11224 (N_11224,N_10956,N_11079);
nor U11225 (N_11225,N_10869,N_10875);
or U11226 (N_11226,N_11007,N_11060);
nor U11227 (N_11227,N_10992,N_11071);
nand U11228 (N_11228,N_11006,N_10854);
or U11229 (N_11229,N_10893,N_10991);
nor U11230 (N_11230,N_11001,N_10909);
or U11231 (N_11231,N_10866,N_11073);
and U11232 (N_11232,N_11053,N_11022);
nor U11233 (N_11233,N_10805,N_11045);
and U11234 (N_11234,N_10832,N_11049);
or U11235 (N_11235,N_10829,N_10879);
nand U11236 (N_11236,N_11092,N_10980);
or U11237 (N_11237,N_10895,N_11021);
xnor U11238 (N_11238,N_10800,N_11091);
nand U11239 (N_11239,N_11088,N_11047);
nand U11240 (N_11240,N_10949,N_10839);
xor U11241 (N_11241,N_11062,N_10900);
or U11242 (N_11242,N_10835,N_10851);
nor U11243 (N_11243,N_11084,N_10910);
xnor U11244 (N_11244,N_11003,N_10872);
and U11245 (N_11245,N_10801,N_10826);
nor U11246 (N_11246,N_10981,N_10857);
or U11247 (N_11247,N_10807,N_10874);
or U11248 (N_11248,N_10914,N_10973);
nor U11249 (N_11249,N_10935,N_10838);
or U11250 (N_11250,N_10826,N_10871);
or U11251 (N_11251,N_10806,N_10867);
and U11252 (N_11252,N_11005,N_10894);
or U11253 (N_11253,N_10824,N_10900);
or U11254 (N_11254,N_11002,N_11036);
nor U11255 (N_11255,N_10977,N_10944);
or U11256 (N_11256,N_11082,N_11071);
xnor U11257 (N_11257,N_10986,N_11066);
nor U11258 (N_11258,N_10981,N_11079);
xor U11259 (N_11259,N_10896,N_10911);
nand U11260 (N_11260,N_11038,N_10978);
or U11261 (N_11261,N_10911,N_10987);
and U11262 (N_11262,N_11020,N_10800);
and U11263 (N_11263,N_10965,N_10906);
nor U11264 (N_11264,N_10950,N_10992);
nand U11265 (N_11265,N_11006,N_10970);
xor U11266 (N_11266,N_10825,N_10857);
and U11267 (N_11267,N_11024,N_11010);
or U11268 (N_11268,N_11051,N_10845);
xnor U11269 (N_11269,N_10925,N_11043);
nor U11270 (N_11270,N_11022,N_10908);
and U11271 (N_11271,N_11074,N_10835);
nand U11272 (N_11272,N_10878,N_10986);
xnor U11273 (N_11273,N_11022,N_11003);
and U11274 (N_11274,N_10913,N_11002);
xnor U11275 (N_11275,N_10906,N_10959);
or U11276 (N_11276,N_10949,N_11078);
or U11277 (N_11277,N_11091,N_10868);
xor U11278 (N_11278,N_11032,N_10874);
xnor U11279 (N_11279,N_10932,N_10834);
and U11280 (N_11280,N_11015,N_10917);
and U11281 (N_11281,N_10851,N_11057);
and U11282 (N_11282,N_10927,N_10991);
xor U11283 (N_11283,N_11080,N_11062);
xor U11284 (N_11284,N_11088,N_11053);
or U11285 (N_11285,N_10943,N_10808);
xor U11286 (N_11286,N_10811,N_10828);
and U11287 (N_11287,N_11021,N_11046);
and U11288 (N_11288,N_11087,N_10972);
nor U11289 (N_11289,N_10916,N_11049);
nor U11290 (N_11290,N_10874,N_11091);
and U11291 (N_11291,N_10909,N_10994);
nand U11292 (N_11292,N_10950,N_10937);
and U11293 (N_11293,N_10821,N_11092);
nand U11294 (N_11294,N_10809,N_10811);
nor U11295 (N_11295,N_10832,N_10829);
nand U11296 (N_11296,N_11006,N_10917);
xor U11297 (N_11297,N_11047,N_10943);
and U11298 (N_11298,N_11082,N_10814);
nand U11299 (N_11299,N_10845,N_10963);
nor U11300 (N_11300,N_10866,N_10985);
and U11301 (N_11301,N_11066,N_10805);
nand U11302 (N_11302,N_10809,N_10918);
and U11303 (N_11303,N_10989,N_10802);
and U11304 (N_11304,N_10839,N_10907);
or U11305 (N_11305,N_10847,N_10856);
xor U11306 (N_11306,N_10933,N_11060);
xnor U11307 (N_11307,N_10813,N_11019);
xnor U11308 (N_11308,N_10883,N_10951);
or U11309 (N_11309,N_10915,N_10980);
xor U11310 (N_11310,N_10931,N_10801);
and U11311 (N_11311,N_10808,N_10803);
xnor U11312 (N_11312,N_10854,N_11085);
nand U11313 (N_11313,N_10836,N_10926);
and U11314 (N_11314,N_10903,N_10892);
and U11315 (N_11315,N_10885,N_11062);
nand U11316 (N_11316,N_10985,N_11062);
nand U11317 (N_11317,N_11065,N_11008);
nand U11318 (N_11318,N_10982,N_11038);
and U11319 (N_11319,N_10996,N_10893);
xor U11320 (N_11320,N_11046,N_10937);
and U11321 (N_11321,N_10834,N_10824);
nand U11322 (N_11322,N_11093,N_11054);
nand U11323 (N_11323,N_11022,N_10918);
xor U11324 (N_11324,N_10851,N_10854);
and U11325 (N_11325,N_10960,N_10883);
nor U11326 (N_11326,N_11029,N_10858);
nor U11327 (N_11327,N_10875,N_11034);
or U11328 (N_11328,N_10846,N_11046);
nand U11329 (N_11329,N_10835,N_10826);
nor U11330 (N_11330,N_10910,N_11054);
xnor U11331 (N_11331,N_10858,N_11083);
or U11332 (N_11332,N_10850,N_10924);
nor U11333 (N_11333,N_11039,N_10920);
or U11334 (N_11334,N_10866,N_11007);
nor U11335 (N_11335,N_10917,N_10837);
nand U11336 (N_11336,N_11012,N_11044);
nor U11337 (N_11337,N_10899,N_10980);
xnor U11338 (N_11338,N_11044,N_11059);
nor U11339 (N_11339,N_10864,N_10815);
or U11340 (N_11340,N_11062,N_10911);
and U11341 (N_11341,N_10982,N_10814);
and U11342 (N_11342,N_11045,N_10837);
nor U11343 (N_11343,N_11033,N_10839);
nand U11344 (N_11344,N_11045,N_11027);
nand U11345 (N_11345,N_10933,N_10843);
xor U11346 (N_11346,N_10915,N_10900);
or U11347 (N_11347,N_10911,N_10891);
nor U11348 (N_11348,N_11005,N_10938);
nand U11349 (N_11349,N_10866,N_10955);
nor U11350 (N_11350,N_10860,N_11047);
xor U11351 (N_11351,N_10814,N_11011);
xor U11352 (N_11352,N_10850,N_10973);
xnor U11353 (N_11353,N_10953,N_11047);
nor U11354 (N_11354,N_10837,N_10852);
nor U11355 (N_11355,N_10885,N_10855);
and U11356 (N_11356,N_10949,N_10983);
or U11357 (N_11357,N_11071,N_11027);
nor U11358 (N_11358,N_10958,N_10927);
nor U11359 (N_11359,N_11094,N_11088);
or U11360 (N_11360,N_10840,N_10872);
nor U11361 (N_11361,N_11038,N_11001);
and U11362 (N_11362,N_10989,N_11096);
nand U11363 (N_11363,N_11094,N_10802);
or U11364 (N_11364,N_10950,N_10848);
xor U11365 (N_11365,N_11006,N_10926);
nand U11366 (N_11366,N_11084,N_11093);
and U11367 (N_11367,N_10836,N_10870);
or U11368 (N_11368,N_10885,N_10815);
or U11369 (N_11369,N_10938,N_11022);
xnor U11370 (N_11370,N_10871,N_10869);
xor U11371 (N_11371,N_10844,N_11068);
and U11372 (N_11372,N_11013,N_10809);
nand U11373 (N_11373,N_10922,N_10930);
nand U11374 (N_11374,N_10920,N_10960);
nor U11375 (N_11375,N_10978,N_11098);
or U11376 (N_11376,N_11079,N_10954);
or U11377 (N_11377,N_10892,N_10829);
or U11378 (N_11378,N_11068,N_11093);
nor U11379 (N_11379,N_11004,N_11005);
nand U11380 (N_11380,N_10961,N_10927);
or U11381 (N_11381,N_10910,N_11040);
and U11382 (N_11382,N_10839,N_10917);
nand U11383 (N_11383,N_10958,N_10957);
and U11384 (N_11384,N_10979,N_10852);
xor U11385 (N_11385,N_11082,N_10819);
or U11386 (N_11386,N_10946,N_10916);
or U11387 (N_11387,N_10972,N_10835);
and U11388 (N_11388,N_10931,N_10920);
nor U11389 (N_11389,N_10810,N_10922);
xnor U11390 (N_11390,N_10818,N_10857);
and U11391 (N_11391,N_10817,N_11019);
nor U11392 (N_11392,N_11097,N_10924);
or U11393 (N_11393,N_10867,N_10974);
nand U11394 (N_11394,N_11002,N_11048);
nor U11395 (N_11395,N_11045,N_10989);
or U11396 (N_11396,N_10876,N_11064);
nor U11397 (N_11397,N_10830,N_10936);
xor U11398 (N_11398,N_11065,N_11096);
or U11399 (N_11399,N_10991,N_11020);
nor U11400 (N_11400,N_11375,N_11309);
and U11401 (N_11401,N_11185,N_11337);
and U11402 (N_11402,N_11217,N_11192);
xnor U11403 (N_11403,N_11108,N_11248);
and U11404 (N_11404,N_11273,N_11176);
and U11405 (N_11405,N_11119,N_11154);
xor U11406 (N_11406,N_11310,N_11268);
nor U11407 (N_11407,N_11172,N_11286);
xnor U11408 (N_11408,N_11346,N_11347);
nand U11409 (N_11409,N_11103,N_11226);
nor U11410 (N_11410,N_11153,N_11137);
xor U11411 (N_11411,N_11323,N_11136);
or U11412 (N_11412,N_11167,N_11304);
nand U11413 (N_11413,N_11160,N_11203);
nand U11414 (N_11414,N_11210,N_11300);
xor U11415 (N_11415,N_11101,N_11275);
or U11416 (N_11416,N_11385,N_11276);
or U11417 (N_11417,N_11123,N_11259);
and U11418 (N_11418,N_11313,N_11311);
or U11419 (N_11419,N_11209,N_11132);
and U11420 (N_11420,N_11205,N_11228);
or U11421 (N_11421,N_11158,N_11324);
xnor U11422 (N_11422,N_11356,N_11229);
xor U11423 (N_11423,N_11339,N_11332);
xnor U11424 (N_11424,N_11283,N_11100);
and U11425 (N_11425,N_11193,N_11117);
xnor U11426 (N_11426,N_11178,N_11340);
xnor U11427 (N_11427,N_11115,N_11186);
or U11428 (N_11428,N_11204,N_11124);
xor U11429 (N_11429,N_11298,N_11317);
or U11430 (N_11430,N_11378,N_11355);
and U11431 (N_11431,N_11107,N_11291);
nor U11432 (N_11432,N_11348,N_11157);
xnor U11433 (N_11433,N_11195,N_11365);
nor U11434 (N_11434,N_11395,N_11327);
nand U11435 (N_11435,N_11263,N_11322);
and U11436 (N_11436,N_11230,N_11345);
nor U11437 (N_11437,N_11338,N_11179);
nand U11438 (N_11438,N_11373,N_11280);
or U11439 (N_11439,N_11211,N_11398);
nor U11440 (N_11440,N_11353,N_11325);
nor U11441 (N_11441,N_11238,N_11125);
and U11442 (N_11442,N_11218,N_11162);
or U11443 (N_11443,N_11381,N_11244);
or U11444 (N_11444,N_11138,N_11223);
or U11445 (N_11445,N_11106,N_11140);
or U11446 (N_11446,N_11155,N_11234);
xor U11447 (N_11447,N_11364,N_11253);
xor U11448 (N_11448,N_11191,N_11301);
and U11449 (N_11449,N_11333,N_11202);
and U11450 (N_11450,N_11299,N_11374);
nand U11451 (N_11451,N_11328,N_11199);
xor U11452 (N_11452,N_11342,N_11251);
xor U11453 (N_11453,N_11190,N_11216);
nor U11454 (N_11454,N_11113,N_11254);
nor U11455 (N_11455,N_11267,N_11261);
or U11456 (N_11456,N_11279,N_11116);
and U11457 (N_11457,N_11366,N_11393);
or U11458 (N_11458,N_11219,N_11330);
xnor U11459 (N_11459,N_11163,N_11145);
and U11460 (N_11460,N_11245,N_11307);
xnor U11461 (N_11461,N_11148,N_11169);
or U11462 (N_11462,N_11387,N_11196);
xnor U11463 (N_11463,N_11128,N_11344);
nor U11464 (N_11464,N_11105,N_11308);
or U11465 (N_11465,N_11319,N_11367);
nand U11466 (N_11466,N_11264,N_11232);
xor U11467 (N_11467,N_11371,N_11239);
and U11468 (N_11468,N_11392,N_11187);
nand U11469 (N_11469,N_11351,N_11326);
xnor U11470 (N_11470,N_11354,N_11135);
or U11471 (N_11471,N_11220,N_11359);
xor U11472 (N_11472,N_11134,N_11201);
xnor U11473 (N_11473,N_11290,N_11151);
nor U11474 (N_11474,N_11177,N_11331);
and U11475 (N_11475,N_11272,N_11156);
nor U11476 (N_11476,N_11255,N_11379);
and U11477 (N_11477,N_11293,N_11233);
nor U11478 (N_11478,N_11215,N_11122);
and U11479 (N_11479,N_11189,N_11181);
and U11480 (N_11480,N_11321,N_11121);
nand U11481 (N_11481,N_11270,N_11109);
xor U11482 (N_11482,N_11399,N_11329);
nand U11483 (N_11483,N_11315,N_11320);
nor U11484 (N_11484,N_11335,N_11242);
nor U11485 (N_11485,N_11287,N_11341);
and U11486 (N_11486,N_11118,N_11237);
and U11487 (N_11487,N_11266,N_11377);
xnor U11488 (N_11488,N_11278,N_11188);
xnor U11489 (N_11489,N_11173,N_11386);
xnor U11490 (N_11490,N_11182,N_11357);
and U11491 (N_11491,N_11164,N_11257);
or U11492 (N_11492,N_11390,N_11152);
and U11493 (N_11493,N_11388,N_11295);
and U11494 (N_11494,N_11197,N_11296);
or U11495 (N_11495,N_11394,N_11144);
or U11496 (N_11496,N_11288,N_11258);
nand U11497 (N_11497,N_11174,N_11363);
or U11498 (N_11498,N_11168,N_11126);
and U11499 (N_11499,N_11284,N_11170);
or U11500 (N_11500,N_11120,N_11235);
nor U11501 (N_11501,N_11246,N_11262);
nand U11502 (N_11502,N_11352,N_11391);
or U11503 (N_11503,N_11360,N_11149);
nand U11504 (N_11504,N_11249,N_11200);
xnor U11505 (N_11505,N_11269,N_11225);
nor U11506 (N_11506,N_11382,N_11133);
xor U11507 (N_11507,N_11396,N_11147);
nand U11508 (N_11508,N_11243,N_11349);
nand U11509 (N_11509,N_11165,N_11343);
nor U11510 (N_11510,N_11104,N_11102);
nor U11511 (N_11511,N_11130,N_11383);
and U11512 (N_11512,N_11368,N_11369);
nor U11513 (N_11513,N_11302,N_11236);
nor U11514 (N_11514,N_11183,N_11376);
and U11515 (N_11515,N_11142,N_11171);
nand U11516 (N_11516,N_11265,N_11362);
xor U11517 (N_11517,N_11334,N_11316);
or U11518 (N_11518,N_11127,N_11141);
nand U11519 (N_11519,N_11252,N_11240);
nor U11520 (N_11520,N_11175,N_11110);
or U11521 (N_11521,N_11282,N_11358);
nand U11522 (N_11522,N_11336,N_11297);
or U11523 (N_11523,N_11274,N_11350);
and U11524 (N_11524,N_11370,N_11389);
and U11525 (N_11525,N_11146,N_11212);
nand U11526 (N_11526,N_11111,N_11114);
or U11527 (N_11527,N_11112,N_11221);
nand U11528 (N_11528,N_11372,N_11198);
and U11529 (N_11529,N_11247,N_11161);
nand U11530 (N_11530,N_11271,N_11285);
nor U11531 (N_11531,N_11131,N_11281);
or U11532 (N_11532,N_11256,N_11312);
or U11533 (N_11533,N_11213,N_11361);
nand U11534 (N_11534,N_11306,N_11305);
and U11535 (N_11535,N_11314,N_11289);
nor U11536 (N_11536,N_11206,N_11384);
nor U11537 (N_11537,N_11260,N_11184);
and U11538 (N_11538,N_11292,N_11139);
xor U11539 (N_11539,N_11303,N_11214);
and U11540 (N_11540,N_11208,N_11143);
nand U11541 (N_11541,N_11380,N_11277);
nand U11542 (N_11542,N_11194,N_11129);
or U11543 (N_11543,N_11150,N_11159);
nor U11544 (N_11544,N_11166,N_11250);
and U11545 (N_11545,N_11227,N_11224);
and U11546 (N_11546,N_11207,N_11318);
nand U11547 (N_11547,N_11180,N_11294);
nor U11548 (N_11548,N_11241,N_11397);
nor U11549 (N_11549,N_11231,N_11222);
nor U11550 (N_11550,N_11297,N_11226);
or U11551 (N_11551,N_11297,N_11306);
nand U11552 (N_11552,N_11374,N_11366);
xor U11553 (N_11553,N_11262,N_11149);
and U11554 (N_11554,N_11118,N_11170);
nor U11555 (N_11555,N_11397,N_11372);
nand U11556 (N_11556,N_11390,N_11176);
or U11557 (N_11557,N_11293,N_11245);
and U11558 (N_11558,N_11308,N_11398);
and U11559 (N_11559,N_11226,N_11236);
xor U11560 (N_11560,N_11284,N_11185);
nor U11561 (N_11561,N_11143,N_11213);
nor U11562 (N_11562,N_11154,N_11352);
and U11563 (N_11563,N_11131,N_11361);
or U11564 (N_11564,N_11318,N_11315);
xor U11565 (N_11565,N_11261,N_11194);
nor U11566 (N_11566,N_11322,N_11292);
nand U11567 (N_11567,N_11138,N_11397);
xor U11568 (N_11568,N_11253,N_11388);
nor U11569 (N_11569,N_11215,N_11262);
or U11570 (N_11570,N_11268,N_11349);
and U11571 (N_11571,N_11212,N_11334);
and U11572 (N_11572,N_11169,N_11267);
and U11573 (N_11573,N_11111,N_11240);
and U11574 (N_11574,N_11382,N_11312);
or U11575 (N_11575,N_11334,N_11115);
xnor U11576 (N_11576,N_11204,N_11307);
nand U11577 (N_11577,N_11319,N_11125);
nor U11578 (N_11578,N_11105,N_11394);
and U11579 (N_11579,N_11327,N_11355);
nand U11580 (N_11580,N_11170,N_11275);
and U11581 (N_11581,N_11308,N_11129);
xor U11582 (N_11582,N_11295,N_11331);
nand U11583 (N_11583,N_11264,N_11287);
and U11584 (N_11584,N_11383,N_11278);
xor U11585 (N_11585,N_11318,N_11122);
nand U11586 (N_11586,N_11347,N_11173);
xnor U11587 (N_11587,N_11149,N_11190);
xor U11588 (N_11588,N_11117,N_11322);
nor U11589 (N_11589,N_11356,N_11176);
nand U11590 (N_11590,N_11190,N_11196);
and U11591 (N_11591,N_11202,N_11339);
or U11592 (N_11592,N_11169,N_11307);
nor U11593 (N_11593,N_11156,N_11381);
and U11594 (N_11594,N_11250,N_11218);
or U11595 (N_11595,N_11133,N_11343);
and U11596 (N_11596,N_11335,N_11156);
nand U11597 (N_11597,N_11211,N_11231);
xor U11598 (N_11598,N_11310,N_11367);
or U11599 (N_11599,N_11246,N_11141);
xor U11600 (N_11600,N_11245,N_11394);
xor U11601 (N_11601,N_11293,N_11392);
or U11602 (N_11602,N_11223,N_11272);
xnor U11603 (N_11603,N_11387,N_11279);
nand U11604 (N_11604,N_11359,N_11207);
or U11605 (N_11605,N_11147,N_11239);
nor U11606 (N_11606,N_11121,N_11343);
and U11607 (N_11607,N_11357,N_11286);
nand U11608 (N_11608,N_11334,N_11331);
xor U11609 (N_11609,N_11342,N_11226);
and U11610 (N_11610,N_11210,N_11192);
nor U11611 (N_11611,N_11366,N_11243);
nand U11612 (N_11612,N_11202,N_11256);
xnor U11613 (N_11613,N_11334,N_11251);
nor U11614 (N_11614,N_11372,N_11175);
or U11615 (N_11615,N_11178,N_11308);
nor U11616 (N_11616,N_11156,N_11220);
or U11617 (N_11617,N_11291,N_11283);
nand U11618 (N_11618,N_11134,N_11256);
and U11619 (N_11619,N_11207,N_11372);
xnor U11620 (N_11620,N_11284,N_11173);
or U11621 (N_11621,N_11240,N_11340);
xor U11622 (N_11622,N_11208,N_11172);
nand U11623 (N_11623,N_11390,N_11233);
and U11624 (N_11624,N_11304,N_11386);
and U11625 (N_11625,N_11279,N_11360);
nand U11626 (N_11626,N_11317,N_11218);
or U11627 (N_11627,N_11336,N_11162);
xor U11628 (N_11628,N_11143,N_11192);
and U11629 (N_11629,N_11182,N_11189);
xor U11630 (N_11630,N_11135,N_11181);
and U11631 (N_11631,N_11206,N_11287);
nand U11632 (N_11632,N_11217,N_11189);
and U11633 (N_11633,N_11260,N_11222);
nand U11634 (N_11634,N_11236,N_11231);
nand U11635 (N_11635,N_11358,N_11383);
nand U11636 (N_11636,N_11164,N_11126);
or U11637 (N_11637,N_11267,N_11159);
or U11638 (N_11638,N_11369,N_11271);
or U11639 (N_11639,N_11329,N_11295);
xnor U11640 (N_11640,N_11299,N_11342);
nand U11641 (N_11641,N_11298,N_11268);
and U11642 (N_11642,N_11147,N_11336);
nand U11643 (N_11643,N_11313,N_11382);
or U11644 (N_11644,N_11310,N_11314);
xnor U11645 (N_11645,N_11292,N_11161);
nand U11646 (N_11646,N_11378,N_11292);
nand U11647 (N_11647,N_11230,N_11228);
nand U11648 (N_11648,N_11274,N_11374);
nor U11649 (N_11649,N_11163,N_11178);
nand U11650 (N_11650,N_11255,N_11118);
or U11651 (N_11651,N_11190,N_11313);
and U11652 (N_11652,N_11336,N_11270);
and U11653 (N_11653,N_11322,N_11392);
and U11654 (N_11654,N_11196,N_11314);
nor U11655 (N_11655,N_11289,N_11255);
xor U11656 (N_11656,N_11352,N_11271);
xnor U11657 (N_11657,N_11387,N_11128);
xor U11658 (N_11658,N_11268,N_11321);
nand U11659 (N_11659,N_11263,N_11159);
nand U11660 (N_11660,N_11262,N_11311);
nand U11661 (N_11661,N_11311,N_11336);
nand U11662 (N_11662,N_11172,N_11388);
nor U11663 (N_11663,N_11265,N_11255);
xnor U11664 (N_11664,N_11214,N_11139);
xor U11665 (N_11665,N_11314,N_11393);
nand U11666 (N_11666,N_11337,N_11323);
nor U11667 (N_11667,N_11174,N_11107);
and U11668 (N_11668,N_11237,N_11267);
nand U11669 (N_11669,N_11236,N_11338);
or U11670 (N_11670,N_11289,N_11166);
and U11671 (N_11671,N_11226,N_11360);
nor U11672 (N_11672,N_11333,N_11102);
nand U11673 (N_11673,N_11276,N_11226);
xnor U11674 (N_11674,N_11373,N_11224);
and U11675 (N_11675,N_11244,N_11170);
xor U11676 (N_11676,N_11380,N_11166);
nand U11677 (N_11677,N_11293,N_11324);
nor U11678 (N_11678,N_11227,N_11391);
xor U11679 (N_11679,N_11335,N_11255);
xor U11680 (N_11680,N_11224,N_11391);
or U11681 (N_11681,N_11334,N_11242);
and U11682 (N_11682,N_11330,N_11125);
and U11683 (N_11683,N_11210,N_11321);
xnor U11684 (N_11684,N_11369,N_11109);
xor U11685 (N_11685,N_11367,N_11315);
xnor U11686 (N_11686,N_11284,N_11176);
xor U11687 (N_11687,N_11236,N_11391);
or U11688 (N_11688,N_11287,N_11197);
xor U11689 (N_11689,N_11371,N_11284);
nand U11690 (N_11690,N_11102,N_11339);
xor U11691 (N_11691,N_11273,N_11278);
nand U11692 (N_11692,N_11111,N_11160);
nand U11693 (N_11693,N_11379,N_11127);
or U11694 (N_11694,N_11222,N_11325);
xnor U11695 (N_11695,N_11309,N_11189);
and U11696 (N_11696,N_11280,N_11128);
or U11697 (N_11697,N_11156,N_11200);
xor U11698 (N_11698,N_11276,N_11315);
and U11699 (N_11699,N_11257,N_11251);
and U11700 (N_11700,N_11685,N_11612);
xnor U11701 (N_11701,N_11515,N_11680);
xnor U11702 (N_11702,N_11644,N_11616);
xor U11703 (N_11703,N_11671,N_11655);
nor U11704 (N_11704,N_11444,N_11578);
and U11705 (N_11705,N_11535,N_11404);
or U11706 (N_11706,N_11467,N_11646);
nand U11707 (N_11707,N_11417,N_11519);
nand U11708 (N_11708,N_11476,N_11419);
xnor U11709 (N_11709,N_11403,N_11422);
nor U11710 (N_11710,N_11654,N_11457);
or U11711 (N_11711,N_11401,N_11672);
or U11712 (N_11712,N_11479,N_11659);
nand U11713 (N_11713,N_11536,N_11562);
and U11714 (N_11714,N_11673,N_11491);
nand U11715 (N_11715,N_11682,N_11584);
nand U11716 (N_11716,N_11617,N_11500);
nor U11717 (N_11717,N_11527,N_11429);
or U11718 (N_11718,N_11495,N_11540);
or U11719 (N_11719,N_11697,N_11549);
and U11720 (N_11720,N_11413,N_11447);
or U11721 (N_11721,N_11624,N_11473);
nand U11722 (N_11722,N_11451,N_11454);
xor U11723 (N_11723,N_11468,N_11516);
and U11724 (N_11724,N_11592,N_11580);
or U11725 (N_11725,N_11640,N_11565);
nor U11726 (N_11726,N_11698,N_11690);
nand U11727 (N_11727,N_11656,N_11475);
and U11728 (N_11728,N_11657,N_11517);
nor U11729 (N_11729,N_11537,N_11525);
nor U11730 (N_11730,N_11554,N_11507);
nor U11731 (N_11731,N_11464,N_11606);
nor U11732 (N_11732,N_11650,N_11570);
nor U11733 (N_11733,N_11689,N_11676);
nor U11734 (N_11734,N_11618,N_11424);
nand U11735 (N_11735,N_11423,N_11414);
xnor U11736 (N_11736,N_11534,N_11684);
and U11737 (N_11737,N_11550,N_11649);
xor U11738 (N_11738,N_11572,N_11552);
nand U11739 (N_11739,N_11492,N_11607);
and U11740 (N_11740,N_11462,N_11437);
nand U11741 (N_11741,N_11501,N_11586);
or U11742 (N_11742,N_11663,N_11566);
nand U11743 (N_11743,N_11555,N_11531);
or U11744 (N_11744,N_11510,N_11440);
or U11745 (N_11745,N_11506,N_11641);
xnor U11746 (N_11746,N_11452,N_11629);
nand U11747 (N_11747,N_11613,N_11508);
nor U11748 (N_11748,N_11483,N_11596);
and U11749 (N_11749,N_11463,N_11493);
and U11750 (N_11750,N_11469,N_11683);
nor U11751 (N_11751,N_11472,N_11605);
and U11752 (N_11752,N_11509,N_11643);
nand U11753 (N_11753,N_11590,N_11518);
nor U11754 (N_11754,N_11427,N_11597);
nand U11755 (N_11755,N_11405,N_11648);
and U11756 (N_11756,N_11577,N_11474);
nor U11757 (N_11757,N_11647,N_11660);
or U11758 (N_11758,N_11695,N_11620);
xor U11759 (N_11759,N_11634,N_11412);
nor U11760 (N_11760,N_11441,N_11528);
nor U11761 (N_11761,N_11511,N_11622);
nand U11762 (N_11762,N_11557,N_11670);
nor U11763 (N_11763,N_11665,N_11686);
nor U11764 (N_11764,N_11445,N_11489);
and U11765 (N_11765,N_11425,N_11579);
and U11766 (N_11766,N_11520,N_11539);
and U11767 (N_11767,N_11521,N_11411);
or U11768 (N_11768,N_11533,N_11679);
nand U11769 (N_11769,N_11594,N_11633);
nand U11770 (N_11770,N_11436,N_11446);
or U11771 (N_11771,N_11547,N_11455);
nand U11772 (N_11772,N_11421,N_11658);
or U11773 (N_11773,N_11443,N_11482);
nor U11774 (N_11774,N_11526,N_11621);
xnor U11775 (N_11775,N_11544,N_11564);
nor U11776 (N_11776,N_11627,N_11573);
and U11777 (N_11777,N_11448,N_11558);
nor U11778 (N_11778,N_11439,N_11639);
nor U11779 (N_11779,N_11691,N_11593);
nor U11780 (N_11780,N_11494,N_11402);
and U11781 (N_11781,N_11611,N_11490);
xor U11782 (N_11782,N_11460,N_11434);
nand U11783 (N_11783,N_11522,N_11466);
nor U11784 (N_11784,N_11487,N_11523);
nand U11785 (N_11785,N_11610,N_11631);
xor U11786 (N_11786,N_11438,N_11688);
nor U11787 (N_11787,N_11503,N_11532);
or U11788 (N_11788,N_11635,N_11693);
nand U11789 (N_11789,N_11585,N_11602);
nor U11790 (N_11790,N_11435,N_11505);
or U11791 (N_11791,N_11677,N_11678);
or U11792 (N_11792,N_11478,N_11553);
xor U11793 (N_11793,N_11645,N_11458);
nor U11794 (N_11794,N_11662,N_11615);
nor U11795 (N_11795,N_11530,N_11433);
nor U11796 (N_11796,N_11407,N_11614);
or U11797 (N_11797,N_11696,N_11582);
nand U11798 (N_11798,N_11496,N_11569);
nand U11799 (N_11799,N_11461,N_11420);
and U11800 (N_11800,N_11588,N_11410);
xor U11801 (N_11801,N_11484,N_11674);
nor U11802 (N_11802,N_11636,N_11603);
nand U11803 (N_11803,N_11485,N_11587);
or U11804 (N_11804,N_11431,N_11668);
nand U11805 (N_11805,N_11524,N_11556);
nand U11806 (N_11806,N_11449,N_11514);
nor U11807 (N_11807,N_11571,N_11669);
nand U11808 (N_11808,N_11651,N_11652);
nor U11809 (N_11809,N_11542,N_11661);
and U11810 (N_11810,N_11513,N_11504);
or U11811 (N_11811,N_11575,N_11546);
or U11812 (N_11812,N_11545,N_11456);
and U11813 (N_11813,N_11459,N_11625);
nand U11814 (N_11814,N_11687,N_11529);
nand U11815 (N_11815,N_11589,N_11400);
nand U11816 (N_11816,N_11664,N_11637);
nor U11817 (N_11817,N_11415,N_11470);
or U11818 (N_11818,N_11595,N_11450);
and U11819 (N_11819,N_11428,N_11653);
nor U11820 (N_11820,N_11626,N_11694);
nand U11821 (N_11821,N_11583,N_11481);
xor U11822 (N_11822,N_11442,N_11416);
nor U11823 (N_11823,N_11609,N_11601);
or U11824 (N_11824,N_11465,N_11608);
or U11825 (N_11825,N_11541,N_11543);
or U11826 (N_11826,N_11551,N_11600);
xor U11827 (N_11827,N_11567,N_11591);
and U11828 (N_11828,N_11430,N_11632);
and U11829 (N_11829,N_11560,N_11408);
or U11830 (N_11830,N_11574,N_11512);
or U11831 (N_11831,N_11628,N_11406);
and U11832 (N_11832,N_11681,N_11502);
or U11833 (N_11833,N_11498,N_11638);
xor U11834 (N_11834,N_11548,N_11561);
nor U11835 (N_11835,N_11599,N_11568);
nor U11836 (N_11836,N_11642,N_11619);
or U11837 (N_11837,N_11563,N_11630);
or U11838 (N_11838,N_11598,N_11418);
and U11839 (N_11839,N_11559,N_11477);
xor U11840 (N_11840,N_11623,N_11486);
nor U11841 (N_11841,N_11604,N_11581);
xor U11842 (N_11842,N_11426,N_11409);
nor U11843 (N_11843,N_11480,N_11453);
xnor U11844 (N_11844,N_11576,N_11499);
or U11845 (N_11845,N_11432,N_11675);
and U11846 (N_11846,N_11666,N_11699);
or U11847 (N_11847,N_11497,N_11538);
or U11848 (N_11848,N_11488,N_11692);
and U11849 (N_11849,N_11471,N_11667);
nor U11850 (N_11850,N_11536,N_11475);
nor U11851 (N_11851,N_11578,N_11454);
and U11852 (N_11852,N_11408,N_11420);
nand U11853 (N_11853,N_11574,N_11481);
or U11854 (N_11854,N_11587,N_11667);
and U11855 (N_11855,N_11582,N_11563);
xnor U11856 (N_11856,N_11520,N_11685);
or U11857 (N_11857,N_11565,N_11490);
and U11858 (N_11858,N_11689,N_11633);
xnor U11859 (N_11859,N_11662,N_11684);
nor U11860 (N_11860,N_11649,N_11402);
nor U11861 (N_11861,N_11464,N_11401);
nand U11862 (N_11862,N_11550,N_11545);
xnor U11863 (N_11863,N_11680,N_11528);
nand U11864 (N_11864,N_11493,N_11496);
or U11865 (N_11865,N_11554,N_11603);
xnor U11866 (N_11866,N_11646,N_11556);
or U11867 (N_11867,N_11531,N_11592);
xor U11868 (N_11868,N_11639,N_11506);
xor U11869 (N_11869,N_11679,N_11573);
xor U11870 (N_11870,N_11592,N_11600);
xor U11871 (N_11871,N_11634,N_11698);
or U11872 (N_11872,N_11554,N_11597);
xor U11873 (N_11873,N_11434,N_11510);
nand U11874 (N_11874,N_11558,N_11679);
and U11875 (N_11875,N_11487,N_11621);
or U11876 (N_11876,N_11592,N_11442);
nand U11877 (N_11877,N_11434,N_11598);
and U11878 (N_11878,N_11629,N_11447);
and U11879 (N_11879,N_11685,N_11445);
and U11880 (N_11880,N_11610,N_11657);
xor U11881 (N_11881,N_11680,N_11467);
and U11882 (N_11882,N_11468,N_11636);
or U11883 (N_11883,N_11459,N_11536);
nor U11884 (N_11884,N_11420,N_11445);
xnor U11885 (N_11885,N_11458,N_11445);
and U11886 (N_11886,N_11519,N_11517);
xor U11887 (N_11887,N_11628,N_11495);
and U11888 (N_11888,N_11447,N_11656);
or U11889 (N_11889,N_11446,N_11573);
nor U11890 (N_11890,N_11572,N_11515);
xor U11891 (N_11891,N_11668,N_11423);
or U11892 (N_11892,N_11444,N_11512);
and U11893 (N_11893,N_11424,N_11488);
xor U11894 (N_11894,N_11665,N_11407);
and U11895 (N_11895,N_11607,N_11426);
xor U11896 (N_11896,N_11653,N_11621);
or U11897 (N_11897,N_11518,N_11695);
nor U11898 (N_11898,N_11586,N_11691);
nand U11899 (N_11899,N_11613,N_11452);
nand U11900 (N_11900,N_11524,N_11544);
or U11901 (N_11901,N_11504,N_11434);
nand U11902 (N_11902,N_11488,N_11570);
nor U11903 (N_11903,N_11444,N_11412);
nand U11904 (N_11904,N_11583,N_11589);
nand U11905 (N_11905,N_11633,N_11471);
nor U11906 (N_11906,N_11536,N_11401);
nor U11907 (N_11907,N_11612,N_11687);
or U11908 (N_11908,N_11646,N_11600);
nand U11909 (N_11909,N_11495,N_11433);
nand U11910 (N_11910,N_11577,N_11476);
or U11911 (N_11911,N_11582,N_11523);
and U11912 (N_11912,N_11472,N_11669);
nand U11913 (N_11913,N_11575,N_11488);
xor U11914 (N_11914,N_11437,N_11535);
and U11915 (N_11915,N_11596,N_11490);
and U11916 (N_11916,N_11600,N_11457);
xor U11917 (N_11917,N_11513,N_11542);
or U11918 (N_11918,N_11681,N_11613);
nor U11919 (N_11919,N_11405,N_11475);
or U11920 (N_11920,N_11453,N_11407);
nand U11921 (N_11921,N_11439,N_11549);
xnor U11922 (N_11922,N_11440,N_11479);
or U11923 (N_11923,N_11622,N_11693);
and U11924 (N_11924,N_11570,N_11514);
nor U11925 (N_11925,N_11482,N_11506);
xor U11926 (N_11926,N_11449,N_11498);
nand U11927 (N_11927,N_11545,N_11471);
xor U11928 (N_11928,N_11440,N_11580);
and U11929 (N_11929,N_11525,N_11468);
nor U11930 (N_11930,N_11633,N_11568);
and U11931 (N_11931,N_11536,N_11586);
or U11932 (N_11932,N_11659,N_11476);
xor U11933 (N_11933,N_11647,N_11436);
xnor U11934 (N_11934,N_11675,N_11413);
or U11935 (N_11935,N_11565,N_11575);
and U11936 (N_11936,N_11524,N_11624);
and U11937 (N_11937,N_11611,N_11687);
nor U11938 (N_11938,N_11463,N_11640);
xor U11939 (N_11939,N_11677,N_11406);
and U11940 (N_11940,N_11473,N_11577);
and U11941 (N_11941,N_11523,N_11415);
nand U11942 (N_11942,N_11409,N_11525);
and U11943 (N_11943,N_11420,N_11493);
xnor U11944 (N_11944,N_11455,N_11555);
nand U11945 (N_11945,N_11401,N_11544);
or U11946 (N_11946,N_11439,N_11569);
nor U11947 (N_11947,N_11654,N_11521);
xnor U11948 (N_11948,N_11634,N_11539);
xnor U11949 (N_11949,N_11605,N_11591);
or U11950 (N_11950,N_11608,N_11686);
nor U11951 (N_11951,N_11635,N_11427);
nand U11952 (N_11952,N_11471,N_11468);
or U11953 (N_11953,N_11457,N_11610);
or U11954 (N_11954,N_11690,N_11446);
nand U11955 (N_11955,N_11479,N_11637);
and U11956 (N_11956,N_11538,N_11625);
or U11957 (N_11957,N_11646,N_11445);
and U11958 (N_11958,N_11532,N_11692);
nor U11959 (N_11959,N_11601,N_11598);
and U11960 (N_11960,N_11452,N_11619);
or U11961 (N_11961,N_11655,N_11446);
xor U11962 (N_11962,N_11505,N_11626);
nand U11963 (N_11963,N_11612,N_11643);
and U11964 (N_11964,N_11522,N_11449);
nor U11965 (N_11965,N_11416,N_11624);
nor U11966 (N_11966,N_11663,N_11447);
and U11967 (N_11967,N_11681,N_11650);
nand U11968 (N_11968,N_11626,N_11485);
and U11969 (N_11969,N_11520,N_11600);
xor U11970 (N_11970,N_11626,N_11634);
xor U11971 (N_11971,N_11484,N_11634);
and U11972 (N_11972,N_11427,N_11577);
nand U11973 (N_11973,N_11450,N_11507);
and U11974 (N_11974,N_11556,N_11500);
nand U11975 (N_11975,N_11622,N_11522);
nor U11976 (N_11976,N_11557,N_11619);
xnor U11977 (N_11977,N_11480,N_11513);
nand U11978 (N_11978,N_11638,N_11476);
xnor U11979 (N_11979,N_11602,N_11539);
xor U11980 (N_11980,N_11529,N_11461);
nand U11981 (N_11981,N_11643,N_11491);
nand U11982 (N_11982,N_11624,N_11512);
nor U11983 (N_11983,N_11498,N_11431);
xor U11984 (N_11984,N_11474,N_11532);
nand U11985 (N_11985,N_11617,N_11591);
and U11986 (N_11986,N_11654,N_11686);
and U11987 (N_11987,N_11589,N_11422);
nand U11988 (N_11988,N_11698,N_11450);
xor U11989 (N_11989,N_11600,N_11447);
or U11990 (N_11990,N_11580,N_11400);
xnor U11991 (N_11991,N_11445,N_11573);
nor U11992 (N_11992,N_11669,N_11604);
xor U11993 (N_11993,N_11484,N_11538);
nand U11994 (N_11994,N_11421,N_11455);
nor U11995 (N_11995,N_11622,N_11521);
or U11996 (N_11996,N_11452,N_11531);
or U11997 (N_11997,N_11607,N_11618);
and U11998 (N_11998,N_11562,N_11476);
xnor U11999 (N_11999,N_11558,N_11591);
nand U12000 (N_12000,N_11874,N_11866);
nor U12001 (N_12001,N_11875,N_11825);
or U12002 (N_12002,N_11770,N_11865);
xor U12003 (N_12003,N_11759,N_11858);
or U12004 (N_12004,N_11753,N_11976);
nor U12005 (N_12005,N_11939,N_11763);
nor U12006 (N_12006,N_11984,N_11715);
xor U12007 (N_12007,N_11931,N_11796);
or U12008 (N_12008,N_11852,N_11749);
or U12009 (N_12009,N_11822,N_11881);
nor U12010 (N_12010,N_11893,N_11913);
nor U12011 (N_12011,N_11803,N_11954);
nand U12012 (N_12012,N_11827,N_11779);
and U12013 (N_12013,N_11879,N_11994);
xor U12014 (N_12014,N_11834,N_11804);
xor U12015 (N_12015,N_11944,N_11772);
and U12016 (N_12016,N_11788,N_11819);
or U12017 (N_12017,N_11938,N_11723);
xor U12018 (N_12018,N_11747,N_11752);
or U12019 (N_12019,N_11761,N_11789);
nor U12020 (N_12020,N_11845,N_11967);
nor U12021 (N_12021,N_11800,N_11754);
and U12022 (N_12022,N_11989,N_11744);
xnor U12023 (N_12023,N_11959,N_11973);
or U12024 (N_12024,N_11783,N_11756);
or U12025 (N_12025,N_11871,N_11907);
nand U12026 (N_12026,N_11705,N_11771);
xor U12027 (N_12027,N_11781,N_11883);
nand U12028 (N_12028,N_11933,N_11988);
xnor U12029 (N_12029,N_11876,N_11785);
nor U12030 (N_12030,N_11709,N_11912);
nor U12031 (N_12031,N_11943,N_11860);
nor U12032 (N_12032,N_11814,N_11710);
nor U12033 (N_12033,N_11963,N_11859);
nand U12034 (N_12034,N_11702,N_11762);
or U12035 (N_12035,N_11884,N_11828);
nor U12036 (N_12036,N_11766,N_11846);
or U12037 (N_12037,N_11918,N_11950);
or U12038 (N_12038,N_11979,N_11835);
nor U12039 (N_12039,N_11873,N_11958);
xnor U12040 (N_12040,N_11991,N_11995);
and U12041 (N_12041,N_11768,N_11798);
nand U12042 (N_12042,N_11707,N_11997);
nand U12043 (N_12043,N_11864,N_11818);
nor U12044 (N_12044,N_11897,N_11712);
nand U12045 (N_12045,N_11731,N_11729);
or U12046 (N_12046,N_11996,N_11849);
nand U12047 (N_12047,N_11955,N_11888);
nand U12048 (N_12048,N_11802,N_11816);
and U12049 (N_12049,N_11823,N_11745);
or U12050 (N_12050,N_11947,N_11894);
nand U12051 (N_12051,N_11930,N_11901);
xnor U12052 (N_12052,N_11850,N_11760);
nand U12053 (N_12053,N_11978,N_11826);
xor U12054 (N_12054,N_11728,N_11869);
xor U12055 (N_12055,N_11778,N_11953);
and U12056 (N_12056,N_11807,N_11808);
xor U12057 (N_12057,N_11957,N_11703);
nand U12058 (N_12058,N_11986,N_11851);
xor U12059 (N_12059,N_11801,N_11946);
nor U12060 (N_12060,N_11926,N_11908);
xor U12061 (N_12061,N_11794,N_11777);
xnor U12062 (N_12062,N_11972,N_11708);
nand U12063 (N_12063,N_11843,N_11964);
and U12064 (N_12064,N_11880,N_11738);
xor U12065 (N_12065,N_11889,N_11962);
nor U12066 (N_12066,N_11837,N_11793);
nand U12067 (N_12067,N_11841,N_11840);
xor U12068 (N_12068,N_11810,N_11700);
nand U12069 (N_12069,N_11868,N_11861);
and U12070 (N_12070,N_11730,N_11820);
nand U12071 (N_12071,N_11790,N_11746);
or U12072 (N_12072,N_11848,N_11891);
nand U12073 (N_12073,N_11706,N_11951);
or U12074 (N_12074,N_11993,N_11878);
nand U12075 (N_12075,N_11758,N_11791);
xnor U12076 (N_12076,N_11928,N_11863);
nand U12077 (N_12077,N_11838,N_11857);
nor U12078 (N_12078,N_11960,N_11795);
and U12079 (N_12079,N_11985,N_11755);
xor U12080 (N_12080,N_11727,N_11915);
and U12081 (N_12081,N_11992,N_11739);
and U12082 (N_12082,N_11922,N_11799);
nor U12083 (N_12083,N_11911,N_11870);
xor U12084 (N_12084,N_11942,N_11900);
nand U12085 (N_12085,N_11975,N_11780);
or U12086 (N_12086,N_11971,N_11899);
nor U12087 (N_12087,N_11896,N_11824);
or U12088 (N_12088,N_11833,N_11853);
nand U12089 (N_12089,N_11941,N_11898);
xor U12090 (N_12090,N_11904,N_11867);
or U12091 (N_12091,N_11914,N_11935);
xor U12092 (N_12092,N_11885,N_11719);
xor U12093 (N_12093,N_11905,N_11811);
or U12094 (N_12094,N_11732,N_11817);
or U12095 (N_12095,N_11736,N_11990);
xor U12096 (N_12096,N_11812,N_11773);
and U12097 (N_12097,N_11981,N_11740);
nor U12098 (N_12098,N_11977,N_11965);
nor U12099 (N_12099,N_11765,N_11815);
nand U12100 (N_12100,N_11895,N_11805);
or U12101 (N_12101,N_11813,N_11919);
nand U12102 (N_12102,N_11970,N_11775);
nand U12103 (N_12103,N_11784,N_11952);
or U12104 (N_12104,N_11733,N_11956);
nand U12105 (N_12105,N_11842,N_11927);
xnor U12106 (N_12106,N_11832,N_11713);
nor U12107 (N_12107,N_11792,N_11724);
and U12108 (N_12108,N_11701,N_11903);
nand U12109 (N_12109,N_11750,N_11821);
and U12110 (N_12110,N_11769,N_11855);
or U12111 (N_12111,N_11776,N_11725);
or U12112 (N_12112,N_11916,N_11717);
nand U12113 (N_12113,N_11945,N_11961);
and U12114 (N_12114,N_11921,N_11839);
nand U12115 (N_12115,N_11999,N_11925);
or U12116 (N_12116,N_11872,N_11704);
or U12117 (N_12117,N_11774,N_11968);
nor U12118 (N_12118,N_11787,N_11902);
and U12119 (N_12119,N_11716,N_11937);
nor U12120 (N_12120,N_11836,N_11909);
nand U12121 (N_12121,N_11726,N_11906);
or U12122 (N_12122,N_11887,N_11735);
or U12123 (N_12123,N_11974,N_11711);
nor U12124 (N_12124,N_11757,N_11934);
xnor U12125 (N_12125,N_11969,N_11714);
or U12126 (N_12126,N_11782,N_11982);
xor U12127 (N_12127,N_11910,N_11809);
nand U12128 (N_12128,N_11847,N_11932);
nor U12129 (N_12129,N_11923,N_11936);
and U12130 (N_12130,N_11854,N_11720);
xnor U12131 (N_12131,N_11830,N_11829);
xor U12132 (N_12132,N_11718,N_11737);
nor U12133 (N_12133,N_11856,N_11949);
nor U12134 (N_12134,N_11844,N_11831);
and U12135 (N_12135,N_11966,N_11983);
nand U12136 (N_12136,N_11741,N_11748);
nor U12137 (N_12137,N_11767,N_11877);
nand U12138 (N_12138,N_11797,N_11722);
xor U12139 (N_12139,N_11998,N_11862);
nand U12140 (N_12140,N_11890,N_11948);
xor U12141 (N_12141,N_11743,N_11940);
nor U12142 (N_12142,N_11917,N_11929);
nor U12143 (N_12143,N_11742,N_11751);
xor U12144 (N_12144,N_11786,N_11806);
xor U12145 (N_12145,N_11892,N_11886);
xnor U12146 (N_12146,N_11987,N_11980);
and U12147 (N_12147,N_11764,N_11721);
or U12148 (N_12148,N_11924,N_11920);
or U12149 (N_12149,N_11882,N_11734);
or U12150 (N_12150,N_11936,N_11834);
nand U12151 (N_12151,N_11725,N_11988);
or U12152 (N_12152,N_11949,N_11773);
xnor U12153 (N_12153,N_11996,N_11919);
nor U12154 (N_12154,N_11790,N_11957);
nand U12155 (N_12155,N_11788,N_11878);
xnor U12156 (N_12156,N_11992,N_11858);
nor U12157 (N_12157,N_11758,N_11909);
and U12158 (N_12158,N_11724,N_11700);
nor U12159 (N_12159,N_11749,N_11899);
xor U12160 (N_12160,N_11782,N_11730);
or U12161 (N_12161,N_11865,N_11726);
or U12162 (N_12162,N_11864,N_11743);
nor U12163 (N_12163,N_11937,N_11830);
nor U12164 (N_12164,N_11762,N_11995);
and U12165 (N_12165,N_11748,N_11925);
xnor U12166 (N_12166,N_11802,N_11922);
nor U12167 (N_12167,N_11877,N_11967);
nand U12168 (N_12168,N_11813,N_11911);
nor U12169 (N_12169,N_11939,N_11821);
xnor U12170 (N_12170,N_11802,N_11838);
nand U12171 (N_12171,N_11989,N_11786);
nand U12172 (N_12172,N_11734,N_11843);
nand U12173 (N_12173,N_11861,N_11968);
and U12174 (N_12174,N_11851,N_11886);
xnor U12175 (N_12175,N_11774,N_11770);
nand U12176 (N_12176,N_11905,N_11763);
and U12177 (N_12177,N_11861,N_11920);
or U12178 (N_12178,N_11790,N_11767);
nor U12179 (N_12179,N_11951,N_11920);
xnor U12180 (N_12180,N_11747,N_11900);
nor U12181 (N_12181,N_11758,N_11722);
or U12182 (N_12182,N_11792,N_11848);
nor U12183 (N_12183,N_11882,N_11999);
nor U12184 (N_12184,N_11768,N_11803);
and U12185 (N_12185,N_11997,N_11778);
nor U12186 (N_12186,N_11995,N_11888);
or U12187 (N_12187,N_11768,N_11714);
and U12188 (N_12188,N_11920,N_11943);
and U12189 (N_12189,N_11763,N_11708);
xnor U12190 (N_12190,N_11714,N_11754);
and U12191 (N_12191,N_11998,N_11900);
xor U12192 (N_12192,N_11746,N_11848);
and U12193 (N_12193,N_11703,N_11971);
nand U12194 (N_12194,N_11700,N_11794);
nor U12195 (N_12195,N_11712,N_11700);
or U12196 (N_12196,N_11756,N_11849);
nand U12197 (N_12197,N_11700,N_11980);
nand U12198 (N_12198,N_11881,N_11762);
nand U12199 (N_12199,N_11764,N_11843);
or U12200 (N_12200,N_11782,N_11766);
and U12201 (N_12201,N_11983,N_11755);
or U12202 (N_12202,N_11813,N_11843);
or U12203 (N_12203,N_11771,N_11780);
nand U12204 (N_12204,N_11764,N_11794);
or U12205 (N_12205,N_11814,N_11733);
xnor U12206 (N_12206,N_11762,N_11965);
xnor U12207 (N_12207,N_11945,N_11842);
or U12208 (N_12208,N_11778,N_11834);
xor U12209 (N_12209,N_11775,N_11717);
nand U12210 (N_12210,N_11967,N_11890);
nor U12211 (N_12211,N_11770,N_11953);
nand U12212 (N_12212,N_11935,N_11740);
nor U12213 (N_12213,N_11869,N_11897);
xnor U12214 (N_12214,N_11801,N_11765);
and U12215 (N_12215,N_11704,N_11874);
nor U12216 (N_12216,N_11716,N_11802);
xnor U12217 (N_12217,N_11970,N_11700);
nand U12218 (N_12218,N_11786,N_11769);
or U12219 (N_12219,N_11829,N_11887);
and U12220 (N_12220,N_11909,N_11926);
and U12221 (N_12221,N_11911,N_11874);
and U12222 (N_12222,N_11755,N_11767);
nand U12223 (N_12223,N_11897,N_11786);
and U12224 (N_12224,N_11998,N_11831);
and U12225 (N_12225,N_11765,N_11846);
nor U12226 (N_12226,N_11920,N_11789);
or U12227 (N_12227,N_11987,N_11924);
or U12228 (N_12228,N_11855,N_11725);
nor U12229 (N_12229,N_11760,N_11837);
or U12230 (N_12230,N_11718,N_11814);
nand U12231 (N_12231,N_11817,N_11830);
nand U12232 (N_12232,N_11883,N_11791);
or U12233 (N_12233,N_11965,N_11901);
nor U12234 (N_12234,N_11896,N_11786);
nand U12235 (N_12235,N_11851,N_11803);
or U12236 (N_12236,N_11729,N_11946);
nor U12237 (N_12237,N_11839,N_11880);
or U12238 (N_12238,N_11947,N_11799);
and U12239 (N_12239,N_11810,N_11974);
nand U12240 (N_12240,N_11703,N_11894);
nand U12241 (N_12241,N_11727,N_11996);
nor U12242 (N_12242,N_11886,N_11805);
and U12243 (N_12243,N_11967,N_11743);
nor U12244 (N_12244,N_11715,N_11982);
xnor U12245 (N_12245,N_11931,N_11926);
or U12246 (N_12246,N_11843,N_11975);
nor U12247 (N_12247,N_11944,N_11806);
xor U12248 (N_12248,N_11982,N_11857);
nor U12249 (N_12249,N_11990,N_11864);
nor U12250 (N_12250,N_11918,N_11979);
or U12251 (N_12251,N_11766,N_11986);
nor U12252 (N_12252,N_11820,N_11920);
and U12253 (N_12253,N_11954,N_11949);
nor U12254 (N_12254,N_11984,N_11713);
nand U12255 (N_12255,N_11986,N_11713);
xnor U12256 (N_12256,N_11701,N_11808);
and U12257 (N_12257,N_11972,N_11827);
and U12258 (N_12258,N_11912,N_11815);
xor U12259 (N_12259,N_11933,N_11756);
nand U12260 (N_12260,N_11947,N_11850);
and U12261 (N_12261,N_11892,N_11950);
or U12262 (N_12262,N_11774,N_11761);
nor U12263 (N_12263,N_11859,N_11982);
and U12264 (N_12264,N_11721,N_11973);
and U12265 (N_12265,N_11941,N_11918);
xor U12266 (N_12266,N_11703,N_11819);
nand U12267 (N_12267,N_11884,N_11763);
or U12268 (N_12268,N_11930,N_11772);
and U12269 (N_12269,N_11920,N_11891);
or U12270 (N_12270,N_11779,N_11867);
nor U12271 (N_12271,N_11880,N_11730);
and U12272 (N_12272,N_11827,N_11856);
and U12273 (N_12273,N_11961,N_11898);
nand U12274 (N_12274,N_11781,N_11857);
and U12275 (N_12275,N_11859,N_11774);
xnor U12276 (N_12276,N_11742,N_11903);
and U12277 (N_12277,N_11811,N_11921);
and U12278 (N_12278,N_11925,N_11841);
nand U12279 (N_12279,N_11933,N_11845);
and U12280 (N_12280,N_11983,N_11778);
nor U12281 (N_12281,N_11752,N_11813);
xor U12282 (N_12282,N_11752,N_11975);
and U12283 (N_12283,N_11793,N_11700);
nand U12284 (N_12284,N_11815,N_11741);
and U12285 (N_12285,N_11853,N_11810);
nand U12286 (N_12286,N_11743,N_11981);
and U12287 (N_12287,N_11927,N_11875);
xnor U12288 (N_12288,N_11960,N_11794);
xnor U12289 (N_12289,N_11797,N_11771);
nor U12290 (N_12290,N_11893,N_11826);
nand U12291 (N_12291,N_11930,N_11974);
or U12292 (N_12292,N_11846,N_11901);
xnor U12293 (N_12293,N_11813,N_11875);
or U12294 (N_12294,N_11972,N_11975);
and U12295 (N_12295,N_11917,N_11840);
xnor U12296 (N_12296,N_11764,N_11781);
or U12297 (N_12297,N_11718,N_11828);
and U12298 (N_12298,N_11949,N_11751);
nand U12299 (N_12299,N_11729,N_11931);
nand U12300 (N_12300,N_12107,N_12097);
nand U12301 (N_12301,N_12200,N_12241);
nand U12302 (N_12302,N_12048,N_12099);
nand U12303 (N_12303,N_12135,N_12050);
xnor U12304 (N_12304,N_12251,N_12081);
and U12305 (N_12305,N_12177,N_12110);
or U12306 (N_12306,N_12210,N_12216);
nor U12307 (N_12307,N_12129,N_12109);
nand U12308 (N_12308,N_12131,N_12270);
and U12309 (N_12309,N_12127,N_12188);
and U12310 (N_12310,N_12062,N_12125);
or U12311 (N_12311,N_12041,N_12174);
nor U12312 (N_12312,N_12195,N_12155);
xor U12313 (N_12313,N_12024,N_12149);
xor U12314 (N_12314,N_12299,N_12017);
nand U12315 (N_12315,N_12186,N_12122);
and U12316 (N_12316,N_12157,N_12243);
or U12317 (N_12317,N_12255,N_12208);
xnor U12318 (N_12318,N_12291,N_12185);
or U12319 (N_12319,N_12284,N_12094);
nand U12320 (N_12320,N_12137,N_12212);
nand U12321 (N_12321,N_12281,N_12068);
xor U12322 (N_12322,N_12134,N_12228);
nand U12323 (N_12323,N_12108,N_12112);
or U12324 (N_12324,N_12114,N_12295);
nand U12325 (N_12325,N_12238,N_12260);
nand U12326 (N_12326,N_12269,N_12267);
and U12327 (N_12327,N_12064,N_12049);
nand U12328 (N_12328,N_12076,N_12214);
and U12329 (N_12329,N_12098,N_12219);
nand U12330 (N_12330,N_12139,N_12215);
nor U12331 (N_12331,N_12169,N_12126);
nor U12332 (N_12332,N_12207,N_12007);
or U12333 (N_12333,N_12170,N_12123);
xnor U12334 (N_12334,N_12147,N_12204);
and U12335 (N_12335,N_12136,N_12248);
nand U12336 (N_12336,N_12013,N_12089);
or U12337 (N_12337,N_12266,N_12156);
xor U12338 (N_12338,N_12060,N_12293);
or U12339 (N_12339,N_12067,N_12254);
or U12340 (N_12340,N_12145,N_12229);
nand U12341 (N_12341,N_12282,N_12113);
nor U12342 (N_12342,N_12033,N_12172);
and U12343 (N_12343,N_12225,N_12040);
or U12344 (N_12344,N_12008,N_12275);
nand U12345 (N_12345,N_12085,N_12015);
and U12346 (N_12346,N_12004,N_12231);
and U12347 (N_12347,N_12002,N_12163);
xnor U12348 (N_12348,N_12096,N_12093);
nor U12349 (N_12349,N_12223,N_12078);
nand U12350 (N_12350,N_12003,N_12262);
nand U12351 (N_12351,N_12237,N_12006);
nand U12352 (N_12352,N_12274,N_12146);
xor U12353 (N_12353,N_12055,N_12294);
nand U12354 (N_12354,N_12246,N_12259);
or U12355 (N_12355,N_12077,N_12190);
or U12356 (N_12356,N_12173,N_12034);
nand U12357 (N_12357,N_12198,N_12245);
or U12358 (N_12358,N_12205,N_12028);
and U12359 (N_12359,N_12199,N_12148);
and U12360 (N_12360,N_12118,N_12117);
or U12361 (N_12361,N_12133,N_12232);
nor U12362 (N_12362,N_12023,N_12263);
nor U12363 (N_12363,N_12106,N_12080);
xor U12364 (N_12364,N_12268,N_12277);
nand U12365 (N_12365,N_12273,N_12193);
xor U12366 (N_12366,N_12289,N_12092);
or U12367 (N_12367,N_12104,N_12162);
and U12368 (N_12368,N_12100,N_12069);
nor U12369 (N_12369,N_12025,N_12022);
nand U12370 (N_12370,N_12253,N_12265);
xor U12371 (N_12371,N_12138,N_12236);
and U12372 (N_12372,N_12063,N_12059);
nor U12373 (N_12373,N_12036,N_12020);
or U12374 (N_12374,N_12038,N_12235);
nand U12375 (N_12375,N_12019,N_12032);
and U12376 (N_12376,N_12280,N_12016);
nor U12377 (N_12377,N_12012,N_12075);
nor U12378 (N_12378,N_12086,N_12161);
nand U12379 (N_12379,N_12070,N_12224);
nor U12380 (N_12380,N_12196,N_12121);
and U12381 (N_12381,N_12296,N_12090);
and U12382 (N_12382,N_12184,N_12227);
xnor U12383 (N_12383,N_12128,N_12014);
xnor U12384 (N_12384,N_12189,N_12230);
and U12385 (N_12385,N_12244,N_12256);
and U12386 (N_12386,N_12175,N_12091);
xor U12387 (N_12387,N_12249,N_12192);
nor U12388 (N_12388,N_12166,N_12058);
nor U12389 (N_12389,N_12165,N_12119);
and U12390 (N_12390,N_12039,N_12018);
nor U12391 (N_12391,N_12221,N_12087);
xor U12392 (N_12392,N_12187,N_12031);
nor U12393 (N_12393,N_12071,N_12181);
xnor U12394 (N_12394,N_12285,N_12000);
and U12395 (N_12395,N_12171,N_12105);
xor U12396 (N_12396,N_12276,N_12292);
xor U12397 (N_12397,N_12178,N_12074);
xor U12398 (N_12398,N_12141,N_12233);
xnor U12399 (N_12399,N_12182,N_12180);
nor U12400 (N_12400,N_12220,N_12240);
or U12401 (N_12401,N_12083,N_12103);
and U12402 (N_12402,N_12079,N_12047);
xor U12403 (N_12403,N_12234,N_12154);
and U12404 (N_12404,N_12026,N_12001);
xor U12405 (N_12405,N_12043,N_12124);
or U12406 (N_12406,N_12046,N_12211);
and U12407 (N_12407,N_12286,N_12052);
nor U12408 (N_12408,N_12258,N_12283);
or U12409 (N_12409,N_12035,N_12250);
and U12410 (N_12410,N_12222,N_12030);
or U12411 (N_12411,N_12088,N_12115);
nor U12412 (N_12412,N_12159,N_12213);
or U12413 (N_12413,N_12045,N_12066);
and U12414 (N_12414,N_12209,N_12179);
and U12415 (N_12415,N_12130,N_12143);
and U12416 (N_12416,N_12167,N_12053);
nand U12417 (N_12417,N_12203,N_12279);
or U12418 (N_12418,N_12239,N_12278);
xor U12419 (N_12419,N_12218,N_12027);
xor U12420 (N_12420,N_12061,N_12264);
nand U12421 (N_12421,N_12054,N_12057);
xnor U12422 (N_12422,N_12176,N_12072);
and U12423 (N_12423,N_12297,N_12164);
and U12424 (N_12424,N_12288,N_12152);
nor U12425 (N_12425,N_12298,N_12183);
nor U12426 (N_12426,N_12120,N_12010);
or U12427 (N_12427,N_12247,N_12132);
nand U12428 (N_12428,N_12158,N_12011);
and U12429 (N_12429,N_12021,N_12194);
xor U12430 (N_12430,N_12242,N_12271);
xor U12431 (N_12431,N_12287,N_12116);
or U12432 (N_12432,N_12153,N_12290);
and U12433 (N_12433,N_12051,N_12029);
or U12434 (N_12434,N_12140,N_12217);
nor U12435 (N_12435,N_12191,N_12073);
nand U12436 (N_12436,N_12197,N_12252);
nor U12437 (N_12437,N_12257,N_12082);
nand U12438 (N_12438,N_12044,N_12150);
nor U12439 (N_12439,N_12084,N_12037);
nand U12440 (N_12440,N_12201,N_12009);
or U12441 (N_12441,N_12151,N_12168);
and U12442 (N_12442,N_12261,N_12065);
nor U12443 (N_12443,N_12111,N_12226);
xor U12444 (N_12444,N_12042,N_12056);
nor U12445 (N_12445,N_12144,N_12102);
nor U12446 (N_12446,N_12272,N_12101);
or U12447 (N_12447,N_12202,N_12095);
nor U12448 (N_12448,N_12206,N_12005);
and U12449 (N_12449,N_12142,N_12160);
nand U12450 (N_12450,N_12266,N_12173);
nand U12451 (N_12451,N_12227,N_12044);
or U12452 (N_12452,N_12229,N_12063);
xor U12453 (N_12453,N_12018,N_12074);
nand U12454 (N_12454,N_12184,N_12231);
xor U12455 (N_12455,N_12205,N_12039);
or U12456 (N_12456,N_12063,N_12165);
and U12457 (N_12457,N_12091,N_12212);
nand U12458 (N_12458,N_12108,N_12268);
and U12459 (N_12459,N_12151,N_12217);
nor U12460 (N_12460,N_12150,N_12259);
xor U12461 (N_12461,N_12197,N_12032);
or U12462 (N_12462,N_12292,N_12019);
xor U12463 (N_12463,N_12088,N_12141);
nand U12464 (N_12464,N_12282,N_12126);
nand U12465 (N_12465,N_12251,N_12150);
nor U12466 (N_12466,N_12033,N_12023);
and U12467 (N_12467,N_12034,N_12258);
nor U12468 (N_12468,N_12171,N_12109);
nor U12469 (N_12469,N_12206,N_12066);
nor U12470 (N_12470,N_12210,N_12123);
nand U12471 (N_12471,N_12064,N_12041);
nand U12472 (N_12472,N_12017,N_12265);
xnor U12473 (N_12473,N_12011,N_12278);
or U12474 (N_12474,N_12232,N_12275);
nand U12475 (N_12475,N_12089,N_12064);
nor U12476 (N_12476,N_12264,N_12199);
nor U12477 (N_12477,N_12062,N_12046);
nand U12478 (N_12478,N_12222,N_12054);
xnor U12479 (N_12479,N_12221,N_12199);
nand U12480 (N_12480,N_12249,N_12271);
nor U12481 (N_12481,N_12016,N_12243);
xor U12482 (N_12482,N_12063,N_12099);
and U12483 (N_12483,N_12041,N_12141);
nand U12484 (N_12484,N_12254,N_12008);
or U12485 (N_12485,N_12010,N_12000);
or U12486 (N_12486,N_12065,N_12092);
or U12487 (N_12487,N_12111,N_12199);
xor U12488 (N_12488,N_12156,N_12007);
xor U12489 (N_12489,N_12167,N_12150);
nor U12490 (N_12490,N_12296,N_12217);
nor U12491 (N_12491,N_12260,N_12154);
or U12492 (N_12492,N_12239,N_12270);
nor U12493 (N_12493,N_12175,N_12176);
nor U12494 (N_12494,N_12021,N_12023);
and U12495 (N_12495,N_12166,N_12282);
and U12496 (N_12496,N_12144,N_12175);
nor U12497 (N_12497,N_12117,N_12045);
and U12498 (N_12498,N_12195,N_12053);
or U12499 (N_12499,N_12079,N_12011);
nand U12500 (N_12500,N_12201,N_12224);
nor U12501 (N_12501,N_12292,N_12125);
or U12502 (N_12502,N_12128,N_12215);
and U12503 (N_12503,N_12035,N_12096);
nor U12504 (N_12504,N_12188,N_12156);
or U12505 (N_12505,N_12071,N_12014);
nor U12506 (N_12506,N_12247,N_12030);
xnor U12507 (N_12507,N_12276,N_12093);
nand U12508 (N_12508,N_12045,N_12091);
nor U12509 (N_12509,N_12186,N_12130);
or U12510 (N_12510,N_12175,N_12021);
and U12511 (N_12511,N_12191,N_12078);
nor U12512 (N_12512,N_12113,N_12170);
or U12513 (N_12513,N_12090,N_12147);
nor U12514 (N_12514,N_12148,N_12035);
nand U12515 (N_12515,N_12144,N_12046);
nand U12516 (N_12516,N_12288,N_12276);
and U12517 (N_12517,N_12087,N_12104);
nand U12518 (N_12518,N_12083,N_12235);
or U12519 (N_12519,N_12003,N_12102);
nand U12520 (N_12520,N_12272,N_12132);
xnor U12521 (N_12521,N_12298,N_12291);
xor U12522 (N_12522,N_12178,N_12221);
or U12523 (N_12523,N_12145,N_12026);
xnor U12524 (N_12524,N_12083,N_12169);
xor U12525 (N_12525,N_12266,N_12032);
nand U12526 (N_12526,N_12121,N_12001);
nand U12527 (N_12527,N_12084,N_12038);
and U12528 (N_12528,N_12105,N_12002);
or U12529 (N_12529,N_12198,N_12224);
and U12530 (N_12530,N_12034,N_12003);
nor U12531 (N_12531,N_12214,N_12071);
nor U12532 (N_12532,N_12141,N_12210);
nor U12533 (N_12533,N_12072,N_12226);
nand U12534 (N_12534,N_12150,N_12152);
nand U12535 (N_12535,N_12211,N_12239);
nand U12536 (N_12536,N_12107,N_12238);
or U12537 (N_12537,N_12225,N_12153);
nand U12538 (N_12538,N_12060,N_12034);
nor U12539 (N_12539,N_12271,N_12244);
nor U12540 (N_12540,N_12244,N_12023);
nand U12541 (N_12541,N_12008,N_12106);
nor U12542 (N_12542,N_12267,N_12123);
xor U12543 (N_12543,N_12011,N_12268);
xnor U12544 (N_12544,N_12219,N_12000);
nand U12545 (N_12545,N_12199,N_12138);
xnor U12546 (N_12546,N_12041,N_12150);
nand U12547 (N_12547,N_12093,N_12293);
xor U12548 (N_12548,N_12039,N_12050);
nand U12549 (N_12549,N_12064,N_12042);
and U12550 (N_12550,N_12105,N_12059);
xnor U12551 (N_12551,N_12039,N_12000);
xnor U12552 (N_12552,N_12084,N_12213);
nand U12553 (N_12553,N_12223,N_12271);
and U12554 (N_12554,N_12127,N_12033);
and U12555 (N_12555,N_12059,N_12172);
or U12556 (N_12556,N_12192,N_12160);
and U12557 (N_12557,N_12129,N_12136);
and U12558 (N_12558,N_12139,N_12164);
nor U12559 (N_12559,N_12278,N_12055);
or U12560 (N_12560,N_12120,N_12299);
xor U12561 (N_12561,N_12049,N_12151);
xnor U12562 (N_12562,N_12205,N_12155);
nor U12563 (N_12563,N_12075,N_12041);
xnor U12564 (N_12564,N_12256,N_12150);
and U12565 (N_12565,N_12130,N_12249);
nand U12566 (N_12566,N_12141,N_12227);
or U12567 (N_12567,N_12221,N_12226);
and U12568 (N_12568,N_12270,N_12205);
xnor U12569 (N_12569,N_12265,N_12234);
nand U12570 (N_12570,N_12295,N_12020);
xor U12571 (N_12571,N_12053,N_12198);
and U12572 (N_12572,N_12247,N_12245);
and U12573 (N_12573,N_12106,N_12181);
and U12574 (N_12574,N_12045,N_12071);
xor U12575 (N_12575,N_12235,N_12049);
xor U12576 (N_12576,N_12258,N_12196);
nor U12577 (N_12577,N_12009,N_12109);
nand U12578 (N_12578,N_12123,N_12124);
nor U12579 (N_12579,N_12295,N_12002);
and U12580 (N_12580,N_12156,N_12213);
nand U12581 (N_12581,N_12068,N_12160);
or U12582 (N_12582,N_12218,N_12166);
nand U12583 (N_12583,N_12130,N_12151);
nor U12584 (N_12584,N_12082,N_12067);
or U12585 (N_12585,N_12174,N_12071);
xnor U12586 (N_12586,N_12207,N_12081);
and U12587 (N_12587,N_12148,N_12219);
nand U12588 (N_12588,N_12139,N_12114);
or U12589 (N_12589,N_12082,N_12207);
or U12590 (N_12590,N_12251,N_12230);
nand U12591 (N_12591,N_12178,N_12131);
xor U12592 (N_12592,N_12237,N_12078);
nand U12593 (N_12593,N_12290,N_12259);
xnor U12594 (N_12594,N_12072,N_12115);
and U12595 (N_12595,N_12225,N_12239);
or U12596 (N_12596,N_12002,N_12035);
xnor U12597 (N_12597,N_12094,N_12154);
and U12598 (N_12598,N_12128,N_12203);
xor U12599 (N_12599,N_12165,N_12190);
nor U12600 (N_12600,N_12533,N_12365);
nand U12601 (N_12601,N_12395,N_12408);
or U12602 (N_12602,N_12593,N_12428);
or U12603 (N_12603,N_12349,N_12421);
nor U12604 (N_12604,N_12401,N_12520);
and U12605 (N_12605,N_12560,N_12339);
or U12606 (N_12606,N_12352,N_12381);
and U12607 (N_12607,N_12334,N_12583);
nor U12608 (N_12608,N_12417,N_12411);
nor U12609 (N_12609,N_12493,N_12391);
or U12610 (N_12610,N_12506,N_12535);
nor U12611 (N_12611,N_12576,N_12549);
and U12612 (N_12612,N_12574,N_12521);
or U12613 (N_12613,N_12434,N_12505);
and U12614 (N_12614,N_12548,N_12579);
nor U12615 (N_12615,N_12324,N_12309);
and U12616 (N_12616,N_12449,N_12597);
or U12617 (N_12617,N_12376,N_12363);
nor U12618 (N_12618,N_12366,N_12302);
and U12619 (N_12619,N_12586,N_12384);
or U12620 (N_12620,N_12319,N_12488);
nor U12621 (N_12621,N_12592,N_12343);
or U12622 (N_12622,N_12466,N_12478);
nand U12623 (N_12623,N_12407,N_12513);
xnor U12624 (N_12624,N_12594,N_12370);
nor U12625 (N_12625,N_12353,N_12371);
xnor U12626 (N_12626,N_12397,N_12356);
or U12627 (N_12627,N_12410,N_12476);
nand U12628 (N_12628,N_12322,N_12373);
xnor U12629 (N_12629,N_12498,N_12490);
nor U12630 (N_12630,N_12458,N_12350);
or U12631 (N_12631,N_12547,N_12569);
nor U12632 (N_12632,N_12345,N_12435);
and U12633 (N_12633,N_12452,N_12389);
nand U12634 (N_12634,N_12387,N_12461);
and U12635 (N_12635,N_12554,N_12374);
and U12636 (N_12636,N_12497,N_12336);
nor U12637 (N_12637,N_12450,N_12300);
or U12638 (N_12638,N_12555,N_12426);
nand U12639 (N_12639,N_12358,N_12534);
or U12640 (N_12640,N_12479,N_12396);
and U12641 (N_12641,N_12443,N_12315);
nor U12642 (N_12642,N_12462,N_12453);
and U12643 (N_12643,N_12551,N_12532);
and U12644 (N_12644,N_12444,N_12424);
and U12645 (N_12645,N_12541,N_12527);
and U12646 (N_12646,N_12509,N_12474);
or U12647 (N_12647,N_12346,N_12321);
or U12648 (N_12648,N_12472,N_12344);
and U12649 (N_12649,N_12330,N_12415);
nor U12650 (N_12650,N_12305,N_12437);
nand U12651 (N_12651,N_12456,N_12399);
and U12652 (N_12652,N_12433,N_12316);
xor U12653 (N_12653,N_12325,N_12465);
nor U12654 (N_12654,N_12328,N_12416);
or U12655 (N_12655,N_12578,N_12524);
xor U12656 (N_12656,N_12369,N_12332);
nor U12657 (N_12657,N_12361,N_12572);
xor U12658 (N_12658,N_12483,N_12459);
and U12659 (N_12659,N_12587,N_12420);
and U12660 (N_12660,N_12357,N_12313);
nand U12661 (N_12661,N_12368,N_12582);
and U12662 (N_12662,N_12556,N_12386);
xnor U12663 (N_12663,N_12499,N_12496);
nand U12664 (N_12664,N_12454,N_12446);
nand U12665 (N_12665,N_12372,N_12335);
and U12666 (N_12666,N_12311,N_12503);
nand U12667 (N_12667,N_12378,N_12337);
or U12668 (N_12668,N_12385,N_12501);
and U12669 (N_12669,N_12557,N_12575);
nor U12670 (N_12670,N_12425,N_12568);
nor U12671 (N_12671,N_12562,N_12355);
or U12672 (N_12672,N_12559,N_12563);
nor U12673 (N_12673,N_12413,N_12537);
or U12674 (N_12674,N_12473,N_12545);
nand U12675 (N_12675,N_12566,N_12451);
or U12676 (N_12676,N_12514,N_12412);
xor U12677 (N_12677,N_12348,N_12494);
xor U12678 (N_12678,N_12418,N_12308);
nor U12679 (N_12679,N_12409,N_12573);
or U12680 (N_12680,N_12404,N_12414);
and U12681 (N_12681,N_12406,N_12477);
nand U12682 (N_12682,N_12317,N_12570);
or U12683 (N_12683,N_12400,N_12340);
nand U12684 (N_12684,N_12436,N_12571);
or U12685 (N_12685,N_12375,N_12538);
xor U12686 (N_12686,N_12312,N_12471);
and U12687 (N_12687,N_12581,N_12360);
xor U12688 (N_12688,N_12565,N_12564);
xor U12689 (N_12689,N_12338,N_12398);
or U12690 (N_12690,N_12543,N_12427);
or U12691 (N_12691,N_12445,N_12530);
nor U12692 (N_12692,N_12591,N_12392);
and U12693 (N_12693,N_12383,N_12439);
nand U12694 (N_12694,N_12333,N_12492);
and U12695 (N_12695,N_12469,N_12516);
or U12696 (N_12696,N_12528,N_12359);
nand U12697 (N_12697,N_12377,N_12326);
nor U12698 (N_12698,N_12596,N_12429);
nand U12699 (N_12699,N_12354,N_12301);
nor U12700 (N_12700,N_12480,N_12405);
and U12701 (N_12701,N_12431,N_12525);
nor U12702 (N_12702,N_12307,N_12342);
or U12703 (N_12703,N_12553,N_12577);
or U12704 (N_12704,N_12588,N_12544);
xnor U12705 (N_12705,N_12519,N_12448);
or U12706 (N_12706,N_12550,N_12475);
nand U12707 (N_12707,N_12511,N_12491);
nand U12708 (N_12708,N_12382,N_12585);
nor U12709 (N_12709,N_12529,N_12487);
and U12710 (N_12710,N_12419,N_12526);
and U12711 (N_12711,N_12507,N_12589);
and U12712 (N_12712,N_12517,N_12460);
nor U12713 (N_12713,N_12430,N_12455);
or U12714 (N_12714,N_12536,N_12489);
nand U12715 (N_12715,N_12341,N_12590);
nand U12716 (N_12716,N_12485,N_12486);
nand U12717 (N_12717,N_12510,N_12599);
nand U12718 (N_12718,N_12432,N_12364);
and U12719 (N_12719,N_12422,N_12310);
nor U12720 (N_12720,N_12495,N_12523);
or U12721 (N_12721,N_12504,N_12380);
nor U12722 (N_12722,N_12467,N_12595);
nor U12723 (N_12723,N_12558,N_12463);
or U12724 (N_12724,N_12440,N_12567);
or U12725 (N_12725,N_12481,N_12484);
nand U12726 (N_12726,N_12584,N_12470);
nand U12727 (N_12727,N_12438,N_12393);
xor U12728 (N_12728,N_12329,N_12327);
xnor U12729 (N_12729,N_12508,N_12598);
and U12730 (N_12730,N_12515,N_12442);
or U12731 (N_12731,N_12522,N_12561);
or U12732 (N_12732,N_12546,N_12390);
and U12733 (N_12733,N_12464,N_12320);
nand U12734 (N_12734,N_12540,N_12552);
and U12735 (N_12735,N_12512,N_12500);
nand U12736 (N_12736,N_12468,N_12394);
or U12737 (N_12737,N_12347,N_12518);
nor U12738 (N_12738,N_12539,N_12306);
nor U12739 (N_12739,N_12351,N_12482);
and U12740 (N_12740,N_12362,N_12379);
and U12741 (N_12741,N_12367,N_12323);
or U12742 (N_12742,N_12423,N_12388);
nor U12743 (N_12743,N_12303,N_12580);
and U12744 (N_12744,N_12402,N_12502);
xor U12745 (N_12745,N_12331,N_12457);
xnor U12746 (N_12746,N_12447,N_12314);
nor U12747 (N_12747,N_12403,N_12531);
nor U12748 (N_12748,N_12318,N_12542);
nand U12749 (N_12749,N_12441,N_12304);
or U12750 (N_12750,N_12557,N_12579);
and U12751 (N_12751,N_12554,N_12444);
and U12752 (N_12752,N_12425,N_12446);
or U12753 (N_12753,N_12303,N_12574);
and U12754 (N_12754,N_12593,N_12390);
nand U12755 (N_12755,N_12398,N_12408);
nand U12756 (N_12756,N_12425,N_12380);
xnor U12757 (N_12757,N_12351,N_12436);
or U12758 (N_12758,N_12374,N_12457);
nor U12759 (N_12759,N_12586,N_12371);
and U12760 (N_12760,N_12499,N_12554);
nor U12761 (N_12761,N_12535,N_12410);
or U12762 (N_12762,N_12510,N_12344);
nor U12763 (N_12763,N_12537,N_12492);
nor U12764 (N_12764,N_12376,N_12359);
or U12765 (N_12765,N_12549,N_12512);
or U12766 (N_12766,N_12410,N_12524);
and U12767 (N_12767,N_12360,N_12317);
and U12768 (N_12768,N_12368,N_12327);
nand U12769 (N_12769,N_12591,N_12399);
nand U12770 (N_12770,N_12386,N_12307);
or U12771 (N_12771,N_12330,N_12486);
xor U12772 (N_12772,N_12544,N_12476);
or U12773 (N_12773,N_12427,N_12572);
nand U12774 (N_12774,N_12346,N_12316);
nand U12775 (N_12775,N_12365,N_12431);
or U12776 (N_12776,N_12530,N_12430);
or U12777 (N_12777,N_12310,N_12323);
nor U12778 (N_12778,N_12331,N_12477);
nand U12779 (N_12779,N_12426,N_12408);
and U12780 (N_12780,N_12438,N_12526);
and U12781 (N_12781,N_12422,N_12544);
and U12782 (N_12782,N_12428,N_12427);
and U12783 (N_12783,N_12458,N_12310);
xor U12784 (N_12784,N_12562,N_12373);
or U12785 (N_12785,N_12415,N_12500);
nor U12786 (N_12786,N_12460,N_12508);
and U12787 (N_12787,N_12535,N_12533);
nand U12788 (N_12788,N_12386,N_12495);
or U12789 (N_12789,N_12351,N_12583);
or U12790 (N_12790,N_12305,N_12416);
and U12791 (N_12791,N_12347,N_12455);
or U12792 (N_12792,N_12446,N_12404);
nand U12793 (N_12793,N_12426,N_12433);
or U12794 (N_12794,N_12542,N_12522);
nor U12795 (N_12795,N_12409,N_12442);
or U12796 (N_12796,N_12331,N_12323);
or U12797 (N_12797,N_12434,N_12551);
or U12798 (N_12798,N_12584,N_12414);
and U12799 (N_12799,N_12366,N_12495);
xnor U12800 (N_12800,N_12497,N_12512);
nand U12801 (N_12801,N_12437,N_12318);
nor U12802 (N_12802,N_12496,N_12489);
nand U12803 (N_12803,N_12533,N_12407);
nor U12804 (N_12804,N_12475,N_12305);
xnor U12805 (N_12805,N_12463,N_12565);
or U12806 (N_12806,N_12467,N_12459);
xor U12807 (N_12807,N_12434,N_12366);
nand U12808 (N_12808,N_12325,N_12395);
nand U12809 (N_12809,N_12593,N_12561);
xor U12810 (N_12810,N_12309,N_12592);
or U12811 (N_12811,N_12483,N_12321);
nor U12812 (N_12812,N_12320,N_12319);
nor U12813 (N_12813,N_12548,N_12363);
nor U12814 (N_12814,N_12333,N_12397);
or U12815 (N_12815,N_12363,N_12393);
and U12816 (N_12816,N_12555,N_12330);
nor U12817 (N_12817,N_12508,N_12530);
nand U12818 (N_12818,N_12487,N_12525);
xnor U12819 (N_12819,N_12310,N_12536);
and U12820 (N_12820,N_12478,N_12534);
or U12821 (N_12821,N_12556,N_12337);
xnor U12822 (N_12822,N_12406,N_12428);
or U12823 (N_12823,N_12548,N_12585);
nor U12824 (N_12824,N_12491,N_12538);
xnor U12825 (N_12825,N_12482,N_12405);
nand U12826 (N_12826,N_12396,N_12529);
and U12827 (N_12827,N_12486,N_12395);
nor U12828 (N_12828,N_12367,N_12495);
nand U12829 (N_12829,N_12382,N_12597);
xnor U12830 (N_12830,N_12459,N_12351);
or U12831 (N_12831,N_12579,N_12464);
nand U12832 (N_12832,N_12460,N_12347);
or U12833 (N_12833,N_12329,N_12406);
nor U12834 (N_12834,N_12509,N_12367);
xor U12835 (N_12835,N_12459,N_12540);
nor U12836 (N_12836,N_12552,N_12375);
nand U12837 (N_12837,N_12382,N_12303);
or U12838 (N_12838,N_12491,N_12534);
nor U12839 (N_12839,N_12331,N_12541);
or U12840 (N_12840,N_12492,N_12321);
and U12841 (N_12841,N_12590,N_12479);
nand U12842 (N_12842,N_12520,N_12451);
nand U12843 (N_12843,N_12530,N_12363);
xor U12844 (N_12844,N_12436,N_12300);
or U12845 (N_12845,N_12411,N_12340);
xor U12846 (N_12846,N_12520,N_12354);
nand U12847 (N_12847,N_12420,N_12578);
nand U12848 (N_12848,N_12585,N_12590);
xor U12849 (N_12849,N_12474,N_12442);
and U12850 (N_12850,N_12419,N_12570);
or U12851 (N_12851,N_12367,N_12328);
xnor U12852 (N_12852,N_12368,N_12580);
nor U12853 (N_12853,N_12464,N_12539);
nor U12854 (N_12854,N_12584,N_12517);
or U12855 (N_12855,N_12456,N_12335);
nand U12856 (N_12856,N_12452,N_12446);
or U12857 (N_12857,N_12477,N_12514);
xnor U12858 (N_12858,N_12450,N_12462);
nand U12859 (N_12859,N_12507,N_12325);
nor U12860 (N_12860,N_12513,N_12449);
nand U12861 (N_12861,N_12459,N_12578);
nor U12862 (N_12862,N_12463,N_12344);
nand U12863 (N_12863,N_12374,N_12429);
nor U12864 (N_12864,N_12581,N_12559);
and U12865 (N_12865,N_12391,N_12406);
nor U12866 (N_12866,N_12346,N_12498);
nor U12867 (N_12867,N_12366,N_12587);
or U12868 (N_12868,N_12545,N_12422);
xnor U12869 (N_12869,N_12515,N_12361);
nand U12870 (N_12870,N_12383,N_12548);
nand U12871 (N_12871,N_12447,N_12549);
nor U12872 (N_12872,N_12562,N_12512);
or U12873 (N_12873,N_12573,N_12443);
xor U12874 (N_12874,N_12531,N_12522);
xnor U12875 (N_12875,N_12379,N_12325);
and U12876 (N_12876,N_12596,N_12445);
nand U12877 (N_12877,N_12391,N_12497);
xor U12878 (N_12878,N_12378,N_12359);
or U12879 (N_12879,N_12338,N_12528);
nand U12880 (N_12880,N_12372,N_12394);
and U12881 (N_12881,N_12460,N_12337);
nor U12882 (N_12882,N_12388,N_12495);
nand U12883 (N_12883,N_12425,N_12352);
nand U12884 (N_12884,N_12493,N_12482);
nand U12885 (N_12885,N_12431,N_12583);
xor U12886 (N_12886,N_12422,N_12373);
and U12887 (N_12887,N_12488,N_12531);
nor U12888 (N_12888,N_12494,N_12367);
nor U12889 (N_12889,N_12455,N_12572);
nor U12890 (N_12890,N_12474,N_12328);
nand U12891 (N_12891,N_12331,N_12441);
nor U12892 (N_12892,N_12599,N_12594);
xor U12893 (N_12893,N_12492,N_12361);
xnor U12894 (N_12894,N_12329,N_12407);
nand U12895 (N_12895,N_12449,N_12335);
or U12896 (N_12896,N_12414,N_12562);
xor U12897 (N_12897,N_12366,N_12323);
xor U12898 (N_12898,N_12550,N_12458);
xor U12899 (N_12899,N_12488,N_12530);
nor U12900 (N_12900,N_12734,N_12614);
or U12901 (N_12901,N_12673,N_12812);
nor U12902 (N_12902,N_12661,N_12674);
xnor U12903 (N_12903,N_12784,N_12692);
xor U12904 (N_12904,N_12702,N_12625);
nor U12905 (N_12905,N_12847,N_12885);
or U12906 (N_12906,N_12735,N_12608);
or U12907 (N_12907,N_12835,N_12670);
and U12908 (N_12908,N_12823,N_12886);
or U12909 (N_12909,N_12752,N_12790);
nor U12910 (N_12910,N_12783,N_12657);
xnor U12911 (N_12911,N_12775,N_12789);
or U12912 (N_12912,N_12758,N_12806);
and U12913 (N_12913,N_12719,N_12642);
xor U12914 (N_12914,N_12894,N_12677);
nor U12915 (N_12915,N_12818,N_12891);
xor U12916 (N_12916,N_12766,N_12792);
xor U12917 (N_12917,N_12620,N_12665);
nor U12918 (N_12918,N_12671,N_12730);
xnor U12919 (N_12919,N_12738,N_12870);
and U12920 (N_12920,N_12769,N_12774);
or U12921 (N_12921,N_12650,N_12816);
or U12922 (N_12922,N_12623,N_12753);
xnor U12923 (N_12923,N_12770,N_12841);
and U12924 (N_12924,N_12828,N_12741);
xnor U12925 (N_12925,N_12646,N_12807);
and U12926 (N_12926,N_12712,N_12703);
xor U12927 (N_12927,N_12706,N_12883);
or U12928 (N_12928,N_12853,N_12887);
nor U12929 (N_12929,N_12678,N_12714);
nor U12930 (N_12930,N_12618,N_12773);
nand U12931 (N_12931,N_12824,N_12662);
and U12932 (N_12932,N_12836,N_12852);
xnor U12933 (N_12933,N_12636,N_12669);
nor U12934 (N_12934,N_12869,N_12867);
and U12935 (N_12935,N_12861,N_12659);
or U12936 (N_12936,N_12781,N_12843);
nand U12937 (N_12937,N_12681,N_12604);
xor U12938 (N_12938,N_12685,N_12821);
and U12939 (N_12939,N_12873,N_12811);
nor U12940 (N_12940,N_12856,N_12667);
and U12941 (N_12941,N_12850,N_12876);
and U12942 (N_12942,N_12645,N_12663);
xor U12943 (N_12943,N_12800,N_12696);
xnor U12944 (N_12944,N_12787,N_12820);
and U12945 (N_12945,N_12763,N_12635);
or U12946 (N_12946,N_12822,N_12672);
nand U12947 (N_12947,N_12704,N_12728);
and U12948 (N_12948,N_12640,N_12866);
nor U12949 (N_12949,N_12854,N_12605);
or U12950 (N_12950,N_12621,N_12690);
xnor U12951 (N_12951,N_12740,N_12842);
xnor U12952 (N_12952,N_12743,N_12855);
or U12953 (N_12953,N_12793,N_12709);
xor U12954 (N_12954,N_12615,N_12797);
and U12955 (N_12955,N_12808,N_12746);
xor U12956 (N_12956,N_12813,N_12759);
or U12957 (N_12957,N_12664,N_12733);
nand U12958 (N_12958,N_12622,N_12871);
nand U12959 (N_12959,N_12760,N_12837);
nand U12960 (N_12960,N_12742,N_12627);
nor U12961 (N_12961,N_12701,N_12831);
and U12962 (N_12962,N_12751,N_12731);
nand U12963 (N_12963,N_12711,N_12654);
or U12964 (N_12964,N_12683,N_12624);
nor U12965 (N_12965,N_12868,N_12827);
nand U12966 (N_12966,N_12691,N_12882);
nor U12967 (N_12967,N_12892,N_12802);
and U12968 (N_12968,N_12647,N_12884);
or U12969 (N_12969,N_12705,N_12680);
nor U12970 (N_12970,N_12641,N_12610);
or U12971 (N_12971,N_12778,N_12767);
nor U12972 (N_12972,N_12632,N_12798);
and U12973 (N_12973,N_12805,N_12780);
nor U12974 (N_12974,N_12757,N_12720);
nand U12975 (N_12975,N_12708,N_12832);
and U12976 (N_12976,N_12717,N_12729);
or U12977 (N_12977,N_12791,N_12795);
xnor U12978 (N_12978,N_12765,N_12803);
nor U12979 (N_12979,N_12637,N_12675);
nand U12980 (N_12980,N_12631,N_12838);
and U12981 (N_12981,N_12893,N_12655);
and U12982 (N_12982,N_12676,N_12602);
nor U12983 (N_12983,N_12679,N_12814);
or U12984 (N_12984,N_12653,N_12737);
and U12985 (N_12985,N_12648,N_12739);
or U12986 (N_12986,N_12609,N_12755);
or U12987 (N_12987,N_12628,N_12688);
nor U12988 (N_12988,N_12693,N_12710);
and U12989 (N_12989,N_12833,N_12682);
nor U12990 (N_12990,N_12629,N_12687);
nand U12991 (N_12991,N_12859,N_12777);
nor U12992 (N_12992,N_12601,N_12723);
nor U12993 (N_12993,N_12699,N_12825);
or U12994 (N_12994,N_12858,N_12889);
nand U12995 (N_12995,N_12736,N_12722);
nor U12996 (N_12996,N_12749,N_12656);
or U12997 (N_12997,N_12762,N_12619);
nand U12998 (N_12998,N_12897,N_12877);
nand U12999 (N_12999,N_12772,N_12606);
nand U13000 (N_13000,N_12694,N_12617);
and U13001 (N_13001,N_12810,N_12768);
nand U13002 (N_13002,N_12689,N_12638);
xnor U13003 (N_13003,N_12698,N_12863);
and U13004 (N_13004,N_12616,N_12639);
xnor U13005 (N_13005,N_12845,N_12754);
xor U13006 (N_13006,N_12668,N_12878);
or U13007 (N_13007,N_12840,N_12874);
xnor U13008 (N_13008,N_12809,N_12695);
or U13009 (N_13009,N_12611,N_12713);
or U13010 (N_13010,N_12651,N_12785);
and U13011 (N_13011,N_12643,N_12819);
xnor U13012 (N_13012,N_12849,N_12815);
nand U13013 (N_13013,N_12875,N_12830);
nand U13014 (N_13014,N_12846,N_12761);
xnor U13015 (N_13015,N_12817,N_12748);
and U13016 (N_13016,N_12851,N_12724);
and U13017 (N_13017,N_12686,N_12839);
nor U13018 (N_13018,N_12633,N_12796);
xor U13019 (N_13019,N_12727,N_12750);
nor U13020 (N_13020,N_12744,N_12786);
nand U13021 (N_13021,N_12794,N_12895);
nand U13022 (N_13022,N_12799,N_12864);
xor U13023 (N_13023,N_12862,N_12776);
nand U13024 (N_13024,N_12652,N_12607);
nor U13025 (N_13025,N_12844,N_12644);
xor U13026 (N_13026,N_12881,N_12718);
nand U13027 (N_13027,N_12603,N_12834);
xnor U13028 (N_13028,N_12879,N_12860);
nor U13029 (N_13029,N_12613,N_12700);
xnor U13030 (N_13030,N_12801,N_12697);
nor U13031 (N_13031,N_12865,N_12899);
or U13032 (N_13032,N_12764,N_12896);
nor U13033 (N_13033,N_12626,N_12721);
and U13034 (N_13034,N_12612,N_12600);
nor U13035 (N_13035,N_12716,N_12782);
nor U13036 (N_13036,N_12779,N_12725);
nor U13037 (N_13037,N_12649,N_12715);
or U13038 (N_13038,N_12726,N_12756);
or U13039 (N_13039,N_12747,N_12732);
nand U13040 (N_13040,N_12872,N_12666);
xor U13041 (N_13041,N_12660,N_12888);
and U13042 (N_13042,N_12771,N_12745);
nor U13043 (N_13043,N_12829,N_12658);
xnor U13044 (N_13044,N_12848,N_12804);
xnor U13045 (N_13045,N_12826,N_12707);
and U13046 (N_13046,N_12788,N_12857);
xnor U13047 (N_13047,N_12890,N_12880);
and U13048 (N_13048,N_12634,N_12630);
or U13049 (N_13049,N_12898,N_12684);
nand U13050 (N_13050,N_12756,N_12616);
xor U13051 (N_13051,N_12896,N_12877);
nor U13052 (N_13052,N_12835,N_12885);
nand U13053 (N_13053,N_12646,N_12723);
and U13054 (N_13054,N_12687,N_12657);
nand U13055 (N_13055,N_12832,N_12848);
nand U13056 (N_13056,N_12798,N_12753);
and U13057 (N_13057,N_12691,N_12664);
and U13058 (N_13058,N_12639,N_12773);
xor U13059 (N_13059,N_12884,N_12682);
nand U13060 (N_13060,N_12867,N_12871);
or U13061 (N_13061,N_12633,N_12659);
and U13062 (N_13062,N_12632,N_12704);
nor U13063 (N_13063,N_12717,N_12744);
and U13064 (N_13064,N_12706,N_12810);
nor U13065 (N_13065,N_12830,N_12772);
nor U13066 (N_13066,N_12677,N_12891);
and U13067 (N_13067,N_12775,N_12689);
nor U13068 (N_13068,N_12762,N_12743);
nor U13069 (N_13069,N_12623,N_12643);
or U13070 (N_13070,N_12664,N_12871);
and U13071 (N_13071,N_12827,N_12705);
nand U13072 (N_13072,N_12631,N_12744);
xnor U13073 (N_13073,N_12798,N_12768);
and U13074 (N_13074,N_12680,N_12656);
xor U13075 (N_13075,N_12729,N_12836);
nor U13076 (N_13076,N_12861,N_12818);
and U13077 (N_13077,N_12762,N_12733);
nand U13078 (N_13078,N_12610,N_12743);
xnor U13079 (N_13079,N_12678,N_12845);
nand U13080 (N_13080,N_12728,N_12612);
xor U13081 (N_13081,N_12799,N_12647);
xnor U13082 (N_13082,N_12719,N_12621);
nand U13083 (N_13083,N_12796,N_12861);
xor U13084 (N_13084,N_12723,N_12800);
nor U13085 (N_13085,N_12674,N_12882);
xor U13086 (N_13086,N_12840,N_12687);
or U13087 (N_13087,N_12737,N_12648);
xor U13088 (N_13088,N_12706,N_12702);
xor U13089 (N_13089,N_12880,N_12666);
nor U13090 (N_13090,N_12766,N_12648);
nor U13091 (N_13091,N_12608,N_12791);
or U13092 (N_13092,N_12729,N_12748);
or U13093 (N_13093,N_12727,N_12852);
xor U13094 (N_13094,N_12634,N_12811);
nand U13095 (N_13095,N_12713,N_12776);
xor U13096 (N_13096,N_12681,N_12620);
or U13097 (N_13097,N_12680,N_12874);
or U13098 (N_13098,N_12665,N_12818);
nor U13099 (N_13099,N_12886,N_12807);
xnor U13100 (N_13100,N_12647,N_12843);
nand U13101 (N_13101,N_12898,N_12762);
nor U13102 (N_13102,N_12604,N_12624);
nor U13103 (N_13103,N_12693,N_12824);
or U13104 (N_13104,N_12847,N_12695);
xnor U13105 (N_13105,N_12661,N_12857);
and U13106 (N_13106,N_12724,N_12679);
and U13107 (N_13107,N_12823,N_12640);
and U13108 (N_13108,N_12757,N_12868);
xor U13109 (N_13109,N_12685,N_12826);
xnor U13110 (N_13110,N_12834,N_12774);
nand U13111 (N_13111,N_12636,N_12784);
or U13112 (N_13112,N_12872,N_12863);
nor U13113 (N_13113,N_12746,N_12789);
or U13114 (N_13114,N_12812,N_12827);
or U13115 (N_13115,N_12878,N_12615);
nor U13116 (N_13116,N_12754,N_12893);
nor U13117 (N_13117,N_12796,N_12754);
nand U13118 (N_13118,N_12713,N_12807);
nand U13119 (N_13119,N_12859,N_12679);
nor U13120 (N_13120,N_12898,N_12823);
xor U13121 (N_13121,N_12685,N_12643);
nand U13122 (N_13122,N_12881,N_12697);
and U13123 (N_13123,N_12879,N_12866);
or U13124 (N_13124,N_12736,N_12616);
and U13125 (N_13125,N_12883,N_12735);
xnor U13126 (N_13126,N_12807,N_12707);
nor U13127 (N_13127,N_12758,N_12682);
nand U13128 (N_13128,N_12681,N_12680);
xnor U13129 (N_13129,N_12604,N_12605);
and U13130 (N_13130,N_12761,N_12829);
xor U13131 (N_13131,N_12818,N_12740);
or U13132 (N_13132,N_12737,N_12741);
and U13133 (N_13133,N_12770,N_12755);
nand U13134 (N_13134,N_12788,N_12763);
and U13135 (N_13135,N_12780,N_12796);
or U13136 (N_13136,N_12684,N_12671);
and U13137 (N_13137,N_12838,N_12628);
or U13138 (N_13138,N_12847,N_12764);
xnor U13139 (N_13139,N_12723,N_12651);
nand U13140 (N_13140,N_12751,N_12872);
and U13141 (N_13141,N_12780,N_12876);
nand U13142 (N_13142,N_12895,N_12820);
xor U13143 (N_13143,N_12799,N_12686);
nor U13144 (N_13144,N_12773,N_12659);
and U13145 (N_13145,N_12651,N_12895);
xnor U13146 (N_13146,N_12662,N_12708);
nor U13147 (N_13147,N_12841,N_12686);
or U13148 (N_13148,N_12694,N_12824);
xor U13149 (N_13149,N_12874,N_12755);
nand U13150 (N_13150,N_12762,N_12610);
or U13151 (N_13151,N_12788,N_12699);
nor U13152 (N_13152,N_12760,N_12768);
or U13153 (N_13153,N_12730,N_12821);
nor U13154 (N_13154,N_12806,N_12673);
or U13155 (N_13155,N_12845,N_12632);
nor U13156 (N_13156,N_12878,N_12728);
or U13157 (N_13157,N_12787,N_12735);
xnor U13158 (N_13158,N_12873,N_12657);
or U13159 (N_13159,N_12859,N_12821);
or U13160 (N_13160,N_12853,N_12870);
xnor U13161 (N_13161,N_12683,N_12796);
and U13162 (N_13162,N_12866,N_12695);
or U13163 (N_13163,N_12856,N_12720);
and U13164 (N_13164,N_12895,N_12780);
nand U13165 (N_13165,N_12816,N_12630);
and U13166 (N_13166,N_12770,N_12790);
nand U13167 (N_13167,N_12811,N_12792);
and U13168 (N_13168,N_12734,N_12704);
or U13169 (N_13169,N_12837,N_12862);
nand U13170 (N_13170,N_12862,N_12623);
or U13171 (N_13171,N_12899,N_12677);
or U13172 (N_13172,N_12844,N_12662);
and U13173 (N_13173,N_12726,N_12777);
xor U13174 (N_13174,N_12629,N_12854);
xnor U13175 (N_13175,N_12763,N_12895);
and U13176 (N_13176,N_12654,N_12612);
nand U13177 (N_13177,N_12899,N_12709);
or U13178 (N_13178,N_12704,N_12813);
and U13179 (N_13179,N_12613,N_12853);
and U13180 (N_13180,N_12619,N_12601);
and U13181 (N_13181,N_12678,N_12865);
nor U13182 (N_13182,N_12761,N_12610);
xnor U13183 (N_13183,N_12749,N_12612);
nor U13184 (N_13184,N_12738,N_12835);
and U13185 (N_13185,N_12604,N_12678);
or U13186 (N_13186,N_12604,N_12668);
or U13187 (N_13187,N_12737,N_12828);
nand U13188 (N_13188,N_12757,N_12743);
nor U13189 (N_13189,N_12743,N_12731);
or U13190 (N_13190,N_12666,N_12699);
and U13191 (N_13191,N_12730,N_12803);
and U13192 (N_13192,N_12899,N_12735);
nor U13193 (N_13193,N_12617,N_12889);
or U13194 (N_13194,N_12677,N_12724);
nand U13195 (N_13195,N_12650,N_12781);
nor U13196 (N_13196,N_12766,N_12778);
or U13197 (N_13197,N_12687,N_12609);
and U13198 (N_13198,N_12634,N_12758);
xor U13199 (N_13199,N_12667,N_12607);
xor U13200 (N_13200,N_13003,N_12923);
and U13201 (N_13201,N_13197,N_13058);
xnor U13202 (N_13202,N_13179,N_13181);
nor U13203 (N_13203,N_13029,N_12988);
and U13204 (N_13204,N_13123,N_13004);
nand U13205 (N_13205,N_13174,N_13195);
or U13206 (N_13206,N_13001,N_12954);
nand U13207 (N_13207,N_12972,N_12986);
nor U13208 (N_13208,N_12936,N_13168);
and U13209 (N_13209,N_13173,N_13180);
xnor U13210 (N_13210,N_13120,N_12960);
nor U13211 (N_13211,N_13060,N_13071);
and U13212 (N_13212,N_13145,N_12966);
or U13213 (N_13213,N_13115,N_13076);
xor U13214 (N_13214,N_13118,N_13089);
xnor U13215 (N_13215,N_12999,N_12927);
nand U13216 (N_13216,N_12944,N_13155);
xnor U13217 (N_13217,N_12953,N_13091);
nor U13218 (N_13218,N_13176,N_13194);
or U13219 (N_13219,N_13038,N_12925);
or U13220 (N_13220,N_13104,N_12942);
and U13221 (N_13221,N_12967,N_13014);
or U13222 (N_13222,N_13010,N_13082);
and U13223 (N_13223,N_13033,N_12955);
nand U13224 (N_13224,N_13070,N_12948);
nor U13225 (N_13225,N_12971,N_13059);
and U13226 (N_13226,N_13093,N_12935);
xnor U13227 (N_13227,N_13077,N_12916);
and U13228 (N_13228,N_12973,N_13011);
xor U13229 (N_13229,N_12996,N_13007);
or U13230 (N_13230,N_12911,N_13121);
nand U13231 (N_13231,N_12984,N_13061);
and U13232 (N_13232,N_13156,N_13040);
or U13233 (N_13233,N_12902,N_13138);
nor U13234 (N_13234,N_13063,N_12909);
nand U13235 (N_13235,N_12932,N_12945);
or U13236 (N_13236,N_13160,N_12982);
and U13237 (N_13237,N_13024,N_13162);
xnor U13238 (N_13238,N_13053,N_13035);
or U13239 (N_13239,N_12900,N_12930);
or U13240 (N_13240,N_13133,N_12946);
nand U13241 (N_13241,N_12961,N_13027);
and U13242 (N_13242,N_13049,N_12993);
and U13243 (N_13243,N_12924,N_12974);
and U13244 (N_13244,N_12949,N_12938);
and U13245 (N_13245,N_13086,N_13094);
nand U13246 (N_13246,N_13039,N_12987);
nand U13247 (N_13247,N_12983,N_13171);
nor U13248 (N_13248,N_13013,N_13129);
nor U13249 (N_13249,N_13128,N_13099);
nor U13250 (N_13250,N_13166,N_13187);
and U13251 (N_13251,N_12964,N_13017);
or U13252 (N_13252,N_12940,N_13054);
nand U13253 (N_13253,N_13127,N_12952);
and U13254 (N_13254,N_13144,N_13066);
and U13255 (N_13255,N_13103,N_13164);
nor U13256 (N_13256,N_13170,N_13012);
nor U13257 (N_13257,N_12912,N_13079);
nor U13258 (N_13258,N_13177,N_13002);
and U13259 (N_13259,N_13008,N_13074);
xnor U13260 (N_13260,N_13126,N_12978);
or U13261 (N_13261,N_13131,N_13030);
and U13262 (N_13262,N_13158,N_13106);
xor U13263 (N_13263,N_13031,N_13041);
xor U13264 (N_13264,N_13167,N_12981);
xnor U13265 (N_13265,N_13186,N_12931);
or U13266 (N_13266,N_13023,N_13134);
and U13267 (N_13267,N_12962,N_13080);
and U13268 (N_13268,N_12970,N_13097);
xnor U13269 (N_13269,N_13119,N_13005);
nand U13270 (N_13270,N_13178,N_13087);
nor U13271 (N_13271,N_12933,N_13078);
or U13272 (N_13272,N_12904,N_12959);
xor U13273 (N_13273,N_12950,N_13062);
nor U13274 (N_13274,N_12926,N_13188);
nor U13275 (N_13275,N_13184,N_13142);
and U13276 (N_13276,N_13015,N_12937);
or U13277 (N_13277,N_12919,N_13048);
xnor U13278 (N_13278,N_13037,N_13009);
nand U13279 (N_13279,N_13175,N_13021);
nand U13280 (N_13280,N_13096,N_13107);
nand U13281 (N_13281,N_13139,N_13148);
nor U13282 (N_13282,N_13032,N_12997);
xor U13283 (N_13283,N_13110,N_13132);
xor U13284 (N_13284,N_12913,N_13075);
and U13285 (N_13285,N_13192,N_13045);
nor U13286 (N_13286,N_12980,N_13057);
nor U13287 (N_13287,N_13137,N_13102);
xor U13288 (N_13288,N_13067,N_13146);
nor U13289 (N_13289,N_12977,N_12975);
nor U13290 (N_13290,N_12963,N_12910);
nor U13291 (N_13291,N_13189,N_12956);
and U13292 (N_13292,N_13199,N_13073);
nor U13293 (N_13293,N_13072,N_13114);
xor U13294 (N_13294,N_13191,N_13163);
and U13295 (N_13295,N_13105,N_13182);
and U13296 (N_13296,N_13055,N_13081);
xnor U13297 (N_13297,N_13151,N_13141);
and U13298 (N_13298,N_13034,N_13028);
xor U13299 (N_13299,N_12907,N_12934);
nand U13300 (N_13300,N_13159,N_12908);
xnor U13301 (N_13301,N_12915,N_13092);
or U13302 (N_13302,N_13095,N_12928);
nor U13303 (N_13303,N_13190,N_13154);
or U13304 (N_13304,N_13064,N_12920);
nor U13305 (N_13305,N_12921,N_13098);
nand U13306 (N_13306,N_12990,N_13016);
nor U13307 (N_13307,N_13196,N_13113);
nor U13308 (N_13308,N_13026,N_13125);
xnor U13309 (N_13309,N_13172,N_13050);
xnor U13310 (N_13310,N_13185,N_13143);
or U13311 (N_13311,N_12939,N_12985);
nand U13312 (N_13312,N_12991,N_12905);
or U13313 (N_13313,N_13036,N_13000);
xor U13314 (N_13314,N_13068,N_13088);
and U13315 (N_13315,N_12922,N_13006);
or U13316 (N_13316,N_13044,N_13124);
and U13317 (N_13317,N_12917,N_12951);
or U13318 (N_13318,N_12906,N_13020);
xor U13319 (N_13319,N_13165,N_13183);
and U13320 (N_13320,N_12994,N_12918);
or U13321 (N_13321,N_13147,N_13108);
and U13322 (N_13322,N_13135,N_12914);
xnor U13323 (N_13323,N_13198,N_13161);
xor U13324 (N_13324,N_13117,N_13018);
xnor U13325 (N_13325,N_13157,N_13065);
xor U13326 (N_13326,N_12958,N_13100);
nand U13327 (N_13327,N_12995,N_13084);
and U13328 (N_13328,N_13111,N_13025);
nand U13329 (N_13329,N_13109,N_13193);
nor U13330 (N_13330,N_13042,N_12979);
xor U13331 (N_13331,N_13101,N_12968);
nor U13332 (N_13332,N_12947,N_13056);
and U13333 (N_13333,N_13085,N_13047);
or U13334 (N_13334,N_13140,N_13043);
nor U13335 (N_13335,N_12976,N_13051);
or U13336 (N_13336,N_12998,N_13122);
nand U13337 (N_13337,N_13069,N_12992);
nor U13338 (N_13338,N_13130,N_13022);
nor U13339 (N_13339,N_12969,N_13150);
xor U13340 (N_13340,N_13052,N_13136);
xnor U13341 (N_13341,N_13090,N_12989);
nand U13342 (N_13342,N_12965,N_13083);
nand U13343 (N_13343,N_13046,N_13153);
xor U13344 (N_13344,N_13116,N_12943);
or U13345 (N_13345,N_13149,N_13169);
or U13346 (N_13346,N_13112,N_12901);
nor U13347 (N_13347,N_12941,N_13152);
xnor U13348 (N_13348,N_12903,N_13019);
or U13349 (N_13349,N_12957,N_12929);
nand U13350 (N_13350,N_13072,N_13002);
nand U13351 (N_13351,N_13052,N_13021);
or U13352 (N_13352,N_12942,N_12917);
nand U13353 (N_13353,N_13180,N_12904);
nor U13354 (N_13354,N_12929,N_13050);
or U13355 (N_13355,N_12933,N_13056);
xor U13356 (N_13356,N_13065,N_12955);
nor U13357 (N_13357,N_12936,N_13135);
nand U13358 (N_13358,N_13089,N_13030);
or U13359 (N_13359,N_13091,N_13079);
and U13360 (N_13360,N_13175,N_13181);
nand U13361 (N_13361,N_12927,N_13070);
and U13362 (N_13362,N_12994,N_12946);
or U13363 (N_13363,N_13079,N_13125);
or U13364 (N_13364,N_13046,N_12997);
or U13365 (N_13365,N_12993,N_13014);
nor U13366 (N_13366,N_13054,N_12999);
and U13367 (N_13367,N_13178,N_12926);
xor U13368 (N_13368,N_13101,N_12983);
xnor U13369 (N_13369,N_12968,N_12996);
and U13370 (N_13370,N_12941,N_12961);
nor U13371 (N_13371,N_13087,N_13147);
or U13372 (N_13372,N_12973,N_13049);
and U13373 (N_13373,N_12933,N_12988);
xnor U13374 (N_13374,N_13078,N_12957);
and U13375 (N_13375,N_13031,N_13048);
nor U13376 (N_13376,N_13048,N_13131);
nand U13377 (N_13377,N_12974,N_12912);
nor U13378 (N_13378,N_13097,N_12974);
nand U13379 (N_13379,N_13120,N_13121);
nor U13380 (N_13380,N_13031,N_13183);
nor U13381 (N_13381,N_13049,N_13174);
xor U13382 (N_13382,N_13078,N_13126);
nor U13383 (N_13383,N_12997,N_13050);
nand U13384 (N_13384,N_13004,N_13064);
xor U13385 (N_13385,N_13182,N_12926);
xor U13386 (N_13386,N_13195,N_13184);
or U13387 (N_13387,N_12936,N_12919);
nor U13388 (N_13388,N_12967,N_13113);
and U13389 (N_13389,N_13060,N_12972);
xnor U13390 (N_13390,N_12925,N_13025);
xor U13391 (N_13391,N_12906,N_13021);
nand U13392 (N_13392,N_13142,N_12992);
nor U13393 (N_13393,N_13111,N_12947);
and U13394 (N_13394,N_13087,N_13115);
or U13395 (N_13395,N_13136,N_13055);
xor U13396 (N_13396,N_13124,N_13117);
nand U13397 (N_13397,N_13073,N_13145);
xor U13398 (N_13398,N_12991,N_12915);
xor U13399 (N_13399,N_13102,N_12970);
nand U13400 (N_13400,N_13161,N_13066);
and U13401 (N_13401,N_12984,N_12974);
and U13402 (N_13402,N_12941,N_13072);
or U13403 (N_13403,N_12996,N_13188);
nand U13404 (N_13404,N_13028,N_13113);
nor U13405 (N_13405,N_13056,N_12951);
and U13406 (N_13406,N_12982,N_12906);
and U13407 (N_13407,N_13046,N_13036);
and U13408 (N_13408,N_13132,N_12984);
nand U13409 (N_13409,N_13048,N_12959);
or U13410 (N_13410,N_13068,N_12991);
or U13411 (N_13411,N_13144,N_13039);
xnor U13412 (N_13412,N_13021,N_12990);
or U13413 (N_13413,N_12901,N_12951);
or U13414 (N_13414,N_13164,N_12970);
and U13415 (N_13415,N_13167,N_13179);
nand U13416 (N_13416,N_13054,N_13053);
nand U13417 (N_13417,N_13187,N_13176);
xor U13418 (N_13418,N_13160,N_13094);
or U13419 (N_13419,N_13022,N_12999);
nor U13420 (N_13420,N_12966,N_13151);
nor U13421 (N_13421,N_13161,N_13186);
or U13422 (N_13422,N_13007,N_12949);
nand U13423 (N_13423,N_13174,N_13173);
nor U13424 (N_13424,N_12969,N_12929);
nand U13425 (N_13425,N_13122,N_13109);
xnor U13426 (N_13426,N_12981,N_13039);
nand U13427 (N_13427,N_13032,N_13164);
and U13428 (N_13428,N_12998,N_13124);
nor U13429 (N_13429,N_13049,N_13056);
nor U13430 (N_13430,N_13041,N_13044);
nand U13431 (N_13431,N_13170,N_13079);
or U13432 (N_13432,N_12981,N_12926);
or U13433 (N_13433,N_13157,N_13027);
and U13434 (N_13434,N_13087,N_12963);
or U13435 (N_13435,N_12997,N_13154);
nor U13436 (N_13436,N_13021,N_13132);
or U13437 (N_13437,N_12968,N_13124);
or U13438 (N_13438,N_12989,N_13188);
xor U13439 (N_13439,N_13027,N_12962);
nand U13440 (N_13440,N_13057,N_13170);
xnor U13441 (N_13441,N_13183,N_12914);
and U13442 (N_13442,N_12930,N_13057);
nor U13443 (N_13443,N_13066,N_13100);
nand U13444 (N_13444,N_12947,N_13155);
and U13445 (N_13445,N_13112,N_12970);
nor U13446 (N_13446,N_13071,N_12920);
xor U13447 (N_13447,N_13190,N_12947);
nand U13448 (N_13448,N_12995,N_13063);
or U13449 (N_13449,N_12912,N_12929);
nor U13450 (N_13450,N_13192,N_13010);
nand U13451 (N_13451,N_13065,N_13190);
xnor U13452 (N_13452,N_12935,N_13166);
or U13453 (N_13453,N_13141,N_13140);
xnor U13454 (N_13454,N_13052,N_13013);
nand U13455 (N_13455,N_12972,N_13048);
and U13456 (N_13456,N_13188,N_13161);
or U13457 (N_13457,N_13087,N_13049);
and U13458 (N_13458,N_13061,N_13141);
or U13459 (N_13459,N_13048,N_12911);
or U13460 (N_13460,N_13169,N_13063);
nand U13461 (N_13461,N_12925,N_13115);
nor U13462 (N_13462,N_12935,N_13142);
xnor U13463 (N_13463,N_13193,N_12949);
xor U13464 (N_13464,N_13007,N_12933);
nor U13465 (N_13465,N_13189,N_12958);
or U13466 (N_13466,N_13177,N_12960);
nand U13467 (N_13467,N_12957,N_13079);
and U13468 (N_13468,N_13116,N_12904);
xor U13469 (N_13469,N_13006,N_12925);
nor U13470 (N_13470,N_13119,N_13093);
nor U13471 (N_13471,N_13187,N_12963);
nand U13472 (N_13472,N_13145,N_13020);
or U13473 (N_13473,N_13051,N_13126);
and U13474 (N_13474,N_13183,N_13023);
xnor U13475 (N_13475,N_13143,N_12990);
and U13476 (N_13476,N_13012,N_13112);
nand U13477 (N_13477,N_13091,N_12922);
xor U13478 (N_13478,N_13160,N_13085);
or U13479 (N_13479,N_12971,N_13166);
xor U13480 (N_13480,N_12922,N_12911);
or U13481 (N_13481,N_12986,N_13132);
xnor U13482 (N_13482,N_13070,N_12922);
nand U13483 (N_13483,N_12988,N_12901);
and U13484 (N_13484,N_12969,N_13170);
nand U13485 (N_13485,N_12933,N_13050);
nand U13486 (N_13486,N_13088,N_13149);
nand U13487 (N_13487,N_12955,N_12979);
and U13488 (N_13488,N_12963,N_12915);
nor U13489 (N_13489,N_13136,N_12964);
nor U13490 (N_13490,N_12921,N_13079);
or U13491 (N_13491,N_13033,N_13100);
or U13492 (N_13492,N_13147,N_13105);
xnor U13493 (N_13493,N_13003,N_12937);
nor U13494 (N_13494,N_13156,N_13172);
nand U13495 (N_13495,N_13012,N_12967);
nor U13496 (N_13496,N_12970,N_12965);
nand U13497 (N_13497,N_12911,N_13189);
or U13498 (N_13498,N_13104,N_12963);
nand U13499 (N_13499,N_13121,N_13003);
nand U13500 (N_13500,N_13200,N_13278);
xnor U13501 (N_13501,N_13381,N_13444);
nand U13502 (N_13502,N_13385,N_13372);
and U13503 (N_13503,N_13399,N_13313);
xnor U13504 (N_13504,N_13447,N_13338);
or U13505 (N_13505,N_13300,N_13465);
nor U13506 (N_13506,N_13449,N_13394);
xor U13507 (N_13507,N_13322,N_13389);
or U13508 (N_13508,N_13224,N_13487);
xnor U13509 (N_13509,N_13467,N_13301);
or U13510 (N_13510,N_13423,N_13493);
nand U13511 (N_13511,N_13247,N_13341);
nand U13512 (N_13512,N_13482,N_13375);
or U13513 (N_13513,N_13284,N_13456);
and U13514 (N_13514,N_13431,N_13489);
nand U13515 (N_13515,N_13239,N_13445);
nor U13516 (N_13516,N_13435,N_13241);
xor U13517 (N_13517,N_13443,N_13327);
nor U13518 (N_13518,N_13472,N_13373);
nand U13519 (N_13519,N_13370,N_13417);
xor U13520 (N_13520,N_13331,N_13347);
xor U13521 (N_13521,N_13228,N_13409);
xnor U13522 (N_13522,N_13433,N_13477);
xor U13523 (N_13523,N_13219,N_13234);
nor U13524 (N_13524,N_13237,N_13216);
nand U13525 (N_13525,N_13274,N_13292);
nand U13526 (N_13526,N_13289,N_13392);
nor U13527 (N_13527,N_13256,N_13201);
and U13528 (N_13528,N_13350,N_13494);
and U13529 (N_13529,N_13383,N_13344);
or U13530 (N_13530,N_13400,N_13458);
or U13531 (N_13531,N_13488,N_13388);
or U13532 (N_13532,N_13242,N_13474);
xnor U13533 (N_13533,N_13215,N_13323);
nor U13534 (N_13534,N_13325,N_13471);
nand U13535 (N_13535,N_13430,N_13238);
xnor U13536 (N_13536,N_13236,N_13280);
or U13537 (N_13537,N_13360,N_13438);
xor U13538 (N_13538,N_13273,N_13211);
nor U13539 (N_13539,N_13229,N_13422);
or U13540 (N_13540,N_13208,N_13426);
or U13541 (N_13541,N_13490,N_13379);
nor U13542 (N_13542,N_13272,N_13315);
and U13543 (N_13543,N_13269,N_13479);
xor U13544 (N_13544,N_13262,N_13218);
or U13545 (N_13545,N_13421,N_13251);
xnor U13546 (N_13546,N_13440,N_13317);
xnor U13547 (N_13547,N_13398,N_13304);
or U13548 (N_13548,N_13222,N_13221);
and U13549 (N_13549,N_13436,N_13408);
and U13550 (N_13550,N_13481,N_13276);
or U13551 (N_13551,N_13265,N_13299);
xor U13552 (N_13552,N_13448,N_13346);
xor U13553 (N_13553,N_13460,N_13281);
nand U13554 (N_13554,N_13419,N_13232);
xnor U13555 (N_13555,N_13285,N_13351);
or U13556 (N_13556,N_13457,N_13478);
or U13557 (N_13557,N_13476,N_13428);
or U13558 (N_13558,N_13204,N_13441);
and U13559 (N_13559,N_13427,N_13283);
nor U13560 (N_13560,N_13453,N_13357);
xnor U13561 (N_13561,N_13459,N_13287);
or U13562 (N_13562,N_13326,N_13290);
and U13563 (N_13563,N_13442,N_13384);
and U13564 (N_13564,N_13295,N_13377);
or U13565 (N_13565,N_13318,N_13393);
nor U13566 (N_13566,N_13291,N_13450);
nor U13567 (N_13567,N_13212,N_13244);
xor U13568 (N_13568,N_13332,N_13374);
nor U13569 (N_13569,N_13258,N_13483);
or U13570 (N_13570,N_13279,N_13312);
xnor U13571 (N_13571,N_13249,N_13252);
or U13572 (N_13572,N_13452,N_13468);
or U13573 (N_13573,N_13412,N_13434);
or U13574 (N_13574,N_13397,N_13402);
and U13575 (N_13575,N_13297,N_13316);
or U13576 (N_13576,N_13491,N_13454);
nand U13577 (N_13577,N_13425,N_13282);
nor U13578 (N_13578,N_13217,N_13210);
or U13579 (N_13579,N_13293,N_13306);
xor U13580 (N_13580,N_13275,N_13432);
or U13581 (N_13581,N_13495,N_13213);
nand U13582 (N_13582,N_13356,N_13206);
nand U13583 (N_13583,N_13387,N_13345);
nor U13584 (N_13584,N_13334,N_13255);
nand U13585 (N_13585,N_13260,N_13473);
nand U13586 (N_13586,N_13266,N_13407);
nand U13587 (N_13587,N_13404,N_13309);
and U13588 (N_13588,N_13314,N_13391);
and U13589 (N_13589,N_13263,N_13461);
or U13590 (N_13590,N_13369,N_13203);
nand U13591 (N_13591,N_13277,N_13390);
and U13592 (N_13592,N_13378,N_13348);
and U13593 (N_13593,N_13340,N_13336);
and U13594 (N_13594,N_13361,N_13451);
and U13595 (N_13595,N_13288,N_13466);
or U13596 (N_13596,N_13376,N_13366);
and U13597 (N_13597,N_13437,N_13416);
xor U13598 (N_13598,N_13358,N_13329);
xor U13599 (N_13599,N_13424,N_13324);
nand U13600 (N_13600,N_13305,N_13268);
nand U13601 (N_13601,N_13270,N_13420);
nor U13602 (N_13602,N_13259,N_13455);
and U13603 (N_13603,N_13342,N_13261);
and U13604 (N_13604,N_13207,N_13253);
or U13605 (N_13605,N_13371,N_13298);
and U13606 (N_13606,N_13202,N_13320);
xor U13607 (N_13607,N_13446,N_13264);
nand U13608 (N_13608,N_13227,N_13248);
and U13609 (N_13609,N_13233,N_13462);
nor U13610 (N_13610,N_13380,N_13496);
and U13611 (N_13611,N_13302,N_13497);
nor U13612 (N_13612,N_13246,N_13359);
or U13613 (N_13613,N_13339,N_13243);
or U13614 (N_13614,N_13245,N_13401);
nor U13615 (N_13615,N_13354,N_13226);
xor U13616 (N_13616,N_13439,N_13418);
nand U13617 (N_13617,N_13230,N_13363);
xnor U13618 (N_13618,N_13209,N_13386);
xnor U13619 (N_13619,N_13220,N_13231);
nor U13620 (N_13620,N_13254,N_13364);
or U13621 (N_13621,N_13365,N_13410);
or U13622 (N_13622,N_13485,N_13406);
nor U13623 (N_13623,N_13337,N_13308);
or U13624 (N_13624,N_13475,N_13403);
nand U13625 (N_13625,N_13480,N_13429);
and U13626 (N_13626,N_13362,N_13250);
nand U13627 (N_13627,N_13469,N_13225);
and U13628 (N_13628,N_13307,N_13311);
xnor U13629 (N_13629,N_13321,N_13240);
nor U13630 (N_13630,N_13319,N_13310);
nand U13631 (N_13631,N_13286,N_13223);
nor U13632 (N_13632,N_13464,N_13352);
or U13633 (N_13633,N_13343,N_13328);
or U13634 (N_13634,N_13294,N_13333);
xor U13635 (N_13635,N_13411,N_13395);
nor U13636 (N_13636,N_13492,N_13267);
nand U13637 (N_13637,N_13214,N_13484);
nor U13638 (N_13638,N_13415,N_13355);
xor U13639 (N_13639,N_13353,N_13486);
xnor U13640 (N_13640,N_13396,N_13470);
nor U13641 (N_13641,N_13296,N_13405);
nor U13642 (N_13642,N_13368,N_13303);
and U13643 (N_13643,N_13499,N_13367);
and U13644 (N_13644,N_13349,N_13235);
xor U13645 (N_13645,N_13257,N_13463);
nand U13646 (N_13646,N_13330,N_13335);
and U13647 (N_13647,N_13413,N_13271);
nand U13648 (N_13648,N_13205,N_13498);
or U13649 (N_13649,N_13382,N_13414);
nand U13650 (N_13650,N_13392,N_13211);
nand U13651 (N_13651,N_13406,N_13349);
and U13652 (N_13652,N_13390,N_13474);
nand U13653 (N_13653,N_13282,N_13446);
nor U13654 (N_13654,N_13229,N_13349);
xor U13655 (N_13655,N_13427,N_13443);
and U13656 (N_13656,N_13235,N_13454);
or U13657 (N_13657,N_13276,N_13349);
or U13658 (N_13658,N_13492,N_13259);
nor U13659 (N_13659,N_13474,N_13233);
or U13660 (N_13660,N_13322,N_13243);
nor U13661 (N_13661,N_13291,N_13281);
and U13662 (N_13662,N_13306,N_13339);
nand U13663 (N_13663,N_13440,N_13229);
nor U13664 (N_13664,N_13488,N_13297);
or U13665 (N_13665,N_13258,N_13409);
xnor U13666 (N_13666,N_13477,N_13424);
and U13667 (N_13667,N_13295,N_13411);
xnor U13668 (N_13668,N_13276,N_13420);
and U13669 (N_13669,N_13345,N_13286);
xnor U13670 (N_13670,N_13423,N_13225);
xor U13671 (N_13671,N_13318,N_13201);
xor U13672 (N_13672,N_13375,N_13499);
nor U13673 (N_13673,N_13353,N_13387);
and U13674 (N_13674,N_13390,N_13438);
nand U13675 (N_13675,N_13440,N_13372);
or U13676 (N_13676,N_13254,N_13260);
xnor U13677 (N_13677,N_13411,N_13231);
and U13678 (N_13678,N_13293,N_13448);
nand U13679 (N_13679,N_13466,N_13380);
or U13680 (N_13680,N_13223,N_13247);
and U13681 (N_13681,N_13292,N_13496);
xnor U13682 (N_13682,N_13489,N_13350);
nor U13683 (N_13683,N_13376,N_13409);
nand U13684 (N_13684,N_13284,N_13373);
nor U13685 (N_13685,N_13427,N_13312);
nor U13686 (N_13686,N_13302,N_13328);
xnor U13687 (N_13687,N_13494,N_13249);
xnor U13688 (N_13688,N_13297,N_13494);
or U13689 (N_13689,N_13427,N_13207);
or U13690 (N_13690,N_13430,N_13473);
xnor U13691 (N_13691,N_13290,N_13315);
nor U13692 (N_13692,N_13207,N_13276);
nor U13693 (N_13693,N_13307,N_13467);
and U13694 (N_13694,N_13368,N_13220);
nor U13695 (N_13695,N_13411,N_13377);
nor U13696 (N_13696,N_13445,N_13498);
and U13697 (N_13697,N_13479,N_13375);
or U13698 (N_13698,N_13377,N_13231);
and U13699 (N_13699,N_13413,N_13372);
and U13700 (N_13700,N_13397,N_13289);
nand U13701 (N_13701,N_13260,N_13456);
or U13702 (N_13702,N_13433,N_13352);
and U13703 (N_13703,N_13416,N_13428);
or U13704 (N_13704,N_13270,N_13296);
nor U13705 (N_13705,N_13297,N_13337);
xor U13706 (N_13706,N_13297,N_13491);
nor U13707 (N_13707,N_13458,N_13303);
and U13708 (N_13708,N_13247,N_13276);
or U13709 (N_13709,N_13285,N_13339);
and U13710 (N_13710,N_13414,N_13476);
or U13711 (N_13711,N_13303,N_13225);
or U13712 (N_13712,N_13321,N_13404);
nand U13713 (N_13713,N_13418,N_13374);
xnor U13714 (N_13714,N_13368,N_13400);
nor U13715 (N_13715,N_13297,N_13279);
xor U13716 (N_13716,N_13319,N_13307);
or U13717 (N_13717,N_13286,N_13295);
or U13718 (N_13718,N_13476,N_13351);
xnor U13719 (N_13719,N_13277,N_13371);
or U13720 (N_13720,N_13309,N_13323);
or U13721 (N_13721,N_13222,N_13203);
nor U13722 (N_13722,N_13418,N_13398);
and U13723 (N_13723,N_13374,N_13429);
nor U13724 (N_13724,N_13453,N_13374);
and U13725 (N_13725,N_13209,N_13266);
xor U13726 (N_13726,N_13298,N_13468);
xnor U13727 (N_13727,N_13206,N_13321);
or U13728 (N_13728,N_13495,N_13216);
nor U13729 (N_13729,N_13458,N_13294);
nand U13730 (N_13730,N_13383,N_13354);
nor U13731 (N_13731,N_13369,N_13459);
or U13732 (N_13732,N_13465,N_13249);
or U13733 (N_13733,N_13328,N_13317);
and U13734 (N_13734,N_13411,N_13330);
or U13735 (N_13735,N_13481,N_13304);
nand U13736 (N_13736,N_13210,N_13251);
nand U13737 (N_13737,N_13370,N_13409);
xnor U13738 (N_13738,N_13385,N_13298);
or U13739 (N_13739,N_13335,N_13320);
nand U13740 (N_13740,N_13498,N_13367);
and U13741 (N_13741,N_13486,N_13434);
nand U13742 (N_13742,N_13340,N_13379);
nor U13743 (N_13743,N_13312,N_13207);
nor U13744 (N_13744,N_13223,N_13260);
or U13745 (N_13745,N_13291,N_13209);
xnor U13746 (N_13746,N_13429,N_13367);
nand U13747 (N_13747,N_13481,N_13417);
nor U13748 (N_13748,N_13360,N_13490);
nand U13749 (N_13749,N_13475,N_13394);
nor U13750 (N_13750,N_13433,N_13359);
and U13751 (N_13751,N_13390,N_13356);
nand U13752 (N_13752,N_13488,N_13260);
nor U13753 (N_13753,N_13247,N_13499);
or U13754 (N_13754,N_13445,N_13327);
or U13755 (N_13755,N_13455,N_13219);
nand U13756 (N_13756,N_13357,N_13293);
nor U13757 (N_13757,N_13466,N_13300);
nor U13758 (N_13758,N_13498,N_13266);
and U13759 (N_13759,N_13290,N_13334);
nor U13760 (N_13760,N_13429,N_13461);
and U13761 (N_13761,N_13398,N_13442);
or U13762 (N_13762,N_13265,N_13464);
or U13763 (N_13763,N_13240,N_13463);
and U13764 (N_13764,N_13391,N_13482);
and U13765 (N_13765,N_13343,N_13276);
nor U13766 (N_13766,N_13226,N_13326);
nor U13767 (N_13767,N_13290,N_13433);
nor U13768 (N_13768,N_13260,N_13367);
nor U13769 (N_13769,N_13326,N_13306);
xor U13770 (N_13770,N_13229,N_13293);
nor U13771 (N_13771,N_13365,N_13374);
xor U13772 (N_13772,N_13389,N_13205);
and U13773 (N_13773,N_13272,N_13258);
or U13774 (N_13774,N_13248,N_13312);
or U13775 (N_13775,N_13309,N_13439);
or U13776 (N_13776,N_13342,N_13305);
and U13777 (N_13777,N_13445,N_13311);
or U13778 (N_13778,N_13394,N_13360);
nor U13779 (N_13779,N_13366,N_13379);
nand U13780 (N_13780,N_13408,N_13457);
nor U13781 (N_13781,N_13367,N_13405);
and U13782 (N_13782,N_13384,N_13303);
nand U13783 (N_13783,N_13402,N_13435);
nor U13784 (N_13784,N_13450,N_13468);
nand U13785 (N_13785,N_13225,N_13373);
xor U13786 (N_13786,N_13237,N_13413);
nor U13787 (N_13787,N_13245,N_13489);
or U13788 (N_13788,N_13362,N_13370);
and U13789 (N_13789,N_13345,N_13450);
or U13790 (N_13790,N_13209,N_13242);
nor U13791 (N_13791,N_13223,N_13388);
nand U13792 (N_13792,N_13345,N_13236);
and U13793 (N_13793,N_13267,N_13323);
nand U13794 (N_13794,N_13238,N_13366);
nor U13795 (N_13795,N_13413,N_13266);
xor U13796 (N_13796,N_13308,N_13285);
nand U13797 (N_13797,N_13446,N_13495);
and U13798 (N_13798,N_13450,N_13346);
xnor U13799 (N_13799,N_13422,N_13455);
or U13800 (N_13800,N_13605,N_13534);
and U13801 (N_13801,N_13540,N_13573);
xnor U13802 (N_13802,N_13570,N_13674);
nor U13803 (N_13803,N_13655,N_13682);
nor U13804 (N_13804,N_13600,N_13771);
and U13805 (N_13805,N_13630,N_13694);
nor U13806 (N_13806,N_13679,N_13724);
and U13807 (N_13807,N_13733,N_13618);
xnor U13808 (N_13808,N_13765,N_13639);
xnor U13809 (N_13809,N_13647,N_13508);
xor U13810 (N_13810,N_13525,N_13744);
xor U13811 (N_13811,N_13637,N_13565);
nor U13812 (N_13812,N_13640,N_13662);
and U13813 (N_13813,N_13753,N_13695);
nor U13814 (N_13814,N_13751,N_13675);
or U13815 (N_13815,N_13793,N_13601);
nand U13816 (N_13816,N_13629,N_13754);
nand U13817 (N_13817,N_13619,N_13726);
nand U13818 (N_13818,N_13773,N_13758);
nand U13819 (N_13819,N_13787,N_13799);
xnor U13820 (N_13820,N_13553,N_13645);
or U13821 (N_13821,N_13579,N_13720);
xnor U13822 (N_13822,N_13721,N_13556);
and U13823 (N_13823,N_13666,N_13652);
nand U13824 (N_13824,N_13578,N_13526);
nor U13825 (N_13825,N_13672,N_13791);
xor U13826 (N_13826,N_13788,N_13580);
and U13827 (N_13827,N_13725,N_13547);
or U13828 (N_13828,N_13745,N_13522);
nand U13829 (N_13829,N_13536,N_13712);
or U13830 (N_13830,N_13641,N_13633);
or U13831 (N_13831,N_13626,N_13557);
nand U13832 (N_13832,N_13700,N_13603);
and U13833 (N_13833,N_13748,N_13648);
xnor U13834 (N_13834,N_13705,N_13692);
nor U13835 (N_13835,N_13616,N_13606);
xor U13836 (N_13836,N_13740,N_13519);
and U13837 (N_13837,N_13713,N_13796);
nand U13838 (N_13838,N_13634,N_13535);
nand U13839 (N_13839,N_13704,N_13584);
nand U13840 (N_13840,N_13504,N_13781);
and U13841 (N_13841,N_13708,N_13714);
nand U13842 (N_13842,N_13577,N_13777);
nor U13843 (N_13843,N_13518,N_13731);
xor U13844 (N_13844,N_13632,N_13715);
or U13845 (N_13845,N_13582,N_13509);
or U13846 (N_13846,N_13520,N_13627);
nand U13847 (N_13847,N_13651,N_13597);
xor U13848 (N_13848,N_13511,N_13538);
xor U13849 (N_13849,N_13596,N_13677);
nor U13850 (N_13850,N_13783,N_13546);
nand U13851 (N_13851,N_13595,N_13515);
nor U13852 (N_13852,N_13779,N_13561);
and U13853 (N_13853,N_13690,N_13707);
xnor U13854 (N_13854,N_13719,N_13687);
nor U13855 (N_13855,N_13757,N_13541);
xor U13856 (N_13856,N_13774,N_13734);
and U13857 (N_13857,N_13680,N_13507);
nor U13858 (N_13858,N_13591,N_13589);
or U13859 (N_13859,N_13587,N_13768);
nor U13860 (N_13860,N_13542,N_13503);
and U13861 (N_13861,N_13717,N_13602);
nand U13862 (N_13862,N_13698,N_13752);
and U13863 (N_13863,N_13759,N_13665);
nand U13864 (N_13864,N_13607,N_13505);
nor U13865 (N_13865,N_13684,N_13555);
or U13866 (N_13866,N_13789,N_13539);
or U13867 (N_13867,N_13583,N_13727);
xnor U13868 (N_13868,N_13750,N_13531);
or U13869 (N_13869,N_13795,N_13610);
nand U13870 (N_13870,N_13529,N_13722);
xor U13871 (N_13871,N_13776,N_13623);
and U13872 (N_13872,N_13767,N_13649);
nand U13873 (N_13873,N_13512,N_13568);
or U13874 (N_13874,N_13537,N_13797);
xnor U13875 (N_13875,N_13576,N_13585);
nand U13876 (N_13876,N_13612,N_13736);
nand U13877 (N_13877,N_13703,N_13760);
or U13878 (N_13878,N_13543,N_13617);
or U13879 (N_13879,N_13738,N_13644);
nor U13880 (N_13880,N_13513,N_13741);
and U13881 (N_13881,N_13658,N_13746);
nor U13882 (N_13882,N_13681,N_13588);
or U13883 (N_13883,N_13699,N_13514);
nor U13884 (N_13884,N_13566,N_13572);
nor U13885 (N_13885,N_13544,N_13659);
and U13886 (N_13886,N_13730,N_13747);
nand U13887 (N_13887,N_13737,N_13500);
nand U13888 (N_13888,N_13706,N_13593);
nand U13889 (N_13889,N_13663,N_13581);
nor U13890 (N_13890,N_13533,N_13711);
xor U13891 (N_13891,N_13770,N_13653);
or U13892 (N_13892,N_13693,N_13669);
and U13893 (N_13893,N_13550,N_13785);
or U13894 (N_13894,N_13749,N_13732);
nand U13895 (N_13895,N_13598,N_13769);
and U13896 (N_13896,N_13563,N_13635);
or U13897 (N_13897,N_13686,N_13564);
or U13898 (N_13898,N_13729,N_13530);
or U13899 (N_13899,N_13524,N_13683);
and U13900 (N_13900,N_13646,N_13671);
nor U13901 (N_13901,N_13689,N_13650);
xor U13902 (N_13902,N_13756,N_13764);
or U13903 (N_13903,N_13798,N_13685);
nand U13904 (N_13904,N_13691,N_13780);
nand U13905 (N_13905,N_13558,N_13710);
nand U13906 (N_13906,N_13622,N_13510);
and U13907 (N_13907,N_13516,N_13755);
or U13908 (N_13908,N_13678,N_13615);
and U13909 (N_13909,N_13701,N_13590);
nand U13910 (N_13910,N_13523,N_13742);
nor U13911 (N_13911,N_13621,N_13766);
and U13912 (N_13912,N_13527,N_13718);
xor U13913 (N_13913,N_13794,N_13608);
or U13914 (N_13914,N_13762,N_13532);
and U13915 (N_13915,N_13574,N_13643);
and U13916 (N_13916,N_13625,N_13501);
nand U13917 (N_13917,N_13661,N_13549);
and U13918 (N_13918,N_13624,N_13548);
or U13919 (N_13919,N_13502,N_13790);
xor U13920 (N_13920,N_13772,N_13614);
or U13921 (N_13921,N_13667,N_13552);
and U13922 (N_13922,N_13696,N_13668);
nand U13923 (N_13923,N_13716,N_13642);
nor U13924 (N_13924,N_13545,N_13709);
nand U13925 (N_13925,N_13571,N_13586);
and U13926 (N_13926,N_13554,N_13567);
nor U13927 (N_13927,N_13506,N_13559);
nand U13928 (N_13928,N_13636,N_13761);
and U13929 (N_13929,N_13562,N_13673);
nor U13930 (N_13930,N_13786,N_13664);
nand U13931 (N_13931,N_13784,N_13528);
or U13932 (N_13932,N_13723,N_13654);
or U13933 (N_13933,N_13782,N_13613);
or U13934 (N_13934,N_13702,N_13743);
xor U13935 (N_13935,N_13551,N_13739);
xnor U13936 (N_13936,N_13656,N_13592);
nor U13937 (N_13937,N_13778,N_13599);
nor U13938 (N_13938,N_13670,N_13631);
or U13939 (N_13939,N_13676,N_13575);
nor U13940 (N_13940,N_13697,N_13560);
nor U13941 (N_13941,N_13688,N_13594);
nor U13942 (N_13942,N_13609,N_13611);
or U13943 (N_13943,N_13569,N_13792);
nor U13944 (N_13944,N_13735,N_13660);
or U13945 (N_13945,N_13657,N_13620);
xnor U13946 (N_13946,N_13638,N_13604);
or U13947 (N_13947,N_13521,N_13763);
nor U13948 (N_13948,N_13775,N_13628);
or U13949 (N_13949,N_13728,N_13517);
nor U13950 (N_13950,N_13696,N_13735);
nor U13951 (N_13951,N_13609,N_13533);
xnor U13952 (N_13952,N_13511,N_13584);
nand U13953 (N_13953,N_13734,N_13758);
nor U13954 (N_13954,N_13612,N_13658);
or U13955 (N_13955,N_13538,N_13642);
nand U13956 (N_13956,N_13625,N_13524);
nor U13957 (N_13957,N_13621,N_13730);
nor U13958 (N_13958,N_13643,N_13787);
nand U13959 (N_13959,N_13762,N_13761);
nor U13960 (N_13960,N_13638,N_13615);
nand U13961 (N_13961,N_13561,N_13674);
and U13962 (N_13962,N_13778,N_13666);
nor U13963 (N_13963,N_13683,N_13646);
xor U13964 (N_13964,N_13634,N_13505);
or U13965 (N_13965,N_13716,N_13507);
nor U13966 (N_13966,N_13746,N_13598);
xnor U13967 (N_13967,N_13566,N_13616);
xnor U13968 (N_13968,N_13655,N_13779);
nor U13969 (N_13969,N_13668,N_13658);
or U13970 (N_13970,N_13545,N_13558);
nand U13971 (N_13971,N_13545,N_13536);
or U13972 (N_13972,N_13763,N_13609);
nor U13973 (N_13973,N_13795,N_13500);
and U13974 (N_13974,N_13694,N_13701);
xor U13975 (N_13975,N_13748,N_13782);
and U13976 (N_13976,N_13729,N_13733);
or U13977 (N_13977,N_13799,N_13636);
or U13978 (N_13978,N_13530,N_13777);
nand U13979 (N_13979,N_13748,N_13545);
or U13980 (N_13980,N_13781,N_13746);
xnor U13981 (N_13981,N_13514,N_13638);
or U13982 (N_13982,N_13772,N_13598);
or U13983 (N_13983,N_13696,N_13750);
nor U13984 (N_13984,N_13788,N_13670);
xnor U13985 (N_13985,N_13745,N_13642);
and U13986 (N_13986,N_13756,N_13606);
nor U13987 (N_13987,N_13664,N_13731);
nand U13988 (N_13988,N_13731,N_13665);
xor U13989 (N_13989,N_13729,N_13627);
and U13990 (N_13990,N_13702,N_13583);
or U13991 (N_13991,N_13628,N_13778);
nand U13992 (N_13992,N_13545,N_13664);
and U13993 (N_13993,N_13569,N_13756);
xor U13994 (N_13994,N_13527,N_13795);
xnor U13995 (N_13995,N_13665,N_13765);
and U13996 (N_13996,N_13736,N_13575);
xnor U13997 (N_13997,N_13756,N_13597);
or U13998 (N_13998,N_13601,N_13684);
nand U13999 (N_13999,N_13778,N_13563);
or U14000 (N_14000,N_13696,N_13595);
and U14001 (N_14001,N_13541,N_13574);
and U14002 (N_14002,N_13513,N_13505);
xor U14003 (N_14003,N_13781,N_13598);
or U14004 (N_14004,N_13557,N_13777);
nand U14005 (N_14005,N_13749,N_13506);
and U14006 (N_14006,N_13586,N_13752);
xnor U14007 (N_14007,N_13799,N_13572);
and U14008 (N_14008,N_13616,N_13713);
nor U14009 (N_14009,N_13660,N_13500);
nand U14010 (N_14010,N_13699,N_13744);
nand U14011 (N_14011,N_13788,N_13724);
xnor U14012 (N_14012,N_13692,N_13647);
or U14013 (N_14013,N_13770,N_13758);
and U14014 (N_14014,N_13528,N_13701);
or U14015 (N_14015,N_13654,N_13658);
xnor U14016 (N_14016,N_13775,N_13691);
and U14017 (N_14017,N_13586,N_13657);
nor U14018 (N_14018,N_13714,N_13553);
and U14019 (N_14019,N_13775,N_13759);
and U14020 (N_14020,N_13547,N_13624);
nor U14021 (N_14021,N_13690,N_13537);
nor U14022 (N_14022,N_13649,N_13605);
and U14023 (N_14023,N_13634,N_13765);
nand U14024 (N_14024,N_13574,N_13775);
nand U14025 (N_14025,N_13701,N_13671);
nand U14026 (N_14026,N_13577,N_13795);
or U14027 (N_14027,N_13635,N_13572);
and U14028 (N_14028,N_13560,N_13685);
nand U14029 (N_14029,N_13713,N_13795);
nand U14030 (N_14030,N_13743,N_13681);
xnor U14031 (N_14031,N_13651,N_13666);
xnor U14032 (N_14032,N_13590,N_13502);
or U14033 (N_14033,N_13644,N_13580);
or U14034 (N_14034,N_13601,N_13750);
nand U14035 (N_14035,N_13778,N_13567);
and U14036 (N_14036,N_13540,N_13630);
xnor U14037 (N_14037,N_13563,N_13774);
nor U14038 (N_14038,N_13543,N_13696);
or U14039 (N_14039,N_13672,N_13560);
or U14040 (N_14040,N_13521,N_13707);
and U14041 (N_14041,N_13615,N_13750);
nor U14042 (N_14042,N_13618,N_13766);
nor U14043 (N_14043,N_13542,N_13790);
and U14044 (N_14044,N_13753,N_13565);
or U14045 (N_14045,N_13621,N_13718);
nor U14046 (N_14046,N_13703,N_13704);
nand U14047 (N_14047,N_13780,N_13500);
and U14048 (N_14048,N_13562,N_13527);
nor U14049 (N_14049,N_13574,N_13735);
nor U14050 (N_14050,N_13774,N_13521);
nand U14051 (N_14051,N_13759,N_13754);
or U14052 (N_14052,N_13700,N_13584);
nand U14053 (N_14053,N_13650,N_13612);
and U14054 (N_14054,N_13593,N_13633);
or U14055 (N_14055,N_13714,N_13616);
nor U14056 (N_14056,N_13678,N_13793);
nor U14057 (N_14057,N_13599,N_13795);
nor U14058 (N_14058,N_13648,N_13777);
and U14059 (N_14059,N_13670,N_13619);
or U14060 (N_14060,N_13539,N_13639);
nand U14061 (N_14061,N_13603,N_13500);
and U14062 (N_14062,N_13630,N_13674);
nand U14063 (N_14063,N_13629,N_13785);
and U14064 (N_14064,N_13543,N_13654);
and U14065 (N_14065,N_13643,N_13619);
xor U14066 (N_14066,N_13699,N_13697);
nand U14067 (N_14067,N_13560,N_13637);
xnor U14068 (N_14068,N_13578,N_13701);
nand U14069 (N_14069,N_13770,N_13775);
or U14070 (N_14070,N_13501,N_13615);
nor U14071 (N_14071,N_13750,N_13598);
and U14072 (N_14072,N_13738,N_13795);
or U14073 (N_14073,N_13536,N_13546);
xnor U14074 (N_14074,N_13623,N_13794);
xor U14075 (N_14075,N_13733,N_13513);
nor U14076 (N_14076,N_13755,N_13620);
nand U14077 (N_14077,N_13622,N_13667);
or U14078 (N_14078,N_13607,N_13651);
or U14079 (N_14079,N_13695,N_13642);
and U14080 (N_14080,N_13746,N_13626);
nand U14081 (N_14081,N_13518,N_13644);
xnor U14082 (N_14082,N_13750,N_13674);
xor U14083 (N_14083,N_13600,N_13509);
xor U14084 (N_14084,N_13645,N_13755);
or U14085 (N_14085,N_13641,N_13756);
xor U14086 (N_14086,N_13643,N_13559);
and U14087 (N_14087,N_13769,N_13786);
nand U14088 (N_14088,N_13729,N_13798);
nand U14089 (N_14089,N_13540,N_13795);
or U14090 (N_14090,N_13519,N_13524);
nor U14091 (N_14091,N_13561,N_13575);
xor U14092 (N_14092,N_13518,N_13714);
xnor U14093 (N_14093,N_13588,N_13759);
nand U14094 (N_14094,N_13508,N_13577);
and U14095 (N_14095,N_13629,N_13740);
nand U14096 (N_14096,N_13505,N_13604);
nor U14097 (N_14097,N_13516,N_13572);
nand U14098 (N_14098,N_13717,N_13734);
and U14099 (N_14099,N_13523,N_13569);
and U14100 (N_14100,N_13983,N_13828);
nor U14101 (N_14101,N_14011,N_13944);
and U14102 (N_14102,N_13973,N_13960);
nor U14103 (N_14103,N_13803,N_13914);
or U14104 (N_14104,N_14054,N_13845);
or U14105 (N_14105,N_14076,N_13825);
and U14106 (N_14106,N_13815,N_14010);
nor U14107 (N_14107,N_14007,N_14087);
and U14108 (N_14108,N_14014,N_14037);
nor U14109 (N_14109,N_13835,N_13996);
and U14110 (N_14110,N_14071,N_13924);
and U14111 (N_14111,N_14079,N_14040);
nand U14112 (N_14112,N_14053,N_14000);
xor U14113 (N_14113,N_14051,N_13904);
nand U14114 (N_14114,N_13892,N_13978);
xnor U14115 (N_14115,N_14091,N_14018);
and U14116 (N_14116,N_14047,N_13863);
or U14117 (N_14117,N_13875,N_13839);
nand U14118 (N_14118,N_13947,N_13844);
or U14119 (N_14119,N_14034,N_13966);
xor U14120 (N_14120,N_14059,N_13956);
xnor U14121 (N_14121,N_13855,N_13985);
or U14122 (N_14122,N_14032,N_13981);
nor U14123 (N_14123,N_13880,N_13932);
or U14124 (N_14124,N_13993,N_13943);
or U14125 (N_14125,N_14046,N_13840);
nand U14126 (N_14126,N_13938,N_14070);
or U14127 (N_14127,N_13858,N_13823);
and U14128 (N_14128,N_14005,N_14050);
or U14129 (N_14129,N_13816,N_13910);
xor U14130 (N_14130,N_14089,N_14001);
and U14131 (N_14131,N_14081,N_14073);
nand U14132 (N_14132,N_13917,N_14082);
and U14133 (N_14133,N_13967,N_13899);
xor U14134 (N_14134,N_13908,N_14092);
and U14135 (N_14135,N_14023,N_13998);
nand U14136 (N_14136,N_13830,N_13814);
xnor U14137 (N_14137,N_14038,N_13991);
and U14138 (N_14138,N_13989,N_13826);
or U14139 (N_14139,N_13953,N_14086);
and U14140 (N_14140,N_13842,N_13854);
nor U14141 (N_14141,N_13866,N_13832);
or U14142 (N_14142,N_13974,N_13911);
nand U14143 (N_14143,N_14002,N_13820);
and U14144 (N_14144,N_14075,N_13879);
nand U14145 (N_14145,N_13817,N_14026);
xnor U14146 (N_14146,N_13902,N_13884);
nand U14147 (N_14147,N_13941,N_13894);
nand U14148 (N_14148,N_14080,N_14063);
and U14149 (N_14149,N_14028,N_13923);
xor U14150 (N_14150,N_13852,N_14004);
and U14151 (N_14151,N_14020,N_13957);
nor U14152 (N_14152,N_13994,N_13963);
xnor U14153 (N_14153,N_13909,N_13882);
xor U14154 (N_14154,N_14088,N_14043);
and U14155 (N_14155,N_13968,N_14098);
or U14156 (N_14156,N_13986,N_13896);
and U14157 (N_14157,N_13868,N_14009);
and U14158 (N_14158,N_14024,N_14083);
xnor U14159 (N_14159,N_14056,N_13915);
nand U14160 (N_14160,N_13903,N_14006);
or U14161 (N_14161,N_13897,N_14003);
nand U14162 (N_14162,N_13999,N_14008);
xnor U14163 (N_14163,N_13888,N_13841);
or U14164 (N_14164,N_14029,N_13886);
and U14165 (N_14165,N_14042,N_13873);
nor U14166 (N_14166,N_13802,N_13819);
nand U14167 (N_14167,N_14044,N_13821);
nand U14168 (N_14168,N_14061,N_13933);
nor U14169 (N_14169,N_13808,N_14093);
nand U14170 (N_14170,N_14074,N_14019);
nor U14171 (N_14171,N_13849,N_13810);
nand U14172 (N_14172,N_14078,N_13846);
or U14173 (N_14173,N_13838,N_13950);
and U14174 (N_14174,N_13876,N_14096);
and U14175 (N_14175,N_13976,N_13959);
or U14176 (N_14176,N_14099,N_13881);
or U14177 (N_14177,N_13889,N_13955);
and U14178 (N_14178,N_13864,N_13848);
and U14179 (N_14179,N_13964,N_13927);
nand U14180 (N_14180,N_14031,N_13946);
nor U14181 (N_14181,N_14052,N_14017);
and U14182 (N_14182,N_14033,N_13861);
xor U14183 (N_14183,N_14057,N_14016);
nand U14184 (N_14184,N_14066,N_13806);
xor U14185 (N_14185,N_13949,N_13857);
xnor U14186 (N_14186,N_14067,N_14041);
nand U14187 (N_14187,N_14094,N_13916);
xnor U14188 (N_14188,N_13977,N_13988);
or U14189 (N_14189,N_13809,N_13940);
xnor U14190 (N_14190,N_14039,N_13860);
nor U14191 (N_14191,N_13979,N_14048);
nand U14192 (N_14192,N_13928,N_13834);
nand U14193 (N_14193,N_13948,N_13906);
or U14194 (N_14194,N_13905,N_13813);
nand U14195 (N_14195,N_13952,N_13939);
xor U14196 (N_14196,N_13995,N_13871);
nand U14197 (N_14197,N_14022,N_13887);
nand U14198 (N_14198,N_14065,N_13827);
nand U14199 (N_14199,N_13992,N_13867);
and U14200 (N_14200,N_13931,N_13912);
nand U14201 (N_14201,N_13865,N_13800);
xor U14202 (N_14202,N_13937,N_13878);
or U14203 (N_14203,N_14013,N_14064);
xor U14204 (N_14204,N_13870,N_13850);
or U14205 (N_14205,N_13843,N_13811);
xnor U14206 (N_14206,N_13930,N_14025);
and U14207 (N_14207,N_14085,N_13975);
nor U14208 (N_14208,N_14049,N_13874);
nor U14209 (N_14209,N_13862,N_13972);
nand U14210 (N_14210,N_13851,N_14060);
nor U14211 (N_14211,N_13807,N_13824);
or U14212 (N_14212,N_13869,N_13970);
nor U14213 (N_14213,N_13837,N_13969);
xnor U14214 (N_14214,N_13890,N_14058);
and U14215 (N_14215,N_13804,N_14068);
nand U14216 (N_14216,N_13859,N_13929);
nand U14217 (N_14217,N_13812,N_13918);
or U14218 (N_14218,N_14077,N_13990);
or U14219 (N_14219,N_14030,N_14072);
or U14220 (N_14220,N_13965,N_13958);
nand U14221 (N_14221,N_13907,N_14012);
or U14222 (N_14222,N_13984,N_14090);
and U14223 (N_14223,N_13997,N_13898);
nand U14224 (N_14224,N_13836,N_13853);
or U14225 (N_14225,N_13801,N_13919);
or U14226 (N_14226,N_13962,N_13926);
nand U14227 (N_14227,N_14062,N_13900);
or U14228 (N_14228,N_13891,N_13942);
and U14229 (N_14229,N_13934,N_13833);
xor U14230 (N_14230,N_13831,N_13877);
xor U14231 (N_14231,N_13954,N_14055);
or U14232 (N_14232,N_13847,N_13922);
and U14233 (N_14233,N_13971,N_13818);
nand U14234 (N_14234,N_13822,N_13829);
xnor U14235 (N_14235,N_14036,N_13872);
and U14236 (N_14236,N_13925,N_13895);
or U14237 (N_14237,N_13885,N_13945);
nand U14238 (N_14238,N_13935,N_14045);
xnor U14239 (N_14239,N_13982,N_14027);
and U14240 (N_14240,N_14097,N_13961);
nand U14241 (N_14241,N_13980,N_13921);
xnor U14242 (N_14242,N_13987,N_13856);
nor U14243 (N_14243,N_13920,N_13913);
nand U14244 (N_14244,N_14095,N_14069);
nand U14245 (N_14245,N_13901,N_14035);
nor U14246 (N_14246,N_13883,N_14021);
nor U14247 (N_14247,N_13893,N_14084);
nor U14248 (N_14248,N_13805,N_14015);
nor U14249 (N_14249,N_13936,N_13951);
or U14250 (N_14250,N_14042,N_14036);
nor U14251 (N_14251,N_14037,N_13820);
or U14252 (N_14252,N_14019,N_14078);
nand U14253 (N_14253,N_14031,N_13933);
nor U14254 (N_14254,N_13847,N_13986);
nand U14255 (N_14255,N_13937,N_13832);
nor U14256 (N_14256,N_13899,N_13986);
xor U14257 (N_14257,N_13918,N_13894);
and U14258 (N_14258,N_14014,N_13956);
nor U14259 (N_14259,N_14025,N_14035);
or U14260 (N_14260,N_13946,N_13872);
nor U14261 (N_14261,N_13991,N_13970);
xnor U14262 (N_14262,N_13856,N_14034);
or U14263 (N_14263,N_13813,N_13972);
nor U14264 (N_14264,N_13817,N_14060);
or U14265 (N_14265,N_14011,N_13895);
or U14266 (N_14266,N_14080,N_13993);
nand U14267 (N_14267,N_14025,N_13981);
nand U14268 (N_14268,N_14062,N_14090);
nor U14269 (N_14269,N_14056,N_13806);
nand U14270 (N_14270,N_14053,N_13852);
xnor U14271 (N_14271,N_13934,N_14040);
xnor U14272 (N_14272,N_14090,N_14098);
nand U14273 (N_14273,N_13983,N_13893);
nor U14274 (N_14274,N_13901,N_13822);
nor U14275 (N_14275,N_14008,N_13983);
and U14276 (N_14276,N_14049,N_13911);
nand U14277 (N_14277,N_14021,N_14095);
nand U14278 (N_14278,N_14057,N_14083);
and U14279 (N_14279,N_13946,N_13961);
nand U14280 (N_14280,N_13932,N_13965);
xor U14281 (N_14281,N_13838,N_13897);
nor U14282 (N_14282,N_13830,N_13953);
nor U14283 (N_14283,N_13984,N_13907);
nand U14284 (N_14284,N_14007,N_13862);
nand U14285 (N_14285,N_13996,N_13861);
xor U14286 (N_14286,N_14018,N_13989);
nand U14287 (N_14287,N_13902,N_13976);
nand U14288 (N_14288,N_14031,N_13822);
and U14289 (N_14289,N_13975,N_14001);
or U14290 (N_14290,N_14018,N_13865);
or U14291 (N_14291,N_13986,N_14026);
nor U14292 (N_14292,N_13926,N_13964);
nand U14293 (N_14293,N_14060,N_14078);
and U14294 (N_14294,N_13967,N_13869);
nor U14295 (N_14295,N_13877,N_13878);
xnor U14296 (N_14296,N_13868,N_13860);
xnor U14297 (N_14297,N_13946,N_13812);
xor U14298 (N_14298,N_13919,N_14007);
nor U14299 (N_14299,N_14030,N_14086);
nor U14300 (N_14300,N_13944,N_14065);
or U14301 (N_14301,N_13822,N_13879);
or U14302 (N_14302,N_13933,N_13837);
nand U14303 (N_14303,N_13896,N_13940);
nand U14304 (N_14304,N_14024,N_14081);
nand U14305 (N_14305,N_13835,N_14022);
or U14306 (N_14306,N_13805,N_14060);
and U14307 (N_14307,N_13807,N_13990);
xor U14308 (N_14308,N_14006,N_14045);
xor U14309 (N_14309,N_13880,N_14088);
xnor U14310 (N_14310,N_13943,N_14024);
xnor U14311 (N_14311,N_14024,N_13898);
nand U14312 (N_14312,N_13881,N_13805);
nand U14313 (N_14313,N_13852,N_13808);
xor U14314 (N_14314,N_13903,N_14033);
nor U14315 (N_14315,N_14051,N_14096);
and U14316 (N_14316,N_14090,N_14060);
and U14317 (N_14317,N_13978,N_13882);
nor U14318 (N_14318,N_14031,N_14058);
xnor U14319 (N_14319,N_14083,N_14054);
or U14320 (N_14320,N_13982,N_13966);
or U14321 (N_14321,N_14082,N_14046);
nor U14322 (N_14322,N_13945,N_13951);
and U14323 (N_14323,N_13969,N_13904);
nor U14324 (N_14324,N_13855,N_13872);
nor U14325 (N_14325,N_13865,N_13962);
and U14326 (N_14326,N_13987,N_13868);
nor U14327 (N_14327,N_13986,N_13982);
or U14328 (N_14328,N_14066,N_13823);
xor U14329 (N_14329,N_14029,N_14091);
nor U14330 (N_14330,N_13868,N_13880);
nand U14331 (N_14331,N_13919,N_14074);
and U14332 (N_14332,N_14080,N_13889);
nand U14333 (N_14333,N_14069,N_13912);
nor U14334 (N_14334,N_13986,N_13924);
nand U14335 (N_14335,N_13814,N_14094);
nor U14336 (N_14336,N_13971,N_14063);
or U14337 (N_14337,N_14023,N_14068);
nand U14338 (N_14338,N_13850,N_13841);
or U14339 (N_14339,N_14065,N_13856);
nor U14340 (N_14340,N_14085,N_13951);
nand U14341 (N_14341,N_14058,N_14044);
nand U14342 (N_14342,N_13861,N_14053);
nor U14343 (N_14343,N_13993,N_13885);
and U14344 (N_14344,N_13862,N_13836);
xor U14345 (N_14345,N_13861,N_14047);
nand U14346 (N_14346,N_13984,N_13880);
xor U14347 (N_14347,N_13850,N_13899);
nand U14348 (N_14348,N_13808,N_14003);
or U14349 (N_14349,N_13814,N_13801);
xnor U14350 (N_14350,N_13854,N_14006);
or U14351 (N_14351,N_13957,N_14059);
xor U14352 (N_14352,N_13822,N_13881);
and U14353 (N_14353,N_13853,N_13832);
and U14354 (N_14354,N_14027,N_13991);
and U14355 (N_14355,N_14033,N_13811);
xor U14356 (N_14356,N_13905,N_14083);
nand U14357 (N_14357,N_13975,N_13806);
nand U14358 (N_14358,N_13824,N_13801);
nand U14359 (N_14359,N_14062,N_14097);
and U14360 (N_14360,N_13805,N_14076);
nand U14361 (N_14361,N_14081,N_13976);
nor U14362 (N_14362,N_13870,N_13862);
nand U14363 (N_14363,N_13880,N_13843);
and U14364 (N_14364,N_13941,N_14097);
or U14365 (N_14365,N_13835,N_13913);
and U14366 (N_14366,N_13994,N_14092);
xnor U14367 (N_14367,N_13905,N_13975);
and U14368 (N_14368,N_13992,N_13962);
or U14369 (N_14369,N_13885,N_13997);
xnor U14370 (N_14370,N_13922,N_13830);
xnor U14371 (N_14371,N_13825,N_14047);
xor U14372 (N_14372,N_14028,N_14068);
and U14373 (N_14373,N_14048,N_13853);
nand U14374 (N_14374,N_13997,N_14080);
nor U14375 (N_14375,N_13830,N_13871);
or U14376 (N_14376,N_14078,N_13814);
xnor U14377 (N_14377,N_13800,N_13977);
or U14378 (N_14378,N_13944,N_14066);
or U14379 (N_14379,N_13930,N_14033);
and U14380 (N_14380,N_14019,N_13859);
xnor U14381 (N_14381,N_13976,N_14056);
or U14382 (N_14382,N_13853,N_14091);
nand U14383 (N_14383,N_13978,N_13951);
xor U14384 (N_14384,N_14090,N_13972);
nand U14385 (N_14385,N_13919,N_13961);
nor U14386 (N_14386,N_13947,N_14041);
nor U14387 (N_14387,N_13935,N_14095);
xnor U14388 (N_14388,N_13825,N_13981);
nand U14389 (N_14389,N_13868,N_13878);
and U14390 (N_14390,N_13826,N_14025);
nor U14391 (N_14391,N_14045,N_14062);
xnor U14392 (N_14392,N_13922,N_14022);
nor U14393 (N_14393,N_13854,N_13832);
and U14394 (N_14394,N_13816,N_14021);
and U14395 (N_14395,N_13933,N_13975);
nor U14396 (N_14396,N_14022,N_14064);
and U14397 (N_14397,N_13847,N_14065);
xor U14398 (N_14398,N_14016,N_13960);
nor U14399 (N_14399,N_13855,N_14082);
nor U14400 (N_14400,N_14359,N_14286);
and U14401 (N_14401,N_14235,N_14113);
nor U14402 (N_14402,N_14250,N_14285);
nor U14403 (N_14403,N_14238,N_14344);
xnor U14404 (N_14404,N_14107,N_14193);
xnor U14405 (N_14405,N_14117,N_14348);
and U14406 (N_14406,N_14248,N_14307);
nor U14407 (N_14407,N_14383,N_14204);
nand U14408 (N_14408,N_14183,N_14349);
xor U14409 (N_14409,N_14379,N_14340);
and U14410 (N_14410,N_14257,N_14280);
and U14411 (N_14411,N_14227,N_14291);
nand U14412 (N_14412,N_14370,N_14276);
or U14413 (N_14413,N_14306,N_14269);
xor U14414 (N_14414,N_14211,N_14317);
nor U14415 (N_14415,N_14293,N_14315);
nor U14416 (N_14416,N_14328,N_14392);
and U14417 (N_14417,N_14199,N_14234);
or U14418 (N_14418,N_14282,N_14301);
xnor U14419 (N_14419,N_14223,N_14166);
nor U14420 (N_14420,N_14397,N_14380);
nand U14421 (N_14421,N_14270,N_14311);
xor U14422 (N_14422,N_14313,N_14220);
xnor U14423 (N_14423,N_14110,N_14396);
and U14424 (N_14424,N_14164,N_14346);
and U14425 (N_14425,N_14224,N_14333);
or U14426 (N_14426,N_14351,N_14368);
xnor U14427 (N_14427,N_14100,N_14316);
xnor U14428 (N_14428,N_14385,N_14127);
nand U14429 (N_14429,N_14165,N_14241);
and U14430 (N_14430,N_14387,N_14366);
xnor U14431 (N_14431,N_14126,N_14135);
xnor U14432 (N_14432,N_14145,N_14207);
nor U14433 (N_14433,N_14255,N_14354);
nor U14434 (N_14434,N_14124,N_14300);
nor U14435 (N_14435,N_14137,N_14203);
nor U14436 (N_14436,N_14281,N_14324);
xnor U14437 (N_14437,N_14148,N_14146);
xnor U14438 (N_14438,N_14198,N_14367);
and U14439 (N_14439,N_14294,N_14239);
nor U14440 (N_14440,N_14159,N_14130);
xor U14441 (N_14441,N_14221,N_14369);
nor U14442 (N_14442,N_14103,N_14247);
nor U14443 (N_14443,N_14395,N_14140);
nor U14444 (N_14444,N_14261,N_14236);
and U14445 (N_14445,N_14125,N_14149);
nor U14446 (N_14446,N_14266,N_14195);
nand U14447 (N_14447,N_14178,N_14129);
nor U14448 (N_14448,N_14288,N_14357);
or U14449 (N_14449,N_14230,N_14295);
or U14450 (N_14450,N_14121,N_14296);
and U14451 (N_14451,N_14258,N_14399);
xor U14452 (N_14452,N_14142,N_14310);
xor U14453 (N_14453,N_14190,N_14196);
and U14454 (N_14454,N_14303,N_14168);
and U14455 (N_14455,N_14342,N_14150);
nor U14456 (N_14456,N_14205,N_14156);
nor U14457 (N_14457,N_14133,N_14364);
or U14458 (N_14458,N_14228,N_14181);
or U14459 (N_14459,N_14352,N_14343);
xor U14460 (N_14460,N_14138,N_14173);
nor U14461 (N_14461,N_14358,N_14186);
nor U14462 (N_14462,N_14171,N_14355);
nor U14463 (N_14463,N_14332,N_14376);
nor U14464 (N_14464,N_14308,N_14284);
xor U14465 (N_14465,N_14322,N_14118);
nand U14466 (N_14466,N_14305,N_14120);
or U14467 (N_14467,N_14243,N_14330);
xor U14468 (N_14468,N_14363,N_14297);
xor U14469 (N_14469,N_14252,N_14391);
or U14470 (N_14470,N_14231,N_14112);
nor U14471 (N_14471,N_14189,N_14350);
nand U14472 (N_14472,N_14323,N_14217);
and U14473 (N_14473,N_14214,N_14141);
nand U14474 (N_14474,N_14304,N_14256);
or U14475 (N_14475,N_14105,N_14263);
nand U14476 (N_14476,N_14184,N_14101);
xnor U14477 (N_14477,N_14382,N_14329);
and U14478 (N_14478,N_14208,N_14191);
nor U14479 (N_14479,N_14160,N_14260);
and U14480 (N_14480,N_14331,N_14188);
and U14481 (N_14481,N_14381,N_14389);
and U14482 (N_14482,N_14213,N_14378);
nor U14483 (N_14483,N_14264,N_14232);
nand U14484 (N_14484,N_14157,N_14242);
xor U14485 (N_14485,N_14334,N_14174);
nand U14486 (N_14486,N_14271,N_14273);
nand U14487 (N_14487,N_14390,N_14128);
xnor U14488 (N_14488,N_14201,N_14233);
nor U14489 (N_14489,N_14339,N_14102);
nand U14490 (N_14490,N_14123,N_14345);
xor U14491 (N_14491,N_14163,N_14254);
and U14492 (N_14492,N_14287,N_14229);
nand U14493 (N_14493,N_14104,N_14283);
nand U14494 (N_14494,N_14398,N_14167);
nor U14495 (N_14495,N_14175,N_14136);
or U14496 (N_14496,N_14319,N_14290);
nor U14497 (N_14497,N_14251,N_14371);
nand U14498 (N_14498,N_14321,N_14298);
and U14499 (N_14499,N_14259,N_14360);
nor U14500 (N_14500,N_14362,N_14206);
nand U14501 (N_14501,N_14212,N_14356);
nor U14502 (N_14502,N_14347,N_14218);
xnor U14503 (N_14503,N_14202,N_14240);
or U14504 (N_14504,N_14265,N_14249);
xnor U14505 (N_14505,N_14336,N_14116);
xor U14506 (N_14506,N_14237,N_14377);
and U14507 (N_14507,N_14161,N_14226);
nand U14508 (N_14508,N_14361,N_14268);
xnor U14509 (N_14509,N_14162,N_14335);
xnor U14510 (N_14510,N_14109,N_14327);
or U14511 (N_14511,N_14172,N_14375);
nand U14512 (N_14512,N_14155,N_14216);
xor U14513 (N_14513,N_14169,N_14292);
and U14514 (N_14514,N_14219,N_14253);
or U14515 (N_14515,N_14122,N_14210);
or U14516 (N_14516,N_14179,N_14151);
or U14517 (N_14517,N_14115,N_14374);
or U14518 (N_14518,N_14274,N_14108);
xor U14519 (N_14519,N_14318,N_14338);
and U14520 (N_14520,N_14353,N_14388);
nor U14521 (N_14521,N_14180,N_14277);
xor U14522 (N_14522,N_14225,N_14114);
or U14523 (N_14523,N_14131,N_14299);
nor U14524 (N_14524,N_14279,N_14170);
nor U14525 (N_14525,N_14209,N_14278);
nand U14526 (N_14526,N_14106,N_14289);
or U14527 (N_14527,N_14177,N_14372);
nand U14528 (N_14528,N_14326,N_14176);
or U14529 (N_14529,N_14309,N_14246);
nand U14530 (N_14530,N_14386,N_14144);
nand U14531 (N_14531,N_14394,N_14215);
and U14532 (N_14532,N_14153,N_14337);
and U14533 (N_14533,N_14245,N_14393);
and U14534 (N_14534,N_14158,N_14132);
nor U14535 (N_14535,N_14314,N_14143);
nor U14536 (N_14536,N_14154,N_14147);
nor U14537 (N_14537,N_14325,N_14244);
nor U14538 (N_14538,N_14267,N_14182);
nand U14539 (N_14539,N_14222,N_14152);
xnor U14540 (N_14540,N_14139,N_14119);
nand U14541 (N_14541,N_14365,N_14384);
and U14542 (N_14542,N_14341,N_14192);
or U14543 (N_14543,N_14275,N_14373);
nor U14544 (N_14544,N_14262,N_14272);
nand U14545 (N_14545,N_14200,N_14312);
or U14546 (N_14546,N_14194,N_14320);
xor U14547 (N_14547,N_14134,N_14185);
xor U14548 (N_14548,N_14187,N_14197);
and U14549 (N_14549,N_14302,N_14111);
nor U14550 (N_14550,N_14217,N_14358);
xor U14551 (N_14551,N_14305,N_14174);
nor U14552 (N_14552,N_14324,N_14119);
and U14553 (N_14553,N_14174,N_14104);
or U14554 (N_14554,N_14198,N_14233);
or U14555 (N_14555,N_14256,N_14254);
or U14556 (N_14556,N_14193,N_14333);
and U14557 (N_14557,N_14339,N_14174);
nand U14558 (N_14558,N_14321,N_14250);
xnor U14559 (N_14559,N_14290,N_14276);
nand U14560 (N_14560,N_14295,N_14335);
nand U14561 (N_14561,N_14248,N_14346);
nor U14562 (N_14562,N_14240,N_14351);
or U14563 (N_14563,N_14311,N_14162);
and U14564 (N_14564,N_14209,N_14143);
and U14565 (N_14565,N_14325,N_14291);
nor U14566 (N_14566,N_14118,N_14127);
xnor U14567 (N_14567,N_14146,N_14344);
and U14568 (N_14568,N_14142,N_14254);
or U14569 (N_14569,N_14264,N_14344);
xor U14570 (N_14570,N_14369,N_14138);
and U14571 (N_14571,N_14201,N_14122);
xnor U14572 (N_14572,N_14253,N_14393);
and U14573 (N_14573,N_14156,N_14289);
nor U14574 (N_14574,N_14245,N_14377);
or U14575 (N_14575,N_14143,N_14104);
or U14576 (N_14576,N_14262,N_14220);
xnor U14577 (N_14577,N_14172,N_14275);
and U14578 (N_14578,N_14165,N_14158);
nand U14579 (N_14579,N_14277,N_14390);
nand U14580 (N_14580,N_14359,N_14200);
and U14581 (N_14581,N_14195,N_14396);
nor U14582 (N_14582,N_14385,N_14341);
nor U14583 (N_14583,N_14309,N_14261);
nor U14584 (N_14584,N_14378,N_14232);
or U14585 (N_14585,N_14166,N_14310);
and U14586 (N_14586,N_14271,N_14175);
xnor U14587 (N_14587,N_14395,N_14361);
nor U14588 (N_14588,N_14194,N_14155);
xor U14589 (N_14589,N_14175,N_14243);
or U14590 (N_14590,N_14220,N_14218);
or U14591 (N_14591,N_14101,N_14171);
nor U14592 (N_14592,N_14106,N_14216);
xnor U14593 (N_14593,N_14205,N_14187);
and U14594 (N_14594,N_14162,N_14319);
xor U14595 (N_14595,N_14114,N_14294);
xor U14596 (N_14596,N_14227,N_14218);
nor U14597 (N_14597,N_14209,N_14181);
or U14598 (N_14598,N_14253,N_14213);
nor U14599 (N_14599,N_14232,N_14394);
xnor U14600 (N_14600,N_14220,N_14288);
or U14601 (N_14601,N_14305,N_14126);
or U14602 (N_14602,N_14114,N_14303);
or U14603 (N_14603,N_14280,N_14374);
nor U14604 (N_14604,N_14238,N_14355);
and U14605 (N_14605,N_14221,N_14346);
nor U14606 (N_14606,N_14330,N_14274);
nor U14607 (N_14607,N_14257,N_14156);
and U14608 (N_14608,N_14386,N_14336);
nor U14609 (N_14609,N_14250,N_14101);
nor U14610 (N_14610,N_14389,N_14114);
xor U14611 (N_14611,N_14347,N_14131);
or U14612 (N_14612,N_14144,N_14138);
nand U14613 (N_14613,N_14374,N_14395);
or U14614 (N_14614,N_14327,N_14126);
nand U14615 (N_14615,N_14335,N_14346);
xnor U14616 (N_14616,N_14102,N_14300);
or U14617 (N_14617,N_14198,N_14338);
nor U14618 (N_14618,N_14337,N_14136);
or U14619 (N_14619,N_14255,N_14256);
and U14620 (N_14620,N_14240,N_14118);
xnor U14621 (N_14621,N_14335,N_14395);
xnor U14622 (N_14622,N_14299,N_14104);
and U14623 (N_14623,N_14149,N_14326);
nor U14624 (N_14624,N_14131,N_14124);
or U14625 (N_14625,N_14249,N_14325);
nor U14626 (N_14626,N_14274,N_14304);
nor U14627 (N_14627,N_14149,N_14107);
xnor U14628 (N_14628,N_14319,N_14146);
xnor U14629 (N_14629,N_14377,N_14316);
xor U14630 (N_14630,N_14152,N_14351);
nor U14631 (N_14631,N_14116,N_14318);
nor U14632 (N_14632,N_14184,N_14379);
nor U14633 (N_14633,N_14261,N_14254);
nor U14634 (N_14634,N_14126,N_14108);
or U14635 (N_14635,N_14367,N_14279);
nor U14636 (N_14636,N_14241,N_14264);
nor U14637 (N_14637,N_14345,N_14375);
or U14638 (N_14638,N_14369,N_14244);
nor U14639 (N_14639,N_14249,N_14396);
nor U14640 (N_14640,N_14167,N_14106);
or U14641 (N_14641,N_14294,N_14159);
nor U14642 (N_14642,N_14185,N_14270);
xnor U14643 (N_14643,N_14300,N_14147);
nand U14644 (N_14644,N_14314,N_14308);
nor U14645 (N_14645,N_14201,N_14136);
and U14646 (N_14646,N_14246,N_14159);
nor U14647 (N_14647,N_14365,N_14143);
nor U14648 (N_14648,N_14325,N_14346);
or U14649 (N_14649,N_14169,N_14364);
nor U14650 (N_14650,N_14386,N_14162);
nor U14651 (N_14651,N_14243,N_14113);
nor U14652 (N_14652,N_14392,N_14176);
and U14653 (N_14653,N_14304,N_14151);
and U14654 (N_14654,N_14211,N_14262);
xnor U14655 (N_14655,N_14251,N_14202);
xnor U14656 (N_14656,N_14248,N_14273);
nand U14657 (N_14657,N_14197,N_14228);
and U14658 (N_14658,N_14329,N_14120);
nor U14659 (N_14659,N_14397,N_14335);
nor U14660 (N_14660,N_14372,N_14340);
and U14661 (N_14661,N_14227,N_14162);
and U14662 (N_14662,N_14388,N_14155);
nand U14663 (N_14663,N_14316,N_14175);
nor U14664 (N_14664,N_14388,N_14292);
and U14665 (N_14665,N_14176,N_14328);
nand U14666 (N_14666,N_14238,N_14322);
nand U14667 (N_14667,N_14264,N_14269);
or U14668 (N_14668,N_14317,N_14229);
and U14669 (N_14669,N_14385,N_14154);
xor U14670 (N_14670,N_14210,N_14348);
xor U14671 (N_14671,N_14340,N_14384);
nand U14672 (N_14672,N_14208,N_14220);
xor U14673 (N_14673,N_14128,N_14219);
and U14674 (N_14674,N_14234,N_14200);
or U14675 (N_14675,N_14246,N_14316);
nand U14676 (N_14676,N_14266,N_14165);
nor U14677 (N_14677,N_14210,N_14175);
nand U14678 (N_14678,N_14249,N_14214);
nor U14679 (N_14679,N_14203,N_14173);
and U14680 (N_14680,N_14284,N_14145);
or U14681 (N_14681,N_14366,N_14122);
nor U14682 (N_14682,N_14220,N_14383);
nand U14683 (N_14683,N_14335,N_14237);
or U14684 (N_14684,N_14183,N_14116);
xnor U14685 (N_14685,N_14324,N_14329);
xnor U14686 (N_14686,N_14367,N_14225);
nand U14687 (N_14687,N_14329,N_14212);
nor U14688 (N_14688,N_14203,N_14155);
nand U14689 (N_14689,N_14271,N_14120);
or U14690 (N_14690,N_14243,N_14392);
and U14691 (N_14691,N_14138,N_14362);
and U14692 (N_14692,N_14190,N_14130);
nor U14693 (N_14693,N_14145,N_14221);
nand U14694 (N_14694,N_14291,N_14266);
or U14695 (N_14695,N_14396,N_14122);
and U14696 (N_14696,N_14363,N_14115);
nor U14697 (N_14697,N_14259,N_14328);
xnor U14698 (N_14698,N_14102,N_14120);
or U14699 (N_14699,N_14334,N_14303);
or U14700 (N_14700,N_14683,N_14424);
nor U14701 (N_14701,N_14658,N_14616);
or U14702 (N_14702,N_14402,N_14547);
or U14703 (N_14703,N_14562,N_14540);
or U14704 (N_14704,N_14520,N_14465);
nor U14705 (N_14705,N_14446,N_14414);
nand U14706 (N_14706,N_14645,N_14571);
and U14707 (N_14707,N_14544,N_14474);
or U14708 (N_14708,N_14515,N_14431);
or U14709 (N_14709,N_14497,N_14549);
and U14710 (N_14710,N_14436,N_14605);
nand U14711 (N_14711,N_14678,N_14509);
or U14712 (N_14712,N_14621,N_14587);
or U14713 (N_14713,N_14419,N_14473);
nand U14714 (N_14714,N_14597,N_14423);
nand U14715 (N_14715,N_14570,N_14532);
and U14716 (N_14716,N_14433,N_14403);
nand U14717 (N_14717,N_14644,N_14652);
nor U14718 (N_14718,N_14684,N_14486);
nor U14719 (N_14719,N_14514,N_14657);
nor U14720 (N_14720,N_14609,N_14650);
xnor U14721 (N_14721,N_14655,N_14619);
nand U14722 (N_14722,N_14524,N_14690);
and U14723 (N_14723,N_14673,N_14416);
and U14724 (N_14724,N_14530,N_14592);
or U14725 (N_14725,N_14620,N_14654);
xnor U14726 (N_14726,N_14693,N_14687);
and U14727 (N_14727,N_14443,N_14674);
and U14728 (N_14728,N_14566,N_14457);
nand U14729 (N_14729,N_14445,N_14479);
and U14730 (N_14730,N_14458,N_14664);
and U14731 (N_14731,N_14594,N_14618);
nor U14732 (N_14732,N_14512,N_14500);
or U14733 (N_14733,N_14579,N_14490);
nor U14734 (N_14734,N_14578,N_14575);
or U14735 (N_14735,N_14613,N_14615);
and U14736 (N_14736,N_14685,N_14545);
nand U14737 (N_14737,N_14607,N_14641);
or U14738 (N_14738,N_14625,N_14430);
or U14739 (N_14739,N_14637,N_14502);
nor U14740 (N_14740,N_14591,N_14634);
nand U14741 (N_14741,N_14437,N_14406);
xnor U14742 (N_14742,N_14588,N_14535);
xor U14743 (N_14743,N_14478,N_14432);
nand U14744 (N_14744,N_14529,N_14614);
xor U14745 (N_14745,N_14438,N_14636);
and U14746 (N_14746,N_14554,N_14464);
and U14747 (N_14747,N_14508,N_14632);
and U14748 (N_14748,N_14483,N_14439);
xor U14749 (N_14749,N_14467,N_14504);
nand U14750 (N_14750,N_14598,N_14519);
and U14751 (N_14751,N_14506,N_14686);
xnor U14752 (N_14752,N_14453,N_14599);
nor U14753 (N_14753,N_14527,N_14469);
nand U14754 (N_14754,N_14600,N_14472);
nand U14755 (N_14755,N_14647,N_14489);
and U14756 (N_14756,N_14428,N_14493);
nand U14757 (N_14757,N_14682,N_14429);
nor U14758 (N_14758,N_14537,N_14447);
nor U14759 (N_14759,N_14480,N_14595);
nor U14760 (N_14760,N_14485,N_14463);
or U14761 (N_14761,N_14548,N_14496);
xnor U14762 (N_14762,N_14534,N_14679);
nor U14763 (N_14763,N_14546,N_14405);
and U14764 (N_14764,N_14553,N_14541);
or U14765 (N_14765,N_14569,N_14503);
xnor U14766 (N_14766,N_14550,N_14404);
xor U14767 (N_14767,N_14400,N_14442);
or U14768 (N_14768,N_14452,N_14501);
nor U14769 (N_14769,N_14656,N_14426);
and U14770 (N_14770,N_14585,N_14680);
nand U14771 (N_14771,N_14677,N_14451);
xor U14772 (N_14772,N_14648,N_14581);
and U14773 (N_14773,N_14676,N_14488);
xor U14774 (N_14774,N_14617,N_14456);
nand U14775 (N_14775,N_14642,N_14539);
nand U14776 (N_14776,N_14521,N_14560);
or U14777 (N_14777,N_14522,N_14696);
nor U14778 (N_14778,N_14510,N_14699);
or U14779 (N_14779,N_14671,N_14582);
nor U14780 (N_14780,N_14440,N_14460);
nor U14781 (N_14781,N_14531,N_14572);
nand U14782 (N_14782,N_14669,N_14586);
and U14783 (N_14783,N_14624,N_14583);
nor U14784 (N_14784,N_14408,N_14574);
xor U14785 (N_14785,N_14563,N_14499);
or U14786 (N_14786,N_14481,N_14612);
nor U14787 (N_14787,N_14455,N_14559);
or U14788 (N_14788,N_14413,N_14420);
nor U14789 (N_14789,N_14577,N_14584);
and U14790 (N_14790,N_14626,N_14412);
or U14791 (N_14791,N_14449,N_14603);
or U14792 (N_14792,N_14665,N_14606);
nand U14793 (N_14793,N_14482,N_14557);
xor U14794 (N_14794,N_14576,N_14681);
and U14795 (N_14795,N_14415,N_14694);
nor U14796 (N_14796,N_14523,N_14409);
and U14797 (N_14797,N_14561,N_14513);
nand U14798 (N_14798,N_14649,N_14695);
xor U14799 (N_14799,N_14494,N_14668);
or U14800 (N_14800,N_14660,N_14511);
xor U14801 (N_14801,N_14471,N_14698);
nand U14802 (N_14802,N_14593,N_14484);
nor U14803 (N_14803,N_14468,N_14697);
or U14804 (N_14804,N_14450,N_14418);
and U14805 (N_14805,N_14454,N_14475);
nor U14806 (N_14806,N_14635,N_14461);
and U14807 (N_14807,N_14629,N_14470);
nor U14808 (N_14808,N_14441,N_14466);
nor U14809 (N_14809,N_14516,N_14492);
xnor U14810 (N_14810,N_14608,N_14422);
and U14811 (N_14811,N_14666,N_14631);
nor U14812 (N_14812,N_14476,N_14567);
nor U14813 (N_14813,N_14551,N_14640);
and U14814 (N_14814,N_14526,N_14670);
and U14815 (N_14815,N_14639,N_14434);
nor U14816 (N_14816,N_14661,N_14633);
xnor U14817 (N_14817,N_14689,N_14622);
xnor U14818 (N_14818,N_14601,N_14643);
or U14819 (N_14819,N_14448,N_14533);
nor U14820 (N_14820,N_14638,N_14611);
nor U14821 (N_14821,N_14425,N_14435);
nor U14822 (N_14822,N_14630,N_14543);
xor U14823 (N_14823,N_14653,N_14421);
and U14824 (N_14824,N_14525,N_14555);
and U14825 (N_14825,N_14604,N_14580);
xor U14826 (N_14826,N_14672,N_14542);
and U14827 (N_14827,N_14688,N_14518);
nor U14828 (N_14828,N_14565,N_14505);
xor U14829 (N_14829,N_14667,N_14517);
or U14830 (N_14830,N_14528,N_14410);
or U14831 (N_14831,N_14651,N_14564);
and U14832 (N_14832,N_14596,N_14462);
and U14833 (N_14833,N_14623,N_14495);
and U14834 (N_14834,N_14556,N_14558);
nor U14835 (N_14835,N_14628,N_14427);
and U14836 (N_14836,N_14627,N_14589);
nor U14837 (N_14837,N_14573,N_14663);
or U14838 (N_14838,N_14477,N_14536);
nor U14839 (N_14839,N_14487,N_14610);
and U14840 (N_14840,N_14568,N_14401);
or U14841 (N_14841,N_14590,N_14407);
or U14842 (N_14842,N_14417,N_14662);
or U14843 (N_14843,N_14659,N_14491);
nand U14844 (N_14844,N_14692,N_14498);
xnor U14845 (N_14845,N_14459,N_14691);
xor U14846 (N_14846,N_14444,N_14411);
xnor U14847 (N_14847,N_14602,N_14646);
xor U14848 (N_14848,N_14538,N_14675);
xor U14849 (N_14849,N_14507,N_14552);
and U14850 (N_14850,N_14452,N_14476);
or U14851 (N_14851,N_14478,N_14487);
xnor U14852 (N_14852,N_14649,N_14536);
or U14853 (N_14853,N_14554,N_14478);
nand U14854 (N_14854,N_14551,N_14645);
and U14855 (N_14855,N_14499,N_14457);
nor U14856 (N_14856,N_14497,N_14617);
or U14857 (N_14857,N_14466,N_14523);
nand U14858 (N_14858,N_14582,N_14487);
nand U14859 (N_14859,N_14430,N_14405);
nor U14860 (N_14860,N_14578,N_14544);
nor U14861 (N_14861,N_14590,N_14495);
nand U14862 (N_14862,N_14429,N_14435);
and U14863 (N_14863,N_14553,N_14491);
xor U14864 (N_14864,N_14565,N_14550);
xor U14865 (N_14865,N_14439,N_14621);
or U14866 (N_14866,N_14606,N_14650);
xor U14867 (N_14867,N_14612,N_14640);
and U14868 (N_14868,N_14605,N_14644);
nor U14869 (N_14869,N_14450,N_14573);
or U14870 (N_14870,N_14404,N_14563);
nor U14871 (N_14871,N_14534,N_14634);
and U14872 (N_14872,N_14571,N_14403);
nand U14873 (N_14873,N_14557,N_14690);
or U14874 (N_14874,N_14634,N_14641);
or U14875 (N_14875,N_14550,N_14602);
nor U14876 (N_14876,N_14578,N_14639);
or U14877 (N_14877,N_14490,N_14606);
nor U14878 (N_14878,N_14688,N_14527);
xor U14879 (N_14879,N_14437,N_14414);
and U14880 (N_14880,N_14624,N_14564);
nand U14881 (N_14881,N_14468,N_14622);
or U14882 (N_14882,N_14493,N_14641);
xor U14883 (N_14883,N_14664,N_14494);
nor U14884 (N_14884,N_14419,N_14558);
and U14885 (N_14885,N_14475,N_14466);
nand U14886 (N_14886,N_14454,N_14466);
nand U14887 (N_14887,N_14513,N_14515);
xor U14888 (N_14888,N_14425,N_14430);
and U14889 (N_14889,N_14684,N_14552);
xor U14890 (N_14890,N_14562,N_14452);
or U14891 (N_14891,N_14470,N_14449);
xor U14892 (N_14892,N_14511,N_14655);
or U14893 (N_14893,N_14440,N_14499);
and U14894 (N_14894,N_14680,N_14520);
nand U14895 (N_14895,N_14439,N_14638);
nor U14896 (N_14896,N_14585,N_14649);
and U14897 (N_14897,N_14583,N_14666);
and U14898 (N_14898,N_14462,N_14662);
nor U14899 (N_14899,N_14527,N_14617);
and U14900 (N_14900,N_14446,N_14488);
nand U14901 (N_14901,N_14406,N_14426);
xnor U14902 (N_14902,N_14622,N_14629);
and U14903 (N_14903,N_14692,N_14545);
and U14904 (N_14904,N_14402,N_14522);
nor U14905 (N_14905,N_14483,N_14622);
nand U14906 (N_14906,N_14524,N_14688);
nand U14907 (N_14907,N_14588,N_14460);
xnor U14908 (N_14908,N_14695,N_14518);
and U14909 (N_14909,N_14437,N_14626);
xnor U14910 (N_14910,N_14611,N_14608);
and U14911 (N_14911,N_14468,N_14577);
or U14912 (N_14912,N_14528,N_14491);
or U14913 (N_14913,N_14656,N_14639);
nor U14914 (N_14914,N_14542,N_14571);
nand U14915 (N_14915,N_14457,N_14506);
nand U14916 (N_14916,N_14671,N_14693);
xnor U14917 (N_14917,N_14562,N_14552);
and U14918 (N_14918,N_14475,N_14451);
or U14919 (N_14919,N_14437,N_14400);
or U14920 (N_14920,N_14570,N_14663);
nand U14921 (N_14921,N_14583,N_14668);
or U14922 (N_14922,N_14535,N_14663);
nand U14923 (N_14923,N_14459,N_14567);
or U14924 (N_14924,N_14673,N_14473);
xor U14925 (N_14925,N_14430,N_14509);
or U14926 (N_14926,N_14506,N_14427);
nand U14927 (N_14927,N_14696,N_14549);
nor U14928 (N_14928,N_14447,N_14601);
or U14929 (N_14929,N_14575,N_14691);
and U14930 (N_14930,N_14462,N_14511);
nand U14931 (N_14931,N_14446,N_14695);
nand U14932 (N_14932,N_14616,N_14609);
xnor U14933 (N_14933,N_14647,N_14444);
and U14934 (N_14934,N_14544,N_14626);
nor U14935 (N_14935,N_14429,N_14416);
or U14936 (N_14936,N_14662,N_14641);
or U14937 (N_14937,N_14503,N_14478);
nor U14938 (N_14938,N_14423,N_14504);
and U14939 (N_14939,N_14622,N_14665);
nor U14940 (N_14940,N_14505,N_14601);
xor U14941 (N_14941,N_14425,N_14572);
or U14942 (N_14942,N_14444,N_14462);
and U14943 (N_14943,N_14659,N_14586);
or U14944 (N_14944,N_14411,N_14505);
nand U14945 (N_14945,N_14447,N_14410);
nor U14946 (N_14946,N_14683,N_14572);
nand U14947 (N_14947,N_14691,N_14637);
and U14948 (N_14948,N_14629,N_14566);
nand U14949 (N_14949,N_14599,N_14476);
nor U14950 (N_14950,N_14406,N_14485);
nor U14951 (N_14951,N_14435,N_14430);
nor U14952 (N_14952,N_14494,N_14479);
or U14953 (N_14953,N_14690,N_14606);
nor U14954 (N_14954,N_14670,N_14577);
nand U14955 (N_14955,N_14532,N_14635);
or U14956 (N_14956,N_14688,N_14574);
nand U14957 (N_14957,N_14488,N_14582);
nand U14958 (N_14958,N_14660,N_14525);
nor U14959 (N_14959,N_14653,N_14400);
xor U14960 (N_14960,N_14654,N_14449);
and U14961 (N_14961,N_14454,N_14496);
nor U14962 (N_14962,N_14597,N_14475);
or U14963 (N_14963,N_14577,N_14467);
nand U14964 (N_14964,N_14667,N_14541);
nand U14965 (N_14965,N_14406,N_14659);
and U14966 (N_14966,N_14643,N_14509);
nor U14967 (N_14967,N_14684,N_14419);
xnor U14968 (N_14968,N_14457,N_14546);
nor U14969 (N_14969,N_14591,N_14533);
xor U14970 (N_14970,N_14503,N_14474);
nand U14971 (N_14971,N_14449,N_14440);
xnor U14972 (N_14972,N_14459,N_14427);
nor U14973 (N_14973,N_14448,N_14483);
or U14974 (N_14974,N_14411,N_14673);
or U14975 (N_14975,N_14462,N_14688);
xnor U14976 (N_14976,N_14550,N_14455);
and U14977 (N_14977,N_14519,N_14579);
xor U14978 (N_14978,N_14620,N_14686);
nor U14979 (N_14979,N_14697,N_14432);
and U14980 (N_14980,N_14538,N_14692);
nand U14981 (N_14981,N_14609,N_14472);
nand U14982 (N_14982,N_14456,N_14460);
xnor U14983 (N_14983,N_14425,N_14517);
xnor U14984 (N_14984,N_14688,N_14682);
xor U14985 (N_14985,N_14418,N_14681);
nand U14986 (N_14986,N_14405,N_14510);
nor U14987 (N_14987,N_14546,N_14474);
nor U14988 (N_14988,N_14611,N_14528);
nor U14989 (N_14989,N_14449,N_14544);
or U14990 (N_14990,N_14656,N_14678);
or U14991 (N_14991,N_14460,N_14559);
and U14992 (N_14992,N_14696,N_14428);
nand U14993 (N_14993,N_14426,N_14409);
nand U14994 (N_14994,N_14608,N_14673);
and U14995 (N_14995,N_14599,N_14530);
xor U14996 (N_14996,N_14458,N_14637);
or U14997 (N_14997,N_14518,N_14582);
and U14998 (N_14998,N_14445,N_14499);
and U14999 (N_14999,N_14645,N_14554);
nand U15000 (N_15000,N_14705,N_14912);
nor U15001 (N_15001,N_14748,N_14770);
and U15002 (N_15002,N_14939,N_14818);
or U15003 (N_15003,N_14765,N_14749);
nand U15004 (N_15004,N_14791,N_14928);
and U15005 (N_15005,N_14958,N_14830);
nor U15006 (N_15006,N_14950,N_14925);
nor U15007 (N_15007,N_14789,N_14784);
or U15008 (N_15008,N_14734,N_14702);
nor U15009 (N_15009,N_14823,N_14898);
nand U15010 (N_15010,N_14817,N_14800);
xor U15011 (N_15011,N_14957,N_14975);
xnor U15012 (N_15012,N_14840,N_14799);
nor U15013 (N_15013,N_14971,N_14965);
or U15014 (N_15014,N_14771,N_14976);
xor U15015 (N_15015,N_14841,N_14948);
nand U15016 (N_15016,N_14719,N_14718);
or U15017 (N_15017,N_14875,N_14760);
nor U15018 (N_15018,N_14804,N_14988);
nor U15019 (N_15019,N_14802,N_14751);
nand U15020 (N_15020,N_14720,N_14932);
or U15021 (N_15021,N_14812,N_14968);
nor U15022 (N_15022,N_14952,N_14981);
and U15023 (N_15023,N_14831,N_14891);
xor U15024 (N_15024,N_14886,N_14710);
and U15025 (N_15025,N_14788,N_14978);
and U15026 (N_15026,N_14908,N_14721);
and U15027 (N_15027,N_14790,N_14838);
or U15028 (N_15028,N_14762,N_14805);
or U15029 (N_15029,N_14743,N_14746);
nand U15030 (N_15030,N_14803,N_14963);
nor U15031 (N_15031,N_14989,N_14938);
nand U15032 (N_15032,N_14973,N_14730);
nor U15033 (N_15033,N_14828,N_14866);
nand U15034 (N_15034,N_14853,N_14846);
nor U15035 (N_15035,N_14844,N_14873);
nor U15036 (N_15036,N_14745,N_14781);
xor U15037 (N_15037,N_14808,N_14763);
xor U15038 (N_15038,N_14826,N_14897);
or U15039 (N_15039,N_14707,N_14909);
and U15040 (N_15040,N_14921,N_14955);
nand U15041 (N_15041,N_14930,N_14915);
nand U15042 (N_15042,N_14813,N_14956);
nor U15043 (N_15043,N_14712,N_14951);
xor U15044 (N_15044,N_14824,N_14913);
xor U15045 (N_15045,N_14755,N_14929);
xnor U15046 (N_15046,N_14836,N_14792);
xnor U15047 (N_15047,N_14741,N_14851);
and U15048 (N_15048,N_14786,N_14994);
and U15049 (N_15049,N_14797,N_14785);
nor U15050 (N_15050,N_14714,N_14920);
nor U15051 (N_15051,N_14814,N_14954);
nand U15052 (N_15052,N_14884,N_14880);
nand U15053 (N_15053,N_14703,N_14991);
or U15054 (N_15054,N_14953,N_14907);
nand U15055 (N_15055,N_14967,N_14758);
and U15056 (N_15056,N_14764,N_14768);
xnor U15057 (N_15057,N_14895,N_14821);
nor U15058 (N_15058,N_14940,N_14737);
nand U15059 (N_15059,N_14827,N_14871);
nor U15060 (N_15060,N_14944,N_14711);
and U15061 (N_15061,N_14927,N_14878);
and U15062 (N_15062,N_14985,N_14924);
xor U15063 (N_15063,N_14782,N_14847);
xor U15064 (N_15064,N_14723,N_14852);
or U15065 (N_15065,N_14961,N_14858);
or U15066 (N_15066,N_14881,N_14704);
nand U15067 (N_15067,N_14761,N_14811);
nor U15068 (N_15068,N_14708,N_14996);
nor U15069 (N_15069,N_14717,N_14816);
and U15070 (N_15070,N_14753,N_14914);
nand U15071 (N_15071,N_14834,N_14835);
nor U15072 (N_15072,N_14807,N_14972);
and U15073 (N_15073,N_14776,N_14937);
nor U15074 (N_15074,N_14859,N_14896);
xnor U15075 (N_15075,N_14868,N_14864);
or U15076 (N_15076,N_14888,N_14740);
xnor U15077 (N_15077,N_14725,N_14713);
nor U15078 (N_15078,N_14874,N_14892);
nor U15079 (N_15079,N_14902,N_14934);
or U15080 (N_15080,N_14949,N_14829);
or U15081 (N_15081,N_14992,N_14845);
nand U15082 (N_15082,N_14867,N_14822);
nand U15083 (N_15083,N_14806,N_14700);
and U15084 (N_15084,N_14923,N_14906);
nand U15085 (N_15085,N_14728,N_14732);
nor U15086 (N_15086,N_14706,N_14890);
nor U15087 (N_15087,N_14879,N_14742);
and U15088 (N_15088,N_14772,N_14942);
xor U15089 (N_15089,N_14837,N_14854);
and U15090 (N_15090,N_14918,N_14872);
nand U15091 (N_15091,N_14987,N_14960);
nand U15092 (N_15092,N_14750,N_14941);
nand U15093 (N_15093,N_14794,N_14919);
and U15094 (N_15094,N_14865,N_14964);
or U15095 (N_15095,N_14795,N_14769);
nor U15096 (N_15096,N_14798,N_14722);
nor U15097 (N_15097,N_14777,N_14999);
xor U15098 (N_15098,N_14860,N_14839);
or U15099 (N_15099,N_14701,N_14820);
nor U15100 (N_15100,N_14778,N_14856);
xnor U15101 (N_15101,N_14855,N_14861);
or U15102 (N_15102,N_14980,N_14849);
and U15103 (N_15103,N_14716,N_14709);
nor U15104 (N_15104,N_14774,N_14984);
nor U15105 (N_15105,N_14773,N_14801);
and U15106 (N_15106,N_14993,N_14810);
nand U15107 (N_15107,N_14756,N_14966);
nand U15108 (N_15108,N_14974,N_14885);
and U15109 (N_15109,N_14889,N_14945);
nand U15110 (N_15110,N_14825,N_14995);
or U15111 (N_15111,N_14910,N_14959);
nand U15112 (N_15112,N_14883,N_14903);
xor U15113 (N_15113,N_14943,N_14744);
xnor U15114 (N_15114,N_14935,N_14809);
xnor U15115 (N_15115,N_14936,N_14848);
nand U15116 (N_15116,N_14979,N_14731);
nor U15117 (N_15117,N_14747,N_14899);
and U15118 (N_15118,N_14986,N_14962);
nor U15119 (N_15119,N_14983,N_14911);
and U15120 (N_15120,N_14922,N_14733);
or U15121 (N_15121,N_14933,N_14982);
nor U15122 (N_15122,N_14931,N_14729);
xnor U15123 (N_15123,N_14775,N_14833);
or U15124 (N_15124,N_14882,N_14726);
nor U15125 (N_15125,N_14904,N_14926);
nand U15126 (N_15126,N_14997,N_14894);
xnor U15127 (N_15127,N_14857,N_14727);
xnor U15128 (N_15128,N_14870,N_14787);
nor U15129 (N_15129,N_14796,N_14832);
xor U15130 (N_15130,N_14752,N_14715);
nor U15131 (N_15131,N_14738,N_14917);
nor U15132 (N_15132,N_14977,N_14893);
xnor U15133 (N_15133,N_14946,N_14759);
or U15134 (N_15134,N_14998,N_14905);
nand U15135 (N_15135,N_14842,N_14735);
and U15136 (N_15136,N_14869,N_14739);
or U15137 (N_15137,N_14916,N_14757);
and U15138 (N_15138,N_14783,N_14947);
xor U15139 (N_15139,N_14819,N_14754);
nand U15140 (N_15140,N_14815,N_14876);
or U15141 (N_15141,N_14887,N_14843);
nor U15142 (N_15142,N_14969,N_14900);
nand U15143 (N_15143,N_14779,N_14736);
nor U15144 (N_15144,N_14766,N_14901);
xor U15145 (N_15145,N_14793,N_14990);
xnor U15146 (N_15146,N_14724,N_14862);
or U15147 (N_15147,N_14780,N_14970);
nor U15148 (N_15148,N_14863,N_14767);
or U15149 (N_15149,N_14877,N_14850);
nand U15150 (N_15150,N_14862,N_14976);
nor U15151 (N_15151,N_14952,N_14822);
xor U15152 (N_15152,N_14969,N_14892);
nor U15153 (N_15153,N_14811,N_14862);
nor U15154 (N_15154,N_14834,N_14927);
xor U15155 (N_15155,N_14860,N_14733);
or U15156 (N_15156,N_14795,N_14985);
nor U15157 (N_15157,N_14766,N_14865);
nand U15158 (N_15158,N_14802,N_14778);
xnor U15159 (N_15159,N_14928,N_14907);
and U15160 (N_15160,N_14765,N_14895);
or U15161 (N_15161,N_14887,N_14738);
nor U15162 (N_15162,N_14957,N_14797);
nor U15163 (N_15163,N_14956,N_14935);
nor U15164 (N_15164,N_14783,N_14989);
nand U15165 (N_15165,N_14713,N_14801);
and U15166 (N_15166,N_14923,N_14937);
nor U15167 (N_15167,N_14806,N_14856);
or U15168 (N_15168,N_14892,N_14794);
nor U15169 (N_15169,N_14761,N_14925);
xor U15170 (N_15170,N_14938,N_14824);
xor U15171 (N_15171,N_14878,N_14962);
or U15172 (N_15172,N_14883,N_14820);
and U15173 (N_15173,N_14849,N_14781);
xor U15174 (N_15174,N_14972,N_14737);
nor U15175 (N_15175,N_14855,N_14808);
xnor U15176 (N_15176,N_14950,N_14904);
and U15177 (N_15177,N_14855,N_14937);
and U15178 (N_15178,N_14890,N_14946);
nand U15179 (N_15179,N_14877,N_14808);
and U15180 (N_15180,N_14812,N_14839);
or U15181 (N_15181,N_14965,N_14901);
xnor U15182 (N_15182,N_14866,N_14963);
xnor U15183 (N_15183,N_14749,N_14810);
nor U15184 (N_15184,N_14970,N_14762);
xnor U15185 (N_15185,N_14947,N_14793);
or U15186 (N_15186,N_14722,N_14896);
nand U15187 (N_15187,N_14845,N_14915);
xnor U15188 (N_15188,N_14970,N_14952);
and U15189 (N_15189,N_14978,N_14962);
nand U15190 (N_15190,N_14748,N_14977);
xor U15191 (N_15191,N_14939,N_14949);
and U15192 (N_15192,N_14746,N_14748);
or U15193 (N_15193,N_14809,N_14831);
or U15194 (N_15194,N_14800,N_14899);
nor U15195 (N_15195,N_14729,N_14751);
or U15196 (N_15196,N_14822,N_14878);
nor U15197 (N_15197,N_14991,N_14752);
or U15198 (N_15198,N_14840,N_14963);
nor U15199 (N_15199,N_14846,N_14821);
xnor U15200 (N_15200,N_14947,N_14823);
or U15201 (N_15201,N_14858,N_14710);
xor U15202 (N_15202,N_14951,N_14881);
nor U15203 (N_15203,N_14998,N_14971);
and U15204 (N_15204,N_14784,N_14979);
or U15205 (N_15205,N_14931,N_14914);
xnor U15206 (N_15206,N_14798,N_14850);
and U15207 (N_15207,N_14873,N_14868);
xnor U15208 (N_15208,N_14802,N_14765);
nand U15209 (N_15209,N_14764,N_14991);
nor U15210 (N_15210,N_14725,N_14743);
or U15211 (N_15211,N_14844,N_14843);
xnor U15212 (N_15212,N_14834,N_14883);
and U15213 (N_15213,N_14764,N_14942);
nor U15214 (N_15214,N_14939,N_14794);
and U15215 (N_15215,N_14813,N_14989);
xor U15216 (N_15216,N_14937,N_14715);
nor U15217 (N_15217,N_14797,N_14760);
xor U15218 (N_15218,N_14845,N_14986);
and U15219 (N_15219,N_14768,N_14834);
and U15220 (N_15220,N_14853,N_14708);
nor U15221 (N_15221,N_14701,N_14722);
and U15222 (N_15222,N_14714,N_14810);
or U15223 (N_15223,N_14788,N_14983);
nor U15224 (N_15224,N_14917,N_14824);
or U15225 (N_15225,N_14851,N_14839);
xnor U15226 (N_15226,N_14787,N_14766);
nand U15227 (N_15227,N_14940,N_14896);
or U15228 (N_15228,N_14832,N_14728);
and U15229 (N_15229,N_14988,N_14837);
xnor U15230 (N_15230,N_14990,N_14863);
and U15231 (N_15231,N_14776,N_14987);
nor U15232 (N_15232,N_14998,N_14715);
xor U15233 (N_15233,N_14984,N_14934);
nor U15234 (N_15234,N_14970,N_14869);
and U15235 (N_15235,N_14776,N_14735);
or U15236 (N_15236,N_14709,N_14805);
nor U15237 (N_15237,N_14841,N_14760);
nor U15238 (N_15238,N_14928,N_14721);
nor U15239 (N_15239,N_14965,N_14984);
nand U15240 (N_15240,N_14886,N_14957);
nor U15241 (N_15241,N_14802,N_14974);
xnor U15242 (N_15242,N_14899,N_14903);
xnor U15243 (N_15243,N_14785,N_14788);
nor U15244 (N_15244,N_14717,N_14982);
nand U15245 (N_15245,N_14856,N_14893);
and U15246 (N_15246,N_14902,N_14724);
nor U15247 (N_15247,N_14985,N_14759);
nor U15248 (N_15248,N_14952,N_14734);
nor U15249 (N_15249,N_14716,N_14914);
xor U15250 (N_15250,N_14995,N_14870);
or U15251 (N_15251,N_14767,N_14898);
or U15252 (N_15252,N_14944,N_14840);
nor U15253 (N_15253,N_14755,N_14904);
nand U15254 (N_15254,N_14883,N_14983);
and U15255 (N_15255,N_14827,N_14768);
nand U15256 (N_15256,N_14746,N_14734);
and U15257 (N_15257,N_14886,N_14989);
or U15258 (N_15258,N_14737,N_14938);
nor U15259 (N_15259,N_14826,N_14849);
nor U15260 (N_15260,N_14785,N_14858);
nor U15261 (N_15261,N_14800,N_14950);
nor U15262 (N_15262,N_14728,N_14778);
and U15263 (N_15263,N_14790,N_14780);
nand U15264 (N_15264,N_14961,N_14718);
and U15265 (N_15265,N_14805,N_14990);
xor U15266 (N_15266,N_14805,N_14753);
nor U15267 (N_15267,N_14775,N_14886);
xnor U15268 (N_15268,N_14713,N_14959);
nor U15269 (N_15269,N_14811,N_14831);
and U15270 (N_15270,N_14712,N_14929);
or U15271 (N_15271,N_14858,N_14849);
nor U15272 (N_15272,N_14742,N_14716);
nor U15273 (N_15273,N_14998,N_14708);
nor U15274 (N_15274,N_14736,N_14812);
nand U15275 (N_15275,N_14736,N_14870);
and U15276 (N_15276,N_14747,N_14827);
and U15277 (N_15277,N_14979,N_14870);
xor U15278 (N_15278,N_14808,N_14724);
nand U15279 (N_15279,N_14895,N_14757);
nor U15280 (N_15280,N_14780,N_14787);
or U15281 (N_15281,N_14908,N_14740);
xor U15282 (N_15282,N_14830,N_14802);
xnor U15283 (N_15283,N_14904,N_14700);
and U15284 (N_15284,N_14833,N_14780);
nor U15285 (N_15285,N_14818,N_14947);
or U15286 (N_15286,N_14847,N_14932);
nand U15287 (N_15287,N_14937,N_14932);
or U15288 (N_15288,N_14920,N_14710);
nand U15289 (N_15289,N_14810,N_14745);
or U15290 (N_15290,N_14834,N_14896);
and U15291 (N_15291,N_14722,N_14805);
or U15292 (N_15292,N_14901,N_14720);
and U15293 (N_15293,N_14724,N_14765);
and U15294 (N_15294,N_14929,N_14985);
and U15295 (N_15295,N_14784,N_14879);
nand U15296 (N_15296,N_14741,N_14731);
or U15297 (N_15297,N_14834,N_14774);
xor U15298 (N_15298,N_14705,N_14916);
or U15299 (N_15299,N_14725,N_14842);
nand U15300 (N_15300,N_15190,N_15277);
and U15301 (N_15301,N_15021,N_15249);
and U15302 (N_15302,N_15083,N_15033);
xnor U15303 (N_15303,N_15215,N_15245);
nand U15304 (N_15304,N_15124,N_15231);
or U15305 (N_15305,N_15278,N_15018);
or U15306 (N_15306,N_15099,N_15123);
and U15307 (N_15307,N_15029,N_15141);
xor U15308 (N_15308,N_15158,N_15267);
nand U15309 (N_15309,N_15187,N_15125);
nand U15310 (N_15310,N_15074,N_15180);
nor U15311 (N_15311,N_15129,N_15292);
xnor U15312 (N_15312,N_15193,N_15241);
nand U15313 (N_15313,N_15214,N_15285);
and U15314 (N_15314,N_15131,N_15096);
or U15315 (N_15315,N_15117,N_15023);
or U15316 (N_15316,N_15203,N_15053);
xnor U15317 (N_15317,N_15163,N_15110);
xor U15318 (N_15318,N_15262,N_15229);
nand U15319 (N_15319,N_15075,N_15050);
xnor U15320 (N_15320,N_15243,N_15031);
xor U15321 (N_15321,N_15042,N_15143);
or U15322 (N_15322,N_15156,N_15005);
xnor U15323 (N_15323,N_15224,N_15258);
nand U15324 (N_15324,N_15233,N_15000);
nand U15325 (N_15325,N_15048,N_15045);
or U15326 (N_15326,N_15162,N_15036);
or U15327 (N_15327,N_15072,N_15259);
nand U15328 (N_15328,N_15264,N_15294);
xnor U15329 (N_15329,N_15127,N_15173);
xnor U15330 (N_15330,N_15228,N_15006);
xor U15331 (N_15331,N_15035,N_15137);
nand U15332 (N_15332,N_15108,N_15236);
nor U15333 (N_15333,N_15254,N_15057);
nand U15334 (N_15334,N_15255,N_15271);
nor U15335 (N_15335,N_15199,N_15116);
nor U15336 (N_15336,N_15211,N_15153);
and U15337 (N_15337,N_15207,N_15183);
and U15338 (N_15338,N_15081,N_15133);
nor U15339 (N_15339,N_15238,N_15280);
xnor U15340 (N_15340,N_15220,N_15273);
nand U15341 (N_15341,N_15253,N_15140);
nor U15342 (N_15342,N_15147,N_15044);
and U15343 (N_15343,N_15232,N_15295);
nor U15344 (N_15344,N_15148,N_15047);
xor U15345 (N_15345,N_15178,N_15296);
nor U15346 (N_15346,N_15136,N_15174);
nand U15347 (N_15347,N_15113,N_15019);
or U15348 (N_15348,N_15168,N_15065);
nand U15349 (N_15349,N_15219,N_15188);
xnor U15350 (N_15350,N_15272,N_15052);
nand U15351 (N_15351,N_15080,N_15145);
xor U15352 (N_15352,N_15161,N_15275);
nor U15353 (N_15353,N_15201,N_15266);
nor U15354 (N_15354,N_15157,N_15028);
or U15355 (N_15355,N_15092,N_15119);
xnor U15356 (N_15356,N_15223,N_15288);
xor U15357 (N_15357,N_15112,N_15287);
xor U15358 (N_15358,N_15009,N_15256);
and U15359 (N_15359,N_15206,N_15059);
and U15360 (N_15360,N_15177,N_15164);
nor U15361 (N_15361,N_15024,N_15134);
xor U15362 (N_15362,N_15251,N_15204);
nand U15363 (N_15363,N_15290,N_15221);
xor U15364 (N_15364,N_15185,N_15093);
nor U15365 (N_15365,N_15195,N_15063);
xnor U15366 (N_15366,N_15212,N_15120);
nand U15367 (N_15367,N_15062,N_15240);
nand U15368 (N_15368,N_15208,N_15008);
nand U15369 (N_15369,N_15181,N_15128);
nor U15370 (N_15370,N_15011,N_15087);
and U15371 (N_15371,N_15122,N_15013);
nand U15372 (N_15372,N_15082,N_15237);
nor U15373 (N_15373,N_15297,N_15291);
xor U15374 (N_15374,N_15091,N_15166);
xnor U15375 (N_15375,N_15084,N_15118);
nor U15376 (N_15376,N_15283,N_15071);
nand U15377 (N_15377,N_15175,N_15234);
nor U15378 (N_15378,N_15076,N_15269);
xor U15379 (N_15379,N_15067,N_15089);
or U15380 (N_15380,N_15126,N_15025);
nor U15381 (N_15381,N_15090,N_15130);
nor U15382 (N_15382,N_15105,N_15061);
and U15383 (N_15383,N_15012,N_15261);
xnor U15384 (N_15384,N_15165,N_15051);
nand U15385 (N_15385,N_15216,N_15289);
or U15386 (N_15386,N_15154,N_15149);
xnor U15387 (N_15387,N_15106,N_15260);
xnor U15388 (N_15388,N_15286,N_15189);
or U15389 (N_15389,N_15152,N_15002);
nand U15390 (N_15390,N_15003,N_15041);
nand U15391 (N_15391,N_15022,N_15194);
or U15392 (N_15392,N_15077,N_15121);
xnor U15393 (N_15393,N_15197,N_15104);
nand U15394 (N_15394,N_15070,N_15046);
nor U15395 (N_15395,N_15274,N_15010);
nor U15396 (N_15396,N_15202,N_15058);
and U15397 (N_15397,N_15226,N_15270);
and U15398 (N_15398,N_15100,N_15094);
and U15399 (N_15399,N_15073,N_15111);
nand U15400 (N_15400,N_15135,N_15184);
xor U15401 (N_15401,N_15169,N_15200);
nor U15402 (N_15402,N_15179,N_15218);
xnor U15403 (N_15403,N_15142,N_15026);
and U15404 (N_15404,N_15244,N_15016);
nand U15405 (N_15405,N_15015,N_15167);
nor U15406 (N_15406,N_15056,N_15066);
or U15407 (N_15407,N_15186,N_15055);
nor U15408 (N_15408,N_15132,N_15176);
xnor U15409 (N_15409,N_15284,N_15034);
nor U15410 (N_15410,N_15032,N_15281);
nor U15411 (N_15411,N_15160,N_15155);
xnor U15412 (N_15412,N_15144,N_15217);
xor U15413 (N_15413,N_15196,N_15151);
nor U15414 (N_15414,N_15230,N_15276);
xor U15415 (N_15415,N_15222,N_15014);
nand U15416 (N_15416,N_15250,N_15268);
or U15417 (N_15417,N_15114,N_15299);
and U15418 (N_15418,N_15054,N_15020);
xor U15419 (N_15419,N_15027,N_15043);
nand U15420 (N_15420,N_15101,N_15263);
or U15421 (N_15421,N_15038,N_15060);
xor U15422 (N_15422,N_15007,N_15192);
nor U15423 (N_15423,N_15248,N_15171);
or U15424 (N_15424,N_15037,N_15064);
nor U15425 (N_15425,N_15039,N_15239);
or U15426 (N_15426,N_15095,N_15227);
and U15427 (N_15427,N_15191,N_15293);
and U15428 (N_15428,N_15138,N_15170);
or U15429 (N_15429,N_15107,N_15150);
xor U15430 (N_15430,N_15235,N_15225);
nand U15431 (N_15431,N_15001,N_15004);
xnor U15432 (N_15432,N_15298,N_15068);
xnor U15433 (N_15433,N_15069,N_15279);
and U15434 (N_15434,N_15242,N_15282);
nand U15435 (N_15435,N_15213,N_15086);
nand U15436 (N_15436,N_15246,N_15079);
xnor U15437 (N_15437,N_15210,N_15146);
nor U15438 (N_15438,N_15030,N_15098);
or U15439 (N_15439,N_15102,N_15049);
nor U15440 (N_15440,N_15078,N_15247);
nor U15441 (N_15441,N_15017,N_15109);
nand U15442 (N_15442,N_15172,N_15097);
nand U15443 (N_15443,N_15209,N_15085);
xor U15444 (N_15444,N_15205,N_15103);
nand U15445 (N_15445,N_15265,N_15040);
nand U15446 (N_15446,N_15088,N_15159);
nor U15447 (N_15447,N_15198,N_15182);
and U15448 (N_15448,N_15115,N_15257);
or U15449 (N_15449,N_15139,N_15252);
or U15450 (N_15450,N_15020,N_15060);
or U15451 (N_15451,N_15140,N_15014);
nand U15452 (N_15452,N_15153,N_15212);
or U15453 (N_15453,N_15224,N_15026);
nor U15454 (N_15454,N_15238,N_15180);
nand U15455 (N_15455,N_15165,N_15076);
xor U15456 (N_15456,N_15285,N_15226);
or U15457 (N_15457,N_15194,N_15265);
nand U15458 (N_15458,N_15201,N_15072);
or U15459 (N_15459,N_15168,N_15111);
or U15460 (N_15460,N_15029,N_15224);
nor U15461 (N_15461,N_15158,N_15107);
nor U15462 (N_15462,N_15073,N_15045);
and U15463 (N_15463,N_15241,N_15256);
or U15464 (N_15464,N_15007,N_15015);
and U15465 (N_15465,N_15102,N_15043);
xor U15466 (N_15466,N_15000,N_15017);
nor U15467 (N_15467,N_15072,N_15210);
nor U15468 (N_15468,N_15117,N_15231);
and U15469 (N_15469,N_15068,N_15135);
xor U15470 (N_15470,N_15250,N_15231);
xor U15471 (N_15471,N_15039,N_15041);
or U15472 (N_15472,N_15061,N_15191);
nor U15473 (N_15473,N_15128,N_15193);
nor U15474 (N_15474,N_15171,N_15261);
nand U15475 (N_15475,N_15161,N_15127);
or U15476 (N_15476,N_15114,N_15101);
nand U15477 (N_15477,N_15187,N_15226);
xor U15478 (N_15478,N_15155,N_15168);
and U15479 (N_15479,N_15192,N_15228);
nor U15480 (N_15480,N_15202,N_15226);
and U15481 (N_15481,N_15260,N_15014);
or U15482 (N_15482,N_15181,N_15249);
and U15483 (N_15483,N_15035,N_15116);
nand U15484 (N_15484,N_15101,N_15276);
and U15485 (N_15485,N_15041,N_15168);
or U15486 (N_15486,N_15016,N_15198);
or U15487 (N_15487,N_15070,N_15055);
or U15488 (N_15488,N_15295,N_15013);
nand U15489 (N_15489,N_15193,N_15037);
or U15490 (N_15490,N_15094,N_15261);
and U15491 (N_15491,N_15022,N_15123);
and U15492 (N_15492,N_15216,N_15159);
nor U15493 (N_15493,N_15028,N_15030);
or U15494 (N_15494,N_15040,N_15076);
or U15495 (N_15495,N_15137,N_15208);
xor U15496 (N_15496,N_15118,N_15264);
xnor U15497 (N_15497,N_15254,N_15234);
nand U15498 (N_15498,N_15195,N_15031);
nor U15499 (N_15499,N_15185,N_15000);
and U15500 (N_15500,N_15093,N_15105);
or U15501 (N_15501,N_15202,N_15006);
nand U15502 (N_15502,N_15199,N_15196);
nor U15503 (N_15503,N_15206,N_15040);
nand U15504 (N_15504,N_15065,N_15061);
and U15505 (N_15505,N_15023,N_15218);
nand U15506 (N_15506,N_15128,N_15268);
nand U15507 (N_15507,N_15038,N_15047);
xnor U15508 (N_15508,N_15091,N_15045);
nand U15509 (N_15509,N_15274,N_15241);
xor U15510 (N_15510,N_15030,N_15175);
nand U15511 (N_15511,N_15008,N_15161);
and U15512 (N_15512,N_15117,N_15124);
or U15513 (N_15513,N_15193,N_15060);
nor U15514 (N_15514,N_15236,N_15016);
nor U15515 (N_15515,N_15115,N_15284);
nand U15516 (N_15516,N_15024,N_15132);
nand U15517 (N_15517,N_15035,N_15070);
nor U15518 (N_15518,N_15143,N_15247);
and U15519 (N_15519,N_15024,N_15056);
or U15520 (N_15520,N_15132,N_15111);
nand U15521 (N_15521,N_15176,N_15133);
and U15522 (N_15522,N_15094,N_15092);
and U15523 (N_15523,N_15298,N_15151);
nor U15524 (N_15524,N_15100,N_15099);
nand U15525 (N_15525,N_15004,N_15204);
nor U15526 (N_15526,N_15055,N_15254);
or U15527 (N_15527,N_15091,N_15080);
xor U15528 (N_15528,N_15080,N_15214);
and U15529 (N_15529,N_15128,N_15046);
nor U15530 (N_15530,N_15026,N_15254);
nand U15531 (N_15531,N_15203,N_15018);
or U15532 (N_15532,N_15052,N_15255);
and U15533 (N_15533,N_15155,N_15145);
xor U15534 (N_15534,N_15147,N_15053);
or U15535 (N_15535,N_15061,N_15101);
and U15536 (N_15536,N_15213,N_15115);
or U15537 (N_15537,N_15042,N_15017);
nand U15538 (N_15538,N_15162,N_15009);
nor U15539 (N_15539,N_15082,N_15102);
or U15540 (N_15540,N_15087,N_15182);
nand U15541 (N_15541,N_15248,N_15040);
nand U15542 (N_15542,N_15256,N_15115);
nand U15543 (N_15543,N_15271,N_15107);
or U15544 (N_15544,N_15039,N_15276);
nand U15545 (N_15545,N_15238,N_15119);
and U15546 (N_15546,N_15202,N_15109);
and U15547 (N_15547,N_15193,N_15243);
and U15548 (N_15548,N_15037,N_15044);
nand U15549 (N_15549,N_15022,N_15172);
nand U15550 (N_15550,N_15228,N_15128);
or U15551 (N_15551,N_15004,N_15017);
nand U15552 (N_15552,N_15101,N_15105);
or U15553 (N_15553,N_15235,N_15106);
xor U15554 (N_15554,N_15251,N_15244);
xor U15555 (N_15555,N_15029,N_15053);
or U15556 (N_15556,N_15120,N_15279);
nand U15557 (N_15557,N_15212,N_15014);
xnor U15558 (N_15558,N_15115,N_15042);
xnor U15559 (N_15559,N_15206,N_15068);
nand U15560 (N_15560,N_15185,N_15206);
nor U15561 (N_15561,N_15138,N_15083);
nor U15562 (N_15562,N_15012,N_15055);
or U15563 (N_15563,N_15261,N_15246);
and U15564 (N_15564,N_15196,N_15214);
xor U15565 (N_15565,N_15041,N_15287);
and U15566 (N_15566,N_15162,N_15264);
and U15567 (N_15567,N_15214,N_15061);
or U15568 (N_15568,N_15180,N_15177);
nor U15569 (N_15569,N_15136,N_15127);
nand U15570 (N_15570,N_15120,N_15127);
and U15571 (N_15571,N_15207,N_15090);
and U15572 (N_15572,N_15011,N_15181);
or U15573 (N_15573,N_15134,N_15040);
or U15574 (N_15574,N_15063,N_15266);
xnor U15575 (N_15575,N_15204,N_15245);
or U15576 (N_15576,N_15283,N_15148);
or U15577 (N_15577,N_15263,N_15230);
nor U15578 (N_15578,N_15147,N_15115);
or U15579 (N_15579,N_15164,N_15054);
xnor U15580 (N_15580,N_15145,N_15019);
xnor U15581 (N_15581,N_15130,N_15047);
xor U15582 (N_15582,N_15048,N_15260);
xnor U15583 (N_15583,N_15003,N_15179);
or U15584 (N_15584,N_15287,N_15176);
xnor U15585 (N_15585,N_15074,N_15175);
or U15586 (N_15586,N_15239,N_15166);
xor U15587 (N_15587,N_15217,N_15173);
and U15588 (N_15588,N_15284,N_15058);
nor U15589 (N_15589,N_15027,N_15154);
nand U15590 (N_15590,N_15140,N_15177);
nor U15591 (N_15591,N_15027,N_15049);
nand U15592 (N_15592,N_15058,N_15236);
or U15593 (N_15593,N_15038,N_15262);
xor U15594 (N_15594,N_15124,N_15045);
nand U15595 (N_15595,N_15209,N_15053);
nand U15596 (N_15596,N_15162,N_15145);
nor U15597 (N_15597,N_15059,N_15212);
xnor U15598 (N_15598,N_15039,N_15031);
xnor U15599 (N_15599,N_15091,N_15081);
nand U15600 (N_15600,N_15377,N_15304);
and U15601 (N_15601,N_15349,N_15347);
xnor U15602 (N_15602,N_15498,N_15523);
xor U15603 (N_15603,N_15301,N_15562);
nor U15604 (N_15604,N_15465,N_15521);
xor U15605 (N_15605,N_15487,N_15309);
nand U15606 (N_15606,N_15356,N_15387);
nand U15607 (N_15607,N_15386,N_15401);
and U15608 (N_15608,N_15431,N_15403);
or U15609 (N_15609,N_15329,N_15569);
xnor U15610 (N_15610,N_15362,N_15322);
xor U15611 (N_15611,N_15565,N_15365);
and U15612 (N_15612,N_15575,N_15508);
nor U15613 (N_15613,N_15528,N_15306);
and U15614 (N_15614,N_15519,N_15328);
nor U15615 (N_15615,N_15504,N_15480);
and U15616 (N_15616,N_15315,N_15564);
nor U15617 (N_15617,N_15570,N_15559);
and U15618 (N_15618,N_15469,N_15422);
and U15619 (N_15619,N_15332,N_15497);
nand U15620 (N_15620,N_15314,N_15448);
xor U15621 (N_15621,N_15444,N_15512);
xor U15622 (N_15622,N_15358,N_15415);
or U15623 (N_15623,N_15320,N_15516);
or U15624 (N_15624,N_15408,N_15539);
or U15625 (N_15625,N_15524,N_15405);
xnor U15626 (N_15626,N_15589,N_15454);
or U15627 (N_15627,N_15360,N_15479);
xnor U15628 (N_15628,N_15433,N_15568);
and U15629 (N_15629,N_15407,N_15493);
and U15630 (N_15630,N_15331,N_15507);
xor U15631 (N_15631,N_15369,N_15544);
or U15632 (N_15632,N_15390,N_15475);
and U15633 (N_15633,N_15492,N_15501);
xor U15634 (N_15634,N_15319,N_15558);
or U15635 (N_15635,N_15513,N_15404);
xnor U15636 (N_15636,N_15580,N_15368);
or U15637 (N_15637,N_15485,N_15346);
nor U15638 (N_15638,N_15579,N_15338);
nor U15639 (N_15639,N_15577,N_15445);
nand U15640 (N_15640,N_15560,N_15550);
xnor U15641 (N_15641,N_15409,N_15423);
and U15642 (N_15642,N_15452,N_15510);
xor U15643 (N_15643,N_15364,N_15416);
and U15644 (N_15644,N_15552,N_15354);
nor U15645 (N_15645,N_15323,N_15476);
nor U15646 (N_15646,N_15527,N_15361);
nor U15647 (N_15647,N_15483,N_15472);
nor U15648 (N_15648,N_15394,N_15583);
and U15649 (N_15649,N_15437,N_15406);
nand U15650 (N_15650,N_15592,N_15532);
or U15651 (N_15651,N_15343,N_15363);
xor U15652 (N_15652,N_15436,N_15514);
nand U15653 (N_15653,N_15491,N_15460);
or U15654 (N_15654,N_15573,N_15378);
xnor U15655 (N_15655,N_15553,N_15556);
or U15656 (N_15656,N_15334,N_15313);
nor U15657 (N_15657,N_15372,N_15353);
and U15658 (N_15658,N_15376,N_15417);
nand U15659 (N_15659,N_15463,N_15312);
nor U15660 (N_15660,N_15587,N_15359);
xor U15661 (N_15661,N_15515,N_15542);
and U15662 (N_15662,N_15549,N_15543);
or U15663 (N_15663,N_15595,N_15490);
and U15664 (N_15664,N_15581,N_15341);
nand U15665 (N_15665,N_15432,N_15438);
and U15666 (N_15666,N_15434,N_15351);
nor U15667 (N_15667,N_15379,N_15590);
or U15668 (N_15668,N_15529,N_15317);
or U15669 (N_15669,N_15461,N_15541);
or U15670 (N_15670,N_15414,N_15427);
or U15671 (N_15671,N_15350,N_15509);
xnor U15672 (N_15672,N_15375,N_15467);
xor U15673 (N_15673,N_15505,N_15447);
and U15674 (N_15674,N_15588,N_15574);
and U15675 (N_15675,N_15392,N_15426);
nor U15676 (N_15676,N_15382,N_15496);
nand U15677 (N_15677,N_15400,N_15591);
nor U15678 (N_15678,N_15450,N_15371);
xnor U15679 (N_15679,N_15473,N_15398);
or U15680 (N_15680,N_15495,N_15596);
nor U15681 (N_15681,N_15458,N_15345);
and U15682 (N_15682,N_15333,N_15525);
xor U15683 (N_15683,N_15411,N_15443);
xor U15684 (N_15684,N_15477,N_15446);
nor U15685 (N_15685,N_15425,N_15385);
nand U15686 (N_15686,N_15468,N_15395);
and U15687 (N_15687,N_15518,N_15388);
nor U15688 (N_15688,N_15462,N_15316);
or U15689 (N_15689,N_15474,N_15488);
or U15690 (N_15690,N_15336,N_15547);
nor U15691 (N_15691,N_15321,N_15537);
nor U15692 (N_15692,N_15344,N_15563);
or U15693 (N_15693,N_15367,N_15453);
or U15694 (N_15694,N_15548,N_15397);
nand U15695 (N_15695,N_15545,N_15486);
nor U15696 (N_15696,N_15418,N_15374);
and U15697 (N_15697,N_15335,N_15307);
and U15698 (N_15698,N_15500,N_15511);
nor U15699 (N_15699,N_15561,N_15326);
nor U15700 (N_15700,N_15484,N_15530);
xnor U15701 (N_15701,N_15370,N_15302);
and U15702 (N_15702,N_15419,N_15534);
or U15703 (N_15703,N_15303,N_15348);
xnor U15704 (N_15704,N_15383,N_15451);
or U15705 (N_15705,N_15526,N_15520);
or U15706 (N_15706,N_15481,N_15435);
nor U15707 (N_15707,N_15311,N_15324);
nand U15708 (N_15708,N_15413,N_15586);
nand U15709 (N_15709,N_15424,N_15554);
xnor U15710 (N_15710,N_15459,N_15381);
nand U15711 (N_15711,N_15399,N_15305);
or U15712 (N_15712,N_15540,N_15566);
or U15713 (N_15713,N_15325,N_15470);
nor U15714 (N_15714,N_15594,N_15522);
nor U15715 (N_15715,N_15502,N_15517);
xnor U15716 (N_15716,N_15355,N_15308);
and U15717 (N_15717,N_15503,N_15430);
or U15718 (N_15718,N_15440,N_15555);
nor U15719 (N_15719,N_15536,N_15593);
xor U15720 (N_15720,N_15535,N_15384);
xor U15721 (N_15721,N_15494,N_15599);
or U15722 (N_15722,N_15340,N_15584);
nor U15723 (N_15723,N_15389,N_15337);
and U15724 (N_15724,N_15538,N_15310);
xnor U15725 (N_15725,N_15533,N_15327);
nor U15726 (N_15726,N_15598,N_15576);
xor U15727 (N_15727,N_15578,N_15489);
and U15728 (N_15728,N_15585,N_15428);
or U15729 (N_15729,N_15420,N_15439);
or U15730 (N_15730,N_15499,N_15366);
and U15731 (N_15731,N_15412,N_15380);
nor U15732 (N_15732,N_15441,N_15357);
or U15733 (N_15733,N_15429,N_15531);
nor U15734 (N_15734,N_15442,N_15402);
and U15735 (N_15735,N_15352,N_15466);
nor U15736 (N_15736,N_15557,N_15391);
or U15737 (N_15737,N_15300,N_15464);
nor U15738 (N_15738,N_15421,N_15546);
xor U15739 (N_15739,N_15373,N_15410);
nor U15740 (N_15740,N_15393,N_15449);
nor U15741 (N_15741,N_15396,N_15572);
xor U15742 (N_15742,N_15339,N_15330);
and U15743 (N_15743,N_15582,N_15342);
nand U15744 (N_15744,N_15455,N_15506);
nand U15745 (N_15745,N_15482,N_15551);
or U15746 (N_15746,N_15567,N_15478);
nand U15747 (N_15747,N_15457,N_15597);
xnor U15748 (N_15748,N_15471,N_15571);
xnor U15749 (N_15749,N_15318,N_15456);
xor U15750 (N_15750,N_15441,N_15375);
or U15751 (N_15751,N_15419,N_15411);
and U15752 (N_15752,N_15366,N_15488);
nand U15753 (N_15753,N_15327,N_15578);
nand U15754 (N_15754,N_15568,N_15360);
xnor U15755 (N_15755,N_15314,N_15454);
or U15756 (N_15756,N_15442,N_15312);
nor U15757 (N_15757,N_15564,N_15537);
xnor U15758 (N_15758,N_15342,N_15591);
or U15759 (N_15759,N_15385,N_15449);
xnor U15760 (N_15760,N_15494,N_15342);
xnor U15761 (N_15761,N_15399,N_15303);
nor U15762 (N_15762,N_15394,N_15461);
nor U15763 (N_15763,N_15573,N_15413);
xor U15764 (N_15764,N_15487,N_15304);
nor U15765 (N_15765,N_15591,N_15403);
xnor U15766 (N_15766,N_15364,N_15459);
and U15767 (N_15767,N_15341,N_15532);
and U15768 (N_15768,N_15397,N_15324);
nor U15769 (N_15769,N_15574,N_15475);
nor U15770 (N_15770,N_15538,N_15495);
or U15771 (N_15771,N_15579,N_15522);
nor U15772 (N_15772,N_15342,N_15531);
or U15773 (N_15773,N_15350,N_15387);
nor U15774 (N_15774,N_15539,N_15315);
xnor U15775 (N_15775,N_15595,N_15565);
nand U15776 (N_15776,N_15411,N_15433);
nand U15777 (N_15777,N_15367,N_15379);
xor U15778 (N_15778,N_15564,N_15588);
nor U15779 (N_15779,N_15398,N_15527);
nand U15780 (N_15780,N_15477,N_15599);
nand U15781 (N_15781,N_15433,N_15544);
nand U15782 (N_15782,N_15389,N_15378);
nand U15783 (N_15783,N_15407,N_15504);
and U15784 (N_15784,N_15317,N_15374);
xor U15785 (N_15785,N_15366,N_15337);
or U15786 (N_15786,N_15372,N_15305);
or U15787 (N_15787,N_15397,N_15589);
or U15788 (N_15788,N_15561,N_15498);
nand U15789 (N_15789,N_15325,N_15563);
and U15790 (N_15790,N_15322,N_15365);
and U15791 (N_15791,N_15306,N_15458);
xnor U15792 (N_15792,N_15477,N_15320);
xnor U15793 (N_15793,N_15479,N_15400);
nand U15794 (N_15794,N_15366,N_15394);
nor U15795 (N_15795,N_15413,N_15306);
xnor U15796 (N_15796,N_15552,N_15313);
nand U15797 (N_15797,N_15493,N_15503);
nand U15798 (N_15798,N_15343,N_15307);
nand U15799 (N_15799,N_15325,N_15466);
or U15800 (N_15800,N_15431,N_15453);
and U15801 (N_15801,N_15502,N_15584);
and U15802 (N_15802,N_15405,N_15408);
nor U15803 (N_15803,N_15495,N_15483);
nand U15804 (N_15804,N_15311,N_15354);
or U15805 (N_15805,N_15316,N_15527);
or U15806 (N_15806,N_15325,N_15592);
nor U15807 (N_15807,N_15580,N_15401);
xnor U15808 (N_15808,N_15446,N_15474);
or U15809 (N_15809,N_15444,N_15456);
xor U15810 (N_15810,N_15592,N_15310);
xor U15811 (N_15811,N_15329,N_15558);
and U15812 (N_15812,N_15431,N_15593);
xor U15813 (N_15813,N_15408,N_15470);
xnor U15814 (N_15814,N_15513,N_15350);
and U15815 (N_15815,N_15459,N_15354);
or U15816 (N_15816,N_15409,N_15502);
nor U15817 (N_15817,N_15337,N_15574);
nor U15818 (N_15818,N_15554,N_15376);
and U15819 (N_15819,N_15592,N_15366);
nand U15820 (N_15820,N_15409,N_15520);
xor U15821 (N_15821,N_15573,N_15589);
nand U15822 (N_15822,N_15308,N_15465);
and U15823 (N_15823,N_15314,N_15396);
xnor U15824 (N_15824,N_15438,N_15571);
nor U15825 (N_15825,N_15391,N_15409);
xnor U15826 (N_15826,N_15575,N_15579);
nand U15827 (N_15827,N_15425,N_15454);
and U15828 (N_15828,N_15340,N_15378);
and U15829 (N_15829,N_15489,N_15548);
or U15830 (N_15830,N_15421,N_15396);
nand U15831 (N_15831,N_15479,N_15446);
nor U15832 (N_15832,N_15540,N_15322);
or U15833 (N_15833,N_15355,N_15354);
or U15834 (N_15834,N_15317,N_15471);
and U15835 (N_15835,N_15574,N_15441);
and U15836 (N_15836,N_15426,N_15485);
xnor U15837 (N_15837,N_15356,N_15481);
xnor U15838 (N_15838,N_15324,N_15346);
or U15839 (N_15839,N_15385,N_15489);
nor U15840 (N_15840,N_15377,N_15567);
or U15841 (N_15841,N_15499,N_15547);
or U15842 (N_15842,N_15494,N_15406);
and U15843 (N_15843,N_15498,N_15510);
xnor U15844 (N_15844,N_15516,N_15489);
nor U15845 (N_15845,N_15540,N_15538);
or U15846 (N_15846,N_15577,N_15517);
and U15847 (N_15847,N_15379,N_15545);
xnor U15848 (N_15848,N_15413,N_15445);
xor U15849 (N_15849,N_15361,N_15388);
nor U15850 (N_15850,N_15525,N_15318);
nor U15851 (N_15851,N_15403,N_15435);
and U15852 (N_15852,N_15425,N_15576);
nor U15853 (N_15853,N_15446,N_15354);
nand U15854 (N_15854,N_15583,N_15421);
nand U15855 (N_15855,N_15442,N_15435);
or U15856 (N_15856,N_15355,N_15436);
xnor U15857 (N_15857,N_15365,N_15449);
and U15858 (N_15858,N_15487,N_15473);
nand U15859 (N_15859,N_15444,N_15599);
or U15860 (N_15860,N_15407,N_15484);
nor U15861 (N_15861,N_15385,N_15381);
nor U15862 (N_15862,N_15442,N_15475);
nand U15863 (N_15863,N_15517,N_15522);
nor U15864 (N_15864,N_15472,N_15380);
nor U15865 (N_15865,N_15525,N_15381);
or U15866 (N_15866,N_15572,N_15443);
nor U15867 (N_15867,N_15416,N_15447);
xnor U15868 (N_15868,N_15461,N_15587);
nand U15869 (N_15869,N_15324,N_15335);
or U15870 (N_15870,N_15444,N_15466);
nor U15871 (N_15871,N_15516,N_15470);
nand U15872 (N_15872,N_15454,N_15328);
nand U15873 (N_15873,N_15533,N_15464);
or U15874 (N_15874,N_15492,N_15498);
nand U15875 (N_15875,N_15454,N_15476);
xnor U15876 (N_15876,N_15369,N_15417);
or U15877 (N_15877,N_15403,N_15384);
or U15878 (N_15878,N_15354,N_15468);
or U15879 (N_15879,N_15565,N_15362);
nand U15880 (N_15880,N_15515,N_15520);
nor U15881 (N_15881,N_15389,N_15533);
nor U15882 (N_15882,N_15321,N_15508);
nand U15883 (N_15883,N_15546,N_15462);
nand U15884 (N_15884,N_15553,N_15430);
xor U15885 (N_15885,N_15518,N_15435);
xnor U15886 (N_15886,N_15446,N_15506);
nor U15887 (N_15887,N_15389,N_15319);
nand U15888 (N_15888,N_15592,N_15400);
nand U15889 (N_15889,N_15561,N_15364);
and U15890 (N_15890,N_15369,N_15466);
or U15891 (N_15891,N_15476,N_15524);
or U15892 (N_15892,N_15591,N_15457);
or U15893 (N_15893,N_15460,N_15464);
and U15894 (N_15894,N_15547,N_15489);
nand U15895 (N_15895,N_15463,N_15452);
nand U15896 (N_15896,N_15547,N_15302);
and U15897 (N_15897,N_15430,N_15392);
or U15898 (N_15898,N_15577,N_15530);
or U15899 (N_15899,N_15547,N_15478);
nor U15900 (N_15900,N_15889,N_15626);
nand U15901 (N_15901,N_15681,N_15818);
and U15902 (N_15902,N_15779,N_15638);
nor U15903 (N_15903,N_15734,N_15697);
and U15904 (N_15904,N_15744,N_15703);
nor U15905 (N_15905,N_15809,N_15774);
xnor U15906 (N_15906,N_15887,N_15643);
xor U15907 (N_15907,N_15775,N_15875);
xnor U15908 (N_15908,N_15789,N_15837);
and U15909 (N_15909,N_15784,N_15659);
nand U15910 (N_15910,N_15780,N_15896);
or U15911 (N_15911,N_15825,N_15814);
and U15912 (N_15912,N_15748,N_15606);
nand U15913 (N_15913,N_15854,N_15841);
nor U15914 (N_15914,N_15838,N_15604);
nor U15915 (N_15915,N_15639,N_15803);
nor U15916 (N_15916,N_15795,N_15674);
nand U15917 (N_15917,N_15759,N_15823);
and U15918 (N_15918,N_15762,N_15684);
nand U15919 (N_15919,N_15724,N_15696);
nor U15920 (N_15920,N_15673,N_15805);
nor U15921 (N_15921,N_15867,N_15702);
xnor U15922 (N_15922,N_15735,N_15758);
and U15923 (N_15923,N_15622,N_15753);
xnor U15924 (N_15924,N_15699,N_15811);
xnor U15925 (N_15925,N_15757,N_15876);
nand U15926 (N_15926,N_15881,N_15668);
xor U15927 (N_15927,N_15806,N_15650);
or U15928 (N_15928,N_15882,N_15609);
and U15929 (N_15929,N_15851,N_15798);
nor U15930 (N_15930,N_15897,N_15625);
nor U15931 (N_15931,N_15615,N_15676);
nand U15932 (N_15932,N_15869,N_15866);
and U15933 (N_15933,N_15862,N_15726);
or U15934 (N_15934,N_15847,N_15729);
or U15935 (N_15935,N_15692,N_15821);
xor U15936 (N_15936,N_15750,N_15845);
nor U15937 (N_15937,N_15898,N_15688);
and U15938 (N_15938,N_15716,N_15880);
xnor U15939 (N_15939,N_15655,N_15623);
or U15940 (N_15940,N_15679,N_15834);
nor U15941 (N_15941,N_15683,N_15883);
and U15942 (N_15942,N_15741,N_15830);
and U15943 (N_15943,N_15872,N_15733);
xnor U15944 (N_15944,N_15871,N_15717);
nor U15945 (N_15945,N_15754,N_15852);
or U15946 (N_15946,N_15819,N_15644);
and U15947 (N_15947,N_15800,N_15893);
nand U15948 (N_15948,N_15895,N_15611);
or U15949 (N_15949,N_15778,N_15846);
and U15950 (N_15950,N_15794,N_15853);
xnor U15951 (N_15951,N_15664,N_15810);
xnor U15952 (N_15952,N_15621,N_15892);
or U15953 (N_15953,N_15685,N_15894);
nor U15954 (N_15954,N_15785,N_15720);
xor U15955 (N_15955,N_15879,N_15788);
nor U15956 (N_15956,N_15637,N_15689);
xnor U15957 (N_15957,N_15817,N_15860);
and U15958 (N_15958,N_15614,N_15767);
nor U15959 (N_15959,N_15712,N_15861);
nor U15960 (N_15960,N_15740,N_15660);
nor U15961 (N_15961,N_15768,N_15886);
nor U15962 (N_15962,N_15840,N_15640);
nor U15963 (N_15963,N_15612,N_15705);
xor U15964 (N_15964,N_15687,N_15710);
and U15965 (N_15965,N_15829,N_15770);
xnor U15966 (N_15966,N_15796,N_15730);
nor U15967 (N_15967,N_15738,N_15630);
nor U15968 (N_15968,N_15657,N_15844);
xor U15969 (N_15969,N_15843,N_15833);
and U15970 (N_15970,N_15694,N_15736);
and U15971 (N_15971,N_15781,N_15666);
and U15972 (N_15972,N_15827,N_15864);
xnor U15973 (N_15973,N_15603,N_15773);
and U15974 (N_15974,N_15715,N_15619);
nand U15975 (N_15975,N_15764,N_15749);
and U15976 (N_15976,N_15665,N_15891);
nor U15977 (N_15977,N_15701,N_15792);
and U15978 (N_15978,N_15824,N_15783);
xor U15979 (N_15979,N_15826,N_15835);
xnor U15980 (N_15980,N_15627,N_15799);
or U15981 (N_15981,N_15690,N_15634);
or U15982 (N_15982,N_15731,N_15686);
nor U15983 (N_15983,N_15760,N_15601);
nor U15984 (N_15984,N_15877,N_15763);
or U15985 (N_15985,N_15878,N_15610);
nor U15986 (N_15986,N_15870,N_15616);
nand U15987 (N_15987,N_15698,N_15801);
and U15988 (N_15988,N_15797,N_15747);
nand U15989 (N_15989,N_15863,N_15714);
and U15990 (N_15990,N_15865,N_15808);
and U15991 (N_15991,N_15761,N_15742);
and U15992 (N_15992,N_15671,N_15802);
xor U15993 (N_15993,N_15654,N_15624);
and U15994 (N_15994,N_15857,N_15652);
or U15995 (N_15995,N_15719,N_15787);
nand U15996 (N_15996,N_15745,N_15790);
or U15997 (N_15997,N_15855,N_15766);
nand U15998 (N_15998,N_15678,N_15832);
nand U15999 (N_15999,N_15859,N_15771);
or U16000 (N_16000,N_15605,N_15663);
nand U16001 (N_16001,N_15617,N_15727);
xnor U16002 (N_16002,N_15658,N_15751);
or U16003 (N_16003,N_15728,N_15633);
nand U16004 (N_16004,N_15700,N_15618);
nand U16005 (N_16005,N_15725,N_15613);
xnor U16006 (N_16006,N_15884,N_15888);
nand U16007 (N_16007,N_15667,N_15756);
nand U16008 (N_16008,N_15856,N_15628);
xor U16009 (N_16009,N_15620,N_15691);
nand U16010 (N_16010,N_15722,N_15651);
nand U16011 (N_16011,N_15656,N_15642);
nor U16012 (N_16012,N_15723,N_15600);
nand U16013 (N_16013,N_15804,N_15670);
xor U16014 (N_16014,N_15890,N_15646);
and U16015 (N_16015,N_15706,N_15842);
or U16016 (N_16016,N_15677,N_15718);
nor U16017 (N_16017,N_15772,N_15831);
xnor U16018 (N_16018,N_15721,N_15873);
and U16019 (N_16019,N_15807,N_15839);
nand U16020 (N_16020,N_15708,N_15885);
and U16021 (N_16021,N_15669,N_15776);
and U16022 (N_16022,N_15899,N_15737);
xnor U16023 (N_16023,N_15791,N_15647);
and U16024 (N_16024,N_15693,N_15608);
xor U16025 (N_16025,N_15695,N_15675);
nor U16026 (N_16026,N_15661,N_15709);
and U16027 (N_16027,N_15793,N_15662);
xnor U16028 (N_16028,N_15711,N_15850);
nand U16029 (N_16029,N_15732,N_15649);
or U16030 (N_16030,N_15815,N_15858);
nand U16031 (N_16031,N_15641,N_15786);
or U16032 (N_16032,N_15822,N_15836);
or U16033 (N_16033,N_15812,N_15820);
xnor U16034 (N_16034,N_15782,N_15653);
and U16035 (N_16035,N_15874,N_15607);
or U16036 (N_16036,N_15765,N_15636);
nand U16037 (N_16037,N_15645,N_15704);
and U16038 (N_16038,N_15752,N_15602);
nand U16039 (N_16039,N_15755,N_15682);
nand U16040 (N_16040,N_15743,N_15868);
or U16041 (N_16041,N_15849,N_15631);
and U16042 (N_16042,N_15746,N_15813);
or U16043 (N_16043,N_15777,N_15648);
xor U16044 (N_16044,N_15848,N_15672);
nand U16045 (N_16045,N_15680,N_15629);
xnor U16046 (N_16046,N_15713,N_15828);
nor U16047 (N_16047,N_15769,N_15635);
nor U16048 (N_16048,N_15816,N_15707);
nand U16049 (N_16049,N_15739,N_15632);
and U16050 (N_16050,N_15694,N_15780);
nor U16051 (N_16051,N_15895,N_15742);
and U16052 (N_16052,N_15768,N_15854);
or U16053 (N_16053,N_15625,N_15603);
or U16054 (N_16054,N_15617,N_15796);
nand U16055 (N_16055,N_15756,N_15693);
nand U16056 (N_16056,N_15880,N_15878);
and U16057 (N_16057,N_15836,N_15672);
nor U16058 (N_16058,N_15867,N_15859);
nand U16059 (N_16059,N_15805,N_15715);
xor U16060 (N_16060,N_15898,N_15881);
nor U16061 (N_16061,N_15776,N_15796);
and U16062 (N_16062,N_15654,N_15736);
nor U16063 (N_16063,N_15795,N_15704);
nor U16064 (N_16064,N_15860,N_15889);
nor U16065 (N_16065,N_15775,N_15613);
or U16066 (N_16066,N_15786,N_15819);
nand U16067 (N_16067,N_15750,N_15875);
nor U16068 (N_16068,N_15693,N_15604);
or U16069 (N_16069,N_15828,N_15623);
xor U16070 (N_16070,N_15648,N_15638);
and U16071 (N_16071,N_15885,N_15859);
xor U16072 (N_16072,N_15690,N_15601);
xor U16073 (N_16073,N_15768,N_15873);
xor U16074 (N_16074,N_15721,N_15735);
nand U16075 (N_16075,N_15893,N_15810);
and U16076 (N_16076,N_15614,N_15831);
and U16077 (N_16077,N_15766,N_15862);
or U16078 (N_16078,N_15898,N_15667);
xor U16079 (N_16079,N_15606,N_15648);
nand U16080 (N_16080,N_15717,N_15833);
nand U16081 (N_16081,N_15797,N_15825);
or U16082 (N_16082,N_15799,N_15899);
or U16083 (N_16083,N_15686,N_15863);
nor U16084 (N_16084,N_15832,N_15686);
nand U16085 (N_16085,N_15646,N_15627);
nor U16086 (N_16086,N_15830,N_15686);
nand U16087 (N_16087,N_15705,N_15786);
and U16088 (N_16088,N_15870,N_15784);
nand U16089 (N_16089,N_15700,N_15669);
and U16090 (N_16090,N_15820,N_15804);
xor U16091 (N_16091,N_15881,N_15656);
xor U16092 (N_16092,N_15861,N_15627);
or U16093 (N_16093,N_15834,N_15712);
and U16094 (N_16094,N_15752,N_15887);
xor U16095 (N_16095,N_15653,N_15815);
nor U16096 (N_16096,N_15745,N_15784);
xor U16097 (N_16097,N_15845,N_15770);
and U16098 (N_16098,N_15653,N_15674);
nor U16099 (N_16099,N_15778,N_15601);
xnor U16100 (N_16100,N_15834,N_15659);
nand U16101 (N_16101,N_15621,N_15836);
nand U16102 (N_16102,N_15764,N_15729);
nor U16103 (N_16103,N_15821,N_15643);
xor U16104 (N_16104,N_15625,N_15658);
nor U16105 (N_16105,N_15721,N_15702);
or U16106 (N_16106,N_15884,N_15769);
or U16107 (N_16107,N_15707,N_15738);
nor U16108 (N_16108,N_15703,N_15814);
or U16109 (N_16109,N_15852,N_15660);
and U16110 (N_16110,N_15824,N_15752);
nand U16111 (N_16111,N_15668,N_15750);
nor U16112 (N_16112,N_15668,N_15820);
or U16113 (N_16113,N_15612,N_15863);
nor U16114 (N_16114,N_15803,N_15899);
or U16115 (N_16115,N_15788,N_15736);
xnor U16116 (N_16116,N_15886,N_15703);
nand U16117 (N_16117,N_15772,N_15672);
xnor U16118 (N_16118,N_15770,N_15603);
nand U16119 (N_16119,N_15610,N_15628);
nand U16120 (N_16120,N_15863,N_15755);
and U16121 (N_16121,N_15840,N_15629);
nand U16122 (N_16122,N_15640,N_15606);
nand U16123 (N_16123,N_15817,N_15897);
nand U16124 (N_16124,N_15867,N_15724);
nor U16125 (N_16125,N_15864,N_15652);
or U16126 (N_16126,N_15680,N_15893);
nand U16127 (N_16127,N_15622,N_15800);
nand U16128 (N_16128,N_15857,N_15749);
nand U16129 (N_16129,N_15689,N_15890);
or U16130 (N_16130,N_15799,N_15730);
or U16131 (N_16131,N_15658,N_15732);
nand U16132 (N_16132,N_15790,N_15773);
xor U16133 (N_16133,N_15735,N_15849);
xor U16134 (N_16134,N_15869,N_15628);
nand U16135 (N_16135,N_15808,N_15768);
and U16136 (N_16136,N_15602,N_15832);
and U16137 (N_16137,N_15668,N_15614);
xnor U16138 (N_16138,N_15766,N_15685);
or U16139 (N_16139,N_15734,N_15798);
or U16140 (N_16140,N_15865,N_15836);
xnor U16141 (N_16141,N_15732,N_15619);
or U16142 (N_16142,N_15652,N_15659);
or U16143 (N_16143,N_15757,N_15788);
nor U16144 (N_16144,N_15617,N_15777);
xor U16145 (N_16145,N_15811,N_15602);
nor U16146 (N_16146,N_15806,N_15770);
or U16147 (N_16147,N_15810,N_15628);
and U16148 (N_16148,N_15783,N_15813);
and U16149 (N_16149,N_15641,N_15752);
or U16150 (N_16150,N_15602,N_15860);
xnor U16151 (N_16151,N_15786,N_15815);
or U16152 (N_16152,N_15681,N_15828);
xnor U16153 (N_16153,N_15677,N_15889);
nand U16154 (N_16154,N_15628,N_15758);
nand U16155 (N_16155,N_15891,N_15893);
nor U16156 (N_16156,N_15660,N_15604);
xor U16157 (N_16157,N_15859,N_15667);
or U16158 (N_16158,N_15821,N_15779);
or U16159 (N_16159,N_15771,N_15633);
nand U16160 (N_16160,N_15638,N_15823);
nor U16161 (N_16161,N_15656,N_15694);
nand U16162 (N_16162,N_15692,N_15853);
nor U16163 (N_16163,N_15634,N_15660);
nor U16164 (N_16164,N_15623,N_15771);
or U16165 (N_16165,N_15808,N_15657);
and U16166 (N_16166,N_15680,N_15782);
nand U16167 (N_16167,N_15757,N_15773);
nand U16168 (N_16168,N_15641,N_15710);
or U16169 (N_16169,N_15800,N_15640);
nand U16170 (N_16170,N_15692,N_15747);
nand U16171 (N_16171,N_15889,N_15855);
nor U16172 (N_16172,N_15730,N_15609);
or U16173 (N_16173,N_15669,N_15741);
and U16174 (N_16174,N_15755,N_15700);
or U16175 (N_16175,N_15756,N_15793);
nor U16176 (N_16176,N_15892,N_15894);
and U16177 (N_16177,N_15682,N_15706);
or U16178 (N_16178,N_15711,N_15689);
nor U16179 (N_16179,N_15839,N_15850);
nor U16180 (N_16180,N_15842,N_15739);
nand U16181 (N_16181,N_15883,N_15638);
nor U16182 (N_16182,N_15814,N_15735);
nand U16183 (N_16183,N_15800,N_15727);
xor U16184 (N_16184,N_15767,N_15688);
and U16185 (N_16185,N_15733,N_15602);
nor U16186 (N_16186,N_15672,N_15806);
nand U16187 (N_16187,N_15884,N_15840);
xnor U16188 (N_16188,N_15882,N_15722);
xnor U16189 (N_16189,N_15828,N_15873);
or U16190 (N_16190,N_15812,N_15725);
or U16191 (N_16191,N_15832,N_15860);
xor U16192 (N_16192,N_15772,N_15730);
xor U16193 (N_16193,N_15817,N_15623);
nor U16194 (N_16194,N_15852,N_15746);
nor U16195 (N_16195,N_15654,N_15828);
xor U16196 (N_16196,N_15787,N_15717);
and U16197 (N_16197,N_15732,N_15774);
or U16198 (N_16198,N_15663,N_15877);
xor U16199 (N_16199,N_15624,N_15673);
nand U16200 (N_16200,N_16087,N_16181);
xnor U16201 (N_16201,N_15919,N_15987);
nand U16202 (N_16202,N_16140,N_16005);
nor U16203 (N_16203,N_16141,N_16178);
and U16204 (N_16204,N_15940,N_16164);
nand U16205 (N_16205,N_16157,N_16028);
nand U16206 (N_16206,N_15944,N_15950);
or U16207 (N_16207,N_16009,N_16018);
or U16208 (N_16208,N_15908,N_16037);
xor U16209 (N_16209,N_15920,N_16114);
nand U16210 (N_16210,N_16046,N_16136);
or U16211 (N_16211,N_16022,N_16083);
or U16212 (N_16212,N_16034,N_16045);
nor U16213 (N_16213,N_15947,N_15985);
or U16214 (N_16214,N_15982,N_15956);
or U16215 (N_16215,N_16082,N_16002);
nand U16216 (N_16216,N_16121,N_16161);
nor U16217 (N_16217,N_15939,N_16133);
xor U16218 (N_16218,N_16016,N_16049);
xor U16219 (N_16219,N_16126,N_16090);
and U16220 (N_16220,N_15998,N_16198);
xor U16221 (N_16221,N_15922,N_16112);
nor U16222 (N_16222,N_16061,N_15931);
or U16223 (N_16223,N_16148,N_16053);
nor U16224 (N_16224,N_16174,N_15973);
nor U16225 (N_16225,N_16194,N_15986);
nand U16226 (N_16226,N_16130,N_16123);
nor U16227 (N_16227,N_16066,N_16195);
nand U16228 (N_16228,N_16150,N_15995);
and U16229 (N_16229,N_16055,N_15914);
or U16230 (N_16230,N_15990,N_16173);
and U16231 (N_16231,N_16091,N_16145);
nor U16232 (N_16232,N_16047,N_15925);
and U16233 (N_16233,N_16056,N_16026);
or U16234 (N_16234,N_16187,N_15984);
nor U16235 (N_16235,N_16007,N_16072);
or U16236 (N_16236,N_16168,N_16177);
or U16237 (N_16237,N_15954,N_16064);
or U16238 (N_16238,N_15941,N_16192);
xnor U16239 (N_16239,N_15911,N_15909);
nor U16240 (N_16240,N_16184,N_16176);
xnor U16241 (N_16241,N_15994,N_16020);
nor U16242 (N_16242,N_16149,N_15942);
and U16243 (N_16243,N_16107,N_16079);
nor U16244 (N_16244,N_16078,N_15946);
nor U16245 (N_16245,N_16180,N_16154);
or U16246 (N_16246,N_16120,N_16160);
xor U16247 (N_16247,N_16131,N_15933);
nor U16248 (N_16248,N_15921,N_15943);
xnor U16249 (N_16249,N_15905,N_15955);
xnor U16250 (N_16250,N_15978,N_16115);
xor U16251 (N_16251,N_15927,N_15977);
nor U16252 (N_16252,N_16013,N_15913);
or U16253 (N_16253,N_16127,N_16146);
xor U16254 (N_16254,N_16170,N_15976);
or U16255 (N_16255,N_15961,N_15930);
xor U16256 (N_16256,N_15962,N_16128);
xor U16257 (N_16257,N_16081,N_15929);
xor U16258 (N_16258,N_15970,N_15964);
xor U16259 (N_16259,N_15952,N_16100);
nand U16260 (N_16260,N_16191,N_15980);
xnor U16261 (N_16261,N_16105,N_16035);
xnor U16262 (N_16262,N_16175,N_15917);
and U16263 (N_16263,N_16033,N_15900);
nor U16264 (N_16264,N_15901,N_16113);
xor U16265 (N_16265,N_16186,N_16092);
or U16266 (N_16266,N_16076,N_16104);
or U16267 (N_16267,N_16137,N_16074);
xor U16268 (N_16268,N_15992,N_16185);
xor U16269 (N_16269,N_16004,N_15949);
or U16270 (N_16270,N_16118,N_15989);
or U16271 (N_16271,N_16065,N_16089);
xor U16272 (N_16272,N_16196,N_16166);
nand U16273 (N_16273,N_16162,N_16155);
nand U16274 (N_16274,N_16071,N_16108);
xnor U16275 (N_16275,N_16171,N_15958);
xor U16276 (N_16276,N_16197,N_15932);
xnor U16277 (N_16277,N_15966,N_15971);
xor U16278 (N_16278,N_16179,N_15934);
or U16279 (N_16279,N_15903,N_16101);
xnor U16280 (N_16280,N_15945,N_16156);
and U16281 (N_16281,N_16017,N_16096);
and U16282 (N_16282,N_15948,N_15979);
nor U16283 (N_16283,N_16099,N_15915);
or U16284 (N_16284,N_15972,N_16051);
xnor U16285 (N_16285,N_16000,N_16152);
or U16286 (N_16286,N_15928,N_16031);
nor U16287 (N_16287,N_15960,N_16159);
and U16288 (N_16288,N_16019,N_16106);
nand U16289 (N_16289,N_15907,N_15988);
and U16290 (N_16290,N_15926,N_16098);
and U16291 (N_16291,N_16036,N_15983);
or U16292 (N_16292,N_15910,N_16058);
or U16293 (N_16293,N_16023,N_16097);
nand U16294 (N_16294,N_16163,N_16015);
xnor U16295 (N_16295,N_16085,N_15924);
nor U16296 (N_16296,N_16062,N_15999);
nor U16297 (N_16297,N_15993,N_16042);
xor U16298 (N_16298,N_15975,N_16080);
nand U16299 (N_16299,N_16129,N_16093);
and U16300 (N_16300,N_15981,N_16029);
xnor U16301 (N_16301,N_15906,N_16103);
or U16302 (N_16302,N_16068,N_16025);
or U16303 (N_16303,N_16088,N_16094);
nand U16304 (N_16304,N_16167,N_16199);
and U16305 (N_16305,N_16038,N_15959);
nor U16306 (N_16306,N_15902,N_15997);
and U16307 (N_16307,N_16117,N_16084);
xor U16308 (N_16308,N_16139,N_16169);
nand U16309 (N_16309,N_16153,N_16183);
or U16310 (N_16310,N_16014,N_16142);
and U16311 (N_16311,N_15935,N_16032);
xor U16312 (N_16312,N_16021,N_15965);
nor U16313 (N_16313,N_16122,N_16003);
or U16314 (N_16314,N_16151,N_16111);
or U16315 (N_16315,N_16102,N_15968);
or U16316 (N_16316,N_15937,N_16024);
and U16317 (N_16317,N_16012,N_16041);
and U16318 (N_16318,N_16010,N_16075);
or U16319 (N_16319,N_15967,N_16132);
xnor U16320 (N_16320,N_16135,N_16172);
and U16321 (N_16321,N_16050,N_15991);
nand U16322 (N_16322,N_16143,N_15957);
or U16323 (N_16323,N_15953,N_16189);
nand U16324 (N_16324,N_15996,N_16124);
nand U16325 (N_16325,N_16086,N_15918);
xor U16326 (N_16326,N_16067,N_16125);
or U16327 (N_16327,N_16109,N_16059);
or U16328 (N_16328,N_16039,N_16043);
xor U16329 (N_16329,N_16060,N_15969);
nor U16330 (N_16330,N_16008,N_16011);
and U16331 (N_16331,N_15936,N_15904);
or U16332 (N_16332,N_16001,N_15963);
nor U16333 (N_16333,N_16048,N_16138);
and U16334 (N_16334,N_16057,N_16188);
and U16335 (N_16335,N_16110,N_16165);
and U16336 (N_16336,N_16119,N_16027);
or U16337 (N_16337,N_16158,N_16147);
xor U16338 (N_16338,N_16052,N_16069);
and U16339 (N_16339,N_16054,N_16144);
and U16340 (N_16340,N_15923,N_16063);
nand U16341 (N_16341,N_15974,N_15951);
and U16342 (N_16342,N_15912,N_16030);
nand U16343 (N_16343,N_16073,N_16044);
or U16344 (N_16344,N_16040,N_16116);
xnor U16345 (N_16345,N_16193,N_16134);
nor U16346 (N_16346,N_15916,N_16006);
nor U16347 (N_16347,N_16070,N_16077);
or U16348 (N_16348,N_16190,N_16095);
nand U16349 (N_16349,N_15938,N_16182);
nor U16350 (N_16350,N_16130,N_15960);
or U16351 (N_16351,N_16179,N_16057);
and U16352 (N_16352,N_16076,N_16026);
or U16353 (N_16353,N_15988,N_16068);
or U16354 (N_16354,N_16149,N_15970);
xor U16355 (N_16355,N_16063,N_16190);
or U16356 (N_16356,N_15986,N_15970);
or U16357 (N_16357,N_16189,N_15919);
nand U16358 (N_16358,N_16005,N_16191);
xor U16359 (N_16359,N_16187,N_16098);
xnor U16360 (N_16360,N_16030,N_15971);
nor U16361 (N_16361,N_16022,N_16102);
or U16362 (N_16362,N_16048,N_15949);
nor U16363 (N_16363,N_16010,N_15909);
xor U16364 (N_16364,N_16066,N_15911);
or U16365 (N_16365,N_16183,N_15979);
xnor U16366 (N_16366,N_16027,N_16144);
nand U16367 (N_16367,N_15931,N_16122);
nand U16368 (N_16368,N_15901,N_16137);
nand U16369 (N_16369,N_15922,N_15998);
nor U16370 (N_16370,N_15923,N_15971);
nor U16371 (N_16371,N_16190,N_15916);
nor U16372 (N_16372,N_16105,N_16189);
and U16373 (N_16373,N_16116,N_16145);
nor U16374 (N_16374,N_16010,N_16179);
xor U16375 (N_16375,N_16008,N_15935);
or U16376 (N_16376,N_15962,N_15933);
nand U16377 (N_16377,N_16194,N_16124);
or U16378 (N_16378,N_16068,N_16178);
nand U16379 (N_16379,N_16100,N_16134);
and U16380 (N_16380,N_16020,N_16061);
and U16381 (N_16381,N_16062,N_15926);
and U16382 (N_16382,N_16043,N_15958);
xor U16383 (N_16383,N_16101,N_16088);
and U16384 (N_16384,N_15927,N_15939);
nor U16385 (N_16385,N_15990,N_16150);
xnor U16386 (N_16386,N_16108,N_15915);
nor U16387 (N_16387,N_16011,N_15924);
xor U16388 (N_16388,N_15942,N_16177);
nand U16389 (N_16389,N_16019,N_15922);
and U16390 (N_16390,N_16094,N_15964);
or U16391 (N_16391,N_16006,N_16115);
nor U16392 (N_16392,N_16129,N_16053);
or U16393 (N_16393,N_15905,N_16199);
and U16394 (N_16394,N_16077,N_16128);
nand U16395 (N_16395,N_15932,N_16023);
or U16396 (N_16396,N_16195,N_16141);
nand U16397 (N_16397,N_16166,N_16194);
xor U16398 (N_16398,N_16026,N_16163);
and U16399 (N_16399,N_15953,N_16171);
nand U16400 (N_16400,N_16119,N_16185);
nand U16401 (N_16401,N_16188,N_16183);
nor U16402 (N_16402,N_16172,N_16100);
xor U16403 (N_16403,N_16014,N_16197);
nor U16404 (N_16404,N_15961,N_15928);
xnor U16405 (N_16405,N_16042,N_15964);
nor U16406 (N_16406,N_16122,N_15944);
and U16407 (N_16407,N_16095,N_15946);
and U16408 (N_16408,N_15970,N_16185);
nor U16409 (N_16409,N_16150,N_16050);
nor U16410 (N_16410,N_16057,N_16083);
and U16411 (N_16411,N_15938,N_16131);
nand U16412 (N_16412,N_15991,N_16105);
nand U16413 (N_16413,N_16100,N_16040);
xor U16414 (N_16414,N_16186,N_16134);
or U16415 (N_16415,N_16136,N_16194);
nor U16416 (N_16416,N_15957,N_15927);
nor U16417 (N_16417,N_16040,N_15962);
and U16418 (N_16418,N_16078,N_15928);
nor U16419 (N_16419,N_16070,N_16194);
xnor U16420 (N_16420,N_15934,N_15981);
xnor U16421 (N_16421,N_16095,N_16193);
and U16422 (N_16422,N_15956,N_16036);
nor U16423 (N_16423,N_16144,N_15927);
or U16424 (N_16424,N_15963,N_16151);
nand U16425 (N_16425,N_16148,N_16098);
or U16426 (N_16426,N_16080,N_15968);
nor U16427 (N_16427,N_16085,N_15971);
nand U16428 (N_16428,N_15945,N_16199);
or U16429 (N_16429,N_15906,N_15930);
nand U16430 (N_16430,N_15990,N_16041);
nand U16431 (N_16431,N_16183,N_16053);
or U16432 (N_16432,N_15988,N_15962);
and U16433 (N_16433,N_16173,N_15907);
and U16434 (N_16434,N_16174,N_16176);
and U16435 (N_16435,N_16140,N_16168);
or U16436 (N_16436,N_16031,N_15936);
and U16437 (N_16437,N_15978,N_16150);
and U16438 (N_16438,N_15906,N_16078);
xor U16439 (N_16439,N_15937,N_16169);
nand U16440 (N_16440,N_16160,N_16197);
nand U16441 (N_16441,N_15974,N_16131);
nand U16442 (N_16442,N_16092,N_16093);
or U16443 (N_16443,N_15997,N_15943);
or U16444 (N_16444,N_16197,N_16103);
nor U16445 (N_16445,N_15912,N_15982);
or U16446 (N_16446,N_15984,N_16086);
nand U16447 (N_16447,N_16083,N_16098);
xnor U16448 (N_16448,N_16104,N_15925);
or U16449 (N_16449,N_15975,N_16092);
or U16450 (N_16450,N_16148,N_16181);
or U16451 (N_16451,N_16076,N_15992);
xor U16452 (N_16452,N_16113,N_16143);
nor U16453 (N_16453,N_15913,N_16158);
xnor U16454 (N_16454,N_16118,N_15932);
or U16455 (N_16455,N_16063,N_16113);
and U16456 (N_16456,N_16009,N_16178);
nor U16457 (N_16457,N_16184,N_16150);
nor U16458 (N_16458,N_16077,N_15979);
nor U16459 (N_16459,N_16152,N_15954);
or U16460 (N_16460,N_16070,N_15979);
nor U16461 (N_16461,N_15972,N_16176);
nand U16462 (N_16462,N_16021,N_16059);
nand U16463 (N_16463,N_16107,N_16004);
and U16464 (N_16464,N_16134,N_16183);
xnor U16465 (N_16465,N_15945,N_16129);
or U16466 (N_16466,N_15976,N_16086);
and U16467 (N_16467,N_16184,N_16157);
or U16468 (N_16468,N_15963,N_16162);
nand U16469 (N_16469,N_16152,N_15938);
or U16470 (N_16470,N_15971,N_16045);
and U16471 (N_16471,N_16032,N_16140);
or U16472 (N_16472,N_16011,N_16140);
xnor U16473 (N_16473,N_16042,N_15931);
or U16474 (N_16474,N_16017,N_16135);
nor U16475 (N_16475,N_16099,N_16156);
nand U16476 (N_16476,N_16058,N_15998);
or U16477 (N_16477,N_15985,N_16066);
and U16478 (N_16478,N_16124,N_16067);
or U16479 (N_16479,N_15994,N_16075);
and U16480 (N_16480,N_16061,N_16093);
and U16481 (N_16481,N_15957,N_15988);
nor U16482 (N_16482,N_15911,N_15913);
nor U16483 (N_16483,N_16080,N_16104);
xnor U16484 (N_16484,N_15997,N_15956);
nand U16485 (N_16485,N_16141,N_16139);
xnor U16486 (N_16486,N_16197,N_16175);
or U16487 (N_16487,N_16137,N_15907);
nor U16488 (N_16488,N_16151,N_16037);
nand U16489 (N_16489,N_16190,N_16093);
nor U16490 (N_16490,N_16040,N_15933);
nand U16491 (N_16491,N_16191,N_15966);
or U16492 (N_16492,N_15931,N_16028);
and U16493 (N_16493,N_16054,N_16074);
nor U16494 (N_16494,N_16049,N_15932);
xor U16495 (N_16495,N_16118,N_15999);
xor U16496 (N_16496,N_16051,N_16116);
nand U16497 (N_16497,N_16003,N_16084);
and U16498 (N_16498,N_15918,N_16091);
or U16499 (N_16499,N_16137,N_16092);
and U16500 (N_16500,N_16368,N_16372);
and U16501 (N_16501,N_16376,N_16389);
nor U16502 (N_16502,N_16377,N_16499);
nand U16503 (N_16503,N_16293,N_16450);
nand U16504 (N_16504,N_16347,N_16215);
xnor U16505 (N_16505,N_16423,N_16221);
nand U16506 (N_16506,N_16283,N_16463);
or U16507 (N_16507,N_16470,N_16395);
nand U16508 (N_16508,N_16338,N_16278);
xnor U16509 (N_16509,N_16286,N_16440);
and U16510 (N_16510,N_16254,N_16447);
xnor U16511 (N_16511,N_16219,N_16412);
nor U16512 (N_16512,N_16252,N_16358);
nor U16513 (N_16513,N_16245,N_16392);
or U16514 (N_16514,N_16437,N_16336);
or U16515 (N_16515,N_16279,N_16244);
and U16516 (N_16516,N_16481,N_16260);
nor U16517 (N_16517,N_16402,N_16489);
or U16518 (N_16518,N_16307,N_16271);
nor U16519 (N_16519,N_16255,N_16427);
nand U16520 (N_16520,N_16216,N_16299);
nand U16521 (N_16521,N_16453,N_16291);
xnor U16522 (N_16522,N_16249,N_16426);
xor U16523 (N_16523,N_16310,N_16485);
and U16524 (N_16524,N_16359,N_16436);
and U16525 (N_16525,N_16298,N_16212);
nor U16526 (N_16526,N_16403,N_16401);
nor U16527 (N_16527,N_16380,N_16367);
or U16528 (N_16528,N_16251,N_16445);
xor U16529 (N_16529,N_16465,N_16207);
or U16530 (N_16530,N_16237,N_16248);
and U16531 (N_16531,N_16408,N_16296);
nor U16532 (N_16532,N_16231,N_16210);
and U16533 (N_16533,N_16461,N_16486);
and U16534 (N_16534,N_16354,N_16484);
and U16535 (N_16535,N_16451,N_16315);
nor U16536 (N_16536,N_16333,N_16295);
nor U16537 (N_16537,N_16261,N_16438);
nand U16538 (N_16538,N_16200,N_16236);
or U16539 (N_16539,N_16439,N_16474);
nand U16540 (N_16540,N_16473,N_16327);
and U16541 (N_16541,N_16430,N_16243);
or U16542 (N_16542,N_16280,N_16443);
nand U16543 (N_16543,N_16203,N_16258);
nor U16544 (N_16544,N_16329,N_16362);
xor U16545 (N_16545,N_16407,N_16413);
xor U16546 (N_16546,N_16361,N_16356);
nand U16547 (N_16547,N_16272,N_16240);
nor U16548 (N_16548,N_16391,N_16218);
nand U16549 (N_16549,N_16331,N_16444);
nand U16550 (N_16550,N_16388,N_16224);
and U16551 (N_16551,N_16289,N_16211);
nand U16552 (N_16552,N_16263,N_16350);
and U16553 (N_16553,N_16234,N_16220);
xnor U16554 (N_16554,N_16309,N_16222);
nand U16555 (N_16555,N_16337,N_16351);
or U16556 (N_16556,N_16277,N_16202);
nand U16557 (N_16557,N_16483,N_16441);
nor U16558 (N_16558,N_16232,N_16493);
nor U16559 (N_16559,N_16382,N_16267);
nand U16560 (N_16560,N_16454,N_16320);
or U16561 (N_16561,N_16206,N_16459);
nor U16562 (N_16562,N_16415,N_16287);
or U16563 (N_16563,N_16400,N_16214);
xor U16564 (N_16564,N_16326,N_16482);
nand U16565 (N_16565,N_16213,N_16360);
and U16566 (N_16566,N_16322,N_16328);
or U16567 (N_16567,N_16209,N_16406);
xnor U16568 (N_16568,N_16311,N_16330);
nand U16569 (N_16569,N_16448,N_16418);
nor U16570 (N_16570,N_16273,N_16480);
xor U16571 (N_16571,N_16313,N_16469);
xor U16572 (N_16572,N_16306,N_16494);
and U16573 (N_16573,N_16409,N_16371);
nor U16574 (N_16574,N_16312,N_16281);
xor U16575 (N_16575,N_16208,N_16460);
or U16576 (N_16576,N_16446,N_16365);
nand U16577 (N_16577,N_16345,N_16458);
nor U16578 (N_16578,N_16225,N_16227);
nor U16579 (N_16579,N_16364,N_16300);
xor U16580 (N_16580,N_16270,N_16471);
nor U16581 (N_16581,N_16269,N_16332);
nor U16582 (N_16582,N_16246,N_16325);
or U16583 (N_16583,N_16229,N_16226);
nor U16584 (N_16584,N_16339,N_16488);
and U16585 (N_16585,N_16414,N_16301);
nor U16586 (N_16586,N_16290,N_16265);
and U16587 (N_16587,N_16398,N_16321);
or U16588 (N_16588,N_16434,N_16496);
xnor U16589 (N_16589,N_16223,N_16428);
and U16590 (N_16590,N_16435,N_16383);
nand U16591 (N_16591,N_16264,N_16390);
nor U16592 (N_16592,N_16381,N_16355);
nor U16593 (N_16593,N_16204,N_16353);
nor U16594 (N_16594,N_16228,N_16343);
nand U16595 (N_16595,N_16495,N_16387);
nand U16596 (N_16596,N_16497,N_16262);
nor U16597 (N_16597,N_16449,N_16217);
xor U16598 (N_16598,N_16319,N_16314);
nor U16599 (N_16599,N_16274,N_16490);
xnor U16600 (N_16600,N_16304,N_16384);
or U16601 (N_16601,N_16373,N_16452);
xor U16602 (N_16602,N_16282,N_16472);
nand U16603 (N_16603,N_16346,N_16241);
and U16604 (N_16604,N_16285,N_16421);
nand U16605 (N_16605,N_16335,N_16467);
nand U16606 (N_16606,N_16477,N_16239);
xnor U16607 (N_16607,N_16344,N_16479);
nand U16608 (N_16608,N_16466,N_16462);
or U16609 (N_16609,N_16257,N_16334);
xor U16610 (N_16610,N_16242,N_16416);
or U16611 (N_16611,N_16491,N_16266);
xnor U16612 (N_16612,N_16316,N_16352);
or U16613 (N_16613,N_16375,N_16405);
nand U16614 (N_16614,N_16341,N_16230);
xor U16615 (N_16615,N_16288,N_16378);
and U16616 (N_16616,N_16292,N_16205);
nand U16617 (N_16617,N_16235,N_16420);
and U16618 (N_16618,N_16468,N_16284);
xnor U16619 (N_16619,N_16456,N_16308);
xnor U16620 (N_16620,N_16305,N_16429);
xnor U16621 (N_16621,N_16433,N_16268);
and U16622 (N_16622,N_16442,N_16492);
nand U16623 (N_16623,N_16317,N_16410);
nand U16624 (N_16624,N_16422,N_16393);
and U16625 (N_16625,N_16275,N_16404);
or U16626 (N_16626,N_16294,N_16318);
or U16627 (N_16627,N_16487,N_16379);
nand U16628 (N_16628,N_16349,N_16324);
nand U16629 (N_16629,N_16276,N_16386);
nand U16630 (N_16630,N_16302,N_16201);
nand U16631 (N_16631,N_16419,N_16363);
nor U16632 (N_16632,N_16478,N_16366);
and U16633 (N_16633,N_16476,N_16455);
or U16634 (N_16634,N_16411,N_16431);
or U16635 (N_16635,N_16498,N_16250);
nor U16636 (N_16636,N_16357,N_16417);
nand U16637 (N_16637,N_16342,N_16396);
and U16638 (N_16638,N_16340,N_16303);
nand U16639 (N_16639,N_16233,N_16348);
xnor U16640 (N_16640,N_16424,N_16247);
nand U16641 (N_16641,N_16256,N_16374);
nor U16642 (N_16642,N_16297,N_16432);
nand U16643 (N_16643,N_16425,N_16259);
or U16644 (N_16644,N_16238,N_16475);
xor U16645 (N_16645,N_16394,N_16397);
nand U16646 (N_16646,N_16457,N_16370);
or U16647 (N_16647,N_16464,N_16253);
nand U16648 (N_16648,N_16385,N_16323);
xor U16649 (N_16649,N_16399,N_16369);
nand U16650 (N_16650,N_16229,N_16491);
or U16651 (N_16651,N_16479,N_16221);
nand U16652 (N_16652,N_16216,N_16364);
and U16653 (N_16653,N_16265,N_16454);
and U16654 (N_16654,N_16336,N_16424);
xor U16655 (N_16655,N_16479,N_16367);
nor U16656 (N_16656,N_16352,N_16381);
and U16657 (N_16657,N_16315,N_16335);
or U16658 (N_16658,N_16204,N_16344);
nor U16659 (N_16659,N_16426,N_16375);
xor U16660 (N_16660,N_16405,N_16359);
nor U16661 (N_16661,N_16423,N_16420);
or U16662 (N_16662,N_16415,N_16271);
and U16663 (N_16663,N_16345,N_16411);
and U16664 (N_16664,N_16260,N_16326);
and U16665 (N_16665,N_16233,N_16224);
or U16666 (N_16666,N_16336,N_16413);
or U16667 (N_16667,N_16424,N_16314);
or U16668 (N_16668,N_16299,N_16366);
or U16669 (N_16669,N_16362,N_16261);
nand U16670 (N_16670,N_16205,N_16322);
and U16671 (N_16671,N_16346,N_16480);
and U16672 (N_16672,N_16463,N_16460);
or U16673 (N_16673,N_16489,N_16285);
nand U16674 (N_16674,N_16488,N_16209);
and U16675 (N_16675,N_16376,N_16309);
or U16676 (N_16676,N_16333,N_16471);
or U16677 (N_16677,N_16322,N_16377);
and U16678 (N_16678,N_16381,N_16475);
and U16679 (N_16679,N_16297,N_16329);
and U16680 (N_16680,N_16436,N_16316);
nor U16681 (N_16681,N_16399,N_16245);
nor U16682 (N_16682,N_16472,N_16397);
nor U16683 (N_16683,N_16380,N_16452);
and U16684 (N_16684,N_16325,N_16229);
xor U16685 (N_16685,N_16449,N_16411);
xnor U16686 (N_16686,N_16326,N_16422);
nand U16687 (N_16687,N_16488,N_16387);
nor U16688 (N_16688,N_16331,N_16309);
nor U16689 (N_16689,N_16374,N_16355);
nor U16690 (N_16690,N_16221,N_16422);
xor U16691 (N_16691,N_16201,N_16286);
or U16692 (N_16692,N_16428,N_16326);
and U16693 (N_16693,N_16256,N_16458);
xor U16694 (N_16694,N_16213,N_16396);
nand U16695 (N_16695,N_16438,N_16202);
or U16696 (N_16696,N_16419,N_16229);
or U16697 (N_16697,N_16417,N_16206);
and U16698 (N_16698,N_16467,N_16209);
nor U16699 (N_16699,N_16222,N_16204);
nand U16700 (N_16700,N_16223,N_16376);
and U16701 (N_16701,N_16290,N_16388);
and U16702 (N_16702,N_16353,N_16321);
nand U16703 (N_16703,N_16489,N_16454);
xor U16704 (N_16704,N_16346,N_16322);
and U16705 (N_16705,N_16325,N_16449);
and U16706 (N_16706,N_16392,N_16437);
or U16707 (N_16707,N_16386,N_16415);
or U16708 (N_16708,N_16415,N_16422);
xor U16709 (N_16709,N_16478,N_16496);
xor U16710 (N_16710,N_16411,N_16361);
nand U16711 (N_16711,N_16485,N_16476);
nor U16712 (N_16712,N_16361,N_16318);
or U16713 (N_16713,N_16357,N_16293);
and U16714 (N_16714,N_16223,N_16455);
and U16715 (N_16715,N_16266,N_16413);
and U16716 (N_16716,N_16388,N_16346);
or U16717 (N_16717,N_16345,N_16438);
nand U16718 (N_16718,N_16212,N_16461);
nand U16719 (N_16719,N_16432,N_16484);
nand U16720 (N_16720,N_16248,N_16339);
nand U16721 (N_16721,N_16395,N_16374);
xor U16722 (N_16722,N_16487,N_16218);
and U16723 (N_16723,N_16400,N_16379);
nor U16724 (N_16724,N_16460,N_16344);
and U16725 (N_16725,N_16364,N_16322);
nand U16726 (N_16726,N_16219,N_16426);
xnor U16727 (N_16727,N_16261,N_16420);
and U16728 (N_16728,N_16330,N_16264);
xor U16729 (N_16729,N_16272,N_16251);
and U16730 (N_16730,N_16364,N_16327);
and U16731 (N_16731,N_16357,N_16351);
xor U16732 (N_16732,N_16351,N_16288);
xnor U16733 (N_16733,N_16252,N_16251);
or U16734 (N_16734,N_16441,N_16351);
xnor U16735 (N_16735,N_16317,N_16247);
or U16736 (N_16736,N_16374,N_16409);
nand U16737 (N_16737,N_16284,N_16423);
nand U16738 (N_16738,N_16283,N_16296);
nor U16739 (N_16739,N_16422,N_16320);
xor U16740 (N_16740,N_16282,N_16467);
or U16741 (N_16741,N_16333,N_16407);
nand U16742 (N_16742,N_16348,N_16440);
nor U16743 (N_16743,N_16237,N_16468);
xnor U16744 (N_16744,N_16381,N_16443);
nand U16745 (N_16745,N_16440,N_16356);
or U16746 (N_16746,N_16248,N_16439);
or U16747 (N_16747,N_16439,N_16273);
nor U16748 (N_16748,N_16272,N_16458);
xor U16749 (N_16749,N_16438,N_16472);
nand U16750 (N_16750,N_16389,N_16405);
and U16751 (N_16751,N_16464,N_16298);
nand U16752 (N_16752,N_16354,N_16258);
nand U16753 (N_16753,N_16418,N_16324);
nor U16754 (N_16754,N_16464,N_16412);
nand U16755 (N_16755,N_16440,N_16457);
nand U16756 (N_16756,N_16291,N_16394);
xor U16757 (N_16757,N_16406,N_16436);
nor U16758 (N_16758,N_16383,N_16283);
xnor U16759 (N_16759,N_16469,N_16387);
and U16760 (N_16760,N_16278,N_16325);
and U16761 (N_16761,N_16257,N_16401);
nor U16762 (N_16762,N_16233,N_16215);
nand U16763 (N_16763,N_16251,N_16292);
xor U16764 (N_16764,N_16333,N_16270);
nor U16765 (N_16765,N_16240,N_16466);
xnor U16766 (N_16766,N_16414,N_16485);
nor U16767 (N_16767,N_16356,N_16237);
nand U16768 (N_16768,N_16436,N_16369);
xnor U16769 (N_16769,N_16386,N_16388);
or U16770 (N_16770,N_16348,N_16372);
nand U16771 (N_16771,N_16217,N_16337);
or U16772 (N_16772,N_16251,N_16382);
and U16773 (N_16773,N_16298,N_16315);
and U16774 (N_16774,N_16403,N_16423);
xor U16775 (N_16775,N_16213,N_16304);
xnor U16776 (N_16776,N_16226,N_16243);
or U16777 (N_16777,N_16351,N_16440);
or U16778 (N_16778,N_16471,N_16426);
nor U16779 (N_16779,N_16463,N_16262);
or U16780 (N_16780,N_16350,N_16304);
nor U16781 (N_16781,N_16420,N_16327);
or U16782 (N_16782,N_16247,N_16246);
or U16783 (N_16783,N_16338,N_16432);
nand U16784 (N_16784,N_16220,N_16382);
xor U16785 (N_16785,N_16363,N_16207);
and U16786 (N_16786,N_16399,N_16466);
xnor U16787 (N_16787,N_16236,N_16277);
and U16788 (N_16788,N_16469,N_16475);
or U16789 (N_16789,N_16484,N_16205);
or U16790 (N_16790,N_16273,N_16454);
nand U16791 (N_16791,N_16428,N_16233);
nand U16792 (N_16792,N_16200,N_16360);
xor U16793 (N_16793,N_16283,N_16248);
xnor U16794 (N_16794,N_16227,N_16288);
or U16795 (N_16795,N_16488,N_16437);
and U16796 (N_16796,N_16313,N_16375);
nor U16797 (N_16797,N_16249,N_16200);
xnor U16798 (N_16798,N_16412,N_16230);
or U16799 (N_16799,N_16425,N_16388);
or U16800 (N_16800,N_16691,N_16723);
and U16801 (N_16801,N_16600,N_16513);
nor U16802 (N_16802,N_16777,N_16563);
or U16803 (N_16803,N_16635,N_16579);
nand U16804 (N_16804,N_16732,N_16690);
or U16805 (N_16805,N_16675,N_16506);
and U16806 (N_16806,N_16741,N_16551);
or U16807 (N_16807,N_16788,N_16689);
and U16808 (N_16808,N_16783,N_16717);
nand U16809 (N_16809,N_16693,N_16668);
and U16810 (N_16810,N_16799,N_16770);
nand U16811 (N_16811,N_16743,N_16583);
and U16812 (N_16812,N_16501,N_16533);
nor U16813 (N_16813,N_16559,N_16613);
xnor U16814 (N_16814,N_16752,N_16699);
xnor U16815 (N_16815,N_16685,N_16784);
nand U16816 (N_16816,N_16779,N_16680);
nor U16817 (N_16817,N_16765,N_16644);
xor U16818 (N_16818,N_16584,N_16591);
nor U16819 (N_16819,N_16536,N_16586);
or U16820 (N_16820,N_16683,N_16603);
nor U16821 (N_16821,N_16522,N_16751);
or U16822 (N_16822,N_16658,N_16764);
and U16823 (N_16823,N_16767,N_16588);
or U16824 (N_16824,N_16669,N_16585);
and U16825 (N_16825,N_16570,N_16518);
or U16826 (N_16826,N_16527,N_16523);
or U16827 (N_16827,N_16581,N_16646);
and U16828 (N_16828,N_16507,N_16692);
and U16829 (N_16829,N_16514,N_16761);
nor U16830 (N_16830,N_16709,N_16617);
and U16831 (N_16831,N_16519,N_16557);
xor U16832 (N_16832,N_16554,N_16508);
nand U16833 (N_16833,N_16758,N_16776);
or U16834 (N_16834,N_16643,N_16636);
xor U16835 (N_16835,N_16597,N_16544);
and U16836 (N_16836,N_16778,N_16534);
and U16837 (N_16837,N_16667,N_16592);
or U16838 (N_16838,N_16549,N_16731);
nand U16839 (N_16839,N_16564,N_16730);
xor U16840 (N_16840,N_16612,N_16638);
or U16841 (N_16841,N_16673,N_16605);
nor U16842 (N_16842,N_16753,N_16678);
and U16843 (N_16843,N_16772,N_16754);
nor U16844 (N_16844,N_16755,N_16676);
nand U16845 (N_16845,N_16571,N_16704);
nand U16846 (N_16846,N_16567,N_16575);
xor U16847 (N_16847,N_16785,N_16653);
nor U16848 (N_16848,N_16759,N_16566);
nor U16849 (N_16849,N_16543,N_16782);
nand U16850 (N_16850,N_16684,N_16781);
xnor U16851 (N_16851,N_16516,N_16548);
or U16852 (N_16852,N_16745,N_16648);
nand U16853 (N_16853,N_16769,N_16798);
or U16854 (N_16854,N_16763,N_16766);
nand U16855 (N_16855,N_16572,N_16705);
xor U16856 (N_16856,N_16526,N_16629);
or U16857 (N_16857,N_16619,N_16512);
and U16858 (N_16858,N_16682,N_16604);
nand U16859 (N_16859,N_16627,N_16774);
and U16860 (N_16860,N_16511,N_16677);
xnor U16861 (N_16861,N_16748,N_16793);
or U16862 (N_16862,N_16504,N_16738);
or U16863 (N_16863,N_16651,N_16594);
nand U16864 (N_16864,N_16742,N_16671);
or U16865 (N_16865,N_16503,N_16568);
and U16866 (N_16866,N_16664,N_16618);
nor U16867 (N_16867,N_16590,N_16560);
and U16868 (N_16868,N_16562,N_16589);
nor U16869 (N_16869,N_16569,N_16724);
nand U16870 (N_16870,N_16598,N_16642);
nor U16871 (N_16871,N_16510,N_16734);
and U16872 (N_16872,N_16700,N_16532);
or U16873 (N_16873,N_16720,N_16707);
nand U16874 (N_16874,N_16609,N_16602);
or U16875 (N_16875,N_16744,N_16737);
and U16876 (N_16876,N_16553,N_16657);
nand U16877 (N_16877,N_16640,N_16735);
nand U16878 (N_16878,N_16726,N_16792);
xnor U16879 (N_16879,N_16686,N_16623);
nand U16880 (N_16880,N_16698,N_16630);
xor U16881 (N_16881,N_16681,N_16546);
and U16882 (N_16882,N_16728,N_16747);
and U16883 (N_16883,N_16580,N_16775);
nand U16884 (N_16884,N_16786,N_16702);
nand U16885 (N_16885,N_16652,N_16538);
or U16886 (N_16886,N_16666,N_16718);
nand U16887 (N_16887,N_16520,N_16521);
nor U16888 (N_16888,N_16573,N_16582);
and U16889 (N_16889,N_16736,N_16595);
xnor U16890 (N_16890,N_16556,N_16639);
or U16891 (N_16891,N_16650,N_16645);
nand U16892 (N_16892,N_16727,N_16708);
or U16893 (N_16893,N_16537,N_16525);
or U16894 (N_16894,N_16773,N_16637);
and U16895 (N_16895,N_16593,N_16626);
xnor U16896 (N_16896,N_16565,N_16714);
or U16897 (N_16897,N_16649,N_16539);
nand U16898 (N_16898,N_16659,N_16663);
nor U16899 (N_16899,N_16535,N_16550);
nor U16900 (N_16900,N_16596,N_16696);
or U16901 (N_16901,N_16515,N_16797);
and U16902 (N_16902,N_16631,N_16694);
or U16903 (N_16903,N_16509,N_16621);
xor U16904 (N_16904,N_16789,N_16502);
xor U16905 (N_16905,N_16787,N_16561);
nor U16906 (N_16906,N_16721,N_16628);
nor U16907 (N_16907,N_16711,N_16746);
and U16908 (N_16908,N_16749,N_16531);
xor U16909 (N_16909,N_16611,N_16796);
xnor U16910 (N_16910,N_16655,N_16713);
nor U16911 (N_16911,N_16587,N_16614);
or U16912 (N_16912,N_16719,N_16606);
nor U16913 (N_16913,N_16712,N_16601);
or U16914 (N_16914,N_16672,N_16624);
and U16915 (N_16915,N_16670,N_16687);
or U16916 (N_16916,N_16703,N_16701);
nand U16917 (N_16917,N_16555,N_16780);
nand U16918 (N_16918,N_16716,N_16654);
and U16919 (N_16919,N_16656,N_16661);
or U16920 (N_16920,N_16610,N_16760);
or U16921 (N_16921,N_16679,N_16608);
or U16922 (N_16922,N_16740,N_16674);
nor U16923 (N_16923,N_16771,N_16620);
xnor U16924 (N_16924,N_16517,N_16622);
nand U16925 (N_16925,N_16662,N_16794);
nor U16926 (N_16926,N_16541,N_16540);
nor U16927 (N_16927,N_16695,N_16733);
or U16928 (N_16928,N_16545,N_16524);
nand U16929 (N_16929,N_16697,N_16576);
nor U16930 (N_16930,N_16688,N_16665);
and U16931 (N_16931,N_16633,N_16725);
and U16932 (N_16932,N_16750,N_16578);
xor U16933 (N_16933,N_16634,N_16722);
nor U16934 (N_16934,N_16641,N_16558);
xnor U16935 (N_16935,N_16505,N_16768);
xor U16936 (N_16936,N_16756,N_16625);
or U16937 (N_16937,N_16616,N_16706);
nor U16938 (N_16938,N_16790,N_16552);
or U16939 (N_16939,N_16574,N_16795);
xnor U16940 (N_16940,N_16710,N_16715);
and U16941 (N_16941,N_16500,N_16577);
nor U16942 (N_16942,N_16757,N_16647);
and U16943 (N_16943,N_16528,N_16660);
nor U16944 (N_16944,N_16615,N_16530);
nor U16945 (N_16945,N_16599,N_16547);
nand U16946 (N_16946,N_16542,N_16739);
and U16947 (N_16947,N_16729,N_16791);
and U16948 (N_16948,N_16529,N_16762);
or U16949 (N_16949,N_16632,N_16607);
xor U16950 (N_16950,N_16631,N_16515);
and U16951 (N_16951,N_16666,N_16545);
and U16952 (N_16952,N_16788,N_16766);
xnor U16953 (N_16953,N_16759,N_16736);
nor U16954 (N_16954,N_16549,N_16612);
and U16955 (N_16955,N_16693,N_16611);
and U16956 (N_16956,N_16560,N_16552);
xnor U16957 (N_16957,N_16574,N_16546);
nand U16958 (N_16958,N_16697,N_16669);
nor U16959 (N_16959,N_16739,N_16683);
or U16960 (N_16960,N_16543,N_16645);
and U16961 (N_16961,N_16628,N_16518);
nand U16962 (N_16962,N_16792,N_16669);
and U16963 (N_16963,N_16550,N_16573);
or U16964 (N_16964,N_16620,N_16631);
nor U16965 (N_16965,N_16776,N_16705);
nand U16966 (N_16966,N_16513,N_16642);
and U16967 (N_16967,N_16618,N_16739);
xnor U16968 (N_16968,N_16514,N_16648);
xor U16969 (N_16969,N_16517,N_16590);
nor U16970 (N_16970,N_16773,N_16728);
xor U16971 (N_16971,N_16630,N_16624);
xor U16972 (N_16972,N_16777,N_16718);
nand U16973 (N_16973,N_16794,N_16536);
and U16974 (N_16974,N_16526,N_16634);
nand U16975 (N_16975,N_16737,N_16646);
xor U16976 (N_16976,N_16700,N_16788);
nand U16977 (N_16977,N_16712,N_16605);
nor U16978 (N_16978,N_16587,N_16736);
nand U16979 (N_16979,N_16549,N_16515);
xor U16980 (N_16980,N_16691,N_16731);
nor U16981 (N_16981,N_16674,N_16666);
xor U16982 (N_16982,N_16656,N_16561);
nor U16983 (N_16983,N_16749,N_16729);
and U16984 (N_16984,N_16622,N_16776);
or U16985 (N_16985,N_16530,N_16650);
nor U16986 (N_16986,N_16743,N_16690);
or U16987 (N_16987,N_16653,N_16515);
xor U16988 (N_16988,N_16539,N_16504);
nand U16989 (N_16989,N_16729,N_16519);
nor U16990 (N_16990,N_16544,N_16615);
or U16991 (N_16991,N_16680,N_16708);
and U16992 (N_16992,N_16576,N_16561);
or U16993 (N_16993,N_16673,N_16600);
and U16994 (N_16994,N_16509,N_16637);
nor U16995 (N_16995,N_16700,N_16724);
xor U16996 (N_16996,N_16591,N_16667);
nor U16997 (N_16997,N_16651,N_16645);
or U16998 (N_16998,N_16508,N_16719);
nand U16999 (N_16999,N_16782,N_16695);
xnor U17000 (N_17000,N_16766,N_16582);
nand U17001 (N_17001,N_16774,N_16540);
nor U17002 (N_17002,N_16738,N_16744);
and U17003 (N_17003,N_16700,N_16530);
nor U17004 (N_17004,N_16681,N_16593);
or U17005 (N_17005,N_16645,N_16517);
nand U17006 (N_17006,N_16744,N_16732);
or U17007 (N_17007,N_16544,N_16683);
or U17008 (N_17008,N_16566,N_16501);
nor U17009 (N_17009,N_16725,N_16745);
nor U17010 (N_17010,N_16697,N_16550);
nor U17011 (N_17011,N_16682,N_16657);
nand U17012 (N_17012,N_16773,N_16557);
and U17013 (N_17013,N_16626,N_16658);
nand U17014 (N_17014,N_16565,N_16547);
xor U17015 (N_17015,N_16769,N_16708);
xnor U17016 (N_17016,N_16558,N_16712);
xor U17017 (N_17017,N_16770,N_16530);
and U17018 (N_17018,N_16789,N_16726);
or U17019 (N_17019,N_16679,N_16535);
and U17020 (N_17020,N_16754,N_16528);
nand U17021 (N_17021,N_16637,N_16724);
nand U17022 (N_17022,N_16660,N_16519);
and U17023 (N_17023,N_16580,N_16689);
nor U17024 (N_17024,N_16642,N_16608);
nor U17025 (N_17025,N_16760,N_16523);
nor U17026 (N_17026,N_16560,N_16672);
nand U17027 (N_17027,N_16581,N_16677);
nor U17028 (N_17028,N_16787,N_16679);
and U17029 (N_17029,N_16636,N_16758);
and U17030 (N_17030,N_16672,N_16756);
xnor U17031 (N_17031,N_16795,N_16750);
nor U17032 (N_17032,N_16503,N_16622);
nor U17033 (N_17033,N_16742,N_16592);
and U17034 (N_17034,N_16635,N_16610);
xor U17035 (N_17035,N_16687,N_16708);
and U17036 (N_17036,N_16784,N_16760);
xnor U17037 (N_17037,N_16634,N_16660);
and U17038 (N_17038,N_16635,N_16771);
nor U17039 (N_17039,N_16710,N_16517);
nor U17040 (N_17040,N_16536,N_16683);
and U17041 (N_17041,N_16609,N_16637);
nand U17042 (N_17042,N_16655,N_16744);
or U17043 (N_17043,N_16717,N_16671);
or U17044 (N_17044,N_16613,N_16561);
and U17045 (N_17045,N_16779,N_16739);
and U17046 (N_17046,N_16761,N_16690);
nor U17047 (N_17047,N_16714,N_16573);
or U17048 (N_17048,N_16691,N_16689);
nor U17049 (N_17049,N_16654,N_16785);
or U17050 (N_17050,N_16761,N_16660);
nand U17051 (N_17051,N_16592,N_16633);
nand U17052 (N_17052,N_16709,N_16649);
xor U17053 (N_17053,N_16560,N_16574);
xor U17054 (N_17054,N_16740,N_16534);
xor U17055 (N_17055,N_16520,N_16618);
and U17056 (N_17056,N_16613,N_16792);
nand U17057 (N_17057,N_16515,N_16548);
and U17058 (N_17058,N_16601,N_16625);
or U17059 (N_17059,N_16726,N_16700);
nor U17060 (N_17060,N_16692,N_16770);
or U17061 (N_17061,N_16673,N_16765);
nor U17062 (N_17062,N_16604,N_16799);
nor U17063 (N_17063,N_16503,N_16590);
nor U17064 (N_17064,N_16628,N_16751);
nor U17065 (N_17065,N_16658,N_16785);
nor U17066 (N_17066,N_16570,N_16668);
nand U17067 (N_17067,N_16579,N_16775);
xnor U17068 (N_17068,N_16634,N_16706);
and U17069 (N_17069,N_16536,N_16753);
nand U17070 (N_17070,N_16523,N_16720);
nand U17071 (N_17071,N_16593,N_16765);
or U17072 (N_17072,N_16713,N_16720);
nand U17073 (N_17073,N_16524,N_16536);
and U17074 (N_17074,N_16547,N_16659);
nand U17075 (N_17075,N_16526,N_16752);
nand U17076 (N_17076,N_16629,N_16788);
xor U17077 (N_17077,N_16553,N_16540);
nor U17078 (N_17078,N_16661,N_16703);
and U17079 (N_17079,N_16556,N_16739);
nor U17080 (N_17080,N_16558,N_16524);
xnor U17081 (N_17081,N_16692,N_16601);
nor U17082 (N_17082,N_16646,N_16666);
xnor U17083 (N_17083,N_16518,N_16749);
nor U17084 (N_17084,N_16602,N_16780);
nor U17085 (N_17085,N_16719,N_16707);
nor U17086 (N_17086,N_16675,N_16623);
or U17087 (N_17087,N_16687,N_16598);
or U17088 (N_17088,N_16787,N_16572);
nand U17089 (N_17089,N_16694,N_16554);
or U17090 (N_17090,N_16594,N_16641);
nor U17091 (N_17091,N_16710,N_16696);
xnor U17092 (N_17092,N_16505,N_16506);
and U17093 (N_17093,N_16523,N_16678);
or U17094 (N_17094,N_16578,N_16743);
nor U17095 (N_17095,N_16638,N_16748);
or U17096 (N_17096,N_16620,N_16637);
and U17097 (N_17097,N_16736,N_16750);
xor U17098 (N_17098,N_16728,N_16626);
and U17099 (N_17099,N_16575,N_16628);
or U17100 (N_17100,N_16960,N_17036);
nand U17101 (N_17101,N_16982,N_16861);
xor U17102 (N_17102,N_16824,N_16964);
or U17103 (N_17103,N_16991,N_16939);
or U17104 (N_17104,N_16979,N_16980);
nand U17105 (N_17105,N_16938,N_16888);
or U17106 (N_17106,N_17029,N_16972);
or U17107 (N_17107,N_16836,N_16987);
nand U17108 (N_17108,N_16838,N_17024);
xor U17109 (N_17109,N_16802,N_17003);
nand U17110 (N_17110,N_16916,N_16818);
or U17111 (N_17111,N_16927,N_17043);
xnor U17112 (N_17112,N_17011,N_17052);
or U17113 (N_17113,N_17055,N_16808);
and U17114 (N_17114,N_17050,N_16833);
or U17115 (N_17115,N_16975,N_17012);
or U17116 (N_17116,N_17006,N_16864);
xnor U17117 (N_17117,N_16950,N_16875);
nand U17118 (N_17118,N_17001,N_17005);
or U17119 (N_17119,N_17078,N_16989);
and U17120 (N_17120,N_17059,N_16966);
nor U17121 (N_17121,N_16856,N_16919);
nor U17122 (N_17122,N_17034,N_16829);
xnor U17123 (N_17123,N_16957,N_16832);
xnor U17124 (N_17124,N_16901,N_17093);
nand U17125 (N_17125,N_17079,N_16896);
xnor U17126 (N_17126,N_16895,N_17083);
and U17127 (N_17127,N_16819,N_16977);
and U17128 (N_17128,N_17032,N_16913);
nor U17129 (N_17129,N_16827,N_16998);
xnor U17130 (N_17130,N_17053,N_16868);
nor U17131 (N_17131,N_17014,N_16915);
nor U17132 (N_17132,N_16910,N_16929);
nor U17133 (N_17133,N_16889,N_16800);
and U17134 (N_17134,N_17021,N_17041);
and U17135 (N_17135,N_17016,N_16962);
and U17136 (N_17136,N_17091,N_16988);
nand U17137 (N_17137,N_16933,N_16995);
xor U17138 (N_17138,N_17070,N_17088);
or U17139 (N_17139,N_16843,N_16924);
and U17140 (N_17140,N_16810,N_16981);
nand U17141 (N_17141,N_17084,N_16955);
and U17142 (N_17142,N_17023,N_16863);
xor U17143 (N_17143,N_17064,N_17010);
nand U17144 (N_17144,N_16958,N_17062);
nor U17145 (N_17145,N_16935,N_16805);
nand U17146 (N_17146,N_16920,N_17013);
nor U17147 (N_17147,N_16934,N_16999);
or U17148 (N_17148,N_17068,N_16961);
nand U17149 (N_17149,N_16816,N_16912);
nand U17150 (N_17150,N_16867,N_16951);
and U17151 (N_17151,N_16897,N_16905);
or U17152 (N_17152,N_16853,N_16874);
or U17153 (N_17153,N_17020,N_17097);
or U17154 (N_17154,N_16954,N_17092);
nor U17155 (N_17155,N_16876,N_17007);
xor U17156 (N_17156,N_17073,N_16963);
and U17157 (N_17157,N_16880,N_17004);
nor U17158 (N_17158,N_16994,N_16893);
nand U17159 (N_17159,N_17042,N_16922);
nor U17160 (N_17160,N_16812,N_16967);
or U17161 (N_17161,N_17089,N_17035);
and U17162 (N_17162,N_17033,N_16907);
or U17163 (N_17163,N_17060,N_17085);
xnor U17164 (N_17164,N_16945,N_16984);
nor U17165 (N_17165,N_16826,N_16930);
or U17166 (N_17166,N_16848,N_17074);
xnor U17167 (N_17167,N_16837,N_16886);
xor U17168 (N_17168,N_16872,N_17075);
or U17169 (N_17169,N_16976,N_16814);
nand U17170 (N_17170,N_16834,N_16918);
nor U17171 (N_17171,N_16801,N_16894);
xnor U17172 (N_17172,N_16909,N_16877);
nand U17173 (N_17173,N_17082,N_16831);
or U17174 (N_17174,N_16925,N_16865);
or U17175 (N_17175,N_17065,N_17000);
nand U17176 (N_17176,N_16936,N_16850);
nor U17177 (N_17177,N_16956,N_16821);
and U17178 (N_17178,N_16996,N_16965);
nand U17179 (N_17179,N_16844,N_16928);
nor U17180 (N_17180,N_16904,N_16873);
xnor U17181 (N_17181,N_16891,N_16835);
xor U17182 (N_17182,N_16804,N_16943);
and U17183 (N_17183,N_16911,N_17038);
xor U17184 (N_17184,N_17009,N_16858);
nand U17185 (N_17185,N_16917,N_16947);
nand U17186 (N_17186,N_16840,N_17094);
xor U17187 (N_17187,N_16898,N_16871);
xor U17188 (N_17188,N_16830,N_16900);
and U17189 (N_17189,N_16878,N_17076);
nand U17190 (N_17190,N_17037,N_16879);
nand U17191 (N_17191,N_16937,N_16903);
and U17192 (N_17192,N_16846,N_17026);
and U17193 (N_17193,N_17044,N_16887);
nor U17194 (N_17194,N_16908,N_17066);
and U17195 (N_17195,N_17045,N_16841);
or U17196 (N_17196,N_17054,N_16986);
or U17197 (N_17197,N_16932,N_16906);
and U17198 (N_17198,N_16931,N_16842);
or U17199 (N_17199,N_16882,N_17049);
or U17200 (N_17200,N_17015,N_16953);
and U17201 (N_17201,N_17051,N_17099);
or U17202 (N_17202,N_16983,N_17039);
or U17203 (N_17203,N_17025,N_16993);
and U17204 (N_17204,N_16883,N_17002);
xnor U17205 (N_17205,N_17030,N_16959);
xor U17206 (N_17206,N_16828,N_16885);
nand U17207 (N_17207,N_16817,N_17080);
and U17208 (N_17208,N_16869,N_16855);
xor U17209 (N_17209,N_16940,N_17067);
xor U17210 (N_17210,N_16854,N_17008);
nand U17211 (N_17211,N_16899,N_16839);
or U17212 (N_17212,N_16921,N_17056);
and U17213 (N_17213,N_17096,N_16825);
and U17214 (N_17214,N_16857,N_16823);
nor U17215 (N_17215,N_16815,N_17028);
and U17216 (N_17216,N_16969,N_16968);
and U17217 (N_17217,N_17040,N_17072);
xor U17218 (N_17218,N_17095,N_16902);
nor U17219 (N_17219,N_16881,N_16926);
nand U17220 (N_17220,N_16870,N_17057);
xnor U17221 (N_17221,N_16884,N_17090);
and U17222 (N_17222,N_16859,N_17031);
nand U17223 (N_17223,N_16892,N_17071);
and U17224 (N_17224,N_16974,N_16862);
and U17225 (N_17225,N_16851,N_16942);
nor U17226 (N_17226,N_16946,N_17081);
or U17227 (N_17227,N_16807,N_16978);
and U17228 (N_17228,N_16860,N_17048);
xor U17229 (N_17229,N_17046,N_16866);
xnor U17230 (N_17230,N_16952,N_17086);
or U17231 (N_17231,N_17087,N_16949);
and U17232 (N_17232,N_17058,N_17047);
and U17233 (N_17233,N_16847,N_16914);
nand U17234 (N_17234,N_16820,N_17061);
or U17235 (N_17235,N_17017,N_17063);
and U17236 (N_17236,N_16822,N_16845);
xor U17237 (N_17237,N_16990,N_16803);
and U17238 (N_17238,N_16970,N_16985);
nand U17239 (N_17239,N_16852,N_17077);
nor U17240 (N_17240,N_16806,N_16813);
nor U17241 (N_17241,N_16973,N_17022);
or U17242 (N_17242,N_16971,N_17018);
or U17243 (N_17243,N_16992,N_16923);
or U17244 (N_17244,N_16849,N_16944);
nor U17245 (N_17245,N_17069,N_16811);
and U17246 (N_17246,N_17019,N_17098);
nand U17247 (N_17247,N_16941,N_16809);
nor U17248 (N_17248,N_16890,N_16948);
nand U17249 (N_17249,N_16997,N_17027);
nand U17250 (N_17250,N_17062,N_16845);
nand U17251 (N_17251,N_16859,N_16840);
nand U17252 (N_17252,N_17095,N_16943);
nor U17253 (N_17253,N_17078,N_16937);
nor U17254 (N_17254,N_17083,N_17021);
nor U17255 (N_17255,N_17070,N_17031);
and U17256 (N_17256,N_16868,N_16898);
nand U17257 (N_17257,N_16861,N_17092);
nand U17258 (N_17258,N_17080,N_17027);
nand U17259 (N_17259,N_16990,N_17082);
nor U17260 (N_17260,N_16821,N_16928);
xnor U17261 (N_17261,N_17016,N_16938);
xor U17262 (N_17262,N_16913,N_16955);
and U17263 (N_17263,N_16976,N_16833);
and U17264 (N_17264,N_16932,N_17042);
or U17265 (N_17265,N_16810,N_17084);
nor U17266 (N_17266,N_16847,N_17066);
nand U17267 (N_17267,N_16878,N_16931);
xnor U17268 (N_17268,N_16910,N_16843);
and U17269 (N_17269,N_17046,N_17088);
or U17270 (N_17270,N_16874,N_16998);
or U17271 (N_17271,N_17015,N_16805);
nor U17272 (N_17272,N_17002,N_17047);
and U17273 (N_17273,N_17047,N_17087);
nand U17274 (N_17274,N_17016,N_16805);
or U17275 (N_17275,N_16813,N_16895);
and U17276 (N_17276,N_16859,N_16997);
xor U17277 (N_17277,N_16885,N_17083);
or U17278 (N_17278,N_16960,N_16983);
and U17279 (N_17279,N_17083,N_16970);
or U17280 (N_17280,N_17047,N_17008);
or U17281 (N_17281,N_16977,N_16831);
or U17282 (N_17282,N_16881,N_16987);
xor U17283 (N_17283,N_16960,N_16873);
nand U17284 (N_17284,N_16814,N_16845);
or U17285 (N_17285,N_16836,N_16936);
nor U17286 (N_17286,N_16920,N_16921);
nand U17287 (N_17287,N_16826,N_16949);
nor U17288 (N_17288,N_17017,N_17052);
xnor U17289 (N_17289,N_16846,N_16826);
and U17290 (N_17290,N_17041,N_16971);
nand U17291 (N_17291,N_16984,N_16940);
nand U17292 (N_17292,N_16851,N_17096);
xnor U17293 (N_17293,N_17005,N_16976);
or U17294 (N_17294,N_17081,N_17014);
or U17295 (N_17295,N_16920,N_16800);
xnor U17296 (N_17296,N_17080,N_16897);
and U17297 (N_17297,N_16856,N_17030);
and U17298 (N_17298,N_17055,N_16834);
or U17299 (N_17299,N_17057,N_16820);
nand U17300 (N_17300,N_16882,N_16817);
and U17301 (N_17301,N_16845,N_17007);
or U17302 (N_17302,N_16942,N_16856);
or U17303 (N_17303,N_16905,N_16914);
xor U17304 (N_17304,N_16820,N_16914);
xor U17305 (N_17305,N_16863,N_16838);
and U17306 (N_17306,N_16843,N_16865);
nor U17307 (N_17307,N_16944,N_16868);
or U17308 (N_17308,N_16884,N_16881);
xnor U17309 (N_17309,N_16979,N_16821);
or U17310 (N_17310,N_16877,N_17024);
and U17311 (N_17311,N_16808,N_17062);
nor U17312 (N_17312,N_17063,N_16922);
xnor U17313 (N_17313,N_17012,N_16820);
or U17314 (N_17314,N_16962,N_16912);
or U17315 (N_17315,N_16941,N_16900);
nor U17316 (N_17316,N_16934,N_16940);
and U17317 (N_17317,N_16910,N_16899);
nand U17318 (N_17318,N_16928,N_16805);
nor U17319 (N_17319,N_16829,N_16871);
xor U17320 (N_17320,N_16924,N_17080);
xnor U17321 (N_17321,N_16848,N_16807);
and U17322 (N_17322,N_17042,N_16908);
and U17323 (N_17323,N_17018,N_17097);
or U17324 (N_17324,N_16995,N_16919);
or U17325 (N_17325,N_16818,N_16815);
and U17326 (N_17326,N_16977,N_17084);
xnor U17327 (N_17327,N_16926,N_16863);
xnor U17328 (N_17328,N_17003,N_16888);
and U17329 (N_17329,N_16855,N_16956);
nor U17330 (N_17330,N_17085,N_16863);
or U17331 (N_17331,N_16859,N_16940);
xnor U17332 (N_17332,N_16974,N_16942);
xor U17333 (N_17333,N_17049,N_16959);
nand U17334 (N_17334,N_16924,N_16867);
or U17335 (N_17335,N_16831,N_16841);
nor U17336 (N_17336,N_16973,N_16888);
nor U17337 (N_17337,N_16945,N_16858);
or U17338 (N_17338,N_16856,N_17027);
xnor U17339 (N_17339,N_16839,N_16987);
nand U17340 (N_17340,N_17086,N_16896);
nor U17341 (N_17341,N_16952,N_17039);
nor U17342 (N_17342,N_17076,N_17073);
xor U17343 (N_17343,N_16999,N_17049);
or U17344 (N_17344,N_16817,N_16908);
nand U17345 (N_17345,N_16905,N_16870);
and U17346 (N_17346,N_17062,N_17098);
nand U17347 (N_17347,N_16978,N_16831);
or U17348 (N_17348,N_16998,N_16939);
or U17349 (N_17349,N_17061,N_16963);
nor U17350 (N_17350,N_16806,N_17096);
nor U17351 (N_17351,N_17047,N_17092);
nand U17352 (N_17352,N_16938,N_16825);
or U17353 (N_17353,N_16930,N_16929);
or U17354 (N_17354,N_16863,N_17067);
or U17355 (N_17355,N_17038,N_16956);
and U17356 (N_17356,N_16945,N_16959);
nor U17357 (N_17357,N_16811,N_17063);
xnor U17358 (N_17358,N_16996,N_16872);
and U17359 (N_17359,N_16930,N_16979);
nor U17360 (N_17360,N_16945,N_17072);
and U17361 (N_17361,N_16936,N_17010);
or U17362 (N_17362,N_17016,N_16896);
and U17363 (N_17363,N_17090,N_16969);
nand U17364 (N_17364,N_16992,N_16835);
or U17365 (N_17365,N_17004,N_17041);
nor U17366 (N_17366,N_17056,N_17043);
and U17367 (N_17367,N_16814,N_16944);
or U17368 (N_17368,N_16918,N_17051);
xnor U17369 (N_17369,N_16928,N_16893);
and U17370 (N_17370,N_16872,N_17057);
or U17371 (N_17371,N_16922,N_17027);
nand U17372 (N_17372,N_17006,N_16878);
and U17373 (N_17373,N_17007,N_16868);
nor U17374 (N_17374,N_16961,N_16801);
nand U17375 (N_17375,N_17026,N_16918);
nand U17376 (N_17376,N_16968,N_16895);
xnor U17377 (N_17377,N_17041,N_16853);
nor U17378 (N_17378,N_16998,N_17016);
nor U17379 (N_17379,N_16810,N_17088);
nand U17380 (N_17380,N_16992,N_16803);
xor U17381 (N_17381,N_16936,N_17085);
nor U17382 (N_17382,N_16996,N_17077);
nand U17383 (N_17383,N_16990,N_16937);
and U17384 (N_17384,N_17046,N_17038);
and U17385 (N_17385,N_17042,N_16947);
nor U17386 (N_17386,N_17038,N_16866);
xnor U17387 (N_17387,N_16907,N_16965);
xnor U17388 (N_17388,N_17076,N_17019);
nor U17389 (N_17389,N_17073,N_16912);
xnor U17390 (N_17390,N_17046,N_16850);
nor U17391 (N_17391,N_16874,N_16820);
nand U17392 (N_17392,N_16960,N_17021);
nor U17393 (N_17393,N_16869,N_16891);
or U17394 (N_17394,N_16898,N_17012);
nand U17395 (N_17395,N_17085,N_17070);
nor U17396 (N_17396,N_16895,N_17003);
or U17397 (N_17397,N_16915,N_16844);
and U17398 (N_17398,N_16958,N_16915);
or U17399 (N_17399,N_16861,N_16954);
xor U17400 (N_17400,N_17308,N_17240);
or U17401 (N_17401,N_17117,N_17154);
xor U17402 (N_17402,N_17113,N_17132);
nor U17403 (N_17403,N_17316,N_17325);
nor U17404 (N_17404,N_17378,N_17287);
xnor U17405 (N_17405,N_17131,N_17291);
and U17406 (N_17406,N_17344,N_17149);
xor U17407 (N_17407,N_17277,N_17341);
xor U17408 (N_17408,N_17207,N_17186);
or U17409 (N_17409,N_17280,N_17255);
or U17410 (N_17410,N_17193,N_17133);
nand U17411 (N_17411,N_17103,N_17336);
xor U17412 (N_17412,N_17122,N_17129);
nand U17413 (N_17413,N_17359,N_17266);
and U17414 (N_17414,N_17357,N_17127);
and U17415 (N_17415,N_17331,N_17296);
nand U17416 (N_17416,N_17295,N_17318);
nand U17417 (N_17417,N_17145,N_17142);
xnor U17418 (N_17418,N_17352,N_17206);
nor U17419 (N_17419,N_17355,N_17302);
nor U17420 (N_17420,N_17115,N_17320);
or U17421 (N_17421,N_17157,N_17164);
and U17422 (N_17422,N_17262,N_17343);
nand U17423 (N_17423,N_17261,N_17274);
nand U17424 (N_17424,N_17246,N_17367);
or U17425 (N_17425,N_17241,N_17156);
or U17426 (N_17426,N_17168,N_17310);
nor U17427 (N_17427,N_17324,N_17214);
and U17428 (N_17428,N_17201,N_17155);
nor U17429 (N_17429,N_17259,N_17312);
nor U17430 (N_17430,N_17353,N_17144);
or U17431 (N_17431,N_17181,N_17249);
nand U17432 (N_17432,N_17363,N_17342);
xor U17433 (N_17433,N_17323,N_17375);
or U17434 (N_17434,N_17313,N_17196);
or U17435 (N_17435,N_17300,N_17118);
or U17436 (N_17436,N_17285,N_17205);
or U17437 (N_17437,N_17260,N_17163);
and U17438 (N_17438,N_17381,N_17385);
nand U17439 (N_17439,N_17368,N_17227);
nor U17440 (N_17440,N_17383,N_17338);
nand U17441 (N_17441,N_17224,N_17101);
and U17442 (N_17442,N_17251,N_17237);
nor U17443 (N_17443,N_17123,N_17172);
nand U17444 (N_17444,N_17140,N_17372);
nand U17445 (N_17445,N_17257,N_17350);
and U17446 (N_17446,N_17263,N_17134);
or U17447 (N_17447,N_17146,N_17126);
nor U17448 (N_17448,N_17100,N_17178);
or U17449 (N_17449,N_17170,N_17198);
and U17450 (N_17450,N_17314,N_17190);
and U17451 (N_17451,N_17119,N_17221);
nand U17452 (N_17452,N_17387,N_17319);
nor U17453 (N_17453,N_17254,N_17309);
and U17454 (N_17454,N_17138,N_17121);
or U17455 (N_17455,N_17223,N_17272);
xnor U17456 (N_17456,N_17374,N_17346);
nand U17457 (N_17457,N_17289,N_17269);
xor U17458 (N_17458,N_17150,N_17361);
nand U17459 (N_17459,N_17199,N_17216);
nor U17460 (N_17460,N_17347,N_17328);
xor U17461 (N_17461,N_17128,N_17107);
nor U17462 (N_17462,N_17398,N_17171);
xor U17463 (N_17463,N_17185,N_17162);
nor U17464 (N_17464,N_17377,N_17130);
nand U17465 (N_17465,N_17340,N_17362);
nor U17466 (N_17466,N_17229,N_17376);
xor U17467 (N_17467,N_17180,N_17332);
and U17468 (N_17468,N_17158,N_17268);
and U17469 (N_17469,N_17384,N_17183);
nor U17470 (N_17470,N_17187,N_17116);
nand U17471 (N_17471,N_17226,N_17258);
nand U17472 (N_17472,N_17165,N_17232);
nor U17473 (N_17473,N_17195,N_17160);
or U17474 (N_17474,N_17151,N_17174);
or U17475 (N_17475,N_17211,N_17311);
nor U17476 (N_17476,N_17239,N_17242);
or U17477 (N_17477,N_17395,N_17124);
nand U17478 (N_17478,N_17369,N_17380);
nand U17479 (N_17479,N_17202,N_17371);
xnor U17480 (N_17480,N_17213,N_17326);
and U17481 (N_17481,N_17109,N_17147);
or U17482 (N_17482,N_17191,N_17348);
nand U17483 (N_17483,N_17243,N_17264);
nor U17484 (N_17484,N_17321,N_17373);
xor U17485 (N_17485,N_17281,N_17386);
or U17486 (N_17486,N_17200,N_17245);
nand U17487 (N_17487,N_17382,N_17188);
nor U17488 (N_17488,N_17365,N_17278);
xor U17489 (N_17489,N_17161,N_17292);
or U17490 (N_17490,N_17339,N_17110);
nand U17491 (N_17491,N_17379,N_17212);
xnor U17492 (N_17492,N_17112,N_17228);
nor U17493 (N_17493,N_17293,N_17286);
and U17494 (N_17494,N_17301,N_17218);
and U17495 (N_17495,N_17279,N_17233);
nand U17496 (N_17496,N_17111,N_17337);
nand U17497 (N_17497,N_17322,N_17217);
xor U17498 (N_17498,N_17210,N_17105);
or U17499 (N_17499,N_17358,N_17219);
xor U17500 (N_17500,N_17139,N_17238);
and U17501 (N_17501,N_17390,N_17177);
nor U17502 (N_17502,N_17152,N_17276);
xor U17503 (N_17503,N_17391,N_17335);
or U17504 (N_17504,N_17333,N_17273);
and U17505 (N_17505,N_17143,N_17225);
or U17506 (N_17506,N_17329,N_17153);
xor U17507 (N_17507,N_17290,N_17370);
and U17508 (N_17508,N_17204,N_17208);
xor U17509 (N_17509,N_17299,N_17288);
or U17510 (N_17510,N_17234,N_17394);
or U17511 (N_17511,N_17197,N_17388);
nand U17512 (N_17512,N_17250,N_17297);
nand U17513 (N_17513,N_17235,N_17192);
or U17514 (N_17514,N_17215,N_17231);
nor U17515 (N_17515,N_17102,N_17351);
and U17516 (N_17516,N_17393,N_17148);
and U17517 (N_17517,N_17270,N_17303);
and U17518 (N_17518,N_17159,N_17298);
nor U17519 (N_17519,N_17167,N_17360);
nand U17520 (N_17520,N_17108,N_17244);
nor U17521 (N_17521,N_17230,N_17248);
xor U17522 (N_17522,N_17236,N_17173);
xnor U17523 (N_17523,N_17120,N_17169);
nor U17524 (N_17524,N_17141,N_17267);
or U17525 (N_17525,N_17399,N_17283);
nor U17526 (N_17526,N_17306,N_17364);
and U17527 (N_17527,N_17317,N_17182);
or U17528 (N_17528,N_17305,N_17203);
nand U17529 (N_17529,N_17354,N_17275);
xnor U17530 (N_17530,N_17252,N_17327);
and U17531 (N_17531,N_17220,N_17282);
nand U17532 (N_17532,N_17209,N_17104);
nand U17533 (N_17533,N_17349,N_17106);
nor U17534 (N_17534,N_17397,N_17271);
nand U17535 (N_17535,N_17176,N_17179);
and U17536 (N_17536,N_17366,N_17284);
and U17537 (N_17537,N_17307,N_17166);
nand U17538 (N_17538,N_17356,N_17253);
nor U17539 (N_17539,N_17189,N_17184);
nor U17540 (N_17540,N_17392,N_17222);
and U17541 (N_17541,N_17137,N_17330);
and U17542 (N_17542,N_17396,N_17345);
nand U17543 (N_17543,N_17334,N_17136);
nand U17544 (N_17544,N_17125,N_17247);
xor U17545 (N_17545,N_17389,N_17135);
nand U17546 (N_17546,N_17315,N_17114);
xnor U17547 (N_17547,N_17304,N_17256);
nor U17548 (N_17548,N_17294,N_17265);
nand U17549 (N_17549,N_17175,N_17194);
nand U17550 (N_17550,N_17146,N_17305);
nand U17551 (N_17551,N_17350,N_17278);
xor U17552 (N_17552,N_17313,N_17280);
nor U17553 (N_17553,N_17143,N_17123);
or U17554 (N_17554,N_17144,N_17106);
nand U17555 (N_17555,N_17318,N_17274);
nand U17556 (N_17556,N_17102,N_17130);
or U17557 (N_17557,N_17275,N_17217);
xor U17558 (N_17558,N_17293,N_17337);
xnor U17559 (N_17559,N_17146,N_17102);
nand U17560 (N_17560,N_17141,N_17328);
and U17561 (N_17561,N_17372,N_17181);
nand U17562 (N_17562,N_17316,N_17237);
nand U17563 (N_17563,N_17340,N_17224);
xnor U17564 (N_17564,N_17258,N_17286);
nand U17565 (N_17565,N_17175,N_17128);
nand U17566 (N_17566,N_17332,N_17266);
nor U17567 (N_17567,N_17136,N_17219);
nor U17568 (N_17568,N_17203,N_17261);
or U17569 (N_17569,N_17240,N_17283);
or U17570 (N_17570,N_17164,N_17347);
and U17571 (N_17571,N_17172,N_17185);
or U17572 (N_17572,N_17369,N_17343);
or U17573 (N_17573,N_17367,N_17286);
nor U17574 (N_17574,N_17252,N_17182);
and U17575 (N_17575,N_17342,N_17112);
xnor U17576 (N_17576,N_17202,N_17348);
and U17577 (N_17577,N_17194,N_17326);
or U17578 (N_17578,N_17257,N_17243);
or U17579 (N_17579,N_17120,N_17326);
and U17580 (N_17580,N_17153,N_17313);
xnor U17581 (N_17581,N_17274,N_17368);
and U17582 (N_17582,N_17164,N_17346);
nor U17583 (N_17583,N_17324,N_17196);
nand U17584 (N_17584,N_17206,N_17340);
nor U17585 (N_17585,N_17331,N_17349);
or U17586 (N_17586,N_17194,N_17196);
xor U17587 (N_17587,N_17147,N_17278);
or U17588 (N_17588,N_17276,N_17349);
nand U17589 (N_17589,N_17158,N_17272);
nand U17590 (N_17590,N_17232,N_17371);
nand U17591 (N_17591,N_17111,N_17154);
or U17592 (N_17592,N_17225,N_17375);
or U17593 (N_17593,N_17360,N_17172);
xor U17594 (N_17594,N_17255,N_17311);
nor U17595 (N_17595,N_17364,N_17203);
nor U17596 (N_17596,N_17117,N_17333);
nand U17597 (N_17597,N_17362,N_17399);
nand U17598 (N_17598,N_17344,N_17168);
xnor U17599 (N_17599,N_17232,N_17267);
nand U17600 (N_17600,N_17293,N_17353);
or U17601 (N_17601,N_17354,N_17140);
nor U17602 (N_17602,N_17159,N_17239);
nand U17603 (N_17603,N_17182,N_17279);
or U17604 (N_17604,N_17172,N_17234);
or U17605 (N_17605,N_17132,N_17395);
nand U17606 (N_17606,N_17146,N_17241);
nand U17607 (N_17607,N_17304,N_17334);
xor U17608 (N_17608,N_17246,N_17281);
and U17609 (N_17609,N_17290,N_17245);
xor U17610 (N_17610,N_17364,N_17288);
nor U17611 (N_17611,N_17141,N_17174);
nand U17612 (N_17612,N_17111,N_17285);
nor U17613 (N_17613,N_17286,N_17294);
xnor U17614 (N_17614,N_17218,N_17384);
xor U17615 (N_17615,N_17257,N_17316);
nand U17616 (N_17616,N_17309,N_17352);
nand U17617 (N_17617,N_17264,N_17149);
or U17618 (N_17618,N_17236,N_17179);
and U17619 (N_17619,N_17321,N_17257);
and U17620 (N_17620,N_17345,N_17192);
nor U17621 (N_17621,N_17344,N_17369);
xor U17622 (N_17622,N_17228,N_17167);
nand U17623 (N_17623,N_17229,N_17380);
nor U17624 (N_17624,N_17311,N_17334);
and U17625 (N_17625,N_17147,N_17315);
nor U17626 (N_17626,N_17246,N_17197);
xor U17627 (N_17627,N_17248,N_17176);
and U17628 (N_17628,N_17152,N_17329);
or U17629 (N_17629,N_17259,N_17106);
xor U17630 (N_17630,N_17165,N_17242);
and U17631 (N_17631,N_17209,N_17223);
nand U17632 (N_17632,N_17387,N_17130);
xnor U17633 (N_17633,N_17378,N_17128);
or U17634 (N_17634,N_17372,N_17132);
nand U17635 (N_17635,N_17289,N_17291);
nand U17636 (N_17636,N_17257,N_17142);
xnor U17637 (N_17637,N_17189,N_17259);
nand U17638 (N_17638,N_17237,N_17175);
xor U17639 (N_17639,N_17354,N_17324);
and U17640 (N_17640,N_17163,N_17216);
nor U17641 (N_17641,N_17350,N_17243);
nand U17642 (N_17642,N_17112,N_17321);
and U17643 (N_17643,N_17145,N_17187);
nand U17644 (N_17644,N_17215,N_17290);
nor U17645 (N_17645,N_17339,N_17263);
xor U17646 (N_17646,N_17301,N_17368);
xor U17647 (N_17647,N_17107,N_17300);
nand U17648 (N_17648,N_17370,N_17376);
nand U17649 (N_17649,N_17222,N_17387);
or U17650 (N_17650,N_17270,N_17197);
nor U17651 (N_17651,N_17138,N_17109);
and U17652 (N_17652,N_17326,N_17156);
nand U17653 (N_17653,N_17226,N_17212);
or U17654 (N_17654,N_17301,N_17243);
nand U17655 (N_17655,N_17283,N_17322);
nor U17656 (N_17656,N_17142,N_17190);
or U17657 (N_17657,N_17295,N_17371);
nand U17658 (N_17658,N_17329,N_17233);
and U17659 (N_17659,N_17268,N_17168);
xor U17660 (N_17660,N_17391,N_17390);
nor U17661 (N_17661,N_17350,N_17337);
nor U17662 (N_17662,N_17293,N_17245);
and U17663 (N_17663,N_17341,N_17362);
nor U17664 (N_17664,N_17211,N_17235);
nor U17665 (N_17665,N_17174,N_17170);
or U17666 (N_17666,N_17186,N_17175);
and U17667 (N_17667,N_17229,N_17365);
nor U17668 (N_17668,N_17231,N_17369);
and U17669 (N_17669,N_17208,N_17137);
nor U17670 (N_17670,N_17334,N_17221);
nor U17671 (N_17671,N_17245,N_17233);
nor U17672 (N_17672,N_17101,N_17106);
nand U17673 (N_17673,N_17203,N_17136);
and U17674 (N_17674,N_17297,N_17317);
or U17675 (N_17675,N_17156,N_17147);
and U17676 (N_17676,N_17367,N_17188);
or U17677 (N_17677,N_17159,N_17320);
nand U17678 (N_17678,N_17323,N_17165);
xnor U17679 (N_17679,N_17394,N_17270);
nor U17680 (N_17680,N_17108,N_17301);
or U17681 (N_17681,N_17264,N_17222);
nor U17682 (N_17682,N_17251,N_17198);
nor U17683 (N_17683,N_17252,N_17306);
and U17684 (N_17684,N_17244,N_17399);
nand U17685 (N_17685,N_17271,N_17327);
nor U17686 (N_17686,N_17212,N_17125);
or U17687 (N_17687,N_17246,N_17277);
nand U17688 (N_17688,N_17269,N_17382);
nor U17689 (N_17689,N_17375,N_17322);
xor U17690 (N_17690,N_17253,N_17194);
nand U17691 (N_17691,N_17165,N_17346);
and U17692 (N_17692,N_17271,N_17368);
xnor U17693 (N_17693,N_17357,N_17175);
or U17694 (N_17694,N_17384,N_17225);
or U17695 (N_17695,N_17200,N_17281);
nand U17696 (N_17696,N_17380,N_17178);
xnor U17697 (N_17697,N_17179,N_17289);
nor U17698 (N_17698,N_17298,N_17223);
nor U17699 (N_17699,N_17180,N_17318);
and U17700 (N_17700,N_17632,N_17580);
or U17701 (N_17701,N_17609,N_17436);
nand U17702 (N_17702,N_17534,N_17590);
and U17703 (N_17703,N_17622,N_17462);
nand U17704 (N_17704,N_17551,N_17434);
xor U17705 (N_17705,N_17600,N_17625);
or U17706 (N_17706,N_17550,N_17473);
nand U17707 (N_17707,N_17628,N_17476);
or U17708 (N_17708,N_17481,N_17682);
xnor U17709 (N_17709,N_17460,N_17468);
nand U17710 (N_17710,N_17688,N_17648);
or U17711 (N_17711,N_17491,N_17588);
and U17712 (N_17712,N_17418,N_17523);
nor U17713 (N_17713,N_17584,N_17664);
and U17714 (N_17714,N_17623,N_17451);
xnor U17715 (N_17715,N_17454,N_17558);
and U17716 (N_17716,N_17440,N_17638);
xnor U17717 (N_17717,N_17533,N_17446);
and U17718 (N_17718,N_17696,N_17575);
or U17719 (N_17719,N_17689,N_17641);
or U17720 (N_17720,N_17576,N_17517);
nand U17721 (N_17721,N_17514,N_17512);
nor U17722 (N_17722,N_17477,N_17643);
nand U17723 (N_17723,N_17634,N_17673);
or U17724 (N_17724,N_17698,N_17614);
or U17725 (N_17725,N_17570,N_17412);
xor U17726 (N_17726,N_17581,N_17408);
nor U17727 (N_17727,N_17589,N_17650);
nor U17728 (N_17728,N_17430,N_17453);
nand U17729 (N_17729,N_17545,N_17487);
or U17730 (N_17730,N_17478,N_17601);
nor U17731 (N_17731,N_17535,N_17630);
and U17732 (N_17732,N_17444,N_17616);
or U17733 (N_17733,N_17578,N_17555);
nor U17734 (N_17734,N_17539,N_17458);
and U17735 (N_17735,N_17680,N_17687);
or U17736 (N_17736,N_17642,N_17456);
nor U17737 (N_17737,N_17699,N_17407);
xnor U17738 (N_17738,N_17656,N_17571);
nor U17739 (N_17739,N_17668,N_17606);
nor U17740 (N_17740,N_17437,N_17654);
or U17741 (N_17741,N_17669,N_17567);
or U17742 (N_17742,N_17672,N_17431);
nand U17743 (N_17743,N_17474,N_17644);
xor U17744 (N_17744,N_17690,N_17537);
nor U17745 (N_17745,N_17646,N_17599);
or U17746 (N_17746,N_17586,N_17624);
nor U17747 (N_17747,N_17546,N_17647);
and U17748 (N_17748,N_17627,N_17611);
nand U17749 (N_17749,N_17679,N_17405);
and U17750 (N_17750,N_17513,N_17465);
xor U17751 (N_17751,N_17496,N_17631);
nor U17752 (N_17752,N_17621,N_17427);
nand U17753 (N_17753,N_17526,N_17694);
xnor U17754 (N_17754,N_17585,N_17564);
xor U17755 (N_17755,N_17484,N_17659);
or U17756 (N_17756,N_17629,N_17433);
xor U17757 (N_17757,N_17422,N_17490);
xor U17758 (N_17758,N_17470,N_17509);
or U17759 (N_17759,N_17489,N_17691);
nor U17760 (N_17760,N_17435,N_17596);
xnor U17761 (N_17761,N_17658,N_17613);
xor U17762 (N_17762,N_17676,N_17604);
nor U17763 (N_17763,N_17525,N_17561);
or U17764 (N_17764,N_17515,N_17665);
xnor U17765 (N_17765,N_17498,N_17423);
nand U17766 (N_17766,N_17442,N_17566);
nand U17767 (N_17767,N_17520,N_17404);
and U17768 (N_17768,N_17529,N_17615);
xor U17769 (N_17769,N_17527,N_17577);
nor U17770 (N_17770,N_17485,N_17602);
or U17771 (N_17771,N_17530,N_17552);
xor U17772 (N_17772,N_17417,N_17495);
nor U17773 (N_17773,N_17522,N_17677);
nand U17774 (N_17774,N_17536,N_17457);
nor U17775 (N_17775,N_17562,N_17544);
and U17776 (N_17776,N_17432,N_17540);
xor U17777 (N_17777,N_17678,N_17524);
nor U17778 (N_17778,N_17568,N_17637);
xnor U17779 (N_17779,N_17450,N_17573);
or U17780 (N_17780,N_17666,N_17508);
or U17781 (N_17781,N_17419,N_17612);
nor U17782 (N_17782,N_17411,N_17519);
and U17783 (N_17783,N_17420,N_17521);
nand U17784 (N_17784,N_17607,N_17582);
or U17785 (N_17785,N_17559,N_17603);
nor U17786 (N_17786,N_17429,N_17574);
xor U17787 (N_17787,N_17511,N_17506);
nor U17788 (N_17788,N_17510,N_17531);
nand U17789 (N_17789,N_17681,N_17488);
or U17790 (N_17790,N_17605,N_17693);
nor U17791 (N_17791,N_17499,N_17425);
nand U17792 (N_17792,N_17655,N_17504);
xnor U17793 (N_17793,N_17518,N_17402);
nand U17794 (N_17794,N_17594,N_17610);
or U17795 (N_17795,N_17501,N_17633);
or U17796 (N_17796,N_17595,N_17409);
nand U17797 (N_17797,N_17608,N_17507);
nand U17798 (N_17798,N_17414,N_17403);
and U17799 (N_17799,N_17572,N_17445);
xnor U17800 (N_17800,N_17439,N_17554);
and U17801 (N_17801,N_17416,N_17553);
and U17802 (N_17802,N_17401,N_17626);
and U17803 (N_17803,N_17466,N_17591);
or U17804 (N_17804,N_17410,N_17652);
and U17805 (N_17805,N_17653,N_17472);
nor U17806 (N_17806,N_17461,N_17593);
and U17807 (N_17807,N_17657,N_17528);
or U17808 (N_17808,N_17620,N_17479);
nor U17809 (N_17809,N_17421,N_17494);
and U17810 (N_17810,N_17547,N_17406);
and U17811 (N_17811,N_17426,N_17670);
or U17812 (N_17812,N_17438,N_17482);
or U17813 (N_17813,N_17449,N_17587);
or U17814 (N_17814,N_17463,N_17400);
or U17815 (N_17815,N_17492,N_17686);
nor U17816 (N_17816,N_17579,N_17549);
xnor U17817 (N_17817,N_17663,N_17471);
nor U17818 (N_17818,N_17480,N_17443);
nor U17819 (N_17819,N_17538,N_17448);
or U17820 (N_17820,N_17467,N_17660);
nor U17821 (N_17821,N_17542,N_17452);
and U17822 (N_17822,N_17532,N_17684);
and U17823 (N_17823,N_17556,N_17661);
nand U17824 (N_17824,N_17619,N_17428);
nor U17825 (N_17825,N_17563,N_17617);
xor U17826 (N_17826,N_17497,N_17685);
nand U17827 (N_17827,N_17635,N_17557);
or U17828 (N_17828,N_17667,N_17475);
or U17829 (N_17829,N_17505,N_17645);
and U17830 (N_17830,N_17565,N_17592);
and U17831 (N_17831,N_17692,N_17695);
or U17832 (N_17832,N_17493,N_17455);
and U17833 (N_17833,N_17483,N_17516);
and U17834 (N_17834,N_17674,N_17464);
nor U17835 (N_17835,N_17636,N_17598);
nand U17836 (N_17836,N_17503,N_17424);
or U17837 (N_17837,N_17469,N_17548);
nor U17838 (N_17838,N_17649,N_17569);
or U17839 (N_17839,N_17486,N_17459);
nor U17840 (N_17840,N_17597,N_17543);
and U17841 (N_17841,N_17671,N_17662);
and U17842 (N_17842,N_17697,N_17415);
xnor U17843 (N_17843,N_17413,N_17683);
nor U17844 (N_17844,N_17640,N_17583);
and U17845 (N_17845,N_17560,N_17541);
nand U17846 (N_17846,N_17500,N_17639);
xor U17847 (N_17847,N_17675,N_17441);
nor U17848 (N_17848,N_17447,N_17651);
nand U17849 (N_17849,N_17618,N_17502);
and U17850 (N_17850,N_17549,N_17530);
xor U17851 (N_17851,N_17643,N_17409);
and U17852 (N_17852,N_17620,N_17652);
and U17853 (N_17853,N_17624,N_17646);
xor U17854 (N_17854,N_17439,N_17657);
and U17855 (N_17855,N_17536,N_17567);
nor U17856 (N_17856,N_17452,N_17527);
or U17857 (N_17857,N_17656,N_17570);
xor U17858 (N_17858,N_17485,N_17498);
and U17859 (N_17859,N_17442,N_17679);
or U17860 (N_17860,N_17630,N_17565);
and U17861 (N_17861,N_17645,N_17551);
xor U17862 (N_17862,N_17666,N_17443);
xnor U17863 (N_17863,N_17538,N_17547);
nor U17864 (N_17864,N_17440,N_17625);
xor U17865 (N_17865,N_17505,N_17507);
nor U17866 (N_17866,N_17654,N_17561);
nor U17867 (N_17867,N_17615,N_17641);
xnor U17868 (N_17868,N_17417,N_17462);
or U17869 (N_17869,N_17688,N_17647);
nor U17870 (N_17870,N_17641,N_17404);
nor U17871 (N_17871,N_17604,N_17569);
nor U17872 (N_17872,N_17519,N_17652);
nand U17873 (N_17873,N_17459,N_17642);
nand U17874 (N_17874,N_17511,N_17406);
and U17875 (N_17875,N_17697,N_17677);
nand U17876 (N_17876,N_17567,N_17404);
or U17877 (N_17877,N_17695,N_17656);
or U17878 (N_17878,N_17526,N_17652);
xnor U17879 (N_17879,N_17643,N_17644);
or U17880 (N_17880,N_17451,N_17496);
or U17881 (N_17881,N_17627,N_17662);
nand U17882 (N_17882,N_17622,N_17570);
or U17883 (N_17883,N_17546,N_17525);
and U17884 (N_17884,N_17667,N_17650);
and U17885 (N_17885,N_17644,N_17601);
nand U17886 (N_17886,N_17629,N_17622);
xor U17887 (N_17887,N_17543,N_17439);
nor U17888 (N_17888,N_17668,N_17494);
and U17889 (N_17889,N_17503,N_17512);
or U17890 (N_17890,N_17696,N_17490);
and U17891 (N_17891,N_17468,N_17604);
nand U17892 (N_17892,N_17582,N_17619);
nor U17893 (N_17893,N_17546,N_17400);
or U17894 (N_17894,N_17449,N_17657);
nand U17895 (N_17895,N_17698,N_17575);
nand U17896 (N_17896,N_17521,N_17662);
and U17897 (N_17897,N_17629,N_17554);
nand U17898 (N_17898,N_17484,N_17554);
nor U17899 (N_17899,N_17576,N_17692);
nand U17900 (N_17900,N_17601,N_17629);
or U17901 (N_17901,N_17693,N_17513);
nor U17902 (N_17902,N_17653,N_17630);
xor U17903 (N_17903,N_17484,N_17439);
and U17904 (N_17904,N_17614,N_17624);
xor U17905 (N_17905,N_17468,N_17538);
and U17906 (N_17906,N_17623,N_17619);
or U17907 (N_17907,N_17643,N_17423);
xor U17908 (N_17908,N_17555,N_17400);
nor U17909 (N_17909,N_17553,N_17578);
and U17910 (N_17910,N_17534,N_17617);
nand U17911 (N_17911,N_17451,N_17412);
nor U17912 (N_17912,N_17685,N_17467);
xnor U17913 (N_17913,N_17505,N_17418);
xnor U17914 (N_17914,N_17532,N_17675);
nand U17915 (N_17915,N_17645,N_17585);
xor U17916 (N_17916,N_17445,N_17497);
and U17917 (N_17917,N_17599,N_17585);
or U17918 (N_17918,N_17557,N_17657);
and U17919 (N_17919,N_17573,N_17697);
nand U17920 (N_17920,N_17489,N_17539);
xnor U17921 (N_17921,N_17408,N_17563);
or U17922 (N_17922,N_17508,N_17676);
and U17923 (N_17923,N_17493,N_17462);
nand U17924 (N_17924,N_17448,N_17529);
nand U17925 (N_17925,N_17657,N_17525);
or U17926 (N_17926,N_17467,N_17684);
nor U17927 (N_17927,N_17400,N_17418);
or U17928 (N_17928,N_17452,N_17671);
or U17929 (N_17929,N_17696,N_17619);
nand U17930 (N_17930,N_17450,N_17605);
or U17931 (N_17931,N_17616,N_17663);
or U17932 (N_17932,N_17589,N_17593);
or U17933 (N_17933,N_17531,N_17675);
nand U17934 (N_17934,N_17611,N_17557);
nand U17935 (N_17935,N_17679,N_17430);
or U17936 (N_17936,N_17424,N_17415);
and U17937 (N_17937,N_17532,N_17448);
nor U17938 (N_17938,N_17458,N_17642);
nor U17939 (N_17939,N_17593,N_17569);
and U17940 (N_17940,N_17486,N_17673);
and U17941 (N_17941,N_17560,N_17645);
or U17942 (N_17942,N_17614,N_17449);
or U17943 (N_17943,N_17606,N_17629);
nor U17944 (N_17944,N_17438,N_17574);
nand U17945 (N_17945,N_17504,N_17503);
nand U17946 (N_17946,N_17400,N_17563);
nand U17947 (N_17947,N_17520,N_17496);
xor U17948 (N_17948,N_17538,N_17459);
xnor U17949 (N_17949,N_17519,N_17511);
or U17950 (N_17950,N_17457,N_17414);
xor U17951 (N_17951,N_17436,N_17502);
or U17952 (N_17952,N_17649,N_17686);
and U17953 (N_17953,N_17482,N_17694);
or U17954 (N_17954,N_17497,N_17627);
nand U17955 (N_17955,N_17540,N_17469);
nor U17956 (N_17956,N_17464,N_17488);
and U17957 (N_17957,N_17434,N_17680);
nand U17958 (N_17958,N_17658,N_17519);
and U17959 (N_17959,N_17628,N_17555);
nor U17960 (N_17960,N_17662,N_17468);
xor U17961 (N_17961,N_17474,N_17555);
xor U17962 (N_17962,N_17658,N_17402);
nand U17963 (N_17963,N_17651,N_17547);
nand U17964 (N_17964,N_17429,N_17683);
and U17965 (N_17965,N_17545,N_17470);
xor U17966 (N_17966,N_17465,N_17563);
xnor U17967 (N_17967,N_17603,N_17518);
nor U17968 (N_17968,N_17551,N_17693);
nor U17969 (N_17969,N_17627,N_17539);
and U17970 (N_17970,N_17569,N_17631);
or U17971 (N_17971,N_17535,N_17686);
and U17972 (N_17972,N_17611,N_17581);
and U17973 (N_17973,N_17450,N_17456);
and U17974 (N_17974,N_17432,N_17682);
and U17975 (N_17975,N_17482,N_17567);
and U17976 (N_17976,N_17653,N_17623);
nor U17977 (N_17977,N_17472,N_17470);
and U17978 (N_17978,N_17543,N_17505);
and U17979 (N_17979,N_17532,N_17582);
nor U17980 (N_17980,N_17555,N_17448);
or U17981 (N_17981,N_17444,N_17539);
nor U17982 (N_17982,N_17631,N_17663);
or U17983 (N_17983,N_17641,N_17585);
or U17984 (N_17984,N_17637,N_17573);
nand U17985 (N_17985,N_17511,N_17473);
nor U17986 (N_17986,N_17613,N_17441);
nand U17987 (N_17987,N_17648,N_17503);
nand U17988 (N_17988,N_17475,N_17699);
or U17989 (N_17989,N_17624,N_17420);
or U17990 (N_17990,N_17661,N_17465);
xnor U17991 (N_17991,N_17528,N_17488);
nor U17992 (N_17992,N_17663,N_17698);
nor U17993 (N_17993,N_17634,N_17455);
or U17994 (N_17994,N_17501,N_17512);
or U17995 (N_17995,N_17539,N_17459);
and U17996 (N_17996,N_17636,N_17594);
nor U17997 (N_17997,N_17614,N_17699);
nand U17998 (N_17998,N_17425,N_17691);
xnor U17999 (N_17999,N_17659,N_17531);
xnor U18000 (N_18000,N_17805,N_17761);
or U18001 (N_18001,N_17791,N_17881);
or U18002 (N_18002,N_17922,N_17891);
and U18003 (N_18003,N_17931,N_17840);
xor U18004 (N_18004,N_17837,N_17726);
xor U18005 (N_18005,N_17818,N_17755);
xnor U18006 (N_18006,N_17720,N_17975);
nand U18007 (N_18007,N_17819,N_17820);
xor U18008 (N_18008,N_17950,N_17816);
xor U18009 (N_18009,N_17776,N_17885);
or U18010 (N_18010,N_17804,N_17844);
and U18011 (N_18011,N_17879,N_17759);
xnor U18012 (N_18012,N_17800,N_17893);
nand U18013 (N_18013,N_17972,N_17809);
xor U18014 (N_18014,N_17769,N_17980);
xnor U18015 (N_18015,N_17849,N_17751);
xnor U18016 (N_18016,N_17926,N_17727);
nor U18017 (N_18017,N_17841,N_17990);
nand U18018 (N_18018,N_17827,N_17864);
or U18019 (N_18019,N_17780,N_17721);
and U18020 (N_18020,N_17803,N_17850);
xnor U18021 (N_18021,N_17875,N_17775);
and U18022 (N_18022,N_17882,N_17843);
or U18023 (N_18023,N_17883,N_17963);
or U18024 (N_18024,N_17758,N_17917);
or U18025 (N_18025,N_17982,N_17874);
and U18026 (N_18026,N_17942,N_17929);
or U18027 (N_18027,N_17734,N_17838);
nand U18028 (N_18028,N_17733,N_17738);
nand U18029 (N_18029,N_17984,N_17872);
nand U18030 (N_18030,N_17862,N_17983);
nand U18031 (N_18031,N_17719,N_17877);
and U18032 (N_18032,N_17953,N_17900);
or U18033 (N_18033,N_17787,N_17810);
xnor U18034 (N_18034,N_17979,N_17814);
and U18035 (N_18035,N_17997,N_17770);
and U18036 (N_18036,N_17924,N_17796);
xor U18037 (N_18037,N_17960,N_17913);
xor U18038 (N_18038,N_17868,N_17940);
nand U18039 (N_18039,N_17936,N_17866);
nand U18040 (N_18040,N_17763,N_17869);
nor U18041 (N_18041,N_17833,N_17895);
and U18042 (N_18042,N_17873,N_17732);
or U18043 (N_18043,N_17836,N_17978);
nor U18044 (N_18044,N_17863,N_17949);
xnor U18045 (N_18045,N_17903,N_17861);
xnor U18046 (N_18046,N_17966,N_17959);
nor U18047 (N_18047,N_17757,N_17899);
nor U18048 (N_18048,N_17944,N_17933);
xor U18049 (N_18049,N_17886,N_17888);
or U18050 (N_18050,N_17789,N_17909);
and U18051 (N_18051,N_17845,N_17867);
xnor U18052 (N_18052,N_17930,N_17773);
nor U18053 (N_18053,N_17858,N_17756);
nor U18054 (N_18054,N_17825,N_17945);
or U18055 (N_18055,N_17928,N_17737);
and U18056 (N_18056,N_17852,N_17829);
nor U18057 (N_18057,N_17961,N_17938);
nor U18058 (N_18058,N_17896,N_17764);
nor U18059 (N_18059,N_17815,N_17923);
or U18060 (N_18060,N_17707,N_17958);
nor U18061 (N_18061,N_17906,N_17907);
xnor U18062 (N_18062,N_17914,N_17817);
xor U18063 (N_18063,N_17854,N_17821);
nor U18064 (N_18064,N_17797,N_17855);
xor U18065 (N_18065,N_17976,N_17918);
nand U18066 (N_18066,N_17932,N_17702);
xnor U18067 (N_18067,N_17740,N_17799);
nor U18068 (N_18068,N_17842,N_17973);
xnor U18069 (N_18069,N_17847,N_17794);
nor U18070 (N_18070,N_17952,N_17880);
and U18071 (N_18071,N_17822,N_17742);
xnor U18072 (N_18072,N_17813,N_17772);
nor U18073 (N_18073,N_17722,N_17736);
nand U18074 (N_18074,N_17934,N_17856);
and U18075 (N_18075,N_17999,N_17743);
xnor U18076 (N_18076,N_17898,N_17714);
or U18077 (N_18077,N_17835,N_17729);
or U18078 (N_18078,N_17920,N_17993);
nor U18079 (N_18079,N_17712,N_17853);
xor U18080 (N_18080,N_17807,N_17746);
and U18081 (N_18081,N_17904,N_17956);
xnor U18082 (N_18082,N_17860,N_17996);
and U18083 (N_18083,N_17705,N_17752);
or U18084 (N_18084,N_17741,N_17781);
or U18085 (N_18085,N_17970,N_17765);
xor U18086 (N_18086,N_17750,N_17901);
and U18087 (N_18087,N_17992,N_17967);
xnor U18088 (N_18088,N_17995,N_17801);
nor U18089 (N_18089,N_17774,N_17778);
nand U18090 (N_18090,N_17859,N_17890);
xnor U18091 (N_18091,N_17725,N_17795);
xor U18092 (N_18092,N_17783,N_17985);
and U18093 (N_18093,N_17782,N_17998);
or U18094 (N_18094,N_17991,N_17784);
nand U18095 (N_18095,N_17941,N_17724);
and U18096 (N_18096,N_17768,N_17710);
and U18097 (N_18097,N_17912,N_17921);
or U18098 (N_18098,N_17925,N_17718);
nor U18099 (N_18099,N_17777,N_17723);
xnor U18100 (N_18100,N_17955,N_17908);
nand U18101 (N_18101,N_17951,N_17897);
xnor U18102 (N_18102,N_17851,N_17968);
or U18103 (N_18103,N_17793,N_17711);
nor U18104 (N_18104,N_17839,N_17911);
and U18105 (N_18105,N_17716,N_17962);
nand U18106 (N_18106,N_17760,N_17971);
and U18107 (N_18107,N_17965,N_17754);
or U18108 (N_18108,N_17703,N_17969);
nor U18109 (N_18109,N_17905,N_17964);
xor U18110 (N_18110,N_17748,N_17876);
nor U18111 (N_18111,N_17808,N_17878);
nand U18112 (N_18112,N_17834,N_17739);
and U18113 (N_18113,N_17954,N_17857);
nor U18114 (N_18114,N_17802,N_17826);
or U18115 (N_18115,N_17828,N_17701);
nand U18116 (N_18116,N_17749,N_17987);
or U18117 (N_18117,N_17846,N_17977);
xnor U18118 (N_18118,N_17700,N_17994);
nand U18119 (N_18119,N_17943,N_17871);
or U18120 (N_18120,N_17715,N_17811);
and U18121 (N_18121,N_17870,N_17766);
xnor U18122 (N_18122,N_17947,N_17989);
and U18123 (N_18123,N_17779,N_17708);
xor U18124 (N_18124,N_17919,N_17824);
nand U18125 (N_18125,N_17704,N_17884);
or U18126 (N_18126,N_17894,N_17798);
or U18127 (N_18127,N_17935,N_17974);
xor U18128 (N_18128,N_17753,N_17910);
nand U18129 (N_18129,N_17713,N_17823);
and U18130 (N_18130,N_17915,N_17788);
xnor U18131 (N_18131,N_17717,N_17986);
or U18132 (N_18132,N_17830,N_17709);
or U18133 (N_18133,N_17939,N_17735);
nor U18134 (N_18134,N_17790,N_17771);
nor U18135 (N_18135,N_17948,N_17731);
or U18136 (N_18136,N_17706,N_17745);
or U18137 (N_18137,N_17937,N_17730);
nor U18138 (N_18138,N_17848,N_17762);
and U18139 (N_18139,N_17767,N_17792);
and U18140 (N_18140,N_17865,N_17887);
xor U18141 (N_18141,N_17744,N_17831);
nand U18142 (N_18142,N_17892,N_17806);
and U18143 (N_18143,N_17988,N_17981);
and U18144 (N_18144,N_17728,N_17902);
nor U18145 (N_18145,N_17957,N_17927);
and U18146 (N_18146,N_17747,N_17916);
nand U18147 (N_18147,N_17946,N_17832);
nor U18148 (N_18148,N_17786,N_17889);
and U18149 (N_18149,N_17785,N_17812);
and U18150 (N_18150,N_17807,N_17725);
and U18151 (N_18151,N_17931,N_17924);
nand U18152 (N_18152,N_17849,N_17760);
nor U18153 (N_18153,N_17877,N_17873);
or U18154 (N_18154,N_17729,N_17952);
or U18155 (N_18155,N_17736,N_17849);
nand U18156 (N_18156,N_17733,N_17776);
and U18157 (N_18157,N_17813,N_17842);
nor U18158 (N_18158,N_17709,N_17715);
nor U18159 (N_18159,N_17735,N_17846);
nor U18160 (N_18160,N_17936,N_17998);
xnor U18161 (N_18161,N_17838,N_17760);
and U18162 (N_18162,N_17999,N_17831);
xnor U18163 (N_18163,N_17997,N_17900);
nor U18164 (N_18164,N_17918,N_17820);
xor U18165 (N_18165,N_17725,N_17836);
nor U18166 (N_18166,N_17794,N_17826);
nor U18167 (N_18167,N_17811,N_17718);
or U18168 (N_18168,N_17725,N_17790);
and U18169 (N_18169,N_17808,N_17783);
xnor U18170 (N_18170,N_17718,N_17829);
and U18171 (N_18171,N_17710,N_17938);
nor U18172 (N_18172,N_17901,N_17707);
nand U18173 (N_18173,N_17789,N_17839);
or U18174 (N_18174,N_17738,N_17976);
nor U18175 (N_18175,N_17765,N_17933);
nand U18176 (N_18176,N_17951,N_17962);
nand U18177 (N_18177,N_17870,N_17989);
or U18178 (N_18178,N_17800,N_17980);
or U18179 (N_18179,N_17939,N_17760);
nand U18180 (N_18180,N_17926,N_17766);
or U18181 (N_18181,N_17971,N_17849);
nand U18182 (N_18182,N_17769,N_17715);
or U18183 (N_18183,N_17816,N_17850);
nor U18184 (N_18184,N_17991,N_17947);
and U18185 (N_18185,N_17735,N_17837);
nand U18186 (N_18186,N_17944,N_17836);
xor U18187 (N_18187,N_17750,N_17852);
and U18188 (N_18188,N_17742,N_17845);
and U18189 (N_18189,N_17705,N_17868);
nor U18190 (N_18190,N_17763,N_17707);
or U18191 (N_18191,N_17952,N_17985);
nor U18192 (N_18192,N_17939,N_17927);
nor U18193 (N_18193,N_17730,N_17978);
xor U18194 (N_18194,N_17970,N_17877);
nand U18195 (N_18195,N_17985,N_17778);
nor U18196 (N_18196,N_17737,N_17900);
nor U18197 (N_18197,N_17917,N_17797);
or U18198 (N_18198,N_17729,N_17807);
or U18199 (N_18199,N_17709,N_17739);
nand U18200 (N_18200,N_17756,N_17853);
nor U18201 (N_18201,N_17873,N_17711);
and U18202 (N_18202,N_17807,N_17799);
or U18203 (N_18203,N_17947,N_17820);
and U18204 (N_18204,N_17952,N_17980);
or U18205 (N_18205,N_17796,N_17704);
nand U18206 (N_18206,N_17715,N_17755);
or U18207 (N_18207,N_17987,N_17865);
nand U18208 (N_18208,N_17777,N_17911);
and U18209 (N_18209,N_17739,N_17991);
nor U18210 (N_18210,N_17957,N_17727);
nor U18211 (N_18211,N_17921,N_17833);
xor U18212 (N_18212,N_17973,N_17717);
and U18213 (N_18213,N_17878,N_17711);
nor U18214 (N_18214,N_17836,N_17893);
xnor U18215 (N_18215,N_17715,N_17784);
xnor U18216 (N_18216,N_17864,N_17917);
and U18217 (N_18217,N_17846,N_17853);
or U18218 (N_18218,N_17979,N_17864);
xor U18219 (N_18219,N_17956,N_17962);
nand U18220 (N_18220,N_17791,N_17931);
or U18221 (N_18221,N_17735,N_17762);
nor U18222 (N_18222,N_17729,N_17997);
nor U18223 (N_18223,N_17904,N_17884);
xor U18224 (N_18224,N_17961,N_17732);
nand U18225 (N_18225,N_17859,N_17711);
xnor U18226 (N_18226,N_17816,N_17776);
xor U18227 (N_18227,N_17855,N_17803);
and U18228 (N_18228,N_17717,N_17731);
nand U18229 (N_18229,N_17898,N_17777);
nand U18230 (N_18230,N_17768,N_17987);
nor U18231 (N_18231,N_17997,N_17941);
and U18232 (N_18232,N_17812,N_17885);
and U18233 (N_18233,N_17711,N_17918);
or U18234 (N_18234,N_17984,N_17750);
or U18235 (N_18235,N_17939,N_17738);
and U18236 (N_18236,N_17734,N_17750);
xnor U18237 (N_18237,N_17929,N_17879);
and U18238 (N_18238,N_17733,N_17990);
xor U18239 (N_18239,N_17783,N_17737);
and U18240 (N_18240,N_17821,N_17870);
or U18241 (N_18241,N_17812,N_17842);
and U18242 (N_18242,N_17852,N_17886);
and U18243 (N_18243,N_17867,N_17943);
or U18244 (N_18244,N_17724,N_17968);
and U18245 (N_18245,N_17976,N_17729);
nor U18246 (N_18246,N_17710,N_17708);
or U18247 (N_18247,N_17854,N_17749);
xnor U18248 (N_18248,N_17797,N_17836);
nor U18249 (N_18249,N_17984,N_17714);
nand U18250 (N_18250,N_17881,N_17730);
xnor U18251 (N_18251,N_17856,N_17700);
and U18252 (N_18252,N_17931,N_17780);
or U18253 (N_18253,N_17737,N_17802);
nor U18254 (N_18254,N_17937,N_17762);
and U18255 (N_18255,N_17763,N_17790);
nand U18256 (N_18256,N_17915,N_17980);
or U18257 (N_18257,N_17913,N_17847);
nand U18258 (N_18258,N_17736,N_17738);
xor U18259 (N_18259,N_17774,N_17927);
xnor U18260 (N_18260,N_17977,N_17747);
or U18261 (N_18261,N_17890,N_17711);
nand U18262 (N_18262,N_17788,N_17787);
nand U18263 (N_18263,N_17951,N_17790);
and U18264 (N_18264,N_17705,N_17884);
nor U18265 (N_18265,N_17800,N_17845);
nand U18266 (N_18266,N_17989,N_17863);
nand U18267 (N_18267,N_17952,N_17827);
xnor U18268 (N_18268,N_17726,N_17788);
nor U18269 (N_18269,N_17753,N_17740);
nand U18270 (N_18270,N_17924,N_17854);
or U18271 (N_18271,N_17884,N_17767);
xor U18272 (N_18272,N_17748,N_17824);
xnor U18273 (N_18273,N_17890,N_17718);
nor U18274 (N_18274,N_17978,N_17718);
nand U18275 (N_18275,N_17905,N_17878);
and U18276 (N_18276,N_17848,N_17733);
and U18277 (N_18277,N_17762,N_17717);
nor U18278 (N_18278,N_17714,N_17873);
nand U18279 (N_18279,N_17794,N_17969);
and U18280 (N_18280,N_17965,N_17955);
nand U18281 (N_18281,N_17823,N_17832);
and U18282 (N_18282,N_17778,N_17787);
and U18283 (N_18283,N_17954,N_17761);
and U18284 (N_18284,N_17922,N_17986);
nand U18285 (N_18285,N_17739,N_17848);
or U18286 (N_18286,N_17807,N_17901);
xnor U18287 (N_18287,N_17918,N_17809);
nor U18288 (N_18288,N_17906,N_17735);
nand U18289 (N_18289,N_17770,N_17976);
nor U18290 (N_18290,N_17997,N_17747);
and U18291 (N_18291,N_17713,N_17717);
or U18292 (N_18292,N_17979,N_17966);
and U18293 (N_18293,N_17906,N_17749);
nand U18294 (N_18294,N_17968,N_17707);
nand U18295 (N_18295,N_17728,N_17999);
and U18296 (N_18296,N_17766,N_17732);
xor U18297 (N_18297,N_17952,N_17783);
nand U18298 (N_18298,N_17944,N_17758);
xor U18299 (N_18299,N_17843,N_17840);
and U18300 (N_18300,N_18069,N_18125);
xnor U18301 (N_18301,N_18131,N_18263);
or U18302 (N_18302,N_18232,N_18193);
nand U18303 (N_18303,N_18240,N_18246);
nand U18304 (N_18304,N_18067,N_18118);
nor U18305 (N_18305,N_18064,N_18105);
nand U18306 (N_18306,N_18128,N_18152);
xnor U18307 (N_18307,N_18165,N_18060);
and U18308 (N_18308,N_18074,N_18268);
or U18309 (N_18309,N_18221,N_18151);
xnor U18310 (N_18310,N_18033,N_18110);
nand U18311 (N_18311,N_18279,N_18146);
and U18312 (N_18312,N_18199,N_18208);
or U18313 (N_18313,N_18140,N_18267);
nand U18314 (N_18314,N_18158,N_18298);
nor U18315 (N_18315,N_18266,N_18088);
or U18316 (N_18316,N_18015,N_18282);
or U18317 (N_18317,N_18028,N_18273);
nand U18318 (N_18318,N_18236,N_18106);
xor U18319 (N_18319,N_18117,N_18008);
xnor U18320 (N_18320,N_18150,N_18260);
nor U18321 (N_18321,N_18197,N_18164);
and U18322 (N_18322,N_18109,N_18253);
nor U18323 (N_18323,N_18233,N_18123);
and U18324 (N_18324,N_18144,N_18274);
nand U18325 (N_18325,N_18114,N_18042);
xor U18326 (N_18326,N_18120,N_18213);
nor U18327 (N_18327,N_18027,N_18061);
xnor U18328 (N_18328,N_18051,N_18284);
nand U18329 (N_18329,N_18133,N_18269);
and U18330 (N_18330,N_18116,N_18288);
and U18331 (N_18331,N_18254,N_18291);
or U18332 (N_18332,N_18024,N_18155);
nor U18333 (N_18333,N_18179,N_18041);
and U18334 (N_18334,N_18251,N_18026);
nand U18335 (N_18335,N_18075,N_18124);
and U18336 (N_18336,N_18135,N_18210);
or U18337 (N_18337,N_18001,N_18203);
or U18338 (N_18338,N_18290,N_18043);
xor U18339 (N_18339,N_18172,N_18245);
xnor U18340 (N_18340,N_18047,N_18270);
nor U18341 (N_18341,N_18002,N_18081);
or U18342 (N_18342,N_18272,N_18059);
or U18343 (N_18343,N_18077,N_18037);
nor U18344 (N_18344,N_18166,N_18091);
xor U18345 (N_18345,N_18046,N_18108);
nand U18346 (N_18346,N_18070,N_18154);
nor U18347 (N_18347,N_18055,N_18147);
or U18348 (N_18348,N_18045,N_18004);
or U18349 (N_18349,N_18080,N_18159);
xor U18350 (N_18350,N_18052,N_18247);
or U18351 (N_18351,N_18198,N_18177);
xnor U18352 (N_18352,N_18084,N_18050);
xnor U18353 (N_18353,N_18227,N_18073);
nand U18354 (N_18354,N_18217,N_18249);
nor U18355 (N_18355,N_18020,N_18185);
or U18356 (N_18356,N_18214,N_18293);
and U18357 (N_18357,N_18182,N_18107);
or U18358 (N_18358,N_18054,N_18286);
or U18359 (N_18359,N_18261,N_18030);
and U18360 (N_18360,N_18163,N_18257);
or U18361 (N_18361,N_18238,N_18053);
or U18362 (N_18362,N_18031,N_18202);
or U18363 (N_18363,N_18295,N_18259);
nor U18364 (N_18364,N_18013,N_18039);
nand U18365 (N_18365,N_18103,N_18014);
xnor U18366 (N_18366,N_18189,N_18100);
nor U18367 (N_18367,N_18289,N_18191);
and U18368 (N_18368,N_18275,N_18023);
or U18369 (N_18369,N_18256,N_18299);
or U18370 (N_18370,N_18048,N_18078);
nor U18371 (N_18371,N_18196,N_18137);
or U18372 (N_18372,N_18102,N_18089);
nand U18373 (N_18373,N_18250,N_18297);
or U18374 (N_18374,N_18220,N_18211);
nor U18375 (N_18375,N_18139,N_18072);
xor U18376 (N_18376,N_18243,N_18122);
nor U18377 (N_18377,N_18138,N_18223);
or U18378 (N_18378,N_18136,N_18248);
nor U18379 (N_18379,N_18255,N_18111);
xor U18380 (N_18380,N_18156,N_18113);
nand U18381 (N_18381,N_18285,N_18098);
nand U18382 (N_18382,N_18280,N_18090);
nor U18383 (N_18383,N_18175,N_18207);
or U18384 (N_18384,N_18206,N_18119);
nand U18385 (N_18385,N_18184,N_18085);
xor U18386 (N_18386,N_18034,N_18003);
xnor U18387 (N_18387,N_18180,N_18044);
xnor U18388 (N_18388,N_18019,N_18265);
xnor U18389 (N_18389,N_18036,N_18225);
and U18390 (N_18390,N_18239,N_18170);
xor U18391 (N_18391,N_18195,N_18230);
nor U18392 (N_18392,N_18021,N_18068);
nor U18393 (N_18393,N_18277,N_18010);
nand U18394 (N_18394,N_18216,N_18276);
xor U18395 (N_18395,N_18215,N_18160);
nor U18396 (N_18396,N_18148,N_18241);
and U18397 (N_18397,N_18174,N_18063);
or U18398 (N_18398,N_18095,N_18173);
and U18399 (N_18399,N_18244,N_18012);
and U18400 (N_18400,N_18000,N_18096);
nor U18401 (N_18401,N_18219,N_18205);
xor U18402 (N_18402,N_18121,N_18056);
or U18403 (N_18403,N_18262,N_18168);
and U18404 (N_18404,N_18129,N_18283);
nand U18405 (N_18405,N_18149,N_18005);
nor U18406 (N_18406,N_18018,N_18076);
or U18407 (N_18407,N_18082,N_18025);
and U18408 (N_18408,N_18192,N_18281);
nand U18409 (N_18409,N_18087,N_18200);
xnor U18410 (N_18410,N_18234,N_18242);
nor U18411 (N_18411,N_18093,N_18235);
nor U18412 (N_18412,N_18161,N_18181);
or U18413 (N_18413,N_18224,N_18186);
nand U18414 (N_18414,N_18127,N_18134);
xnor U18415 (N_18415,N_18141,N_18264);
nand U18416 (N_18416,N_18062,N_18058);
nor U18417 (N_18417,N_18112,N_18294);
nand U18418 (N_18418,N_18237,N_18066);
nand U18419 (N_18419,N_18097,N_18222);
and U18420 (N_18420,N_18083,N_18115);
and U18421 (N_18421,N_18187,N_18209);
or U18422 (N_18422,N_18029,N_18104);
and U18423 (N_18423,N_18292,N_18153);
or U18424 (N_18424,N_18201,N_18079);
or U18425 (N_18425,N_18065,N_18169);
or U18426 (N_18426,N_18092,N_18212);
and U18427 (N_18427,N_18218,N_18142);
nor U18428 (N_18428,N_18049,N_18130);
xor U18429 (N_18429,N_18162,N_18143);
xnor U18430 (N_18430,N_18094,N_18007);
nor U18431 (N_18431,N_18011,N_18229);
and U18432 (N_18432,N_18171,N_18017);
and U18433 (N_18433,N_18057,N_18016);
or U18434 (N_18434,N_18101,N_18271);
nor U18435 (N_18435,N_18157,N_18167);
nand U18436 (N_18436,N_18204,N_18178);
or U18437 (N_18437,N_18132,N_18190);
nand U18438 (N_18438,N_18258,N_18099);
or U18439 (N_18439,N_18022,N_18296);
or U18440 (N_18440,N_18086,N_18040);
nor U18441 (N_18441,N_18126,N_18252);
nand U18442 (N_18442,N_18009,N_18226);
nand U18443 (N_18443,N_18287,N_18231);
nor U18444 (N_18444,N_18278,N_18194);
nand U18445 (N_18445,N_18145,N_18183);
nor U18446 (N_18446,N_18188,N_18006);
xnor U18447 (N_18447,N_18176,N_18228);
xor U18448 (N_18448,N_18038,N_18071);
or U18449 (N_18449,N_18032,N_18035);
xnor U18450 (N_18450,N_18148,N_18209);
nor U18451 (N_18451,N_18128,N_18154);
nand U18452 (N_18452,N_18200,N_18101);
nand U18453 (N_18453,N_18115,N_18165);
and U18454 (N_18454,N_18207,N_18297);
xor U18455 (N_18455,N_18210,N_18077);
and U18456 (N_18456,N_18088,N_18046);
xor U18457 (N_18457,N_18019,N_18260);
nor U18458 (N_18458,N_18044,N_18177);
xor U18459 (N_18459,N_18069,N_18062);
or U18460 (N_18460,N_18182,N_18267);
nand U18461 (N_18461,N_18016,N_18284);
nor U18462 (N_18462,N_18055,N_18013);
nand U18463 (N_18463,N_18041,N_18280);
nand U18464 (N_18464,N_18205,N_18278);
xnor U18465 (N_18465,N_18003,N_18246);
nand U18466 (N_18466,N_18275,N_18026);
and U18467 (N_18467,N_18043,N_18194);
and U18468 (N_18468,N_18262,N_18008);
nor U18469 (N_18469,N_18271,N_18153);
or U18470 (N_18470,N_18122,N_18142);
nor U18471 (N_18471,N_18253,N_18288);
nand U18472 (N_18472,N_18113,N_18143);
and U18473 (N_18473,N_18251,N_18081);
xnor U18474 (N_18474,N_18293,N_18166);
and U18475 (N_18475,N_18144,N_18119);
or U18476 (N_18476,N_18286,N_18140);
or U18477 (N_18477,N_18014,N_18115);
or U18478 (N_18478,N_18013,N_18095);
nor U18479 (N_18479,N_18018,N_18202);
or U18480 (N_18480,N_18177,N_18235);
or U18481 (N_18481,N_18086,N_18275);
nor U18482 (N_18482,N_18265,N_18013);
xnor U18483 (N_18483,N_18138,N_18275);
nor U18484 (N_18484,N_18038,N_18215);
nor U18485 (N_18485,N_18055,N_18260);
or U18486 (N_18486,N_18179,N_18085);
or U18487 (N_18487,N_18176,N_18257);
nor U18488 (N_18488,N_18086,N_18206);
nand U18489 (N_18489,N_18034,N_18266);
nor U18490 (N_18490,N_18232,N_18069);
and U18491 (N_18491,N_18139,N_18171);
xor U18492 (N_18492,N_18266,N_18031);
xor U18493 (N_18493,N_18240,N_18260);
nand U18494 (N_18494,N_18176,N_18171);
and U18495 (N_18495,N_18288,N_18008);
nor U18496 (N_18496,N_18257,N_18195);
and U18497 (N_18497,N_18286,N_18275);
and U18498 (N_18498,N_18054,N_18240);
nor U18499 (N_18499,N_18237,N_18115);
and U18500 (N_18500,N_18227,N_18033);
and U18501 (N_18501,N_18275,N_18099);
or U18502 (N_18502,N_18198,N_18023);
or U18503 (N_18503,N_18013,N_18269);
nor U18504 (N_18504,N_18157,N_18103);
nand U18505 (N_18505,N_18125,N_18124);
nor U18506 (N_18506,N_18262,N_18134);
nor U18507 (N_18507,N_18124,N_18056);
xnor U18508 (N_18508,N_18099,N_18236);
nor U18509 (N_18509,N_18150,N_18096);
nand U18510 (N_18510,N_18054,N_18079);
and U18511 (N_18511,N_18232,N_18073);
nor U18512 (N_18512,N_18035,N_18052);
xnor U18513 (N_18513,N_18015,N_18250);
and U18514 (N_18514,N_18082,N_18213);
nor U18515 (N_18515,N_18191,N_18257);
xor U18516 (N_18516,N_18220,N_18099);
or U18517 (N_18517,N_18189,N_18185);
xnor U18518 (N_18518,N_18030,N_18086);
nand U18519 (N_18519,N_18215,N_18089);
nor U18520 (N_18520,N_18114,N_18235);
nand U18521 (N_18521,N_18055,N_18221);
or U18522 (N_18522,N_18201,N_18130);
nand U18523 (N_18523,N_18084,N_18091);
nand U18524 (N_18524,N_18118,N_18072);
and U18525 (N_18525,N_18189,N_18222);
and U18526 (N_18526,N_18080,N_18140);
or U18527 (N_18527,N_18007,N_18109);
nand U18528 (N_18528,N_18206,N_18298);
xnor U18529 (N_18529,N_18298,N_18100);
and U18530 (N_18530,N_18127,N_18226);
and U18531 (N_18531,N_18089,N_18063);
and U18532 (N_18532,N_18170,N_18225);
xnor U18533 (N_18533,N_18169,N_18211);
nor U18534 (N_18534,N_18267,N_18206);
xnor U18535 (N_18535,N_18164,N_18226);
or U18536 (N_18536,N_18170,N_18115);
and U18537 (N_18537,N_18050,N_18204);
and U18538 (N_18538,N_18026,N_18004);
and U18539 (N_18539,N_18277,N_18230);
xnor U18540 (N_18540,N_18217,N_18294);
nor U18541 (N_18541,N_18132,N_18162);
and U18542 (N_18542,N_18236,N_18223);
and U18543 (N_18543,N_18182,N_18098);
xor U18544 (N_18544,N_18132,N_18006);
or U18545 (N_18545,N_18009,N_18098);
nand U18546 (N_18546,N_18131,N_18108);
xor U18547 (N_18547,N_18185,N_18023);
nand U18548 (N_18548,N_18200,N_18076);
nor U18549 (N_18549,N_18252,N_18288);
nand U18550 (N_18550,N_18054,N_18209);
or U18551 (N_18551,N_18221,N_18059);
nand U18552 (N_18552,N_18153,N_18043);
nor U18553 (N_18553,N_18131,N_18140);
xnor U18554 (N_18554,N_18030,N_18178);
xnor U18555 (N_18555,N_18250,N_18201);
and U18556 (N_18556,N_18261,N_18134);
nor U18557 (N_18557,N_18248,N_18239);
nand U18558 (N_18558,N_18179,N_18116);
and U18559 (N_18559,N_18181,N_18091);
or U18560 (N_18560,N_18064,N_18107);
nor U18561 (N_18561,N_18056,N_18192);
and U18562 (N_18562,N_18284,N_18115);
nor U18563 (N_18563,N_18193,N_18046);
nor U18564 (N_18564,N_18107,N_18004);
or U18565 (N_18565,N_18266,N_18273);
and U18566 (N_18566,N_18155,N_18199);
nand U18567 (N_18567,N_18269,N_18076);
and U18568 (N_18568,N_18170,N_18180);
or U18569 (N_18569,N_18275,N_18098);
and U18570 (N_18570,N_18100,N_18082);
nand U18571 (N_18571,N_18118,N_18165);
xor U18572 (N_18572,N_18038,N_18015);
or U18573 (N_18573,N_18078,N_18132);
nand U18574 (N_18574,N_18178,N_18044);
nand U18575 (N_18575,N_18126,N_18032);
and U18576 (N_18576,N_18140,N_18218);
nor U18577 (N_18577,N_18013,N_18136);
xnor U18578 (N_18578,N_18107,N_18017);
and U18579 (N_18579,N_18130,N_18283);
xor U18580 (N_18580,N_18108,N_18283);
and U18581 (N_18581,N_18121,N_18123);
xnor U18582 (N_18582,N_18060,N_18270);
xnor U18583 (N_18583,N_18202,N_18102);
and U18584 (N_18584,N_18192,N_18193);
or U18585 (N_18585,N_18007,N_18044);
xor U18586 (N_18586,N_18095,N_18277);
nor U18587 (N_18587,N_18077,N_18082);
and U18588 (N_18588,N_18194,N_18002);
or U18589 (N_18589,N_18152,N_18201);
nor U18590 (N_18590,N_18257,N_18197);
nor U18591 (N_18591,N_18094,N_18204);
or U18592 (N_18592,N_18171,N_18222);
nor U18593 (N_18593,N_18092,N_18094);
nor U18594 (N_18594,N_18075,N_18120);
nor U18595 (N_18595,N_18270,N_18214);
xor U18596 (N_18596,N_18245,N_18088);
nor U18597 (N_18597,N_18193,N_18178);
or U18598 (N_18598,N_18126,N_18219);
nor U18599 (N_18599,N_18277,N_18023);
xnor U18600 (N_18600,N_18310,N_18303);
nand U18601 (N_18601,N_18319,N_18324);
xnor U18602 (N_18602,N_18387,N_18366);
nor U18603 (N_18603,N_18540,N_18521);
xnor U18604 (N_18604,N_18526,N_18318);
nor U18605 (N_18605,N_18321,N_18472);
and U18606 (N_18606,N_18300,N_18409);
or U18607 (N_18607,N_18452,N_18333);
xor U18608 (N_18608,N_18550,N_18408);
or U18609 (N_18609,N_18492,N_18523);
nand U18610 (N_18610,N_18505,N_18512);
nor U18611 (N_18611,N_18444,N_18528);
or U18612 (N_18612,N_18425,N_18468);
and U18613 (N_18613,N_18322,N_18500);
and U18614 (N_18614,N_18520,N_18377);
or U18615 (N_18615,N_18481,N_18384);
or U18616 (N_18616,N_18546,N_18317);
nand U18617 (N_18617,N_18419,N_18422);
and U18618 (N_18618,N_18595,N_18599);
nand U18619 (N_18619,N_18326,N_18517);
nand U18620 (N_18620,N_18421,N_18502);
or U18621 (N_18621,N_18372,N_18340);
or U18622 (N_18622,N_18399,N_18577);
and U18623 (N_18623,N_18455,N_18533);
or U18624 (N_18624,N_18557,N_18401);
or U18625 (N_18625,N_18510,N_18446);
xnor U18626 (N_18626,N_18493,N_18587);
nand U18627 (N_18627,N_18593,N_18436);
xnor U18628 (N_18628,N_18598,N_18487);
nand U18629 (N_18629,N_18556,N_18351);
xor U18630 (N_18630,N_18572,N_18494);
nor U18631 (N_18631,N_18416,N_18544);
or U18632 (N_18632,N_18365,N_18359);
nand U18633 (N_18633,N_18383,N_18462);
and U18634 (N_18634,N_18412,N_18463);
nand U18635 (N_18635,N_18323,N_18568);
nor U18636 (N_18636,N_18570,N_18552);
nand U18637 (N_18637,N_18439,N_18561);
and U18638 (N_18638,N_18539,N_18334);
nor U18639 (N_18639,N_18480,N_18591);
nand U18640 (N_18640,N_18543,N_18378);
xor U18641 (N_18641,N_18578,N_18508);
nor U18642 (N_18642,N_18574,N_18457);
or U18643 (N_18643,N_18414,N_18567);
nor U18644 (N_18644,N_18368,N_18315);
nand U18645 (N_18645,N_18395,N_18464);
and U18646 (N_18646,N_18306,N_18353);
and U18647 (N_18647,N_18375,N_18475);
nand U18648 (N_18648,N_18536,N_18537);
nor U18649 (N_18649,N_18553,N_18381);
and U18650 (N_18650,N_18542,N_18518);
nand U18651 (N_18651,N_18586,N_18346);
nand U18652 (N_18652,N_18435,N_18562);
and U18653 (N_18653,N_18428,N_18519);
nand U18654 (N_18654,N_18527,N_18358);
or U18655 (N_18655,N_18458,N_18332);
or U18656 (N_18656,N_18460,N_18573);
xnor U18657 (N_18657,N_18445,N_18491);
and U18658 (N_18658,N_18547,N_18569);
or U18659 (N_18659,N_18380,N_18382);
xnor U18660 (N_18660,N_18371,N_18486);
nor U18661 (N_18661,N_18459,N_18415);
nand U18662 (N_18662,N_18559,N_18476);
nand U18663 (N_18663,N_18406,N_18388);
and U18664 (N_18664,N_18427,N_18349);
nor U18665 (N_18665,N_18347,N_18585);
or U18666 (N_18666,N_18554,N_18442);
and U18667 (N_18667,N_18506,N_18563);
and U18668 (N_18668,N_18385,N_18434);
or U18669 (N_18669,N_18407,N_18311);
xor U18670 (N_18670,N_18483,N_18454);
nand U18671 (N_18671,N_18474,N_18379);
nand U18672 (N_18672,N_18431,N_18555);
nor U18673 (N_18673,N_18488,N_18529);
or U18674 (N_18674,N_18565,N_18350);
nand U18675 (N_18675,N_18558,N_18504);
and U18676 (N_18676,N_18440,N_18370);
xor U18677 (N_18677,N_18447,N_18309);
nor U18678 (N_18678,N_18496,N_18404);
xnor U18679 (N_18679,N_18479,N_18511);
and U18680 (N_18680,N_18339,N_18420);
and U18681 (N_18681,N_18551,N_18453);
nor U18682 (N_18682,N_18410,N_18451);
and U18683 (N_18683,N_18534,N_18423);
and U18684 (N_18684,N_18374,N_18352);
or U18685 (N_18685,N_18594,N_18345);
and U18686 (N_18686,N_18525,N_18413);
xor U18687 (N_18687,N_18485,N_18301);
nand U18688 (N_18688,N_18307,N_18325);
nor U18689 (N_18689,N_18432,N_18448);
xnor U18690 (N_18690,N_18582,N_18397);
and U18691 (N_18691,N_18348,N_18426);
nor U18692 (N_18692,N_18499,N_18584);
or U18693 (N_18693,N_18588,N_18418);
and U18694 (N_18694,N_18367,N_18336);
and U18695 (N_18695,N_18545,N_18361);
or U18696 (N_18696,N_18441,N_18342);
xor U18697 (N_18697,N_18597,N_18589);
nor U18698 (N_18698,N_18530,N_18338);
or U18699 (N_18699,N_18390,N_18386);
nand U18700 (N_18700,N_18327,N_18524);
nand U18701 (N_18701,N_18398,N_18564);
and U18702 (N_18702,N_18355,N_18514);
nand U18703 (N_18703,N_18424,N_18443);
nor U18704 (N_18704,N_18337,N_18509);
or U18705 (N_18705,N_18400,N_18373);
nor U18706 (N_18706,N_18531,N_18471);
nand U18707 (N_18707,N_18501,N_18590);
or U18708 (N_18708,N_18490,N_18362);
nor U18709 (N_18709,N_18579,N_18389);
or U18710 (N_18710,N_18391,N_18437);
or U18711 (N_18711,N_18308,N_18357);
xor U18712 (N_18712,N_18596,N_18592);
and U18713 (N_18713,N_18376,N_18576);
and U18714 (N_18714,N_18478,N_18438);
nor U18715 (N_18715,N_18394,N_18344);
or U18716 (N_18716,N_18302,N_18470);
nand U18717 (N_18717,N_18433,N_18417);
nand U18718 (N_18718,N_18316,N_18331);
nand U18719 (N_18719,N_18495,N_18360);
nor U18720 (N_18720,N_18330,N_18497);
and U18721 (N_18721,N_18449,N_18450);
nor U18722 (N_18722,N_18354,N_18364);
nor U18723 (N_18723,N_18484,N_18304);
and U18724 (N_18724,N_18467,N_18363);
xor U18725 (N_18725,N_18538,N_18393);
and U18726 (N_18726,N_18580,N_18411);
nand U18727 (N_18727,N_18305,N_18405);
or U18728 (N_18728,N_18516,N_18320);
or U18729 (N_18729,N_18313,N_18402);
or U18730 (N_18730,N_18403,N_18581);
nand U18731 (N_18731,N_18560,N_18312);
xor U18732 (N_18732,N_18532,N_18369);
nand U18733 (N_18733,N_18456,N_18548);
or U18734 (N_18734,N_18566,N_18461);
nand U18735 (N_18735,N_18515,N_18469);
and U18736 (N_18736,N_18477,N_18575);
nand U18737 (N_18737,N_18328,N_18507);
nand U18738 (N_18738,N_18356,N_18535);
nor U18739 (N_18739,N_18341,N_18335);
nor U18740 (N_18740,N_18473,N_18343);
nor U18741 (N_18741,N_18329,N_18498);
or U18742 (N_18742,N_18522,N_18466);
and U18743 (N_18743,N_18513,N_18541);
nand U18744 (N_18744,N_18482,N_18392);
and U18745 (N_18745,N_18396,N_18549);
or U18746 (N_18746,N_18314,N_18571);
nand U18747 (N_18747,N_18465,N_18430);
and U18748 (N_18748,N_18503,N_18489);
nand U18749 (N_18749,N_18583,N_18429);
and U18750 (N_18750,N_18416,N_18408);
and U18751 (N_18751,N_18368,N_18516);
nand U18752 (N_18752,N_18560,N_18398);
nor U18753 (N_18753,N_18447,N_18444);
and U18754 (N_18754,N_18412,N_18388);
and U18755 (N_18755,N_18499,N_18303);
nand U18756 (N_18756,N_18356,N_18504);
and U18757 (N_18757,N_18328,N_18409);
xnor U18758 (N_18758,N_18553,N_18508);
nand U18759 (N_18759,N_18430,N_18584);
or U18760 (N_18760,N_18501,N_18447);
or U18761 (N_18761,N_18328,N_18382);
and U18762 (N_18762,N_18358,N_18488);
xnor U18763 (N_18763,N_18549,N_18413);
or U18764 (N_18764,N_18559,N_18331);
and U18765 (N_18765,N_18536,N_18331);
nor U18766 (N_18766,N_18494,N_18396);
nand U18767 (N_18767,N_18597,N_18573);
or U18768 (N_18768,N_18581,N_18521);
or U18769 (N_18769,N_18535,N_18370);
and U18770 (N_18770,N_18491,N_18310);
or U18771 (N_18771,N_18334,N_18340);
nand U18772 (N_18772,N_18542,N_18599);
xor U18773 (N_18773,N_18466,N_18318);
nor U18774 (N_18774,N_18559,N_18585);
and U18775 (N_18775,N_18566,N_18353);
nand U18776 (N_18776,N_18376,N_18345);
nor U18777 (N_18777,N_18446,N_18440);
xnor U18778 (N_18778,N_18496,N_18543);
nand U18779 (N_18779,N_18409,N_18526);
or U18780 (N_18780,N_18306,N_18479);
xor U18781 (N_18781,N_18367,N_18352);
or U18782 (N_18782,N_18593,N_18451);
and U18783 (N_18783,N_18516,N_18558);
nand U18784 (N_18784,N_18358,N_18336);
xor U18785 (N_18785,N_18513,N_18301);
or U18786 (N_18786,N_18415,N_18377);
nand U18787 (N_18787,N_18446,N_18349);
and U18788 (N_18788,N_18345,N_18538);
and U18789 (N_18789,N_18325,N_18489);
or U18790 (N_18790,N_18420,N_18337);
and U18791 (N_18791,N_18329,N_18437);
nand U18792 (N_18792,N_18420,N_18511);
nand U18793 (N_18793,N_18441,N_18489);
nand U18794 (N_18794,N_18346,N_18356);
nand U18795 (N_18795,N_18484,N_18394);
nand U18796 (N_18796,N_18570,N_18487);
and U18797 (N_18797,N_18465,N_18354);
or U18798 (N_18798,N_18445,N_18312);
nor U18799 (N_18799,N_18510,N_18458);
nor U18800 (N_18800,N_18493,N_18597);
or U18801 (N_18801,N_18544,N_18494);
xor U18802 (N_18802,N_18572,N_18569);
or U18803 (N_18803,N_18504,N_18349);
xnor U18804 (N_18804,N_18590,N_18300);
nand U18805 (N_18805,N_18530,N_18353);
or U18806 (N_18806,N_18330,N_18381);
or U18807 (N_18807,N_18320,N_18401);
nor U18808 (N_18808,N_18356,N_18495);
nand U18809 (N_18809,N_18544,N_18503);
or U18810 (N_18810,N_18514,N_18361);
nor U18811 (N_18811,N_18412,N_18387);
or U18812 (N_18812,N_18499,N_18419);
and U18813 (N_18813,N_18508,N_18373);
and U18814 (N_18814,N_18552,N_18527);
nand U18815 (N_18815,N_18518,N_18544);
nand U18816 (N_18816,N_18590,N_18371);
or U18817 (N_18817,N_18374,N_18514);
xnor U18818 (N_18818,N_18394,N_18445);
or U18819 (N_18819,N_18543,N_18421);
nor U18820 (N_18820,N_18596,N_18477);
xor U18821 (N_18821,N_18446,N_18421);
or U18822 (N_18822,N_18319,N_18330);
and U18823 (N_18823,N_18571,N_18573);
nand U18824 (N_18824,N_18301,N_18328);
nor U18825 (N_18825,N_18412,N_18329);
nor U18826 (N_18826,N_18323,N_18437);
nand U18827 (N_18827,N_18420,N_18318);
nor U18828 (N_18828,N_18564,N_18510);
xnor U18829 (N_18829,N_18333,N_18495);
nand U18830 (N_18830,N_18322,N_18305);
or U18831 (N_18831,N_18490,N_18418);
xor U18832 (N_18832,N_18483,N_18418);
and U18833 (N_18833,N_18457,N_18414);
xnor U18834 (N_18834,N_18390,N_18548);
or U18835 (N_18835,N_18485,N_18591);
and U18836 (N_18836,N_18564,N_18368);
xnor U18837 (N_18837,N_18409,N_18540);
xnor U18838 (N_18838,N_18499,N_18358);
xor U18839 (N_18839,N_18349,N_18557);
nor U18840 (N_18840,N_18514,N_18496);
and U18841 (N_18841,N_18461,N_18487);
nand U18842 (N_18842,N_18441,N_18414);
nand U18843 (N_18843,N_18372,N_18344);
nand U18844 (N_18844,N_18592,N_18573);
or U18845 (N_18845,N_18446,N_18462);
or U18846 (N_18846,N_18347,N_18504);
nor U18847 (N_18847,N_18319,N_18471);
nand U18848 (N_18848,N_18501,N_18491);
xnor U18849 (N_18849,N_18548,N_18531);
xnor U18850 (N_18850,N_18560,N_18321);
and U18851 (N_18851,N_18444,N_18517);
nand U18852 (N_18852,N_18495,N_18346);
or U18853 (N_18853,N_18544,N_18469);
nor U18854 (N_18854,N_18326,N_18593);
nor U18855 (N_18855,N_18440,N_18360);
nor U18856 (N_18856,N_18423,N_18512);
nor U18857 (N_18857,N_18454,N_18373);
or U18858 (N_18858,N_18486,N_18482);
nor U18859 (N_18859,N_18344,N_18477);
nand U18860 (N_18860,N_18385,N_18345);
or U18861 (N_18861,N_18499,N_18466);
nand U18862 (N_18862,N_18513,N_18329);
nor U18863 (N_18863,N_18542,N_18480);
xnor U18864 (N_18864,N_18514,N_18426);
or U18865 (N_18865,N_18568,N_18500);
nor U18866 (N_18866,N_18527,N_18508);
xnor U18867 (N_18867,N_18515,N_18327);
nor U18868 (N_18868,N_18446,N_18410);
nor U18869 (N_18869,N_18429,N_18513);
nor U18870 (N_18870,N_18598,N_18471);
or U18871 (N_18871,N_18375,N_18302);
nor U18872 (N_18872,N_18502,N_18483);
nand U18873 (N_18873,N_18466,N_18463);
and U18874 (N_18874,N_18480,N_18433);
and U18875 (N_18875,N_18423,N_18396);
nand U18876 (N_18876,N_18597,N_18324);
xor U18877 (N_18877,N_18336,N_18570);
nor U18878 (N_18878,N_18371,N_18317);
or U18879 (N_18879,N_18563,N_18455);
xor U18880 (N_18880,N_18525,N_18498);
or U18881 (N_18881,N_18351,N_18542);
xnor U18882 (N_18882,N_18537,N_18524);
or U18883 (N_18883,N_18409,N_18437);
or U18884 (N_18884,N_18435,N_18355);
xnor U18885 (N_18885,N_18341,N_18348);
xnor U18886 (N_18886,N_18417,N_18325);
nor U18887 (N_18887,N_18399,N_18461);
nand U18888 (N_18888,N_18354,N_18462);
nor U18889 (N_18889,N_18481,N_18477);
and U18890 (N_18890,N_18590,N_18442);
and U18891 (N_18891,N_18392,N_18595);
xor U18892 (N_18892,N_18452,N_18449);
or U18893 (N_18893,N_18496,N_18570);
nand U18894 (N_18894,N_18553,N_18380);
nand U18895 (N_18895,N_18396,N_18485);
or U18896 (N_18896,N_18465,N_18486);
and U18897 (N_18897,N_18326,N_18300);
and U18898 (N_18898,N_18499,N_18420);
and U18899 (N_18899,N_18325,N_18526);
nor U18900 (N_18900,N_18784,N_18754);
or U18901 (N_18901,N_18771,N_18666);
and U18902 (N_18902,N_18787,N_18781);
and U18903 (N_18903,N_18821,N_18839);
nor U18904 (N_18904,N_18723,N_18841);
xor U18905 (N_18905,N_18664,N_18794);
or U18906 (N_18906,N_18637,N_18792);
nor U18907 (N_18907,N_18670,N_18716);
xor U18908 (N_18908,N_18634,N_18659);
and U18909 (N_18909,N_18882,N_18777);
and U18910 (N_18910,N_18818,N_18898);
xor U18911 (N_18911,N_18865,N_18826);
and U18912 (N_18912,N_18843,N_18791);
nand U18913 (N_18913,N_18662,N_18786);
or U18914 (N_18914,N_18851,N_18809);
nand U18915 (N_18915,N_18609,N_18628);
or U18916 (N_18916,N_18710,N_18744);
nor U18917 (N_18917,N_18601,N_18790);
nor U18918 (N_18918,N_18665,N_18864);
nor U18919 (N_18919,N_18735,N_18813);
and U18920 (N_18920,N_18630,N_18803);
and U18921 (N_18921,N_18772,N_18881);
or U18922 (N_18922,N_18890,N_18761);
nand U18923 (N_18923,N_18873,N_18859);
or U18924 (N_18924,N_18880,N_18681);
and U18925 (N_18925,N_18604,N_18731);
xnor U18926 (N_18926,N_18615,N_18708);
nand U18927 (N_18927,N_18696,N_18808);
nor U18928 (N_18928,N_18835,N_18600);
nor U18929 (N_18929,N_18752,N_18774);
nor U18930 (N_18930,N_18663,N_18636);
or U18931 (N_18931,N_18686,N_18698);
nor U18932 (N_18932,N_18769,N_18779);
nor U18933 (N_18933,N_18640,N_18718);
nand U18934 (N_18934,N_18825,N_18763);
and U18935 (N_18935,N_18672,N_18680);
xor U18936 (N_18936,N_18707,N_18610);
xnor U18937 (N_18937,N_18805,N_18627);
nor U18938 (N_18938,N_18837,N_18811);
or U18939 (N_18939,N_18776,N_18883);
nand U18940 (N_18940,N_18846,N_18678);
nand U18941 (N_18941,N_18612,N_18695);
xnor U18942 (N_18942,N_18651,N_18715);
and U18943 (N_18943,N_18667,N_18857);
or U18944 (N_18944,N_18607,N_18878);
and U18945 (N_18945,N_18732,N_18650);
nor U18946 (N_18946,N_18868,N_18709);
nor U18947 (N_18947,N_18747,N_18829);
nand U18948 (N_18948,N_18850,N_18814);
nand U18949 (N_18949,N_18861,N_18620);
nand U18950 (N_18950,N_18849,N_18757);
xnor U18951 (N_18951,N_18658,N_18778);
or U18952 (N_18952,N_18780,N_18720);
xor U18953 (N_18953,N_18797,N_18743);
nor U18954 (N_18954,N_18832,N_18783);
xnor U18955 (N_18955,N_18669,N_18704);
xnor U18956 (N_18956,N_18644,N_18834);
or U18957 (N_18957,N_18893,N_18891);
nand U18958 (N_18958,N_18674,N_18764);
nand U18959 (N_18959,N_18886,N_18828);
nand U18960 (N_18960,N_18657,N_18799);
or U18961 (N_18961,N_18765,N_18632);
and U18962 (N_18962,N_18758,N_18760);
and U18963 (N_18963,N_18848,N_18625);
nand U18964 (N_18964,N_18618,N_18817);
nand U18965 (N_18965,N_18639,N_18854);
nand U18966 (N_18966,N_18694,N_18894);
nor U18967 (N_18967,N_18616,N_18702);
nor U18968 (N_18968,N_18688,N_18840);
nor U18969 (N_18969,N_18654,N_18719);
nand U18970 (N_18970,N_18812,N_18671);
and U18971 (N_18971,N_18713,N_18806);
and U18972 (N_18972,N_18633,N_18673);
nand U18973 (N_18973,N_18860,N_18692);
xnor U18974 (N_18974,N_18833,N_18693);
or U18975 (N_18975,N_18807,N_18819);
or U18976 (N_18976,N_18823,N_18874);
xor U18977 (N_18977,N_18729,N_18802);
nor U18978 (N_18978,N_18676,N_18876);
xor U18979 (N_18979,N_18824,N_18721);
xor U18980 (N_18980,N_18816,N_18870);
xnor U18981 (N_18981,N_18614,N_18725);
nor U18982 (N_18982,N_18653,N_18888);
and U18983 (N_18983,N_18863,N_18796);
nor U18984 (N_18984,N_18629,N_18838);
nand U18985 (N_18985,N_18712,N_18768);
nor U18986 (N_18986,N_18800,N_18685);
and U18987 (N_18987,N_18603,N_18852);
or U18988 (N_18988,N_18897,N_18742);
and U18989 (N_18989,N_18617,N_18801);
and U18990 (N_18990,N_18677,N_18635);
and U18991 (N_18991,N_18879,N_18730);
nand U18992 (N_18992,N_18722,N_18741);
and U18993 (N_18993,N_18690,N_18853);
or U18994 (N_18994,N_18875,N_18782);
and U18995 (N_18995,N_18656,N_18668);
xnor U18996 (N_18996,N_18728,N_18645);
xnor U18997 (N_18997,N_18738,N_18682);
xor U18998 (N_18998,N_18827,N_18687);
xnor U18999 (N_18999,N_18711,N_18795);
nor U19000 (N_19000,N_18767,N_18844);
xnor U19001 (N_19001,N_18727,N_18847);
nand U19002 (N_19002,N_18641,N_18647);
and U19003 (N_19003,N_18867,N_18714);
nand U19004 (N_19004,N_18626,N_18624);
nand U19005 (N_19005,N_18749,N_18726);
and U19006 (N_19006,N_18788,N_18775);
and U19007 (N_19007,N_18745,N_18734);
xnor U19008 (N_19008,N_18798,N_18724);
or U19009 (N_19009,N_18820,N_18773);
and U19010 (N_19010,N_18733,N_18611);
and U19011 (N_19011,N_18700,N_18622);
or U19012 (N_19012,N_18691,N_18877);
and U19013 (N_19013,N_18643,N_18740);
xor U19014 (N_19014,N_18866,N_18871);
xor U19015 (N_19015,N_18646,N_18619);
and U19016 (N_19016,N_18856,N_18739);
and U19017 (N_19017,N_18648,N_18862);
nand U19018 (N_19018,N_18896,N_18751);
and U19019 (N_19019,N_18701,N_18683);
xnor U19020 (N_19020,N_18679,N_18815);
or U19021 (N_19021,N_18830,N_18705);
or U19022 (N_19022,N_18855,N_18858);
nand U19023 (N_19023,N_18613,N_18606);
or U19024 (N_19024,N_18810,N_18789);
and U19025 (N_19025,N_18785,N_18766);
nor U19026 (N_19026,N_18623,N_18621);
and U19027 (N_19027,N_18675,N_18869);
and U19028 (N_19028,N_18889,N_18884);
and U19029 (N_19029,N_18762,N_18697);
nor U19030 (N_19030,N_18699,N_18895);
xnor U19031 (N_19031,N_18887,N_18661);
xnor U19032 (N_19032,N_18649,N_18793);
nand U19033 (N_19033,N_18753,N_18605);
nand U19034 (N_19034,N_18842,N_18652);
or U19035 (N_19035,N_18885,N_18638);
xnor U19036 (N_19036,N_18759,N_18631);
nor U19037 (N_19037,N_18822,N_18736);
xor U19038 (N_19038,N_18750,N_18872);
or U19039 (N_19039,N_18703,N_18831);
or U19040 (N_19040,N_18737,N_18845);
nand U19041 (N_19041,N_18706,N_18642);
or U19042 (N_19042,N_18746,N_18756);
or U19043 (N_19043,N_18684,N_18804);
and U19044 (N_19044,N_18655,N_18755);
xnor U19045 (N_19045,N_18770,N_18892);
xnor U19046 (N_19046,N_18608,N_18689);
or U19047 (N_19047,N_18660,N_18717);
xnor U19048 (N_19048,N_18836,N_18748);
xnor U19049 (N_19049,N_18899,N_18602);
nand U19050 (N_19050,N_18844,N_18665);
or U19051 (N_19051,N_18789,N_18727);
or U19052 (N_19052,N_18824,N_18615);
nand U19053 (N_19053,N_18667,N_18825);
nor U19054 (N_19054,N_18729,N_18732);
nand U19055 (N_19055,N_18627,N_18658);
or U19056 (N_19056,N_18778,N_18846);
and U19057 (N_19057,N_18889,N_18612);
or U19058 (N_19058,N_18617,N_18711);
nand U19059 (N_19059,N_18854,N_18603);
nand U19060 (N_19060,N_18786,N_18790);
or U19061 (N_19061,N_18767,N_18635);
nor U19062 (N_19062,N_18868,N_18763);
nor U19063 (N_19063,N_18633,N_18702);
xnor U19064 (N_19064,N_18893,N_18682);
or U19065 (N_19065,N_18618,N_18699);
nand U19066 (N_19066,N_18897,N_18778);
nor U19067 (N_19067,N_18607,N_18742);
nand U19068 (N_19068,N_18753,N_18731);
xor U19069 (N_19069,N_18892,N_18876);
xor U19070 (N_19070,N_18646,N_18710);
xnor U19071 (N_19071,N_18702,N_18676);
xor U19072 (N_19072,N_18812,N_18869);
xnor U19073 (N_19073,N_18867,N_18835);
or U19074 (N_19074,N_18716,N_18867);
nor U19075 (N_19075,N_18845,N_18686);
and U19076 (N_19076,N_18803,N_18742);
xor U19077 (N_19077,N_18835,N_18877);
xnor U19078 (N_19078,N_18819,N_18788);
nor U19079 (N_19079,N_18767,N_18860);
xor U19080 (N_19080,N_18769,N_18768);
and U19081 (N_19081,N_18786,N_18645);
and U19082 (N_19082,N_18876,N_18617);
nor U19083 (N_19083,N_18886,N_18691);
nor U19084 (N_19084,N_18609,N_18860);
nor U19085 (N_19085,N_18836,N_18621);
nor U19086 (N_19086,N_18674,N_18754);
xnor U19087 (N_19087,N_18760,N_18668);
xor U19088 (N_19088,N_18665,N_18663);
nor U19089 (N_19089,N_18613,N_18886);
and U19090 (N_19090,N_18660,N_18645);
or U19091 (N_19091,N_18789,N_18833);
nor U19092 (N_19092,N_18783,N_18704);
and U19093 (N_19093,N_18655,N_18874);
nor U19094 (N_19094,N_18844,N_18840);
xnor U19095 (N_19095,N_18851,N_18844);
and U19096 (N_19096,N_18834,N_18709);
nand U19097 (N_19097,N_18766,N_18730);
and U19098 (N_19098,N_18624,N_18788);
nand U19099 (N_19099,N_18741,N_18672);
nor U19100 (N_19100,N_18689,N_18812);
or U19101 (N_19101,N_18820,N_18703);
xnor U19102 (N_19102,N_18644,N_18609);
and U19103 (N_19103,N_18878,N_18807);
nand U19104 (N_19104,N_18828,N_18743);
nand U19105 (N_19105,N_18779,N_18677);
nor U19106 (N_19106,N_18717,N_18821);
or U19107 (N_19107,N_18853,N_18606);
nand U19108 (N_19108,N_18606,N_18678);
or U19109 (N_19109,N_18772,N_18644);
nor U19110 (N_19110,N_18890,N_18618);
and U19111 (N_19111,N_18898,N_18617);
xor U19112 (N_19112,N_18781,N_18849);
nor U19113 (N_19113,N_18852,N_18736);
xor U19114 (N_19114,N_18675,N_18670);
nor U19115 (N_19115,N_18787,N_18637);
and U19116 (N_19116,N_18637,N_18706);
nand U19117 (N_19117,N_18874,N_18681);
or U19118 (N_19118,N_18806,N_18663);
or U19119 (N_19119,N_18838,N_18688);
nand U19120 (N_19120,N_18617,N_18699);
or U19121 (N_19121,N_18646,N_18888);
xnor U19122 (N_19122,N_18767,N_18770);
and U19123 (N_19123,N_18621,N_18693);
nor U19124 (N_19124,N_18702,N_18625);
nand U19125 (N_19125,N_18605,N_18869);
nand U19126 (N_19126,N_18757,N_18749);
xor U19127 (N_19127,N_18711,N_18612);
nor U19128 (N_19128,N_18685,N_18846);
nand U19129 (N_19129,N_18857,N_18751);
nor U19130 (N_19130,N_18742,N_18711);
nor U19131 (N_19131,N_18867,N_18666);
nand U19132 (N_19132,N_18896,N_18690);
and U19133 (N_19133,N_18786,N_18711);
or U19134 (N_19134,N_18799,N_18865);
nor U19135 (N_19135,N_18838,N_18871);
xnor U19136 (N_19136,N_18668,N_18735);
or U19137 (N_19137,N_18770,N_18817);
and U19138 (N_19138,N_18811,N_18890);
xor U19139 (N_19139,N_18657,N_18737);
nor U19140 (N_19140,N_18801,N_18695);
and U19141 (N_19141,N_18656,N_18846);
and U19142 (N_19142,N_18706,N_18624);
and U19143 (N_19143,N_18740,N_18700);
nor U19144 (N_19144,N_18807,N_18881);
and U19145 (N_19145,N_18664,N_18707);
and U19146 (N_19146,N_18813,N_18682);
nor U19147 (N_19147,N_18647,N_18719);
or U19148 (N_19148,N_18702,N_18609);
or U19149 (N_19149,N_18739,N_18755);
xor U19150 (N_19150,N_18663,N_18716);
or U19151 (N_19151,N_18691,N_18658);
or U19152 (N_19152,N_18744,N_18814);
xor U19153 (N_19153,N_18732,N_18764);
nor U19154 (N_19154,N_18661,N_18796);
nor U19155 (N_19155,N_18838,N_18858);
or U19156 (N_19156,N_18731,N_18624);
nor U19157 (N_19157,N_18733,N_18787);
xnor U19158 (N_19158,N_18787,N_18838);
xor U19159 (N_19159,N_18872,N_18617);
nor U19160 (N_19160,N_18773,N_18613);
or U19161 (N_19161,N_18798,N_18888);
nor U19162 (N_19162,N_18828,N_18824);
and U19163 (N_19163,N_18893,N_18707);
and U19164 (N_19164,N_18809,N_18886);
and U19165 (N_19165,N_18827,N_18865);
xor U19166 (N_19166,N_18845,N_18657);
or U19167 (N_19167,N_18793,N_18740);
nor U19168 (N_19168,N_18658,N_18690);
or U19169 (N_19169,N_18751,N_18713);
nor U19170 (N_19170,N_18709,N_18623);
and U19171 (N_19171,N_18668,N_18817);
nand U19172 (N_19172,N_18866,N_18751);
xnor U19173 (N_19173,N_18835,N_18651);
nand U19174 (N_19174,N_18728,N_18659);
and U19175 (N_19175,N_18650,N_18811);
nand U19176 (N_19176,N_18648,N_18659);
xnor U19177 (N_19177,N_18895,N_18793);
nor U19178 (N_19178,N_18690,N_18726);
nor U19179 (N_19179,N_18738,N_18890);
and U19180 (N_19180,N_18730,N_18867);
xor U19181 (N_19181,N_18800,N_18756);
nand U19182 (N_19182,N_18813,N_18696);
and U19183 (N_19183,N_18873,N_18653);
or U19184 (N_19184,N_18756,N_18788);
or U19185 (N_19185,N_18642,N_18662);
xnor U19186 (N_19186,N_18792,N_18823);
nand U19187 (N_19187,N_18756,N_18833);
or U19188 (N_19188,N_18876,N_18702);
xor U19189 (N_19189,N_18841,N_18752);
or U19190 (N_19190,N_18890,N_18603);
nand U19191 (N_19191,N_18867,N_18601);
xnor U19192 (N_19192,N_18602,N_18747);
nor U19193 (N_19193,N_18646,N_18739);
nand U19194 (N_19194,N_18722,N_18683);
and U19195 (N_19195,N_18653,N_18879);
nor U19196 (N_19196,N_18887,N_18664);
and U19197 (N_19197,N_18746,N_18764);
xor U19198 (N_19198,N_18736,N_18691);
nor U19199 (N_19199,N_18710,N_18732);
and U19200 (N_19200,N_18996,N_19013);
or U19201 (N_19201,N_18974,N_19009);
nand U19202 (N_19202,N_19158,N_18904);
or U19203 (N_19203,N_19105,N_19197);
nand U19204 (N_19204,N_19154,N_19094);
nor U19205 (N_19205,N_18972,N_18931);
nand U19206 (N_19206,N_19079,N_19004);
nor U19207 (N_19207,N_19115,N_19199);
xor U19208 (N_19208,N_19135,N_19058);
xnor U19209 (N_19209,N_19119,N_18963);
or U19210 (N_19210,N_19090,N_18993);
and U19211 (N_19211,N_19137,N_18955);
or U19212 (N_19212,N_18915,N_19003);
nand U19213 (N_19213,N_19084,N_19081);
xor U19214 (N_19214,N_18927,N_19122);
or U19215 (N_19215,N_18939,N_18909);
nor U19216 (N_19216,N_18934,N_19172);
or U19217 (N_19217,N_19114,N_19026);
xnor U19218 (N_19218,N_19175,N_19053);
nor U19219 (N_19219,N_18924,N_18917);
nor U19220 (N_19220,N_19107,N_19121);
or U19221 (N_19221,N_19189,N_19022);
nor U19222 (N_19222,N_19169,N_19118);
nand U19223 (N_19223,N_19012,N_19076);
or U19224 (N_19224,N_19016,N_18947);
xnor U19225 (N_19225,N_19092,N_19178);
nor U19226 (N_19226,N_19007,N_18985);
and U19227 (N_19227,N_19136,N_18964);
nand U19228 (N_19228,N_19101,N_19164);
nand U19229 (N_19229,N_19177,N_18932);
xor U19230 (N_19230,N_19069,N_19075);
or U19231 (N_19231,N_19098,N_19071);
or U19232 (N_19232,N_18905,N_18921);
nor U19233 (N_19233,N_19063,N_19100);
nand U19234 (N_19234,N_18942,N_19174);
and U19235 (N_19235,N_19171,N_19049);
xor U19236 (N_19236,N_19152,N_19088);
nand U19237 (N_19237,N_19157,N_19041);
nand U19238 (N_19238,N_19198,N_18918);
and U19239 (N_19239,N_19073,N_18945);
nor U19240 (N_19240,N_19196,N_19042);
xor U19241 (N_19241,N_19035,N_18978);
nand U19242 (N_19242,N_19110,N_19173);
nand U19243 (N_19243,N_18913,N_19129);
nor U19244 (N_19244,N_18975,N_19179);
and U19245 (N_19245,N_19176,N_19166);
or U19246 (N_19246,N_18980,N_19162);
or U19247 (N_19247,N_19056,N_19047);
xor U19248 (N_19248,N_18928,N_18948);
xnor U19249 (N_19249,N_19143,N_19032);
nand U19250 (N_19250,N_19052,N_19034);
nor U19251 (N_19251,N_19167,N_18973);
and U19252 (N_19252,N_19062,N_19077);
xor U19253 (N_19253,N_19148,N_19153);
nand U19254 (N_19254,N_19165,N_19161);
or U19255 (N_19255,N_19147,N_19018);
or U19256 (N_19256,N_19020,N_18914);
and U19257 (N_19257,N_19168,N_19044);
and U19258 (N_19258,N_19111,N_19061);
xnor U19259 (N_19259,N_19030,N_19127);
nor U19260 (N_19260,N_18991,N_19039);
or U19261 (N_19261,N_19060,N_18984);
xnor U19262 (N_19262,N_18912,N_18946);
nand U19263 (N_19263,N_18935,N_18990);
or U19264 (N_19264,N_18979,N_18910);
xor U19265 (N_19265,N_19057,N_19093);
nor U19266 (N_19266,N_18994,N_18937);
or U19267 (N_19267,N_19108,N_19000);
nand U19268 (N_19268,N_18919,N_18992);
nand U19269 (N_19269,N_18951,N_18981);
xnor U19270 (N_19270,N_19195,N_19065);
nor U19271 (N_19271,N_18950,N_19170);
and U19272 (N_19272,N_18911,N_18998);
nand U19273 (N_19273,N_19085,N_18965);
or U19274 (N_19274,N_18976,N_18933);
and U19275 (N_19275,N_18941,N_19190);
or U19276 (N_19276,N_19043,N_18968);
and U19277 (N_19277,N_19054,N_19078);
or U19278 (N_19278,N_18900,N_18938);
nor U19279 (N_19279,N_18962,N_18906);
or U19280 (N_19280,N_19028,N_19074);
nor U19281 (N_19281,N_19117,N_19017);
and U19282 (N_19282,N_18957,N_18920);
nor U19283 (N_19283,N_19124,N_18925);
nand U19284 (N_19284,N_18995,N_18908);
nor U19285 (N_19285,N_18944,N_19045);
and U19286 (N_19286,N_19040,N_19021);
nor U19287 (N_19287,N_19091,N_18940);
or U19288 (N_19288,N_19019,N_19095);
or U19289 (N_19289,N_19038,N_19145);
or U19290 (N_19290,N_19008,N_19097);
xnor U19291 (N_19291,N_19001,N_19087);
nand U19292 (N_19292,N_19006,N_18999);
or U19293 (N_19293,N_18977,N_18986);
nand U19294 (N_19294,N_18988,N_19024);
nor U19295 (N_19295,N_19144,N_19086);
nor U19296 (N_19296,N_19066,N_19031);
nand U19297 (N_19297,N_18958,N_19113);
and U19298 (N_19298,N_19025,N_19180);
or U19299 (N_19299,N_18956,N_19141);
xor U19300 (N_19300,N_19184,N_18970);
nor U19301 (N_19301,N_18961,N_19067);
nand U19302 (N_19302,N_19186,N_18907);
nor U19303 (N_19303,N_19033,N_18952);
nor U19304 (N_19304,N_19181,N_19096);
or U19305 (N_19305,N_19126,N_18971);
nor U19306 (N_19306,N_18923,N_19104);
or U19307 (N_19307,N_19192,N_18901);
nand U19308 (N_19308,N_18903,N_19134);
and U19309 (N_19309,N_18966,N_18916);
xnor U19310 (N_19310,N_19183,N_19156);
or U19311 (N_19311,N_18953,N_19083);
or U19312 (N_19312,N_18960,N_19131);
xnor U19313 (N_19313,N_18929,N_19150);
or U19314 (N_19314,N_18902,N_19015);
nor U19315 (N_19315,N_19023,N_19149);
nand U19316 (N_19316,N_19029,N_19146);
nor U19317 (N_19317,N_19103,N_19070);
xor U19318 (N_19318,N_19046,N_19125);
or U19319 (N_19319,N_19102,N_19193);
or U19320 (N_19320,N_19050,N_18983);
xor U19321 (N_19321,N_18936,N_19099);
nand U19322 (N_19322,N_19182,N_19011);
or U19323 (N_19323,N_19051,N_19187);
nor U19324 (N_19324,N_19002,N_18926);
and U19325 (N_19325,N_18982,N_19128);
nor U19326 (N_19326,N_19132,N_19142);
or U19327 (N_19327,N_19109,N_18997);
or U19328 (N_19328,N_19139,N_18922);
xor U19329 (N_19329,N_19036,N_19010);
nand U19330 (N_19330,N_19188,N_19112);
nor U19331 (N_19331,N_19116,N_19106);
or U19332 (N_19332,N_19120,N_19185);
and U19333 (N_19333,N_19082,N_18949);
xor U19334 (N_19334,N_18954,N_19089);
xor U19335 (N_19335,N_19163,N_19138);
nor U19336 (N_19336,N_19080,N_19140);
xnor U19337 (N_19337,N_18987,N_19151);
and U19338 (N_19338,N_19123,N_19160);
and U19339 (N_19339,N_18930,N_18969);
nor U19340 (N_19340,N_19048,N_19159);
nor U19341 (N_19341,N_18959,N_19059);
nand U19342 (N_19342,N_19064,N_18989);
xor U19343 (N_19343,N_19072,N_19005);
and U19344 (N_19344,N_19194,N_19055);
nand U19345 (N_19345,N_19014,N_19130);
nor U19346 (N_19346,N_19037,N_18967);
and U19347 (N_19347,N_19133,N_19191);
xnor U19348 (N_19348,N_18943,N_19155);
xnor U19349 (N_19349,N_19068,N_19027);
nand U19350 (N_19350,N_18943,N_19034);
xor U19351 (N_19351,N_18949,N_19103);
xor U19352 (N_19352,N_19104,N_19176);
nand U19353 (N_19353,N_18928,N_18949);
xnor U19354 (N_19354,N_19028,N_18900);
nand U19355 (N_19355,N_19085,N_19100);
or U19356 (N_19356,N_19195,N_19087);
and U19357 (N_19357,N_19004,N_19111);
nand U19358 (N_19358,N_18934,N_18946);
or U19359 (N_19359,N_18933,N_18992);
or U19360 (N_19360,N_19159,N_19019);
xor U19361 (N_19361,N_18939,N_19153);
and U19362 (N_19362,N_18927,N_19170);
or U19363 (N_19363,N_18904,N_19109);
or U19364 (N_19364,N_18928,N_18983);
xor U19365 (N_19365,N_18926,N_19165);
nor U19366 (N_19366,N_19063,N_19117);
and U19367 (N_19367,N_19182,N_18944);
or U19368 (N_19368,N_19055,N_19124);
or U19369 (N_19369,N_19123,N_19040);
or U19370 (N_19370,N_19029,N_19023);
or U19371 (N_19371,N_19098,N_19091);
xnor U19372 (N_19372,N_19125,N_18943);
xnor U19373 (N_19373,N_19154,N_19156);
nand U19374 (N_19374,N_19007,N_19036);
nand U19375 (N_19375,N_19083,N_19029);
or U19376 (N_19376,N_18954,N_19165);
xnor U19377 (N_19377,N_19133,N_19088);
and U19378 (N_19378,N_18936,N_19037);
xor U19379 (N_19379,N_19110,N_18907);
or U19380 (N_19380,N_18999,N_19083);
nor U19381 (N_19381,N_18975,N_19158);
nand U19382 (N_19382,N_18999,N_19197);
or U19383 (N_19383,N_18923,N_19145);
and U19384 (N_19384,N_19052,N_18945);
xor U19385 (N_19385,N_19172,N_18984);
nor U19386 (N_19386,N_18981,N_19184);
nand U19387 (N_19387,N_19170,N_19052);
nor U19388 (N_19388,N_19169,N_18979);
xor U19389 (N_19389,N_19111,N_19169);
xor U19390 (N_19390,N_19002,N_19157);
and U19391 (N_19391,N_19189,N_18950);
nand U19392 (N_19392,N_19121,N_19126);
nor U19393 (N_19393,N_19019,N_19122);
xnor U19394 (N_19394,N_19154,N_19031);
nand U19395 (N_19395,N_19178,N_18964);
nand U19396 (N_19396,N_19150,N_19149);
nor U19397 (N_19397,N_19043,N_19108);
or U19398 (N_19398,N_19146,N_19108);
or U19399 (N_19399,N_19146,N_19042);
nor U19400 (N_19400,N_18990,N_19004);
nor U19401 (N_19401,N_18973,N_19127);
nor U19402 (N_19402,N_18931,N_19138);
xor U19403 (N_19403,N_18947,N_18962);
and U19404 (N_19404,N_19139,N_18982);
nand U19405 (N_19405,N_19157,N_18955);
and U19406 (N_19406,N_19030,N_18938);
and U19407 (N_19407,N_18931,N_18967);
and U19408 (N_19408,N_19019,N_18925);
and U19409 (N_19409,N_18905,N_19149);
xnor U19410 (N_19410,N_19087,N_18942);
and U19411 (N_19411,N_19081,N_18931);
nor U19412 (N_19412,N_19128,N_18952);
nor U19413 (N_19413,N_19152,N_18941);
nor U19414 (N_19414,N_19017,N_19135);
nand U19415 (N_19415,N_18936,N_19074);
nor U19416 (N_19416,N_18950,N_19151);
nand U19417 (N_19417,N_19026,N_19080);
and U19418 (N_19418,N_19120,N_19172);
or U19419 (N_19419,N_19099,N_19008);
nor U19420 (N_19420,N_18971,N_18948);
xnor U19421 (N_19421,N_18917,N_18914);
xor U19422 (N_19422,N_19135,N_18962);
nor U19423 (N_19423,N_19033,N_19170);
nor U19424 (N_19424,N_18996,N_19189);
nand U19425 (N_19425,N_18948,N_19053);
or U19426 (N_19426,N_18903,N_19034);
or U19427 (N_19427,N_19138,N_18912);
nor U19428 (N_19428,N_18983,N_19120);
nand U19429 (N_19429,N_19003,N_19030);
or U19430 (N_19430,N_19100,N_18900);
xnor U19431 (N_19431,N_18941,N_18953);
xnor U19432 (N_19432,N_19099,N_18951);
nand U19433 (N_19433,N_19112,N_19008);
or U19434 (N_19434,N_19031,N_19015);
xor U19435 (N_19435,N_18925,N_18944);
nor U19436 (N_19436,N_19162,N_18999);
nand U19437 (N_19437,N_19095,N_18929);
nand U19438 (N_19438,N_18996,N_19094);
nor U19439 (N_19439,N_19172,N_18901);
and U19440 (N_19440,N_18924,N_18955);
and U19441 (N_19441,N_19119,N_18956);
nand U19442 (N_19442,N_19121,N_19055);
nand U19443 (N_19443,N_19007,N_19097);
or U19444 (N_19444,N_19125,N_18909);
nor U19445 (N_19445,N_19188,N_19144);
xnor U19446 (N_19446,N_19026,N_19168);
xnor U19447 (N_19447,N_19097,N_19069);
nand U19448 (N_19448,N_19146,N_19078);
nand U19449 (N_19449,N_19106,N_19053);
or U19450 (N_19450,N_19197,N_18967);
and U19451 (N_19451,N_18912,N_19026);
nor U19452 (N_19452,N_19185,N_19066);
and U19453 (N_19453,N_18947,N_18936);
nand U19454 (N_19454,N_18932,N_19085);
xnor U19455 (N_19455,N_19008,N_18955);
and U19456 (N_19456,N_19144,N_18948);
nor U19457 (N_19457,N_19122,N_19095);
nor U19458 (N_19458,N_19044,N_19008);
and U19459 (N_19459,N_18937,N_18914);
xnor U19460 (N_19460,N_19095,N_18923);
nand U19461 (N_19461,N_19045,N_19028);
or U19462 (N_19462,N_19068,N_18919);
xor U19463 (N_19463,N_19135,N_19134);
nor U19464 (N_19464,N_19066,N_19036);
and U19465 (N_19465,N_19145,N_18962);
nand U19466 (N_19466,N_19083,N_18964);
nor U19467 (N_19467,N_18977,N_18968);
nor U19468 (N_19468,N_19023,N_18984);
and U19469 (N_19469,N_18969,N_18951);
nor U19470 (N_19470,N_19107,N_19073);
or U19471 (N_19471,N_18900,N_18989);
nor U19472 (N_19472,N_19189,N_19185);
nor U19473 (N_19473,N_19061,N_18986);
nand U19474 (N_19474,N_19116,N_19110);
or U19475 (N_19475,N_19094,N_19056);
and U19476 (N_19476,N_19175,N_19156);
xnor U19477 (N_19477,N_19097,N_19156);
nor U19478 (N_19478,N_18978,N_19136);
nor U19479 (N_19479,N_19033,N_19021);
and U19480 (N_19480,N_18910,N_19192);
nor U19481 (N_19481,N_19126,N_19151);
or U19482 (N_19482,N_18932,N_19170);
xor U19483 (N_19483,N_18956,N_18951);
and U19484 (N_19484,N_18915,N_18907);
and U19485 (N_19485,N_19050,N_19136);
nor U19486 (N_19486,N_19158,N_18977);
and U19487 (N_19487,N_18991,N_19147);
and U19488 (N_19488,N_19189,N_18926);
xnor U19489 (N_19489,N_19162,N_19031);
and U19490 (N_19490,N_19180,N_19150);
xnor U19491 (N_19491,N_19099,N_19190);
or U19492 (N_19492,N_19107,N_18902);
nand U19493 (N_19493,N_19152,N_18970);
and U19494 (N_19494,N_19013,N_18909);
nor U19495 (N_19495,N_18909,N_19197);
nand U19496 (N_19496,N_19019,N_19140);
nand U19497 (N_19497,N_19142,N_19149);
nand U19498 (N_19498,N_18962,N_18956);
or U19499 (N_19499,N_19121,N_19187);
and U19500 (N_19500,N_19296,N_19444);
or U19501 (N_19501,N_19340,N_19452);
xor U19502 (N_19502,N_19201,N_19266);
or U19503 (N_19503,N_19220,N_19247);
xor U19504 (N_19504,N_19403,N_19473);
and U19505 (N_19505,N_19227,N_19350);
and U19506 (N_19506,N_19382,N_19251);
nand U19507 (N_19507,N_19469,N_19229);
nor U19508 (N_19508,N_19427,N_19391);
xor U19509 (N_19509,N_19388,N_19485);
xnor U19510 (N_19510,N_19438,N_19453);
nor U19511 (N_19511,N_19298,N_19205);
nor U19512 (N_19512,N_19499,N_19317);
nand U19513 (N_19513,N_19377,N_19475);
nor U19514 (N_19514,N_19404,N_19398);
and U19515 (N_19515,N_19419,N_19304);
nor U19516 (N_19516,N_19365,N_19378);
xnor U19517 (N_19517,N_19488,N_19496);
and U19518 (N_19518,N_19487,N_19372);
nor U19519 (N_19519,N_19206,N_19215);
or U19520 (N_19520,N_19231,N_19217);
nor U19521 (N_19521,N_19439,N_19308);
xor U19522 (N_19522,N_19356,N_19320);
xor U19523 (N_19523,N_19284,N_19417);
and U19524 (N_19524,N_19423,N_19346);
or U19525 (N_19525,N_19491,N_19449);
xor U19526 (N_19526,N_19384,N_19315);
nand U19527 (N_19527,N_19457,N_19337);
xor U19528 (N_19528,N_19376,N_19326);
nand U19529 (N_19529,N_19322,N_19450);
nor U19530 (N_19530,N_19361,N_19349);
nor U19531 (N_19531,N_19250,N_19425);
and U19532 (N_19532,N_19360,N_19219);
or U19533 (N_19533,N_19244,N_19275);
and U19534 (N_19534,N_19324,N_19413);
xor U19535 (N_19535,N_19328,N_19310);
xor U19536 (N_19536,N_19292,N_19258);
xnor U19537 (N_19537,N_19448,N_19218);
xor U19538 (N_19538,N_19397,N_19273);
nor U19539 (N_19539,N_19462,N_19354);
nand U19540 (N_19540,N_19478,N_19463);
xnor U19541 (N_19541,N_19392,N_19339);
xor U19542 (N_19542,N_19305,N_19238);
xor U19543 (N_19543,N_19494,N_19470);
and U19544 (N_19544,N_19431,N_19207);
or U19545 (N_19545,N_19264,N_19375);
or U19546 (N_19546,N_19233,N_19430);
nor U19547 (N_19547,N_19271,N_19293);
or U19548 (N_19548,N_19249,N_19210);
or U19549 (N_19549,N_19393,N_19368);
or U19550 (N_19550,N_19236,N_19331);
or U19551 (N_19551,N_19486,N_19465);
nor U19552 (N_19552,N_19259,N_19254);
nor U19553 (N_19553,N_19440,N_19385);
xor U19554 (N_19554,N_19325,N_19367);
nor U19555 (N_19555,N_19243,N_19480);
nor U19556 (N_19556,N_19255,N_19460);
and U19557 (N_19557,N_19260,N_19295);
and U19558 (N_19558,N_19389,N_19228);
or U19559 (N_19559,N_19287,N_19262);
and U19560 (N_19560,N_19409,N_19471);
xor U19561 (N_19561,N_19224,N_19222);
nand U19562 (N_19562,N_19467,N_19371);
or U19563 (N_19563,N_19234,N_19290);
and U19564 (N_19564,N_19373,N_19272);
xnor U19565 (N_19565,N_19357,N_19242);
nor U19566 (N_19566,N_19241,N_19351);
or U19567 (N_19567,N_19434,N_19380);
nand U19568 (N_19568,N_19202,N_19297);
or U19569 (N_19569,N_19355,N_19497);
and U19570 (N_19570,N_19447,N_19212);
and U19571 (N_19571,N_19239,N_19395);
and U19572 (N_19572,N_19407,N_19461);
and U19573 (N_19573,N_19265,N_19267);
xor U19574 (N_19574,N_19476,N_19416);
nor U19575 (N_19575,N_19223,N_19256);
and U19576 (N_19576,N_19410,N_19301);
nand U19577 (N_19577,N_19443,N_19402);
nand U19578 (N_19578,N_19268,N_19221);
and U19579 (N_19579,N_19263,N_19436);
xnor U19580 (N_19580,N_19422,N_19386);
nor U19581 (N_19581,N_19394,N_19442);
nand U19582 (N_19582,N_19232,N_19466);
and U19583 (N_19583,N_19342,N_19369);
nand U19584 (N_19584,N_19323,N_19455);
or U19585 (N_19585,N_19314,N_19278);
and U19586 (N_19586,N_19279,N_19341);
nor U19587 (N_19587,N_19399,N_19362);
nand U19588 (N_19588,N_19344,N_19329);
or U19589 (N_19589,N_19387,N_19370);
nor U19590 (N_19590,N_19490,N_19379);
nor U19591 (N_19591,N_19336,N_19225);
nand U19592 (N_19592,N_19433,N_19408);
and U19593 (N_19593,N_19319,N_19456);
and U19594 (N_19594,N_19454,N_19281);
nor U19595 (N_19595,N_19445,N_19451);
and U19596 (N_19596,N_19432,N_19214);
and U19597 (N_19597,N_19400,N_19321);
nor U19598 (N_19598,N_19401,N_19498);
nand U19599 (N_19599,N_19235,N_19489);
xnor U19600 (N_19600,N_19472,N_19333);
or U19601 (N_19601,N_19484,N_19343);
or U19602 (N_19602,N_19300,N_19311);
or U19603 (N_19603,N_19390,N_19381);
nand U19604 (N_19604,N_19240,N_19359);
xnor U19605 (N_19605,N_19213,N_19426);
and U19606 (N_19606,N_19330,N_19316);
and U19607 (N_19607,N_19338,N_19313);
and U19608 (N_19608,N_19307,N_19209);
nand U19609 (N_19609,N_19446,N_19282);
or U19610 (N_19610,N_19327,N_19257);
and U19611 (N_19611,N_19347,N_19479);
nand U19612 (N_19612,N_19274,N_19294);
nand U19613 (N_19613,N_19334,N_19441);
nor U19614 (N_19614,N_19252,N_19374);
nand U19615 (N_19615,N_19289,N_19200);
xnor U19616 (N_19616,N_19332,N_19481);
or U19617 (N_19617,N_19435,N_19358);
nor U19618 (N_19618,N_19352,N_19428);
nor U19619 (N_19619,N_19364,N_19424);
and U19620 (N_19620,N_19230,N_19303);
and U19621 (N_19621,N_19437,N_19226);
nand U19622 (N_19622,N_19283,N_19474);
or U19623 (N_19623,N_19291,N_19468);
or U19624 (N_19624,N_19406,N_19208);
nor U19625 (N_19625,N_19203,N_19204);
or U19626 (N_19626,N_19415,N_19348);
and U19627 (N_19627,N_19285,N_19414);
xor U19628 (N_19628,N_19245,N_19216);
nor U19629 (N_19629,N_19345,N_19261);
and U19630 (N_19630,N_19299,N_19269);
xor U19631 (N_19631,N_19482,N_19418);
nand U19632 (N_19632,N_19492,N_19366);
and U19633 (N_19633,N_19277,N_19411);
nor U19634 (N_19634,N_19280,N_19493);
xnor U19635 (N_19635,N_19405,N_19495);
nand U19636 (N_19636,N_19353,N_19302);
nor U19637 (N_19637,N_19318,N_19421);
nand U19638 (N_19638,N_19483,N_19306);
nand U19639 (N_19639,N_19464,N_19335);
nor U19640 (N_19640,N_19429,N_19237);
nand U19641 (N_19641,N_19288,N_19458);
or U19642 (N_19642,N_19459,N_19211);
xor U19643 (N_19643,N_19248,N_19312);
nor U19644 (N_19644,N_19420,N_19396);
nor U19645 (N_19645,N_19270,N_19309);
xor U19646 (N_19646,N_19253,N_19246);
and U19647 (N_19647,N_19276,N_19286);
nand U19648 (N_19648,N_19383,N_19363);
nor U19649 (N_19649,N_19412,N_19477);
xnor U19650 (N_19650,N_19475,N_19374);
xor U19651 (N_19651,N_19243,N_19283);
nor U19652 (N_19652,N_19382,N_19211);
nand U19653 (N_19653,N_19428,N_19453);
nand U19654 (N_19654,N_19386,N_19420);
or U19655 (N_19655,N_19211,N_19247);
or U19656 (N_19656,N_19303,N_19478);
nor U19657 (N_19657,N_19450,N_19442);
or U19658 (N_19658,N_19201,N_19254);
or U19659 (N_19659,N_19258,N_19442);
or U19660 (N_19660,N_19424,N_19339);
nand U19661 (N_19661,N_19298,N_19352);
xnor U19662 (N_19662,N_19243,N_19214);
xnor U19663 (N_19663,N_19324,N_19206);
nor U19664 (N_19664,N_19329,N_19267);
nor U19665 (N_19665,N_19271,N_19471);
and U19666 (N_19666,N_19468,N_19353);
nor U19667 (N_19667,N_19470,N_19462);
or U19668 (N_19668,N_19329,N_19237);
nor U19669 (N_19669,N_19422,N_19236);
or U19670 (N_19670,N_19379,N_19445);
nor U19671 (N_19671,N_19264,N_19400);
xnor U19672 (N_19672,N_19229,N_19344);
or U19673 (N_19673,N_19370,N_19464);
and U19674 (N_19674,N_19241,N_19341);
or U19675 (N_19675,N_19251,N_19436);
or U19676 (N_19676,N_19473,N_19283);
nor U19677 (N_19677,N_19345,N_19275);
nand U19678 (N_19678,N_19284,N_19410);
or U19679 (N_19679,N_19497,N_19261);
nand U19680 (N_19680,N_19213,N_19252);
nor U19681 (N_19681,N_19345,N_19276);
xor U19682 (N_19682,N_19498,N_19217);
nand U19683 (N_19683,N_19431,N_19225);
or U19684 (N_19684,N_19443,N_19407);
nor U19685 (N_19685,N_19337,N_19283);
or U19686 (N_19686,N_19233,N_19467);
xnor U19687 (N_19687,N_19234,N_19278);
or U19688 (N_19688,N_19200,N_19305);
nand U19689 (N_19689,N_19393,N_19212);
and U19690 (N_19690,N_19270,N_19235);
nand U19691 (N_19691,N_19348,N_19240);
nand U19692 (N_19692,N_19333,N_19427);
and U19693 (N_19693,N_19411,N_19490);
nor U19694 (N_19694,N_19346,N_19299);
xnor U19695 (N_19695,N_19432,N_19331);
and U19696 (N_19696,N_19460,N_19270);
and U19697 (N_19697,N_19206,N_19410);
nand U19698 (N_19698,N_19391,N_19251);
or U19699 (N_19699,N_19227,N_19347);
nor U19700 (N_19700,N_19494,N_19442);
nor U19701 (N_19701,N_19371,N_19374);
and U19702 (N_19702,N_19436,N_19347);
or U19703 (N_19703,N_19448,N_19309);
xor U19704 (N_19704,N_19480,N_19252);
nor U19705 (N_19705,N_19318,N_19499);
nand U19706 (N_19706,N_19393,N_19459);
and U19707 (N_19707,N_19485,N_19359);
or U19708 (N_19708,N_19275,N_19486);
nand U19709 (N_19709,N_19471,N_19469);
and U19710 (N_19710,N_19259,N_19300);
nand U19711 (N_19711,N_19338,N_19294);
or U19712 (N_19712,N_19279,N_19315);
xor U19713 (N_19713,N_19343,N_19482);
or U19714 (N_19714,N_19492,N_19456);
and U19715 (N_19715,N_19321,N_19247);
nand U19716 (N_19716,N_19269,N_19278);
and U19717 (N_19717,N_19225,N_19468);
and U19718 (N_19718,N_19444,N_19211);
and U19719 (N_19719,N_19452,N_19356);
or U19720 (N_19720,N_19290,N_19209);
or U19721 (N_19721,N_19378,N_19393);
xnor U19722 (N_19722,N_19439,N_19380);
or U19723 (N_19723,N_19462,N_19246);
nor U19724 (N_19724,N_19318,N_19416);
and U19725 (N_19725,N_19376,N_19450);
or U19726 (N_19726,N_19250,N_19474);
nand U19727 (N_19727,N_19401,N_19234);
and U19728 (N_19728,N_19242,N_19286);
nand U19729 (N_19729,N_19381,N_19313);
or U19730 (N_19730,N_19463,N_19452);
or U19731 (N_19731,N_19345,N_19212);
nand U19732 (N_19732,N_19436,N_19262);
nor U19733 (N_19733,N_19423,N_19416);
or U19734 (N_19734,N_19452,N_19374);
and U19735 (N_19735,N_19395,N_19292);
and U19736 (N_19736,N_19380,N_19378);
or U19737 (N_19737,N_19238,N_19271);
or U19738 (N_19738,N_19379,N_19314);
xnor U19739 (N_19739,N_19265,N_19364);
xnor U19740 (N_19740,N_19487,N_19396);
nand U19741 (N_19741,N_19448,N_19395);
nor U19742 (N_19742,N_19356,N_19326);
or U19743 (N_19743,N_19479,N_19381);
and U19744 (N_19744,N_19265,N_19380);
xor U19745 (N_19745,N_19439,N_19292);
xnor U19746 (N_19746,N_19261,N_19228);
nor U19747 (N_19747,N_19291,N_19470);
and U19748 (N_19748,N_19280,N_19356);
or U19749 (N_19749,N_19264,N_19213);
or U19750 (N_19750,N_19408,N_19458);
nand U19751 (N_19751,N_19257,N_19335);
xnor U19752 (N_19752,N_19321,N_19356);
and U19753 (N_19753,N_19215,N_19348);
xnor U19754 (N_19754,N_19376,N_19422);
nand U19755 (N_19755,N_19491,N_19203);
nand U19756 (N_19756,N_19499,N_19379);
and U19757 (N_19757,N_19228,N_19251);
and U19758 (N_19758,N_19420,N_19333);
or U19759 (N_19759,N_19398,N_19458);
and U19760 (N_19760,N_19474,N_19288);
and U19761 (N_19761,N_19384,N_19253);
nand U19762 (N_19762,N_19333,N_19361);
nor U19763 (N_19763,N_19268,N_19200);
and U19764 (N_19764,N_19330,N_19411);
nand U19765 (N_19765,N_19334,N_19432);
nand U19766 (N_19766,N_19311,N_19307);
nor U19767 (N_19767,N_19379,N_19423);
or U19768 (N_19768,N_19428,N_19332);
nand U19769 (N_19769,N_19266,N_19371);
xnor U19770 (N_19770,N_19374,N_19343);
or U19771 (N_19771,N_19347,N_19249);
nor U19772 (N_19772,N_19452,N_19237);
and U19773 (N_19773,N_19208,N_19335);
or U19774 (N_19774,N_19376,N_19254);
xor U19775 (N_19775,N_19331,N_19278);
nand U19776 (N_19776,N_19445,N_19310);
or U19777 (N_19777,N_19482,N_19246);
and U19778 (N_19778,N_19263,N_19409);
xor U19779 (N_19779,N_19424,N_19262);
or U19780 (N_19780,N_19458,N_19477);
nand U19781 (N_19781,N_19378,N_19443);
or U19782 (N_19782,N_19265,N_19347);
xor U19783 (N_19783,N_19479,N_19329);
nor U19784 (N_19784,N_19413,N_19276);
nor U19785 (N_19785,N_19493,N_19378);
nor U19786 (N_19786,N_19471,N_19234);
nand U19787 (N_19787,N_19275,N_19287);
nor U19788 (N_19788,N_19242,N_19354);
nor U19789 (N_19789,N_19422,N_19221);
or U19790 (N_19790,N_19348,N_19474);
nand U19791 (N_19791,N_19321,N_19351);
nand U19792 (N_19792,N_19301,N_19228);
nand U19793 (N_19793,N_19498,N_19415);
xor U19794 (N_19794,N_19227,N_19403);
nand U19795 (N_19795,N_19402,N_19463);
xor U19796 (N_19796,N_19405,N_19451);
nor U19797 (N_19797,N_19255,N_19336);
or U19798 (N_19798,N_19322,N_19261);
nor U19799 (N_19799,N_19481,N_19492);
nand U19800 (N_19800,N_19664,N_19533);
or U19801 (N_19801,N_19569,N_19797);
or U19802 (N_19802,N_19783,N_19679);
nand U19803 (N_19803,N_19763,N_19656);
or U19804 (N_19804,N_19760,N_19681);
or U19805 (N_19805,N_19554,N_19748);
or U19806 (N_19806,N_19701,N_19649);
and U19807 (N_19807,N_19615,N_19546);
nor U19808 (N_19808,N_19594,N_19511);
or U19809 (N_19809,N_19575,N_19683);
and U19810 (N_19810,N_19504,N_19631);
xnor U19811 (N_19811,N_19609,N_19704);
nand U19812 (N_19812,N_19650,N_19567);
or U19813 (N_19813,N_19582,N_19700);
nand U19814 (N_19814,N_19688,N_19677);
nand U19815 (N_19815,N_19675,N_19727);
and U19816 (N_19816,N_19785,N_19782);
xor U19817 (N_19817,N_19709,N_19661);
xor U19818 (N_19818,N_19577,N_19795);
or U19819 (N_19819,N_19672,N_19562);
nand U19820 (N_19820,N_19508,N_19728);
or U19821 (N_19821,N_19738,N_19680);
nor U19822 (N_19822,N_19604,N_19684);
xor U19823 (N_19823,N_19669,N_19520);
nand U19824 (N_19824,N_19674,N_19509);
and U19825 (N_19825,N_19524,N_19695);
nor U19826 (N_19826,N_19587,N_19799);
nor U19827 (N_19827,N_19570,N_19761);
or U19828 (N_19828,N_19741,N_19777);
xor U19829 (N_19829,N_19647,N_19692);
nand U19830 (N_19830,N_19721,N_19781);
xnor U19831 (N_19831,N_19666,N_19667);
nor U19832 (N_19832,N_19643,N_19529);
nand U19833 (N_19833,N_19564,N_19694);
nor U19834 (N_19834,N_19521,N_19746);
xor U19835 (N_19835,N_19710,N_19780);
and U19836 (N_19836,N_19718,N_19640);
and U19837 (N_19837,N_19628,N_19552);
and U19838 (N_19838,N_19734,N_19762);
nand U19839 (N_19839,N_19703,N_19623);
xor U19840 (N_19840,N_19531,N_19597);
xnor U19841 (N_19841,N_19580,N_19589);
nor U19842 (N_19842,N_19723,N_19586);
nand U19843 (N_19843,N_19660,N_19715);
or U19844 (N_19844,N_19774,N_19638);
or U19845 (N_19845,N_19523,N_19503);
nor U19846 (N_19846,N_19540,N_19561);
nand U19847 (N_19847,N_19670,N_19616);
and U19848 (N_19848,N_19553,N_19685);
nor U19849 (N_19849,N_19654,N_19798);
nand U19850 (N_19850,N_19513,N_19527);
xnor U19851 (N_19851,N_19653,N_19500);
or U19852 (N_19852,N_19550,N_19543);
xor U19853 (N_19853,N_19689,N_19784);
xnor U19854 (N_19854,N_19563,N_19574);
xnor U19855 (N_19855,N_19599,N_19505);
and U19856 (N_19856,N_19705,N_19572);
nand U19857 (N_19857,N_19779,N_19751);
and U19858 (N_19858,N_19771,N_19592);
nand U19859 (N_19859,N_19637,N_19755);
nor U19860 (N_19860,N_19636,N_19790);
or U19861 (N_19861,N_19633,N_19750);
or U19862 (N_19862,N_19698,N_19730);
or U19863 (N_19863,N_19548,N_19642);
nand U19864 (N_19864,N_19516,N_19625);
and U19865 (N_19865,N_19530,N_19506);
xor U19866 (N_19866,N_19722,N_19632);
nor U19867 (N_19867,N_19566,N_19585);
or U19868 (N_19868,N_19515,N_19644);
nand U19869 (N_19869,N_19758,N_19534);
or U19870 (N_19870,N_19613,N_19665);
nand U19871 (N_19871,N_19568,N_19612);
or U19872 (N_19872,N_19600,N_19547);
nand U19873 (N_19873,N_19769,N_19745);
nand U19874 (N_19874,N_19652,N_19560);
nor U19875 (N_19875,N_19742,N_19571);
nand U19876 (N_19876,N_19622,N_19602);
nor U19877 (N_19877,N_19711,N_19687);
xnor U19878 (N_19878,N_19682,N_19603);
or U19879 (N_19879,N_19772,N_19608);
and U19880 (N_19880,N_19645,N_19536);
or U19881 (N_19881,N_19686,N_19598);
or U19882 (N_19882,N_19526,N_19634);
and U19883 (N_19883,N_19794,N_19590);
and U19884 (N_19884,N_19696,N_19537);
nand U19885 (N_19885,N_19678,N_19658);
nand U19886 (N_19886,N_19627,N_19729);
and U19887 (N_19887,N_19588,N_19714);
nor U19888 (N_19888,N_19576,N_19764);
xnor U19889 (N_19889,N_19732,N_19535);
xnor U19890 (N_19890,N_19736,N_19557);
xor U19891 (N_19891,N_19707,N_19502);
xnor U19892 (N_19892,N_19757,N_19551);
or U19893 (N_19893,N_19791,N_19651);
and U19894 (N_19894,N_19716,N_19744);
or U19895 (N_19895,N_19659,N_19786);
and U19896 (N_19896,N_19514,N_19691);
nor U19897 (N_19897,N_19773,N_19573);
nand U19898 (N_19898,N_19641,N_19743);
nor U19899 (N_19899,N_19778,N_19578);
and U19900 (N_19900,N_19699,N_19737);
and U19901 (N_19901,N_19541,N_19630);
xor U19902 (N_19902,N_19617,N_19655);
or U19903 (N_19903,N_19671,N_19646);
and U19904 (N_19904,N_19756,N_19789);
or U19905 (N_19905,N_19614,N_19593);
nand U19906 (N_19906,N_19584,N_19512);
nor U19907 (N_19907,N_19766,N_19605);
nand U19908 (N_19908,N_19713,N_19648);
nand U19909 (N_19909,N_19538,N_19595);
xnor U19910 (N_19910,N_19559,N_19525);
xnor U19911 (N_19911,N_19510,N_19558);
xor U19912 (N_19912,N_19775,N_19793);
xnor U19913 (N_19913,N_19752,N_19624);
nor U19914 (N_19914,N_19759,N_19708);
xnor U19915 (N_19915,N_19754,N_19629);
and U19916 (N_19916,N_19740,N_19776);
and U19917 (N_19917,N_19528,N_19676);
xnor U19918 (N_19918,N_19663,N_19768);
nand U19919 (N_19919,N_19731,N_19507);
xnor U19920 (N_19920,N_19626,N_19610);
or U19921 (N_19921,N_19690,N_19747);
nor U19922 (N_19922,N_19668,N_19717);
or U19923 (N_19923,N_19770,N_19673);
or U19924 (N_19924,N_19726,N_19539);
nand U19925 (N_19925,N_19735,N_19544);
and U19926 (N_19926,N_19620,N_19635);
nand U19927 (N_19927,N_19501,N_19725);
nor U19928 (N_19928,N_19522,N_19545);
or U19929 (N_19929,N_19787,N_19796);
and U19930 (N_19930,N_19724,N_19549);
xnor U19931 (N_19931,N_19556,N_19621);
nor U19932 (N_19932,N_19618,N_19583);
nand U19933 (N_19933,N_19733,N_19767);
or U19934 (N_19934,N_19712,N_19706);
nor U19935 (N_19935,N_19720,N_19753);
or U19936 (N_19936,N_19555,N_19532);
and U19937 (N_19937,N_19657,N_19719);
and U19938 (N_19938,N_19581,N_19662);
nor U19939 (N_19939,N_19591,N_19702);
xnor U19940 (N_19940,N_19517,N_19749);
and U19941 (N_19941,N_19611,N_19606);
or U19942 (N_19942,N_19788,N_19639);
xnor U19943 (N_19943,N_19607,N_19565);
nor U19944 (N_19944,N_19601,N_19518);
xnor U19945 (N_19945,N_19619,N_19542);
xnor U19946 (N_19946,N_19693,N_19519);
nor U19947 (N_19947,N_19579,N_19697);
or U19948 (N_19948,N_19765,N_19596);
or U19949 (N_19949,N_19792,N_19739);
xnor U19950 (N_19950,N_19607,N_19633);
nand U19951 (N_19951,N_19765,N_19557);
and U19952 (N_19952,N_19750,N_19536);
nor U19953 (N_19953,N_19740,N_19676);
and U19954 (N_19954,N_19641,N_19670);
nor U19955 (N_19955,N_19766,N_19549);
xor U19956 (N_19956,N_19584,N_19641);
and U19957 (N_19957,N_19722,N_19763);
xnor U19958 (N_19958,N_19758,N_19668);
and U19959 (N_19959,N_19704,N_19555);
nand U19960 (N_19960,N_19700,N_19547);
and U19961 (N_19961,N_19532,N_19791);
nand U19962 (N_19962,N_19563,N_19699);
or U19963 (N_19963,N_19532,N_19713);
and U19964 (N_19964,N_19585,N_19755);
or U19965 (N_19965,N_19699,N_19501);
nand U19966 (N_19966,N_19781,N_19543);
and U19967 (N_19967,N_19683,N_19577);
or U19968 (N_19968,N_19700,N_19548);
nor U19969 (N_19969,N_19527,N_19785);
xnor U19970 (N_19970,N_19798,N_19701);
nand U19971 (N_19971,N_19534,N_19578);
and U19972 (N_19972,N_19794,N_19626);
nor U19973 (N_19973,N_19664,N_19703);
xor U19974 (N_19974,N_19713,N_19530);
and U19975 (N_19975,N_19614,N_19608);
xnor U19976 (N_19976,N_19591,N_19708);
nand U19977 (N_19977,N_19653,N_19519);
nand U19978 (N_19978,N_19734,N_19584);
nand U19979 (N_19979,N_19508,N_19658);
nor U19980 (N_19980,N_19524,N_19637);
xnor U19981 (N_19981,N_19705,N_19623);
nand U19982 (N_19982,N_19669,N_19742);
nor U19983 (N_19983,N_19788,N_19591);
and U19984 (N_19984,N_19667,N_19766);
xor U19985 (N_19985,N_19534,N_19675);
and U19986 (N_19986,N_19566,N_19710);
or U19987 (N_19987,N_19654,N_19663);
and U19988 (N_19988,N_19508,N_19543);
xnor U19989 (N_19989,N_19782,N_19573);
or U19990 (N_19990,N_19555,N_19605);
nand U19991 (N_19991,N_19567,N_19525);
nand U19992 (N_19992,N_19698,N_19544);
nand U19993 (N_19993,N_19563,N_19780);
xnor U19994 (N_19994,N_19735,N_19587);
or U19995 (N_19995,N_19513,N_19723);
or U19996 (N_19996,N_19609,N_19694);
nand U19997 (N_19997,N_19760,N_19535);
or U19998 (N_19998,N_19787,N_19771);
nand U19999 (N_19999,N_19743,N_19733);
xnor U20000 (N_20000,N_19713,N_19695);
or U20001 (N_20001,N_19668,N_19607);
nand U20002 (N_20002,N_19515,N_19679);
nand U20003 (N_20003,N_19713,N_19699);
or U20004 (N_20004,N_19730,N_19784);
or U20005 (N_20005,N_19526,N_19720);
xor U20006 (N_20006,N_19619,N_19734);
nand U20007 (N_20007,N_19576,N_19536);
xnor U20008 (N_20008,N_19549,N_19570);
nand U20009 (N_20009,N_19549,N_19568);
nand U20010 (N_20010,N_19751,N_19626);
xor U20011 (N_20011,N_19538,N_19722);
nor U20012 (N_20012,N_19643,N_19679);
xor U20013 (N_20013,N_19774,N_19648);
nor U20014 (N_20014,N_19632,N_19623);
and U20015 (N_20015,N_19644,N_19578);
nand U20016 (N_20016,N_19554,N_19778);
and U20017 (N_20017,N_19622,N_19547);
nand U20018 (N_20018,N_19712,N_19747);
nand U20019 (N_20019,N_19675,N_19544);
or U20020 (N_20020,N_19684,N_19783);
nor U20021 (N_20021,N_19679,N_19530);
and U20022 (N_20022,N_19709,N_19603);
nor U20023 (N_20023,N_19728,N_19780);
nand U20024 (N_20024,N_19586,N_19656);
xor U20025 (N_20025,N_19774,N_19506);
and U20026 (N_20026,N_19528,N_19566);
or U20027 (N_20027,N_19723,N_19691);
xnor U20028 (N_20028,N_19544,N_19601);
nand U20029 (N_20029,N_19729,N_19719);
xor U20030 (N_20030,N_19611,N_19564);
nand U20031 (N_20031,N_19569,N_19757);
nand U20032 (N_20032,N_19702,N_19722);
nand U20033 (N_20033,N_19747,N_19744);
nand U20034 (N_20034,N_19544,N_19534);
nor U20035 (N_20035,N_19544,N_19569);
nor U20036 (N_20036,N_19535,N_19741);
or U20037 (N_20037,N_19627,N_19645);
or U20038 (N_20038,N_19552,N_19775);
nand U20039 (N_20039,N_19694,N_19710);
xor U20040 (N_20040,N_19568,N_19504);
nand U20041 (N_20041,N_19562,N_19755);
xor U20042 (N_20042,N_19660,N_19628);
nand U20043 (N_20043,N_19679,N_19675);
xnor U20044 (N_20044,N_19586,N_19619);
xnor U20045 (N_20045,N_19666,N_19728);
xor U20046 (N_20046,N_19712,N_19505);
and U20047 (N_20047,N_19716,N_19724);
nor U20048 (N_20048,N_19699,N_19721);
nor U20049 (N_20049,N_19558,N_19746);
and U20050 (N_20050,N_19797,N_19558);
or U20051 (N_20051,N_19759,N_19715);
and U20052 (N_20052,N_19712,N_19672);
and U20053 (N_20053,N_19736,N_19664);
nor U20054 (N_20054,N_19788,N_19686);
xor U20055 (N_20055,N_19786,N_19523);
nand U20056 (N_20056,N_19684,N_19510);
or U20057 (N_20057,N_19512,N_19676);
nand U20058 (N_20058,N_19796,N_19706);
or U20059 (N_20059,N_19531,N_19555);
nand U20060 (N_20060,N_19545,N_19619);
or U20061 (N_20061,N_19726,N_19528);
and U20062 (N_20062,N_19784,N_19632);
xnor U20063 (N_20063,N_19697,N_19688);
or U20064 (N_20064,N_19534,N_19690);
or U20065 (N_20065,N_19758,N_19579);
xnor U20066 (N_20066,N_19759,N_19761);
xor U20067 (N_20067,N_19565,N_19592);
nand U20068 (N_20068,N_19562,N_19689);
nand U20069 (N_20069,N_19766,N_19708);
xor U20070 (N_20070,N_19568,N_19753);
nor U20071 (N_20071,N_19731,N_19557);
xor U20072 (N_20072,N_19586,N_19561);
or U20073 (N_20073,N_19632,N_19586);
or U20074 (N_20074,N_19628,N_19546);
nor U20075 (N_20075,N_19554,N_19702);
and U20076 (N_20076,N_19502,N_19568);
nor U20077 (N_20077,N_19546,N_19578);
nand U20078 (N_20078,N_19763,N_19786);
nand U20079 (N_20079,N_19543,N_19707);
nand U20080 (N_20080,N_19546,N_19761);
nand U20081 (N_20081,N_19636,N_19547);
xnor U20082 (N_20082,N_19627,N_19726);
or U20083 (N_20083,N_19599,N_19622);
xor U20084 (N_20084,N_19635,N_19784);
and U20085 (N_20085,N_19784,N_19569);
or U20086 (N_20086,N_19516,N_19693);
xor U20087 (N_20087,N_19549,N_19569);
nand U20088 (N_20088,N_19577,N_19798);
nand U20089 (N_20089,N_19630,N_19770);
nor U20090 (N_20090,N_19692,N_19766);
nor U20091 (N_20091,N_19724,N_19664);
nand U20092 (N_20092,N_19644,N_19650);
and U20093 (N_20093,N_19618,N_19633);
or U20094 (N_20094,N_19655,N_19711);
xnor U20095 (N_20095,N_19604,N_19747);
nor U20096 (N_20096,N_19617,N_19658);
xnor U20097 (N_20097,N_19569,N_19541);
or U20098 (N_20098,N_19658,N_19580);
or U20099 (N_20099,N_19537,N_19527);
or U20100 (N_20100,N_19917,N_19973);
and U20101 (N_20101,N_19865,N_19854);
nor U20102 (N_20102,N_19825,N_19999);
xor U20103 (N_20103,N_19855,N_19897);
nand U20104 (N_20104,N_20097,N_19988);
and U20105 (N_20105,N_19919,N_19976);
xor U20106 (N_20106,N_19926,N_19851);
xnor U20107 (N_20107,N_19890,N_19995);
nor U20108 (N_20108,N_19831,N_19885);
or U20109 (N_20109,N_19869,N_19801);
xnor U20110 (N_20110,N_19994,N_19847);
or U20111 (N_20111,N_19992,N_19998);
nor U20112 (N_20112,N_19892,N_19985);
nor U20113 (N_20113,N_19809,N_19900);
nor U20114 (N_20114,N_19958,N_19806);
xor U20115 (N_20115,N_20063,N_20086);
xnor U20116 (N_20116,N_20024,N_19981);
xnor U20117 (N_20117,N_19975,N_20070);
xor U20118 (N_20118,N_19874,N_19977);
or U20119 (N_20119,N_20098,N_19932);
or U20120 (N_20120,N_19841,N_19949);
nor U20121 (N_20121,N_20002,N_19818);
xnor U20122 (N_20122,N_19898,N_19912);
or U20123 (N_20123,N_20045,N_19907);
and U20124 (N_20124,N_19996,N_20042);
or U20125 (N_20125,N_20017,N_19884);
nor U20126 (N_20126,N_19808,N_19930);
and U20127 (N_20127,N_19853,N_20049);
or U20128 (N_20128,N_19813,N_19812);
nand U20129 (N_20129,N_20038,N_20039);
xor U20130 (N_20130,N_19840,N_20014);
xnor U20131 (N_20131,N_20074,N_19941);
nand U20132 (N_20132,N_19833,N_19993);
nor U20133 (N_20133,N_20062,N_20075);
nor U20134 (N_20134,N_19934,N_19879);
nand U20135 (N_20135,N_20099,N_20010);
or U20136 (N_20136,N_19911,N_20079);
nand U20137 (N_20137,N_19811,N_19957);
or U20138 (N_20138,N_19972,N_19942);
nor U20139 (N_20139,N_19914,N_19936);
xnor U20140 (N_20140,N_20061,N_20025);
and U20141 (N_20141,N_19979,N_19887);
or U20142 (N_20142,N_19895,N_19873);
and U20143 (N_20143,N_19815,N_20067);
nand U20144 (N_20144,N_19928,N_20084);
xor U20145 (N_20145,N_19987,N_19844);
or U20146 (N_20146,N_19944,N_19959);
or U20147 (N_20147,N_19901,N_19970);
nand U20148 (N_20148,N_19878,N_19894);
or U20149 (N_20149,N_20081,N_19962);
nor U20150 (N_20150,N_20069,N_19868);
nand U20151 (N_20151,N_20068,N_20044);
or U20152 (N_20152,N_19816,N_19923);
nor U20153 (N_20153,N_19902,N_20043);
nand U20154 (N_20154,N_19933,N_19814);
xnor U20155 (N_20155,N_20020,N_19807);
nor U20156 (N_20156,N_19938,N_20065);
xor U20157 (N_20157,N_20015,N_19839);
nand U20158 (N_20158,N_19866,N_19950);
xnor U20159 (N_20159,N_19916,N_20001);
nand U20160 (N_20160,N_20057,N_19948);
or U20161 (N_20161,N_20047,N_19955);
or U20162 (N_20162,N_19945,N_19828);
or U20163 (N_20163,N_20093,N_19827);
nor U20164 (N_20164,N_19838,N_19889);
nor U20165 (N_20165,N_19964,N_19997);
or U20166 (N_20166,N_19984,N_20013);
and U20167 (N_20167,N_20056,N_19935);
nor U20168 (N_20168,N_20051,N_19872);
nand U20169 (N_20169,N_20004,N_19804);
nor U20170 (N_20170,N_20046,N_20019);
nor U20171 (N_20171,N_20009,N_20008);
xnor U20172 (N_20172,N_19960,N_20083);
nor U20173 (N_20173,N_20090,N_20022);
and U20174 (N_20174,N_19849,N_19820);
and U20175 (N_20175,N_20023,N_19990);
or U20176 (N_20176,N_19823,N_20021);
xnor U20177 (N_20177,N_20040,N_19858);
or U20178 (N_20178,N_20050,N_19924);
and U20179 (N_20179,N_19826,N_19830);
nand U20180 (N_20180,N_20037,N_19871);
and U20181 (N_20181,N_20058,N_19822);
and U20182 (N_20182,N_19867,N_19899);
nor U20183 (N_20183,N_20030,N_20082);
xnor U20184 (N_20184,N_19842,N_20092);
and U20185 (N_20185,N_19877,N_20088);
nand U20186 (N_20186,N_19802,N_20032);
or U20187 (N_20187,N_19946,N_20089);
xnor U20188 (N_20188,N_19963,N_19870);
nor U20189 (N_20189,N_19939,N_20035);
nand U20190 (N_20190,N_20085,N_19856);
nor U20191 (N_20191,N_20076,N_19925);
or U20192 (N_20192,N_19986,N_20053);
and U20193 (N_20193,N_20054,N_19881);
xor U20194 (N_20194,N_19835,N_19846);
nand U20195 (N_20195,N_19819,N_19832);
nand U20196 (N_20196,N_19824,N_20016);
nand U20197 (N_20197,N_19857,N_19921);
nand U20198 (N_20198,N_19876,N_20003);
nand U20199 (N_20199,N_20087,N_20000);
xnor U20200 (N_20200,N_19810,N_19953);
nand U20201 (N_20201,N_19805,N_20073);
xnor U20202 (N_20202,N_19845,N_19834);
xor U20203 (N_20203,N_19880,N_20096);
nor U20204 (N_20204,N_20007,N_19891);
nor U20205 (N_20205,N_20055,N_19980);
nor U20206 (N_20206,N_20012,N_19910);
nand U20207 (N_20207,N_19956,N_19918);
and U20208 (N_20208,N_20011,N_19837);
nor U20209 (N_20209,N_19883,N_20064);
nor U20210 (N_20210,N_20034,N_19913);
nand U20211 (N_20211,N_19940,N_19836);
xor U20212 (N_20212,N_19908,N_19967);
nand U20213 (N_20213,N_20059,N_19821);
xor U20214 (N_20214,N_20027,N_20041);
nor U20215 (N_20215,N_19893,N_19947);
and U20216 (N_20216,N_19920,N_20033);
xnor U20217 (N_20217,N_20095,N_19803);
and U20218 (N_20218,N_19966,N_20094);
nand U20219 (N_20219,N_20006,N_19982);
and U20220 (N_20220,N_20036,N_19852);
or U20221 (N_20221,N_19991,N_20091);
xor U20222 (N_20222,N_19886,N_20029);
nand U20223 (N_20223,N_20071,N_19906);
nor U20224 (N_20224,N_20080,N_19909);
nand U20225 (N_20225,N_20048,N_19931);
nor U20226 (N_20226,N_19800,N_19829);
nor U20227 (N_20227,N_19843,N_19954);
or U20228 (N_20228,N_19888,N_19859);
or U20229 (N_20229,N_19864,N_20052);
xnor U20230 (N_20230,N_19951,N_19961);
and U20231 (N_20231,N_19965,N_20072);
and U20232 (N_20232,N_20026,N_19915);
or U20233 (N_20233,N_20018,N_19943);
and U20234 (N_20234,N_20077,N_19978);
or U20235 (N_20235,N_19904,N_20005);
nand U20236 (N_20236,N_20078,N_19817);
nand U20237 (N_20237,N_19862,N_19974);
or U20238 (N_20238,N_19905,N_19952);
nor U20239 (N_20239,N_19922,N_20028);
nand U20240 (N_20240,N_20066,N_19850);
or U20241 (N_20241,N_19861,N_19929);
xor U20242 (N_20242,N_19989,N_19882);
or U20243 (N_20243,N_19863,N_19903);
and U20244 (N_20244,N_20031,N_19860);
or U20245 (N_20245,N_19848,N_19875);
xnor U20246 (N_20246,N_19971,N_19896);
or U20247 (N_20247,N_19968,N_19927);
and U20248 (N_20248,N_19937,N_19969);
xor U20249 (N_20249,N_20060,N_19983);
nor U20250 (N_20250,N_19829,N_19933);
or U20251 (N_20251,N_20078,N_19804);
nand U20252 (N_20252,N_19993,N_19841);
xor U20253 (N_20253,N_20091,N_20058);
nor U20254 (N_20254,N_20010,N_19923);
xnor U20255 (N_20255,N_19952,N_19920);
nor U20256 (N_20256,N_19864,N_20083);
and U20257 (N_20257,N_20024,N_19802);
xor U20258 (N_20258,N_19870,N_19987);
and U20259 (N_20259,N_20036,N_20074);
nand U20260 (N_20260,N_19868,N_19997);
xor U20261 (N_20261,N_19859,N_19957);
nand U20262 (N_20262,N_19913,N_20046);
or U20263 (N_20263,N_19958,N_20081);
nand U20264 (N_20264,N_20090,N_19993);
and U20265 (N_20265,N_19852,N_19902);
and U20266 (N_20266,N_19898,N_19829);
xor U20267 (N_20267,N_19947,N_20031);
nor U20268 (N_20268,N_19907,N_19990);
nor U20269 (N_20269,N_20014,N_19879);
or U20270 (N_20270,N_20028,N_19903);
and U20271 (N_20271,N_20088,N_19959);
xnor U20272 (N_20272,N_19947,N_19836);
or U20273 (N_20273,N_20092,N_19927);
xor U20274 (N_20274,N_20094,N_19901);
or U20275 (N_20275,N_20095,N_20096);
nor U20276 (N_20276,N_19917,N_20004);
xor U20277 (N_20277,N_20070,N_20067);
nor U20278 (N_20278,N_19946,N_19860);
and U20279 (N_20279,N_19824,N_19839);
or U20280 (N_20280,N_19899,N_19888);
or U20281 (N_20281,N_20054,N_19973);
and U20282 (N_20282,N_20095,N_19845);
nor U20283 (N_20283,N_19972,N_20069);
and U20284 (N_20284,N_20086,N_19972);
nand U20285 (N_20285,N_19846,N_20085);
and U20286 (N_20286,N_19984,N_20018);
and U20287 (N_20287,N_19817,N_20055);
and U20288 (N_20288,N_20083,N_19827);
and U20289 (N_20289,N_19912,N_19985);
or U20290 (N_20290,N_19814,N_20012);
nand U20291 (N_20291,N_20038,N_19852);
nor U20292 (N_20292,N_19967,N_19832);
nor U20293 (N_20293,N_19995,N_19804);
and U20294 (N_20294,N_19808,N_19948);
and U20295 (N_20295,N_19852,N_19851);
nand U20296 (N_20296,N_20072,N_20001);
and U20297 (N_20297,N_20056,N_19882);
nor U20298 (N_20298,N_19846,N_19942);
xnor U20299 (N_20299,N_20047,N_20004);
xor U20300 (N_20300,N_20082,N_20025);
nor U20301 (N_20301,N_19851,N_20087);
or U20302 (N_20302,N_20085,N_19976);
xor U20303 (N_20303,N_19985,N_20059);
nand U20304 (N_20304,N_20083,N_20089);
xnor U20305 (N_20305,N_19914,N_19883);
and U20306 (N_20306,N_19826,N_19898);
and U20307 (N_20307,N_20007,N_20034);
and U20308 (N_20308,N_19966,N_19951);
or U20309 (N_20309,N_20028,N_19881);
nor U20310 (N_20310,N_19801,N_20084);
nand U20311 (N_20311,N_20041,N_19813);
xnor U20312 (N_20312,N_19871,N_20041);
and U20313 (N_20313,N_19972,N_20050);
nand U20314 (N_20314,N_20030,N_19978);
nor U20315 (N_20315,N_19948,N_19871);
and U20316 (N_20316,N_19991,N_20056);
or U20317 (N_20317,N_19942,N_19959);
xnor U20318 (N_20318,N_19911,N_19917);
or U20319 (N_20319,N_19836,N_19948);
or U20320 (N_20320,N_20049,N_19928);
nand U20321 (N_20321,N_19973,N_20003);
or U20322 (N_20322,N_20066,N_19891);
nand U20323 (N_20323,N_19944,N_20063);
nand U20324 (N_20324,N_20049,N_20071);
and U20325 (N_20325,N_20045,N_19937);
xor U20326 (N_20326,N_19876,N_20031);
and U20327 (N_20327,N_19820,N_20088);
nand U20328 (N_20328,N_19912,N_19940);
or U20329 (N_20329,N_20097,N_19992);
or U20330 (N_20330,N_19847,N_19979);
or U20331 (N_20331,N_19965,N_20022);
or U20332 (N_20332,N_19839,N_20043);
xor U20333 (N_20333,N_19837,N_19875);
xor U20334 (N_20334,N_19930,N_19946);
and U20335 (N_20335,N_19989,N_19947);
or U20336 (N_20336,N_20087,N_20055);
xor U20337 (N_20337,N_19874,N_19863);
nand U20338 (N_20338,N_20086,N_19880);
xor U20339 (N_20339,N_19859,N_19868);
and U20340 (N_20340,N_20044,N_19832);
and U20341 (N_20341,N_19824,N_20028);
nand U20342 (N_20342,N_20026,N_20050);
nor U20343 (N_20343,N_19845,N_19801);
xor U20344 (N_20344,N_19981,N_19913);
nand U20345 (N_20345,N_19955,N_20045);
or U20346 (N_20346,N_19869,N_19977);
and U20347 (N_20347,N_19865,N_20063);
xnor U20348 (N_20348,N_19978,N_20040);
or U20349 (N_20349,N_19831,N_20083);
nand U20350 (N_20350,N_20016,N_20088);
or U20351 (N_20351,N_19966,N_19964);
nand U20352 (N_20352,N_20080,N_19853);
xnor U20353 (N_20353,N_19942,N_20009);
and U20354 (N_20354,N_20067,N_19914);
or U20355 (N_20355,N_19878,N_19866);
nor U20356 (N_20356,N_19946,N_20022);
xnor U20357 (N_20357,N_19968,N_19939);
nor U20358 (N_20358,N_19953,N_20069);
nor U20359 (N_20359,N_19818,N_19811);
or U20360 (N_20360,N_20095,N_20082);
or U20361 (N_20361,N_19874,N_19813);
and U20362 (N_20362,N_19886,N_19949);
and U20363 (N_20363,N_19867,N_19984);
or U20364 (N_20364,N_20094,N_19958);
xnor U20365 (N_20365,N_20042,N_20033);
xor U20366 (N_20366,N_20007,N_19903);
and U20367 (N_20367,N_19811,N_19911);
or U20368 (N_20368,N_19803,N_19939);
and U20369 (N_20369,N_20048,N_20097);
nand U20370 (N_20370,N_19872,N_20006);
nor U20371 (N_20371,N_19923,N_20036);
or U20372 (N_20372,N_19951,N_19932);
or U20373 (N_20373,N_19950,N_20029);
and U20374 (N_20374,N_20079,N_19949);
and U20375 (N_20375,N_19869,N_19888);
xor U20376 (N_20376,N_19936,N_19821);
and U20377 (N_20377,N_19830,N_20066);
nand U20378 (N_20378,N_20036,N_20089);
and U20379 (N_20379,N_19868,N_20057);
nand U20380 (N_20380,N_20076,N_19816);
or U20381 (N_20381,N_20067,N_19948);
nand U20382 (N_20382,N_19813,N_19821);
xnor U20383 (N_20383,N_19964,N_19830);
xor U20384 (N_20384,N_19818,N_20006);
nor U20385 (N_20385,N_19827,N_19981);
nand U20386 (N_20386,N_19868,N_19938);
or U20387 (N_20387,N_20006,N_19898);
and U20388 (N_20388,N_19825,N_19934);
xnor U20389 (N_20389,N_19943,N_19911);
nor U20390 (N_20390,N_19814,N_20013);
nand U20391 (N_20391,N_19927,N_20028);
nand U20392 (N_20392,N_19869,N_19804);
nor U20393 (N_20393,N_19998,N_20018);
nand U20394 (N_20394,N_19910,N_19905);
nand U20395 (N_20395,N_19915,N_20033);
xor U20396 (N_20396,N_19808,N_20080);
nor U20397 (N_20397,N_19840,N_19807);
and U20398 (N_20398,N_19908,N_20091);
or U20399 (N_20399,N_19890,N_20080);
and U20400 (N_20400,N_20302,N_20155);
xor U20401 (N_20401,N_20392,N_20337);
xnor U20402 (N_20402,N_20169,N_20166);
and U20403 (N_20403,N_20248,N_20103);
nor U20404 (N_20404,N_20238,N_20151);
and U20405 (N_20405,N_20129,N_20213);
or U20406 (N_20406,N_20358,N_20193);
nor U20407 (N_20407,N_20265,N_20240);
or U20408 (N_20408,N_20121,N_20305);
nand U20409 (N_20409,N_20175,N_20397);
or U20410 (N_20410,N_20219,N_20139);
and U20411 (N_20411,N_20297,N_20114);
or U20412 (N_20412,N_20122,N_20320);
nand U20413 (N_20413,N_20314,N_20235);
xnor U20414 (N_20414,N_20131,N_20108);
nor U20415 (N_20415,N_20264,N_20192);
nand U20416 (N_20416,N_20229,N_20279);
nand U20417 (N_20417,N_20367,N_20321);
and U20418 (N_20418,N_20256,N_20333);
or U20419 (N_20419,N_20323,N_20211);
nand U20420 (N_20420,N_20171,N_20247);
nand U20421 (N_20421,N_20212,N_20249);
xor U20422 (N_20422,N_20126,N_20109);
or U20423 (N_20423,N_20142,N_20383);
or U20424 (N_20424,N_20174,N_20143);
nor U20425 (N_20425,N_20257,N_20361);
or U20426 (N_20426,N_20276,N_20391);
or U20427 (N_20427,N_20290,N_20325);
nand U20428 (N_20428,N_20286,N_20241);
or U20429 (N_20429,N_20348,N_20373);
or U20430 (N_20430,N_20246,N_20170);
xor U20431 (N_20431,N_20124,N_20288);
nand U20432 (N_20432,N_20224,N_20269);
nand U20433 (N_20433,N_20304,N_20387);
nor U20434 (N_20434,N_20398,N_20385);
nor U20435 (N_20435,N_20365,N_20376);
xnor U20436 (N_20436,N_20313,N_20234);
xor U20437 (N_20437,N_20394,N_20230);
and U20438 (N_20438,N_20153,N_20243);
and U20439 (N_20439,N_20217,N_20285);
or U20440 (N_20440,N_20141,N_20366);
nand U20441 (N_20441,N_20233,N_20355);
nor U20442 (N_20442,N_20226,N_20118);
nor U20443 (N_20443,N_20210,N_20360);
xnor U20444 (N_20444,N_20251,N_20364);
and U20445 (N_20445,N_20307,N_20278);
and U20446 (N_20446,N_20389,N_20135);
and U20447 (N_20447,N_20150,N_20318);
nand U20448 (N_20448,N_20316,N_20195);
nor U20449 (N_20449,N_20197,N_20329);
nand U20450 (N_20450,N_20395,N_20223);
nand U20451 (N_20451,N_20301,N_20106);
or U20452 (N_20452,N_20375,N_20322);
nand U20453 (N_20453,N_20270,N_20262);
and U20454 (N_20454,N_20294,N_20134);
xnor U20455 (N_20455,N_20271,N_20228);
nand U20456 (N_20456,N_20245,N_20130);
and U20457 (N_20457,N_20184,N_20298);
xnor U20458 (N_20458,N_20146,N_20253);
nand U20459 (N_20459,N_20277,N_20119);
and U20460 (N_20460,N_20393,N_20208);
or U20461 (N_20461,N_20396,N_20180);
xnor U20462 (N_20462,N_20202,N_20371);
nor U20463 (N_20463,N_20273,N_20368);
nor U20464 (N_20464,N_20352,N_20237);
nand U20465 (N_20465,N_20149,N_20254);
xnor U20466 (N_20466,N_20312,N_20147);
nor U20467 (N_20467,N_20133,N_20207);
xor U20468 (N_20468,N_20140,N_20105);
and U20469 (N_20469,N_20284,N_20287);
xnor U20470 (N_20470,N_20145,N_20158);
xor U20471 (N_20471,N_20381,N_20116);
nor U20472 (N_20472,N_20292,N_20120);
or U20473 (N_20473,N_20282,N_20199);
nor U20474 (N_20474,N_20369,N_20216);
nand U20475 (N_20475,N_20188,N_20344);
and U20476 (N_20476,N_20160,N_20183);
xor U20477 (N_20477,N_20177,N_20300);
nor U20478 (N_20478,N_20345,N_20379);
and U20479 (N_20479,N_20165,N_20252);
or U20480 (N_20480,N_20363,N_20125);
nand U20481 (N_20481,N_20346,N_20161);
and U20482 (N_20482,N_20283,N_20341);
or U20483 (N_20483,N_20236,N_20162);
or U20484 (N_20484,N_20201,N_20359);
or U20485 (N_20485,N_20222,N_20220);
and U20486 (N_20486,N_20187,N_20176);
and U20487 (N_20487,N_20315,N_20261);
or U20488 (N_20488,N_20388,N_20168);
and U20489 (N_20489,N_20186,N_20113);
nand U20490 (N_20490,N_20221,N_20340);
nor U20491 (N_20491,N_20343,N_20382);
nand U20492 (N_20492,N_20159,N_20112);
or U20493 (N_20493,N_20268,N_20123);
nor U20494 (N_20494,N_20136,N_20384);
nor U20495 (N_20495,N_20328,N_20347);
nor U20496 (N_20496,N_20214,N_20196);
nor U20497 (N_20497,N_20100,N_20231);
or U20498 (N_20498,N_20308,N_20293);
nor U20499 (N_20499,N_20157,N_20306);
nor U20500 (N_20500,N_20203,N_20370);
and U20501 (N_20501,N_20357,N_20335);
or U20502 (N_20502,N_20339,N_20319);
xnor U20503 (N_20503,N_20110,N_20331);
xnor U20504 (N_20504,N_20326,N_20349);
or U20505 (N_20505,N_20336,N_20167);
and U20506 (N_20506,N_20353,N_20239);
nor U20507 (N_20507,N_20372,N_20148);
xor U20508 (N_20508,N_20362,N_20152);
nor U20509 (N_20509,N_20275,N_20266);
nor U20510 (N_20510,N_20334,N_20350);
xnor U20511 (N_20511,N_20225,N_20356);
nor U20512 (N_20512,N_20327,N_20104);
and U20513 (N_20513,N_20204,N_20399);
and U20514 (N_20514,N_20242,N_20227);
xnor U20515 (N_20515,N_20190,N_20332);
or U20516 (N_20516,N_20138,N_20132);
and U20517 (N_20517,N_20128,N_20181);
xor U20518 (N_20518,N_20107,N_20115);
nor U20519 (N_20519,N_20232,N_20172);
nor U20520 (N_20520,N_20218,N_20380);
xnor U20521 (N_20521,N_20274,N_20291);
nor U20522 (N_20522,N_20378,N_20374);
nor U20523 (N_20523,N_20198,N_20296);
nor U20524 (N_20524,N_20127,N_20189);
nand U20525 (N_20525,N_20154,N_20215);
nor U20526 (N_20526,N_20137,N_20200);
and U20527 (N_20527,N_20280,N_20295);
and U20528 (N_20528,N_20342,N_20102);
or U20529 (N_20529,N_20338,N_20259);
nand U20530 (N_20530,N_20281,N_20179);
or U20531 (N_20531,N_20311,N_20244);
or U20532 (N_20532,N_20191,N_20205);
or U20533 (N_20533,N_20101,N_20309);
or U20534 (N_20534,N_20303,N_20255);
nand U20535 (N_20535,N_20354,N_20209);
nand U20536 (N_20536,N_20164,N_20178);
nor U20537 (N_20537,N_20111,N_20377);
xor U20538 (N_20538,N_20258,N_20182);
nor U20539 (N_20539,N_20390,N_20260);
xnor U20540 (N_20540,N_20144,N_20156);
nor U20541 (N_20541,N_20163,N_20173);
nand U20542 (N_20542,N_20310,N_20185);
or U20543 (N_20543,N_20330,N_20299);
nor U20544 (N_20544,N_20272,N_20263);
nor U20545 (N_20545,N_20351,N_20206);
or U20546 (N_20546,N_20386,N_20317);
or U20547 (N_20547,N_20324,N_20289);
or U20548 (N_20548,N_20194,N_20117);
nor U20549 (N_20549,N_20267,N_20250);
nand U20550 (N_20550,N_20204,N_20172);
or U20551 (N_20551,N_20152,N_20354);
xnor U20552 (N_20552,N_20205,N_20321);
or U20553 (N_20553,N_20273,N_20180);
xnor U20554 (N_20554,N_20214,N_20243);
nor U20555 (N_20555,N_20236,N_20129);
nand U20556 (N_20556,N_20263,N_20318);
nand U20557 (N_20557,N_20365,N_20128);
xor U20558 (N_20558,N_20151,N_20140);
and U20559 (N_20559,N_20339,N_20221);
and U20560 (N_20560,N_20116,N_20152);
or U20561 (N_20561,N_20336,N_20241);
or U20562 (N_20562,N_20164,N_20149);
xor U20563 (N_20563,N_20253,N_20124);
or U20564 (N_20564,N_20219,N_20247);
or U20565 (N_20565,N_20335,N_20339);
nor U20566 (N_20566,N_20229,N_20124);
or U20567 (N_20567,N_20330,N_20226);
and U20568 (N_20568,N_20158,N_20204);
nand U20569 (N_20569,N_20188,N_20371);
nor U20570 (N_20570,N_20281,N_20216);
nand U20571 (N_20571,N_20149,N_20219);
nand U20572 (N_20572,N_20153,N_20151);
or U20573 (N_20573,N_20351,N_20190);
or U20574 (N_20574,N_20127,N_20232);
nor U20575 (N_20575,N_20112,N_20278);
and U20576 (N_20576,N_20376,N_20272);
nor U20577 (N_20577,N_20336,N_20204);
or U20578 (N_20578,N_20136,N_20377);
xor U20579 (N_20579,N_20223,N_20384);
nand U20580 (N_20580,N_20262,N_20310);
or U20581 (N_20581,N_20310,N_20369);
xor U20582 (N_20582,N_20385,N_20145);
nor U20583 (N_20583,N_20341,N_20329);
nand U20584 (N_20584,N_20182,N_20165);
nand U20585 (N_20585,N_20272,N_20235);
and U20586 (N_20586,N_20319,N_20321);
nand U20587 (N_20587,N_20232,N_20168);
xor U20588 (N_20588,N_20151,N_20321);
or U20589 (N_20589,N_20154,N_20279);
and U20590 (N_20590,N_20169,N_20304);
nor U20591 (N_20591,N_20340,N_20252);
and U20592 (N_20592,N_20281,N_20211);
or U20593 (N_20593,N_20297,N_20140);
nand U20594 (N_20594,N_20257,N_20177);
xor U20595 (N_20595,N_20384,N_20168);
nor U20596 (N_20596,N_20130,N_20353);
and U20597 (N_20597,N_20195,N_20331);
xnor U20598 (N_20598,N_20257,N_20323);
nor U20599 (N_20599,N_20143,N_20141);
and U20600 (N_20600,N_20169,N_20222);
nor U20601 (N_20601,N_20106,N_20343);
or U20602 (N_20602,N_20342,N_20387);
nor U20603 (N_20603,N_20342,N_20174);
or U20604 (N_20604,N_20289,N_20210);
xnor U20605 (N_20605,N_20240,N_20335);
nor U20606 (N_20606,N_20356,N_20121);
nand U20607 (N_20607,N_20389,N_20230);
xnor U20608 (N_20608,N_20183,N_20133);
xor U20609 (N_20609,N_20269,N_20196);
or U20610 (N_20610,N_20263,N_20350);
xnor U20611 (N_20611,N_20231,N_20244);
nand U20612 (N_20612,N_20147,N_20371);
or U20613 (N_20613,N_20196,N_20105);
xnor U20614 (N_20614,N_20174,N_20234);
nand U20615 (N_20615,N_20357,N_20393);
or U20616 (N_20616,N_20224,N_20225);
or U20617 (N_20617,N_20208,N_20308);
or U20618 (N_20618,N_20326,N_20316);
xor U20619 (N_20619,N_20380,N_20148);
nor U20620 (N_20620,N_20320,N_20310);
and U20621 (N_20621,N_20263,N_20161);
xor U20622 (N_20622,N_20328,N_20298);
nor U20623 (N_20623,N_20361,N_20307);
and U20624 (N_20624,N_20378,N_20161);
xor U20625 (N_20625,N_20398,N_20332);
or U20626 (N_20626,N_20175,N_20244);
nor U20627 (N_20627,N_20215,N_20396);
and U20628 (N_20628,N_20258,N_20303);
xnor U20629 (N_20629,N_20301,N_20361);
or U20630 (N_20630,N_20172,N_20321);
xor U20631 (N_20631,N_20314,N_20326);
and U20632 (N_20632,N_20391,N_20177);
nand U20633 (N_20633,N_20273,N_20156);
or U20634 (N_20634,N_20289,N_20323);
nor U20635 (N_20635,N_20334,N_20237);
and U20636 (N_20636,N_20305,N_20148);
and U20637 (N_20637,N_20208,N_20226);
nor U20638 (N_20638,N_20191,N_20381);
nor U20639 (N_20639,N_20175,N_20334);
and U20640 (N_20640,N_20259,N_20285);
nor U20641 (N_20641,N_20270,N_20366);
or U20642 (N_20642,N_20119,N_20267);
and U20643 (N_20643,N_20305,N_20225);
xor U20644 (N_20644,N_20171,N_20349);
or U20645 (N_20645,N_20113,N_20303);
nand U20646 (N_20646,N_20250,N_20311);
xnor U20647 (N_20647,N_20307,N_20142);
or U20648 (N_20648,N_20332,N_20215);
nor U20649 (N_20649,N_20354,N_20257);
or U20650 (N_20650,N_20342,N_20339);
nor U20651 (N_20651,N_20152,N_20134);
or U20652 (N_20652,N_20174,N_20321);
nor U20653 (N_20653,N_20336,N_20318);
nor U20654 (N_20654,N_20339,N_20134);
or U20655 (N_20655,N_20132,N_20295);
or U20656 (N_20656,N_20323,N_20369);
nor U20657 (N_20657,N_20142,N_20232);
and U20658 (N_20658,N_20148,N_20315);
or U20659 (N_20659,N_20260,N_20315);
and U20660 (N_20660,N_20223,N_20376);
nand U20661 (N_20661,N_20243,N_20335);
xnor U20662 (N_20662,N_20101,N_20124);
and U20663 (N_20663,N_20376,N_20312);
nor U20664 (N_20664,N_20116,N_20303);
nor U20665 (N_20665,N_20287,N_20301);
xor U20666 (N_20666,N_20238,N_20216);
nand U20667 (N_20667,N_20168,N_20344);
or U20668 (N_20668,N_20139,N_20257);
and U20669 (N_20669,N_20272,N_20305);
xor U20670 (N_20670,N_20246,N_20334);
nor U20671 (N_20671,N_20210,N_20205);
nand U20672 (N_20672,N_20303,N_20190);
xnor U20673 (N_20673,N_20170,N_20147);
or U20674 (N_20674,N_20206,N_20137);
xnor U20675 (N_20675,N_20336,N_20206);
or U20676 (N_20676,N_20313,N_20209);
nand U20677 (N_20677,N_20166,N_20235);
xnor U20678 (N_20678,N_20135,N_20204);
nand U20679 (N_20679,N_20337,N_20313);
nor U20680 (N_20680,N_20123,N_20201);
nor U20681 (N_20681,N_20255,N_20392);
nand U20682 (N_20682,N_20113,N_20125);
nor U20683 (N_20683,N_20339,N_20273);
xnor U20684 (N_20684,N_20157,N_20235);
xnor U20685 (N_20685,N_20154,N_20177);
or U20686 (N_20686,N_20232,N_20395);
and U20687 (N_20687,N_20322,N_20145);
nand U20688 (N_20688,N_20193,N_20285);
xnor U20689 (N_20689,N_20229,N_20210);
or U20690 (N_20690,N_20193,N_20230);
xnor U20691 (N_20691,N_20278,N_20180);
xor U20692 (N_20692,N_20120,N_20155);
or U20693 (N_20693,N_20366,N_20262);
xor U20694 (N_20694,N_20274,N_20255);
or U20695 (N_20695,N_20264,N_20351);
nor U20696 (N_20696,N_20388,N_20320);
and U20697 (N_20697,N_20298,N_20215);
xor U20698 (N_20698,N_20373,N_20152);
or U20699 (N_20699,N_20358,N_20251);
and U20700 (N_20700,N_20435,N_20457);
nand U20701 (N_20701,N_20577,N_20535);
and U20702 (N_20702,N_20657,N_20611);
xnor U20703 (N_20703,N_20616,N_20588);
or U20704 (N_20704,N_20447,N_20520);
and U20705 (N_20705,N_20496,N_20424);
xor U20706 (N_20706,N_20692,N_20574);
or U20707 (N_20707,N_20487,N_20515);
or U20708 (N_20708,N_20458,N_20656);
nor U20709 (N_20709,N_20471,N_20501);
nand U20710 (N_20710,N_20680,N_20412);
or U20711 (N_20711,N_20585,N_20538);
nand U20712 (N_20712,N_20512,N_20420);
nand U20713 (N_20713,N_20419,N_20400);
nand U20714 (N_20714,N_20417,N_20662);
or U20715 (N_20715,N_20498,N_20483);
nand U20716 (N_20716,N_20600,N_20664);
and U20717 (N_20717,N_20497,N_20413);
nand U20718 (N_20718,N_20409,N_20591);
nand U20719 (N_20719,N_20423,N_20672);
or U20720 (N_20720,N_20540,N_20661);
nor U20721 (N_20721,N_20500,N_20602);
nor U20722 (N_20722,N_20517,N_20623);
xor U20723 (N_20723,N_20652,N_20605);
and U20724 (N_20724,N_20627,N_20618);
nand U20725 (N_20725,N_20418,N_20509);
xor U20726 (N_20726,N_20474,N_20674);
xnor U20727 (N_20727,N_20530,N_20405);
nand U20728 (N_20728,N_20628,N_20679);
and U20729 (N_20729,N_20556,N_20546);
and U20730 (N_20730,N_20451,N_20690);
nor U20731 (N_20731,N_20619,N_20570);
nor U20732 (N_20732,N_20699,N_20449);
nor U20733 (N_20733,N_20408,N_20508);
and U20734 (N_20734,N_20432,N_20572);
and U20735 (N_20735,N_20518,N_20595);
or U20736 (N_20736,N_20693,N_20641);
nor U20737 (N_20737,N_20650,N_20454);
and U20738 (N_20738,N_20678,N_20523);
nor U20739 (N_20739,N_20583,N_20475);
xnor U20740 (N_20740,N_20507,N_20527);
nor U20741 (N_20741,N_20511,N_20548);
nand U20742 (N_20742,N_20613,N_20609);
nor U20743 (N_20743,N_20582,N_20545);
and U20744 (N_20744,N_20436,N_20649);
and U20745 (N_20745,N_20478,N_20614);
or U20746 (N_20746,N_20644,N_20407);
and U20747 (N_20747,N_20456,N_20437);
xnor U20748 (N_20748,N_20594,N_20562);
xor U20749 (N_20749,N_20643,N_20593);
or U20750 (N_20750,N_20668,N_20505);
or U20751 (N_20751,N_20428,N_20414);
nor U20752 (N_20752,N_20544,N_20617);
xor U20753 (N_20753,N_20427,N_20606);
nand U20754 (N_20754,N_20599,N_20687);
xnor U20755 (N_20755,N_20640,N_20670);
or U20756 (N_20756,N_20622,N_20462);
nand U20757 (N_20757,N_20658,N_20421);
and U20758 (N_20758,N_20467,N_20689);
xor U20759 (N_20759,N_20485,N_20470);
nor U20760 (N_20760,N_20607,N_20586);
xnor U20761 (N_20761,N_20442,N_20502);
nand U20762 (N_20762,N_20601,N_20559);
or U20763 (N_20763,N_20560,N_20528);
nand U20764 (N_20764,N_20571,N_20655);
and U20765 (N_20765,N_20539,N_20637);
xnor U20766 (N_20766,N_20682,N_20604);
xnor U20767 (N_20767,N_20525,N_20532);
nor U20768 (N_20768,N_20506,N_20603);
or U20769 (N_20769,N_20529,N_20433);
xor U20770 (N_20770,N_20557,N_20634);
nand U20771 (N_20771,N_20510,N_20410);
nand U20772 (N_20772,N_20446,N_20491);
nand U20773 (N_20773,N_20621,N_20667);
and U20774 (N_20774,N_20479,N_20635);
nand U20775 (N_20775,N_20561,N_20473);
or U20776 (N_20776,N_20434,N_20665);
and U20777 (N_20777,N_20463,N_20533);
or U20778 (N_20778,N_20555,N_20445);
and U20779 (N_20779,N_20406,N_20653);
nor U20780 (N_20780,N_20565,N_20566);
and U20781 (N_20781,N_20587,N_20631);
or U20782 (N_20782,N_20675,N_20639);
xnor U20783 (N_20783,N_20581,N_20576);
and U20784 (N_20784,N_20489,N_20450);
and U20785 (N_20785,N_20550,N_20426);
and U20786 (N_20786,N_20660,N_20551);
xor U20787 (N_20787,N_20615,N_20549);
nor U20788 (N_20788,N_20563,N_20513);
nor U20789 (N_20789,N_20575,N_20696);
nand U20790 (N_20790,N_20677,N_20597);
xor U20791 (N_20791,N_20620,N_20633);
xnor U20792 (N_20792,N_20610,N_20466);
nand U20793 (N_20793,N_20547,N_20695);
nor U20794 (N_20794,N_20542,N_20534);
and U20795 (N_20795,N_20686,N_20484);
and U20796 (N_20796,N_20691,N_20671);
xor U20797 (N_20797,N_20480,N_20647);
or U20798 (N_20798,N_20531,N_20464);
and U20799 (N_20799,N_20698,N_20608);
and U20800 (N_20800,N_20552,N_20584);
and U20801 (N_20801,N_20654,N_20688);
or U20802 (N_20802,N_20429,N_20537);
and U20803 (N_20803,N_20573,N_20625);
nand U20804 (N_20804,N_20460,N_20469);
and U20805 (N_20805,N_20673,N_20642);
nor U20806 (N_20806,N_20543,N_20461);
nand U20807 (N_20807,N_20567,N_20536);
and U20808 (N_20808,N_20401,N_20488);
and U20809 (N_20809,N_20438,N_20638);
or U20810 (N_20810,N_20404,N_20425);
nand U20811 (N_20811,N_20481,N_20453);
and U20812 (N_20812,N_20486,N_20465);
nand U20813 (N_20813,N_20411,N_20632);
nand U20814 (N_20814,N_20503,N_20403);
nor U20815 (N_20815,N_20681,N_20430);
or U20816 (N_20816,N_20499,N_20663);
or U20817 (N_20817,N_20495,N_20504);
nand U20818 (N_20818,N_20564,N_20580);
xor U20819 (N_20819,N_20592,N_20630);
nor U20820 (N_20820,N_20589,N_20443);
or U20821 (N_20821,N_20472,N_20476);
xor U20822 (N_20822,N_20493,N_20659);
and U20823 (N_20823,N_20444,N_20514);
or U20824 (N_20824,N_20558,N_20553);
xor U20825 (N_20825,N_20648,N_20440);
nand U20826 (N_20826,N_20519,N_20624);
nor U20827 (N_20827,N_20448,N_20402);
nand U20828 (N_20828,N_20651,N_20415);
nor U20829 (N_20829,N_20526,N_20468);
nor U20830 (N_20830,N_20459,N_20439);
nor U20831 (N_20831,N_20697,N_20522);
xnor U20832 (N_20832,N_20685,N_20590);
or U20833 (N_20833,N_20521,N_20598);
nor U20834 (N_20834,N_20636,N_20524);
nand U20835 (N_20835,N_20554,N_20455);
or U20836 (N_20836,N_20645,N_20612);
nand U20837 (N_20837,N_20416,N_20669);
or U20838 (N_20838,N_20579,N_20568);
xnor U20839 (N_20839,N_20694,N_20431);
and U20840 (N_20840,N_20490,N_20541);
nor U20841 (N_20841,N_20477,N_20646);
nor U20842 (N_20842,N_20683,N_20596);
or U20843 (N_20843,N_20578,N_20452);
nor U20844 (N_20844,N_20569,N_20494);
and U20845 (N_20845,N_20441,N_20422);
and U20846 (N_20846,N_20629,N_20482);
nor U20847 (N_20847,N_20684,N_20492);
and U20848 (N_20848,N_20666,N_20626);
nand U20849 (N_20849,N_20676,N_20516);
nand U20850 (N_20850,N_20550,N_20622);
xor U20851 (N_20851,N_20606,N_20500);
nor U20852 (N_20852,N_20532,N_20542);
nor U20853 (N_20853,N_20622,N_20624);
xor U20854 (N_20854,N_20582,N_20638);
or U20855 (N_20855,N_20598,N_20426);
xor U20856 (N_20856,N_20562,N_20435);
xnor U20857 (N_20857,N_20514,N_20628);
nand U20858 (N_20858,N_20599,N_20508);
or U20859 (N_20859,N_20570,N_20659);
or U20860 (N_20860,N_20671,N_20497);
and U20861 (N_20861,N_20687,N_20492);
and U20862 (N_20862,N_20656,N_20634);
xnor U20863 (N_20863,N_20561,N_20483);
nand U20864 (N_20864,N_20587,N_20505);
xnor U20865 (N_20865,N_20647,N_20675);
xnor U20866 (N_20866,N_20405,N_20668);
nor U20867 (N_20867,N_20532,N_20674);
xnor U20868 (N_20868,N_20486,N_20699);
xnor U20869 (N_20869,N_20648,N_20669);
nand U20870 (N_20870,N_20460,N_20536);
nor U20871 (N_20871,N_20577,N_20533);
xor U20872 (N_20872,N_20549,N_20613);
nor U20873 (N_20873,N_20631,N_20422);
xnor U20874 (N_20874,N_20448,N_20456);
and U20875 (N_20875,N_20645,N_20559);
or U20876 (N_20876,N_20603,N_20595);
xor U20877 (N_20877,N_20580,N_20535);
nand U20878 (N_20878,N_20611,N_20402);
nor U20879 (N_20879,N_20601,N_20495);
or U20880 (N_20880,N_20635,N_20643);
xnor U20881 (N_20881,N_20633,N_20634);
nor U20882 (N_20882,N_20405,N_20556);
nand U20883 (N_20883,N_20582,N_20521);
nor U20884 (N_20884,N_20494,N_20556);
or U20885 (N_20885,N_20598,N_20497);
nand U20886 (N_20886,N_20403,N_20690);
or U20887 (N_20887,N_20544,N_20575);
xnor U20888 (N_20888,N_20660,N_20684);
nand U20889 (N_20889,N_20641,N_20614);
nand U20890 (N_20890,N_20599,N_20594);
and U20891 (N_20891,N_20424,N_20647);
nor U20892 (N_20892,N_20503,N_20464);
nor U20893 (N_20893,N_20573,N_20537);
or U20894 (N_20894,N_20498,N_20691);
or U20895 (N_20895,N_20585,N_20452);
or U20896 (N_20896,N_20592,N_20608);
xnor U20897 (N_20897,N_20693,N_20594);
and U20898 (N_20898,N_20467,N_20410);
nor U20899 (N_20899,N_20555,N_20466);
xnor U20900 (N_20900,N_20526,N_20527);
xor U20901 (N_20901,N_20502,N_20581);
nand U20902 (N_20902,N_20651,N_20573);
and U20903 (N_20903,N_20664,N_20598);
and U20904 (N_20904,N_20511,N_20637);
nand U20905 (N_20905,N_20543,N_20566);
or U20906 (N_20906,N_20437,N_20497);
and U20907 (N_20907,N_20586,N_20530);
or U20908 (N_20908,N_20440,N_20613);
or U20909 (N_20909,N_20698,N_20548);
and U20910 (N_20910,N_20590,N_20406);
nand U20911 (N_20911,N_20619,N_20669);
or U20912 (N_20912,N_20441,N_20448);
xor U20913 (N_20913,N_20696,N_20597);
or U20914 (N_20914,N_20690,N_20609);
xor U20915 (N_20915,N_20675,N_20561);
nor U20916 (N_20916,N_20674,N_20586);
and U20917 (N_20917,N_20450,N_20411);
nand U20918 (N_20918,N_20623,N_20659);
and U20919 (N_20919,N_20585,N_20657);
or U20920 (N_20920,N_20529,N_20495);
nor U20921 (N_20921,N_20608,N_20447);
nor U20922 (N_20922,N_20628,N_20564);
xnor U20923 (N_20923,N_20547,N_20671);
nand U20924 (N_20924,N_20601,N_20535);
and U20925 (N_20925,N_20692,N_20695);
nor U20926 (N_20926,N_20470,N_20649);
xnor U20927 (N_20927,N_20536,N_20620);
nor U20928 (N_20928,N_20496,N_20555);
or U20929 (N_20929,N_20518,N_20636);
nand U20930 (N_20930,N_20548,N_20425);
nor U20931 (N_20931,N_20527,N_20692);
and U20932 (N_20932,N_20687,N_20402);
or U20933 (N_20933,N_20688,N_20527);
or U20934 (N_20934,N_20410,N_20560);
or U20935 (N_20935,N_20625,N_20550);
nand U20936 (N_20936,N_20484,N_20409);
nand U20937 (N_20937,N_20482,N_20466);
xor U20938 (N_20938,N_20404,N_20478);
nand U20939 (N_20939,N_20500,N_20660);
nor U20940 (N_20940,N_20404,N_20561);
and U20941 (N_20941,N_20428,N_20560);
xnor U20942 (N_20942,N_20583,N_20405);
nand U20943 (N_20943,N_20433,N_20689);
and U20944 (N_20944,N_20558,N_20403);
and U20945 (N_20945,N_20468,N_20659);
nor U20946 (N_20946,N_20554,N_20411);
or U20947 (N_20947,N_20639,N_20664);
or U20948 (N_20948,N_20581,N_20635);
or U20949 (N_20949,N_20570,N_20622);
or U20950 (N_20950,N_20672,N_20674);
or U20951 (N_20951,N_20484,N_20592);
xor U20952 (N_20952,N_20582,N_20459);
nand U20953 (N_20953,N_20619,N_20461);
and U20954 (N_20954,N_20576,N_20469);
xor U20955 (N_20955,N_20428,N_20630);
and U20956 (N_20956,N_20464,N_20506);
nand U20957 (N_20957,N_20482,N_20513);
or U20958 (N_20958,N_20681,N_20686);
xnor U20959 (N_20959,N_20642,N_20569);
nor U20960 (N_20960,N_20561,N_20567);
nand U20961 (N_20961,N_20463,N_20585);
nor U20962 (N_20962,N_20453,N_20414);
nor U20963 (N_20963,N_20402,N_20679);
or U20964 (N_20964,N_20681,N_20420);
or U20965 (N_20965,N_20429,N_20554);
and U20966 (N_20966,N_20532,N_20683);
and U20967 (N_20967,N_20481,N_20486);
nand U20968 (N_20968,N_20648,N_20591);
or U20969 (N_20969,N_20500,N_20472);
nor U20970 (N_20970,N_20691,N_20454);
and U20971 (N_20971,N_20504,N_20650);
nor U20972 (N_20972,N_20564,N_20578);
nand U20973 (N_20973,N_20659,N_20697);
xor U20974 (N_20974,N_20554,N_20589);
and U20975 (N_20975,N_20445,N_20562);
nand U20976 (N_20976,N_20445,N_20631);
nor U20977 (N_20977,N_20482,N_20448);
nor U20978 (N_20978,N_20632,N_20627);
nor U20979 (N_20979,N_20655,N_20432);
nand U20980 (N_20980,N_20698,N_20659);
nand U20981 (N_20981,N_20592,N_20446);
and U20982 (N_20982,N_20576,N_20505);
nor U20983 (N_20983,N_20665,N_20698);
xor U20984 (N_20984,N_20493,N_20574);
and U20985 (N_20985,N_20679,N_20647);
and U20986 (N_20986,N_20459,N_20476);
nor U20987 (N_20987,N_20605,N_20598);
and U20988 (N_20988,N_20492,N_20498);
or U20989 (N_20989,N_20688,N_20509);
nor U20990 (N_20990,N_20671,N_20643);
and U20991 (N_20991,N_20682,N_20689);
nor U20992 (N_20992,N_20630,N_20439);
and U20993 (N_20993,N_20613,N_20466);
nand U20994 (N_20994,N_20637,N_20597);
nor U20995 (N_20995,N_20578,N_20508);
xor U20996 (N_20996,N_20441,N_20676);
nor U20997 (N_20997,N_20463,N_20428);
nor U20998 (N_20998,N_20443,N_20551);
nor U20999 (N_20999,N_20557,N_20593);
or U21000 (N_21000,N_20938,N_20910);
xnor U21001 (N_21001,N_20976,N_20706);
and U21002 (N_21002,N_20839,N_20806);
nand U21003 (N_21003,N_20876,N_20838);
and U21004 (N_21004,N_20749,N_20871);
or U21005 (N_21005,N_20966,N_20834);
xnor U21006 (N_21006,N_20993,N_20799);
nand U21007 (N_21007,N_20944,N_20802);
xnor U21008 (N_21008,N_20874,N_20848);
or U21009 (N_21009,N_20737,N_20942);
nand U21010 (N_21010,N_20721,N_20967);
nand U21011 (N_21011,N_20812,N_20969);
nor U21012 (N_21012,N_20979,N_20972);
nand U21013 (N_21013,N_20723,N_20758);
xor U21014 (N_21014,N_20958,N_20740);
nand U21015 (N_21015,N_20870,N_20890);
and U21016 (N_21016,N_20869,N_20866);
and U21017 (N_21017,N_20902,N_20922);
xor U21018 (N_21018,N_20710,N_20735);
xor U21019 (N_21019,N_20790,N_20939);
xor U21020 (N_21020,N_20864,N_20726);
nor U21021 (N_21021,N_20813,N_20985);
xor U21022 (N_21022,N_20945,N_20775);
nor U21023 (N_21023,N_20982,N_20903);
or U21024 (N_21024,N_20947,N_20745);
nand U21025 (N_21025,N_20765,N_20808);
and U21026 (N_21026,N_20893,N_20889);
nor U21027 (N_21027,N_20828,N_20840);
and U21028 (N_21028,N_20786,N_20729);
or U21029 (N_21029,N_20955,N_20803);
xnor U21030 (N_21030,N_20717,N_20776);
xor U21031 (N_21031,N_20724,N_20901);
or U21032 (N_21032,N_20843,N_20957);
or U21033 (N_21033,N_20912,N_20998);
nand U21034 (N_21034,N_20914,N_20741);
or U21035 (N_21035,N_20851,N_20907);
and U21036 (N_21036,N_20960,N_20904);
nor U21037 (N_21037,N_20733,N_20925);
nor U21038 (N_21038,N_20727,N_20963);
xor U21039 (N_21039,N_20849,N_20973);
and U21040 (N_21040,N_20825,N_20846);
or U21041 (N_21041,N_20926,N_20984);
and U21042 (N_21042,N_20730,N_20766);
nand U21043 (N_21043,N_20923,N_20816);
nor U21044 (N_21044,N_20714,N_20935);
and U21045 (N_21045,N_20784,N_20928);
xnor U21046 (N_21046,N_20995,N_20791);
xnor U21047 (N_21047,N_20800,N_20858);
nor U21048 (N_21048,N_20720,N_20789);
or U21049 (N_21049,N_20769,N_20990);
nor U21050 (N_21050,N_20718,N_20905);
nor U21051 (N_21051,N_20951,N_20762);
and U21052 (N_21052,N_20814,N_20801);
nor U21053 (N_21053,N_20763,N_20748);
and U21054 (N_21054,N_20725,N_20886);
nand U21055 (N_21055,N_20844,N_20946);
or U21056 (N_21056,N_20987,N_20921);
nand U21057 (N_21057,N_20865,N_20949);
or U21058 (N_21058,N_20768,N_20971);
xnor U21059 (N_21059,N_20950,N_20961);
nor U21060 (N_21060,N_20879,N_20777);
xor U21061 (N_21061,N_20761,N_20796);
and U21062 (N_21062,N_20897,N_20756);
or U21063 (N_21063,N_20867,N_20708);
nor U21064 (N_21064,N_20739,N_20892);
nand U21065 (N_21065,N_20919,N_20875);
or U21066 (N_21066,N_20988,N_20752);
xor U21067 (N_21067,N_20747,N_20750);
xor U21068 (N_21068,N_20932,N_20978);
and U21069 (N_21069,N_20953,N_20852);
and U21070 (N_21070,N_20927,N_20770);
and U21071 (N_21071,N_20872,N_20703);
nor U21072 (N_21072,N_20918,N_20836);
nor U21073 (N_21073,N_20716,N_20983);
nand U21074 (N_21074,N_20884,N_20991);
or U21075 (N_21075,N_20911,N_20772);
nand U21076 (N_21076,N_20952,N_20778);
nand U21077 (N_21077,N_20712,N_20794);
nand U21078 (N_21078,N_20916,N_20764);
and U21079 (N_21079,N_20894,N_20823);
xor U21080 (N_21080,N_20797,N_20742);
and U21081 (N_21081,N_20837,N_20989);
xnor U21082 (N_21082,N_20917,N_20826);
or U21083 (N_21083,N_20832,N_20705);
or U21084 (N_21084,N_20807,N_20833);
nand U21085 (N_21085,N_20713,N_20888);
xor U21086 (N_21086,N_20855,N_20974);
nand U21087 (N_21087,N_20835,N_20930);
or U21088 (N_21088,N_20743,N_20931);
xor U21089 (N_21089,N_20829,N_20954);
nor U21090 (N_21090,N_20788,N_20899);
xnor U21091 (N_21091,N_20734,N_20707);
nand U21092 (N_21092,N_20811,N_20885);
nand U21093 (N_21093,N_20785,N_20975);
nor U21094 (N_21094,N_20738,N_20857);
nand U21095 (N_21095,N_20936,N_20906);
or U21096 (N_21096,N_20937,N_20817);
xnor U21097 (N_21097,N_20962,N_20895);
nand U21098 (N_21098,N_20700,N_20964);
xor U21099 (N_21099,N_20856,N_20850);
nand U21100 (N_21100,N_20854,N_20878);
nand U21101 (N_21101,N_20809,N_20818);
nor U21102 (N_21102,N_20948,N_20986);
nand U21103 (N_21103,N_20992,N_20760);
or U21104 (N_21104,N_20798,N_20732);
nand U21105 (N_21105,N_20771,N_20793);
nor U21106 (N_21106,N_20736,N_20731);
and U21107 (N_21107,N_20996,N_20744);
and U21108 (N_21108,N_20795,N_20711);
and U21109 (N_21109,N_20860,N_20868);
or U21110 (N_21110,N_20863,N_20831);
xor U21111 (N_21111,N_20722,N_20965);
nor U21112 (N_21112,N_20968,N_20891);
nor U21113 (N_21113,N_20887,N_20841);
and U21114 (N_21114,N_20847,N_20781);
or U21115 (N_21115,N_20767,N_20804);
xor U21116 (N_21116,N_20981,N_20827);
and U21117 (N_21117,N_20819,N_20859);
or U21118 (N_21118,N_20883,N_20805);
nand U21119 (N_21119,N_20929,N_20728);
and U21120 (N_21120,N_20822,N_20754);
nor U21121 (N_21121,N_20704,N_20997);
or U21122 (N_21122,N_20880,N_20821);
xnor U21123 (N_21123,N_20943,N_20994);
nand U21124 (N_21124,N_20862,N_20780);
nand U21125 (N_21125,N_20881,N_20877);
nor U21126 (N_21126,N_20956,N_20924);
and U21127 (N_21127,N_20787,N_20909);
nand U21128 (N_21128,N_20702,N_20773);
nor U21129 (N_21129,N_20824,N_20751);
xnor U21130 (N_21130,N_20845,N_20701);
nor U21131 (N_21131,N_20757,N_20861);
nor U21132 (N_21132,N_20810,N_20959);
xor U21133 (N_21133,N_20746,N_20882);
xnor U21134 (N_21134,N_20977,N_20940);
and U21135 (N_21135,N_20755,N_20759);
xor U21136 (N_21136,N_20934,N_20913);
or U21137 (N_21137,N_20999,N_20774);
xnor U21138 (N_21138,N_20820,N_20941);
nand U21139 (N_21139,N_20920,N_20908);
nor U21140 (N_21140,N_20792,N_20980);
nor U21141 (N_21141,N_20782,N_20970);
and U21142 (N_21142,N_20715,N_20900);
or U21143 (N_21143,N_20779,N_20853);
and U21144 (N_21144,N_20719,N_20873);
nor U21145 (N_21145,N_20896,N_20915);
xnor U21146 (N_21146,N_20783,N_20830);
nand U21147 (N_21147,N_20815,N_20933);
and U21148 (N_21148,N_20842,N_20753);
or U21149 (N_21149,N_20898,N_20709);
xor U21150 (N_21150,N_20747,N_20973);
nand U21151 (N_21151,N_20768,N_20985);
nand U21152 (N_21152,N_20815,N_20734);
nand U21153 (N_21153,N_20866,N_20727);
xor U21154 (N_21154,N_20940,N_20922);
xor U21155 (N_21155,N_20839,N_20771);
or U21156 (N_21156,N_20754,N_20809);
or U21157 (N_21157,N_20864,N_20937);
and U21158 (N_21158,N_20890,N_20926);
nand U21159 (N_21159,N_20811,N_20981);
or U21160 (N_21160,N_20953,N_20723);
xnor U21161 (N_21161,N_20988,N_20978);
nand U21162 (N_21162,N_20717,N_20894);
and U21163 (N_21163,N_20986,N_20770);
xor U21164 (N_21164,N_20864,N_20989);
or U21165 (N_21165,N_20921,N_20781);
xnor U21166 (N_21166,N_20904,N_20917);
nor U21167 (N_21167,N_20860,N_20816);
or U21168 (N_21168,N_20705,N_20908);
nand U21169 (N_21169,N_20754,N_20863);
xnor U21170 (N_21170,N_20829,N_20828);
or U21171 (N_21171,N_20948,N_20765);
and U21172 (N_21172,N_20782,N_20764);
or U21173 (N_21173,N_20924,N_20968);
nor U21174 (N_21174,N_20837,N_20986);
and U21175 (N_21175,N_20768,N_20846);
nor U21176 (N_21176,N_20806,N_20720);
or U21177 (N_21177,N_20912,N_20868);
nor U21178 (N_21178,N_20831,N_20970);
nand U21179 (N_21179,N_20963,N_20905);
xor U21180 (N_21180,N_20777,N_20961);
or U21181 (N_21181,N_20746,N_20911);
and U21182 (N_21182,N_20772,N_20776);
nand U21183 (N_21183,N_20924,N_20758);
nand U21184 (N_21184,N_20760,N_20996);
and U21185 (N_21185,N_20876,N_20891);
nor U21186 (N_21186,N_20853,N_20928);
nor U21187 (N_21187,N_20800,N_20889);
xnor U21188 (N_21188,N_20968,N_20991);
nor U21189 (N_21189,N_20757,N_20793);
or U21190 (N_21190,N_20879,N_20898);
xnor U21191 (N_21191,N_20708,N_20974);
or U21192 (N_21192,N_20788,N_20910);
xnor U21193 (N_21193,N_20746,N_20866);
or U21194 (N_21194,N_20982,N_20905);
nor U21195 (N_21195,N_20790,N_20779);
nor U21196 (N_21196,N_20724,N_20970);
xor U21197 (N_21197,N_20990,N_20992);
and U21198 (N_21198,N_20849,N_20799);
xor U21199 (N_21199,N_20912,N_20890);
or U21200 (N_21200,N_20818,N_20916);
xnor U21201 (N_21201,N_20760,N_20953);
nor U21202 (N_21202,N_20973,N_20972);
or U21203 (N_21203,N_20924,N_20907);
nand U21204 (N_21204,N_20712,N_20919);
and U21205 (N_21205,N_20749,N_20839);
nand U21206 (N_21206,N_20984,N_20873);
or U21207 (N_21207,N_20987,N_20947);
or U21208 (N_21208,N_20879,N_20710);
nor U21209 (N_21209,N_20969,N_20765);
and U21210 (N_21210,N_20896,N_20989);
nand U21211 (N_21211,N_20954,N_20828);
or U21212 (N_21212,N_20839,N_20801);
nand U21213 (N_21213,N_20823,N_20841);
nand U21214 (N_21214,N_20755,N_20789);
nand U21215 (N_21215,N_20782,N_20778);
xor U21216 (N_21216,N_20888,N_20871);
xnor U21217 (N_21217,N_20982,N_20918);
or U21218 (N_21218,N_20910,N_20968);
or U21219 (N_21219,N_20994,N_20885);
or U21220 (N_21220,N_20808,N_20896);
nand U21221 (N_21221,N_20743,N_20813);
or U21222 (N_21222,N_20796,N_20989);
xnor U21223 (N_21223,N_20919,N_20853);
xnor U21224 (N_21224,N_20808,N_20921);
xnor U21225 (N_21225,N_20787,N_20776);
xor U21226 (N_21226,N_20971,N_20719);
xor U21227 (N_21227,N_20823,N_20721);
xor U21228 (N_21228,N_20700,N_20818);
xnor U21229 (N_21229,N_20826,N_20719);
xor U21230 (N_21230,N_20751,N_20876);
and U21231 (N_21231,N_20930,N_20885);
and U21232 (N_21232,N_20950,N_20704);
nand U21233 (N_21233,N_20711,N_20864);
nand U21234 (N_21234,N_20891,N_20847);
xnor U21235 (N_21235,N_20807,N_20868);
nand U21236 (N_21236,N_20748,N_20877);
nand U21237 (N_21237,N_20741,N_20878);
nor U21238 (N_21238,N_20716,N_20881);
nor U21239 (N_21239,N_20743,N_20963);
and U21240 (N_21240,N_20704,N_20969);
and U21241 (N_21241,N_20762,N_20815);
or U21242 (N_21242,N_20921,N_20853);
and U21243 (N_21243,N_20712,N_20882);
nor U21244 (N_21244,N_20861,N_20772);
nor U21245 (N_21245,N_20860,N_20882);
nor U21246 (N_21246,N_20812,N_20889);
nand U21247 (N_21247,N_20902,N_20909);
xnor U21248 (N_21248,N_20776,N_20767);
xor U21249 (N_21249,N_20810,N_20971);
xor U21250 (N_21250,N_20902,N_20764);
xor U21251 (N_21251,N_20791,N_20730);
or U21252 (N_21252,N_20790,N_20894);
nor U21253 (N_21253,N_20896,N_20718);
or U21254 (N_21254,N_20897,N_20783);
nand U21255 (N_21255,N_20968,N_20725);
nor U21256 (N_21256,N_20837,N_20992);
nor U21257 (N_21257,N_20948,N_20995);
nor U21258 (N_21258,N_20957,N_20781);
xnor U21259 (N_21259,N_20897,N_20892);
xor U21260 (N_21260,N_20986,N_20769);
nor U21261 (N_21261,N_20895,N_20727);
or U21262 (N_21262,N_20799,N_20764);
nor U21263 (N_21263,N_20827,N_20890);
xor U21264 (N_21264,N_20733,N_20927);
nor U21265 (N_21265,N_20872,N_20802);
xor U21266 (N_21266,N_20869,N_20739);
nand U21267 (N_21267,N_20860,N_20749);
or U21268 (N_21268,N_20802,N_20904);
or U21269 (N_21269,N_20865,N_20819);
and U21270 (N_21270,N_20711,N_20750);
and U21271 (N_21271,N_20754,N_20715);
or U21272 (N_21272,N_20781,N_20907);
nand U21273 (N_21273,N_20993,N_20741);
xnor U21274 (N_21274,N_20724,N_20767);
nand U21275 (N_21275,N_20866,N_20993);
and U21276 (N_21276,N_20756,N_20840);
nand U21277 (N_21277,N_20705,N_20947);
nand U21278 (N_21278,N_20896,N_20737);
and U21279 (N_21279,N_20910,N_20750);
nor U21280 (N_21280,N_20741,N_20880);
xor U21281 (N_21281,N_20800,N_20801);
nand U21282 (N_21282,N_20883,N_20761);
and U21283 (N_21283,N_20778,N_20847);
nand U21284 (N_21284,N_20763,N_20898);
and U21285 (N_21285,N_20746,N_20725);
nor U21286 (N_21286,N_20711,N_20965);
nor U21287 (N_21287,N_20714,N_20753);
xor U21288 (N_21288,N_20737,N_20814);
or U21289 (N_21289,N_20813,N_20805);
xnor U21290 (N_21290,N_20941,N_20986);
nand U21291 (N_21291,N_20822,N_20865);
nor U21292 (N_21292,N_20872,N_20824);
and U21293 (N_21293,N_20959,N_20901);
xnor U21294 (N_21294,N_20769,N_20897);
nand U21295 (N_21295,N_20702,N_20850);
nand U21296 (N_21296,N_20742,N_20926);
xor U21297 (N_21297,N_20930,N_20782);
or U21298 (N_21298,N_20937,N_20777);
nand U21299 (N_21299,N_20988,N_20945);
and U21300 (N_21300,N_21158,N_21058);
nor U21301 (N_21301,N_21039,N_21219);
and U21302 (N_21302,N_21184,N_21253);
nand U21303 (N_21303,N_21147,N_21157);
nor U21304 (N_21304,N_21141,N_21212);
nand U21305 (N_21305,N_21074,N_21086);
and U21306 (N_21306,N_21062,N_21026);
nand U21307 (N_21307,N_21188,N_21270);
nor U21308 (N_21308,N_21137,N_21131);
nor U21309 (N_21309,N_21136,N_21056);
and U21310 (N_21310,N_21229,N_21071);
nand U21311 (N_21311,N_21012,N_21292);
nand U21312 (N_21312,N_21268,N_21140);
or U21313 (N_21313,N_21132,N_21087);
nand U21314 (N_21314,N_21149,N_21159);
or U21315 (N_21315,N_21207,N_21231);
nor U21316 (N_21316,N_21028,N_21284);
nand U21317 (N_21317,N_21198,N_21075);
nor U21318 (N_21318,N_21218,N_21000);
nand U21319 (N_21319,N_21102,N_21034);
nand U21320 (N_21320,N_21023,N_21274);
and U21321 (N_21321,N_21122,N_21264);
nand U21322 (N_21322,N_21142,N_21020);
nor U21323 (N_21323,N_21276,N_21155);
xor U21324 (N_21324,N_21024,N_21234);
or U21325 (N_21325,N_21297,N_21106);
or U21326 (N_21326,N_21008,N_21230);
or U21327 (N_21327,N_21232,N_21088);
or U21328 (N_21328,N_21053,N_21279);
xor U21329 (N_21329,N_21113,N_21240);
and U21330 (N_21330,N_21293,N_21070);
or U21331 (N_21331,N_21180,N_21041);
and U21332 (N_21332,N_21258,N_21045);
nand U21333 (N_21333,N_21164,N_21003);
or U21334 (N_21334,N_21223,N_21037);
or U21335 (N_21335,N_21126,N_21153);
and U21336 (N_21336,N_21295,N_21171);
and U21337 (N_21337,N_21195,N_21022);
xnor U21338 (N_21338,N_21162,N_21151);
xnor U21339 (N_21339,N_21092,N_21044);
or U21340 (N_21340,N_21260,N_21254);
nand U21341 (N_21341,N_21204,N_21046);
xor U21342 (N_21342,N_21108,N_21049);
and U21343 (N_21343,N_21082,N_21233);
nor U21344 (N_21344,N_21063,N_21201);
nor U21345 (N_21345,N_21123,N_21291);
nand U21346 (N_21346,N_21081,N_21133);
nor U21347 (N_21347,N_21093,N_21181);
nor U21348 (N_21348,N_21249,N_21226);
or U21349 (N_21349,N_21047,N_21196);
xnor U21350 (N_21350,N_21298,N_21269);
nand U21351 (N_21351,N_21006,N_21121);
xnor U21352 (N_21352,N_21128,N_21032);
and U21353 (N_21353,N_21169,N_21160);
nor U21354 (N_21354,N_21222,N_21239);
and U21355 (N_21355,N_21055,N_21064);
xor U21356 (N_21356,N_21257,N_21124);
nor U21357 (N_21357,N_21031,N_21144);
nand U21358 (N_21358,N_21210,N_21033);
xnor U21359 (N_21359,N_21192,N_21067);
nor U21360 (N_21360,N_21060,N_21101);
xnor U21361 (N_21361,N_21110,N_21073);
and U21362 (N_21362,N_21085,N_21005);
or U21363 (N_21363,N_21263,N_21294);
nor U21364 (N_21364,N_21089,N_21272);
or U21365 (N_21365,N_21130,N_21256);
nand U21366 (N_21366,N_21217,N_21095);
or U21367 (N_21367,N_21096,N_21245);
nand U21368 (N_21368,N_21127,N_21115);
nor U21369 (N_21369,N_21135,N_21007);
xor U21370 (N_21370,N_21134,N_21271);
nand U21371 (N_21371,N_21100,N_21083);
xnor U21372 (N_21372,N_21069,N_21167);
and U21373 (N_21373,N_21038,N_21154);
nor U21374 (N_21374,N_21072,N_21139);
nand U21375 (N_21375,N_21287,N_21103);
nor U21376 (N_21376,N_21027,N_21138);
or U21377 (N_21377,N_21221,N_21199);
nor U21378 (N_21378,N_21161,N_21237);
xnor U21379 (N_21379,N_21191,N_21225);
nand U21380 (N_21380,N_21143,N_21211);
nor U21381 (N_21381,N_21048,N_21009);
xor U21382 (N_21382,N_21277,N_21014);
and U21383 (N_21383,N_21290,N_21107);
or U21384 (N_21384,N_21275,N_21116);
xnor U21385 (N_21385,N_21203,N_21059);
nor U21386 (N_21386,N_21112,N_21261);
nor U21387 (N_21387,N_21016,N_21120);
or U21388 (N_21388,N_21266,N_21068);
nand U21389 (N_21389,N_21241,N_21090);
nor U21390 (N_21390,N_21285,N_21170);
nand U21391 (N_21391,N_21235,N_21145);
or U21392 (N_21392,N_21015,N_21118);
xnor U21393 (N_21393,N_21104,N_21019);
nand U21394 (N_21394,N_21078,N_21246);
or U21395 (N_21395,N_21156,N_21238);
or U21396 (N_21396,N_21057,N_21010);
and U21397 (N_21397,N_21148,N_21187);
nand U21398 (N_21398,N_21030,N_21267);
or U21399 (N_21399,N_21172,N_21215);
and U21400 (N_21400,N_21111,N_21066);
nand U21401 (N_21401,N_21176,N_21175);
or U21402 (N_21402,N_21043,N_21190);
xor U21403 (N_21403,N_21146,N_21098);
xor U21404 (N_21404,N_21163,N_21165);
nand U21405 (N_21405,N_21150,N_21105);
and U21406 (N_21406,N_21109,N_21174);
nand U21407 (N_21407,N_21202,N_21099);
and U21408 (N_21408,N_21243,N_21252);
nand U21409 (N_21409,N_21004,N_21017);
nand U21410 (N_21410,N_21236,N_21193);
or U21411 (N_21411,N_21227,N_21050);
nand U21412 (N_21412,N_21025,N_21255);
xnor U21413 (N_21413,N_21280,N_21296);
xor U21414 (N_21414,N_21054,N_21248);
xor U21415 (N_21415,N_21189,N_21289);
nand U21416 (N_21416,N_21094,N_21288);
nor U21417 (N_21417,N_21011,N_21042);
nand U21418 (N_21418,N_21278,N_21018);
nor U21419 (N_21419,N_21200,N_21080);
or U21420 (N_21420,N_21065,N_21265);
and U21421 (N_21421,N_21051,N_21299);
xnor U21422 (N_21422,N_21077,N_21129);
nor U21423 (N_21423,N_21168,N_21117);
nor U21424 (N_21424,N_21282,N_21262);
xnor U21425 (N_21425,N_21179,N_21040);
nor U21426 (N_21426,N_21247,N_21224);
or U21427 (N_21427,N_21213,N_21084);
nand U21428 (N_21428,N_21205,N_21021);
xor U21429 (N_21429,N_21125,N_21061);
and U21430 (N_21430,N_21197,N_21029);
nand U21431 (N_21431,N_21283,N_21182);
nand U21432 (N_21432,N_21250,N_21001);
and U21433 (N_21433,N_21242,N_21097);
and U21434 (N_21434,N_21002,N_21206);
and U21435 (N_21435,N_21185,N_21152);
nor U21436 (N_21436,N_21183,N_21251);
nor U21437 (N_21437,N_21209,N_21220);
nand U21438 (N_21438,N_21035,N_21208);
nor U21439 (N_21439,N_21036,N_21194);
or U21440 (N_21440,N_21114,N_21281);
nand U21441 (N_21441,N_21013,N_21178);
nor U21442 (N_21442,N_21177,N_21186);
xnor U21443 (N_21443,N_21216,N_21052);
and U21444 (N_21444,N_21173,N_21091);
and U21445 (N_21445,N_21273,N_21214);
xnor U21446 (N_21446,N_21119,N_21079);
and U21447 (N_21447,N_21244,N_21286);
nor U21448 (N_21448,N_21259,N_21228);
and U21449 (N_21449,N_21076,N_21166);
nand U21450 (N_21450,N_21270,N_21261);
and U21451 (N_21451,N_21299,N_21278);
and U21452 (N_21452,N_21169,N_21212);
nor U21453 (N_21453,N_21239,N_21035);
xor U21454 (N_21454,N_21289,N_21266);
and U21455 (N_21455,N_21118,N_21045);
and U21456 (N_21456,N_21169,N_21126);
xor U21457 (N_21457,N_21233,N_21155);
xor U21458 (N_21458,N_21258,N_21041);
xor U21459 (N_21459,N_21290,N_21219);
nand U21460 (N_21460,N_21178,N_21248);
nor U21461 (N_21461,N_21286,N_21102);
xor U21462 (N_21462,N_21287,N_21120);
nor U21463 (N_21463,N_21132,N_21013);
or U21464 (N_21464,N_21026,N_21295);
xnor U21465 (N_21465,N_21018,N_21216);
nor U21466 (N_21466,N_21288,N_21065);
nand U21467 (N_21467,N_21063,N_21106);
xor U21468 (N_21468,N_21238,N_21031);
or U21469 (N_21469,N_21077,N_21144);
or U21470 (N_21470,N_21242,N_21137);
or U21471 (N_21471,N_21000,N_21281);
and U21472 (N_21472,N_21229,N_21203);
or U21473 (N_21473,N_21180,N_21010);
nand U21474 (N_21474,N_21012,N_21279);
nor U21475 (N_21475,N_21046,N_21111);
xnor U21476 (N_21476,N_21144,N_21176);
or U21477 (N_21477,N_21176,N_21285);
and U21478 (N_21478,N_21052,N_21059);
xnor U21479 (N_21479,N_21297,N_21027);
nand U21480 (N_21480,N_21280,N_21216);
and U21481 (N_21481,N_21255,N_21136);
nor U21482 (N_21482,N_21232,N_21097);
nor U21483 (N_21483,N_21291,N_21134);
and U21484 (N_21484,N_21021,N_21222);
nand U21485 (N_21485,N_21132,N_21269);
nand U21486 (N_21486,N_21046,N_21047);
or U21487 (N_21487,N_21125,N_21076);
nor U21488 (N_21488,N_21000,N_21010);
nor U21489 (N_21489,N_21291,N_21129);
xor U21490 (N_21490,N_21217,N_21299);
xor U21491 (N_21491,N_21056,N_21235);
and U21492 (N_21492,N_21245,N_21233);
xor U21493 (N_21493,N_21115,N_21262);
and U21494 (N_21494,N_21005,N_21167);
xor U21495 (N_21495,N_21288,N_21081);
nor U21496 (N_21496,N_21278,N_21106);
nor U21497 (N_21497,N_21205,N_21108);
nor U21498 (N_21498,N_21124,N_21136);
xnor U21499 (N_21499,N_21280,N_21247);
xnor U21500 (N_21500,N_21007,N_21182);
and U21501 (N_21501,N_21097,N_21052);
xor U21502 (N_21502,N_21271,N_21109);
and U21503 (N_21503,N_21057,N_21238);
nand U21504 (N_21504,N_21092,N_21233);
nor U21505 (N_21505,N_21294,N_21111);
or U21506 (N_21506,N_21010,N_21178);
nand U21507 (N_21507,N_21095,N_21182);
or U21508 (N_21508,N_21286,N_21105);
or U21509 (N_21509,N_21212,N_21281);
and U21510 (N_21510,N_21240,N_21297);
nand U21511 (N_21511,N_21132,N_21121);
nand U21512 (N_21512,N_21003,N_21137);
nor U21513 (N_21513,N_21204,N_21167);
nor U21514 (N_21514,N_21084,N_21161);
and U21515 (N_21515,N_21269,N_21085);
nand U21516 (N_21516,N_21255,N_21016);
nor U21517 (N_21517,N_21264,N_21179);
and U21518 (N_21518,N_21128,N_21003);
nand U21519 (N_21519,N_21269,N_21070);
nor U21520 (N_21520,N_21280,N_21090);
nor U21521 (N_21521,N_21071,N_21007);
nand U21522 (N_21522,N_21046,N_21276);
nor U21523 (N_21523,N_21046,N_21153);
and U21524 (N_21524,N_21083,N_21030);
or U21525 (N_21525,N_21180,N_21159);
or U21526 (N_21526,N_21282,N_21098);
or U21527 (N_21527,N_21254,N_21019);
nor U21528 (N_21528,N_21243,N_21255);
nand U21529 (N_21529,N_21191,N_21164);
and U21530 (N_21530,N_21079,N_21216);
xor U21531 (N_21531,N_21220,N_21073);
nand U21532 (N_21532,N_21181,N_21296);
or U21533 (N_21533,N_21296,N_21165);
nor U21534 (N_21534,N_21245,N_21123);
xor U21535 (N_21535,N_21253,N_21043);
or U21536 (N_21536,N_21133,N_21027);
and U21537 (N_21537,N_21206,N_21154);
or U21538 (N_21538,N_21149,N_21059);
and U21539 (N_21539,N_21186,N_21248);
nor U21540 (N_21540,N_21263,N_21284);
nand U21541 (N_21541,N_21205,N_21296);
and U21542 (N_21542,N_21062,N_21148);
xor U21543 (N_21543,N_21235,N_21271);
and U21544 (N_21544,N_21164,N_21206);
xnor U21545 (N_21545,N_21102,N_21190);
nand U21546 (N_21546,N_21106,N_21190);
nor U21547 (N_21547,N_21070,N_21020);
nor U21548 (N_21548,N_21229,N_21234);
or U21549 (N_21549,N_21006,N_21199);
nor U21550 (N_21550,N_21088,N_21086);
nor U21551 (N_21551,N_21285,N_21273);
or U21552 (N_21552,N_21253,N_21002);
nor U21553 (N_21553,N_21247,N_21137);
xor U21554 (N_21554,N_21298,N_21167);
nor U21555 (N_21555,N_21109,N_21298);
nand U21556 (N_21556,N_21296,N_21081);
nor U21557 (N_21557,N_21017,N_21252);
nor U21558 (N_21558,N_21147,N_21012);
or U21559 (N_21559,N_21257,N_21153);
or U21560 (N_21560,N_21207,N_21180);
or U21561 (N_21561,N_21105,N_21017);
nor U21562 (N_21562,N_21222,N_21140);
or U21563 (N_21563,N_21098,N_21193);
nor U21564 (N_21564,N_21147,N_21017);
or U21565 (N_21565,N_21249,N_21205);
nor U21566 (N_21566,N_21106,N_21041);
and U21567 (N_21567,N_21041,N_21164);
nand U21568 (N_21568,N_21034,N_21064);
and U21569 (N_21569,N_21173,N_21277);
and U21570 (N_21570,N_21133,N_21146);
nor U21571 (N_21571,N_21280,N_21226);
xnor U21572 (N_21572,N_21045,N_21295);
nor U21573 (N_21573,N_21163,N_21258);
and U21574 (N_21574,N_21002,N_21031);
nand U21575 (N_21575,N_21178,N_21103);
or U21576 (N_21576,N_21156,N_21039);
and U21577 (N_21577,N_21079,N_21016);
nor U21578 (N_21578,N_21204,N_21147);
nor U21579 (N_21579,N_21236,N_21249);
xor U21580 (N_21580,N_21080,N_21204);
xnor U21581 (N_21581,N_21288,N_21178);
xor U21582 (N_21582,N_21239,N_21200);
or U21583 (N_21583,N_21178,N_21093);
xor U21584 (N_21584,N_21203,N_21032);
xnor U21585 (N_21585,N_21045,N_21086);
or U21586 (N_21586,N_21138,N_21040);
nor U21587 (N_21587,N_21252,N_21273);
xor U21588 (N_21588,N_21264,N_21185);
xor U21589 (N_21589,N_21230,N_21135);
nor U21590 (N_21590,N_21141,N_21224);
xnor U21591 (N_21591,N_21055,N_21181);
xnor U21592 (N_21592,N_21248,N_21139);
or U21593 (N_21593,N_21048,N_21127);
xnor U21594 (N_21594,N_21275,N_21288);
or U21595 (N_21595,N_21124,N_21229);
or U21596 (N_21596,N_21240,N_21122);
nand U21597 (N_21597,N_21263,N_21135);
and U21598 (N_21598,N_21011,N_21120);
xor U21599 (N_21599,N_21118,N_21084);
xor U21600 (N_21600,N_21363,N_21575);
xnor U21601 (N_21601,N_21342,N_21588);
xor U21602 (N_21602,N_21541,N_21311);
nor U21603 (N_21603,N_21386,N_21312);
xnor U21604 (N_21604,N_21550,N_21561);
xor U21605 (N_21605,N_21430,N_21548);
nand U21606 (N_21606,N_21437,N_21562);
nor U21607 (N_21607,N_21338,N_21416);
xnor U21608 (N_21608,N_21354,N_21489);
nor U21609 (N_21609,N_21343,N_21563);
xor U21610 (N_21610,N_21525,N_21579);
nand U21611 (N_21611,N_21301,N_21493);
xnor U21612 (N_21612,N_21320,N_21411);
and U21613 (N_21613,N_21417,N_21572);
nand U21614 (N_21614,N_21467,N_21487);
xnor U21615 (N_21615,N_21332,N_21536);
nand U21616 (N_21616,N_21454,N_21351);
nor U21617 (N_21617,N_21452,N_21466);
xnor U21618 (N_21618,N_21389,N_21453);
or U21619 (N_21619,N_21341,N_21462);
and U21620 (N_21620,N_21500,N_21576);
and U21621 (N_21621,N_21323,N_21414);
nand U21622 (N_21622,N_21427,N_21463);
xor U21623 (N_21623,N_21506,N_21584);
nand U21624 (N_21624,N_21551,N_21420);
nor U21625 (N_21625,N_21365,N_21438);
xnor U21626 (N_21626,N_21574,N_21464);
nand U21627 (N_21627,N_21486,N_21549);
nor U21628 (N_21628,N_21499,N_21415);
nor U21629 (N_21629,N_21592,N_21508);
nor U21630 (N_21630,N_21564,N_21393);
nor U21631 (N_21631,N_21359,N_21475);
xnor U21632 (N_21632,N_21520,N_21306);
nand U21633 (N_21633,N_21317,N_21587);
nor U21634 (N_21634,N_21374,N_21378);
nand U21635 (N_21635,N_21503,N_21510);
and U21636 (N_21636,N_21322,N_21367);
or U21637 (N_21637,N_21349,N_21529);
or U21638 (N_21638,N_21325,N_21539);
xnor U21639 (N_21639,N_21441,N_21540);
xnor U21640 (N_21640,N_21511,N_21522);
and U21641 (N_21641,N_21350,N_21461);
nand U21642 (N_21642,N_21329,N_21364);
or U21643 (N_21643,N_21469,N_21410);
nand U21644 (N_21644,N_21566,N_21392);
or U21645 (N_21645,N_21305,N_21412);
or U21646 (N_21646,N_21482,N_21335);
and U21647 (N_21647,N_21308,N_21568);
nand U21648 (N_21648,N_21483,N_21547);
nor U21649 (N_21649,N_21560,N_21362);
xnor U21650 (N_21650,N_21396,N_21593);
or U21651 (N_21651,N_21513,N_21450);
nor U21652 (N_21652,N_21456,N_21418);
or U21653 (N_21653,N_21528,N_21388);
nand U21654 (N_21654,N_21553,N_21451);
nor U21655 (N_21655,N_21490,N_21316);
and U21656 (N_21656,N_21457,N_21569);
or U21657 (N_21657,N_21470,N_21313);
or U21658 (N_21658,N_21433,N_21431);
nor U21659 (N_21659,N_21491,N_21533);
and U21660 (N_21660,N_21479,N_21333);
nor U21661 (N_21661,N_21434,N_21399);
xnor U21662 (N_21662,N_21358,N_21385);
nand U21663 (N_21663,N_21556,N_21406);
and U21664 (N_21664,N_21543,N_21442);
xor U21665 (N_21665,N_21555,N_21348);
nor U21666 (N_21666,N_21360,N_21402);
or U21667 (N_21667,N_21355,N_21405);
xor U21668 (N_21668,N_21518,N_21580);
xnor U21669 (N_21669,N_21315,N_21419);
and U21670 (N_21670,N_21379,N_21391);
or U21671 (N_21671,N_21460,N_21435);
xor U21672 (N_21672,N_21368,N_21559);
or U21673 (N_21673,N_21309,N_21492);
xor U21674 (N_21674,N_21570,N_21484);
or U21675 (N_21675,N_21408,N_21404);
nor U21676 (N_21676,N_21326,N_21449);
and U21677 (N_21677,N_21459,N_21573);
nor U21678 (N_21678,N_21524,N_21577);
or U21679 (N_21679,N_21432,N_21502);
xnor U21680 (N_21680,N_21595,N_21465);
xor U21681 (N_21681,N_21447,N_21324);
nor U21682 (N_21682,N_21585,N_21421);
nand U21683 (N_21683,N_21303,N_21425);
or U21684 (N_21684,N_21331,N_21497);
nand U21685 (N_21685,N_21599,N_21527);
and U21686 (N_21686,N_21485,N_21477);
xor U21687 (N_21687,N_21336,N_21407);
and U21688 (N_21688,N_21554,N_21480);
or U21689 (N_21689,N_21488,N_21346);
and U21690 (N_21690,N_21302,N_21481);
nand U21691 (N_21691,N_21304,N_21376);
or U21692 (N_21692,N_21429,N_21307);
or U21693 (N_21693,N_21443,N_21413);
nor U21694 (N_21694,N_21353,N_21591);
and U21695 (N_21695,N_21571,N_21590);
nand U21696 (N_21696,N_21321,N_21337);
and U21697 (N_21697,N_21496,N_21468);
or U21698 (N_21698,N_21340,N_21426);
nor U21699 (N_21699,N_21546,N_21361);
or U21700 (N_21700,N_21501,N_21531);
nor U21701 (N_21701,N_21319,N_21330);
and U21702 (N_21702,N_21473,N_21381);
and U21703 (N_21703,N_21448,N_21370);
nor U21704 (N_21704,N_21589,N_21474);
xor U21705 (N_21705,N_21395,N_21383);
nor U21706 (N_21706,N_21565,N_21398);
and U21707 (N_21707,N_21310,N_21345);
or U21708 (N_21708,N_21538,N_21422);
and U21709 (N_21709,N_21428,N_21424);
nor U21710 (N_21710,N_21517,N_21382);
nand U21711 (N_21711,N_21523,N_21444);
nand U21712 (N_21712,N_21458,N_21401);
nand U21713 (N_21713,N_21400,N_21446);
xnor U21714 (N_21714,N_21472,N_21544);
nand U21715 (N_21715,N_21471,N_21372);
and U21716 (N_21716,N_21476,N_21515);
and U21717 (N_21717,N_21594,N_21334);
nor U21718 (N_21718,N_21439,N_21534);
or U21719 (N_21719,N_21567,N_21328);
nor U21720 (N_21720,N_21318,N_21445);
nor U21721 (N_21721,N_21526,N_21380);
nand U21722 (N_21722,N_21586,N_21558);
and U21723 (N_21723,N_21516,N_21582);
nand U21724 (N_21724,N_21514,N_21300);
xor U21725 (N_21725,N_21583,N_21519);
nand U21726 (N_21726,N_21581,N_21403);
nand U21727 (N_21727,N_21498,N_21545);
and U21728 (N_21728,N_21507,N_21505);
and U21729 (N_21729,N_21596,N_21532);
or U21730 (N_21730,N_21535,N_21352);
nor U21731 (N_21731,N_21356,N_21598);
nand U21732 (N_21732,N_21377,N_21357);
nor U21733 (N_21733,N_21436,N_21530);
nor U21734 (N_21734,N_21455,N_21597);
or U21735 (N_21735,N_21339,N_21423);
nand U21736 (N_21736,N_21390,N_21521);
nor U21737 (N_21737,N_21394,N_21552);
nand U21738 (N_21738,N_21542,N_21347);
and U21739 (N_21739,N_21557,N_21375);
xnor U21740 (N_21740,N_21504,N_21495);
nand U21741 (N_21741,N_21509,N_21409);
and U21742 (N_21742,N_21369,N_21512);
or U21743 (N_21743,N_21371,N_21366);
and U21744 (N_21744,N_21314,N_21327);
xor U21745 (N_21745,N_21494,N_21578);
nand U21746 (N_21746,N_21344,N_21478);
or U21747 (N_21747,N_21397,N_21373);
or U21748 (N_21748,N_21387,N_21440);
nand U21749 (N_21749,N_21537,N_21384);
nand U21750 (N_21750,N_21440,N_21490);
or U21751 (N_21751,N_21406,N_21347);
and U21752 (N_21752,N_21545,N_21310);
nand U21753 (N_21753,N_21358,N_21304);
nand U21754 (N_21754,N_21598,N_21369);
or U21755 (N_21755,N_21419,N_21597);
xor U21756 (N_21756,N_21556,N_21483);
or U21757 (N_21757,N_21463,N_21337);
xor U21758 (N_21758,N_21589,N_21439);
and U21759 (N_21759,N_21388,N_21336);
nand U21760 (N_21760,N_21358,N_21390);
nand U21761 (N_21761,N_21335,N_21470);
and U21762 (N_21762,N_21403,N_21503);
xnor U21763 (N_21763,N_21451,N_21446);
nand U21764 (N_21764,N_21445,N_21593);
nand U21765 (N_21765,N_21495,N_21355);
nand U21766 (N_21766,N_21326,N_21405);
or U21767 (N_21767,N_21570,N_21514);
xor U21768 (N_21768,N_21565,N_21406);
nand U21769 (N_21769,N_21516,N_21344);
or U21770 (N_21770,N_21387,N_21360);
nor U21771 (N_21771,N_21473,N_21492);
nand U21772 (N_21772,N_21425,N_21317);
nor U21773 (N_21773,N_21353,N_21364);
nand U21774 (N_21774,N_21445,N_21349);
nor U21775 (N_21775,N_21405,N_21544);
and U21776 (N_21776,N_21471,N_21301);
and U21777 (N_21777,N_21565,N_21429);
xnor U21778 (N_21778,N_21317,N_21429);
nand U21779 (N_21779,N_21569,N_21363);
nand U21780 (N_21780,N_21580,N_21569);
and U21781 (N_21781,N_21585,N_21339);
xnor U21782 (N_21782,N_21448,N_21355);
and U21783 (N_21783,N_21558,N_21410);
xor U21784 (N_21784,N_21590,N_21387);
nor U21785 (N_21785,N_21545,N_21469);
nor U21786 (N_21786,N_21564,N_21336);
and U21787 (N_21787,N_21592,N_21567);
nor U21788 (N_21788,N_21474,N_21590);
nor U21789 (N_21789,N_21489,N_21517);
nand U21790 (N_21790,N_21590,N_21456);
nor U21791 (N_21791,N_21576,N_21388);
nor U21792 (N_21792,N_21508,N_21589);
nand U21793 (N_21793,N_21466,N_21580);
nand U21794 (N_21794,N_21349,N_21355);
and U21795 (N_21795,N_21504,N_21342);
and U21796 (N_21796,N_21465,N_21542);
xnor U21797 (N_21797,N_21529,N_21365);
or U21798 (N_21798,N_21408,N_21419);
nor U21799 (N_21799,N_21451,N_21483);
or U21800 (N_21800,N_21582,N_21424);
nor U21801 (N_21801,N_21449,N_21324);
nand U21802 (N_21802,N_21324,N_21576);
xnor U21803 (N_21803,N_21491,N_21504);
xor U21804 (N_21804,N_21570,N_21311);
xnor U21805 (N_21805,N_21356,N_21316);
nor U21806 (N_21806,N_21599,N_21329);
xnor U21807 (N_21807,N_21409,N_21390);
and U21808 (N_21808,N_21327,N_21561);
nor U21809 (N_21809,N_21496,N_21321);
or U21810 (N_21810,N_21426,N_21368);
and U21811 (N_21811,N_21597,N_21303);
and U21812 (N_21812,N_21440,N_21441);
and U21813 (N_21813,N_21349,N_21557);
nand U21814 (N_21814,N_21345,N_21515);
and U21815 (N_21815,N_21534,N_21472);
nor U21816 (N_21816,N_21417,N_21332);
and U21817 (N_21817,N_21489,N_21582);
or U21818 (N_21818,N_21519,N_21395);
xnor U21819 (N_21819,N_21557,N_21393);
and U21820 (N_21820,N_21420,N_21321);
or U21821 (N_21821,N_21426,N_21417);
xnor U21822 (N_21822,N_21305,N_21489);
nor U21823 (N_21823,N_21516,N_21433);
or U21824 (N_21824,N_21438,N_21449);
xnor U21825 (N_21825,N_21588,N_21542);
nor U21826 (N_21826,N_21402,N_21332);
nand U21827 (N_21827,N_21522,N_21308);
nor U21828 (N_21828,N_21457,N_21578);
nor U21829 (N_21829,N_21552,N_21568);
or U21830 (N_21830,N_21419,N_21345);
and U21831 (N_21831,N_21498,N_21591);
nand U21832 (N_21832,N_21366,N_21437);
nand U21833 (N_21833,N_21511,N_21454);
or U21834 (N_21834,N_21355,N_21367);
and U21835 (N_21835,N_21527,N_21464);
nor U21836 (N_21836,N_21397,N_21370);
nand U21837 (N_21837,N_21324,N_21550);
nand U21838 (N_21838,N_21432,N_21364);
and U21839 (N_21839,N_21490,N_21576);
nor U21840 (N_21840,N_21399,N_21307);
or U21841 (N_21841,N_21331,N_21599);
nor U21842 (N_21842,N_21346,N_21307);
nor U21843 (N_21843,N_21458,N_21377);
xor U21844 (N_21844,N_21410,N_21505);
nor U21845 (N_21845,N_21307,N_21488);
nor U21846 (N_21846,N_21484,N_21411);
xor U21847 (N_21847,N_21339,N_21576);
nor U21848 (N_21848,N_21394,N_21594);
nand U21849 (N_21849,N_21486,N_21577);
nor U21850 (N_21850,N_21327,N_21508);
xnor U21851 (N_21851,N_21325,N_21424);
nor U21852 (N_21852,N_21450,N_21309);
xnor U21853 (N_21853,N_21530,N_21451);
or U21854 (N_21854,N_21516,N_21412);
and U21855 (N_21855,N_21416,N_21400);
or U21856 (N_21856,N_21408,N_21492);
and U21857 (N_21857,N_21463,N_21343);
nor U21858 (N_21858,N_21340,N_21532);
nand U21859 (N_21859,N_21484,N_21424);
nor U21860 (N_21860,N_21593,N_21494);
or U21861 (N_21861,N_21581,N_21523);
or U21862 (N_21862,N_21449,N_21510);
xnor U21863 (N_21863,N_21385,N_21391);
or U21864 (N_21864,N_21319,N_21489);
nand U21865 (N_21865,N_21550,N_21394);
nand U21866 (N_21866,N_21321,N_21345);
or U21867 (N_21867,N_21322,N_21474);
nand U21868 (N_21868,N_21475,N_21328);
and U21869 (N_21869,N_21507,N_21536);
xnor U21870 (N_21870,N_21394,N_21333);
or U21871 (N_21871,N_21536,N_21554);
and U21872 (N_21872,N_21304,N_21452);
or U21873 (N_21873,N_21540,N_21514);
or U21874 (N_21874,N_21492,N_21439);
or U21875 (N_21875,N_21447,N_21479);
nand U21876 (N_21876,N_21345,N_21499);
or U21877 (N_21877,N_21487,N_21503);
xnor U21878 (N_21878,N_21456,N_21526);
nand U21879 (N_21879,N_21406,N_21472);
or U21880 (N_21880,N_21404,N_21569);
xnor U21881 (N_21881,N_21436,N_21478);
xnor U21882 (N_21882,N_21449,N_21506);
nand U21883 (N_21883,N_21574,N_21587);
nand U21884 (N_21884,N_21403,N_21435);
nand U21885 (N_21885,N_21564,N_21545);
xor U21886 (N_21886,N_21413,N_21379);
xor U21887 (N_21887,N_21444,N_21599);
xnor U21888 (N_21888,N_21558,N_21477);
and U21889 (N_21889,N_21548,N_21593);
and U21890 (N_21890,N_21593,N_21481);
or U21891 (N_21891,N_21361,N_21529);
nor U21892 (N_21892,N_21413,N_21373);
nor U21893 (N_21893,N_21302,N_21471);
nand U21894 (N_21894,N_21450,N_21470);
nor U21895 (N_21895,N_21537,N_21425);
nor U21896 (N_21896,N_21552,N_21381);
and U21897 (N_21897,N_21565,N_21443);
or U21898 (N_21898,N_21525,N_21415);
or U21899 (N_21899,N_21438,N_21531);
or U21900 (N_21900,N_21695,N_21625);
and U21901 (N_21901,N_21634,N_21828);
or U21902 (N_21902,N_21795,N_21839);
xnor U21903 (N_21903,N_21787,N_21838);
or U21904 (N_21904,N_21774,N_21629);
nor U21905 (N_21905,N_21706,N_21790);
xnor U21906 (N_21906,N_21678,N_21740);
nor U21907 (N_21907,N_21844,N_21652);
and U21908 (N_21908,N_21733,N_21889);
nand U21909 (N_21909,N_21679,N_21748);
xor U21910 (N_21910,N_21776,N_21744);
xnor U21911 (N_21911,N_21779,N_21618);
or U21912 (N_21912,N_21653,N_21707);
nor U21913 (N_21913,N_21681,N_21785);
nor U21914 (N_21914,N_21723,N_21871);
or U21915 (N_21915,N_21860,N_21818);
and U21916 (N_21916,N_21743,N_21645);
or U21917 (N_21917,N_21633,N_21700);
or U21918 (N_21918,N_21879,N_21736);
and U21919 (N_21919,N_21869,N_21865);
or U21920 (N_21920,N_21713,N_21853);
nor U21921 (N_21921,N_21686,N_21682);
xnor U21922 (N_21922,N_21665,N_21848);
and U21923 (N_21923,N_21797,N_21624);
or U21924 (N_21924,N_21655,N_21701);
xor U21925 (N_21925,N_21773,N_21676);
xnor U21926 (N_21926,N_21843,N_21887);
nand U21927 (N_21927,N_21882,N_21711);
and U21928 (N_21928,N_21780,N_21886);
nor U21929 (N_21929,N_21670,N_21883);
nor U21930 (N_21930,N_21662,N_21609);
or U21931 (N_21931,N_21636,N_21750);
and U21932 (N_21932,N_21829,N_21866);
and U21933 (N_21933,N_21824,N_21666);
nor U21934 (N_21934,N_21896,N_21661);
nand U21935 (N_21935,N_21817,N_21643);
or U21936 (N_21936,N_21672,N_21697);
and U21937 (N_21937,N_21635,N_21751);
or U21938 (N_21938,N_21893,N_21877);
or U21939 (N_21939,N_21745,N_21777);
xor U21940 (N_21940,N_21832,N_21669);
nor U21941 (N_21941,N_21644,N_21607);
nand U21942 (N_21942,N_21814,N_21830);
or U21943 (N_21943,N_21720,N_21771);
nor U21944 (N_21944,N_21630,N_21621);
and U21945 (N_21945,N_21891,N_21764);
nand U21946 (N_21946,N_21845,N_21606);
nand U21947 (N_21947,N_21738,N_21874);
or U21948 (N_21948,N_21759,N_21673);
nor U21949 (N_21949,N_21762,N_21802);
xor U21950 (N_21950,N_21619,N_21820);
nand U21951 (N_21951,N_21731,N_21693);
or U21952 (N_21952,N_21873,N_21812);
nand U21953 (N_21953,N_21852,N_21858);
nand U21954 (N_21954,N_21854,N_21729);
nand U21955 (N_21955,N_21794,N_21641);
and U21956 (N_21956,N_21716,N_21760);
or U21957 (N_21957,N_21604,N_21819);
or U21958 (N_21958,N_21647,N_21677);
nand U21959 (N_21959,N_21810,N_21847);
nor U21960 (N_21960,N_21737,N_21602);
xnor U21961 (N_21961,N_21851,N_21868);
nor U21962 (N_21962,N_21660,N_21876);
nor U21963 (N_21963,N_21742,N_21793);
nand U21964 (N_21964,N_21698,N_21657);
and U21965 (N_21965,N_21768,N_21714);
nand U21966 (N_21966,N_21754,N_21692);
or U21967 (N_21967,N_21833,N_21863);
and U21968 (N_21968,N_21849,N_21765);
nor U21969 (N_21969,N_21658,N_21724);
xor U21970 (N_21970,N_21781,N_21649);
and U21971 (N_21971,N_21667,N_21735);
xor U21972 (N_21972,N_21642,N_21664);
xnor U21973 (N_21973,N_21640,N_21622);
nor U21974 (N_21974,N_21837,N_21864);
nor U21975 (N_21975,N_21675,N_21628);
xor U21976 (N_21976,N_21718,N_21668);
or U21977 (N_21977,N_21811,N_21709);
or U21978 (N_21978,N_21603,N_21763);
or U21979 (N_21979,N_21778,N_21694);
and U21980 (N_21980,N_21796,N_21739);
nor U21981 (N_21981,N_21827,N_21789);
nand U21982 (N_21982,N_21687,N_21788);
and U21983 (N_21983,N_21825,N_21704);
and U21984 (N_21984,N_21826,N_21758);
or U21985 (N_21985,N_21783,N_21722);
and U21986 (N_21986,N_21834,N_21637);
xnor U21987 (N_21987,N_21683,N_21798);
xnor U21988 (N_21988,N_21836,N_21631);
nand U21989 (N_21989,N_21699,N_21861);
xor U21990 (N_21990,N_21813,N_21888);
nand U21991 (N_21991,N_21616,N_21884);
and U21992 (N_21992,N_21890,N_21684);
xor U21993 (N_21993,N_21855,N_21749);
and U21994 (N_21994,N_21856,N_21689);
xor U21995 (N_21995,N_21772,N_21757);
nor U21996 (N_21996,N_21808,N_21805);
xnor U21997 (N_21997,N_21804,N_21691);
nand U21998 (N_21998,N_21842,N_21638);
xnor U21999 (N_21999,N_21835,N_21680);
nand U22000 (N_22000,N_21807,N_21727);
or U22001 (N_22001,N_21755,N_21775);
nand U22002 (N_22002,N_21894,N_21867);
nor U22003 (N_22003,N_21620,N_21734);
and U22004 (N_22004,N_21786,N_21726);
and U22005 (N_22005,N_21850,N_21746);
and U22006 (N_22006,N_21715,N_21690);
nand U22007 (N_22007,N_21761,N_21791);
nor U22008 (N_22008,N_21656,N_21895);
xnor U22009 (N_22009,N_21840,N_21717);
and U22010 (N_22010,N_21702,N_21623);
nor U22011 (N_22011,N_21752,N_21632);
and U22012 (N_22012,N_21605,N_21610);
and U22013 (N_22013,N_21741,N_21612);
nor U22014 (N_22014,N_21872,N_21823);
and U22015 (N_22015,N_21859,N_21870);
or U22016 (N_22016,N_21654,N_21892);
and U22017 (N_22017,N_21784,N_21721);
nor U22018 (N_22018,N_21608,N_21857);
xor U22019 (N_22019,N_21725,N_21816);
nor U22020 (N_22020,N_21615,N_21626);
nand U22021 (N_22021,N_21862,N_21747);
nand U22022 (N_22022,N_21617,N_21769);
nor U22023 (N_22023,N_21821,N_21792);
nand U22024 (N_22024,N_21809,N_21611);
and U22025 (N_22025,N_21897,N_21732);
and U22026 (N_22026,N_21803,N_21822);
and U22027 (N_22027,N_21627,N_21756);
xor U22028 (N_22028,N_21648,N_21898);
nand U22029 (N_22029,N_21688,N_21730);
or U22030 (N_22030,N_21650,N_21696);
xor U22031 (N_22031,N_21646,N_21601);
xnor U22032 (N_22032,N_21600,N_21831);
nand U22033 (N_22033,N_21770,N_21880);
nand U22034 (N_22034,N_21767,N_21878);
nand U22035 (N_22035,N_21671,N_21881);
nand U22036 (N_22036,N_21846,N_21728);
and U22037 (N_22037,N_21815,N_21719);
xnor U22038 (N_22038,N_21766,N_21801);
nor U22039 (N_22039,N_21710,N_21708);
and U22040 (N_22040,N_21703,N_21651);
nor U22041 (N_22041,N_21614,N_21885);
nand U22042 (N_22042,N_21685,N_21705);
xor U22043 (N_22043,N_21753,N_21712);
xor U22044 (N_22044,N_21613,N_21899);
or U22045 (N_22045,N_21800,N_21806);
or U22046 (N_22046,N_21841,N_21875);
and U22047 (N_22047,N_21782,N_21659);
nand U22048 (N_22048,N_21639,N_21799);
xor U22049 (N_22049,N_21674,N_21663);
xnor U22050 (N_22050,N_21623,N_21767);
nor U22051 (N_22051,N_21888,N_21848);
or U22052 (N_22052,N_21860,N_21838);
nor U22053 (N_22053,N_21877,N_21638);
and U22054 (N_22054,N_21740,N_21889);
nand U22055 (N_22055,N_21682,N_21769);
or U22056 (N_22056,N_21742,N_21746);
nor U22057 (N_22057,N_21863,N_21658);
and U22058 (N_22058,N_21824,N_21605);
xor U22059 (N_22059,N_21798,N_21885);
and U22060 (N_22060,N_21783,N_21683);
and U22061 (N_22061,N_21777,N_21894);
nand U22062 (N_22062,N_21822,N_21838);
nand U22063 (N_22063,N_21693,N_21838);
or U22064 (N_22064,N_21668,N_21711);
xnor U22065 (N_22065,N_21746,N_21790);
xnor U22066 (N_22066,N_21876,N_21881);
nor U22067 (N_22067,N_21863,N_21621);
xnor U22068 (N_22068,N_21864,N_21789);
nor U22069 (N_22069,N_21782,N_21654);
nand U22070 (N_22070,N_21839,N_21895);
nand U22071 (N_22071,N_21844,N_21775);
nor U22072 (N_22072,N_21796,N_21611);
or U22073 (N_22073,N_21875,N_21601);
or U22074 (N_22074,N_21770,N_21857);
nor U22075 (N_22075,N_21824,N_21748);
and U22076 (N_22076,N_21604,N_21719);
nand U22077 (N_22077,N_21709,N_21694);
nor U22078 (N_22078,N_21736,N_21848);
nor U22079 (N_22079,N_21720,N_21850);
nor U22080 (N_22080,N_21701,N_21827);
xnor U22081 (N_22081,N_21725,N_21639);
nor U22082 (N_22082,N_21743,N_21884);
xor U22083 (N_22083,N_21766,N_21836);
or U22084 (N_22084,N_21862,N_21701);
or U22085 (N_22085,N_21827,N_21745);
xnor U22086 (N_22086,N_21765,N_21616);
nand U22087 (N_22087,N_21767,N_21888);
and U22088 (N_22088,N_21668,N_21832);
nor U22089 (N_22089,N_21738,N_21623);
xor U22090 (N_22090,N_21896,N_21854);
nand U22091 (N_22091,N_21811,N_21790);
or U22092 (N_22092,N_21801,N_21805);
nand U22093 (N_22093,N_21844,N_21751);
nor U22094 (N_22094,N_21849,N_21846);
or U22095 (N_22095,N_21772,N_21668);
xnor U22096 (N_22096,N_21670,N_21780);
and U22097 (N_22097,N_21697,N_21837);
nor U22098 (N_22098,N_21869,N_21778);
xnor U22099 (N_22099,N_21600,N_21815);
and U22100 (N_22100,N_21810,N_21688);
nand U22101 (N_22101,N_21643,N_21792);
or U22102 (N_22102,N_21602,N_21654);
xnor U22103 (N_22103,N_21854,N_21783);
nor U22104 (N_22104,N_21806,N_21895);
xnor U22105 (N_22105,N_21885,N_21839);
nand U22106 (N_22106,N_21638,N_21616);
nand U22107 (N_22107,N_21877,N_21661);
and U22108 (N_22108,N_21749,N_21671);
nand U22109 (N_22109,N_21815,N_21656);
nand U22110 (N_22110,N_21844,N_21834);
nor U22111 (N_22111,N_21620,N_21853);
or U22112 (N_22112,N_21785,N_21694);
and U22113 (N_22113,N_21640,N_21849);
and U22114 (N_22114,N_21680,N_21839);
xor U22115 (N_22115,N_21836,N_21667);
nor U22116 (N_22116,N_21806,N_21860);
or U22117 (N_22117,N_21852,N_21785);
nand U22118 (N_22118,N_21798,N_21790);
or U22119 (N_22119,N_21859,N_21866);
nor U22120 (N_22120,N_21601,N_21884);
nor U22121 (N_22121,N_21686,N_21873);
or U22122 (N_22122,N_21622,N_21652);
and U22123 (N_22123,N_21689,N_21649);
nand U22124 (N_22124,N_21762,N_21798);
or U22125 (N_22125,N_21833,N_21736);
and U22126 (N_22126,N_21765,N_21610);
or U22127 (N_22127,N_21835,N_21693);
and U22128 (N_22128,N_21831,N_21819);
xor U22129 (N_22129,N_21736,N_21758);
nand U22130 (N_22130,N_21812,N_21806);
nor U22131 (N_22131,N_21875,N_21709);
nor U22132 (N_22132,N_21820,N_21782);
or U22133 (N_22133,N_21746,N_21733);
nor U22134 (N_22134,N_21662,N_21889);
xor U22135 (N_22135,N_21783,N_21681);
xnor U22136 (N_22136,N_21726,N_21869);
nand U22137 (N_22137,N_21708,N_21882);
nor U22138 (N_22138,N_21671,N_21890);
or U22139 (N_22139,N_21618,N_21634);
or U22140 (N_22140,N_21753,N_21889);
or U22141 (N_22141,N_21820,N_21664);
xnor U22142 (N_22142,N_21844,N_21856);
xnor U22143 (N_22143,N_21856,N_21624);
and U22144 (N_22144,N_21823,N_21663);
nand U22145 (N_22145,N_21883,N_21609);
and U22146 (N_22146,N_21630,N_21793);
xnor U22147 (N_22147,N_21622,N_21890);
and U22148 (N_22148,N_21765,N_21865);
or U22149 (N_22149,N_21870,N_21602);
nand U22150 (N_22150,N_21710,N_21824);
xor U22151 (N_22151,N_21773,N_21810);
xnor U22152 (N_22152,N_21857,N_21895);
nand U22153 (N_22153,N_21881,N_21833);
xnor U22154 (N_22154,N_21641,N_21721);
nor U22155 (N_22155,N_21805,N_21867);
xnor U22156 (N_22156,N_21704,N_21864);
xnor U22157 (N_22157,N_21778,N_21754);
or U22158 (N_22158,N_21720,N_21621);
nor U22159 (N_22159,N_21642,N_21890);
and U22160 (N_22160,N_21662,N_21852);
and U22161 (N_22161,N_21821,N_21842);
nor U22162 (N_22162,N_21792,N_21896);
xnor U22163 (N_22163,N_21859,N_21783);
xor U22164 (N_22164,N_21671,N_21648);
and U22165 (N_22165,N_21734,N_21725);
and U22166 (N_22166,N_21769,N_21832);
and U22167 (N_22167,N_21697,N_21891);
nand U22168 (N_22168,N_21621,N_21884);
nor U22169 (N_22169,N_21674,N_21614);
or U22170 (N_22170,N_21713,N_21635);
xor U22171 (N_22171,N_21798,N_21816);
or U22172 (N_22172,N_21699,N_21715);
xnor U22173 (N_22173,N_21875,N_21702);
xor U22174 (N_22174,N_21740,N_21716);
nand U22175 (N_22175,N_21840,N_21716);
xor U22176 (N_22176,N_21774,N_21894);
xor U22177 (N_22177,N_21728,N_21761);
or U22178 (N_22178,N_21851,N_21629);
and U22179 (N_22179,N_21763,N_21715);
or U22180 (N_22180,N_21619,N_21741);
nand U22181 (N_22181,N_21624,N_21623);
or U22182 (N_22182,N_21811,N_21600);
nand U22183 (N_22183,N_21630,N_21693);
nor U22184 (N_22184,N_21826,N_21843);
or U22185 (N_22185,N_21791,N_21781);
nor U22186 (N_22186,N_21680,N_21669);
or U22187 (N_22187,N_21828,N_21636);
nor U22188 (N_22188,N_21668,N_21815);
or U22189 (N_22189,N_21790,N_21755);
or U22190 (N_22190,N_21880,N_21745);
xor U22191 (N_22191,N_21812,N_21843);
or U22192 (N_22192,N_21684,N_21750);
nand U22193 (N_22193,N_21679,N_21757);
xnor U22194 (N_22194,N_21779,N_21793);
xnor U22195 (N_22195,N_21739,N_21661);
and U22196 (N_22196,N_21813,N_21895);
nor U22197 (N_22197,N_21759,N_21786);
or U22198 (N_22198,N_21813,N_21751);
nor U22199 (N_22199,N_21886,N_21758);
nand U22200 (N_22200,N_22109,N_22070);
and U22201 (N_22201,N_22064,N_22069);
nand U22202 (N_22202,N_22013,N_21917);
or U22203 (N_22203,N_21938,N_22143);
nor U22204 (N_22204,N_22006,N_22009);
and U22205 (N_22205,N_22146,N_22130);
nand U22206 (N_22206,N_22191,N_21986);
xnor U22207 (N_22207,N_22063,N_22118);
nor U22208 (N_22208,N_21948,N_22124);
or U22209 (N_22209,N_21920,N_22022);
nand U22210 (N_22210,N_22010,N_22199);
and U22211 (N_22211,N_22040,N_22004);
nor U22212 (N_22212,N_21942,N_22189);
or U22213 (N_22213,N_22145,N_22086);
xor U22214 (N_22214,N_22018,N_22148);
xor U22215 (N_22215,N_22133,N_22157);
nand U22216 (N_22216,N_22046,N_22147);
or U22217 (N_22217,N_22101,N_22182);
nand U22218 (N_22218,N_22042,N_22067);
xnor U22219 (N_22219,N_22080,N_21907);
nor U22220 (N_22220,N_22075,N_22115);
and U22221 (N_22221,N_22072,N_21963);
nand U22222 (N_22222,N_22048,N_22073);
xor U22223 (N_22223,N_22151,N_21930);
xnor U22224 (N_22224,N_22102,N_22071);
or U22225 (N_22225,N_21919,N_22176);
nor U22226 (N_22226,N_22029,N_22195);
nor U22227 (N_22227,N_22056,N_22052);
and U22228 (N_22228,N_21925,N_21987);
xor U22229 (N_22229,N_21915,N_21961);
nor U22230 (N_22230,N_22152,N_21971);
nand U22231 (N_22231,N_22186,N_21947);
nor U22232 (N_22232,N_22132,N_22104);
or U22233 (N_22233,N_22091,N_22081);
or U22234 (N_22234,N_22110,N_22055);
and U22235 (N_22235,N_22165,N_22164);
or U22236 (N_22236,N_21967,N_22078);
and U22237 (N_22237,N_21937,N_21982);
xor U22238 (N_22238,N_22139,N_22028);
or U22239 (N_22239,N_22015,N_22066);
nand U22240 (N_22240,N_22196,N_22161);
nand U22241 (N_22241,N_22194,N_22041);
or U22242 (N_22242,N_22065,N_22012);
and U22243 (N_22243,N_21914,N_22134);
nor U22244 (N_22244,N_22023,N_22051);
or U22245 (N_22245,N_22011,N_21927);
nand U22246 (N_22246,N_21902,N_22180);
nor U22247 (N_22247,N_21988,N_21904);
nand U22248 (N_22248,N_22000,N_21905);
xor U22249 (N_22249,N_22008,N_22007);
nand U22250 (N_22250,N_21989,N_22096);
and U22251 (N_22251,N_22149,N_22098);
nand U22252 (N_22252,N_22049,N_22021);
nand U22253 (N_22253,N_21977,N_22127);
or U22254 (N_22254,N_22083,N_22184);
or U22255 (N_22255,N_22061,N_21949);
nor U22256 (N_22256,N_22137,N_21936);
xor U22257 (N_22257,N_22126,N_21995);
or U22258 (N_22258,N_21954,N_22154);
xnor U22259 (N_22259,N_22033,N_22177);
nand U22260 (N_22260,N_22076,N_22035);
and U22261 (N_22261,N_22153,N_22087);
and U22262 (N_22262,N_22045,N_21908);
nand U22263 (N_22263,N_22128,N_21952);
nand U22264 (N_22264,N_22100,N_22155);
nor U22265 (N_22265,N_21958,N_21990);
nand U22266 (N_22266,N_21912,N_21901);
nand U22267 (N_22267,N_22060,N_22020);
and U22268 (N_22268,N_21955,N_22172);
xnor U22269 (N_22269,N_22187,N_21976);
xor U22270 (N_22270,N_22003,N_21972);
nand U22271 (N_22271,N_21932,N_22197);
and U22272 (N_22272,N_22125,N_22039);
nor U22273 (N_22273,N_22173,N_22112);
xor U22274 (N_22274,N_21910,N_21994);
and U22275 (N_22275,N_22043,N_21964);
nor U22276 (N_22276,N_21940,N_21953);
nand U22277 (N_22277,N_22183,N_22097);
or U22278 (N_22278,N_21943,N_21965);
nand U22279 (N_22279,N_22036,N_21926);
and U22280 (N_22280,N_22142,N_21993);
and U22281 (N_22281,N_21968,N_22068);
or U22282 (N_22282,N_21956,N_22121);
nand U22283 (N_22283,N_21911,N_22082);
nor U22284 (N_22284,N_21962,N_22108);
nand U22285 (N_22285,N_21959,N_21903);
and U22286 (N_22286,N_22119,N_22037);
or U22287 (N_22287,N_22167,N_22141);
nor U22288 (N_22288,N_22158,N_21983);
nor U22289 (N_22289,N_22111,N_22129);
xor U22290 (N_22290,N_21960,N_22014);
xor U22291 (N_22291,N_22156,N_22090);
nor U22292 (N_22292,N_22001,N_22074);
nor U22293 (N_22293,N_22131,N_22166);
nand U22294 (N_22294,N_22088,N_22024);
xor U22295 (N_22295,N_22106,N_22193);
nor U22296 (N_22296,N_21973,N_22058);
nor U22297 (N_22297,N_22026,N_21999);
or U22298 (N_22298,N_21991,N_21997);
nor U22299 (N_22299,N_21998,N_21945);
or U22300 (N_22300,N_22034,N_21941);
and U22301 (N_22301,N_22144,N_21928);
or U22302 (N_22302,N_22027,N_21946);
and U22303 (N_22303,N_22175,N_21985);
xnor U22304 (N_22304,N_21979,N_22114);
nor U22305 (N_22305,N_22038,N_22059);
and U22306 (N_22306,N_21980,N_22168);
nand U22307 (N_22307,N_22092,N_22116);
and U22308 (N_22308,N_21974,N_21934);
xnor U22309 (N_22309,N_22062,N_21921);
and U22310 (N_22310,N_22084,N_21984);
nor U22311 (N_22311,N_21957,N_22094);
nor U22312 (N_22312,N_22016,N_22017);
nor U22313 (N_22313,N_22050,N_21923);
and U22314 (N_22314,N_22077,N_21900);
or U22315 (N_22315,N_22136,N_21933);
nand U22316 (N_22316,N_22047,N_22135);
nand U22317 (N_22317,N_21996,N_21913);
nand U22318 (N_22318,N_22162,N_22002);
nand U22319 (N_22319,N_22179,N_22120);
nand U22320 (N_22320,N_22181,N_22169);
and U22321 (N_22321,N_22160,N_21939);
nand U22322 (N_22322,N_22107,N_22085);
and U22323 (N_22323,N_22053,N_22188);
nor U22324 (N_22324,N_21992,N_22190);
nor U22325 (N_22325,N_22025,N_22099);
and U22326 (N_22326,N_22044,N_22095);
xnor U22327 (N_22327,N_22103,N_22089);
or U22328 (N_22328,N_21906,N_21924);
nor U22329 (N_22329,N_22150,N_21966);
xor U22330 (N_22330,N_22117,N_22032);
or U22331 (N_22331,N_22079,N_21978);
or U22332 (N_22332,N_21981,N_21918);
nand U22333 (N_22333,N_21970,N_21951);
nand U22334 (N_22334,N_22113,N_22178);
or U22335 (N_22335,N_21916,N_22174);
and U22336 (N_22336,N_22122,N_21950);
nor U22337 (N_22337,N_22057,N_21931);
and U22338 (N_22338,N_21922,N_22123);
xnor U22339 (N_22339,N_22054,N_22105);
nor U22340 (N_22340,N_22192,N_22093);
nand U22341 (N_22341,N_21975,N_22198);
xor U22342 (N_22342,N_21909,N_22170);
or U22343 (N_22343,N_22019,N_21944);
and U22344 (N_22344,N_22031,N_22140);
and U22345 (N_22345,N_21929,N_22163);
nand U22346 (N_22346,N_22171,N_22005);
xor U22347 (N_22347,N_22030,N_22159);
nand U22348 (N_22348,N_21969,N_21935);
nand U22349 (N_22349,N_22185,N_22138);
xor U22350 (N_22350,N_21994,N_22196);
and U22351 (N_22351,N_21981,N_22154);
and U22352 (N_22352,N_21908,N_21981);
or U22353 (N_22353,N_22071,N_22045);
and U22354 (N_22354,N_22101,N_22073);
nand U22355 (N_22355,N_21940,N_22126);
nand U22356 (N_22356,N_21909,N_22075);
and U22357 (N_22357,N_21948,N_21957);
xor U22358 (N_22358,N_22142,N_22083);
nor U22359 (N_22359,N_22155,N_21996);
or U22360 (N_22360,N_21943,N_21915);
xor U22361 (N_22361,N_22100,N_22071);
nor U22362 (N_22362,N_21958,N_21921);
nand U22363 (N_22363,N_21940,N_22078);
xor U22364 (N_22364,N_22139,N_22041);
nor U22365 (N_22365,N_22051,N_22017);
nand U22366 (N_22366,N_22015,N_22044);
or U22367 (N_22367,N_22036,N_21984);
xnor U22368 (N_22368,N_22033,N_22116);
xnor U22369 (N_22369,N_21983,N_21917);
nor U22370 (N_22370,N_22188,N_22164);
xor U22371 (N_22371,N_21986,N_22063);
or U22372 (N_22372,N_22114,N_22059);
nor U22373 (N_22373,N_22062,N_21910);
xor U22374 (N_22374,N_22188,N_22079);
or U22375 (N_22375,N_21955,N_21956);
and U22376 (N_22376,N_22022,N_22186);
nand U22377 (N_22377,N_22151,N_22144);
xnor U22378 (N_22378,N_21980,N_21930);
nor U22379 (N_22379,N_22138,N_22027);
xnor U22380 (N_22380,N_21934,N_21968);
nand U22381 (N_22381,N_21931,N_21907);
or U22382 (N_22382,N_22022,N_22051);
nor U22383 (N_22383,N_22152,N_21995);
nand U22384 (N_22384,N_22054,N_22150);
and U22385 (N_22385,N_22157,N_21932);
and U22386 (N_22386,N_22189,N_21928);
and U22387 (N_22387,N_22123,N_21990);
xor U22388 (N_22388,N_21988,N_21960);
nand U22389 (N_22389,N_22163,N_22091);
or U22390 (N_22390,N_21961,N_22160);
or U22391 (N_22391,N_22106,N_21936);
and U22392 (N_22392,N_22046,N_22178);
nand U22393 (N_22393,N_22051,N_21954);
xor U22394 (N_22394,N_22149,N_22143);
xor U22395 (N_22395,N_21929,N_22124);
or U22396 (N_22396,N_22126,N_21960);
nor U22397 (N_22397,N_22061,N_21959);
or U22398 (N_22398,N_21926,N_21948);
or U22399 (N_22399,N_21994,N_21927);
nor U22400 (N_22400,N_22179,N_22106);
nor U22401 (N_22401,N_22127,N_22138);
nand U22402 (N_22402,N_22093,N_22087);
nor U22403 (N_22403,N_22013,N_21931);
and U22404 (N_22404,N_22060,N_22016);
nor U22405 (N_22405,N_21925,N_21917);
nor U22406 (N_22406,N_22141,N_21959);
nand U22407 (N_22407,N_21964,N_22092);
and U22408 (N_22408,N_22035,N_22053);
xor U22409 (N_22409,N_21914,N_22163);
xor U22410 (N_22410,N_21961,N_22171);
or U22411 (N_22411,N_22126,N_22015);
nor U22412 (N_22412,N_21933,N_21968);
xnor U22413 (N_22413,N_22005,N_22031);
nor U22414 (N_22414,N_22108,N_22141);
and U22415 (N_22415,N_22146,N_22064);
and U22416 (N_22416,N_21958,N_22130);
nand U22417 (N_22417,N_22053,N_21980);
xor U22418 (N_22418,N_21995,N_22180);
xnor U22419 (N_22419,N_22060,N_21990);
nor U22420 (N_22420,N_22001,N_22125);
nor U22421 (N_22421,N_22122,N_22071);
and U22422 (N_22422,N_22112,N_21985);
xor U22423 (N_22423,N_22176,N_22041);
nand U22424 (N_22424,N_22173,N_21972);
and U22425 (N_22425,N_22062,N_21905);
nand U22426 (N_22426,N_22107,N_22020);
or U22427 (N_22427,N_22105,N_22153);
xnor U22428 (N_22428,N_22050,N_22039);
nor U22429 (N_22429,N_22085,N_22150);
nor U22430 (N_22430,N_22097,N_22156);
and U22431 (N_22431,N_22082,N_22145);
xnor U22432 (N_22432,N_22013,N_22009);
nor U22433 (N_22433,N_22006,N_21901);
nor U22434 (N_22434,N_22088,N_22081);
nand U22435 (N_22435,N_22189,N_22197);
nor U22436 (N_22436,N_22011,N_22137);
nand U22437 (N_22437,N_22165,N_22026);
nand U22438 (N_22438,N_21944,N_21914);
nor U22439 (N_22439,N_22105,N_22172);
xnor U22440 (N_22440,N_22183,N_21958);
nor U22441 (N_22441,N_22136,N_22154);
or U22442 (N_22442,N_22071,N_21937);
nor U22443 (N_22443,N_22079,N_22197);
nor U22444 (N_22444,N_22058,N_21953);
or U22445 (N_22445,N_22046,N_22027);
nor U22446 (N_22446,N_22033,N_22010);
nand U22447 (N_22447,N_21975,N_22166);
and U22448 (N_22448,N_22041,N_22048);
nand U22449 (N_22449,N_22118,N_22081);
nand U22450 (N_22450,N_22003,N_22148);
or U22451 (N_22451,N_22082,N_22177);
nor U22452 (N_22452,N_21955,N_21987);
nand U22453 (N_22453,N_22159,N_22146);
nand U22454 (N_22454,N_22090,N_21966);
nand U22455 (N_22455,N_22084,N_22097);
nor U22456 (N_22456,N_22187,N_22014);
nand U22457 (N_22457,N_22029,N_22111);
or U22458 (N_22458,N_22018,N_22172);
nand U22459 (N_22459,N_22088,N_21925);
and U22460 (N_22460,N_22029,N_22079);
or U22461 (N_22461,N_22126,N_21958);
nand U22462 (N_22462,N_22002,N_22190);
nand U22463 (N_22463,N_22108,N_22029);
xnor U22464 (N_22464,N_22069,N_22112);
nor U22465 (N_22465,N_21900,N_22171);
nand U22466 (N_22466,N_21980,N_22001);
nand U22467 (N_22467,N_22036,N_22034);
and U22468 (N_22468,N_22157,N_21901);
and U22469 (N_22469,N_22047,N_22087);
nand U22470 (N_22470,N_22132,N_22055);
or U22471 (N_22471,N_22157,N_22063);
nor U22472 (N_22472,N_21958,N_22152);
or U22473 (N_22473,N_22044,N_21909);
nand U22474 (N_22474,N_22007,N_22147);
nand U22475 (N_22475,N_22194,N_21971);
and U22476 (N_22476,N_22085,N_22177);
nor U22477 (N_22477,N_22129,N_21976);
or U22478 (N_22478,N_21961,N_21903);
xor U22479 (N_22479,N_22158,N_22033);
and U22480 (N_22480,N_22159,N_22132);
or U22481 (N_22481,N_21931,N_22111);
and U22482 (N_22482,N_22180,N_21975);
xnor U22483 (N_22483,N_21961,N_21941);
nor U22484 (N_22484,N_22088,N_21980);
or U22485 (N_22485,N_22194,N_22162);
and U22486 (N_22486,N_21947,N_21931);
nand U22487 (N_22487,N_22188,N_21932);
and U22488 (N_22488,N_22190,N_22112);
xnor U22489 (N_22489,N_22066,N_22011);
or U22490 (N_22490,N_21903,N_21986);
or U22491 (N_22491,N_21915,N_21908);
nor U22492 (N_22492,N_22043,N_22138);
or U22493 (N_22493,N_22068,N_22141);
or U22494 (N_22494,N_22006,N_21971);
xnor U22495 (N_22495,N_22136,N_22013);
xnor U22496 (N_22496,N_21921,N_22117);
xor U22497 (N_22497,N_22164,N_22150);
xor U22498 (N_22498,N_21933,N_22104);
nor U22499 (N_22499,N_22003,N_22021);
nor U22500 (N_22500,N_22442,N_22427);
xnor U22501 (N_22501,N_22489,N_22472);
nor U22502 (N_22502,N_22312,N_22470);
nor U22503 (N_22503,N_22492,N_22200);
or U22504 (N_22504,N_22202,N_22259);
and U22505 (N_22505,N_22416,N_22417);
or U22506 (N_22506,N_22475,N_22361);
and U22507 (N_22507,N_22347,N_22272);
xor U22508 (N_22508,N_22295,N_22222);
nand U22509 (N_22509,N_22438,N_22236);
and U22510 (N_22510,N_22443,N_22284);
xnor U22511 (N_22511,N_22223,N_22451);
or U22512 (N_22512,N_22363,N_22399);
nand U22513 (N_22513,N_22359,N_22478);
and U22514 (N_22514,N_22429,N_22233);
nor U22515 (N_22515,N_22425,N_22433);
nor U22516 (N_22516,N_22420,N_22206);
xor U22517 (N_22517,N_22299,N_22344);
or U22518 (N_22518,N_22238,N_22216);
or U22519 (N_22519,N_22217,N_22260);
xnor U22520 (N_22520,N_22471,N_22249);
xor U22521 (N_22521,N_22481,N_22356);
nor U22522 (N_22522,N_22257,N_22209);
nand U22523 (N_22523,N_22230,N_22211);
nor U22524 (N_22524,N_22483,N_22245);
nor U22525 (N_22525,N_22498,N_22331);
nand U22526 (N_22526,N_22456,N_22221);
or U22527 (N_22527,N_22403,N_22266);
nor U22528 (N_22528,N_22374,N_22410);
nand U22529 (N_22529,N_22204,N_22386);
or U22530 (N_22530,N_22353,N_22394);
or U22531 (N_22531,N_22212,N_22321);
nand U22532 (N_22532,N_22404,N_22400);
xnor U22533 (N_22533,N_22407,N_22460);
nand U22534 (N_22534,N_22298,N_22373);
nor U22535 (N_22535,N_22465,N_22474);
nor U22536 (N_22536,N_22307,N_22402);
or U22537 (N_22537,N_22301,N_22463);
nand U22538 (N_22538,N_22459,N_22235);
xor U22539 (N_22539,N_22302,N_22324);
and U22540 (N_22540,N_22305,N_22358);
or U22541 (N_22541,N_22285,N_22319);
nor U22542 (N_22542,N_22293,N_22248);
or U22543 (N_22543,N_22458,N_22300);
xnor U22544 (N_22544,N_22218,N_22452);
nand U22545 (N_22545,N_22335,N_22247);
nand U22546 (N_22546,N_22279,N_22468);
and U22547 (N_22547,N_22387,N_22303);
nor U22548 (N_22548,N_22390,N_22445);
and U22549 (N_22549,N_22213,N_22393);
xor U22550 (N_22550,N_22367,N_22219);
xnor U22551 (N_22551,N_22304,N_22328);
and U22552 (N_22552,N_22336,N_22326);
and U22553 (N_22553,N_22318,N_22224);
nand U22554 (N_22554,N_22381,N_22482);
nor U22555 (N_22555,N_22428,N_22294);
xnor U22556 (N_22556,N_22430,N_22265);
and U22557 (N_22557,N_22243,N_22447);
and U22558 (N_22558,N_22225,N_22497);
or U22559 (N_22559,N_22330,N_22395);
nand U22560 (N_22560,N_22286,N_22352);
nand U22561 (N_22561,N_22268,N_22412);
xor U22562 (N_22562,N_22466,N_22389);
nor U22563 (N_22563,N_22343,N_22431);
or U22564 (N_22564,N_22296,N_22480);
nand U22565 (N_22565,N_22411,N_22437);
or U22566 (N_22566,N_22435,N_22227);
xnor U22567 (N_22567,N_22271,N_22369);
xnor U22568 (N_22568,N_22306,N_22231);
nor U22569 (N_22569,N_22340,N_22383);
or U22570 (N_22570,N_22372,N_22364);
nand U22571 (N_22571,N_22276,N_22316);
and U22572 (N_22572,N_22337,N_22309);
or U22573 (N_22573,N_22270,N_22378);
nand U22574 (N_22574,N_22362,N_22229);
nor U22575 (N_22575,N_22280,N_22253);
nand U22576 (N_22576,N_22287,N_22487);
nand U22577 (N_22577,N_22205,N_22338);
and U22578 (N_22578,N_22333,N_22461);
nor U22579 (N_22579,N_22244,N_22291);
xnor U22580 (N_22580,N_22453,N_22365);
xnor U22581 (N_22581,N_22491,N_22308);
nand U22582 (N_22582,N_22485,N_22495);
nand U22583 (N_22583,N_22269,N_22457);
or U22584 (N_22584,N_22391,N_22220);
nor U22585 (N_22585,N_22440,N_22467);
xor U22586 (N_22586,N_22469,N_22486);
or U22587 (N_22587,N_22310,N_22346);
and U22588 (N_22588,N_22208,N_22366);
nor U22589 (N_22589,N_22449,N_22250);
nand U22590 (N_22590,N_22256,N_22292);
and U22591 (N_22591,N_22341,N_22329);
nand U22592 (N_22592,N_22436,N_22476);
nor U22593 (N_22593,N_22210,N_22494);
or U22594 (N_22594,N_22289,N_22255);
nand U22595 (N_22595,N_22332,N_22448);
xnor U22596 (N_22596,N_22251,N_22325);
or U22597 (N_22597,N_22370,N_22345);
nand U22598 (N_22598,N_22405,N_22488);
or U22599 (N_22599,N_22267,N_22264);
or U22600 (N_22600,N_22357,N_22464);
and U22601 (N_22601,N_22479,N_22368);
or U22602 (N_22602,N_22434,N_22377);
nand U22603 (N_22603,N_22297,N_22273);
or U22604 (N_22604,N_22314,N_22320);
and U22605 (N_22605,N_22462,N_22414);
xor U22606 (N_22606,N_22406,N_22484);
or U22607 (N_22607,N_22203,N_22288);
xnor U22608 (N_22608,N_22348,N_22254);
nor U22609 (N_22609,N_22422,N_22441);
and U22610 (N_22610,N_22385,N_22473);
xor U22611 (N_22611,N_22263,N_22283);
nor U22612 (N_22612,N_22376,N_22388);
nand U22613 (N_22613,N_22392,N_22351);
nand U22614 (N_22614,N_22281,N_22232);
nand U22615 (N_22615,N_22490,N_22432);
xnor U22616 (N_22616,N_22415,N_22382);
nor U22617 (N_22617,N_22496,N_22342);
nand U22618 (N_22618,N_22277,N_22282);
or U22619 (N_22619,N_22401,N_22242);
and U22620 (N_22620,N_22215,N_22252);
xor U22621 (N_22621,N_22424,N_22214);
nor U22622 (N_22622,N_22397,N_22290);
nor U22623 (N_22623,N_22234,N_22439);
nand U22624 (N_22624,N_22421,N_22207);
or U22625 (N_22625,N_22311,N_22262);
xnor U22626 (N_22626,N_22379,N_22313);
or U22627 (N_22627,N_22315,N_22454);
xnor U22628 (N_22628,N_22446,N_22246);
nor U22629 (N_22629,N_22275,N_22258);
nor U22630 (N_22630,N_22226,N_22354);
xnor U22631 (N_22631,N_22334,N_22261);
nor U22632 (N_22632,N_22493,N_22413);
nor U22633 (N_22633,N_22278,N_22239);
xor U22634 (N_22634,N_22323,N_22398);
and U22635 (N_22635,N_22499,N_22237);
or U22636 (N_22636,N_22419,N_22322);
nor U22637 (N_22637,N_22409,N_22418);
xor U22638 (N_22638,N_22444,N_22360);
and U22639 (N_22639,N_22423,N_22349);
nor U22640 (N_22640,N_22396,N_22455);
nor U22641 (N_22641,N_22375,N_22327);
nand U22642 (N_22642,N_22355,N_22408);
xor U22643 (N_22643,N_22241,N_22350);
nor U22644 (N_22644,N_22228,N_22317);
and U22645 (N_22645,N_22477,N_22450);
nand U22646 (N_22646,N_22240,N_22380);
and U22647 (N_22647,N_22201,N_22339);
nor U22648 (N_22648,N_22371,N_22426);
and U22649 (N_22649,N_22274,N_22384);
and U22650 (N_22650,N_22401,N_22233);
or U22651 (N_22651,N_22438,N_22259);
or U22652 (N_22652,N_22283,N_22348);
xnor U22653 (N_22653,N_22330,N_22205);
xnor U22654 (N_22654,N_22390,N_22264);
nor U22655 (N_22655,N_22397,N_22274);
nor U22656 (N_22656,N_22230,N_22460);
nand U22657 (N_22657,N_22252,N_22294);
and U22658 (N_22658,N_22436,N_22351);
xnor U22659 (N_22659,N_22253,N_22291);
nor U22660 (N_22660,N_22338,N_22237);
nor U22661 (N_22661,N_22498,N_22312);
or U22662 (N_22662,N_22421,N_22310);
nor U22663 (N_22663,N_22476,N_22344);
and U22664 (N_22664,N_22417,N_22204);
or U22665 (N_22665,N_22406,N_22214);
xnor U22666 (N_22666,N_22297,N_22405);
xor U22667 (N_22667,N_22309,N_22424);
and U22668 (N_22668,N_22231,N_22334);
or U22669 (N_22669,N_22433,N_22218);
and U22670 (N_22670,N_22467,N_22261);
and U22671 (N_22671,N_22235,N_22391);
nor U22672 (N_22672,N_22324,N_22212);
or U22673 (N_22673,N_22453,N_22330);
and U22674 (N_22674,N_22365,N_22410);
nor U22675 (N_22675,N_22356,N_22418);
or U22676 (N_22676,N_22293,N_22269);
or U22677 (N_22677,N_22484,N_22441);
nor U22678 (N_22678,N_22263,N_22210);
nor U22679 (N_22679,N_22386,N_22283);
nand U22680 (N_22680,N_22404,N_22407);
and U22681 (N_22681,N_22280,N_22353);
and U22682 (N_22682,N_22498,N_22375);
nand U22683 (N_22683,N_22337,N_22267);
and U22684 (N_22684,N_22254,N_22347);
and U22685 (N_22685,N_22277,N_22315);
nand U22686 (N_22686,N_22434,N_22361);
xor U22687 (N_22687,N_22246,N_22424);
xor U22688 (N_22688,N_22438,N_22436);
xor U22689 (N_22689,N_22227,N_22482);
xnor U22690 (N_22690,N_22232,N_22425);
or U22691 (N_22691,N_22388,N_22495);
nand U22692 (N_22692,N_22358,N_22215);
xnor U22693 (N_22693,N_22393,N_22246);
xor U22694 (N_22694,N_22367,N_22482);
nor U22695 (N_22695,N_22446,N_22372);
nand U22696 (N_22696,N_22214,N_22257);
nand U22697 (N_22697,N_22475,N_22205);
nand U22698 (N_22698,N_22270,N_22439);
and U22699 (N_22699,N_22394,N_22444);
nand U22700 (N_22700,N_22412,N_22362);
and U22701 (N_22701,N_22463,N_22443);
and U22702 (N_22702,N_22208,N_22446);
and U22703 (N_22703,N_22498,N_22421);
or U22704 (N_22704,N_22439,N_22488);
and U22705 (N_22705,N_22341,N_22439);
nand U22706 (N_22706,N_22337,N_22433);
or U22707 (N_22707,N_22468,N_22482);
and U22708 (N_22708,N_22396,N_22404);
nor U22709 (N_22709,N_22298,N_22369);
and U22710 (N_22710,N_22404,N_22430);
or U22711 (N_22711,N_22473,N_22327);
xor U22712 (N_22712,N_22450,N_22496);
or U22713 (N_22713,N_22497,N_22359);
nor U22714 (N_22714,N_22425,N_22253);
nor U22715 (N_22715,N_22259,N_22423);
nor U22716 (N_22716,N_22315,N_22298);
and U22717 (N_22717,N_22276,N_22470);
xnor U22718 (N_22718,N_22419,N_22467);
or U22719 (N_22719,N_22302,N_22387);
nand U22720 (N_22720,N_22444,N_22470);
or U22721 (N_22721,N_22216,N_22449);
and U22722 (N_22722,N_22315,N_22409);
xor U22723 (N_22723,N_22223,N_22368);
nor U22724 (N_22724,N_22305,N_22421);
nor U22725 (N_22725,N_22394,N_22216);
or U22726 (N_22726,N_22437,N_22284);
nand U22727 (N_22727,N_22205,N_22292);
or U22728 (N_22728,N_22254,N_22341);
xnor U22729 (N_22729,N_22275,N_22294);
xor U22730 (N_22730,N_22263,N_22464);
and U22731 (N_22731,N_22324,N_22486);
and U22732 (N_22732,N_22421,N_22238);
and U22733 (N_22733,N_22264,N_22388);
xor U22734 (N_22734,N_22326,N_22408);
and U22735 (N_22735,N_22249,N_22352);
nand U22736 (N_22736,N_22388,N_22276);
xnor U22737 (N_22737,N_22475,N_22286);
nand U22738 (N_22738,N_22200,N_22427);
and U22739 (N_22739,N_22392,N_22285);
and U22740 (N_22740,N_22361,N_22445);
and U22741 (N_22741,N_22218,N_22252);
nand U22742 (N_22742,N_22269,N_22284);
nand U22743 (N_22743,N_22242,N_22345);
nor U22744 (N_22744,N_22498,N_22296);
nor U22745 (N_22745,N_22245,N_22368);
xor U22746 (N_22746,N_22460,N_22440);
and U22747 (N_22747,N_22266,N_22376);
nand U22748 (N_22748,N_22293,N_22211);
and U22749 (N_22749,N_22371,N_22429);
and U22750 (N_22750,N_22451,N_22341);
and U22751 (N_22751,N_22288,N_22243);
nand U22752 (N_22752,N_22379,N_22294);
and U22753 (N_22753,N_22451,N_22436);
or U22754 (N_22754,N_22494,N_22267);
nor U22755 (N_22755,N_22334,N_22400);
or U22756 (N_22756,N_22220,N_22299);
and U22757 (N_22757,N_22441,N_22490);
xnor U22758 (N_22758,N_22349,N_22302);
nor U22759 (N_22759,N_22214,N_22452);
nand U22760 (N_22760,N_22353,N_22331);
nand U22761 (N_22761,N_22268,N_22487);
and U22762 (N_22762,N_22453,N_22211);
xor U22763 (N_22763,N_22449,N_22242);
nand U22764 (N_22764,N_22216,N_22315);
nand U22765 (N_22765,N_22498,N_22288);
and U22766 (N_22766,N_22320,N_22394);
or U22767 (N_22767,N_22249,N_22379);
and U22768 (N_22768,N_22434,N_22250);
nor U22769 (N_22769,N_22361,N_22275);
and U22770 (N_22770,N_22427,N_22283);
and U22771 (N_22771,N_22232,N_22369);
and U22772 (N_22772,N_22498,N_22415);
or U22773 (N_22773,N_22387,N_22451);
or U22774 (N_22774,N_22241,N_22347);
nor U22775 (N_22775,N_22391,N_22403);
and U22776 (N_22776,N_22386,N_22273);
nor U22777 (N_22777,N_22379,N_22494);
nor U22778 (N_22778,N_22433,N_22371);
xor U22779 (N_22779,N_22264,N_22424);
nor U22780 (N_22780,N_22497,N_22365);
xnor U22781 (N_22781,N_22330,N_22206);
nor U22782 (N_22782,N_22354,N_22320);
nand U22783 (N_22783,N_22359,N_22442);
xnor U22784 (N_22784,N_22378,N_22202);
and U22785 (N_22785,N_22430,N_22314);
and U22786 (N_22786,N_22417,N_22437);
or U22787 (N_22787,N_22303,N_22450);
or U22788 (N_22788,N_22226,N_22425);
nand U22789 (N_22789,N_22444,N_22308);
xor U22790 (N_22790,N_22371,N_22241);
nand U22791 (N_22791,N_22406,N_22353);
nor U22792 (N_22792,N_22309,N_22238);
or U22793 (N_22793,N_22359,N_22312);
nor U22794 (N_22794,N_22231,N_22466);
or U22795 (N_22795,N_22206,N_22223);
or U22796 (N_22796,N_22299,N_22432);
nand U22797 (N_22797,N_22353,N_22377);
and U22798 (N_22798,N_22470,N_22408);
and U22799 (N_22799,N_22397,N_22385);
and U22800 (N_22800,N_22736,N_22598);
nor U22801 (N_22801,N_22593,N_22766);
nor U22802 (N_22802,N_22606,N_22573);
nand U22803 (N_22803,N_22665,N_22678);
nand U22804 (N_22804,N_22539,N_22611);
or U22805 (N_22805,N_22756,N_22647);
nand U22806 (N_22806,N_22641,N_22667);
xor U22807 (N_22807,N_22660,N_22741);
nand U22808 (N_22808,N_22698,N_22786);
nand U22809 (N_22809,N_22779,N_22623);
or U22810 (N_22810,N_22592,N_22735);
nor U22811 (N_22811,N_22501,N_22694);
xor U22812 (N_22812,N_22674,N_22575);
nand U22813 (N_22813,N_22625,N_22513);
nand U22814 (N_22814,N_22675,N_22719);
xnor U22815 (N_22815,N_22682,N_22572);
nor U22816 (N_22816,N_22703,N_22522);
or U22817 (N_22817,N_22765,N_22517);
or U22818 (N_22818,N_22595,N_22714);
nor U22819 (N_22819,N_22755,N_22791);
xnor U22820 (N_22820,N_22596,N_22732);
nand U22821 (N_22821,N_22689,N_22559);
or U22822 (N_22822,N_22567,N_22734);
nand U22823 (N_22823,N_22781,N_22551);
nor U22824 (N_22824,N_22507,N_22650);
and U22825 (N_22825,N_22688,N_22785);
nor U22826 (N_22826,N_22696,N_22670);
xnor U22827 (N_22827,N_22654,N_22643);
xnor U22828 (N_22828,N_22731,N_22629);
and U22829 (N_22829,N_22776,N_22799);
and U22830 (N_22830,N_22740,N_22789);
and U22831 (N_22831,N_22686,N_22767);
or U22832 (N_22832,N_22639,N_22697);
xor U22833 (N_22833,N_22750,N_22742);
nand U22834 (N_22834,N_22608,N_22603);
nand U22835 (N_22835,N_22653,N_22531);
xnor U22836 (N_22836,N_22502,N_22536);
nor U22837 (N_22837,N_22628,N_22524);
nand U22838 (N_22838,N_22617,N_22797);
or U22839 (N_22839,N_22587,N_22630);
or U22840 (N_22840,N_22514,N_22687);
nand U22841 (N_22841,N_22622,N_22646);
nor U22842 (N_22842,N_22684,N_22645);
or U22843 (N_22843,N_22535,N_22683);
nor U22844 (N_22844,N_22768,N_22597);
xnor U22845 (N_22845,N_22508,N_22605);
nand U22846 (N_22846,N_22761,N_22612);
xnor U22847 (N_22847,N_22542,N_22792);
or U22848 (N_22848,N_22588,N_22538);
and U22849 (N_22849,N_22685,N_22614);
nand U22850 (N_22850,N_22574,N_22635);
nand U22851 (N_22851,N_22532,N_22648);
nand U22852 (N_22852,N_22525,N_22657);
and U22853 (N_22853,N_22631,N_22730);
nor U22854 (N_22854,N_22794,N_22726);
nand U22855 (N_22855,N_22744,N_22533);
xnor U22856 (N_22856,N_22618,N_22724);
nand U22857 (N_22857,N_22748,N_22621);
or U22858 (N_22858,N_22590,N_22519);
nor U22859 (N_22859,N_22527,N_22552);
and U22860 (N_22860,N_22661,N_22638);
nand U22861 (N_22861,N_22775,N_22560);
or U22862 (N_22862,N_22770,N_22619);
nor U22863 (N_22863,N_22585,N_22634);
nand U22864 (N_22864,N_22652,N_22745);
xor U22865 (N_22865,N_22782,N_22672);
and U22866 (N_22866,N_22566,N_22721);
nor U22867 (N_22867,N_22757,N_22795);
and U22868 (N_22868,N_22610,N_22700);
nand U22869 (N_22869,N_22568,N_22570);
or U22870 (N_22870,N_22743,N_22576);
nor U22871 (N_22871,N_22722,N_22707);
or U22872 (N_22872,N_22505,N_22582);
nand U22873 (N_22873,N_22717,N_22540);
and U22874 (N_22874,N_22788,N_22562);
nand U22875 (N_22875,N_22777,N_22579);
nand U22876 (N_22876,N_22746,N_22725);
and U22877 (N_22877,N_22520,N_22772);
nand U22878 (N_22878,N_22602,N_22710);
xnor U22879 (N_22879,N_22787,N_22589);
or U22880 (N_22880,N_22708,N_22681);
xor U22881 (N_22881,N_22695,N_22547);
and U22882 (N_22882,N_22626,N_22565);
and U22883 (N_22883,N_22556,N_22546);
or U22884 (N_22884,N_22764,N_22680);
nor U22885 (N_22885,N_22558,N_22754);
or U22886 (N_22886,N_22506,N_22604);
nand U22887 (N_22887,N_22600,N_22516);
xnor U22888 (N_22888,N_22543,N_22671);
xor U22889 (N_22889,N_22711,N_22561);
or U22890 (N_22890,N_22702,N_22774);
nand U22891 (N_22891,N_22500,N_22583);
nor U22892 (N_22892,N_22580,N_22658);
nor U22893 (N_22893,N_22607,N_22594);
and U22894 (N_22894,N_22541,N_22727);
xnor U22895 (N_22895,N_22769,N_22728);
xor U22896 (N_22896,N_22581,N_22503);
xnor U22897 (N_22897,N_22762,N_22712);
nor U22898 (N_22898,N_22557,N_22571);
or U22899 (N_22899,N_22749,N_22518);
or U22900 (N_22900,N_22627,N_22550);
nand U22901 (N_22901,N_22729,N_22705);
nor U22902 (N_22902,N_22739,N_22663);
xnor U22903 (N_22903,N_22763,N_22668);
xor U22904 (N_22904,N_22511,N_22656);
and U22905 (N_22905,N_22793,N_22640);
nand U22906 (N_22906,N_22528,N_22758);
nand U22907 (N_22907,N_22677,N_22632);
nor U22908 (N_22908,N_22718,N_22615);
nand U22909 (N_22909,N_22549,N_22624);
nand U22910 (N_22910,N_22796,N_22798);
or U22911 (N_22911,N_22530,N_22752);
and U22912 (N_22912,N_22642,N_22704);
xnor U22913 (N_22913,N_22780,N_22523);
or U22914 (N_22914,N_22679,N_22716);
nand U22915 (N_22915,N_22751,N_22690);
nand U22916 (N_22916,N_22578,N_22673);
and U22917 (N_22917,N_22521,N_22599);
nor U22918 (N_22918,N_22644,N_22633);
and U22919 (N_22919,N_22555,N_22509);
nor U22920 (N_22920,N_22586,N_22691);
or U22921 (N_22921,N_22738,N_22655);
nor U22922 (N_22922,N_22737,N_22537);
nor U22923 (N_22923,N_22591,N_22620);
xnor U22924 (N_22924,N_22783,N_22659);
nor U22925 (N_22925,N_22693,N_22613);
or U22926 (N_22926,N_22601,N_22664);
and U22927 (N_22927,N_22699,N_22720);
nor U22928 (N_22928,N_22713,N_22577);
xor U22929 (N_22929,N_22616,N_22747);
and U22930 (N_22930,N_22649,N_22676);
and U22931 (N_22931,N_22692,N_22760);
and U22932 (N_22932,N_22545,N_22669);
nor U22933 (N_22933,N_22564,N_22569);
and U22934 (N_22934,N_22504,N_22584);
and U22935 (N_22935,N_22790,N_22771);
xor U22936 (N_22936,N_22709,N_22515);
nand U22937 (N_22937,N_22666,N_22510);
nand U22938 (N_22938,N_22637,N_22701);
xor U22939 (N_22939,N_22778,N_22544);
or U22940 (N_22940,N_22534,N_22784);
nor U22941 (N_22941,N_22636,N_22553);
and U22942 (N_22942,N_22526,N_22609);
xor U22943 (N_22943,N_22723,N_22753);
nor U22944 (N_22944,N_22759,N_22662);
and U22945 (N_22945,N_22706,N_22512);
xor U22946 (N_22946,N_22733,N_22554);
nor U22947 (N_22947,N_22651,N_22529);
and U22948 (N_22948,N_22715,N_22563);
nor U22949 (N_22949,N_22773,N_22548);
nor U22950 (N_22950,N_22728,N_22790);
xor U22951 (N_22951,N_22624,N_22758);
nor U22952 (N_22952,N_22640,N_22567);
or U22953 (N_22953,N_22658,N_22585);
xor U22954 (N_22954,N_22740,N_22576);
nand U22955 (N_22955,N_22619,N_22620);
and U22956 (N_22956,N_22793,N_22612);
nor U22957 (N_22957,N_22764,N_22732);
and U22958 (N_22958,N_22549,N_22726);
nor U22959 (N_22959,N_22634,N_22750);
and U22960 (N_22960,N_22596,N_22738);
xnor U22961 (N_22961,N_22637,N_22564);
nor U22962 (N_22962,N_22631,N_22604);
or U22963 (N_22963,N_22610,N_22736);
or U22964 (N_22964,N_22765,N_22544);
nor U22965 (N_22965,N_22655,N_22649);
or U22966 (N_22966,N_22540,N_22703);
or U22967 (N_22967,N_22670,N_22549);
or U22968 (N_22968,N_22611,N_22515);
and U22969 (N_22969,N_22682,N_22579);
and U22970 (N_22970,N_22715,N_22610);
xnor U22971 (N_22971,N_22644,N_22773);
xnor U22972 (N_22972,N_22723,N_22554);
nand U22973 (N_22973,N_22551,N_22542);
or U22974 (N_22974,N_22630,N_22504);
xnor U22975 (N_22975,N_22528,N_22572);
xor U22976 (N_22976,N_22580,N_22749);
xnor U22977 (N_22977,N_22570,N_22767);
nand U22978 (N_22978,N_22552,N_22665);
nor U22979 (N_22979,N_22617,N_22691);
xor U22980 (N_22980,N_22778,N_22599);
nor U22981 (N_22981,N_22504,N_22730);
or U22982 (N_22982,N_22726,N_22682);
xnor U22983 (N_22983,N_22554,N_22694);
nor U22984 (N_22984,N_22711,N_22675);
and U22985 (N_22985,N_22696,N_22743);
xnor U22986 (N_22986,N_22777,N_22689);
nand U22987 (N_22987,N_22704,N_22693);
nor U22988 (N_22988,N_22717,N_22524);
and U22989 (N_22989,N_22728,N_22701);
nand U22990 (N_22990,N_22572,N_22757);
xnor U22991 (N_22991,N_22511,N_22698);
nand U22992 (N_22992,N_22692,N_22538);
nand U22993 (N_22993,N_22620,N_22579);
xnor U22994 (N_22994,N_22641,N_22758);
and U22995 (N_22995,N_22666,N_22594);
xor U22996 (N_22996,N_22706,N_22520);
or U22997 (N_22997,N_22636,N_22526);
nor U22998 (N_22998,N_22681,N_22697);
nor U22999 (N_22999,N_22794,N_22561);
nor U23000 (N_23000,N_22597,N_22640);
xnor U23001 (N_23001,N_22509,N_22527);
xnor U23002 (N_23002,N_22683,N_22792);
or U23003 (N_23003,N_22537,N_22678);
nand U23004 (N_23004,N_22569,N_22696);
xor U23005 (N_23005,N_22702,N_22748);
nor U23006 (N_23006,N_22798,N_22715);
or U23007 (N_23007,N_22749,N_22791);
xor U23008 (N_23008,N_22611,N_22546);
nand U23009 (N_23009,N_22718,N_22747);
xnor U23010 (N_23010,N_22771,N_22599);
and U23011 (N_23011,N_22722,N_22587);
or U23012 (N_23012,N_22545,N_22556);
nor U23013 (N_23013,N_22617,N_22679);
or U23014 (N_23014,N_22781,N_22503);
xnor U23015 (N_23015,N_22573,N_22567);
nor U23016 (N_23016,N_22722,N_22765);
nor U23017 (N_23017,N_22565,N_22634);
and U23018 (N_23018,N_22543,N_22609);
and U23019 (N_23019,N_22782,N_22637);
and U23020 (N_23020,N_22769,N_22542);
nor U23021 (N_23021,N_22595,N_22519);
or U23022 (N_23022,N_22706,N_22569);
xnor U23023 (N_23023,N_22516,N_22788);
nor U23024 (N_23024,N_22566,N_22734);
nor U23025 (N_23025,N_22644,N_22733);
nor U23026 (N_23026,N_22790,N_22549);
nor U23027 (N_23027,N_22715,N_22642);
nor U23028 (N_23028,N_22569,N_22766);
nand U23029 (N_23029,N_22634,N_22524);
nor U23030 (N_23030,N_22575,N_22502);
and U23031 (N_23031,N_22525,N_22661);
nor U23032 (N_23032,N_22596,N_22529);
or U23033 (N_23033,N_22663,N_22646);
or U23034 (N_23034,N_22768,N_22716);
or U23035 (N_23035,N_22682,N_22693);
xnor U23036 (N_23036,N_22743,N_22787);
nor U23037 (N_23037,N_22622,N_22775);
nand U23038 (N_23038,N_22618,N_22756);
nor U23039 (N_23039,N_22589,N_22768);
and U23040 (N_23040,N_22580,N_22746);
or U23041 (N_23041,N_22525,N_22776);
xnor U23042 (N_23042,N_22704,N_22787);
nor U23043 (N_23043,N_22633,N_22606);
nand U23044 (N_23044,N_22513,N_22543);
and U23045 (N_23045,N_22525,N_22780);
or U23046 (N_23046,N_22659,N_22791);
nand U23047 (N_23047,N_22775,N_22556);
xnor U23048 (N_23048,N_22507,N_22563);
nand U23049 (N_23049,N_22552,N_22521);
xnor U23050 (N_23050,N_22565,N_22522);
nor U23051 (N_23051,N_22663,N_22743);
nor U23052 (N_23052,N_22780,N_22770);
nand U23053 (N_23053,N_22792,N_22722);
and U23054 (N_23054,N_22555,N_22536);
nand U23055 (N_23055,N_22642,N_22793);
nor U23056 (N_23056,N_22635,N_22647);
nor U23057 (N_23057,N_22520,N_22727);
and U23058 (N_23058,N_22695,N_22667);
or U23059 (N_23059,N_22656,N_22615);
nor U23060 (N_23060,N_22657,N_22759);
and U23061 (N_23061,N_22570,N_22653);
xor U23062 (N_23062,N_22504,N_22698);
nor U23063 (N_23063,N_22578,N_22790);
nand U23064 (N_23064,N_22678,N_22561);
xnor U23065 (N_23065,N_22721,N_22599);
or U23066 (N_23066,N_22762,N_22624);
or U23067 (N_23067,N_22747,N_22562);
nand U23068 (N_23068,N_22688,N_22677);
nor U23069 (N_23069,N_22506,N_22735);
nand U23070 (N_23070,N_22725,N_22560);
nor U23071 (N_23071,N_22748,N_22761);
nor U23072 (N_23072,N_22661,N_22722);
and U23073 (N_23073,N_22718,N_22523);
nand U23074 (N_23074,N_22609,N_22633);
nand U23075 (N_23075,N_22753,N_22590);
xnor U23076 (N_23076,N_22723,N_22523);
xnor U23077 (N_23077,N_22642,N_22739);
xnor U23078 (N_23078,N_22672,N_22764);
nand U23079 (N_23079,N_22613,N_22649);
or U23080 (N_23080,N_22534,N_22517);
xnor U23081 (N_23081,N_22600,N_22551);
xnor U23082 (N_23082,N_22610,N_22526);
nand U23083 (N_23083,N_22692,N_22718);
xnor U23084 (N_23084,N_22723,N_22575);
and U23085 (N_23085,N_22671,N_22501);
nand U23086 (N_23086,N_22776,N_22780);
xor U23087 (N_23087,N_22514,N_22675);
nand U23088 (N_23088,N_22633,N_22574);
or U23089 (N_23089,N_22711,N_22589);
or U23090 (N_23090,N_22509,N_22537);
and U23091 (N_23091,N_22546,N_22562);
xor U23092 (N_23092,N_22632,N_22748);
and U23093 (N_23093,N_22654,N_22655);
or U23094 (N_23094,N_22724,N_22512);
nand U23095 (N_23095,N_22639,N_22642);
and U23096 (N_23096,N_22738,N_22641);
and U23097 (N_23097,N_22559,N_22520);
xor U23098 (N_23098,N_22764,N_22582);
and U23099 (N_23099,N_22711,N_22610);
nand U23100 (N_23100,N_23006,N_22816);
and U23101 (N_23101,N_22813,N_22914);
nor U23102 (N_23102,N_23095,N_22908);
nand U23103 (N_23103,N_22889,N_22828);
and U23104 (N_23104,N_22948,N_23036);
and U23105 (N_23105,N_23069,N_22852);
xor U23106 (N_23106,N_22976,N_22903);
xnor U23107 (N_23107,N_22917,N_23055);
xor U23108 (N_23108,N_22910,N_22974);
and U23109 (N_23109,N_22977,N_22878);
or U23110 (N_23110,N_22832,N_23063);
nor U23111 (N_23111,N_23079,N_22823);
and U23112 (N_23112,N_22909,N_23005);
nor U23113 (N_23113,N_23098,N_22811);
or U23114 (N_23114,N_22869,N_22807);
or U23115 (N_23115,N_23059,N_22947);
xor U23116 (N_23116,N_23047,N_22956);
xor U23117 (N_23117,N_22839,N_22965);
or U23118 (N_23118,N_22980,N_23011);
nor U23119 (N_23119,N_22942,N_22997);
nor U23120 (N_23120,N_23058,N_22949);
or U23121 (N_23121,N_22944,N_23066);
and U23122 (N_23122,N_22919,N_23082);
and U23123 (N_23123,N_23039,N_22911);
and U23124 (N_23124,N_22945,N_22985);
nor U23125 (N_23125,N_23057,N_22900);
nor U23126 (N_23126,N_22935,N_23031);
nor U23127 (N_23127,N_23083,N_23026);
xnor U23128 (N_23128,N_22814,N_23075);
or U23129 (N_23129,N_22931,N_22955);
xor U23130 (N_23130,N_23099,N_22926);
and U23131 (N_23131,N_22891,N_22859);
nor U23132 (N_23132,N_23056,N_22975);
and U23133 (N_23133,N_22915,N_23061);
nand U23134 (N_23134,N_22970,N_22898);
nand U23135 (N_23135,N_23091,N_22809);
xor U23136 (N_23136,N_22857,N_22888);
and U23137 (N_23137,N_22817,N_23040);
xor U23138 (N_23138,N_23096,N_22899);
and U23139 (N_23139,N_22879,N_22993);
nor U23140 (N_23140,N_22834,N_23089);
and U23141 (N_23141,N_22907,N_22983);
nor U23142 (N_23142,N_22886,N_22841);
nand U23143 (N_23143,N_22925,N_23092);
and U23144 (N_23144,N_23019,N_22962);
nor U23145 (N_23145,N_22966,N_22822);
xnor U23146 (N_23146,N_22961,N_22906);
and U23147 (N_23147,N_23086,N_22860);
xnor U23148 (N_23148,N_22881,N_22991);
nand U23149 (N_23149,N_22994,N_23032);
nand U23150 (N_23150,N_23008,N_22831);
xor U23151 (N_23151,N_22835,N_22981);
xor U23152 (N_23152,N_22920,N_22842);
xnor U23153 (N_23153,N_23045,N_22856);
or U23154 (N_23154,N_22896,N_22957);
or U23155 (N_23155,N_22953,N_22854);
and U23156 (N_23156,N_23070,N_22850);
or U23157 (N_23157,N_23009,N_22904);
nor U23158 (N_23158,N_22868,N_22912);
or U23159 (N_23159,N_22923,N_22876);
nand U23160 (N_23160,N_23085,N_23018);
nor U23161 (N_23161,N_22996,N_22825);
and U23162 (N_23162,N_23020,N_22936);
nand U23163 (N_23163,N_23012,N_22826);
and U23164 (N_23164,N_22838,N_22928);
nor U23165 (N_23165,N_22837,N_23010);
nand U23166 (N_23166,N_22855,N_23080);
xor U23167 (N_23167,N_23021,N_22801);
xnor U23168 (N_23168,N_22890,N_22901);
nand U23169 (N_23169,N_23071,N_22853);
nand U23170 (N_23170,N_22951,N_22916);
nand U23171 (N_23171,N_22845,N_22821);
nand U23172 (N_23172,N_22973,N_22893);
or U23173 (N_23173,N_22865,N_22918);
nor U23174 (N_23174,N_22851,N_23028);
and U23175 (N_23175,N_22885,N_23077);
nor U23176 (N_23176,N_22932,N_23024);
xnor U23177 (N_23177,N_22963,N_22964);
nor U23178 (N_23178,N_22972,N_23043);
nor U23179 (N_23179,N_22810,N_23003);
nand U23180 (N_23180,N_22806,N_22938);
and U23181 (N_23181,N_22830,N_22802);
and U23182 (N_23182,N_22874,N_22897);
nand U23183 (N_23183,N_23060,N_23052);
or U23184 (N_23184,N_23054,N_23065);
nor U23185 (N_23185,N_23041,N_23027);
and U23186 (N_23186,N_22844,N_22892);
nor U23187 (N_23187,N_23094,N_23081);
and U23188 (N_23188,N_23044,N_22954);
xor U23189 (N_23189,N_23048,N_23087);
nor U23190 (N_23190,N_22847,N_22827);
nand U23191 (N_23191,N_22934,N_22987);
nor U23192 (N_23192,N_22969,N_23042);
and U23193 (N_23193,N_22863,N_22984);
and U23194 (N_23194,N_23034,N_23013);
nor U23195 (N_23195,N_22986,N_22982);
and U23196 (N_23196,N_22819,N_22927);
and U23197 (N_23197,N_22967,N_22992);
nor U23198 (N_23198,N_22941,N_23067);
or U23199 (N_23199,N_22833,N_22999);
nor U23200 (N_23200,N_23062,N_22894);
xor U23201 (N_23201,N_23016,N_22959);
nor U23202 (N_23202,N_23051,N_22820);
xnor U23203 (N_23203,N_22871,N_23014);
nor U23204 (N_23204,N_23076,N_22978);
or U23205 (N_23205,N_22943,N_22924);
or U23206 (N_23206,N_22905,N_22808);
xnor U23207 (N_23207,N_22968,N_23023);
xnor U23208 (N_23208,N_22960,N_22922);
or U23209 (N_23209,N_23035,N_22858);
and U23210 (N_23210,N_23053,N_22861);
nand U23211 (N_23211,N_22846,N_23073);
and U23212 (N_23212,N_23001,N_22979);
or U23213 (N_23213,N_23072,N_23000);
and U23214 (N_23214,N_23068,N_22872);
xnor U23215 (N_23215,N_22836,N_23090);
or U23216 (N_23216,N_22989,N_22882);
xnor U23217 (N_23217,N_22902,N_23084);
nor U23218 (N_23218,N_22933,N_22812);
nand U23219 (N_23219,N_22913,N_22829);
nand U23220 (N_23220,N_22803,N_22873);
or U23221 (N_23221,N_22921,N_22877);
and U23222 (N_23222,N_22946,N_23022);
nand U23223 (N_23223,N_22815,N_22990);
or U23224 (N_23224,N_22883,N_23029);
or U23225 (N_23225,N_22805,N_23097);
nor U23226 (N_23226,N_22866,N_22995);
xnor U23227 (N_23227,N_22880,N_22958);
nor U23228 (N_23228,N_23025,N_22939);
nor U23229 (N_23229,N_22840,N_22875);
or U23230 (N_23230,N_23049,N_23074);
nor U23231 (N_23231,N_23093,N_22929);
or U23232 (N_23232,N_22804,N_22849);
and U23233 (N_23233,N_23038,N_23050);
nor U23234 (N_23234,N_22864,N_23046);
nor U23235 (N_23235,N_23033,N_22998);
and U23236 (N_23236,N_23064,N_22843);
or U23237 (N_23237,N_23078,N_23088);
or U23238 (N_23238,N_22937,N_22870);
nor U23239 (N_23239,N_23015,N_23007);
nor U23240 (N_23240,N_22940,N_22848);
nand U23241 (N_23241,N_22988,N_22800);
xor U23242 (N_23242,N_22971,N_22884);
or U23243 (N_23243,N_22824,N_23004);
or U23244 (N_23244,N_22818,N_22867);
nor U23245 (N_23245,N_23030,N_22930);
and U23246 (N_23246,N_22895,N_22950);
nor U23247 (N_23247,N_22862,N_23017);
and U23248 (N_23248,N_23037,N_23002);
or U23249 (N_23249,N_22952,N_22887);
nand U23250 (N_23250,N_23024,N_22921);
nor U23251 (N_23251,N_22938,N_22802);
xnor U23252 (N_23252,N_22835,N_22862);
nor U23253 (N_23253,N_22835,N_22938);
nand U23254 (N_23254,N_23050,N_22846);
xnor U23255 (N_23255,N_22981,N_22968);
xor U23256 (N_23256,N_23078,N_23018);
or U23257 (N_23257,N_22998,N_22904);
xor U23258 (N_23258,N_22965,N_22957);
xnor U23259 (N_23259,N_23008,N_22829);
nor U23260 (N_23260,N_22826,N_23043);
nand U23261 (N_23261,N_22838,N_23049);
xor U23262 (N_23262,N_22878,N_22824);
nand U23263 (N_23263,N_23072,N_22945);
nor U23264 (N_23264,N_22922,N_23070);
nor U23265 (N_23265,N_22984,N_22832);
nand U23266 (N_23266,N_22870,N_22892);
nor U23267 (N_23267,N_22974,N_22879);
xor U23268 (N_23268,N_23064,N_22997);
nand U23269 (N_23269,N_22977,N_23006);
xnor U23270 (N_23270,N_22998,N_22927);
nor U23271 (N_23271,N_23069,N_22802);
nor U23272 (N_23272,N_22897,N_22927);
nor U23273 (N_23273,N_22987,N_22937);
or U23274 (N_23274,N_23030,N_22994);
and U23275 (N_23275,N_23059,N_22876);
and U23276 (N_23276,N_22816,N_22944);
xor U23277 (N_23277,N_22803,N_23050);
xor U23278 (N_23278,N_22989,N_22820);
and U23279 (N_23279,N_22893,N_22866);
nor U23280 (N_23280,N_22819,N_22865);
nand U23281 (N_23281,N_22810,N_23064);
or U23282 (N_23282,N_23082,N_22992);
xor U23283 (N_23283,N_23038,N_22824);
xnor U23284 (N_23284,N_23060,N_23072);
or U23285 (N_23285,N_22949,N_22908);
xnor U23286 (N_23286,N_23076,N_22996);
nand U23287 (N_23287,N_22989,N_23022);
nand U23288 (N_23288,N_23046,N_22990);
nor U23289 (N_23289,N_23067,N_22883);
nand U23290 (N_23290,N_22905,N_23014);
nor U23291 (N_23291,N_23093,N_23021);
nand U23292 (N_23292,N_22928,N_22941);
and U23293 (N_23293,N_23090,N_22993);
xor U23294 (N_23294,N_22832,N_22964);
or U23295 (N_23295,N_22966,N_22811);
nor U23296 (N_23296,N_22908,N_22938);
nand U23297 (N_23297,N_22835,N_22980);
xor U23298 (N_23298,N_23045,N_23083);
xnor U23299 (N_23299,N_23070,N_23075);
xor U23300 (N_23300,N_23017,N_23060);
and U23301 (N_23301,N_23033,N_22944);
or U23302 (N_23302,N_22875,N_22979);
xnor U23303 (N_23303,N_22803,N_22847);
nand U23304 (N_23304,N_22910,N_22866);
and U23305 (N_23305,N_22853,N_22925);
or U23306 (N_23306,N_22820,N_23070);
and U23307 (N_23307,N_22809,N_22997);
or U23308 (N_23308,N_22955,N_22806);
xnor U23309 (N_23309,N_22888,N_22908);
or U23310 (N_23310,N_22895,N_23037);
xnor U23311 (N_23311,N_23021,N_22980);
xor U23312 (N_23312,N_23052,N_22942);
xor U23313 (N_23313,N_22954,N_22852);
xnor U23314 (N_23314,N_22967,N_22938);
nand U23315 (N_23315,N_23060,N_22858);
xnor U23316 (N_23316,N_22872,N_22848);
nand U23317 (N_23317,N_22923,N_23007);
nand U23318 (N_23318,N_23019,N_22913);
and U23319 (N_23319,N_22845,N_23016);
and U23320 (N_23320,N_22912,N_22852);
nand U23321 (N_23321,N_22901,N_22975);
nor U23322 (N_23322,N_22977,N_22881);
nand U23323 (N_23323,N_22985,N_22862);
nor U23324 (N_23324,N_22983,N_22894);
or U23325 (N_23325,N_22914,N_22936);
and U23326 (N_23326,N_22913,N_22897);
and U23327 (N_23327,N_22951,N_23061);
xnor U23328 (N_23328,N_23007,N_22876);
or U23329 (N_23329,N_23092,N_23088);
xnor U23330 (N_23330,N_22944,N_22886);
and U23331 (N_23331,N_22837,N_23056);
and U23332 (N_23332,N_22816,N_23001);
nand U23333 (N_23333,N_22810,N_22906);
nand U23334 (N_23334,N_23071,N_22839);
or U23335 (N_23335,N_23087,N_22820);
xor U23336 (N_23336,N_22939,N_23059);
xor U23337 (N_23337,N_22934,N_22808);
nor U23338 (N_23338,N_23064,N_22912);
nand U23339 (N_23339,N_22895,N_22901);
or U23340 (N_23340,N_22858,N_22922);
nor U23341 (N_23341,N_22803,N_22855);
or U23342 (N_23342,N_23060,N_22864);
nand U23343 (N_23343,N_23072,N_22888);
xnor U23344 (N_23344,N_23087,N_22953);
nand U23345 (N_23345,N_22855,N_22880);
nor U23346 (N_23346,N_22883,N_23046);
and U23347 (N_23347,N_22882,N_22944);
nand U23348 (N_23348,N_22900,N_22864);
or U23349 (N_23349,N_22937,N_23096);
and U23350 (N_23350,N_22876,N_22865);
nand U23351 (N_23351,N_22824,N_22854);
and U23352 (N_23352,N_22842,N_22815);
or U23353 (N_23353,N_22942,N_22821);
or U23354 (N_23354,N_22873,N_22998);
or U23355 (N_23355,N_22897,N_22846);
and U23356 (N_23356,N_22929,N_22958);
or U23357 (N_23357,N_22970,N_23052);
nor U23358 (N_23358,N_23097,N_22979);
nand U23359 (N_23359,N_23010,N_22804);
nor U23360 (N_23360,N_22990,N_22857);
or U23361 (N_23361,N_22803,N_22845);
and U23362 (N_23362,N_22928,N_23098);
or U23363 (N_23363,N_23018,N_22990);
nor U23364 (N_23364,N_23035,N_22976);
or U23365 (N_23365,N_23060,N_22963);
and U23366 (N_23366,N_23052,N_23028);
and U23367 (N_23367,N_22973,N_22811);
nor U23368 (N_23368,N_22999,N_22869);
nor U23369 (N_23369,N_23082,N_22891);
xnor U23370 (N_23370,N_23013,N_22917);
and U23371 (N_23371,N_22812,N_23045);
nand U23372 (N_23372,N_22960,N_22876);
nand U23373 (N_23373,N_23069,N_22953);
nand U23374 (N_23374,N_22958,N_22941);
or U23375 (N_23375,N_22972,N_22854);
nand U23376 (N_23376,N_22856,N_22812);
and U23377 (N_23377,N_22909,N_23096);
xnor U23378 (N_23378,N_22985,N_22817);
nand U23379 (N_23379,N_22899,N_23054);
or U23380 (N_23380,N_23065,N_22984);
or U23381 (N_23381,N_23027,N_22929);
nand U23382 (N_23382,N_22804,N_23075);
nor U23383 (N_23383,N_22980,N_22876);
or U23384 (N_23384,N_23083,N_22914);
and U23385 (N_23385,N_22954,N_22877);
xnor U23386 (N_23386,N_22827,N_22858);
and U23387 (N_23387,N_22919,N_23021);
xnor U23388 (N_23388,N_22889,N_22998);
nor U23389 (N_23389,N_22858,N_22823);
nand U23390 (N_23390,N_23083,N_22947);
nand U23391 (N_23391,N_22924,N_22820);
nand U23392 (N_23392,N_22942,N_22959);
xor U23393 (N_23393,N_22901,N_22931);
nor U23394 (N_23394,N_22998,N_22865);
xnor U23395 (N_23395,N_23029,N_22967);
nand U23396 (N_23396,N_22852,N_22925);
nand U23397 (N_23397,N_22951,N_22935);
and U23398 (N_23398,N_22806,N_22986);
or U23399 (N_23399,N_23008,N_23047);
or U23400 (N_23400,N_23206,N_23367);
xor U23401 (N_23401,N_23167,N_23321);
nand U23402 (N_23402,N_23198,N_23165);
and U23403 (N_23403,N_23288,N_23391);
and U23404 (N_23404,N_23223,N_23107);
or U23405 (N_23405,N_23247,N_23205);
and U23406 (N_23406,N_23369,N_23377);
or U23407 (N_23407,N_23358,N_23149);
nor U23408 (N_23408,N_23300,N_23246);
xor U23409 (N_23409,N_23309,N_23118);
nor U23410 (N_23410,N_23155,N_23383);
and U23411 (N_23411,N_23217,N_23325);
and U23412 (N_23412,N_23259,N_23251);
nand U23413 (N_23413,N_23131,N_23177);
and U23414 (N_23414,N_23101,N_23228);
nand U23415 (N_23415,N_23237,N_23194);
xor U23416 (N_23416,N_23153,N_23121);
nand U23417 (N_23417,N_23276,N_23241);
nand U23418 (N_23418,N_23388,N_23371);
and U23419 (N_23419,N_23179,N_23133);
xnor U23420 (N_23420,N_23141,N_23227);
nand U23421 (N_23421,N_23307,N_23170);
nor U23422 (N_23422,N_23310,N_23176);
nor U23423 (N_23423,N_23320,N_23122);
nand U23424 (N_23424,N_23266,N_23372);
nand U23425 (N_23425,N_23108,N_23392);
xor U23426 (N_23426,N_23350,N_23336);
or U23427 (N_23427,N_23314,N_23202);
xor U23428 (N_23428,N_23352,N_23190);
xor U23429 (N_23429,N_23154,N_23346);
nor U23430 (N_23430,N_23306,N_23337);
or U23431 (N_23431,N_23362,N_23329);
xnor U23432 (N_23432,N_23215,N_23220);
nor U23433 (N_23433,N_23342,N_23347);
nand U23434 (N_23434,N_23114,N_23263);
and U23435 (N_23435,N_23102,N_23393);
nand U23436 (N_23436,N_23229,N_23315);
or U23437 (N_23437,N_23104,N_23399);
nand U23438 (N_23438,N_23210,N_23373);
xor U23439 (N_23439,N_23117,N_23250);
nand U23440 (N_23440,N_23270,N_23232);
and U23441 (N_23441,N_23389,N_23258);
nor U23442 (N_23442,N_23111,N_23208);
and U23443 (N_23443,N_23380,N_23302);
and U23444 (N_23444,N_23376,N_23226);
xor U23445 (N_23445,N_23191,N_23368);
xor U23446 (N_23446,N_23152,N_23254);
nand U23447 (N_23447,N_23283,N_23284);
xnor U23448 (N_23448,N_23299,N_23142);
nand U23449 (N_23449,N_23249,N_23338);
nor U23450 (N_23450,N_23242,N_23116);
nor U23451 (N_23451,N_23305,N_23100);
nor U23452 (N_23452,N_23356,N_23292);
nor U23453 (N_23453,N_23304,N_23290);
xor U23454 (N_23454,N_23124,N_23230);
nor U23455 (N_23455,N_23221,N_23178);
xnor U23456 (N_23456,N_23162,N_23113);
nor U23457 (N_23457,N_23192,N_23378);
or U23458 (N_23458,N_23134,N_23274);
xnor U23459 (N_23459,N_23382,N_23253);
xor U23460 (N_23460,N_23390,N_23126);
nor U23461 (N_23461,N_23252,N_23257);
nor U23462 (N_23462,N_23218,N_23161);
xnor U23463 (N_23463,N_23261,N_23197);
and U23464 (N_23464,N_23301,N_23151);
nand U23465 (N_23465,N_23278,N_23319);
or U23466 (N_23466,N_23282,N_23243);
nor U23467 (N_23467,N_23156,N_23384);
and U23468 (N_23468,N_23354,N_23199);
nor U23469 (N_23469,N_23169,N_23289);
and U23470 (N_23470,N_23203,N_23180);
and U23471 (N_23471,N_23385,N_23398);
or U23472 (N_23472,N_23109,N_23333);
nor U23473 (N_23473,N_23244,N_23201);
nor U23474 (N_23474,N_23387,N_23264);
nand U23475 (N_23475,N_23394,N_23328);
or U23476 (N_23476,N_23164,N_23163);
nand U23477 (N_23477,N_23291,N_23150);
or U23478 (N_23478,N_23360,N_23119);
or U23479 (N_23479,N_23211,N_23129);
and U23480 (N_23480,N_23312,N_23331);
and U23481 (N_23481,N_23255,N_23365);
or U23482 (N_23482,N_23269,N_23132);
and U23483 (N_23483,N_23157,N_23359);
and U23484 (N_23484,N_23240,N_23143);
and U23485 (N_23485,N_23195,N_23125);
xnor U23486 (N_23486,N_23245,N_23193);
and U23487 (N_23487,N_23224,N_23137);
nor U23488 (N_23488,N_23375,N_23330);
or U23489 (N_23489,N_23322,N_23268);
xor U23490 (N_23490,N_23366,N_23106);
or U23491 (N_23491,N_23207,N_23339);
nand U23492 (N_23492,N_23138,N_23172);
nor U23493 (N_23493,N_23334,N_23363);
and U23494 (N_23494,N_23222,N_23140);
or U23495 (N_23495,N_23216,N_23265);
and U23496 (N_23496,N_23135,N_23213);
xor U23497 (N_23497,N_23386,N_23145);
or U23498 (N_23498,N_23357,N_23335);
and U23499 (N_23499,N_23209,N_23296);
nor U23500 (N_23500,N_23271,N_23341);
nand U23501 (N_23501,N_23311,N_23295);
nor U23502 (N_23502,N_23395,N_23238);
or U23503 (N_23503,N_23281,N_23214);
or U23504 (N_23504,N_23256,N_23234);
and U23505 (N_23505,N_23146,N_23317);
xor U23506 (N_23506,N_23260,N_23148);
xnor U23507 (N_23507,N_23351,N_23147);
xor U23508 (N_23508,N_23287,N_23316);
and U23509 (N_23509,N_23158,N_23188);
nand U23510 (N_23510,N_23231,N_23168);
nand U23511 (N_23511,N_23381,N_23103);
and U23512 (N_23512,N_23323,N_23204);
nor U23513 (N_23513,N_23189,N_23267);
or U23514 (N_23514,N_23279,N_23343);
xor U23515 (N_23515,N_23313,N_23123);
nand U23516 (N_23516,N_23318,N_23173);
nand U23517 (N_23517,N_23326,N_23349);
and U23518 (N_23518,N_23159,N_23340);
or U23519 (N_23519,N_23308,N_23127);
xor U23520 (N_23520,N_23286,N_23181);
xor U23521 (N_23521,N_23105,N_23186);
or U23522 (N_23522,N_23171,N_23370);
nor U23523 (N_23523,N_23353,N_23187);
nor U23524 (N_23524,N_23219,N_23348);
nor U23525 (N_23525,N_23160,N_23112);
nand U23526 (N_23526,N_23361,N_23297);
nand U23527 (N_23527,N_23396,N_23294);
and U23528 (N_23528,N_23277,N_23184);
nand U23529 (N_23529,N_23212,N_23293);
and U23530 (N_23530,N_23397,N_23262);
nor U23531 (N_23531,N_23225,N_23332);
nand U23532 (N_23532,N_23239,N_23120);
and U23533 (N_23533,N_23327,N_23175);
and U23534 (N_23534,N_23183,N_23136);
nand U23535 (N_23535,N_23128,N_23355);
xor U23536 (N_23536,N_23233,N_23130);
or U23537 (N_23537,N_23275,N_23364);
xor U23538 (N_23538,N_23110,N_23139);
nor U23539 (N_23539,N_23324,N_23298);
xnor U23540 (N_23540,N_23285,N_23236);
nor U23541 (N_23541,N_23200,N_23182);
xor U23542 (N_23542,N_23248,N_23303);
xor U23543 (N_23543,N_23344,N_23166);
and U23544 (N_23544,N_23272,N_23235);
nand U23545 (N_23545,N_23174,N_23115);
xor U23546 (N_23546,N_23196,N_23374);
and U23547 (N_23547,N_23280,N_23345);
nor U23548 (N_23548,N_23379,N_23185);
and U23549 (N_23549,N_23273,N_23144);
or U23550 (N_23550,N_23265,N_23252);
nor U23551 (N_23551,N_23245,N_23158);
or U23552 (N_23552,N_23367,N_23222);
nor U23553 (N_23553,N_23189,N_23131);
xnor U23554 (N_23554,N_23149,N_23392);
and U23555 (N_23555,N_23235,N_23337);
nor U23556 (N_23556,N_23134,N_23205);
nor U23557 (N_23557,N_23152,N_23115);
and U23558 (N_23558,N_23220,N_23200);
and U23559 (N_23559,N_23367,N_23331);
or U23560 (N_23560,N_23329,N_23189);
nor U23561 (N_23561,N_23311,N_23324);
nand U23562 (N_23562,N_23268,N_23314);
or U23563 (N_23563,N_23390,N_23265);
nor U23564 (N_23564,N_23223,N_23171);
xor U23565 (N_23565,N_23367,N_23274);
xnor U23566 (N_23566,N_23328,N_23325);
nor U23567 (N_23567,N_23307,N_23117);
nor U23568 (N_23568,N_23277,N_23175);
nand U23569 (N_23569,N_23376,N_23274);
nand U23570 (N_23570,N_23145,N_23284);
nor U23571 (N_23571,N_23230,N_23272);
xor U23572 (N_23572,N_23155,N_23141);
nor U23573 (N_23573,N_23264,N_23332);
xor U23574 (N_23574,N_23228,N_23121);
nand U23575 (N_23575,N_23253,N_23321);
xor U23576 (N_23576,N_23236,N_23159);
or U23577 (N_23577,N_23175,N_23270);
or U23578 (N_23578,N_23277,N_23205);
and U23579 (N_23579,N_23189,N_23351);
and U23580 (N_23580,N_23136,N_23308);
nand U23581 (N_23581,N_23362,N_23317);
or U23582 (N_23582,N_23101,N_23325);
or U23583 (N_23583,N_23294,N_23218);
xnor U23584 (N_23584,N_23129,N_23119);
and U23585 (N_23585,N_23355,N_23321);
and U23586 (N_23586,N_23158,N_23241);
xnor U23587 (N_23587,N_23364,N_23251);
nor U23588 (N_23588,N_23368,N_23255);
or U23589 (N_23589,N_23350,N_23242);
nand U23590 (N_23590,N_23233,N_23333);
or U23591 (N_23591,N_23235,N_23232);
or U23592 (N_23592,N_23138,N_23392);
xor U23593 (N_23593,N_23255,N_23145);
nor U23594 (N_23594,N_23346,N_23128);
nand U23595 (N_23595,N_23150,N_23188);
nor U23596 (N_23596,N_23254,N_23334);
xnor U23597 (N_23597,N_23126,N_23202);
xor U23598 (N_23598,N_23208,N_23132);
and U23599 (N_23599,N_23198,N_23170);
nor U23600 (N_23600,N_23303,N_23305);
and U23601 (N_23601,N_23286,N_23379);
or U23602 (N_23602,N_23355,N_23169);
xnor U23603 (N_23603,N_23191,N_23398);
or U23604 (N_23604,N_23101,N_23160);
nand U23605 (N_23605,N_23138,N_23117);
nand U23606 (N_23606,N_23359,N_23326);
nor U23607 (N_23607,N_23296,N_23316);
nand U23608 (N_23608,N_23192,N_23277);
and U23609 (N_23609,N_23200,N_23164);
nand U23610 (N_23610,N_23204,N_23180);
and U23611 (N_23611,N_23278,N_23114);
xnor U23612 (N_23612,N_23314,N_23191);
nand U23613 (N_23613,N_23231,N_23372);
nand U23614 (N_23614,N_23155,N_23154);
nand U23615 (N_23615,N_23275,N_23220);
xor U23616 (N_23616,N_23268,N_23187);
or U23617 (N_23617,N_23358,N_23275);
nor U23618 (N_23618,N_23195,N_23379);
or U23619 (N_23619,N_23291,N_23397);
or U23620 (N_23620,N_23148,N_23334);
xor U23621 (N_23621,N_23107,N_23268);
nand U23622 (N_23622,N_23239,N_23166);
or U23623 (N_23623,N_23385,N_23278);
nor U23624 (N_23624,N_23204,N_23221);
and U23625 (N_23625,N_23171,N_23102);
nand U23626 (N_23626,N_23232,N_23152);
xor U23627 (N_23627,N_23305,N_23341);
nand U23628 (N_23628,N_23355,N_23245);
xor U23629 (N_23629,N_23153,N_23358);
nand U23630 (N_23630,N_23309,N_23356);
nor U23631 (N_23631,N_23115,N_23172);
nor U23632 (N_23632,N_23368,N_23307);
xor U23633 (N_23633,N_23211,N_23292);
or U23634 (N_23634,N_23368,N_23183);
nand U23635 (N_23635,N_23233,N_23278);
nor U23636 (N_23636,N_23383,N_23319);
and U23637 (N_23637,N_23249,N_23245);
xnor U23638 (N_23638,N_23315,N_23119);
nand U23639 (N_23639,N_23255,N_23310);
or U23640 (N_23640,N_23262,N_23336);
nor U23641 (N_23641,N_23151,N_23318);
nand U23642 (N_23642,N_23323,N_23159);
and U23643 (N_23643,N_23105,N_23333);
xor U23644 (N_23644,N_23353,N_23343);
nor U23645 (N_23645,N_23257,N_23357);
nor U23646 (N_23646,N_23307,N_23318);
nand U23647 (N_23647,N_23125,N_23131);
xor U23648 (N_23648,N_23367,N_23357);
and U23649 (N_23649,N_23237,N_23120);
or U23650 (N_23650,N_23192,N_23135);
xnor U23651 (N_23651,N_23281,N_23273);
xor U23652 (N_23652,N_23327,N_23341);
nand U23653 (N_23653,N_23186,N_23332);
nor U23654 (N_23654,N_23278,N_23309);
xnor U23655 (N_23655,N_23317,N_23287);
or U23656 (N_23656,N_23343,N_23135);
and U23657 (N_23657,N_23276,N_23131);
nand U23658 (N_23658,N_23121,N_23365);
nor U23659 (N_23659,N_23318,N_23340);
and U23660 (N_23660,N_23225,N_23263);
nand U23661 (N_23661,N_23370,N_23344);
and U23662 (N_23662,N_23248,N_23302);
or U23663 (N_23663,N_23298,N_23230);
xor U23664 (N_23664,N_23235,N_23255);
nand U23665 (N_23665,N_23267,N_23241);
or U23666 (N_23666,N_23369,N_23167);
nor U23667 (N_23667,N_23190,N_23392);
and U23668 (N_23668,N_23376,N_23303);
xnor U23669 (N_23669,N_23298,N_23257);
nor U23670 (N_23670,N_23383,N_23274);
nand U23671 (N_23671,N_23300,N_23156);
nand U23672 (N_23672,N_23200,N_23234);
nand U23673 (N_23673,N_23280,N_23110);
nand U23674 (N_23674,N_23303,N_23363);
or U23675 (N_23675,N_23318,N_23273);
nor U23676 (N_23676,N_23178,N_23194);
or U23677 (N_23677,N_23262,N_23392);
nor U23678 (N_23678,N_23160,N_23237);
xnor U23679 (N_23679,N_23129,N_23272);
nand U23680 (N_23680,N_23317,N_23226);
nor U23681 (N_23681,N_23131,N_23104);
nand U23682 (N_23682,N_23116,N_23154);
nor U23683 (N_23683,N_23337,N_23325);
and U23684 (N_23684,N_23322,N_23106);
nor U23685 (N_23685,N_23209,N_23261);
nand U23686 (N_23686,N_23128,N_23213);
xnor U23687 (N_23687,N_23194,N_23267);
xnor U23688 (N_23688,N_23317,N_23329);
and U23689 (N_23689,N_23117,N_23190);
and U23690 (N_23690,N_23129,N_23110);
nor U23691 (N_23691,N_23303,N_23290);
xor U23692 (N_23692,N_23246,N_23161);
nand U23693 (N_23693,N_23199,N_23161);
or U23694 (N_23694,N_23269,N_23260);
or U23695 (N_23695,N_23370,N_23346);
and U23696 (N_23696,N_23232,N_23272);
xor U23697 (N_23697,N_23367,N_23363);
or U23698 (N_23698,N_23307,N_23197);
xor U23699 (N_23699,N_23197,N_23396);
nand U23700 (N_23700,N_23654,N_23693);
and U23701 (N_23701,N_23673,N_23537);
xnor U23702 (N_23702,N_23425,N_23414);
or U23703 (N_23703,N_23439,N_23564);
nor U23704 (N_23704,N_23600,N_23554);
nand U23705 (N_23705,N_23543,N_23659);
and U23706 (N_23706,N_23490,N_23410);
nor U23707 (N_23707,N_23502,N_23677);
xor U23708 (N_23708,N_23456,N_23506);
xnor U23709 (N_23709,N_23696,N_23463);
or U23710 (N_23710,N_23427,N_23687);
and U23711 (N_23711,N_23531,N_23408);
or U23712 (N_23712,N_23624,N_23460);
and U23713 (N_23713,N_23539,N_23405);
and U23714 (N_23714,N_23694,N_23528);
nand U23715 (N_23715,N_23446,N_23606);
and U23716 (N_23716,N_23524,N_23611);
or U23717 (N_23717,N_23499,N_23598);
nand U23718 (N_23718,N_23535,N_23665);
xor U23719 (N_23719,N_23594,N_23447);
xor U23720 (N_23720,N_23587,N_23457);
nor U23721 (N_23721,N_23464,N_23678);
nand U23722 (N_23722,N_23666,N_23503);
nor U23723 (N_23723,N_23417,N_23581);
nand U23724 (N_23724,N_23510,N_23612);
or U23725 (N_23725,N_23605,N_23400);
nand U23726 (N_23726,N_23650,N_23567);
xnor U23727 (N_23727,N_23527,N_23618);
or U23728 (N_23728,N_23538,N_23630);
or U23729 (N_23729,N_23631,N_23416);
nand U23730 (N_23730,N_23652,N_23511);
and U23731 (N_23731,N_23488,N_23476);
xnor U23732 (N_23732,N_23435,N_23608);
and U23733 (N_23733,N_23613,N_23471);
xor U23734 (N_23734,N_23485,N_23625);
nor U23735 (N_23735,N_23566,N_23619);
xor U23736 (N_23736,N_23420,N_23640);
and U23737 (N_23737,N_23402,N_23655);
or U23738 (N_23738,N_23526,N_23532);
or U23739 (N_23739,N_23604,N_23575);
and U23740 (N_23740,N_23418,N_23513);
nor U23741 (N_23741,N_23621,N_23592);
nor U23742 (N_23742,N_23628,N_23649);
nor U23743 (N_23743,N_23498,N_23449);
nand U23744 (N_23744,N_23582,N_23656);
or U23745 (N_23745,N_23648,N_23634);
xnor U23746 (N_23746,N_23660,N_23595);
nor U23747 (N_23747,N_23579,N_23597);
xor U23748 (N_23748,N_23433,N_23686);
or U23749 (N_23749,N_23679,N_23627);
and U23750 (N_23750,N_23413,N_23590);
xnor U23751 (N_23751,N_23637,N_23521);
nor U23752 (N_23752,N_23657,N_23469);
xor U23753 (N_23753,N_23541,N_23475);
xor U23754 (N_23754,N_23481,N_23482);
nand U23755 (N_23755,N_23635,N_23601);
nand U23756 (N_23756,N_23504,N_23542);
nor U23757 (N_23757,N_23599,N_23681);
and U23758 (N_23758,N_23699,N_23536);
or U23759 (N_23759,N_23478,N_23629);
xor U23760 (N_23760,N_23695,N_23658);
nand U23761 (N_23761,N_23403,N_23492);
or U23762 (N_23762,N_23517,N_23563);
nand U23763 (N_23763,N_23530,N_23662);
nand U23764 (N_23764,N_23495,N_23443);
or U23765 (N_23765,N_23429,N_23451);
and U23766 (N_23766,N_23642,N_23448);
xor U23767 (N_23767,N_23620,N_23646);
and U23768 (N_23768,N_23486,N_23578);
and U23769 (N_23769,N_23419,N_23663);
and U23770 (N_23770,N_23500,N_23515);
nor U23771 (N_23771,N_23674,N_23467);
nor U23772 (N_23772,N_23638,N_23562);
nor U23773 (N_23773,N_23483,N_23548);
nor U23774 (N_23774,N_23442,N_23661);
xor U23775 (N_23775,N_23491,N_23430);
and U23776 (N_23776,N_23445,N_23438);
nand U23777 (N_23777,N_23428,N_23639);
nand U23778 (N_23778,N_23576,N_23422);
or U23779 (N_23779,N_23603,N_23667);
and U23780 (N_23780,N_23470,N_23653);
nor U23781 (N_23781,N_23450,N_23669);
or U23782 (N_23782,N_23523,N_23549);
nand U23783 (N_23783,N_23568,N_23558);
and U23784 (N_23784,N_23487,N_23676);
nor U23785 (N_23785,N_23584,N_23509);
and U23786 (N_23786,N_23671,N_23545);
nor U23787 (N_23787,N_23680,N_23643);
or U23788 (N_23788,N_23547,N_23645);
nand U23789 (N_23789,N_23670,N_23689);
nor U23790 (N_23790,N_23574,N_23609);
xnor U23791 (N_23791,N_23633,N_23489);
nor U23792 (N_23792,N_23551,N_23626);
or U23793 (N_23793,N_23493,N_23426);
xor U23794 (N_23794,N_23685,N_23644);
and U23795 (N_23795,N_23434,N_23474);
nor U23796 (N_23796,N_23623,N_23572);
and U23797 (N_23797,N_23580,N_23550);
nor U23798 (N_23798,N_23610,N_23691);
and U23799 (N_23799,N_23465,N_23440);
nand U23800 (N_23800,N_23570,N_23494);
nor U23801 (N_23801,N_23675,N_23444);
or U23802 (N_23802,N_23454,N_23404);
nand U23803 (N_23803,N_23571,N_23466);
and U23804 (N_23804,N_23533,N_23505);
nand U23805 (N_23805,N_23622,N_23602);
or U23806 (N_23806,N_23692,N_23552);
or U23807 (N_23807,N_23682,N_23589);
xor U23808 (N_23808,N_23688,N_23651);
or U23809 (N_23809,N_23501,N_23529);
nor U23810 (N_23810,N_23591,N_23424);
nand U23811 (N_23811,N_23569,N_23401);
or U23812 (N_23812,N_23432,N_23617);
or U23813 (N_23813,N_23596,N_23462);
nor U23814 (N_23814,N_23525,N_23518);
and U23815 (N_23815,N_23468,N_23672);
nand U23816 (N_23816,N_23593,N_23522);
xnor U23817 (N_23817,N_23647,N_23556);
xor U23818 (N_23818,N_23409,N_23477);
and U23819 (N_23819,N_23508,N_23514);
and U23820 (N_23820,N_23683,N_23480);
and U23821 (N_23821,N_23455,N_23684);
nor U23822 (N_23822,N_23421,N_23586);
and U23823 (N_23823,N_23516,N_23544);
xnor U23824 (N_23824,N_23473,N_23565);
nand U23825 (N_23825,N_23507,N_23472);
nor U23826 (N_23826,N_23583,N_23540);
or U23827 (N_23827,N_23664,N_23577);
xor U23828 (N_23828,N_23546,N_23461);
and U23829 (N_23829,N_23406,N_23697);
nand U23830 (N_23830,N_23555,N_23561);
or U23831 (N_23831,N_23479,N_23559);
nor U23832 (N_23832,N_23557,N_23453);
and U23833 (N_23833,N_23534,N_23512);
or U23834 (N_23834,N_23436,N_23458);
and U23835 (N_23835,N_23698,N_23616);
nand U23836 (N_23836,N_23411,N_23573);
nor U23837 (N_23837,N_23407,N_23641);
and U23838 (N_23838,N_23519,N_23459);
nand U23839 (N_23839,N_23585,N_23437);
nand U23840 (N_23840,N_23520,N_23632);
xnor U23841 (N_23841,N_23452,N_23560);
nor U23842 (N_23842,N_23412,N_23553);
nor U23843 (N_23843,N_23588,N_23636);
or U23844 (N_23844,N_23615,N_23431);
and U23845 (N_23845,N_23496,N_23614);
or U23846 (N_23846,N_23484,N_23668);
and U23847 (N_23847,N_23497,N_23607);
xnor U23848 (N_23848,N_23690,N_23415);
and U23849 (N_23849,N_23441,N_23423);
nand U23850 (N_23850,N_23555,N_23616);
xnor U23851 (N_23851,N_23578,N_23625);
and U23852 (N_23852,N_23603,N_23400);
and U23853 (N_23853,N_23415,N_23597);
nor U23854 (N_23854,N_23467,N_23648);
xor U23855 (N_23855,N_23689,N_23439);
nand U23856 (N_23856,N_23548,N_23640);
nand U23857 (N_23857,N_23504,N_23627);
or U23858 (N_23858,N_23694,N_23649);
nand U23859 (N_23859,N_23620,N_23537);
nand U23860 (N_23860,N_23617,N_23423);
and U23861 (N_23861,N_23692,N_23653);
nor U23862 (N_23862,N_23555,N_23582);
and U23863 (N_23863,N_23636,N_23477);
nor U23864 (N_23864,N_23697,N_23404);
or U23865 (N_23865,N_23515,N_23437);
nor U23866 (N_23866,N_23546,N_23620);
or U23867 (N_23867,N_23681,N_23522);
xnor U23868 (N_23868,N_23458,N_23565);
xor U23869 (N_23869,N_23439,N_23413);
nor U23870 (N_23870,N_23642,N_23452);
xnor U23871 (N_23871,N_23454,N_23650);
nor U23872 (N_23872,N_23401,N_23411);
nor U23873 (N_23873,N_23699,N_23652);
nand U23874 (N_23874,N_23486,N_23527);
nand U23875 (N_23875,N_23565,N_23456);
nand U23876 (N_23876,N_23523,N_23476);
nand U23877 (N_23877,N_23625,N_23604);
or U23878 (N_23878,N_23444,N_23424);
nor U23879 (N_23879,N_23575,N_23569);
nand U23880 (N_23880,N_23569,N_23439);
or U23881 (N_23881,N_23605,N_23527);
or U23882 (N_23882,N_23595,N_23674);
nor U23883 (N_23883,N_23417,N_23490);
nand U23884 (N_23884,N_23564,N_23630);
nor U23885 (N_23885,N_23617,N_23604);
nand U23886 (N_23886,N_23685,N_23562);
and U23887 (N_23887,N_23438,N_23613);
nor U23888 (N_23888,N_23514,N_23638);
and U23889 (N_23889,N_23407,N_23629);
nand U23890 (N_23890,N_23516,N_23417);
or U23891 (N_23891,N_23683,N_23509);
xor U23892 (N_23892,N_23587,N_23450);
nand U23893 (N_23893,N_23653,N_23583);
xor U23894 (N_23894,N_23673,N_23568);
or U23895 (N_23895,N_23474,N_23471);
xor U23896 (N_23896,N_23542,N_23679);
nor U23897 (N_23897,N_23597,N_23539);
or U23898 (N_23898,N_23475,N_23451);
nor U23899 (N_23899,N_23693,N_23696);
and U23900 (N_23900,N_23408,N_23464);
nand U23901 (N_23901,N_23573,N_23406);
xor U23902 (N_23902,N_23563,N_23419);
xnor U23903 (N_23903,N_23458,N_23442);
and U23904 (N_23904,N_23531,N_23505);
and U23905 (N_23905,N_23556,N_23600);
and U23906 (N_23906,N_23490,N_23441);
nand U23907 (N_23907,N_23654,N_23565);
xor U23908 (N_23908,N_23532,N_23553);
nand U23909 (N_23909,N_23699,N_23640);
nor U23910 (N_23910,N_23613,N_23665);
nand U23911 (N_23911,N_23554,N_23582);
nand U23912 (N_23912,N_23437,N_23494);
nand U23913 (N_23913,N_23526,N_23607);
nand U23914 (N_23914,N_23502,N_23685);
and U23915 (N_23915,N_23474,N_23570);
and U23916 (N_23916,N_23630,N_23504);
and U23917 (N_23917,N_23448,N_23630);
xor U23918 (N_23918,N_23552,N_23549);
nor U23919 (N_23919,N_23623,N_23439);
and U23920 (N_23920,N_23472,N_23510);
or U23921 (N_23921,N_23533,N_23687);
and U23922 (N_23922,N_23503,N_23605);
or U23923 (N_23923,N_23679,N_23698);
nand U23924 (N_23924,N_23684,N_23570);
and U23925 (N_23925,N_23475,N_23539);
nand U23926 (N_23926,N_23488,N_23553);
or U23927 (N_23927,N_23639,N_23637);
or U23928 (N_23928,N_23496,N_23651);
or U23929 (N_23929,N_23693,N_23670);
nor U23930 (N_23930,N_23498,N_23650);
nand U23931 (N_23931,N_23695,N_23521);
or U23932 (N_23932,N_23459,N_23457);
or U23933 (N_23933,N_23409,N_23429);
and U23934 (N_23934,N_23612,N_23461);
and U23935 (N_23935,N_23472,N_23435);
nor U23936 (N_23936,N_23501,N_23488);
xor U23937 (N_23937,N_23532,N_23537);
and U23938 (N_23938,N_23589,N_23585);
or U23939 (N_23939,N_23616,N_23474);
xor U23940 (N_23940,N_23470,N_23433);
nor U23941 (N_23941,N_23610,N_23422);
xor U23942 (N_23942,N_23610,N_23603);
and U23943 (N_23943,N_23479,N_23505);
nand U23944 (N_23944,N_23634,N_23478);
xor U23945 (N_23945,N_23567,N_23479);
xor U23946 (N_23946,N_23519,N_23404);
nand U23947 (N_23947,N_23598,N_23464);
and U23948 (N_23948,N_23445,N_23491);
nor U23949 (N_23949,N_23439,N_23561);
xor U23950 (N_23950,N_23529,N_23663);
nand U23951 (N_23951,N_23629,N_23487);
and U23952 (N_23952,N_23631,N_23429);
nand U23953 (N_23953,N_23486,N_23541);
xor U23954 (N_23954,N_23558,N_23442);
nor U23955 (N_23955,N_23420,N_23402);
nand U23956 (N_23956,N_23590,N_23469);
and U23957 (N_23957,N_23408,N_23559);
nor U23958 (N_23958,N_23420,N_23526);
and U23959 (N_23959,N_23601,N_23495);
and U23960 (N_23960,N_23492,N_23526);
nor U23961 (N_23961,N_23619,N_23559);
xor U23962 (N_23962,N_23415,N_23684);
nand U23963 (N_23963,N_23558,N_23549);
xor U23964 (N_23964,N_23567,N_23563);
and U23965 (N_23965,N_23612,N_23489);
nand U23966 (N_23966,N_23581,N_23502);
and U23967 (N_23967,N_23487,N_23444);
nand U23968 (N_23968,N_23462,N_23595);
nor U23969 (N_23969,N_23548,N_23460);
xor U23970 (N_23970,N_23495,N_23532);
and U23971 (N_23971,N_23484,N_23435);
nand U23972 (N_23972,N_23550,N_23566);
and U23973 (N_23973,N_23682,N_23501);
and U23974 (N_23974,N_23595,N_23598);
nor U23975 (N_23975,N_23413,N_23461);
xor U23976 (N_23976,N_23500,N_23467);
nor U23977 (N_23977,N_23592,N_23406);
xnor U23978 (N_23978,N_23423,N_23573);
xnor U23979 (N_23979,N_23527,N_23593);
xor U23980 (N_23980,N_23631,N_23459);
nor U23981 (N_23981,N_23482,N_23623);
and U23982 (N_23982,N_23627,N_23543);
nor U23983 (N_23983,N_23479,N_23605);
or U23984 (N_23984,N_23511,N_23422);
and U23985 (N_23985,N_23693,N_23448);
xor U23986 (N_23986,N_23591,N_23695);
and U23987 (N_23987,N_23592,N_23566);
xnor U23988 (N_23988,N_23505,N_23621);
nand U23989 (N_23989,N_23424,N_23484);
nor U23990 (N_23990,N_23543,N_23561);
xnor U23991 (N_23991,N_23590,N_23490);
xnor U23992 (N_23992,N_23646,N_23618);
and U23993 (N_23993,N_23537,N_23622);
or U23994 (N_23994,N_23537,N_23434);
or U23995 (N_23995,N_23412,N_23521);
or U23996 (N_23996,N_23597,N_23591);
nor U23997 (N_23997,N_23654,N_23420);
nor U23998 (N_23998,N_23615,N_23620);
or U23999 (N_23999,N_23493,N_23574);
or U24000 (N_24000,N_23746,N_23789);
nor U24001 (N_24001,N_23794,N_23736);
and U24002 (N_24002,N_23713,N_23804);
or U24003 (N_24003,N_23731,N_23823);
xor U24004 (N_24004,N_23830,N_23962);
and U24005 (N_24005,N_23898,N_23972);
nand U24006 (N_24006,N_23956,N_23841);
and U24007 (N_24007,N_23880,N_23910);
or U24008 (N_24008,N_23905,N_23990);
nor U24009 (N_24009,N_23983,N_23803);
and U24010 (N_24010,N_23978,N_23901);
xnor U24011 (N_24011,N_23927,N_23848);
xor U24012 (N_24012,N_23745,N_23963);
nor U24013 (N_24013,N_23870,N_23786);
nand U24014 (N_24014,N_23872,N_23931);
and U24015 (N_24015,N_23752,N_23776);
or U24016 (N_24016,N_23950,N_23806);
xor U24017 (N_24017,N_23784,N_23826);
nor U24018 (N_24018,N_23850,N_23976);
xnor U24019 (N_24019,N_23829,N_23721);
nor U24020 (N_24020,N_23722,N_23857);
or U24021 (N_24021,N_23986,N_23723);
xnor U24022 (N_24022,N_23926,N_23838);
and U24023 (N_24023,N_23997,N_23903);
nor U24024 (N_24024,N_23874,N_23795);
nor U24025 (N_24025,N_23840,N_23788);
nor U24026 (N_24026,N_23989,N_23727);
nand U24027 (N_24027,N_23937,N_23980);
nor U24028 (N_24028,N_23994,N_23856);
or U24029 (N_24029,N_23875,N_23991);
nand U24030 (N_24030,N_23711,N_23894);
nand U24031 (N_24031,N_23720,N_23953);
nand U24032 (N_24032,N_23779,N_23923);
nor U24033 (N_24033,N_23750,N_23887);
nand U24034 (N_24034,N_23900,N_23807);
xnor U24035 (N_24035,N_23966,N_23724);
nand U24036 (N_24036,N_23932,N_23888);
nand U24037 (N_24037,N_23785,N_23941);
or U24038 (N_24038,N_23877,N_23917);
and U24039 (N_24039,N_23704,N_23867);
nor U24040 (N_24040,N_23868,N_23973);
nand U24041 (N_24041,N_23984,N_23952);
or U24042 (N_24042,N_23708,N_23717);
nor U24043 (N_24043,N_23732,N_23974);
xnor U24044 (N_24044,N_23812,N_23992);
or U24045 (N_24045,N_23706,N_23774);
or U24046 (N_24046,N_23749,N_23742);
or U24047 (N_24047,N_23998,N_23781);
nor U24048 (N_24048,N_23897,N_23833);
and U24049 (N_24049,N_23861,N_23819);
or U24050 (N_24050,N_23863,N_23949);
and U24051 (N_24051,N_23911,N_23712);
or U24052 (N_24052,N_23800,N_23922);
nand U24053 (N_24053,N_23822,N_23768);
and U24054 (N_24054,N_23882,N_23961);
nor U24055 (N_24055,N_23959,N_23718);
or U24056 (N_24056,N_23960,N_23754);
or U24057 (N_24057,N_23797,N_23946);
xnor U24058 (N_24058,N_23738,N_23740);
nor U24059 (N_24059,N_23790,N_23940);
xnor U24060 (N_24060,N_23993,N_23860);
nand U24061 (N_24061,N_23853,N_23824);
nand U24062 (N_24062,N_23747,N_23753);
and U24063 (N_24063,N_23787,N_23739);
nand U24064 (N_24064,N_23930,N_23816);
xnor U24065 (N_24065,N_23866,N_23879);
and U24066 (N_24066,N_23808,N_23700);
or U24067 (N_24067,N_23726,N_23999);
xnor U24068 (N_24068,N_23773,N_23968);
xor U24069 (N_24069,N_23743,N_23777);
or U24070 (N_24070,N_23873,N_23884);
xor U24071 (N_24071,N_23886,N_23728);
and U24072 (N_24072,N_23707,N_23762);
nor U24073 (N_24073,N_23907,N_23835);
xnor U24074 (N_24074,N_23764,N_23985);
nand U24075 (N_24075,N_23844,N_23958);
nor U24076 (N_24076,N_23802,N_23895);
nor U24077 (N_24077,N_23855,N_23703);
nor U24078 (N_24078,N_23915,N_23847);
xor U24079 (N_24079,N_23805,N_23842);
or U24080 (N_24080,N_23741,N_23821);
nand U24081 (N_24081,N_23859,N_23965);
or U24082 (N_24082,N_23995,N_23815);
nand U24083 (N_24083,N_23893,N_23921);
and U24084 (N_24084,N_23920,N_23818);
nor U24085 (N_24085,N_23827,N_23935);
or U24086 (N_24086,N_23828,N_23970);
xnor U24087 (N_24087,N_23846,N_23878);
and U24088 (N_24088,N_23782,N_23792);
and U24089 (N_24089,N_23996,N_23889);
or U24090 (N_24090,N_23843,N_23948);
and U24091 (N_24091,N_23979,N_23928);
xor U24092 (N_24092,N_23801,N_23714);
nand U24093 (N_24093,N_23765,N_23769);
nand U24094 (N_24094,N_23793,N_23730);
nor U24095 (N_24095,N_23876,N_23988);
nand U24096 (N_24096,N_23817,N_23854);
xnor U24097 (N_24097,N_23982,N_23869);
nor U24098 (N_24098,N_23918,N_23933);
nor U24099 (N_24099,N_23904,N_23820);
nor U24100 (N_24100,N_23947,N_23929);
xnor U24101 (N_24101,N_23852,N_23758);
or U24102 (N_24102,N_23734,N_23913);
xor U24103 (N_24103,N_23836,N_23957);
or U24104 (N_24104,N_23881,N_23906);
nand U24105 (N_24105,N_23759,N_23810);
xnor U24106 (N_24106,N_23755,N_23813);
and U24107 (N_24107,N_23936,N_23916);
or U24108 (N_24108,N_23967,N_23899);
nand U24109 (N_24109,N_23751,N_23891);
and U24110 (N_24110,N_23981,N_23778);
nand U24111 (N_24111,N_23825,N_23709);
or U24112 (N_24112,N_23902,N_23744);
and U24113 (N_24113,N_23766,N_23851);
nor U24114 (N_24114,N_23939,N_23925);
or U24115 (N_24115,N_23733,N_23885);
and U24116 (N_24116,N_23890,N_23954);
nand U24117 (N_24117,N_23969,N_23938);
or U24118 (N_24118,N_23710,N_23791);
or U24119 (N_24119,N_23832,N_23705);
nand U24120 (N_24120,N_23767,N_23799);
xor U24121 (N_24121,N_23763,N_23845);
xor U24122 (N_24122,N_23761,N_23735);
or U24123 (N_24123,N_23912,N_23770);
nand U24124 (N_24124,N_23862,N_23971);
nor U24125 (N_24125,N_23896,N_23849);
nand U24126 (N_24126,N_23837,N_23871);
or U24127 (N_24127,N_23858,N_23955);
and U24128 (N_24128,N_23748,N_23864);
xnor U24129 (N_24129,N_23919,N_23944);
nand U24130 (N_24130,N_23839,N_23783);
nor U24131 (N_24131,N_23977,N_23987);
and U24132 (N_24132,N_23892,N_23934);
or U24133 (N_24133,N_23809,N_23942);
and U24134 (N_24134,N_23831,N_23865);
xor U24135 (N_24135,N_23914,N_23737);
nand U24136 (N_24136,N_23951,N_23909);
xnor U24137 (N_24137,N_23796,N_23756);
nor U24138 (N_24138,N_23760,N_23814);
nor U24139 (N_24139,N_23924,N_23775);
and U24140 (N_24140,N_23729,N_23701);
or U24141 (N_24141,N_23883,N_23943);
and U24142 (N_24142,N_23975,N_23702);
and U24143 (N_24143,N_23771,N_23834);
or U24144 (N_24144,N_23715,N_23908);
nor U24145 (N_24145,N_23964,N_23945);
or U24146 (N_24146,N_23725,N_23772);
nand U24147 (N_24147,N_23811,N_23716);
nand U24148 (N_24148,N_23757,N_23798);
nor U24149 (N_24149,N_23780,N_23719);
nand U24150 (N_24150,N_23901,N_23951);
and U24151 (N_24151,N_23955,N_23838);
nor U24152 (N_24152,N_23893,N_23856);
or U24153 (N_24153,N_23925,N_23799);
or U24154 (N_24154,N_23836,N_23928);
nor U24155 (N_24155,N_23726,N_23918);
nor U24156 (N_24156,N_23999,N_23793);
and U24157 (N_24157,N_23768,N_23780);
xnor U24158 (N_24158,N_23930,N_23935);
xor U24159 (N_24159,N_23741,N_23969);
or U24160 (N_24160,N_23824,N_23768);
xnor U24161 (N_24161,N_23953,N_23829);
nor U24162 (N_24162,N_23722,N_23975);
and U24163 (N_24163,N_23769,N_23813);
xor U24164 (N_24164,N_23949,N_23832);
nor U24165 (N_24165,N_23762,N_23801);
and U24166 (N_24166,N_23885,N_23717);
or U24167 (N_24167,N_23817,N_23720);
xor U24168 (N_24168,N_23878,N_23998);
nor U24169 (N_24169,N_23702,N_23735);
and U24170 (N_24170,N_23778,N_23781);
and U24171 (N_24171,N_23702,N_23800);
xnor U24172 (N_24172,N_23844,N_23893);
or U24173 (N_24173,N_23830,N_23763);
xnor U24174 (N_24174,N_23798,N_23801);
or U24175 (N_24175,N_23978,N_23872);
nor U24176 (N_24176,N_23734,N_23725);
or U24177 (N_24177,N_23984,N_23796);
nor U24178 (N_24178,N_23896,N_23893);
or U24179 (N_24179,N_23969,N_23874);
nand U24180 (N_24180,N_23968,N_23992);
nand U24181 (N_24181,N_23969,N_23899);
xor U24182 (N_24182,N_23817,N_23809);
nand U24183 (N_24183,N_23751,N_23707);
nor U24184 (N_24184,N_23980,N_23710);
nor U24185 (N_24185,N_23717,N_23928);
xor U24186 (N_24186,N_23798,N_23959);
and U24187 (N_24187,N_23916,N_23802);
xnor U24188 (N_24188,N_23786,N_23841);
xnor U24189 (N_24189,N_23897,N_23799);
nor U24190 (N_24190,N_23813,N_23914);
nor U24191 (N_24191,N_23753,N_23854);
nand U24192 (N_24192,N_23757,N_23933);
or U24193 (N_24193,N_23770,N_23937);
and U24194 (N_24194,N_23838,N_23903);
nor U24195 (N_24195,N_23944,N_23766);
and U24196 (N_24196,N_23801,N_23833);
nand U24197 (N_24197,N_23947,N_23970);
nand U24198 (N_24198,N_23967,N_23861);
nor U24199 (N_24199,N_23862,N_23718);
nor U24200 (N_24200,N_23905,N_23776);
and U24201 (N_24201,N_23927,N_23878);
xor U24202 (N_24202,N_23960,N_23859);
xnor U24203 (N_24203,N_23827,N_23924);
nand U24204 (N_24204,N_23826,N_23847);
nand U24205 (N_24205,N_23718,N_23908);
nand U24206 (N_24206,N_23967,N_23944);
and U24207 (N_24207,N_23785,N_23780);
xor U24208 (N_24208,N_23783,N_23981);
and U24209 (N_24209,N_23965,N_23745);
nor U24210 (N_24210,N_23724,N_23806);
or U24211 (N_24211,N_23994,N_23986);
nor U24212 (N_24212,N_23898,N_23893);
or U24213 (N_24213,N_23841,N_23914);
xnor U24214 (N_24214,N_23937,N_23752);
nand U24215 (N_24215,N_23751,N_23899);
xor U24216 (N_24216,N_23761,N_23936);
and U24217 (N_24217,N_23998,N_23977);
nor U24218 (N_24218,N_23809,N_23834);
and U24219 (N_24219,N_23872,N_23999);
nand U24220 (N_24220,N_23789,N_23720);
nand U24221 (N_24221,N_23974,N_23707);
xnor U24222 (N_24222,N_23834,N_23887);
xor U24223 (N_24223,N_23721,N_23928);
nand U24224 (N_24224,N_23882,N_23907);
nor U24225 (N_24225,N_23999,N_23879);
and U24226 (N_24226,N_23821,N_23921);
or U24227 (N_24227,N_23942,N_23742);
xor U24228 (N_24228,N_23866,N_23801);
or U24229 (N_24229,N_23722,N_23956);
xor U24230 (N_24230,N_23994,N_23823);
nand U24231 (N_24231,N_23866,N_23913);
and U24232 (N_24232,N_23723,N_23751);
and U24233 (N_24233,N_23753,N_23935);
nand U24234 (N_24234,N_23995,N_23766);
or U24235 (N_24235,N_23966,N_23851);
and U24236 (N_24236,N_23800,N_23810);
and U24237 (N_24237,N_23984,N_23829);
xnor U24238 (N_24238,N_23955,N_23729);
xnor U24239 (N_24239,N_23887,N_23974);
nand U24240 (N_24240,N_23877,N_23989);
or U24241 (N_24241,N_23846,N_23898);
and U24242 (N_24242,N_23913,N_23794);
and U24243 (N_24243,N_23888,N_23907);
nand U24244 (N_24244,N_23727,N_23706);
nor U24245 (N_24245,N_23755,N_23758);
nand U24246 (N_24246,N_23969,N_23925);
nor U24247 (N_24247,N_23737,N_23817);
or U24248 (N_24248,N_23899,N_23877);
and U24249 (N_24249,N_23977,N_23999);
xnor U24250 (N_24250,N_23746,N_23998);
or U24251 (N_24251,N_23811,N_23879);
and U24252 (N_24252,N_23886,N_23777);
xor U24253 (N_24253,N_23850,N_23802);
xor U24254 (N_24254,N_23930,N_23856);
nand U24255 (N_24255,N_23992,N_23866);
nand U24256 (N_24256,N_23915,N_23791);
and U24257 (N_24257,N_23992,N_23916);
xnor U24258 (N_24258,N_23960,N_23913);
or U24259 (N_24259,N_23845,N_23796);
or U24260 (N_24260,N_23998,N_23824);
xor U24261 (N_24261,N_23900,N_23797);
xor U24262 (N_24262,N_23916,N_23949);
nor U24263 (N_24263,N_23817,N_23897);
nand U24264 (N_24264,N_23883,N_23790);
and U24265 (N_24265,N_23922,N_23929);
nand U24266 (N_24266,N_23823,N_23891);
nand U24267 (N_24267,N_23763,N_23917);
and U24268 (N_24268,N_23802,N_23756);
xnor U24269 (N_24269,N_23960,N_23999);
and U24270 (N_24270,N_23906,N_23747);
nand U24271 (N_24271,N_23919,N_23818);
nor U24272 (N_24272,N_23803,N_23856);
nor U24273 (N_24273,N_23794,N_23744);
nand U24274 (N_24274,N_23962,N_23968);
xnor U24275 (N_24275,N_23725,N_23702);
nor U24276 (N_24276,N_23889,N_23944);
nand U24277 (N_24277,N_23852,N_23821);
and U24278 (N_24278,N_23966,N_23921);
xnor U24279 (N_24279,N_23942,N_23916);
xnor U24280 (N_24280,N_23743,N_23834);
and U24281 (N_24281,N_23745,N_23952);
and U24282 (N_24282,N_23800,N_23774);
and U24283 (N_24283,N_23805,N_23711);
or U24284 (N_24284,N_23815,N_23941);
or U24285 (N_24285,N_23989,N_23805);
nand U24286 (N_24286,N_23935,N_23787);
nor U24287 (N_24287,N_23955,N_23793);
nor U24288 (N_24288,N_23984,N_23950);
xor U24289 (N_24289,N_23790,N_23784);
or U24290 (N_24290,N_23976,N_23994);
xor U24291 (N_24291,N_23957,N_23837);
or U24292 (N_24292,N_23881,N_23747);
and U24293 (N_24293,N_23965,N_23860);
nand U24294 (N_24294,N_23832,N_23704);
nor U24295 (N_24295,N_23814,N_23883);
or U24296 (N_24296,N_23909,N_23714);
or U24297 (N_24297,N_23762,N_23894);
or U24298 (N_24298,N_23865,N_23828);
and U24299 (N_24299,N_23855,N_23976);
nor U24300 (N_24300,N_24236,N_24177);
nand U24301 (N_24301,N_24213,N_24124);
nand U24302 (N_24302,N_24030,N_24243);
xor U24303 (N_24303,N_24281,N_24076);
xor U24304 (N_24304,N_24110,N_24275);
xor U24305 (N_24305,N_24205,N_24077);
and U24306 (N_24306,N_24268,N_24218);
xnor U24307 (N_24307,N_24078,N_24014);
and U24308 (N_24308,N_24228,N_24021);
and U24309 (N_24309,N_24016,N_24181);
or U24310 (N_24310,N_24237,N_24135);
xnor U24311 (N_24311,N_24131,N_24020);
and U24312 (N_24312,N_24035,N_24234);
and U24313 (N_24313,N_24250,N_24291);
nor U24314 (N_24314,N_24132,N_24231);
xor U24315 (N_24315,N_24107,N_24264);
and U24316 (N_24316,N_24062,N_24039);
xor U24317 (N_24317,N_24157,N_24003);
nand U24318 (N_24318,N_24079,N_24024);
and U24319 (N_24319,N_24261,N_24258);
and U24320 (N_24320,N_24084,N_24155);
xor U24321 (N_24321,N_24278,N_24125);
nand U24322 (N_24322,N_24004,N_24096);
or U24323 (N_24323,N_24115,N_24064);
and U24324 (N_24324,N_24019,N_24173);
xnor U24325 (N_24325,N_24253,N_24288);
or U24326 (N_24326,N_24012,N_24127);
or U24327 (N_24327,N_24036,N_24182);
nor U24328 (N_24328,N_24289,N_24190);
nor U24329 (N_24329,N_24145,N_24153);
or U24330 (N_24330,N_24252,N_24154);
and U24331 (N_24331,N_24010,N_24255);
or U24332 (N_24332,N_24242,N_24071);
xor U24333 (N_24333,N_24058,N_24294);
or U24334 (N_24334,N_24249,N_24054);
and U24335 (N_24335,N_24279,N_24098);
or U24336 (N_24336,N_24007,N_24144);
nor U24337 (N_24337,N_24290,N_24065);
and U24338 (N_24338,N_24285,N_24284);
nand U24339 (N_24339,N_24299,N_24056);
xnor U24340 (N_24340,N_24262,N_24101);
and U24341 (N_24341,N_24171,N_24260);
or U24342 (N_24342,N_24158,N_24027);
or U24343 (N_24343,N_24130,N_24106);
nand U24344 (N_24344,N_24123,N_24043);
or U24345 (N_24345,N_24227,N_24109);
xnor U24346 (N_24346,N_24188,N_24025);
or U24347 (N_24347,N_24201,N_24067);
nand U24348 (N_24348,N_24099,N_24179);
nand U24349 (N_24349,N_24093,N_24169);
and U24350 (N_24350,N_24295,N_24053);
nor U24351 (N_24351,N_24142,N_24298);
xnor U24352 (N_24352,N_24229,N_24164);
or U24353 (N_24353,N_24051,N_24167);
nand U24354 (N_24354,N_24176,N_24293);
nand U24355 (N_24355,N_24046,N_24152);
and U24356 (N_24356,N_24097,N_24208);
nand U24357 (N_24357,N_24070,N_24066);
or U24358 (N_24358,N_24042,N_24159);
nor U24359 (N_24359,N_24011,N_24015);
xor U24360 (N_24360,N_24283,N_24002);
xor U24361 (N_24361,N_24033,N_24270);
or U24362 (N_24362,N_24001,N_24138);
xor U24363 (N_24363,N_24189,N_24055);
and U24364 (N_24364,N_24089,N_24112);
xnor U24365 (N_24365,N_24140,N_24120);
nor U24366 (N_24366,N_24220,N_24150);
xor U24367 (N_24367,N_24251,N_24184);
nand U24368 (N_24368,N_24221,N_24224);
nor U24369 (N_24369,N_24160,N_24063);
and U24370 (N_24370,N_24017,N_24119);
or U24371 (N_24371,N_24246,N_24257);
xor U24372 (N_24372,N_24126,N_24094);
or U24373 (N_24373,N_24200,N_24223);
xor U24374 (N_24374,N_24045,N_24018);
or U24375 (N_24375,N_24100,N_24122);
and U24376 (N_24376,N_24280,N_24128);
or U24377 (N_24377,N_24183,N_24296);
nand U24378 (N_24378,N_24207,N_24068);
and U24379 (N_24379,N_24116,N_24286);
nor U24380 (N_24380,N_24256,N_24180);
xor U24381 (N_24381,N_24090,N_24248);
nand U24382 (N_24382,N_24031,N_24187);
and U24383 (N_24383,N_24166,N_24037);
nand U24384 (N_24384,N_24165,N_24163);
xor U24385 (N_24385,N_24297,N_24102);
or U24386 (N_24386,N_24271,N_24195);
and U24387 (N_24387,N_24212,N_24210);
or U24388 (N_24388,N_24060,N_24244);
or U24389 (N_24389,N_24121,N_24108);
nand U24390 (N_24390,N_24083,N_24240);
nand U24391 (N_24391,N_24292,N_24215);
nand U24392 (N_24392,N_24272,N_24129);
nand U24393 (N_24393,N_24052,N_24203);
or U24394 (N_24394,N_24172,N_24174);
xor U24395 (N_24395,N_24194,N_24222);
nor U24396 (N_24396,N_24023,N_24117);
nand U24397 (N_24397,N_24082,N_24239);
nand U24398 (N_24398,N_24143,N_24162);
nand U24399 (N_24399,N_24191,N_24081);
or U24400 (N_24400,N_24086,N_24134);
xnor U24401 (N_24401,N_24137,N_24266);
or U24402 (N_24402,N_24273,N_24057);
xor U24403 (N_24403,N_24032,N_24059);
nand U24404 (N_24404,N_24217,N_24006);
or U24405 (N_24405,N_24075,N_24232);
nor U24406 (N_24406,N_24034,N_24050);
and U24407 (N_24407,N_24274,N_24147);
or U24408 (N_24408,N_24204,N_24139);
or U24409 (N_24409,N_24193,N_24041);
or U24410 (N_24410,N_24196,N_24247);
nor U24411 (N_24411,N_24091,N_24073);
nand U24412 (N_24412,N_24209,N_24022);
xnor U24413 (N_24413,N_24185,N_24047);
nor U24414 (N_24414,N_24175,N_24005);
nor U24415 (N_24415,N_24214,N_24061);
nand U24416 (N_24416,N_24267,N_24265);
or U24417 (N_24417,N_24085,N_24199);
xnor U24418 (N_24418,N_24044,N_24048);
or U24419 (N_24419,N_24254,N_24105);
nand U24420 (N_24420,N_24168,N_24235);
nand U24421 (N_24421,N_24269,N_24111);
xor U24422 (N_24422,N_24026,N_24088);
nor U24423 (N_24423,N_24211,N_24241);
nor U24424 (N_24424,N_24136,N_24287);
xor U24425 (N_24425,N_24259,N_24113);
xor U24426 (N_24426,N_24149,N_24049);
nor U24427 (N_24427,N_24146,N_24141);
and U24428 (N_24428,N_24118,N_24186);
or U24429 (N_24429,N_24080,N_24103);
nand U24430 (N_24430,N_24156,N_24277);
or U24431 (N_24431,N_24038,N_24161);
and U24432 (N_24432,N_24013,N_24238);
xor U24433 (N_24433,N_24170,N_24233);
nand U24434 (N_24434,N_24151,N_24072);
xnor U24435 (N_24435,N_24219,N_24009);
and U24436 (N_24436,N_24092,N_24074);
xor U24437 (N_24437,N_24008,N_24198);
or U24438 (N_24438,N_24148,N_24202);
nand U24439 (N_24439,N_24028,N_24197);
and U24440 (N_24440,N_24263,N_24282);
or U24441 (N_24441,N_24245,N_24087);
nor U24442 (N_24442,N_24069,N_24095);
xnor U24443 (N_24443,N_24276,N_24104);
or U24444 (N_24444,N_24192,N_24216);
and U24445 (N_24445,N_24178,N_24040);
nand U24446 (N_24446,N_24206,N_24114);
nand U24447 (N_24447,N_24029,N_24230);
nand U24448 (N_24448,N_24225,N_24133);
xor U24449 (N_24449,N_24000,N_24226);
or U24450 (N_24450,N_24245,N_24235);
and U24451 (N_24451,N_24182,N_24227);
nor U24452 (N_24452,N_24061,N_24268);
and U24453 (N_24453,N_24082,N_24107);
or U24454 (N_24454,N_24079,N_24262);
nand U24455 (N_24455,N_24201,N_24155);
and U24456 (N_24456,N_24115,N_24257);
or U24457 (N_24457,N_24247,N_24013);
nor U24458 (N_24458,N_24194,N_24154);
nor U24459 (N_24459,N_24274,N_24162);
and U24460 (N_24460,N_24117,N_24115);
nor U24461 (N_24461,N_24120,N_24296);
and U24462 (N_24462,N_24172,N_24119);
or U24463 (N_24463,N_24061,N_24022);
xnor U24464 (N_24464,N_24174,N_24101);
xnor U24465 (N_24465,N_24100,N_24130);
nand U24466 (N_24466,N_24046,N_24067);
or U24467 (N_24467,N_24089,N_24059);
nor U24468 (N_24468,N_24088,N_24262);
nand U24469 (N_24469,N_24125,N_24140);
and U24470 (N_24470,N_24158,N_24260);
xor U24471 (N_24471,N_24122,N_24139);
nor U24472 (N_24472,N_24279,N_24172);
nand U24473 (N_24473,N_24078,N_24279);
xor U24474 (N_24474,N_24275,N_24182);
or U24475 (N_24475,N_24059,N_24141);
nand U24476 (N_24476,N_24108,N_24094);
and U24477 (N_24477,N_24276,N_24132);
or U24478 (N_24478,N_24266,N_24125);
nand U24479 (N_24479,N_24011,N_24055);
nor U24480 (N_24480,N_24055,N_24187);
and U24481 (N_24481,N_24164,N_24127);
nor U24482 (N_24482,N_24159,N_24185);
xnor U24483 (N_24483,N_24133,N_24141);
or U24484 (N_24484,N_24190,N_24007);
and U24485 (N_24485,N_24122,N_24248);
xnor U24486 (N_24486,N_24222,N_24109);
and U24487 (N_24487,N_24066,N_24166);
and U24488 (N_24488,N_24116,N_24191);
or U24489 (N_24489,N_24249,N_24176);
nor U24490 (N_24490,N_24108,N_24095);
or U24491 (N_24491,N_24280,N_24222);
xor U24492 (N_24492,N_24211,N_24178);
or U24493 (N_24493,N_24261,N_24297);
and U24494 (N_24494,N_24269,N_24093);
and U24495 (N_24495,N_24190,N_24006);
xor U24496 (N_24496,N_24139,N_24261);
nor U24497 (N_24497,N_24030,N_24202);
xor U24498 (N_24498,N_24291,N_24292);
nor U24499 (N_24499,N_24228,N_24152);
nand U24500 (N_24500,N_24056,N_24178);
xnor U24501 (N_24501,N_24265,N_24061);
xnor U24502 (N_24502,N_24037,N_24246);
xor U24503 (N_24503,N_24160,N_24279);
or U24504 (N_24504,N_24090,N_24072);
or U24505 (N_24505,N_24271,N_24253);
xnor U24506 (N_24506,N_24160,N_24035);
xnor U24507 (N_24507,N_24217,N_24248);
and U24508 (N_24508,N_24275,N_24200);
or U24509 (N_24509,N_24030,N_24162);
nand U24510 (N_24510,N_24163,N_24035);
nor U24511 (N_24511,N_24227,N_24185);
or U24512 (N_24512,N_24177,N_24191);
xor U24513 (N_24513,N_24143,N_24198);
or U24514 (N_24514,N_24211,N_24056);
nor U24515 (N_24515,N_24207,N_24190);
or U24516 (N_24516,N_24095,N_24043);
nor U24517 (N_24517,N_24202,N_24162);
and U24518 (N_24518,N_24298,N_24214);
or U24519 (N_24519,N_24095,N_24212);
and U24520 (N_24520,N_24010,N_24009);
xor U24521 (N_24521,N_24159,N_24125);
or U24522 (N_24522,N_24009,N_24088);
xor U24523 (N_24523,N_24016,N_24298);
nor U24524 (N_24524,N_24298,N_24219);
xor U24525 (N_24525,N_24216,N_24183);
nor U24526 (N_24526,N_24026,N_24090);
nand U24527 (N_24527,N_24159,N_24173);
or U24528 (N_24528,N_24195,N_24040);
nand U24529 (N_24529,N_24215,N_24159);
nand U24530 (N_24530,N_24103,N_24185);
nor U24531 (N_24531,N_24129,N_24285);
and U24532 (N_24532,N_24142,N_24104);
and U24533 (N_24533,N_24260,N_24179);
and U24534 (N_24534,N_24273,N_24115);
xor U24535 (N_24535,N_24101,N_24069);
nand U24536 (N_24536,N_24191,N_24215);
and U24537 (N_24537,N_24028,N_24042);
nand U24538 (N_24538,N_24256,N_24214);
nor U24539 (N_24539,N_24286,N_24173);
nand U24540 (N_24540,N_24127,N_24280);
or U24541 (N_24541,N_24216,N_24271);
and U24542 (N_24542,N_24258,N_24107);
or U24543 (N_24543,N_24091,N_24268);
xor U24544 (N_24544,N_24097,N_24258);
and U24545 (N_24545,N_24276,N_24232);
nor U24546 (N_24546,N_24261,N_24029);
and U24547 (N_24547,N_24246,N_24209);
and U24548 (N_24548,N_24259,N_24262);
and U24549 (N_24549,N_24298,N_24136);
or U24550 (N_24550,N_24022,N_24152);
or U24551 (N_24551,N_24153,N_24206);
nor U24552 (N_24552,N_24065,N_24244);
and U24553 (N_24553,N_24034,N_24230);
xnor U24554 (N_24554,N_24220,N_24088);
nor U24555 (N_24555,N_24037,N_24282);
nor U24556 (N_24556,N_24279,N_24134);
nand U24557 (N_24557,N_24182,N_24012);
xor U24558 (N_24558,N_24244,N_24032);
nor U24559 (N_24559,N_24170,N_24092);
or U24560 (N_24560,N_24168,N_24187);
nand U24561 (N_24561,N_24123,N_24034);
nor U24562 (N_24562,N_24265,N_24225);
nor U24563 (N_24563,N_24216,N_24012);
and U24564 (N_24564,N_24230,N_24185);
nand U24565 (N_24565,N_24059,N_24248);
or U24566 (N_24566,N_24123,N_24018);
xor U24567 (N_24567,N_24038,N_24140);
or U24568 (N_24568,N_24089,N_24132);
nor U24569 (N_24569,N_24033,N_24213);
xor U24570 (N_24570,N_24298,N_24127);
and U24571 (N_24571,N_24015,N_24215);
nor U24572 (N_24572,N_24240,N_24131);
xor U24573 (N_24573,N_24131,N_24206);
nand U24574 (N_24574,N_24110,N_24166);
or U24575 (N_24575,N_24264,N_24143);
and U24576 (N_24576,N_24282,N_24120);
or U24577 (N_24577,N_24142,N_24011);
xnor U24578 (N_24578,N_24152,N_24113);
nor U24579 (N_24579,N_24235,N_24008);
and U24580 (N_24580,N_24293,N_24216);
and U24581 (N_24581,N_24014,N_24214);
or U24582 (N_24582,N_24185,N_24157);
or U24583 (N_24583,N_24278,N_24120);
xnor U24584 (N_24584,N_24217,N_24014);
nand U24585 (N_24585,N_24119,N_24249);
and U24586 (N_24586,N_24258,N_24067);
and U24587 (N_24587,N_24166,N_24078);
nor U24588 (N_24588,N_24279,N_24206);
and U24589 (N_24589,N_24276,N_24241);
and U24590 (N_24590,N_24157,N_24194);
or U24591 (N_24591,N_24127,N_24150);
and U24592 (N_24592,N_24071,N_24077);
and U24593 (N_24593,N_24266,N_24278);
and U24594 (N_24594,N_24286,N_24104);
nand U24595 (N_24595,N_24048,N_24208);
and U24596 (N_24596,N_24191,N_24054);
nand U24597 (N_24597,N_24261,N_24269);
or U24598 (N_24598,N_24297,N_24255);
nand U24599 (N_24599,N_24068,N_24193);
or U24600 (N_24600,N_24451,N_24492);
nand U24601 (N_24601,N_24402,N_24468);
or U24602 (N_24602,N_24343,N_24311);
xor U24603 (N_24603,N_24308,N_24458);
or U24604 (N_24604,N_24326,N_24426);
xor U24605 (N_24605,N_24578,N_24482);
xor U24606 (N_24606,N_24556,N_24309);
and U24607 (N_24607,N_24407,N_24406);
nor U24608 (N_24608,N_24507,N_24584);
nor U24609 (N_24609,N_24307,N_24412);
nand U24610 (N_24610,N_24488,N_24440);
nand U24611 (N_24611,N_24504,N_24521);
nand U24612 (N_24612,N_24337,N_24471);
nor U24613 (N_24613,N_24486,N_24405);
xor U24614 (N_24614,N_24335,N_24457);
nor U24615 (N_24615,N_24439,N_24494);
and U24616 (N_24616,N_24347,N_24385);
nand U24617 (N_24617,N_24590,N_24354);
nand U24618 (N_24618,N_24365,N_24339);
nand U24619 (N_24619,N_24522,N_24340);
or U24620 (N_24620,N_24540,N_24384);
xnor U24621 (N_24621,N_24364,N_24532);
nand U24622 (N_24622,N_24397,N_24596);
or U24623 (N_24623,N_24304,N_24353);
nand U24624 (N_24624,N_24533,N_24403);
nand U24625 (N_24625,N_24387,N_24376);
nor U24626 (N_24626,N_24508,N_24489);
and U24627 (N_24627,N_24324,N_24310);
xnor U24628 (N_24628,N_24421,N_24470);
xor U24629 (N_24629,N_24573,N_24373);
nand U24630 (N_24630,N_24417,N_24534);
and U24631 (N_24631,N_24328,N_24467);
and U24632 (N_24632,N_24483,N_24448);
or U24633 (N_24633,N_24375,N_24429);
xnor U24634 (N_24634,N_24513,N_24502);
or U24635 (N_24635,N_24475,N_24436);
and U24636 (N_24636,N_24520,N_24314);
nand U24637 (N_24637,N_24333,N_24581);
nor U24638 (N_24638,N_24322,N_24320);
nand U24639 (N_24639,N_24415,N_24390);
and U24640 (N_24640,N_24577,N_24349);
xnor U24641 (N_24641,N_24554,N_24505);
nor U24642 (N_24642,N_24549,N_24386);
nor U24643 (N_24643,N_24569,N_24449);
nor U24644 (N_24644,N_24346,N_24591);
xnor U24645 (N_24645,N_24465,N_24543);
nor U24646 (N_24646,N_24352,N_24416);
nand U24647 (N_24647,N_24538,N_24332);
nor U24648 (N_24648,N_24418,N_24338);
nor U24649 (N_24649,N_24321,N_24301);
nor U24650 (N_24650,N_24455,N_24372);
and U24651 (N_24651,N_24366,N_24481);
or U24652 (N_24652,N_24317,N_24472);
xnor U24653 (N_24653,N_24565,N_24500);
and U24654 (N_24654,N_24551,N_24348);
xor U24655 (N_24655,N_24497,N_24393);
and U24656 (N_24656,N_24531,N_24318);
and U24657 (N_24657,N_24329,N_24312);
nor U24658 (N_24658,N_24535,N_24562);
and U24659 (N_24659,N_24527,N_24359);
or U24660 (N_24660,N_24460,N_24441);
nor U24661 (N_24661,N_24341,N_24501);
nor U24662 (N_24662,N_24392,N_24526);
nor U24663 (N_24663,N_24443,N_24399);
and U24664 (N_24664,N_24388,N_24345);
or U24665 (N_24665,N_24401,N_24360);
nand U24666 (N_24666,N_24567,N_24325);
nor U24667 (N_24667,N_24453,N_24529);
nor U24668 (N_24668,N_24411,N_24599);
nand U24669 (N_24669,N_24377,N_24424);
nor U24670 (N_24670,N_24342,N_24514);
xnor U24671 (N_24671,N_24461,N_24408);
and U24672 (N_24672,N_24552,N_24331);
nand U24673 (N_24673,N_24469,N_24548);
xnor U24674 (N_24674,N_24383,N_24400);
and U24675 (N_24675,N_24357,N_24541);
or U24676 (N_24676,N_24560,N_24445);
nand U24677 (N_24677,N_24546,N_24545);
nand U24678 (N_24678,N_24595,N_24361);
nand U24679 (N_24679,N_24477,N_24442);
nand U24680 (N_24680,N_24517,N_24355);
xor U24681 (N_24681,N_24446,N_24413);
xnor U24682 (N_24682,N_24300,N_24369);
xor U24683 (N_24683,N_24447,N_24575);
nor U24684 (N_24684,N_24409,N_24438);
xor U24685 (N_24685,N_24553,N_24572);
and U24686 (N_24686,N_24585,N_24557);
and U24687 (N_24687,N_24589,N_24323);
nor U24688 (N_24688,N_24499,N_24420);
and U24689 (N_24689,N_24370,N_24398);
nand U24690 (N_24690,N_24450,N_24380);
or U24691 (N_24691,N_24493,N_24559);
and U24692 (N_24692,N_24586,N_24485);
or U24693 (N_24693,N_24305,N_24498);
and U24694 (N_24694,N_24381,N_24433);
nor U24695 (N_24695,N_24484,N_24480);
nand U24696 (N_24696,N_24583,N_24593);
xor U24697 (N_24697,N_24563,N_24422);
and U24698 (N_24698,N_24368,N_24452);
or U24699 (N_24699,N_24555,N_24313);
and U24700 (N_24700,N_24479,N_24378);
nor U24701 (N_24701,N_24454,N_24568);
nor U24702 (N_24702,N_24435,N_24444);
nand U24703 (N_24703,N_24512,N_24537);
nand U24704 (N_24704,N_24358,N_24503);
nand U24705 (N_24705,N_24404,N_24395);
and U24706 (N_24706,N_24428,N_24410);
or U24707 (N_24707,N_24389,N_24356);
and U24708 (N_24708,N_24434,N_24574);
nand U24709 (N_24709,N_24487,N_24518);
and U24710 (N_24710,N_24437,N_24476);
and U24711 (N_24711,N_24334,N_24597);
nand U24712 (N_24712,N_24536,N_24425);
or U24713 (N_24713,N_24466,N_24363);
and U24714 (N_24714,N_24371,N_24506);
xor U24715 (N_24715,N_24509,N_24580);
nand U24716 (N_24716,N_24511,N_24432);
xnor U24717 (N_24717,N_24316,N_24523);
xor U24718 (N_24718,N_24516,N_24391);
xnor U24719 (N_24719,N_24464,N_24315);
and U24720 (N_24720,N_24561,N_24544);
xor U24721 (N_24721,N_24592,N_24576);
nand U24722 (N_24722,N_24571,N_24374);
or U24723 (N_24723,N_24570,N_24528);
or U24724 (N_24724,N_24490,N_24495);
or U24725 (N_24725,N_24473,N_24564);
nor U24726 (N_24726,N_24558,N_24582);
or U24727 (N_24727,N_24456,N_24542);
and U24728 (N_24728,N_24427,N_24496);
and U24729 (N_24729,N_24382,N_24474);
and U24730 (N_24730,N_24414,N_24362);
or U24731 (N_24731,N_24594,N_24302);
xnor U24732 (N_24732,N_24587,N_24491);
xor U24733 (N_24733,N_24430,N_24367);
nor U24734 (N_24734,N_24588,N_24598);
nor U24735 (N_24735,N_24350,N_24396);
and U24736 (N_24736,N_24550,N_24566);
or U24737 (N_24737,N_24303,N_24394);
and U24738 (N_24738,N_24579,N_24327);
nor U24739 (N_24739,N_24319,N_24547);
nor U24740 (N_24740,N_24431,N_24423);
nor U24741 (N_24741,N_24510,N_24524);
xnor U24742 (N_24742,N_24419,N_24306);
nor U24743 (N_24743,N_24539,N_24344);
nor U24744 (N_24744,N_24462,N_24336);
or U24745 (N_24745,N_24519,N_24525);
nor U24746 (N_24746,N_24459,N_24330);
or U24747 (N_24747,N_24478,N_24515);
or U24748 (N_24748,N_24351,N_24530);
nor U24749 (N_24749,N_24463,N_24379);
and U24750 (N_24750,N_24339,N_24335);
xor U24751 (N_24751,N_24568,N_24440);
xnor U24752 (N_24752,N_24568,N_24333);
nor U24753 (N_24753,N_24393,N_24488);
and U24754 (N_24754,N_24344,N_24365);
nor U24755 (N_24755,N_24449,N_24589);
xor U24756 (N_24756,N_24463,N_24330);
nand U24757 (N_24757,N_24423,N_24529);
or U24758 (N_24758,N_24596,N_24417);
nand U24759 (N_24759,N_24513,N_24520);
xnor U24760 (N_24760,N_24321,N_24334);
and U24761 (N_24761,N_24560,N_24390);
or U24762 (N_24762,N_24550,N_24407);
xnor U24763 (N_24763,N_24461,N_24592);
or U24764 (N_24764,N_24321,N_24305);
nand U24765 (N_24765,N_24379,N_24360);
or U24766 (N_24766,N_24303,N_24440);
nand U24767 (N_24767,N_24329,N_24396);
xor U24768 (N_24768,N_24530,N_24572);
nor U24769 (N_24769,N_24311,N_24487);
xor U24770 (N_24770,N_24314,N_24391);
nand U24771 (N_24771,N_24598,N_24567);
or U24772 (N_24772,N_24550,N_24482);
or U24773 (N_24773,N_24557,N_24510);
nand U24774 (N_24774,N_24315,N_24312);
xor U24775 (N_24775,N_24302,N_24303);
xnor U24776 (N_24776,N_24320,N_24573);
nor U24777 (N_24777,N_24539,N_24374);
or U24778 (N_24778,N_24468,N_24368);
and U24779 (N_24779,N_24446,N_24420);
or U24780 (N_24780,N_24528,N_24554);
and U24781 (N_24781,N_24499,N_24427);
xor U24782 (N_24782,N_24472,N_24301);
xor U24783 (N_24783,N_24324,N_24549);
nor U24784 (N_24784,N_24516,N_24474);
or U24785 (N_24785,N_24561,N_24580);
and U24786 (N_24786,N_24409,N_24331);
nand U24787 (N_24787,N_24561,N_24340);
nand U24788 (N_24788,N_24422,N_24451);
or U24789 (N_24789,N_24369,N_24422);
xor U24790 (N_24790,N_24448,N_24471);
and U24791 (N_24791,N_24368,N_24458);
or U24792 (N_24792,N_24437,N_24508);
nand U24793 (N_24793,N_24447,N_24389);
nand U24794 (N_24794,N_24545,N_24481);
and U24795 (N_24795,N_24597,N_24463);
nor U24796 (N_24796,N_24317,N_24469);
and U24797 (N_24797,N_24555,N_24584);
nand U24798 (N_24798,N_24530,N_24391);
nor U24799 (N_24799,N_24590,N_24329);
or U24800 (N_24800,N_24301,N_24528);
xor U24801 (N_24801,N_24408,N_24413);
or U24802 (N_24802,N_24552,N_24393);
nor U24803 (N_24803,N_24482,N_24328);
xnor U24804 (N_24804,N_24391,N_24379);
xnor U24805 (N_24805,N_24384,N_24588);
and U24806 (N_24806,N_24412,N_24419);
nand U24807 (N_24807,N_24355,N_24319);
or U24808 (N_24808,N_24558,N_24407);
and U24809 (N_24809,N_24571,N_24522);
xor U24810 (N_24810,N_24424,N_24416);
nand U24811 (N_24811,N_24463,N_24517);
nor U24812 (N_24812,N_24458,N_24388);
and U24813 (N_24813,N_24523,N_24589);
nand U24814 (N_24814,N_24384,N_24476);
or U24815 (N_24815,N_24460,N_24582);
xnor U24816 (N_24816,N_24361,N_24577);
nor U24817 (N_24817,N_24554,N_24372);
nor U24818 (N_24818,N_24470,N_24390);
nand U24819 (N_24819,N_24549,N_24446);
nand U24820 (N_24820,N_24471,N_24580);
and U24821 (N_24821,N_24485,N_24446);
and U24822 (N_24822,N_24512,N_24538);
and U24823 (N_24823,N_24476,N_24387);
nor U24824 (N_24824,N_24457,N_24501);
or U24825 (N_24825,N_24551,N_24483);
xor U24826 (N_24826,N_24556,N_24469);
nor U24827 (N_24827,N_24470,N_24385);
nor U24828 (N_24828,N_24454,N_24456);
and U24829 (N_24829,N_24531,N_24441);
and U24830 (N_24830,N_24415,N_24540);
xor U24831 (N_24831,N_24428,N_24329);
nand U24832 (N_24832,N_24411,N_24508);
nor U24833 (N_24833,N_24467,N_24582);
or U24834 (N_24834,N_24515,N_24472);
xor U24835 (N_24835,N_24548,N_24400);
nor U24836 (N_24836,N_24590,N_24309);
nand U24837 (N_24837,N_24501,N_24514);
xor U24838 (N_24838,N_24457,N_24535);
nand U24839 (N_24839,N_24353,N_24423);
nor U24840 (N_24840,N_24407,N_24384);
nand U24841 (N_24841,N_24310,N_24521);
nand U24842 (N_24842,N_24595,N_24558);
nand U24843 (N_24843,N_24412,N_24327);
or U24844 (N_24844,N_24451,N_24513);
nor U24845 (N_24845,N_24441,N_24487);
xnor U24846 (N_24846,N_24525,N_24498);
nor U24847 (N_24847,N_24399,N_24547);
or U24848 (N_24848,N_24444,N_24581);
xor U24849 (N_24849,N_24493,N_24401);
or U24850 (N_24850,N_24521,N_24366);
and U24851 (N_24851,N_24348,N_24372);
nor U24852 (N_24852,N_24408,N_24354);
nor U24853 (N_24853,N_24364,N_24301);
nand U24854 (N_24854,N_24310,N_24517);
xnor U24855 (N_24855,N_24312,N_24583);
nor U24856 (N_24856,N_24334,N_24419);
nand U24857 (N_24857,N_24482,N_24469);
nor U24858 (N_24858,N_24444,N_24520);
xnor U24859 (N_24859,N_24592,N_24492);
nand U24860 (N_24860,N_24530,N_24347);
nor U24861 (N_24861,N_24393,N_24540);
and U24862 (N_24862,N_24557,N_24351);
or U24863 (N_24863,N_24597,N_24353);
nor U24864 (N_24864,N_24469,N_24593);
nor U24865 (N_24865,N_24355,N_24436);
or U24866 (N_24866,N_24537,N_24453);
and U24867 (N_24867,N_24330,N_24363);
and U24868 (N_24868,N_24380,N_24371);
or U24869 (N_24869,N_24457,N_24557);
nand U24870 (N_24870,N_24493,N_24504);
nand U24871 (N_24871,N_24585,N_24594);
nor U24872 (N_24872,N_24317,N_24594);
nor U24873 (N_24873,N_24390,N_24333);
nand U24874 (N_24874,N_24387,N_24544);
nand U24875 (N_24875,N_24349,N_24307);
nor U24876 (N_24876,N_24307,N_24444);
xnor U24877 (N_24877,N_24498,N_24330);
nand U24878 (N_24878,N_24395,N_24386);
nand U24879 (N_24879,N_24462,N_24494);
nor U24880 (N_24880,N_24409,N_24398);
or U24881 (N_24881,N_24432,N_24473);
or U24882 (N_24882,N_24443,N_24522);
and U24883 (N_24883,N_24337,N_24317);
or U24884 (N_24884,N_24359,N_24354);
or U24885 (N_24885,N_24408,N_24334);
nand U24886 (N_24886,N_24307,N_24375);
and U24887 (N_24887,N_24578,N_24462);
or U24888 (N_24888,N_24552,N_24597);
or U24889 (N_24889,N_24356,N_24503);
or U24890 (N_24890,N_24586,N_24518);
nand U24891 (N_24891,N_24598,N_24494);
nor U24892 (N_24892,N_24361,N_24344);
xor U24893 (N_24893,N_24578,N_24486);
or U24894 (N_24894,N_24467,N_24370);
nor U24895 (N_24895,N_24495,N_24361);
or U24896 (N_24896,N_24428,N_24588);
xor U24897 (N_24897,N_24504,N_24595);
nor U24898 (N_24898,N_24344,N_24553);
nand U24899 (N_24899,N_24455,N_24497);
nand U24900 (N_24900,N_24854,N_24747);
nor U24901 (N_24901,N_24651,N_24859);
or U24902 (N_24902,N_24807,N_24842);
nand U24903 (N_24903,N_24753,N_24796);
and U24904 (N_24904,N_24690,N_24660);
and U24905 (N_24905,N_24686,N_24869);
xor U24906 (N_24906,N_24888,N_24821);
and U24907 (N_24907,N_24832,N_24865);
nor U24908 (N_24908,N_24876,N_24727);
or U24909 (N_24909,N_24734,N_24799);
nor U24910 (N_24910,N_24801,N_24626);
xnor U24911 (N_24911,N_24836,N_24872);
nor U24912 (N_24912,N_24749,N_24856);
nor U24913 (N_24913,N_24630,N_24895);
nor U24914 (N_24914,N_24769,N_24713);
and U24915 (N_24915,N_24861,N_24719);
xnor U24916 (N_24916,N_24634,N_24815);
and U24917 (N_24917,N_24656,N_24826);
nand U24918 (N_24918,N_24616,N_24720);
nand U24919 (N_24919,N_24893,N_24863);
nor U24920 (N_24920,N_24709,N_24728);
nand U24921 (N_24921,N_24664,N_24890);
or U24922 (N_24922,N_24721,N_24676);
nand U24923 (N_24923,N_24857,N_24666);
or U24924 (N_24924,N_24804,N_24657);
xnor U24925 (N_24925,N_24897,N_24705);
nor U24926 (N_24926,N_24795,N_24603);
or U24927 (N_24927,N_24623,N_24862);
xor U24928 (N_24928,N_24787,N_24699);
or U24929 (N_24929,N_24885,N_24833);
nor U24930 (N_24930,N_24752,N_24622);
nor U24931 (N_24931,N_24881,N_24810);
or U24932 (N_24932,N_24655,N_24688);
and U24933 (N_24933,N_24687,N_24866);
and U24934 (N_24934,N_24673,N_24641);
nand U24935 (N_24935,N_24612,N_24695);
or U24936 (N_24936,N_24678,N_24868);
and U24937 (N_24937,N_24644,N_24786);
and U24938 (N_24938,N_24646,N_24736);
or U24939 (N_24939,N_24710,N_24723);
xor U24940 (N_24940,N_24889,N_24892);
xnor U24941 (N_24941,N_24700,N_24648);
and U24942 (N_24942,N_24702,N_24798);
xor U24943 (N_24943,N_24877,N_24886);
xor U24944 (N_24944,N_24611,N_24731);
nor U24945 (N_24945,N_24742,N_24671);
xor U24946 (N_24946,N_24697,N_24781);
nor U24947 (N_24947,N_24820,N_24670);
and U24948 (N_24948,N_24755,N_24779);
nor U24949 (N_24949,N_24640,N_24760);
nor U24950 (N_24950,N_24668,N_24629);
and U24951 (N_24951,N_24770,N_24793);
nand U24952 (N_24952,N_24610,N_24777);
nand U24953 (N_24953,N_24637,N_24733);
nand U24954 (N_24954,N_24726,N_24771);
or U24955 (N_24955,N_24732,N_24825);
xnor U24956 (N_24956,N_24649,N_24792);
xor U24957 (N_24957,N_24600,N_24766);
and U24958 (N_24958,N_24858,N_24812);
nand U24959 (N_24959,N_24669,N_24840);
nor U24960 (N_24960,N_24887,N_24844);
or U24961 (N_24961,N_24891,N_24797);
nor U24962 (N_24962,N_24837,N_24718);
nor U24963 (N_24963,N_24704,N_24808);
nor U24964 (N_24964,N_24794,N_24619);
xor U24965 (N_24965,N_24850,N_24659);
and U24966 (N_24966,N_24703,N_24636);
or U24967 (N_24967,N_24604,N_24739);
and U24968 (N_24968,N_24730,N_24849);
or U24969 (N_24969,N_24722,N_24838);
nor U24970 (N_24970,N_24682,N_24707);
xnor U24971 (N_24971,N_24624,N_24628);
xor U24972 (N_24972,N_24607,N_24767);
nand U24973 (N_24973,N_24784,N_24741);
nand U24974 (N_24974,N_24737,N_24652);
xnor U24975 (N_24975,N_24831,N_24803);
xnor U24976 (N_24976,N_24745,N_24693);
and U24977 (N_24977,N_24882,N_24675);
and U24978 (N_24978,N_24638,N_24661);
xor U24979 (N_24979,N_24608,N_24874);
xnor U24980 (N_24980,N_24658,N_24871);
nand U24981 (N_24981,N_24883,N_24650);
and U24982 (N_24982,N_24879,N_24653);
and U24983 (N_24983,N_24791,N_24667);
xor U24984 (N_24984,N_24692,N_24814);
and U24985 (N_24985,N_24751,N_24609);
nand U24986 (N_24986,N_24717,N_24824);
or U24987 (N_24987,N_24813,N_24899);
xnor U24988 (N_24988,N_24743,N_24870);
or U24989 (N_24989,N_24818,N_24768);
and U24990 (N_24990,N_24677,N_24756);
or U24991 (N_24991,N_24631,N_24715);
nor U24992 (N_24992,N_24694,N_24776);
nand U24993 (N_24993,N_24606,N_24816);
xnor U24994 (N_24994,N_24860,N_24613);
nand U24995 (N_24995,N_24746,N_24775);
nor U24996 (N_24996,N_24829,N_24763);
nor U24997 (N_24997,N_24851,N_24625);
xor U24998 (N_24998,N_24639,N_24839);
and U24999 (N_24999,N_24873,N_24685);
and U25000 (N_25000,N_24620,N_24642);
or U25001 (N_25001,N_24773,N_24696);
xnor U25002 (N_25002,N_24762,N_24841);
xor U25003 (N_25003,N_24615,N_24674);
or U25004 (N_25004,N_24701,N_24802);
nand U25005 (N_25005,N_24847,N_24698);
nor U25006 (N_25006,N_24822,N_24774);
or U25007 (N_25007,N_24627,N_24665);
nand U25008 (N_25008,N_24867,N_24789);
xor U25009 (N_25009,N_24601,N_24788);
and U25010 (N_25010,N_24617,N_24683);
xnor U25011 (N_25011,N_24689,N_24778);
nand U25012 (N_25012,N_24819,N_24602);
and U25013 (N_25013,N_24898,N_24855);
nor U25014 (N_25014,N_24830,N_24684);
or U25015 (N_25015,N_24706,N_24765);
xor U25016 (N_25016,N_24759,N_24754);
xnor U25017 (N_25017,N_24724,N_24852);
nor U25018 (N_25018,N_24894,N_24811);
and U25019 (N_25019,N_24785,N_24809);
xor U25020 (N_25020,N_24735,N_24663);
xor U25021 (N_25021,N_24843,N_24823);
and U25022 (N_25022,N_24672,N_24681);
nor U25023 (N_25023,N_24679,N_24647);
nor U25024 (N_25024,N_24878,N_24729);
nor U25025 (N_25025,N_24654,N_24662);
xor U25026 (N_25026,N_24632,N_24790);
nor U25027 (N_25027,N_24884,N_24848);
and U25028 (N_25028,N_24740,N_24880);
or U25029 (N_25029,N_24761,N_24783);
nor U25030 (N_25030,N_24645,N_24643);
nand U25031 (N_25031,N_24605,N_24757);
nand U25032 (N_25032,N_24714,N_24725);
nor U25033 (N_25033,N_24614,N_24875);
and U25034 (N_25034,N_24750,N_24817);
nor U25035 (N_25035,N_24800,N_24835);
and U25036 (N_25036,N_24708,N_24680);
xor U25037 (N_25037,N_24711,N_24712);
nor U25038 (N_25038,N_24758,N_24845);
or U25039 (N_25039,N_24764,N_24780);
or U25040 (N_25040,N_24744,N_24635);
xnor U25041 (N_25041,N_24772,N_24806);
nor U25042 (N_25042,N_24896,N_24846);
nor U25043 (N_25043,N_24716,N_24828);
or U25044 (N_25044,N_24633,N_24782);
nand U25045 (N_25045,N_24834,N_24827);
xor U25046 (N_25046,N_24621,N_24748);
nor U25047 (N_25047,N_24805,N_24853);
xnor U25048 (N_25048,N_24618,N_24738);
and U25049 (N_25049,N_24864,N_24691);
nor U25050 (N_25050,N_24774,N_24688);
or U25051 (N_25051,N_24820,N_24622);
and U25052 (N_25052,N_24777,N_24689);
xor U25053 (N_25053,N_24837,N_24807);
nand U25054 (N_25054,N_24795,N_24616);
nor U25055 (N_25055,N_24614,N_24698);
xnor U25056 (N_25056,N_24685,N_24837);
nor U25057 (N_25057,N_24612,N_24634);
and U25058 (N_25058,N_24898,N_24845);
and U25059 (N_25059,N_24685,N_24741);
nor U25060 (N_25060,N_24822,N_24659);
and U25061 (N_25061,N_24656,N_24807);
nor U25062 (N_25062,N_24806,N_24798);
and U25063 (N_25063,N_24647,N_24734);
nand U25064 (N_25064,N_24851,N_24760);
or U25065 (N_25065,N_24635,N_24672);
nor U25066 (N_25066,N_24821,N_24692);
nand U25067 (N_25067,N_24633,N_24891);
and U25068 (N_25068,N_24606,N_24724);
xnor U25069 (N_25069,N_24677,N_24673);
xor U25070 (N_25070,N_24880,N_24765);
nand U25071 (N_25071,N_24620,N_24838);
or U25072 (N_25072,N_24798,N_24773);
nor U25073 (N_25073,N_24650,N_24673);
nor U25074 (N_25074,N_24837,N_24746);
and U25075 (N_25075,N_24629,N_24798);
nand U25076 (N_25076,N_24825,N_24668);
nor U25077 (N_25077,N_24817,N_24818);
and U25078 (N_25078,N_24634,N_24825);
or U25079 (N_25079,N_24690,N_24735);
nand U25080 (N_25080,N_24835,N_24874);
xnor U25081 (N_25081,N_24615,N_24854);
nor U25082 (N_25082,N_24869,N_24655);
or U25083 (N_25083,N_24868,N_24770);
xor U25084 (N_25084,N_24755,N_24796);
nand U25085 (N_25085,N_24845,N_24806);
nand U25086 (N_25086,N_24670,N_24864);
and U25087 (N_25087,N_24872,N_24784);
nand U25088 (N_25088,N_24606,N_24878);
nor U25089 (N_25089,N_24655,N_24853);
nor U25090 (N_25090,N_24882,N_24650);
and U25091 (N_25091,N_24612,N_24730);
and U25092 (N_25092,N_24696,N_24737);
xor U25093 (N_25093,N_24865,N_24801);
and U25094 (N_25094,N_24605,N_24621);
xnor U25095 (N_25095,N_24779,N_24837);
nand U25096 (N_25096,N_24641,N_24605);
nor U25097 (N_25097,N_24782,N_24645);
xnor U25098 (N_25098,N_24796,N_24721);
xor U25099 (N_25099,N_24601,N_24817);
nor U25100 (N_25100,N_24847,N_24641);
and U25101 (N_25101,N_24834,N_24614);
or U25102 (N_25102,N_24731,N_24815);
nand U25103 (N_25103,N_24742,N_24854);
or U25104 (N_25104,N_24894,N_24883);
and U25105 (N_25105,N_24764,N_24846);
or U25106 (N_25106,N_24704,N_24830);
nand U25107 (N_25107,N_24781,N_24862);
or U25108 (N_25108,N_24746,N_24887);
and U25109 (N_25109,N_24768,N_24702);
nor U25110 (N_25110,N_24709,N_24781);
and U25111 (N_25111,N_24887,N_24777);
xor U25112 (N_25112,N_24766,N_24626);
nor U25113 (N_25113,N_24685,N_24733);
nand U25114 (N_25114,N_24759,N_24671);
and U25115 (N_25115,N_24796,N_24785);
nand U25116 (N_25116,N_24811,N_24606);
xnor U25117 (N_25117,N_24764,N_24614);
nand U25118 (N_25118,N_24772,N_24725);
and U25119 (N_25119,N_24655,N_24852);
and U25120 (N_25120,N_24679,N_24745);
xor U25121 (N_25121,N_24803,N_24637);
and U25122 (N_25122,N_24855,N_24857);
and U25123 (N_25123,N_24838,N_24806);
nor U25124 (N_25124,N_24619,N_24866);
or U25125 (N_25125,N_24870,N_24842);
nor U25126 (N_25126,N_24817,N_24641);
nand U25127 (N_25127,N_24753,N_24624);
nand U25128 (N_25128,N_24713,N_24858);
or U25129 (N_25129,N_24763,N_24750);
and U25130 (N_25130,N_24882,N_24810);
xnor U25131 (N_25131,N_24664,N_24753);
nand U25132 (N_25132,N_24652,N_24792);
xor U25133 (N_25133,N_24640,N_24685);
or U25134 (N_25134,N_24703,N_24695);
or U25135 (N_25135,N_24654,N_24890);
nand U25136 (N_25136,N_24689,N_24676);
xnor U25137 (N_25137,N_24817,N_24874);
or U25138 (N_25138,N_24795,N_24754);
nor U25139 (N_25139,N_24695,N_24801);
or U25140 (N_25140,N_24725,N_24885);
and U25141 (N_25141,N_24709,N_24685);
nor U25142 (N_25142,N_24726,N_24863);
xnor U25143 (N_25143,N_24775,N_24899);
and U25144 (N_25144,N_24896,N_24743);
xnor U25145 (N_25145,N_24736,N_24768);
and U25146 (N_25146,N_24722,N_24854);
or U25147 (N_25147,N_24870,N_24636);
nor U25148 (N_25148,N_24694,N_24816);
xor U25149 (N_25149,N_24718,N_24663);
or U25150 (N_25150,N_24862,N_24858);
nor U25151 (N_25151,N_24798,N_24899);
nand U25152 (N_25152,N_24793,N_24603);
xor U25153 (N_25153,N_24729,N_24627);
nor U25154 (N_25154,N_24781,N_24788);
xor U25155 (N_25155,N_24856,N_24809);
nand U25156 (N_25156,N_24676,N_24790);
nor U25157 (N_25157,N_24635,N_24790);
and U25158 (N_25158,N_24668,N_24622);
xnor U25159 (N_25159,N_24669,N_24751);
nor U25160 (N_25160,N_24851,N_24663);
nor U25161 (N_25161,N_24837,N_24847);
or U25162 (N_25162,N_24873,N_24684);
xor U25163 (N_25163,N_24620,N_24892);
or U25164 (N_25164,N_24889,N_24784);
or U25165 (N_25165,N_24889,N_24638);
and U25166 (N_25166,N_24708,N_24757);
xnor U25167 (N_25167,N_24777,N_24663);
or U25168 (N_25168,N_24602,N_24826);
nand U25169 (N_25169,N_24829,N_24677);
xor U25170 (N_25170,N_24795,N_24865);
or U25171 (N_25171,N_24823,N_24668);
and U25172 (N_25172,N_24820,N_24826);
or U25173 (N_25173,N_24636,N_24753);
or U25174 (N_25174,N_24680,N_24667);
or U25175 (N_25175,N_24761,N_24860);
xnor U25176 (N_25176,N_24778,N_24815);
and U25177 (N_25177,N_24803,N_24664);
and U25178 (N_25178,N_24757,N_24626);
nor U25179 (N_25179,N_24782,N_24676);
and U25180 (N_25180,N_24833,N_24814);
nor U25181 (N_25181,N_24789,N_24632);
xor U25182 (N_25182,N_24698,N_24822);
nor U25183 (N_25183,N_24775,N_24841);
and U25184 (N_25184,N_24804,N_24654);
xor U25185 (N_25185,N_24693,N_24760);
nor U25186 (N_25186,N_24887,N_24827);
and U25187 (N_25187,N_24785,N_24626);
and U25188 (N_25188,N_24849,N_24865);
nor U25189 (N_25189,N_24854,N_24662);
nand U25190 (N_25190,N_24739,N_24684);
xor U25191 (N_25191,N_24605,N_24611);
nand U25192 (N_25192,N_24763,N_24883);
and U25193 (N_25193,N_24754,N_24771);
or U25194 (N_25194,N_24748,N_24787);
nor U25195 (N_25195,N_24650,N_24819);
or U25196 (N_25196,N_24855,N_24737);
nand U25197 (N_25197,N_24692,N_24813);
nand U25198 (N_25198,N_24717,N_24749);
nand U25199 (N_25199,N_24737,N_24742);
nor U25200 (N_25200,N_25130,N_25108);
or U25201 (N_25201,N_25049,N_24906);
or U25202 (N_25202,N_25158,N_25177);
nand U25203 (N_25203,N_25168,N_25037);
nand U25204 (N_25204,N_24903,N_24953);
or U25205 (N_25205,N_25007,N_25090);
nor U25206 (N_25206,N_24927,N_25070);
nand U25207 (N_25207,N_25123,N_24980);
or U25208 (N_25208,N_24968,N_25197);
nor U25209 (N_25209,N_25086,N_24902);
and U25210 (N_25210,N_25011,N_25003);
nor U25211 (N_25211,N_25085,N_24954);
nor U25212 (N_25212,N_25028,N_24928);
nand U25213 (N_25213,N_25182,N_24922);
nor U25214 (N_25214,N_25116,N_24999);
xnor U25215 (N_25215,N_25072,N_25171);
nor U25216 (N_25216,N_25034,N_25196);
or U25217 (N_25217,N_24981,N_25138);
and U25218 (N_25218,N_25187,N_24915);
nand U25219 (N_25219,N_24951,N_25092);
xor U25220 (N_25220,N_25036,N_25170);
and U25221 (N_25221,N_25080,N_25060);
or U25222 (N_25222,N_25193,N_25115);
nand U25223 (N_25223,N_25008,N_25127);
xor U25224 (N_25224,N_25169,N_25073);
nor U25225 (N_25225,N_25048,N_25061);
nand U25226 (N_25226,N_25179,N_25054);
and U25227 (N_25227,N_25091,N_24992);
and U25228 (N_25228,N_24930,N_25063);
and U25229 (N_25229,N_25083,N_25192);
and U25230 (N_25230,N_25121,N_25096);
or U25231 (N_25231,N_24923,N_25174);
nor U25232 (N_25232,N_24971,N_25032);
nor U25233 (N_25233,N_24982,N_24996);
or U25234 (N_25234,N_25033,N_25058);
xor U25235 (N_25235,N_24918,N_25173);
and U25236 (N_25236,N_24944,N_24946);
nor U25237 (N_25237,N_24914,N_25125);
nand U25238 (N_25238,N_25052,N_24958);
or U25239 (N_25239,N_25064,N_24900);
xor U25240 (N_25240,N_25142,N_25134);
or U25241 (N_25241,N_24936,N_25057);
and U25242 (N_25242,N_25135,N_24939);
xor U25243 (N_25243,N_24907,N_24934);
xor U25244 (N_25244,N_24962,N_24937);
or U25245 (N_25245,N_25044,N_24935);
and U25246 (N_25246,N_25189,N_25159);
nor U25247 (N_25247,N_25199,N_25014);
nand U25248 (N_25248,N_25103,N_24976);
and U25249 (N_25249,N_24908,N_24977);
and U25250 (N_25250,N_25129,N_25066);
nand U25251 (N_25251,N_25065,N_25078);
xor U25252 (N_25252,N_25013,N_24941);
or U25253 (N_25253,N_24912,N_25143);
xnor U25254 (N_25254,N_25109,N_25190);
nand U25255 (N_25255,N_25153,N_25157);
nor U25256 (N_25256,N_25162,N_25149);
or U25257 (N_25257,N_24955,N_25039);
and U25258 (N_25258,N_25104,N_24917);
or U25259 (N_25259,N_25046,N_24959);
nand U25260 (N_25260,N_24921,N_24929);
and U25261 (N_25261,N_25185,N_25110);
xnor U25262 (N_25262,N_24964,N_24905);
and U25263 (N_25263,N_24949,N_25015);
nand U25264 (N_25264,N_25082,N_25035);
nor U25265 (N_25265,N_25006,N_25016);
nor U25266 (N_25266,N_25042,N_25178);
nand U25267 (N_25267,N_25088,N_25126);
xor U25268 (N_25268,N_25040,N_25183);
nand U25269 (N_25269,N_25020,N_24950);
nand U25270 (N_25270,N_25136,N_24988);
nor U25271 (N_25271,N_24938,N_24926);
nand U25272 (N_25272,N_24952,N_25074);
nand U25273 (N_25273,N_25155,N_25120);
nor U25274 (N_25274,N_24970,N_25075);
nand U25275 (N_25275,N_25027,N_24972);
nand U25276 (N_25276,N_25195,N_24910);
and U25277 (N_25277,N_25053,N_25194);
nand U25278 (N_25278,N_25002,N_25191);
nor U25279 (N_25279,N_24979,N_25026);
and U25280 (N_25280,N_25150,N_25087);
and U25281 (N_25281,N_24932,N_25102);
and U25282 (N_25282,N_24986,N_24933);
nand U25283 (N_25283,N_25146,N_25068);
nor U25284 (N_25284,N_25176,N_24963);
xor U25285 (N_25285,N_25012,N_25009);
or U25286 (N_25286,N_24931,N_24960);
xor U25287 (N_25287,N_25100,N_25081);
or U25288 (N_25288,N_25180,N_25163);
xor U25289 (N_25289,N_25119,N_25045);
nor U25290 (N_25290,N_24983,N_24956);
nand U25291 (N_25291,N_25132,N_25079);
and U25292 (N_25292,N_25019,N_25167);
nor U25293 (N_25293,N_25041,N_25114);
and U25294 (N_25294,N_25144,N_25118);
nor U25295 (N_25295,N_25017,N_25106);
or U25296 (N_25296,N_24966,N_25067);
nor U25297 (N_25297,N_25055,N_25165);
nor U25298 (N_25298,N_25122,N_25181);
and U25299 (N_25299,N_25128,N_25147);
nand U25300 (N_25300,N_24920,N_24967);
xor U25301 (N_25301,N_24985,N_25095);
nor U25302 (N_25302,N_25071,N_25145);
and U25303 (N_25303,N_25076,N_24916);
xnor U25304 (N_25304,N_24924,N_24948);
and U25305 (N_25305,N_24973,N_25161);
xor U25306 (N_25306,N_25022,N_25077);
xor U25307 (N_25307,N_25164,N_25031);
or U25308 (N_25308,N_24993,N_24997);
nand U25309 (N_25309,N_25188,N_25137);
xor U25310 (N_25310,N_25154,N_24961);
nand U25311 (N_25311,N_25050,N_25160);
xnor U25312 (N_25312,N_25024,N_25148);
or U25313 (N_25313,N_24909,N_25141);
nor U25314 (N_25314,N_25133,N_25139);
nor U25315 (N_25315,N_25117,N_25084);
and U25316 (N_25316,N_25098,N_25059);
nand U25317 (N_25317,N_25062,N_25111);
and U25318 (N_25318,N_25140,N_24911);
xor U25319 (N_25319,N_25000,N_24901);
nor U25320 (N_25320,N_25186,N_25152);
xor U25321 (N_25321,N_24942,N_24998);
nor U25322 (N_25322,N_25001,N_25038);
and U25323 (N_25323,N_25131,N_25166);
and U25324 (N_25324,N_24974,N_25101);
nor U25325 (N_25325,N_24943,N_25029);
or U25326 (N_25326,N_24947,N_25093);
xnor U25327 (N_25327,N_25156,N_24989);
nor U25328 (N_25328,N_25043,N_24984);
or U25329 (N_25329,N_25018,N_24987);
nand U25330 (N_25330,N_25004,N_25025);
or U25331 (N_25331,N_25056,N_24919);
and U25332 (N_25332,N_24975,N_24957);
nand U25333 (N_25333,N_24965,N_24913);
xnor U25334 (N_25334,N_25021,N_25105);
nor U25335 (N_25335,N_24978,N_25069);
nand U25336 (N_25336,N_25097,N_24969);
nand U25337 (N_25337,N_25094,N_25010);
and U25338 (N_25338,N_24991,N_24904);
xnor U25339 (N_25339,N_24990,N_25099);
nor U25340 (N_25340,N_24925,N_25124);
or U25341 (N_25341,N_25112,N_25047);
nor U25342 (N_25342,N_25113,N_25151);
or U25343 (N_25343,N_24995,N_25184);
xnor U25344 (N_25344,N_25051,N_25172);
nand U25345 (N_25345,N_25107,N_25030);
xnor U25346 (N_25346,N_25005,N_25175);
or U25347 (N_25347,N_24940,N_25198);
or U25348 (N_25348,N_25089,N_24945);
nand U25349 (N_25349,N_24994,N_25023);
and U25350 (N_25350,N_24988,N_25195);
nor U25351 (N_25351,N_25075,N_24906);
or U25352 (N_25352,N_25140,N_25151);
xor U25353 (N_25353,N_25031,N_24980);
or U25354 (N_25354,N_25076,N_24903);
nor U25355 (N_25355,N_24931,N_25033);
nor U25356 (N_25356,N_24940,N_25136);
xor U25357 (N_25357,N_25109,N_25107);
nor U25358 (N_25358,N_25026,N_25175);
nand U25359 (N_25359,N_25075,N_24904);
xnor U25360 (N_25360,N_25165,N_25143);
nand U25361 (N_25361,N_24919,N_25125);
nand U25362 (N_25362,N_25102,N_24959);
nand U25363 (N_25363,N_25017,N_25123);
nand U25364 (N_25364,N_24988,N_25116);
xor U25365 (N_25365,N_25088,N_25018);
nand U25366 (N_25366,N_24966,N_25100);
and U25367 (N_25367,N_25060,N_25122);
nand U25368 (N_25368,N_25176,N_25188);
or U25369 (N_25369,N_25113,N_25078);
or U25370 (N_25370,N_24924,N_24987);
xnor U25371 (N_25371,N_25014,N_24965);
xor U25372 (N_25372,N_25070,N_25082);
or U25373 (N_25373,N_25078,N_25134);
nand U25374 (N_25374,N_25149,N_25107);
nor U25375 (N_25375,N_24988,N_24907);
xnor U25376 (N_25376,N_25015,N_25053);
xnor U25377 (N_25377,N_24932,N_24926);
nor U25378 (N_25378,N_25106,N_24924);
and U25379 (N_25379,N_25054,N_25011);
nor U25380 (N_25380,N_25071,N_25117);
or U25381 (N_25381,N_25129,N_25075);
xnor U25382 (N_25382,N_25094,N_25135);
nand U25383 (N_25383,N_24917,N_24949);
xor U25384 (N_25384,N_24987,N_25055);
and U25385 (N_25385,N_25139,N_25081);
nor U25386 (N_25386,N_25058,N_25119);
nand U25387 (N_25387,N_24982,N_25021);
or U25388 (N_25388,N_25079,N_25116);
or U25389 (N_25389,N_25110,N_25121);
and U25390 (N_25390,N_25097,N_25096);
or U25391 (N_25391,N_24965,N_25090);
xnor U25392 (N_25392,N_24965,N_24971);
nor U25393 (N_25393,N_25145,N_24951);
nor U25394 (N_25394,N_25092,N_25026);
nor U25395 (N_25395,N_24998,N_25196);
nor U25396 (N_25396,N_25166,N_25179);
and U25397 (N_25397,N_25096,N_24943);
xor U25398 (N_25398,N_25183,N_25012);
and U25399 (N_25399,N_24950,N_25137);
nand U25400 (N_25400,N_25103,N_25101);
nor U25401 (N_25401,N_24925,N_25040);
nand U25402 (N_25402,N_24913,N_25039);
or U25403 (N_25403,N_24974,N_24922);
xor U25404 (N_25404,N_25089,N_25077);
xor U25405 (N_25405,N_25089,N_25058);
xor U25406 (N_25406,N_24901,N_24968);
or U25407 (N_25407,N_25185,N_25089);
nand U25408 (N_25408,N_25179,N_25119);
nor U25409 (N_25409,N_24931,N_24990);
xor U25410 (N_25410,N_24929,N_25119);
nor U25411 (N_25411,N_24936,N_24994);
xnor U25412 (N_25412,N_25121,N_25046);
and U25413 (N_25413,N_25157,N_25014);
nand U25414 (N_25414,N_25021,N_25110);
or U25415 (N_25415,N_24977,N_25045);
and U25416 (N_25416,N_25040,N_25056);
nand U25417 (N_25417,N_24901,N_24954);
or U25418 (N_25418,N_24923,N_24956);
xnor U25419 (N_25419,N_25178,N_25193);
or U25420 (N_25420,N_25176,N_25093);
or U25421 (N_25421,N_24942,N_24908);
nor U25422 (N_25422,N_25098,N_24911);
or U25423 (N_25423,N_25007,N_25165);
xnor U25424 (N_25424,N_24933,N_24972);
xnor U25425 (N_25425,N_25128,N_25071);
or U25426 (N_25426,N_25082,N_25159);
or U25427 (N_25427,N_24914,N_25139);
and U25428 (N_25428,N_25103,N_24972);
nand U25429 (N_25429,N_25139,N_25105);
and U25430 (N_25430,N_25167,N_25182);
or U25431 (N_25431,N_25011,N_24911);
and U25432 (N_25432,N_25018,N_24985);
and U25433 (N_25433,N_24959,N_25038);
nand U25434 (N_25434,N_25168,N_25005);
nor U25435 (N_25435,N_25176,N_24903);
nor U25436 (N_25436,N_25030,N_25144);
nand U25437 (N_25437,N_25097,N_25022);
nor U25438 (N_25438,N_25061,N_24902);
nand U25439 (N_25439,N_25102,N_24921);
or U25440 (N_25440,N_24988,N_25065);
or U25441 (N_25441,N_25166,N_25153);
nor U25442 (N_25442,N_24948,N_25006);
and U25443 (N_25443,N_25175,N_25090);
xor U25444 (N_25444,N_24935,N_25053);
nor U25445 (N_25445,N_25110,N_24998);
nand U25446 (N_25446,N_24991,N_25146);
nand U25447 (N_25447,N_24968,N_25116);
xor U25448 (N_25448,N_24925,N_25016);
nand U25449 (N_25449,N_24925,N_25162);
nor U25450 (N_25450,N_25055,N_25056);
or U25451 (N_25451,N_25191,N_25058);
and U25452 (N_25452,N_25151,N_25036);
xnor U25453 (N_25453,N_25014,N_25028);
xnor U25454 (N_25454,N_25052,N_24900);
nor U25455 (N_25455,N_25024,N_25054);
xor U25456 (N_25456,N_24965,N_25156);
or U25457 (N_25457,N_25171,N_24953);
xnor U25458 (N_25458,N_25121,N_25068);
xnor U25459 (N_25459,N_24997,N_24948);
and U25460 (N_25460,N_24948,N_25183);
nand U25461 (N_25461,N_25166,N_25097);
nor U25462 (N_25462,N_25116,N_25175);
and U25463 (N_25463,N_25014,N_25127);
xnor U25464 (N_25464,N_25071,N_24957);
nand U25465 (N_25465,N_25160,N_24916);
xor U25466 (N_25466,N_25017,N_25177);
or U25467 (N_25467,N_25084,N_25056);
or U25468 (N_25468,N_25179,N_24986);
nor U25469 (N_25469,N_25137,N_24918);
or U25470 (N_25470,N_24907,N_24928);
nor U25471 (N_25471,N_25004,N_25041);
nand U25472 (N_25472,N_25189,N_24942);
and U25473 (N_25473,N_25045,N_25072);
and U25474 (N_25474,N_25143,N_25115);
xor U25475 (N_25475,N_25060,N_25018);
nor U25476 (N_25476,N_25191,N_25183);
or U25477 (N_25477,N_25157,N_25103);
and U25478 (N_25478,N_25057,N_25019);
nor U25479 (N_25479,N_25106,N_25059);
and U25480 (N_25480,N_25106,N_25131);
and U25481 (N_25481,N_25133,N_24983);
or U25482 (N_25482,N_25030,N_25053);
and U25483 (N_25483,N_24905,N_24902);
xnor U25484 (N_25484,N_25082,N_25067);
nand U25485 (N_25485,N_24907,N_25190);
nor U25486 (N_25486,N_25137,N_24928);
and U25487 (N_25487,N_25029,N_24963);
nand U25488 (N_25488,N_25110,N_25048);
or U25489 (N_25489,N_25112,N_25101);
or U25490 (N_25490,N_25108,N_25035);
nor U25491 (N_25491,N_24999,N_25036);
xnor U25492 (N_25492,N_25079,N_25064);
nand U25493 (N_25493,N_25177,N_25170);
or U25494 (N_25494,N_25027,N_25058);
and U25495 (N_25495,N_25149,N_25043);
nand U25496 (N_25496,N_25009,N_25084);
nand U25497 (N_25497,N_24969,N_25036);
and U25498 (N_25498,N_25172,N_25160);
or U25499 (N_25499,N_24989,N_25110);
nor U25500 (N_25500,N_25203,N_25348);
nand U25501 (N_25501,N_25351,N_25398);
and U25502 (N_25502,N_25336,N_25202);
and U25503 (N_25503,N_25280,N_25232);
nor U25504 (N_25504,N_25380,N_25426);
nand U25505 (N_25505,N_25282,N_25272);
or U25506 (N_25506,N_25328,N_25381);
xor U25507 (N_25507,N_25448,N_25352);
nand U25508 (N_25508,N_25230,N_25439);
nor U25509 (N_25509,N_25362,N_25333);
nand U25510 (N_25510,N_25223,N_25413);
nor U25511 (N_25511,N_25214,N_25461);
and U25512 (N_25512,N_25329,N_25371);
nor U25513 (N_25513,N_25251,N_25377);
xnor U25514 (N_25514,N_25240,N_25309);
nor U25515 (N_25515,N_25313,N_25338);
xnor U25516 (N_25516,N_25421,N_25497);
and U25517 (N_25517,N_25295,N_25496);
or U25518 (N_25518,N_25482,N_25479);
nand U25519 (N_25519,N_25318,N_25498);
nand U25520 (N_25520,N_25345,N_25226);
and U25521 (N_25521,N_25473,N_25443);
xor U25522 (N_25522,N_25215,N_25363);
nor U25523 (N_25523,N_25359,N_25216);
xor U25524 (N_25524,N_25291,N_25499);
and U25525 (N_25525,N_25211,N_25387);
nor U25526 (N_25526,N_25383,N_25449);
nand U25527 (N_25527,N_25365,N_25423);
and U25528 (N_25528,N_25407,N_25281);
and U25529 (N_25529,N_25428,N_25430);
nor U25530 (N_25530,N_25323,N_25257);
and U25531 (N_25531,N_25289,N_25389);
nor U25532 (N_25532,N_25297,N_25401);
nor U25533 (N_25533,N_25206,N_25431);
nand U25534 (N_25534,N_25285,N_25258);
nand U25535 (N_25535,N_25422,N_25264);
and U25536 (N_25536,N_25486,N_25343);
xnor U25537 (N_25537,N_25469,N_25265);
xnor U25538 (N_25538,N_25330,N_25459);
nor U25539 (N_25539,N_25332,N_25484);
and U25540 (N_25540,N_25491,N_25435);
nand U25541 (N_25541,N_25236,N_25267);
xnor U25542 (N_25542,N_25445,N_25494);
xnor U25543 (N_25543,N_25229,N_25488);
and U25544 (N_25544,N_25235,N_25405);
nor U25545 (N_25545,N_25299,N_25460);
or U25546 (N_25546,N_25386,N_25485);
xor U25547 (N_25547,N_25324,N_25385);
and U25548 (N_25548,N_25477,N_25286);
nor U25549 (N_25549,N_25391,N_25288);
or U25550 (N_25550,N_25438,N_25481);
or U25551 (N_25551,N_25255,N_25261);
nor U25552 (N_25552,N_25246,N_25266);
nor U25553 (N_25553,N_25478,N_25274);
xnor U25554 (N_25554,N_25409,N_25315);
xnor U25555 (N_25555,N_25369,N_25326);
xor U25556 (N_25556,N_25487,N_25370);
nor U25557 (N_25557,N_25356,N_25447);
nand U25558 (N_25558,N_25321,N_25366);
or U25559 (N_25559,N_25213,N_25204);
nand U25560 (N_25560,N_25278,N_25340);
or U25561 (N_25561,N_25271,N_25283);
and U25562 (N_25562,N_25450,N_25209);
xnor U25563 (N_25563,N_25222,N_25399);
nand U25564 (N_25564,N_25303,N_25200);
nor U25565 (N_25565,N_25411,N_25293);
and U25566 (N_25566,N_25316,N_25375);
or U25567 (N_25567,N_25312,N_25397);
xnor U25568 (N_25568,N_25228,N_25260);
nand U25569 (N_25569,N_25331,N_25437);
or U25570 (N_25570,N_25440,N_25433);
or U25571 (N_25571,N_25360,N_25350);
or U25572 (N_25572,N_25396,N_25256);
and U25573 (N_25573,N_25254,N_25242);
nor U25574 (N_25574,N_25467,N_25452);
nand U25575 (N_25575,N_25400,N_25493);
and U25576 (N_25576,N_25243,N_25495);
and U25577 (N_25577,N_25406,N_25208);
or U25578 (N_25578,N_25201,N_25234);
and U25579 (N_25579,N_25304,N_25263);
xnor U25580 (N_25580,N_25458,N_25474);
nand U25581 (N_25581,N_25403,N_25390);
and U25582 (N_25582,N_25319,N_25361);
nor U25583 (N_25583,N_25444,N_25489);
xnor U25584 (N_25584,N_25250,N_25429);
and U25585 (N_25585,N_25492,N_25298);
xnor U25586 (N_25586,N_25219,N_25424);
and U25587 (N_25587,N_25314,N_25410);
nand U25588 (N_25588,N_25466,N_25418);
or U25589 (N_25589,N_25320,N_25453);
nand U25590 (N_25590,N_25262,N_25376);
xnor U25591 (N_25591,N_25294,N_25412);
xnor U25592 (N_25592,N_25302,N_25357);
xor U25593 (N_25593,N_25308,N_25279);
and U25594 (N_25594,N_25358,N_25344);
nand U25595 (N_25595,N_25305,N_25420);
xnor U25596 (N_25596,N_25212,N_25220);
xor U25597 (N_25597,N_25379,N_25434);
nand U25598 (N_25598,N_25227,N_25205);
nor U25599 (N_25599,N_25373,N_25284);
or U25600 (N_25600,N_25432,N_25207);
nand U25601 (N_25601,N_25354,N_25404);
xnor U25602 (N_25602,N_25290,N_25245);
or U25603 (N_25603,N_25311,N_25382);
or U25604 (N_25604,N_25277,N_25342);
nor U25605 (N_25605,N_25327,N_25335);
nor U25606 (N_25606,N_25337,N_25468);
and U25607 (N_25607,N_25269,N_25462);
and U25608 (N_25608,N_25210,N_25237);
xnor U25609 (N_25609,N_25241,N_25441);
and U25610 (N_25610,N_25276,N_25300);
nor U25611 (N_25611,N_25217,N_25252);
xor U25612 (N_25612,N_25483,N_25393);
xor U25613 (N_25613,N_25417,N_25317);
nand U25614 (N_25614,N_25347,N_25472);
and U25615 (N_25615,N_25292,N_25425);
nor U25616 (N_25616,N_25378,N_25427);
nand U25617 (N_25617,N_25414,N_25310);
and U25618 (N_25618,N_25322,N_25451);
nand U25619 (N_25619,N_25353,N_25480);
and U25620 (N_25620,N_25239,N_25454);
and U25621 (N_25621,N_25233,N_25334);
and U25622 (N_25622,N_25490,N_25287);
nor U25623 (N_25623,N_25268,N_25275);
nor U25624 (N_25624,N_25476,N_25465);
nand U25625 (N_25625,N_25436,N_25442);
nand U25626 (N_25626,N_25419,N_25464);
and U25627 (N_25627,N_25416,N_25307);
nor U25628 (N_25628,N_25392,N_25270);
nand U25629 (N_25629,N_25247,N_25388);
or U25630 (N_25630,N_25225,N_25224);
and U25631 (N_25631,N_25394,N_25415);
or U25632 (N_25632,N_25306,N_25249);
and U25633 (N_25633,N_25457,N_25374);
and U25634 (N_25634,N_25402,N_25339);
or U25635 (N_25635,N_25341,N_25367);
nand U25636 (N_25636,N_25368,N_25221);
nand U25637 (N_25637,N_25273,N_25248);
nor U25638 (N_25638,N_25395,N_25475);
and U25639 (N_25639,N_25238,N_25218);
or U25640 (N_25640,N_25471,N_25372);
nor U25641 (N_25641,N_25325,N_25470);
nand U25642 (N_25642,N_25446,N_25346);
nand U25643 (N_25643,N_25231,N_25355);
or U25644 (N_25644,N_25301,N_25259);
or U25645 (N_25645,N_25244,N_25349);
xor U25646 (N_25646,N_25463,N_25296);
xor U25647 (N_25647,N_25364,N_25253);
nor U25648 (N_25648,N_25408,N_25455);
and U25649 (N_25649,N_25384,N_25456);
and U25650 (N_25650,N_25357,N_25225);
or U25651 (N_25651,N_25459,N_25268);
or U25652 (N_25652,N_25471,N_25473);
xor U25653 (N_25653,N_25437,N_25356);
nand U25654 (N_25654,N_25339,N_25414);
or U25655 (N_25655,N_25499,N_25219);
xor U25656 (N_25656,N_25261,N_25362);
nand U25657 (N_25657,N_25223,N_25264);
and U25658 (N_25658,N_25458,N_25227);
nor U25659 (N_25659,N_25276,N_25481);
xor U25660 (N_25660,N_25304,N_25211);
and U25661 (N_25661,N_25499,N_25424);
and U25662 (N_25662,N_25444,N_25338);
and U25663 (N_25663,N_25303,N_25207);
nor U25664 (N_25664,N_25461,N_25397);
xnor U25665 (N_25665,N_25483,N_25319);
or U25666 (N_25666,N_25369,N_25445);
nor U25667 (N_25667,N_25314,N_25252);
nand U25668 (N_25668,N_25453,N_25234);
nand U25669 (N_25669,N_25302,N_25339);
and U25670 (N_25670,N_25471,N_25303);
or U25671 (N_25671,N_25222,N_25329);
xor U25672 (N_25672,N_25429,N_25492);
xor U25673 (N_25673,N_25445,N_25412);
nand U25674 (N_25674,N_25300,N_25208);
and U25675 (N_25675,N_25439,N_25329);
nor U25676 (N_25676,N_25286,N_25423);
xor U25677 (N_25677,N_25233,N_25228);
or U25678 (N_25678,N_25225,N_25202);
xor U25679 (N_25679,N_25349,N_25396);
nor U25680 (N_25680,N_25345,N_25395);
nor U25681 (N_25681,N_25225,N_25336);
and U25682 (N_25682,N_25429,N_25311);
nor U25683 (N_25683,N_25201,N_25311);
and U25684 (N_25684,N_25348,N_25202);
and U25685 (N_25685,N_25457,N_25288);
xor U25686 (N_25686,N_25469,N_25316);
nand U25687 (N_25687,N_25224,N_25264);
xor U25688 (N_25688,N_25406,N_25489);
nor U25689 (N_25689,N_25467,N_25495);
or U25690 (N_25690,N_25346,N_25281);
and U25691 (N_25691,N_25416,N_25425);
nor U25692 (N_25692,N_25263,N_25295);
or U25693 (N_25693,N_25396,N_25323);
nor U25694 (N_25694,N_25423,N_25340);
nand U25695 (N_25695,N_25427,N_25316);
or U25696 (N_25696,N_25413,N_25433);
and U25697 (N_25697,N_25357,N_25340);
xor U25698 (N_25698,N_25273,N_25202);
and U25699 (N_25699,N_25321,N_25447);
or U25700 (N_25700,N_25269,N_25428);
nor U25701 (N_25701,N_25205,N_25414);
and U25702 (N_25702,N_25265,N_25253);
nand U25703 (N_25703,N_25446,N_25456);
nor U25704 (N_25704,N_25294,N_25267);
or U25705 (N_25705,N_25253,N_25209);
nand U25706 (N_25706,N_25405,N_25296);
nand U25707 (N_25707,N_25249,N_25449);
nor U25708 (N_25708,N_25209,N_25303);
and U25709 (N_25709,N_25385,N_25410);
or U25710 (N_25710,N_25450,N_25206);
and U25711 (N_25711,N_25382,N_25307);
nand U25712 (N_25712,N_25477,N_25350);
and U25713 (N_25713,N_25480,N_25359);
and U25714 (N_25714,N_25243,N_25275);
nand U25715 (N_25715,N_25487,N_25322);
xor U25716 (N_25716,N_25461,N_25236);
and U25717 (N_25717,N_25204,N_25469);
nor U25718 (N_25718,N_25434,N_25211);
and U25719 (N_25719,N_25481,N_25434);
or U25720 (N_25720,N_25420,N_25362);
or U25721 (N_25721,N_25308,N_25416);
nor U25722 (N_25722,N_25431,N_25303);
or U25723 (N_25723,N_25455,N_25401);
nor U25724 (N_25724,N_25277,N_25374);
nor U25725 (N_25725,N_25432,N_25405);
nand U25726 (N_25726,N_25402,N_25332);
nor U25727 (N_25727,N_25248,N_25494);
nand U25728 (N_25728,N_25428,N_25327);
nor U25729 (N_25729,N_25279,N_25304);
or U25730 (N_25730,N_25275,N_25224);
nor U25731 (N_25731,N_25392,N_25433);
or U25732 (N_25732,N_25476,N_25383);
or U25733 (N_25733,N_25398,N_25206);
nor U25734 (N_25734,N_25230,N_25357);
or U25735 (N_25735,N_25267,N_25347);
xor U25736 (N_25736,N_25366,N_25318);
nand U25737 (N_25737,N_25298,N_25479);
nor U25738 (N_25738,N_25474,N_25347);
nor U25739 (N_25739,N_25244,N_25464);
xor U25740 (N_25740,N_25453,N_25427);
nor U25741 (N_25741,N_25447,N_25410);
nand U25742 (N_25742,N_25421,N_25444);
and U25743 (N_25743,N_25241,N_25408);
or U25744 (N_25744,N_25449,N_25338);
xor U25745 (N_25745,N_25225,N_25497);
nand U25746 (N_25746,N_25232,N_25373);
and U25747 (N_25747,N_25238,N_25350);
xnor U25748 (N_25748,N_25208,N_25346);
or U25749 (N_25749,N_25211,N_25309);
xor U25750 (N_25750,N_25374,N_25306);
xor U25751 (N_25751,N_25292,N_25251);
xnor U25752 (N_25752,N_25446,N_25384);
xor U25753 (N_25753,N_25220,N_25378);
nor U25754 (N_25754,N_25257,N_25200);
or U25755 (N_25755,N_25263,N_25326);
xnor U25756 (N_25756,N_25477,N_25311);
or U25757 (N_25757,N_25353,N_25287);
nor U25758 (N_25758,N_25420,N_25471);
or U25759 (N_25759,N_25236,N_25332);
xor U25760 (N_25760,N_25287,N_25224);
nor U25761 (N_25761,N_25210,N_25225);
nor U25762 (N_25762,N_25329,N_25470);
nand U25763 (N_25763,N_25227,N_25287);
or U25764 (N_25764,N_25470,N_25416);
nand U25765 (N_25765,N_25206,N_25478);
and U25766 (N_25766,N_25255,N_25386);
nor U25767 (N_25767,N_25498,N_25213);
nand U25768 (N_25768,N_25487,N_25461);
nand U25769 (N_25769,N_25201,N_25382);
nor U25770 (N_25770,N_25295,N_25340);
and U25771 (N_25771,N_25294,N_25208);
and U25772 (N_25772,N_25424,N_25496);
nand U25773 (N_25773,N_25307,N_25200);
or U25774 (N_25774,N_25259,N_25321);
nor U25775 (N_25775,N_25458,N_25303);
nand U25776 (N_25776,N_25481,N_25351);
or U25777 (N_25777,N_25461,N_25395);
xor U25778 (N_25778,N_25416,N_25402);
and U25779 (N_25779,N_25424,N_25256);
or U25780 (N_25780,N_25478,N_25329);
and U25781 (N_25781,N_25313,N_25236);
xor U25782 (N_25782,N_25237,N_25247);
or U25783 (N_25783,N_25249,N_25465);
or U25784 (N_25784,N_25292,N_25236);
and U25785 (N_25785,N_25393,N_25427);
nor U25786 (N_25786,N_25240,N_25304);
xor U25787 (N_25787,N_25485,N_25360);
and U25788 (N_25788,N_25428,N_25367);
xor U25789 (N_25789,N_25368,N_25336);
and U25790 (N_25790,N_25452,N_25299);
or U25791 (N_25791,N_25273,N_25348);
nor U25792 (N_25792,N_25227,N_25217);
nor U25793 (N_25793,N_25344,N_25390);
nor U25794 (N_25794,N_25450,N_25284);
xnor U25795 (N_25795,N_25227,N_25499);
and U25796 (N_25796,N_25280,N_25447);
or U25797 (N_25797,N_25282,N_25442);
or U25798 (N_25798,N_25389,N_25443);
nor U25799 (N_25799,N_25309,N_25297);
nand U25800 (N_25800,N_25770,N_25597);
or U25801 (N_25801,N_25548,N_25626);
and U25802 (N_25802,N_25538,N_25603);
xnor U25803 (N_25803,N_25577,N_25753);
nand U25804 (N_25804,N_25572,N_25585);
nand U25805 (N_25805,N_25765,N_25644);
nand U25806 (N_25806,N_25788,N_25576);
and U25807 (N_25807,N_25612,N_25732);
nor U25808 (N_25808,N_25710,N_25535);
or U25809 (N_25809,N_25558,N_25615);
or U25810 (N_25810,N_25718,N_25557);
or U25811 (N_25811,N_25506,N_25648);
nor U25812 (N_25812,N_25617,N_25503);
nor U25813 (N_25813,N_25532,N_25759);
and U25814 (N_25814,N_25652,N_25790);
nand U25815 (N_25815,N_25573,N_25758);
and U25816 (N_25816,N_25781,N_25594);
and U25817 (N_25817,N_25688,N_25614);
or U25818 (N_25818,N_25541,N_25709);
nor U25819 (N_25819,N_25708,N_25655);
xor U25820 (N_25820,N_25663,N_25675);
and U25821 (N_25821,N_25681,N_25504);
nor U25822 (N_25822,N_25703,N_25613);
xnor U25823 (N_25823,N_25764,N_25780);
or U25824 (N_25824,N_25665,N_25555);
nand U25825 (N_25825,N_25734,N_25658);
nor U25826 (N_25826,N_25656,N_25598);
and U25827 (N_25827,N_25638,N_25537);
and U25828 (N_25828,N_25720,N_25768);
and U25829 (N_25829,N_25608,N_25642);
or U25830 (N_25830,N_25698,N_25775);
xnor U25831 (N_25831,N_25755,N_25629);
or U25832 (N_25832,N_25702,N_25729);
or U25833 (N_25833,N_25735,N_25578);
and U25834 (N_25834,N_25673,N_25674);
xor U25835 (N_25835,N_25623,N_25667);
and U25836 (N_25836,N_25550,N_25528);
or U25837 (N_25837,N_25630,N_25697);
xnor U25838 (N_25838,N_25501,N_25502);
or U25839 (N_25839,N_25782,N_25592);
nor U25840 (N_25840,N_25736,N_25602);
nor U25841 (N_25841,N_25590,N_25717);
nor U25842 (N_25842,N_25647,N_25583);
nand U25843 (N_25843,N_25515,N_25624);
xor U25844 (N_25844,N_25591,N_25679);
or U25845 (N_25845,N_25611,N_25536);
nand U25846 (N_25846,N_25547,N_25713);
or U25847 (N_25847,N_25793,N_25518);
nand U25848 (N_25848,N_25527,N_25634);
xnor U25849 (N_25849,N_25659,N_25600);
nor U25850 (N_25850,N_25726,N_25760);
xnor U25851 (N_25851,N_25566,N_25798);
and U25852 (N_25852,N_25771,N_25563);
or U25853 (N_25853,N_25582,N_25737);
xor U25854 (N_25854,N_25721,N_25749);
nand U25855 (N_25855,N_25625,N_25797);
nand U25856 (N_25856,N_25526,N_25523);
xnor U25857 (N_25857,N_25680,N_25514);
or U25858 (N_25858,N_25744,N_25776);
and U25859 (N_25859,N_25530,N_25787);
or U25860 (N_25860,N_25773,N_25699);
or U25861 (N_25861,N_25540,N_25564);
xnor U25862 (N_25862,N_25605,N_25641);
nor U25863 (N_25863,N_25618,N_25789);
and U25864 (N_25864,N_25524,N_25549);
xnor U25865 (N_25865,N_25546,N_25619);
nand U25866 (N_25866,N_25724,N_25531);
and U25867 (N_25867,N_25731,N_25669);
nor U25868 (N_25868,N_25685,N_25589);
or U25869 (N_25869,N_25728,N_25742);
and U25870 (N_25870,N_25701,N_25645);
nand U25871 (N_25871,N_25763,N_25580);
or U25872 (N_25872,N_25571,N_25521);
and U25873 (N_25873,N_25695,N_25568);
or U25874 (N_25874,N_25604,N_25750);
and U25875 (N_25875,N_25693,N_25637);
and U25876 (N_25876,N_25607,N_25762);
xor U25877 (N_25877,N_25616,N_25743);
xor U25878 (N_25878,N_25539,N_25554);
xnor U25879 (N_25879,N_25653,N_25640);
nand U25880 (N_25880,N_25766,N_25767);
nand U25881 (N_25881,N_25761,N_25574);
nor U25882 (N_25882,N_25622,N_25551);
or U25883 (N_25883,N_25687,N_25643);
xor U25884 (N_25884,N_25715,N_25633);
nor U25885 (N_25885,N_25684,N_25786);
xnor U25886 (N_25886,N_25741,N_25799);
or U25887 (N_25887,N_25654,N_25586);
nand U25888 (N_25888,N_25544,N_25757);
and U25889 (N_25889,N_25696,N_25769);
xnor U25890 (N_25890,N_25716,N_25785);
xnor U25891 (N_25891,N_25509,N_25778);
nand U25892 (N_25892,N_25683,N_25575);
nor U25893 (N_25893,N_25632,N_25661);
nor U25894 (N_25894,N_25529,N_25746);
nand U25895 (N_25895,N_25651,N_25584);
or U25896 (N_25896,N_25784,N_25588);
nand U25897 (N_25897,N_25533,N_25631);
nor U25898 (N_25898,N_25723,N_25690);
nor U25899 (N_25899,N_25794,N_25507);
or U25900 (N_25900,N_25620,N_25796);
or U25901 (N_25901,N_25738,N_25739);
and U25902 (N_25902,N_25567,N_25672);
xnor U25903 (N_25903,N_25593,N_25649);
or U25904 (N_25904,N_25595,N_25581);
or U25905 (N_25905,N_25639,N_25561);
and U25906 (N_25906,N_25610,N_25560);
nor U25907 (N_25907,N_25609,N_25512);
or U25908 (N_25908,N_25792,N_25727);
and U25909 (N_25909,N_25606,N_25748);
or U25910 (N_25910,N_25601,N_25756);
xnor U25911 (N_25911,N_25635,N_25714);
or U25912 (N_25912,N_25500,N_25516);
and U25913 (N_25913,N_25627,N_25508);
xnor U25914 (N_25914,N_25543,N_25691);
and U25915 (N_25915,N_25587,N_25562);
nand U25916 (N_25916,N_25772,N_25522);
or U25917 (N_25917,N_25678,N_25525);
xor U25918 (N_25918,N_25570,N_25777);
nor U25919 (N_25919,N_25556,N_25689);
nand U25920 (N_25920,N_25664,N_25711);
or U25921 (N_25921,N_25552,N_25725);
and U25922 (N_25922,N_25650,N_25682);
or U25923 (N_25923,N_25666,N_25704);
nor U25924 (N_25924,N_25706,N_25686);
nand U25925 (N_25925,N_25677,N_25621);
nand U25926 (N_25926,N_25660,N_25545);
or U25927 (N_25927,N_25505,N_25754);
and U25928 (N_25928,N_25692,N_25745);
xnor U25929 (N_25929,N_25795,N_25740);
and U25930 (N_25930,N_25553,N_25694);
and U25931 (N_25931,N_25599,N_25534);
nand U25932 (N_25932,N_25705,N_25559);
nand U25933 (N_25933,N_25520,N_25668);
nor U25934 (N_25934,N_25712,N_25662);
and U25935 (N_25935,N_25628,N_25700);
and U25936 (N_25936,N_25751,N_25783);
and U25937 (N_25937,N_25719,N_25519);
or U25938 (N_25938,N_25670,N_25646);
nor U25939 (N_25939,N_25752,N_25774);
xnor U25940 (N_25940,N_25722,N_25747);
and U25941 (N_25941,N_25707,N_25510);
nor U25942 (N_25942,N_25569,N_25779);
and U25943 (N_25943,N_25579,N_25671);
or U25944 (N_25944,N_25791,N_25657);
or U25945 (N_25945,N_25733,N_25636);
nand U25946 (N_25946,N_25596,N_25517);
xnor U25947 (N_25947,N_25676,N_25730);
or U25948 (N_25948,N_25565,N_25542);
nor U25949 (N_25949,N_25513,N_25511);
nand U25950 (N_25950,N_25728,N_25739);
or U25951 (N_25951,N_25780,N_25537);
or U25952 (N_25952,N_25774,N_25632);
or U25953 (N_25953,N_25601,N_25567);
or U25954 (N_25954,N_25756,N_25702);
and U25955 (N_25955,N_25606,N_25576);
or U25956 (N_25956,N_25568,N_25785);
and U25957 (N_25957,N_25750,N_25587);
and U25958 (N_25958,N_25675,N_25531);
or U25959 (N_25959,N_25600,N_25769);
and U25960 (N_25960,N_25501,N_25759);
nor U25961 (N_25961,N_25663,N_25733);
or U25962 (N_25962,N_25736,N_25544);
nor U25963 (N_25963,N_25780,N_25674);
xor U25964 (N_25964,N_25765,N_25721);
and U25965 (N_25965,N_25693,N_25753);
nand U25966 (N_25966,N_25535,N_25703);
and U25967 (N_25967,N_25742,N_25690);
xnor U25968 (N_25968,N_25712,N_25774);
xor U25969 (N_25969,N_25506,N_25520);
xnor U25970 (N_25970,N_25594,N_25538);
and U25971 (N_25971,N_25762,N_25505);
nand U25972 (N_25972,N_25758,N_25508);
nor U25973 (N_25973,N_25655,N_25665);
nand U25974 (N_25974,N_25521,N_25694);
and U25975 (N_25975,N_25545,N_25694);
nand U25976 (N_25976,N_25697,N_25512);
nor U25977 (N_25977,N_25707,N_25690);
nand U25978 (N_25978,N_25753,N_25727);
nor U25979 (N_25979,N_25565,N_25612);
nand U25980 (N_25980,N_25799,N_25569);
and U25981 (N_25981,N_25585,N_25655);
and U25982 (N_25982,N_25745,N_25646);
or U25983 (N_25983,N_25548,N_25604);
nor U25984 (N_25984,N_25618,N_25759);
nand U25985 (N_25985,N_25599,N_25793);
nand U25986 (N_25986,N_25597,N_25532);
nand U25987 (N_25987,N_25502,N_25710);
xnor U25988 (N_25988,N_25722,N_25761);
xnor U25989 (N_25989,N_25653,N_25750);
and U25990 (N_25990,N_25604,N_25675);
xnor U25991 (N_25991,N_25785,N_25672);
nand U25992 (N_25992,N_25517,N_25541);
xor U25993 (N_25993,N_25775,N_25772);
nand U25994 (N_25994,N_25571,N_25755);
nand U25995 (N_25995,N_25655,N_25576);
and U25996 (N_25996,N_25531,N_25685);
and U25997 (N_25997,N_25669,N_25555);
or U25998 (N_25998,N_25570,N_25524);
nor U25999 (N_25999,N_25576,N_25507);
and U26000 (N_26000,N_25608,N_25772);
and U26001 (N_26001,N_25662,N_25586);
nor U26002 (N_26002,N_25695,N_25592);
or U26003 (N_26003,N_25547,N_25593);
nor U26004 (N_26004,N_25716,N_25723);
nor U26005 (N_26005,N_25723,N_25522);
xnor U26006 (N_26006,N_25579,N_25766);
nand U26007 (N_26007,N_25785,N_25505);
or U26008 (N_26008,N_25525,N_25704);
or U26009 (N_26009,N_25567,N_25667);
xor U26010 (N_26010,N_25608,N_25525);
or U26011 (N_26011,N_25552,N_25698);
xnor U26012 (N_26012,N_25704,N_25721);
nor U26013 (N_26013,N_25508,N_25596);
and U26014 (N_26014,N_25662,N_25762);
and U26015 (N_26015,N_25540,N_25503);
and U26016 (N_26016,N_25798,N_25570);
and U26017 (N_26017,N_25719,N_25767);
nand U26018 (N_26018,N_25670,N_25664);
nor U26019 (N_26019,N_25537,N_25593);
or U26020 (N_26020,N_25637,N_25607);
nand U26021 (N_26021,N_25655,N_25700);
and U26022 (N_26022,N_25528,N_25592);
or U26023 (N_26023,N_25606,N_25658);
nor U26024 (N_26024,N_25763,N_25782);
or U26025 (N_26025,N_25676,N_25639);
or U26026 (N_26026,N_25738,N_25564);
xor U26027 (N_26027,N_25617,N_25551);
nand U26028 (N_26028,N_25625,N_25771);
nand U26029 (N_26029,N_25749,N_25543);
nand U26030 (N_26030,N_25639,N_25547);
and U26031 (N_26031,N_25641,N_25612);
and U26032 (N_26032,N_25542,N_25695);
and U26033 (N_26033,N_25762,N_25559);
nand U26034 (N_26034,N_25590,N_25767);
or U26035 (N_26035,N_25748,N_25656);
and U26036 (N_26036,N_25535,N_25619);
nor U26037 (N_26037,N_25791,N_25626);
nor U26038 (N_26038,N_25767,N_25570);
nand U26039 (N_26039,N_25533,N_25754);
and U26040 (N_26040,N_25618,N_25588);
and U26041 (N_26041,N_25704,N_25512);
or U26042 (N_26042,N_25595,N_25542);
and U26043 (N_26043,N_25534,N_25792);
nand U26044 (N_26044,N_25705,N_25697);
or U26045 (N_26045,N_25764,N_25613);
and U26046 (N_26046,N_25776,N_25520);
nand U26047 (N_26047,N_25716,N_25741);
or U26048 (N_26048,N_25777,N_25684);
or U26049 (N_26049,N_25760,N_25566);
xor U26050 (N_26050,N_25546,N_25527);
and U26051 (N_26051,N_25730,N_25682);
nor U26052 (N_26052,N_25565,N_25586);
and U26053 (N_26053,N_25558,N_25598);
xor U26054 (N_26054,N_25780,N_25586);
xnor U26055 (N_26055,N_25606,N_25778);
and U26056 (N_26056,N_25616,N_25598);
or U26057 (N_26057,N_25694,N_25759);
or U26058 (N_26058,N_25667,N_25515);
nand U26059 (N_26059,N_25666,N_25618);
nand U26060 (N_26060,N_25521,N_25561);
nand U26061 (N_26061,N_25689,N_25661);
nor U26062 (N_26062,N_25613,N_25717);
xnor U26063 (N_26063,N_25534,N_25563);
and U26064 (N_26064,N_25532,N_25664);
nand U26065 (N_26065,N_25712,N_25758);
nand U26066 (N_26066,N_25799,N_25742);
nand U26067 (N_26067,N_25602,N_25684);
or U26068 (N_26068,N_25729,N_25680);
nor U26069 (N_26069,N_25664,N_25698);
nor U26070 (N_26070,N_25792,N_25783);
and U26071 (N_26071,N_25758,N_25745);
or U26072 (N_26072,N_25769,N_25786);
nand U26073 (N_26073,N_25659,N_25533);
nor U26074 (N_26074,N_25678,N_25772);
xnor U26075 (N_26075,N_25780,N_25781);
xnor U26076 (N_26076,N_25561,N_25709);
nand U26077 (N_26077,N_25549,N_25643);
or U26078 (N_26078,N_25740,N_25532);
nor U26079 (N_26079,N_25642,N_25671);
nor U26080 (N_26080,N_25689,N_25786);
and U26081 (N_26081,N_25603,N_25718);
nand U26082 (N_26082,N_25541,N_25726);
or U26083 (N_26083,N_25734,N_25559);
xor U26084 (N_26084,N_25596,N_25593);
or U26085 (N_26085,N_25783,N_25550);
xor U26086 (N_26086,N_25616,N_25560);
xnor U26087 (N_26087,N_25729,N_25634);
and U26088 (N_26088,N_25530,N_25697);
and U26089 (N_26089,N_25726,N_25616);
and U26090 (N_26090,N_25523,N_25577);
or U26091 (N_26091,N_25663,N_25794);
or U26092 (N_26092,N_25500,N_25618);
nor U26093 (N_26093,N_25611,N_25547);
nand U26094 (N_26094,N_25505,N_25578);
and U26095 (N_26095,N_25695,N_25650);
nand U26096 (N_26096,N_25648,N_25556);
or U26097 (N_26097,N_25632,N_25619);
and U26098 (N_26098,N_25693,N_25724);
nor U26099 (N_26099,N_25511,N_25723);
and U26100 (N_26100,N_25830,N_25950);
or U26101 (N_26101,N_25871,N_25937);
or U26102 (N_26102,N_25823,N_25898);
xnor U26103 (N_26103,N_26075,N_25897);
nor U26104 (N_26104,N_26097,N_25826);
nor U26105 (N_26105,N_25902,N_25940);
xor U26106 (N_26106,N_26064,N_26099);
nand U26107 (N_26107,N_25925,N_26028);
nor U26108 (N_26108,N_25883,N_26083);
and U26109 (N_26109,N_26005,N_25843);
xnor U26110 (N_26110,N_25936,N_26069);
nor U26111 (N_26111,N_26037,N_26041);
xor U26112 (N_26112,N_26022,N_26065);
xor U26113 (N_26113,N_25904,N_25921);
xnor U26114 (N_26114,N_25948,N_25913);
xnor U26115 (N_26115,N_25828,N_25879);
or U26116 (N_26116,N_25842,N_25837);
xnor U26117 (N_26117,N_25814,N_25896);
and U26118 (N_26118,N_25803,N_25806);
or U26119 (N_26119,N_25875,N_25822);
and U26120 (N_26120,N_25919,N_25846);
nand U26121 (N_26121,N_25858,N_25972);
nor U26122 (N_26122,N_25911,N_25848);
or U26123 (N_26123,N_25918,N_25833);
nand U26124 (N_26124,N_25861,N_26093);
xor U26125 (N_26125,N_26098,N_25965);
nor U26126 (N_26126,N_25800,N_25834);
and U26127 (N_26127,N_26011,N_26010);
nand U26128 (N_26128,N_25981,N_25817);
and U26129 (N_26129,N_25844,N_25939);
and U26130 (N_26130,N_26077,N_25841);
xnor U26131 (N_26131,N_26040,N_25889);
xnor U26132 (N_26132,N_26092,N_25983);
and U26133 (N_26133,N_26076,N_26034);
or U26134 (N_26134,N_25851,N_25960);
nand U26135 (N_26135,N_26004,N_25984);
xnor U26136 (N_26136,N_25990,N_25856);
nand U26137 (N_26137,N_26045,N_26017);
xor U26138 (N_26138,N_26029,N_26059);
nor U26139 (N_26139,N_25845,N_25964);
nand U26140 (N_26140,N_25912,N_25980);
nor U26141 (N_26141,N_26082,N_25931);
or U26142 (N_26142,N_26055,N_25963);
and U26143 (N_26143,N_25971,N_25829);
and U26144 (N_26144,N_25909,N_26057);
nor U26145 (N_26145,N_25863,N_26095);
and U26146 (N_26146,N_25891,N_26087);
nand U26147 (N_26147,N_26036,N_25838);
or U26148 (N_26148,N_26058,N_26033);
and U26149 (N_26149,N_25872,N_25975);
xor U26150 (N_26150,N_25914,N_25878);
nand U26151 (N_26151,N_26044,N_25951);
nand U26152 (N_26152,N_26047,N_26009);
nand U26153 (N_26153,N_25840,N_25991);
xnor U26154 (N_26154,N_25957,N_26062);
nand U26155 (N_26155,N_25922,N_25938);
nand U26156 (N_26156,N_26084,N_25825);
or U26157 (N_26157,N_25813,N_25827);
xor U26158 (N_26158,N_25893,N_26050);
and U26159 (N_26159,N_25873,N_25993);
xnor U26160 (N_26160,N_26026,N_25862);
and U26161 (N_26161,N_25974,N_25966);
nand U26162 (N_26162,N_25880,N_26070);
nor U26163 (N_26163,N_25962,N_25824);
xnor U26164 (N_26164,N_25866,N_25887);
or U26165 (N_26165,N_26013,N_25989);
nor U26166 (N_26166,N_25901,N_25969);
or U26167 (N_26167,N_25839,N_25850);
or U26168 (N_26168,N_25946,N_25930);
nand U26169 (N_26169,N_25832,N_26088);
or U26170 (N_26170,N_25885,N_25920);
nor U26171 (N_26171,N_25855,N_26003);
xor U26172 (N_26172,N_26079,N_25831);
xnor U26173 (N_26173,N_26002,N_25810);
nor U26174 (N_26174,N_25905,N_26015);
nor U26175 (N_26175,N_25952,N_25935);
nor U26176 (N_26176,N_25994,N_26089);
or U26177 (N_26177,N_26001,N_26007);
and U26178 (N_26178,N_25821,N_25819);
and U26179 (N_26179,N_25811,N_26073);
nand U26180 (N_26180,N_26043,N_26071);
or U26181 (N_26181,N_25992,N_25998);
nand U26182 (N_26182,N_25854,N_26031);
nor U26183 (N_26183,N_26042,N_25941);
and U26184 (N_26184,N_25876,N_25956);
and U26185 (N_26185,N_26078,N_25976);
nor U26186 (N_26186,N_25867,N_26056);
xor U26187 (N_26187,N_25884,N_25886);
nor U26188 (N_26188,N_25982,N_25967);
nor U26189 (N_26189,N_26018,N_26051);
nand U26190 (N_26190,N_26035,N_26060);
or U26191 (N_26191,N_25888,N_26066);
xnor U26192 (N_26192,N_26038,N_25970);
nand U26193 (N_26193,N_26052,N_26023);
xor U26194 (N_26194,N_25932,N_25815);
and U26195 (N_26195,N_25916,N_26091);
xor U26196 (N_26196,N_25818,N_25977);
or U26197 (N_26197,N_26081,N_25973);
nand U26198 (N_26198,N_26008,N_26096);
and U26199 (N_26199,N_26000,N_25928);
and U26200 (N_26200,N_25853,N_25869);
and U26201 (N_26201,N_25801,N_25835);
and U26202 (N_26202,N_25809,N_25874);
xor U26203 (N_26203,N_25852,N_25915);
and U26204 (N_26204,N_26030,N_26068);
nor U26205 (N_26205,N_25870,N_26014);
nand U26206 (N_26206,N_26061,N_25882);
and U26207 (N_26207,N_25999,N_26025);
xnor U26208 (N_26208,N_26020,N_25988);
nor U26209 (N_26209,N_25808,N_25812);
xnor U26210 (N_26210,N_26012,N_26063);
or U26211 (N_26211,N_26054,N_25986);
and U26212 (N_26212,N_25908,N_25860);
or U26213 (N_26213,N_26024,N_25943);
nor U26214 (N_26214,N_25996,N_25959);
or U26215 (N_26215,N_25985,N_25933);
xor U26216 (N_26216,N_25961,N_25847);
xor U26217 (N_26217,N_25804,N_25894);
and U26218 (N_26218,N_25895,N_26027);
or U26219 (N_26219,N_25917,N_25890);
xor U26220 (N_26220,N_25926,N_25978);
nand U26221 (N_26221,N_26074,N_25968);
or U26222 (N_26222,N_25924,N_26019);
xnor U26223 (N_26223,N_25900,N_25955);
or U26224 (N_26224,N_25859,N_25949);
nor U26225 (N_26225,N_25997,N_26086);
xor U26226 (N_26226,N_25987,N_25944);
nand U26227 (N_26227,N_25903,N_26072);
or U26228 (N_26228,N_25945,N_25942);
nor U26229 (N_26229,N_25995,N_25906);
and U26230 (N_26230,N_25807,N_25923);
or U26231 (N_26231,N_26016,N_26039);
nor U26232 (N_26232,N_25805,N_26006);
xnor U26233 (N_26233,N_26048,N_26049);
nand U26234 (N_26234,N_25910,N_26067);
or U26235 (N_26235,N_25802,N_25892);
or U26236 (N_26236,N_25849,N_26080);
and U26237 (N_26237,N_25927,N_25877);
nor U26238 (N_26238,N_26046,N_25836);
nor U26239 (N_26239,N_25958,N_26021);
and U26240 (N_26240,N_25868,N_25954);
and U26241 (N_26241,N_25953,N_25865);
nand U26242 (N_26242,N_25864,N_25899);
and U26243 (N_26243,N_25820,N_25816);
xor U26244 (N_26244,N_25979,N_26090);
xor U26245 (N_26245,N_26053,N_26085);
nor U26246 (N_26246,N_26094,N_25857);
or U26247 (N_26247,N_25907,N_25934);
and U26248 (N_26248,N_26032,N_25929);
nand U26249 (N_26249,N_25947,N_25881);
or U26250 (N_26250,N_26031,N_26065);
and U26251 (N_26251,N_26069,N_25956);
and U26252 (N_26252,N_26064,N_25949);
nand U26253 (N_26253,N_26007,N_25961);
nor U26254 (N_26254,N_25860,N_25867);
xnor U26255 (N_26255,N_26055,N_25931);
nand U26256 (N_26256,N_25941,N_25914);
xor U26257 (N_26257,N_25948,N_26065);
xnor U26258 (N_26258,N_25992,N_26048);
and U26259 (N_26259,N_26076,N_25870);
or U26260 (N_26260,N_25897,N_25962);
nand U26261 (N_26261,N_25965,N_26049);
xnor U26262 (N_26262,N_25939,N_26034);
and U26263 (N_26263,N_26096,N_25944);
or U26264 (N_26264,N_25864,N_25805);
nor U26265 (N_26265,N_26094,N_25865);
or U26266 (N_26266,N_26020,N_26098);
and U26267 (N_26267,N_25964,N_25976);
nand U26268 (N_26268,N_25868,N_25887);
or U26269 (N_26269,N_25809,N_25850);
nor U26270 (N_26270,N_25925,N_25995);
and U26271 (N_26271,N_25822,N_26078);
nand U26272 (N_26272,N_25994,N_25897);
and U26273 (N_26273,N_26052,N_26017);
or U26274 (N_26274,N_25961,N_26025);
and U26275 (N_26275,N_26055,N_25809);
or U26276 (N_26276,N_26001,N_25895);
nand U26277 (N_26277,N_25877,N_25955);
nor U26278 (N_26278,N_26037,N_25861);
and U26279 (N_26279,N_25892,N_26004);
nand U26280 (N_26280,N_25888,N_25960);
and U26281 (N_26281,N_25979,N_25934);
or U26282 (N_26282,N_26050,N_26080);
or U26283 (N_26283,N_25939,N_25899);
and U26284 (N_26284,N_26037,N_26087);
nor U26285 (N_26285,N_26023,N_25933);
or U26286 (N_26286,N_25972,N_25804);
nor U26287 (N_26287,N_26019,N_25998);
nor U26288 (N_26288,N_26091,N_26083);
and U26289 (N_26289,N_25974,N_26014);
and U26290 (N_26290,N_25961,N_25962);
or U26291 (N_26291,N_25949,N_26057);
xnor U26292 (N_26292,N_26032,N_25973);
xor U26293 (N_26293,N_25926,N_25949);
and U26294 (N_26294,N_25909,N_25840);
nor U26295 (N_26295,N_26050,N_25899);
nand U26296 (N_26296,N_25923,N_25973);
nand U26297 (N_26297,N_25800,N_26094);
or U26298 (N_26298,N_25934,N_25909);
or U26299 (N_26299,N_25912,N_25940);
xnor U26300 (N_26300,N_25860,N_25817);
nor U26301 (N_26301,N_25968,N_25954);
or U26302 (N_26302,N_25909,N_25914);
nor U26303 (N_26303,N_25914,N_25802);
nand U26304 (N_26304,N_25943,N_26015);
nand U26305 (N_26305,N_25940,N_25971);
xor U26306 (N_26306,N_25998,N_25945);
nand U26307 (N_26307,N_25940,N_25848);
nand U26308 (N_26308,N_25999,N_25942);
and U26309 (N_26309,N_26033,N_25930);
nor U26310 (N_26310,N_25840,N_25864);
nand U26311 (N_26311,N_25828,N_26012);
nor U26312 (N_26312,N_26070,N_25918);
or U26313 (N_26313,N_25906,N_25948);
xnor U26314 (N_26314,N_25947,N_25960);
and U26315 (N_26315,N_25953,N_26017);
xnor U26316 (N_26316,N_25893,N_25922);
xnor U26317 (N_26317,N_25848,N_25947);
and U26318 (N_26318,N_26022,N_26085);
or U26319 (N_26319,N_26046,N_26016);
nand U26320 (N_26320,N_25814,N_26082);
nor U26321 (N_26321,N_25830,N_25842);
nor U26322 (N_26322,N_25801,N_25896);
nor U26323 (N_26323,N_25924,N_25965);
nor U26324 (N_26324,N_25929,N_25933);
nor U26325 (N_26325,N_25946,N_25923);
nand U26326 (N_26326,N_26036,N_25862);
nand U26327 (N_26327,N_26069,N_26030);
and U26328 (N_26328,N_26080,N_26023);
nand U26329 (N_26329,N_26058,N_25842);
or U26330 (N_26330,N_25833,N_25851);
nand U26331 (N_26331,N_25836,N_25986);
nand U26332 (N_26332,N_25889,N_25910);
xnor U26333 (N_26333,N_26030,N_26024);
or U26334 (N_26334,N_25881,N_25889);
nor U26335 (N_26335,N_25978,N_25867);
nor U26336 (N_26336,N_25808,N_25948);
and U26337 (N_26337,N_25877,N_26056);
nand U26338 (N_26338,N_26063,N_25963);
xnor U26339 (N_26339,N_26031,N_26062);
xnor U26340 (N_26340,N_25851,N_25941);
xnor U26341 (N_26341,N_25826,N_25908);
xor U26342 (N_26342,N_25811,N_26021);
or U26343 (N_26343,N_25840,N_26004);
or U26344 (N_26344,N_26072,N_26097);
or U26345 (N_26345,N_25995,N_26047);
xor U26346 (N_26346,N_25984,N_25938);
nand U26347 (N_26347,N_25853,N_25816);
and U26348 (N_26348,N_25977,N_25997);
nand U26349 (N_26349,N_26097,N_25935);
and U26350 (N_26350,N_25865,N_25956);
or U26351 (N_26351,N_26034,N_25970);
xnor U26352 (N_26352,N_25848,N_25842);
nor U26353 (N_26353,N_25901,N_25995);
or U26354 (N_26354,N_26022,N_25825);
and U26355 (N_26355,N_25946,N_25925);
or U26356 (N_26356,N_26099,N_25818);
xor U26357 (N_26357,N_26019,N_25811);
nor U26358 (N_26358,N_26056,N_25811);
or U26359 (N_26359,N_25829,N_25870);
or U26360 (N_26360,N_25830,N_26052);
and U26361 (N_26361,N_26068,N_26052);
nor U26362 (N_26362,N_25923,N_25878);
and U26363 (N_26363,N_25999,N_26049);
nor U26364 (N_26364,N_25864,N_25967);
nand U26365 (N_26365,N_25995,N_25882);
nand U26366 (N_26366,N_25923,N_25977);
xor U26367 (N_26367,N_26011,N_25869);
and U26368 (N_26368,N_25973,N_25847);
and U26369 (N_26369,N_25993,N_25871);
or U26370 (N_26370,N_25910,N_25911);
or U26371 (N_26371,N_26039,N_25804);
and U26372 (N_26372,N_25877,N_25920);
nor U26373 (N_26373,N_25938,N_26062);
or U26374 (N_26374,N_25878,N_26054);
xor U26375 (N_26375,N_26035,N_25843);
nor U26376 (N_26376,N_25896,N_25982);
xor U26377 (N_26377,N_25941,N_25814);
nand U26378 (N_26378,N_25884,N_26017);
and U26379 (N_26379,N_25811,N_26020);
nor U26380 (N_26380,N_25812,N_25937);
xnor U26381 (N_26381,N_25903,N_25914);
and U26382 (N_26382,N_26023,N_25900);
or U26383 (N_26383,N_26039,N_25922);
nor U26384 (N_26384,N_25929,N_25851);
xnor U26385 (N_26385,N_26090,N_26033);
or U26386 (N_26386,N_25876,N_26033);
or U26387 (N_26387,N_25897,N_25928);
nand U26388 (N_26388,N_25814,N_26003);
xnor U26389 (N_26389,N_25945,N_26058);
xor U26390 (N_26390,N_26097,N_26096);
nor U26391 (N_26391,N_26061,N_25855);
nor U26392 (N_26392,N_25987,N_25966);
nor U26393 (N_26393,N_25975,N_25912);
nand U26394 (N_26394,N_25992,N_25806);
or U26395 (N_26395,N_25866,N_25891);
and U26396 (N_26396,N_25860,N_25950);
and U26397 (N_26397,N_26070,N_26014);
or U26398 (N_26398,N_25974,N_25990);
and U26399 (N_26399,N_26000,N_25982);
and U26400 (N_26400,N_26264,N_26139);
and U26401 (N_26401,N_26358,N_26321);
and U26402 (N_26402,N_26380,N_26303);
or U26403 (N_26403,N_26147,N_26235);
xnor U26404 (N_26404,N_26308,N_26111);
nand U26405 (N_26405,N_26337,N_26288);
or U26406 (N_26406,N_26226,N_26311);
xor U26407 (N_26407,N_26141,N_26307);
nor U26408 (N_26408,N_26172,N_26353);
and U26409 (N_26409,N_26394,N_26151);
and U26410 (N_26410,N_26241,N_26315);
nand U26411 (N_26411,N_26287,N_26290);
or U26412 (N_26412,N_26224,N_26312);
or U26413 (N_26413,N_26359,N_26239);
or U26414 (N_26414,N_26188,N_26165);
nor U26415 (N_26415,N_26360,N_26197);
nand U26416 (N_26416,N_26297,N_26325);
nor U26417 (N_26417,N_26101,N_26318);
or U26418 (N_26418,N_26142,N_26397);
nand U26419 (N_26419,N_26191,N_26250);
or U26420 (N_26420,N_26135,N_26374);
or U26421 (N_26421,N_26381,N_26334);
xnor U26422 (N_26422,N_26181,N_26278);
nand U26423 (N_26423,N_26301,N_26137);
xor U26424 (N_26424,N_26228,N_26396);
nand U26425 (N_26425,N_26193,N_26279);
and U26426 (N_26426,N_26116,N_26261);
and U26427 (N_26427,N_26236,N_26194);
xnor U26428 (N_26428,N_26268,N_26254);
or U26429 (N_26429,N_26158,N_26306);
xnor U26430 (N_26430,N_26136,N_26245);
nor U26431 (N_26431,N_26175,N_26146);
or U26432 (N_26432,N_26342,N_26190);
and U26433 (N_26433,N_26154,N_26294);
nand U26434 (N_26434,N_26187,N_26258);
xnor U26435 (N_26435,N_26350,N_26282);
nand U26436 (N_26436,N_26122,N_26382);
nor U26437 (N_26437,N_26300,N_26369);
and U26438 (N_26438,N_26157,N_26164);
and U26439 (N_26439,N_26395,N_26348);
xnor U26440 (N_26440,N_26257,N_26384);
nor U26441 (N_26441,N_26319,N_26199);
or U26442 (N_26442,N_26339,N_26206);
xnor U26443 (N_26443,N_26143,N_26133);
nor U26444 (N_26444,N_26285,N_26212);
nor U26445 (N_26445,N_26292,N_26159);
xnor U26446 (N_26446,N_26134,N_26113);
xor U26447 (N_26447,N_26115,N_26385);
nor U26448 (N_26448,N_26126,N_26262);
xnor U26449 (N_26449,N_26365,N_26291);
xnor U26450 (N_26450,N_26220,N_26232);
xor U26451 (N_26451,N_26244,N_26249);
xor U26452 (N_26452,N_26240,N_26148);
and U26453 (N_26453,N_26121,N_26336);
nand U26454 (N_26454,N_26377,N_26138);
nor U26455 (N_26455,N_26344,N_26209);
or U26456 (N_26456,N_26251,N_26378);
or U26457 (N_26457,N_26386,N_26296);
and U26458 (N_26458,N_26248,N_26345);
xnor U26459 (N_26459,N_26203,N_26373);
and U26460 (N_26460,N_26356,N_26320);
and U26461 (N_26461,N_26354,N_26340);
and U26462 (N_26462,N_26144,N_26218);
nor U26463 (N_26463,N_26332,N_26343);
or U26464 (N_26464,N_26280,N_26265);
and U26465 (N_26465,N_26202,N_26184);
nor U26466 (N_26466,N_26341,N_26119);
xnor U26467 (N_26467,N_26317,N_26379);
nor U26468 (N_26468,N_26346,N_26305);
nor U26469 (N_26469,N_26364,N_26120);
nor U26470 (N_26470,N_26256,N_26233);
xnor U26471 (N_26471,N_26140,N_26331);
xnor U26472 (N_26472,N_26326,N_26277);
nor U26473 (N_26473,N_26372,N_26180);
and U26474 (N_26474,N_26150,N_26329);
and U26475 (N_26475,N_26237,N_26231);
nor U26476 (N_26476,N_26129,N_26376);
nor U26477 (N_26477,N_26114,N_26309);
nand U26478 (N_26478,N_26182,N_26281);
and U26479 (N_26479,N_26189,N_26162);
and U26480 (N_26480,N_26124,N_26234);
nand U26481 (N_26481,N_26271,N_26152);
and U26482 (N_26482,N_26349,N_26272);
xnor U26483 (N_26483,N_26330,N_26351);
and U26484 (N_26484,N_26389,N_26263);
nor U26485 (N_26485,N_26167,N_26302);
or U26486 (N_26486,N_26171,N_26383);
nand U26487 (N_26487,N_26276,N_26183);
and U26488 (N_26488,N_26118,N_26217);
and U26489 (N_26489,N_26399,N_26112);
and U26490 (N_26490,N_26204,N_26156);
xor U26491 (N_26491,N_26253,N_26255);
nand U26492 (N_26492,N_26357,N_26108);
and U26493 (N_26493,N_26310,N_26299);
nor U26494 (N_26494,N_26392,N_26195);
nand U26495 (N_26495,N_26211,N_26117);
nor U26496 (N_26496,N_26375,N_26333);
and U26497 (N_26497,N_26313,N_26328);
or U26498 (N_26498,N_26273,N_26275);
or U26499 (N_26499,N_26100,N_26269);
nor U26500 (N_26500,N_26335,N_26252);
and U26501 (N_26501,N_26283,N_26106);
nor U26502 (N_26502,N_26366,N_26196);
nor U26503 (N_26503,N_26221,N_26208);
nand U26504 (N_26504,N_26390,N_26205);
nand U26505 (N_26505,N_26213,N_26223);
xnor U26506 (N_26506,N_26102,N_26131);
nand U26507 (N_26507,N_26370,N_26324);
xor U26508 (N_26508,N_26105,N_26127);
or U26509 (N_26509,N_26247,N_26214);
or U26510 (N_26510,N_26166,N_26266);
and U26511 (N_26511,N_26270,N_26179);
nor U26512 (N_26512,N_26145,N_26289);
xor U26513 (N_26513,N_26216,N_26323);
xnor U26514 (N_26514,N_26393,N_26125);
and U26515 (N_26515,N_26186,N_26178);
nand U26516 (N_26516,N_26243,N_26230);
or U26517 (N_26517,N_26293,N_26109);
xnor U26518 (N_26518,N_26173,N_26163);
or U26519 (N_26519,N_26314,N_26267);
and U26520 (N_26520,N_26185,N_26210);
and U26521 (N_26521,N_26123,N_26110);
nor U26522 (N_26522,N_26368,N_26170);
xnor U26523 (N_26523,N_26207,N_26169);
or U26524 (N_26524,N_26174,N_26362);
and U26525 (N_26525,N_26295,N_26192);
and U26526 (N_26526,N_26284,N_26388);
and U26527 (N_26527,N_26176,N_26149);
nand U26528 (N_26528,N_26227,N_26347);
and U26529 (N_26529,N_26316,N_26367);
nand U26530 (N_26530,N_26201,N_26215);
xor U26531 (N_26531,N_26161,N_26200);
nor U26532 (N_26532,N_26104,N_26198);
or U26533 (N_26533,N_26371,N_26177);
xnor U26534 (N_26534,N_26322,N_26355);
nor U26535 (N_26535,N_26260,N_26238);
nand U26536 (N_26536,N_26132,N_26363);
nor U26537 (N_26537,N_26387,N_26286);
and U26538 (N_26538,N_26160,N_26298);
nand U26539 (N_26539,N_26168,N_26274);
nand U26540 (N_26540,N_26361,N_26153);
or U26541 (N_26541,N_26391,N_26107);
xnor U26542 (N_26542,N_26219,N_26352);
and U26543 (N_26543,N_26246,N_26155);
xor U26544 (N_26544,N_26242,N_26128);
nand U26545 (N_26545,N_26222,N_26398);
xnor U26546 (N_26546,N_26103,N_26225);
nor U26547 (N_26547,N_26259,N_26304);
or U26548 (N_26548,N_26338,N_26327);
nor U26549 (N_26549,N_26130,N_26229);
or U26550 (N_26550,N_26297,N_26191);
or U26551 (N_26551,N_26122,N_26168);
and U26552 (N_26552,N_26126,N_26182);
nand U26553 (N_26553,N_26328,N_26398);
or U26554 (N_26554,N_26221,N_26381);
nand U26555 (N_26555,N_26188,N_26131);
nand U26556 (N_26556,N_26245,N_26379);
xor U26557 (N_26557,N_26355,N_26282);
or U26558 (N_26558,N_26160,N_26143);
nand U26559 (N_26559,N_26199,N_26355);
nand U26560 (N_26560,N_26166,N_26376);
and U26561 (N_26561,N_26271,N_26229);
or U26562 (N_26562,N_26386,N_26308);
or U26563 (N_26563,N_26161,N_26155);
and U26564 (N_26564,N_26292,N_26387);
nand U26565 (N_26565,N_26114,N_26233);
xnor U26566 (N_26566,N_26299,N_26385);
nor U26567 (N_26567,N_26230,N_26111);
and U26568 (N_26568,N_26160,N_26285);
xnor U26569 (N_26569,N_26109,N_26198);
and U26570 (N_26570,N_26108,N_26261);
nand U26571 (N_26571,N_26194,N_26337);
and U26572 (N_26572,N_26280,N_26328);
or U26573 (N_26573,N_26128,N_26250);
and U26574 (N_26574,N_26243,N_26303);
nand U26575 (N_26575,N_26387,N_26211);
nor U26576 (N_26576,N_26304,N_26217);
xor U26577 (N_26577,N_26394,N_26391);
nor U26578 (N_26578,N_26158,N_26398);
and U26579 (N_26579,N_26292,N_26319);
nor U26580 (N_26580,N_26287,N_26344);
nor U26581 (N_26581,N_26301,N_26326);
nor U26582 (N_26582,N_26369,N_26185);
nor U26583 (N_26583,N_26139,N_26165);
nor U26584 (N_26584,N_26254,N_26186);
xnor U26585 (N_26585,N_26144,N_26195);
and U26586 (N_26586,N_26334,N_26383);
xnor U26587 (N_26587,N_26333,N_26136);
nand U26588 (N_26588,N_26325,N_26267);
xor U26589 (N_26589,N_26220,N_26301);
nor U26590 (N_26590,N_26117,N_26185);
and U26591 (N_26591,N_26177,N_26220);
or U26592 (N_26592,N_26293,N_26180);
or U26593 (N_26593,N_26259,N_26265);
nand U26594 (N_26594,N_26187,N_26334);
xor U26595 (N_26595,N_26297,N_26117);
and U26596 (N_26596,N_26271,N_26325);
and U26597 (N_26597,N_26198,N_26295);
nor U26598 (N_26598,N_26182,N_26300);
xor U26599 (N_26599,N_26154,N_26135);
and U26600 (N_26600,N_26323,N_26349);
or U26601 (N_26601,N_26390,N_26392);
nor U26602 (N_26602,N_26307,N_26161);
nand U26603 (N_26603,N_26185,N_26172);
and U26604 (N_26604,N_26278,N_26129);
or U26605 (N_26605,N_26103,N_26117);
and U26606 (N_26606,N_26270,N_26353);
nand U26607 (N_26607,N_26296,N_26234);
or U26608 (N_26608,N_26148,N_26325);
and U26609 (N_26609,N_26132,N_26137);
nand U26610 (N_26610,N_26292,N_26196);
nand U26611 (N_26611,N_26156,N_26285);
nor U26612 (N_26612,N_26369,N_26200);
and U26613 (N_26613,N_26341,N_26333);
xor U26614 (N_26614,N_26330,N_26179);
or U26615 (N_26615,N_26260,N_26143);
or U26616 (N_26616,N_26185,N_26345);
or U26617 (N_26617,N_26278,N_26257);
xor U26618 (N_26618,N_26136,N_26131);
xnor U26619 (N_26619,N_26356,N_26228);
nor U26620 (N_26620,N_26309,N_26159);
or U26621 (N_26621,N_26351,N_26263);
xor U26622 (N_26622,N_26257,N_26123);
nor U26623 (N_26623,N_26336,N_26316);
and U26624 (N_26624,N_26188,N_26129);
nand U26625 (N_26625,N_26363,N_26339);
nand U26626 (N_26626,N_26345,N_26127);
and U26627 (N_26627,N_26265,N_26281);
xor U26628 (N_26628,N_26207,N_26242);
nor U26629 (N_26629,N_26266,N_26370);
xnor U26630 (N_26630,N_26138,N_26317);
nand U26631 (N_26631,N_26170,N_26306);
or U26632 (N_26632,N_26262,N_26245);
or U26633 (N_26633,N_26269,N_26274);
or U26634 (N_26634,N_26247,N_26125);
nand U26635 (N_26635,N_26240,N_26233);
or U26636 (N_26636,N_26133,N_26346);
and U26637 (N_26637,N_26282,N_26246);
or U26638 (N_26638,N_26295,N_26113);
nand U26639 (N_26639,N_26227,N_26373);
nand U26640 (N_26640,N_26131,N_26145);
nor U26641 (N_26641,N_26306,N_26395);
xnor U26642 (N_26642,N_26262,N_26382);
or U26643 (N_26643,N_26306,N_26264);
and U26644 (N_26644,N_26378,N_26380);
and U26645 (N_26645,N_26111,N_26156);
and U26646 (N_26646,N_26232,N_26124);
nand U26647 (N_26647,N_26127,N_26199);
xnor U26648 (N_26648,N_26138,N_26119);
and U26649 (N_26649,N_26193,N_26259);
nor U26650 (N_26650,N_26367,N_26305);
and U26651 (N_26651,N_26111,N_26344);
xnor U26652 (N_26652,N_26335,N_26379);
or U26653 (N_26653,N_26300,N_26363);
and U26654 (N_26654,N_26171,N_26390);
nand U26655 (N_26655,N_26360,N_26202);
or U26656 (N_26656,N_26342,N_26343);
nor U26657 (N_26657,N_26240,N_26336);
or U26658 (N_26658,N_26314,N_26108);
nand U26659 (N_26659,N_26208,N_26258);
or U26660 (N_26660,N_26203,N_26228);
and U26661 (N_26661,N_26376,N_26314);
xor U26662 (N_26662,N_26104,N_26263);
nand U26663 (N_26663,N_26241,N_26351);
xnor U26664 (N_26664,N_26358,N_26211);
nor U26665 (N_26665,N_26130,N_26294);
xnor U26666 (N_26666,N_26175,N_26108);
nand U26667 (N_26667,N_26194,N_26144);
nor U26668 (N_26668,N_26183,N_26358);
xnor U26669 (N_26669,N_26204,N_26308);
nand U26670 (N_26670,N_26352,N_26185);
and U26671 (N_26671,N_26235,N_26395);
or U26672 (N_26672,N_26194,N_26126);
or U26673 (N_26673,N_26324,N_26260);
and U26674 (N_26674,N_26293,N_26313);
nor U26675 (N_26675,N_26370,N_26373);
and U26676 (N_26676,N_26302,N_26385);
xor U26677 (N_26677,N_26358,N_26210);
nor U26678 (N_26678,N_26290,N_26271);
nor U26679 (N_26679,N_26222,N_26274);
nand U26680 (N_26680,N_26112,N_26288);
and U26681 (N_26681,N_26245,N_26200);
nor U26682 (N_26682,N_26150,N_26357);
and U26683 (N_26683,N_26276,N_26208);
or U26684 (N_26684,N_26382,N_26211);
nand U26685 (N_26685,N_26354,N_26328);
nor U26686 (N_26686,N_26348,N_26270);
nor U26687 (N_26687,N_26157,N_26188);
nand U26688 (N_26688,N_26185,N_26120);
nor U26689 (N_26689,N_26182,N_26313);
and U26690 (N_26690,N_26310,N_26236);
nor U26691 (N_26691,N_26338,N_26337);
xor U26692 (N_26692,N_26198,N_26312);
nor U26693 (N_26693,N_26326,N_26161);
nand U26694 (N_26694,N_26321,N_26263);
nand U26695 (N_26695,N_26353,N_26276);
nor U26696 (N_26696,N_26319,N_26356);
nand U26697 (N_26697,N_26219,N_26242);
or U26698 (N_26698,N_26213,N_26225);
nor U26699 (N_26699,N_26272,N_26274);
xor U26700 (N_26700,N_26665,N_26475);
nand U26701 (N_26701,N_26448,N_26485);
xnor U26702 (N_26702,N_26577,N_26453);
xor U26703 (N_26703,N_26596,N_26530);
xnor U26704 (N_26704,N_26604,N_26552);
and U26705 (N_26705,N_26652,N_26614);
xor U26706 (N_26706,N_26408,N_26633);
nor U26707 (N_26707,N_26463,N_26600);
nor U26708 (N_26708,N_26431,N_26519);
and U26709 (N_26709,N_26477,N_26660);
and U26710 (N_26710,N_26698,N_26570);
nand U26711 (N_26711,N_26677,N_26646);
nand U26712 (N_26712,N_26578,N_26581);
nand U26713 (N_26713,N_26502,N_26464);
xor U26714 (N_26714,N_26543,N_26678);
or U26715 (N_26715,N_26637,N_26617);
nor U26716 (N_26716,N_26440,N_26655);
nand U26717 (N_26717,N_26508,N_26610);
nand U26718 (N_26718,N_26564,N_26681);
and U26719 (N_26719,N_26631,N_26602);
nor U26720 (N_26720,N_26685,N_26683);
and U26721 (N_26721,N_26585,N_26662);
xnor U26722 (N_26722,N_26635,N_26470);
xnor U26723 (N_26723,N_26435,N_26620);
or U26724 (N_26724,N_26692,N_26471);
nand U26725 (N_26725,N_26406,N_26642);
and U26726 (N_26726,N_26480,N_26561);
and U26727 (N_26727,N_26673,N_26454);
or U26728 (N_26728,N_26414,N_26571);
nor U26729 (N_26729,N_26588,N_26648);
and U26730 (N_26730,N_26669,N_26419);
and U26731 (N_26731,N_26422,N_26627);
xnor U26732 (N_26732,N_26567,N_26636);
nand U26733 (N_26733,N_26534,N_26458);
xor U26734 (N_26734,N_26447,N_26616);
nand U26735 (N_26735,N_26659,N_26443);
xnor U26736 (N_26736,N_26533,N_26686);
nor U26737 (N_26737,N_26521,N_26695);
nand U26738 (N_26738,N_26689,N_26580);
nand U26739 (N_26739,N_26501,N_26668);
or U26740 (N_26740,N_26544,N_26489);
or U26741 (N_26741,N_26412,N_26444);
xor U26742 (N_26742,N_26615,N_26663);
xnor U26743 (N_26743,N_26514,N_26505);
xor U26744 (N_26744,N_26650,N_26675);
or U26745 (N_26745,N_26441,N_26584);
xor U26746 (N_26746,N_26640,N_26490);
nand U26747 (N_26747,N_26557,N_26476);
nor U26748 (N_26748,N_26403,N_26517);
xor U26749 (N_26749,N_26606,N_26539);
nand U26750 (N_26750,N_26455,N_26697);
and U26751 (N_26751,N_26432,N_26540);
and U26752 (N_26752,N_26638,N_26416);
or U26753 (N_26753,N_26449,N_26424);
xnor U26754 (N_26754,N_26528,N_26586);
and U26755 (N_26755,N_26644,N_26487);
nand U26756 (N_26756,N_26672,N_26522);
nand U26757 (N_26757,N_26684,N_26488);
nor U26758 (N_26758,N_26493,N_26651);
nor U26759 (N_26759,N_26495,N_26630);
and U26760 (N_26760,N_26647,N_26516);
and U26761 (N_26761,N_26503,N_26460);
or U26762 (N_26762,N_26573,N_26639);
or U26763 (N_26763,N_26601,N_26587);
or U26764 (N_26764,N_26507,N_26413);
xor U26765 (N_26765,N_26404,N_26434);
and U26766 (N_26766,N_26400,N_26468);
xor U26767 (N_26767,N_26452,N_26560);
nor U26768 (N_26768,N_26624,N_26531);
or U26769 (N_26769,N_26466,N_26520);
xor U26770 (N_26770,N_26595,N_26438);
xor U26771 (N_26771,N_26625,N_26559);
nor U26772 (N_26772,N_26538,N_26426);
and U26773 (N_26773,N_26603,N_26529);
nand U26774 (N_26774,N_26558,N_26696);
or U26775 (N_26775,N_26575,N_26457);
or U26776 (N_26776,N_26481,N_26688);
xnor U26777 (N_26777,N_26478,N_26591);
and U26778 (N_26778,N_26420,N_26609);
nand U26779 (N_26779,N_26428,N_26666);
nor U26780 (N_26780,N_26506,N_26445);
nand U26781 (N_26781,N_26486,N_26605);
or U26782 (N_26782,N_26437,N_26618);
nor U26783 (N_26783,N_26421,N_26459);
nand U26784 (N_26784,N_26546,N_26699);
nor U26785 (N_26785,N_26442,N_26583);
and U26786 (N_26786,N_26612,N_26439);
nor U26787 (N_26787,N_26563,N_26515);
nand U26788 (N_26788,N_26641,N_26497);
xor U26789 (N_26789,N_26611,N_26542);
xor U26790 (N_26790,N_26512,N_26430);
nand U26791 (N_26791,N_26411,N_26461);
nor U26792 (N_26792,N_26527,N_26518);
or U26793 (N_26793,N_26687,N_26425);
xor U26794 (N_26794,N_26451,N_26405);
xor U26795 (N_26795,N_26670,N_26550);
xor U26796 (N_26796,N_26579,N_26679);
or U26797 (N_26797,N_26491,N_26450);
and U26798 (N_26798,N_26417,N_26479);
and U26799 (N_26799,N_26654,N_26598);
xor U26800 (N_26800,N_26626,N_26658);
xnor U26801 (N_26801,N_26613,N_26496);
nand U26802 (N_26802,N_26657,N_26674);
or U26803 (N_26803,N_26467,N_26436);
xor U26804 (N_26804,N_26427,N_26694);
xnor U26805 (N_26805,N_26623,N_26525);
or U26806 (N_26806,N_26526,N_26593);
nand U26807 (N_26807,N_26597,N_26629);
nand U26808 (N_26808,N_26643,N_26667);
nor U26809 (N_26809,N_26645,N_26621);
nand U26810 (N_26810,N_26499,N_26498);
and U26811 (N_26811,N_26462,N_26511);
nor U26812 (N_26812,N_26682,N_26482);
and U26813 (N_26813,N_26649,N_26500);
or U26814 (N_26814,N_26456,N_26555);
xor U26815 (N_26815,N_26537,N_26566);
nor U26816 (N_26816,N_26628,N_26608);
xnor U26817 (N_26817,N_26509,N_26446);
nand U26818 (N_26818,N_26535,N_26599);
xor U26819 (N_26819,N_26569,N_26676);
and U26820 (N_26820,N_26553,N_26524);
xnor U26821 (N_26821,N_26590,N_26513);
xor U26822 (N_26822,N_26680,N_26619);
xor U26823 (N_26823,N_26474,N_26484);
or U26824 (N_26824,N_26661,N_26504);
or U26825 (N_26825,N_26592,N_26693);
nand U26826 (N_26826,N_26634,N_26473);
or U26827 (N_26827,N_26572,N_26589);
xnor U26828 (N_26828,N_26545,N_26691);
xnor U26829 (N_26829,N_26402,N_26418);
or U26830 (N_26830,N_26536,N_26532);
or U26831 (N_26831,N_26429,N_26469);
or U26832 (N_26832,N_26433,N_26656);
nand U26833 (N_26833,N_26548,N_26562);
nand U26834 (N_26834,N_26594,N_26410);
and U26835 (N_26835,N_26565,N_26492);
xor U26836 (N_26836,N_26554,N_26690);
nor U26837 (N_26837,N_26407,N_26494);
or U26838 (N_26838,N_26549,N_26551);
nand U26839 (N_26839,N_26576,N_26523);
or U26840 (N_26840,N_26664,N_26472);
and U26841 (N_26841,N_26582,N_26568);
nor U26842 (N_26842,N_26423,N_26653);
nor U26843 (N_26843,N_26547,N_26483);
nor U26844 (N_26844,N_26415,N_26574);
xnor U26845 (N_26845,N_26622,N_26556);
xnor U26846 (N_26846,N_26541,N_26607);
or U26847 (N_26847,N_26510,N_26401);
nor U26848 (N_26848,N_26465,N_26671);
xnor U26849 (N_26849,N_26632,N_26409);
nor U26850 (N_26850,N_26537,N_26447);
and U26851 (N_26851,N_26579,N_26564);
xor U26852 (N_26852,N_26608,N_26488);
nand U26853 (N_26853,N_26550,N_26598);
nor U26854 (N_26854,N_26624,N_26688);
nor U26855 (N_26855,N_26609,N_26496);
xor U26856 (N_26856,N_26564,N_26625);
nand U26857 (N_26857,N_26695,N_26417);
nor U26858 (N_26858,N_26535,N_26530);
nand U26859 (N_26859,N_26442,N_26511);
or U26860 (N_26860,N_26660,N_26441);
or U26861 (N_26861,N_26581,N_26523);
xor U26862 (N_26862,N_26535,N_26492);
xnor U26863 (N_26863,N_26670,N_26501);
xor U26864 (N_26864,N_26619,N_26413);
or U26865 (N_26865,N_26439,N_26533);
nand U26866 (N_26866,N_26442,N_26514);
nor U26867 (N_26867,N_26538,N_26683);
and U26868 (N_26868,N_26514,N_26664);
nand U26869 (N_26869,N_26532,N_26501);
nand U26870 (N_26870,N_26614,N_26431);
or U26871 (N_26871,N_26476,N_26559);
or U26872 (N_26872,N_26423,N_26475);
nor U26873 (N_26873,N_26453,N_26502);
nand U26874 (N_26874,N_26457,N_26439);
and U26875 (N_26875,N_26617,N_26433);
nand U26876 (N_26876,N_26419,N_26421);
xnor U26877 (N_26877,N_26585,N_26586);
nor U26878 (N_26878,N_26479,N_26411);
nand U26879 (N_26879,N_26637,N_26517);
or U26880 (N_26880,N_26424,N_26441);
nor U26881 (N_26881,N_26585,N_26618);
or U26882 (N_26882,N_26538,N_26478);
nand U26883 (N_26883,N_26621,N_26692);
xnor U26884 (N_26884,N_26555,N_26649);
nand U26885 (N_26885,N_26422,N_26536);
xnor U26886 (N_26886,N_26437,N_26538);
xor U26887 (N_26887,N_26515,N_26492);
nor U26888 (N_26888,N_26460,N_26607);
xor U26889 (N_26889,N_26600,N_26693);
or U26890 (N_26890,N_26675,N_26500);
xor U26891 (N_26891,N_26547,N_26419);
or U26892 (N_26892,N_26539,N_26595);
and U26893 (N_26893,N_26527,N_26456);
xnor U26894 (N_26894,N_26434,N_26483);
and U26895 (N_26895,N_26686,N_26637);
and U26896 (N_26896,N_26434,N_26417);
or U26897 (N_26897,N_26577,N_26558);
or U26898 (N_26898,N_26659,N_26668);
nor U26899 (N_26899,N_26623,N_26556);
nand U26900 (N_26900,N_26588,N_26463);
nand U26901 (N_26901,N_26473,N_26618);
xnor U26902 (N_26902,N_26544,N_26603);
nor U26903 (N_26903,N_26585,N_26563);
and U26904 (N_26904,N_26687,N_26567);
xor U26905 (N_26905,N_26494,N_26669);
xor U26906 (N_26906,N_26470,N_26614);
nand U26907 (N_26907,N_26670,N_26544);
or U26908 (N_26908,N_26523,N_26634);
and U26909 (N_26909,N_26604,N_26581);
or U26910 (N_26910,N_26528,N_26493);
nor U26911 (N_26911,N_26652,N_26622);
and U26912 (N_26912,N_26530,N_26683);
or U26913 (N_26913,N_26621,N_26580);
and U26914 (N_26914,N_26511,N_26422);
and U26915 (N_26915,N_26511,N_26519);
nand U26916 (N_26916,N_26590,N_26517);
nor U26917 (N_26917,N_26689,N_26631);
and U26918 (N_26918,N_26690,N_26406);
nor U26919 (N_26919,N_26504,N_26469);
or U26920 (N_26920,N_26608,N_26577);
or U26921 (N_26921,N_26446,N_26465);
nand U26922 (N_26922,N_26514,N_26609);
xor U26923 (N_26923,N_26433,N_26462);
xor U26924 (N_26924,N_26526,N_26642);
xor U26925 (N_26925,N_26527,N_26595);
or U26926 (N_26926,N_26410,N_26559);
and U26927 (N_26927,N_26657,N_26551);
nor U26928 (N_26928,N_26453,N_26673);
nand U26929 (N_26929,N_26456,N_26592);
xor U26930 (N_26930,N_26668,N_26642);
and U26931 (N_26931,N_26459,N_26597);
and U26932 (N_26932,N_26554,N_26600);
nand U26933 (N_26933,N_26650,N_26410);
nand U26934 (N_26934,N_26556,N_26592);
xor U26935 (N_26935,N_26414,N_26577);
or U26936 (N_26936,N_26590,N_26658);
nor U26937 (N_26937,N_26671,N_26525);
nor U26938 (N_26938,N_26672,N_26464);
nor U26939 (N_26939,N_26461,N_26522);
or U26940 (N_26940,N_26416,N_26685);
and U26941 (N_26941,N_26639,N_26490);
nand U26942 (N_26942,N_26628,N_26638);
xnor U26943 (N_26943,N_26585,N_26505);
nor U26944 (N_26944,N_26676,N_26656);
and U26945 (N_26945,N_26479,N_26673);
xnor U26946 (N_26946,N_26504,N_26520);
or U26947 (N_26947,N_26444,N_26445);
and U26948 (N_26948,N_26469,N_26534);
nand U26949 (N_26949,N_26438,N_26529);
xor U26950 (N_26950,N_26558,N_26576);
nand U26951 (N_26951,N_26605,N_26649);
and U26952 (N_26952,N_26585,N_26683);
and U26953 (N_26953,N_26687,N_26647);
nand U26954 (N_26954,N_26411,N_26664);
or U26955 (N_26955,N_26698,N_26687);
xnor U26956 (N_26956,N_26405,N_26442);
nor U26957 (N_26957,N_26648,N_26541);
nand U26958 (N_26958,N_26572,N_26674);
nor U26959 (N_26959,N_26446,N_26597);
or U26960 (N_26960,N_26408,N_26569);
or U26961 (N_26961,N_26418,N_26644);
nand U26962 (N_26962,N_26466,N_26690);
xnor U26963 (N_26963,N_26440,N_26651);
xor U26964 (N_26964,N_26524,N_26503);
xnor U26965 (N_26965,N_26596,N_26603);
nor U26966 (N_26966,N_26458,N_26484);
nor U26967 (N_26967,N_26680,N_26408);
nand U26968 (N_26968,N_26579,N_26572);
and U26969 (N_26969,N_26564,N_26476);
or U26970 (N_26970,N_26465,N_26546);
or U26971 (N_26971,N_26451,N_26642);
or U26972 (N_26972,N_26694,N_26487);
nor U26973 (N_26973,N_26533,N_26610);
nor U26974 (N_26974,N_26640,N_26592);
or U26975 (N_26975,N_26400,N_26625);
or U26976 (N_26976,N_26510,N_26429);
and U26977 (N_26977,N_26668,N_26686);
xnor U26978 (N_26978,N_26578,N_26556);
nor U26979 (N_26979,N_26516,N_26654);
or U26980 (N_26980,N_26477,N_26488);
or U26981 (N_26981,N_26459,N_26625);
and U26982 (N_26982,N_26502,N_26622);
nand U26983 (N_26983,N_26585,N_26555);
and U26984 (N_26984,N_26637,N_26586);
nor U26985 (N_26985,N_26402,N_26411);
nand U26986 (N_26986,N_26627,N_26461);
and U26987 (N_26987,N_26668,N_26685);
and U26988 (N_26988,N_26672,N_26539);
nand U26989 (N_26989,N_26692,N_26458);
nor U26990 (N_26990,N_26424,N_26446);
and U26991 (N_26991,N_26630,N_26509);
or U26992 (N_26992,N_26452,N_26651);
nor U26993 (N_26993,N_26567,N_26542);
nor U26994 (N_26994,N_26491,N_26667);
nor U26995 (N_26995,N_26694,N_26534);
nor U26996 (N_26996,N_26402,N_26538);
xor U26997 (N_26997,N_26475,N_26484);
xnor U26998 (N_26998,N_26621,N_26505);
nor U26999 (N_26999,N_26604,N_26658);
xnor U27000 (N_27000,N_26891,N_26755);
xor U27001 (N_27001,N_26995,N_26788);
or U27002 (N_27002,N_26779,N_26929);
xor U27003 (N_27003,N_26766,N_26876);
and U27004 (N_27004,N_26709,N_26863);
nor U27005 (N_27005,N_26729,N_26922);
and U27006 (N_27006,N_26809,N_26810);
nor U27007 (N_27007,N_26880,N_26912);
or U27008 (N_27008,N_26921,N_26910);
or U27009 (N_27009,N_26741,N_26881);
nand U27010 (N_27010,N_26996,N_26738);
nor U27011 (N_27011,N_26936,N_26923);
and U27012 (N_27012,N_26791,N_26903);
xor U27013 (N_27013,N_26953,N_26976);
or U27014 (N_27014,N_26890,N_26957);
and U27015 (N_27015,N_26836,N_26839);
nand U27016 (N_27016,N_26768,N_26928);
and U27017 (N_27017,N_26715,N_26843);
nand U27018 (N_27018,N_26799,N_26816);
xor U27019 (N_27019,N_26783,N_26900);
xor U27020 (N_27020,N_26974,N_26735);
xor U27021 (N_27021,N_26723,N_26968);
nand U27022 (N_27022,N_26823,N_26819);
nand U27023 (N_27023,N_26747,N_26972);
and U27024 (N_27024,N_26861,N_26961);
or U27025 (N_27025,N_26814,N_26800);
or U27026 (N_27026,N_26940,N_26776);
nand U27027 (N_27027,N_26969,N_26717);
or U27028 (N_27028,N_26785,N_26934);
or U27029 (N_27029,N_26721,N_26925);
and U27030 (N_27030,N_26727,N_26980);
nor U27031 (N_27031,N_26870,N_26857);
nor U27032 (N_27032,N_26872,N_26983);
nor U27033 (N_27033,N_26758,N_26999);
xnor U27034 (N_27034,N_26796,N_26885);
and U27035 (N_27035,N_26713,N_26977);
nor U27036 (N_27036,N_26984,N_26844);
xnor U27037 (N_27037,N_26965,N_26782);
xor U27038 (N_27038,N_26834,N_26896);
and U27039 (N_27039,N_26884,N_26720);
and U27040 (N_27040,N_26982,N_26949);
xnor U27041 (N_27041,N_26835,N_26798);
nor U27042 (N_27042,N_26710,N_26860);
and U27043 (N_27043,N_26726,N_26701);
xor U27044 (N_27044,N_26784,N_26750);
and U27045 (N_27045,N_26771,N_26821);
nor U27046 (N_27046,N_26852,N_26764);
or U27047 (N_27047,N_26963,N_26829);
or U27048 (N_27048,N_26842,N_26990);
or U27049 (N_27049,N_26793,N_26946);
or U27050 (N_27050,N_26743,N_26840);
or U27051 (N_27051,N_26975,N_26704);
or U27052 (N_27052,N_26959,N_26770);
or U27053 (N_27053,N_26989,N_26956);
xor U27054 (N_27054,N_26744,N_26892);
nand U27055 (N_27055,N_26952,N_26786);
and U27056 (N_27056,N_26871,N_26966);
xnor U27057 (N_27057,N_26873,N_26898);
xnor U27058 (N_27058,N_26858,N_26790);
nor U27059 (N_27059,N_26734,N_26932);
nand U27060 (N_27060,N_26967,N_26998);
xnor U27061 (N_27061,N_26777,N_26824);
xor U27062 (N_27062,N_26705,N_26894);
xor U27063 (N_27063,N_26862,N_26794);
xnor U27064 (N_27064,N_26825,N_26986);
nand U27065 (N_27065,N_26875,N_26907);
or U27066 (N_27066,N_26826,N_26933);
nor U27067 (N_27067,N_26981,N_26948);
nand U27068 (N_27068,N_26917,N_26935);
and U27069 (N_27069,N_26739,N_26908);
and U27070 (N_27070,N_26931,N_26728);
nor U27071 (N_27071,N_26769,N_26774);
nor U27072 (N_27072,N_26805,N_26702);
nor U27073 (N_27073,N_26937,N_26915);
xnor U27074 (N_27074,N_26848,N_26831);
nand U27075 (N_27075,N_26926,N_26781);
xor U27076 (N_27076,N_26939,N_26864);
or U27077 (N_27077,N_26944,N_26994);
xor U27078 (N_27078,N_26978,N_26869);
nand U27079 (N_27079,N_26817,N_26801);
xor U27080 (N_27080,N_26924,N_26751);
nor U27081 (N_27081,N_26833,N_26971);
nor U27082 (N_27082,N_26778,N_26979);
and U27083 (N_27083,N_26802,N_26792);
or U27084 (N_27084,N_26988,N_26754);
nand U27085 (N_27085,N_26832,N_26733);
nand U27086 (N_27086,N_26855,N_26913);
nand U27087 (N_27087,N_26893,N_26806);
nand U27088 (N_27088,N_26759,N_26987);
nand U27089 (N_27089,N_26901,N_26916);
nor U27090 (N_27090,N_26736,N_26760);
nor U27091 (N_27091,N_26943,N_26958);
nand U27092 (N_27092,N_26897,N_26945);
xnor U27093 (N_27093,N_26973,N_26828);
xor U27094 (N_27094,N_26763,N_26879);
nand U27095 (N_27095,N_26745,N_26938);
and U27096 (N_27096,N_26773,N_26849);
nand U27097 (N_27097,N_26712,N_26919);
xor U27098 (N_27098,N_26820,N_26740);
xor U27099 (N_27099,N_26950,N_26847);
nand U27100 (N_27100,N_26942,N_26737);
or U27101 (N_27101,N_26795,N_26889);
nor U27102 (N_27102,N_26748,N_26895);
nand U27103 (N_27103,N_26909,N_26762);
and U27104 (N_27104,N_26850,N_26882);
and U27105 (N_27105,N_26753,N_26993);
nor U27106 (N_27106,N_26811,N_26997);
or U27107 (N_27107,N_26886,N_26845);
or U27108 (N_27108,N_26808,N_26930);
xnor U27109 (N_27109,N_26731,N_26902);
nand U27110 (N_27110,N_26887,N_26920);
nor U27111 (N_27111,N_26964,N_26718);
xnor U27112 (N_27112,N_26724,N_26756);
or U27113 (N_27113,N_26991,N_26807);
or U27114 (N_27114,N_26767,N_26859);
xnor U27115 (N_27115,N_26866,N_26708);
nand U27116 (N_27116,N_26703,N_26761);
nand U27117 (N_27117,N_26877,N_26742);
and U27118 (N_27118,N_26927,N_26911);
xor U27119 (N_27119,N_26854,N_26706);
nand U27120 (N_27120,N_26757,N_26960);
nor U27121 (N_27121,N_26822,N_26904);
nand U27122 (N_27122,N_26780,N_26846);
nor U27123 (N_27123,N_26918,N_26837);
and U27124 (N_27124,N_26906,N_26730);
or U27125 (N_27125,N_26707,N_26700);
nand U27126 (N_27126,N_26874,N_26787);
or U27127 (N_27127,N_26827,N_26992);
and U27128 (N_27128,N_26841,N_26803);
or U27129 (N_27129,N_26804,N_26722);
nor U27130 (N_27130,N_26716,N_26789);
and U27131 (N_27131,N_26772,N_26732);
or U27132 (N_27132,N_26815,N_26954);
nand U27133 (N_27133,N_26725,N_26765);
or U27134 (N_27134,N_26818,N_26867);
nand U27135 (N_27135,N_26853,N_26714);
xor U27136 (N_27136,N_26941,N_26899);
nand U27137 (N_27137,N_26905,N_26962);
or U27138 (N_27138,N_26838,N_26856);
xor U27139 (N_27139,N_26947,N_26719);
or U27140 (N_27140,N_26746,N_26888);
and U27141 (N_27141,N_26812,N_26851);
nor U27142 (N_27142,N_26797,N_26775);
nor U27143 (N_27143,N_26914,N_26749);
or U27144 (N_27144,N_26830,N_26970);
and U27145 (N_27145,N_26865,N_26883);
and U27146 (N_27146,N_26813,N_26955);
and U27147 (N_27147,N_26878,N_26868);
or U27148 (N_27148,N_26752,N_26951);
nor U27149 (N_27149,N_26711,N_26985);
xnor U27150 (N_27150,N_26920,N_26791);
and U27151 (N_27151,N_26986,N_26922);
xor U27152 (N_27152,N_26942,N_26716);
and U27153 (N_27153,N_26853,N_26918);
xor U27154 (N_27154,N_26921,N_26760);
nor U27155 (N_27155,N_26919,N_26928);
or U27156 (N_27156,N_26706,N_26882);
and U27157 (N_27157,N_26869,N_26800);
nand U27158 (N_27158,N_26965,N_26960);
nor U27159 (N_27159,N_26750,N_26944);
nor U27160 (N_27160,N_26792,N_26975);
nand U27161 (N_27161,N_26781,N_26711);
nor U27162 (N_27162,N_26876,N_26924);
nor U27163 (N_27163,N_26716,N_26916);
nand U27164 (N_27164,N_26747,N_26845);
xnor U27165 (N_27165,N_26875,N_26845);
or U27166 (N_27166,N_26821,N_26924);
or U27167 (N_27167,N_26759,N_26852);
and U27168 (N_27168,N_26965,N_26700);
nor U27169 (N_27169,N_26775,N_26764);
nor U27170 (N_27170,N_26719,N_26761);
nand U27171 (N_27171,N_26713,N_26874);
nor U27172 (N_27172,N_26889,N_26727);
nand U27173 (N_27173,N_26849,N_26889);
nand U27174 (N_27174,N_26805,N_26874);
nor U27175 (N_27175,N_26948,N_26808);
xor U27176 (N_27176,N_26772,N_26962);
nand U27177 (N_27177,N_26987,N_26926);
xor U27178 (N_27178,N_26783,N_26749);
nand U27179 (N_27179,N_26870,N_26804);
nor U27180 (N_27180,N_26810,N_26874);
nor U27181 (N_27181,N_26984,N_26986);
and U27182 (N_27182,N_26779,N_26962);
xor U27183 (N_27183,N_26973,N_26781);
nand U27184 (N_27184,N_26783,N_26748);
or U27185 (N_27185,N_26727,N_26770);
and U27186 (N_27186,N_26745,N_26865);
nand U27187 (N_27187,N_26802,N_26930);
xor U27188 (N_27188,N_26986,N_26930);
or U27189 (N_27189,N_26741,N_26836);
xor U27190 (N_27190,N_26917,N_26746);
and U27191 (N_27191,N_26892,N_26770);
nor U27192 (N_27192,N_26898,N_26989);
nand U27193 (N_27193,N_26845,N_26918);
and U27194 (N_27194,N_26749,N_26983);
nand U27195 (N_27195,N_26799,N_26925);
and U27196 (N_27196,N_26841,N_26739);
nand U27197 (N_27197,N_26839,N_26947);
and U27198 (N_27198,N_26886,N_26940);
and U27199 (N_27199,N_26741,N_26964);
nor U27200 (N_27200,N_26949,N_26793);
xnor U27201 (N_27201,N_26801,N_26888);
or U27202 (N_27202,N_26776,N_26937);
and U27203 (N_27203,N_26887,N_26916);
nor U27204 (N_27204,N_26967,N_26843);
nand U27205 (N_27205,N_26874,N_26946);
nand U27206 (N_27206,N_26753,N_26889);
nand U27207 (N_27207,N_26858,N_26872);
nor U27208 (N_27208,N_26866,N_26795);
xor U27209 (N_27209,N_26838,N_26758);
xor U27210 (N_27210,N_26812,N_26901);
and U27211 (N_27211,N_26958,N_26723);
nor U27212 (N_27212,N_26759,N_26789);
and U27213 (N_27213,N_26782,N_26978);
and U27214 (N_27214,N_26776,N_26898);
nand U27215 (N_27215,N_26765,N_26999);
nor U27216 (N_27216,N_26906,N_26761);
xor U27217 (N_27217,N_26965,N_26815);
xnor U27218 (N_27218,N_26830,N_26899);
or U27219 (N_27219,N_26924,N_26954);
xor U27220 (N_27220,N_26864,N_26753);
nand U27221 (N_27221,N_26859,N_26889);
xnor U27222 (N_27222,N_26913,N_26917);
and U27223 (N_27223,N_26951,N_26974);
nor U27224 (N_27224,N_26897,N_26921);
and U27225 (N_27225,N_26904,N_26907);
xnor U27226 (N_27226,N_26863,N_26935);
or U27227 (N_27227,N_26920,N_26948);
nor U27228 (N_27228,N_26765,N_26745);
xnor U27229 (N_27229,N_26910,N_26856);
nand U27230 (N_27230,N_26969,N_26900);
xnor U27231 (N_27231,N_26833,N_26738);
nand U27232 (N_27232,N_26893,N_26984);
xor U27233 (N_27233,N_26990,N_26947);
xor U27234 (N_27234,N_26704,N_26868);
nor U27235 (N_27235,N_26974,N_26834);
xnor U27236 (N_27236,N_26836,N_26936);
nand U27237 (N_27237,N_26889,N_26950);
nand U27238 (N_27238,N_26713,N_26980);
or U27239 (N_27239,N_26844,N_26812);
nand U27240 (N_27240,N_26798,N_26706);
nand U27241 (N_27241,N_26765,N_26851);
and U27242 (N_27242,N_26721,N_26778);
nor U27243 (N_27243,N_26871,N_26769);
and U27244 (N_27244,N_26869,N_26936);
and U27245 (N_27245,N_26704,N_26852);
and U27246 (N_27246,N_26798,N_26803);
nand U27247 (N_27247,N_26853,N_26998);
nor U27248 (N_27248,N_26828,N_26809);
or U27249 (N_27249,N_26839,N_26881);
nand U27250 (N_27250,N_26848,N_26815);
xor U27251 (N_27251,N_26807,N_26769);
nor U27252 (N_27252,N_26955,N_26863);
nor U27253 (N_27253,N_26852,N_26831);
and U27254 (N_27254,N_26894,N_26980);
xnor U27255 (N_27255,N_26770,N_26914);
nor U27256 (N_27256,N_26991,N_26781);
and U27257 (N_27257,N_26969,N_26975);
or U27258 (N_27258,N_26893,N_26745);
nor U27259 (N_27259,N_26723,N_26805);
nor U27260 (N_27260,N_26707,N_26956);
nand U27261 (N_27261,N_26967,N_26996);
and U27262 (N_27262,N_26910,N_26768);
nor U27263 (N_27263,N_26943,N_26969);
and U27264 (N_27264,N_26822,N_26781);
xnor U27265 (N_27265,N_26975,N_26765);
xor U27266 (N_27266,N_26751,N_26899);
nand U27267 (N_27267,N_26745,N_26719);
and U27268 (N_27268,N_26857,N_26954);
or U27269 (N_27269,N_26713,N_26701);
nor U27270 (N_27270,N_26911,N_26989);
or U27271 (N_27271,N_26921,N_26935);
xor U27272 (N_27272,N_26934,N_26945);
xnor U27273 (N_27273,N_26884,N_26843);
nor U27274 (N_27274,N_26835,N_26913);
xor U27275 (N_27275,N_26787,N_26955);
xnor U27276 (N_27276,N_26921,N_26920);
or U27277 (N_27277,N_26702,N_26920);
nand U27278 (N_27278,N_26820,N_26968);
or U27279 (N_27279,N_26758,N_26945);
nor U27280 (N_27280,N_26937,N_26770);
and U27281 (N_27281,N_26968,N_26894);
nand U27282 (N_27282,N_26828,N_26743);
or U27283 (N_27283,N_26976,N_26752);
nor U27284 (N_27284,N_26978,N_26824);
or U27285 (N_27285,N_26948,N_26850);
xor U27286 (N_27286,N_26710,N_26953);
nand U27287 (N_27287,N_26781,N_26813);
and U27288 (N_27288,N_26924,N_26893);
xor U27289 (N_27289,N_26935,N_26868);
nor U27290 (N_27290,N_26969,N_26868);
or U27291 (N_27291,N_26868,N_26785);
nand U27292 (N_27292,N_26824,N_26965);
nand U27293 (N_27293,N_26768,N_26740);
or U27294 (N_27294,N_26824,N_26759);
and U27295 (N_27295,N_26825,N_26720);
xnor U27296 (N_27296,N_26761,N_26878);
xnor U27297 (N_27297,N_26828,N_26908);
nand U27298 (N_27298,N_26863,N_26741);
xor U27299 (N_27299,N_26989,N_26831);
and U27300 (N_27300,N_27111,N_27092);
nand U27301 (N_27301,N_27235,N_27025);
nand U27302 (N_27302,N_27272,N_27236);
nor U27303 (N_27303,N_27043,N_27081);
and U27304 (N_27304,N_27223,N_27296);
nand U27305 (N_27305,N_27060,N_27156);
xor U27306 (N_27306,N_27159,N_27200);
or U27307 (N_27307,N_27281,N_27102);
nor U27308 (N_27308,N_27196,N_27105);
nand U27309 (N_27309,N_27153,N_27085);
nor U27310 (N_27310,N_27206,N_27001);
and U27311 (N_27311,N_27163,N_27195);
or U27312 (N_27312,N_27276,N_27101);
and U27313 (N_27313,N_27000,N_27120);
nor U27314 (N_27314,N_27160,N_27286);
and U27315 (N_27315,N_27169,N_27215);
or U27316 (N_27316,N_27263,N_27265);
and U27317 (N_27317,N_27173,N_27007);
nand U27318 (N_27318,N_27142,N_27044);
nor U27319 (N_27319,N_27175,N_27230);
xnor U27320 (N_27320,N_27192,N_27246);
nor U27321 (N_27321,N_27069,N_27259);
or U27322 (N_27322,N_27010,N_27190);
and U27323 (N_27323,N_27139,N_27151);
and U27324 (N_27324,N_27182,N_27046);
or U27325 (N_27325,N_27034,N_27017);
nand U27326 (N_27326,N_27002,N_27035);
xnor U27327 (N_27327,N_27213,N_27064);
and U27328 (N_27328,N_27157,N_27149);
and U27329 (N_27329,N_27199,N_27298);
xor U27330 (N_27330,N_27185,N_27146);
or U27331 (N_27331,N_27077,N_27197);
nor U27332 (N_27332,N_27242,N_27261);
and U27333 (N_27333,N_27042,N_27022);
and U27334 (N_27334,N_27125,N_27019);
nor U27335 (N_27335,N_27250,N_27198);
nand U27336 (N_27336,N_27145,N_27273);
or U27337 (N_27337,N_27073,N_27088);
and U27338 (N_27338,N_27245,N_27112);
nor U27339 (N_27339,N_27224,N_27015);
nor U27340 (N_27340,N_27264,N_27154);
xnor U27341 (N_27341,N_27033,N_27098);
nor U27342 (N_27342,N_27288,N_27084);
xor U27343 (N_27343,N_27283,N_27114);
and U27344 (N_27344,N_27205,N_27058);
or U27345 (N_27345,N_27030,N_27228);
xnor U27346 (N_27346,N_27227,N_27082);
or U27347 (N_27347,N_27152,N_27179);
or U27348 (N_27348,N_27115,N_27277);
nor U27349 (N_27349,N_27251,N_27148);
nand U27350 (N_27350,N_27067,N_27091);
nand U27351 (N_27351,N_27018,N_27027);
xor U27352 (N_27352,N_27109,N_27248);
xor U27353 (N_27353,N_27123,N_27254);
or U27354 (N_27354,N_27055,N_27278);
and U27355 (N_27355,N_27141,N_27008);
nor U27356 (N_27356,N_27217,N_27174);
or U27357 (N_27357,N_27255,N_27048);
xor U27358 (N_27358,N_27121,N_27041);
or U27359 (N_27359,N_27134,N_27078);
nand U27360 (N_27360,N_27062,N_27188);
nor U27361 (N_27361,N_27292,N_27130);
xor U27362 (N_27362,N_27032,N_27066);
and U27363 (N_27363,N_27194,N_27012);
or U27364 (N_27364,N_27118,N_27260);
xnor U27365 (N_27365,N_27257,N_27222);
nand U27366 (N_27366,N_27168,N_27210);
nor U27367 (N_27367,N_27214,N_27167);
nor U27368 (N_27368,N_27226,N_27268);
and U27369 (N_27369,N_27212,N_27221);
nand U27370 (N_27370,N_27014,N_27143);
nand U27371 (N_27371,N_27104,N_27056);
xnor U27372 (N_27372,N_27119,N_27057);
and U27373 (N_27373,N_27220,N_27158);
nor U27374 (N_27374,N_27021,N_27285);
nand U27375 (N_27375,N_27295,N_27150);
nor U27376 (N_27376,N_27216,N_27280);
xnor U27377 (N_27377,N_27171,N_27234);
nand U27378 (N_27378,N_27103,N_27016);
xnor U27379 (N_27379,N_27093,N_27170);
nor U27380 (N_27380,N_27207,N_27100);
or U27381 (N_27381,N_27026,N_27229);
nor U27382 (N_27382,N_27036,N_27079);
xnor U27383 (N_27383,N_27178,N_27266);
and U27384 (N_27384,N_27039,N_27267);
nor U27385 (N_27385,N_27133,N_27045);
xor U27386 (N_27386,N_27193,N_27040);
and U27387 (N_27387,N_27244,N_27166);
and U27388 (N_27388,N_27291,N_27243);
xnor U27389 (N_27389,N_27061,N_27049);
and U27390 (N_27390,N_27051,N_27128);
and U27391 (N_27391,N_27090,N_27293);
and U27392 (N_27392,N_27024,N_27172);
nor U27393 (N_27393,N_27071,N_27053);
nor U27394 (N_27394,N_27063,N_27252);
and U27395 (N_27395,N_27209,N_27225);
nor U27396 (N_27396,N_27155,N_27237);
nor U27397 (N_27397,N_27116,N_27097);
and U27398 (N_27398,N_27106,N_27140);
or U27399 (N_27399,N_27031,N_27136);
nand U27400 (N_27400,N_27165,N_27003);
or U27401 (N_27401,N_27274,N_27023);
nor U27402 (N_27402,N_27191,N_27038);
or U27403 (N_27403,N_27147,N_27270);
nor U27404 (N_27404,N_27284,N_27068);
nor U27405 (N_27405,N_27240,N_27122);
and U27406 (N_27406,N_27028,N_27294);
or U27407 (N_27407,N_27181,N_27287);
nor U27408 (N_27408,N_27297,N_27162);
and U27409 (N_27409,N_27074,N_27211);
or U27410 (N_27410,N_27177,N_27013);
or U27411 (N_27411,N_27059,N_27087);
xor U27412 (N_27412,N_27117,N_27131);
and U27413 (N_27413,N_27204,N_27164);
or U27414 (N_27414,N_27258,N_27075);
xnor U27415 (N_27415,N_27233,N_27269);
xnor U27416 (N_27416,N_27011,N_27138);
nand U27417 (N_27417,N_27020,N_27072);
or U27418 (N_27418,N_27203,N_27065);
or U27419 (N_27419,N_27275,N_27232);
nor U27420 (N_27420,N_27247,N_27189);
and U27421 (N_27421,N_27187,N_27253);
or U27422 (N_27422,N_27184,N_27107);
nand U27423 (N_27423,N_27004,N_27201);
nand U27424 (N_27424,N_27238,N_27108);
nand U27425 (N_27425,N_27070,N_27099);
and U27426 (N_27426,N_27239,N_27262);
and U27427 (N_27427,N_27290,N_27129);
xor U27428 (N_27428,N_27132,N_27289);
or U27429 (N_27429,N_27127,N_27096);
xor U27430 (N_27430,N_27202,N_27110);
nor U27431 (N_27431,N_27208,N_27126);
or U27432 (N_27432,N_27249,N_27135);
nand U27433 (N_27433,N_27029,N_27089);
or U27434 (N_27434,N_27271,N_27095);
or U27435 (N_27435,N_27218,N_27094);
nor U27436 (N_27436,N_27054,N_27047);
xnor U27437 (N_27437,N_27006,N_27144);
and U27438 (N_27438,N_27076,N_27005);
and U27439 (N_27439,N_27050,N_27183);
xor U27440 (N_27440,N_27009,N_27113);
and U27441 (N_27441,N_27186,N_27052);
nor U27442 (N_27442,N_27241,N_27086);
nand U27443 (N_27443,N_27137,N_27219);
or U27444 (N_27444,N_27180,N_27083);
nor U27445 (N_27445,N_27124,N_27176);
nor U27446 (N_27446,N_27080,N_27161);
and U27447 (N_27447,N_27279,N_27256);
nor U27448 (N_27448,N_27231,N_27299);
nor U27449 (N_27449,N_27282,N_27037);
nand U27450 (N_27450,N_27227,N_27253);
xor U27451 (N_27451,N_27179,N_27070);
or U27452 (N_27452,N_27062,N_27224);
nor U27453 (N_27453,N_27057,N_27031);
and U27454 (N_27454,N_27217,N_27092);
nor U27455 (N_27455,N_27131,N_27129);
nor U27456 (N_27456,N_27094,N_27102);
and U27457 (N_27457,N_27227,N_27097);
xnor U27458 (N_27458,N_27238,N_27098);
and U27459 (N_27459,N_27119,N_27156);
nor U27460 (N_27460,N_27182,N_27130);
and U27461 (N_27461,N_27247,N_27120);
nor U27462 (N_27462,N_27101,N_27024);
and U27463 (N_27463,N_27200,N_27038);
xnor U27464 (N_27464,N_27096,N_27289);
and U27465 (N_27465,N_27060,N_27280);
nor U27466 (N_27466,N_27226,N_27125);
xnor U27467 (N_27467,N_27119,N_27012);
and U27468 (N_27468,N_27217,N_27003);
nor U27469 (N_27469,N_27221,N_27162);
xnor U27470 (N_27470,N_27004,N_27103);
and U27471 (N_27471,N_27262,N_27172);
and U27472 (N_27472,N_27244,N_27071);
xor U27473 (N_27473,N_27210,N_27033);
nor U27474 (N_27474,N_27087,N_27134);
nor U27475 (N_27475,N_27003,N_27016);
xnor U27476 (N_27476,N_27040,N_27226);
and U27477 (N_27477,N_27194,N_27037);
nor U27478 (N_27478,N_27254,N_27050);
or U27479 (N_27479,N_27158,N_27078);
nand U27480 (N_27480,N_27074,N_27158);
nor U27481 (N_27481,N_27021,N_27075);
and U27482 (N_27482,N_27176,N_27033);
xnor U27483 (N_27483,N_27295,N_27117);
or U27484 (N_27484,N_27043,N_27072);
xnor U27485 (N_27485,N_27185,N_27067);
xnor U27486 (N_27486,N_27150,N_27267);
xnor U27487 (N_27487,N_27291,N_27081);
xnor U27488 (N_27488,N_27189,N_27282);
xor U27489 (N_27489,N_27224,N_27172);
or U27490 (N_27490,N_27076,N_27145);
nand U27491 (N_27491,N_27081,N_27064);
nand U27492 (N_27492,N_27201,N_27187);
nor U27493 (N_27493,N_27085,N_27002);
and U27494 (N_27494,N_27018,N_27262);
and U27495 (N_27495,N_27010,N_27297);
xor U27496 (N_27496,N_27299,N_27289);
nor U27497 (N_27497,N_27136,N_27115);
and U27498 (N_27498,N_27010,N_27113);
nand U27499 (N_27499,N_27231,N_27062);
nand U27500 (N_27500,N_27234,N_27260);
xor U27501 (N_27501,N_27202,N_27178);
and U27502 (N_27502,N_27080,N_27198);
nor U27503 (N_27503,N_27160,N_27240);
nand U27504 (N_27504,N_27119,N_27125);
nor U27505 (N_27505,N_27207,N_27180);
or U27506 (N_27506,N_27248,N_27205);
nor U27507 (N_27507,N_27175,N_27234);
nor U27508 (N_27508,N_27295,N_27163);
xor U27509 (N_27509,N_27235,N_27049);
xor U27510 (N_27510,N_27268,N_27293);
xor U27511 (N_27511,N_27029,N_27150);
or U27512 (N_27512,N_27280,N_27045);
nand U27513 (N_27513,N_27225,N_27182);
nand U27514 (N_27514,N_27221,N_27176);
nor U27515 (N_27515,N_27032,N_27101);
nor U27516 (N_27516,N_27093,N_27240);
and U27517 (N_27517,N_27286,N_27176);
xor U27518 (N_27518,N_27239,N_27057);
xor U27519 (N_27519,N_27040,N_27130);
or U27520 (N_27520,N_27031,N_27083);
or U27521 (N_27521,N_27206,N_27096);
nand U27522 (N_27522,N_27267,N_27250);
xor U27523 (N_27523,N_27223,N_27146);
nor U27524 (N_27524,N_27141,N_27220);
nand U27525 (N_27525,N_27197,N_27142);
or U27526 (N_27526,N_27205,N_27172);
or U27527 (N_27527,N_27173,N_27240);
or U27528 (N_27528,N_27256,N_27054);
nand U27529 (N_27529,N_27144,N_27272);
nand U27530 (N_27530,N_27019,N_27219);
nor U27531 (N_27531,N_27011,N_27246);
nor U27532 (N_27532,N_27137,N_27035);
or U27533 (N_27533,N_27088,N_27142);
or U27534 (N_27534,N_27111,N_27219);
nand U27535 (N_27535,N_27030,N_27248);
or U27536 (N_27536,N_27013,N_27032);
xnor U27537 (N_27537,N_27040,N_27147);
and U27538 (N_27538,N_27178,N_27113);
nand U27539 (N_27539,N_27267,N_27035);
nor U27540 (N_27540,N_27187,N_27016);
nor U27541 (N_27541,N_27290,N_27108);
nor U27542 (N_27542,N_27062,N_27261);
nand U27543 (N_27543,N_27130,N_27000);
nor U27544 (N_27544,N_27008,N_27137);
nand U27545 (N_27545,N_27089,N_27002);
or U27546 (N_27546,N_27200,N_27287);
nand U27547 (N_27547,N_27009,N_27058);
xnor U27548 (N_27548,N_27157,N_27003);
xnor U27549 (N_27549,N_27220,N_27249);
or U27550 (N_27550,N_27077,N_27248);
xor U27551 (N_27551,N_27155,N_27083);
xor U27552 (N_27552,N_27009,N_27028);
nor U27553 (N_27553,N_27268,N_27013);
nand U27554 (N_27554,N_27177,N_27112);
nand U27555 (N_27555,N_27115,N_27198);
or U27556 (N_27556,N_27188,N_27091);
xnor U27557 (N_27557,N_27269,N_27059);
or U27558 (N_27558,N_27279,N_27152);
or U27559 (N_27559,N_27123,N_27019);
and U27560 (N_27560,N_27229,N_27261);
nand U27561 (N_27561,N_27177,N_27187);
xnor U27562 (N_27562,N_27233,N_27140);
nand U27563 (N_27563,N_27233,N_27262);
xor U27564 (N_27564,N_27202,N_27191);
nand U27565 (N_27565,N_27197,N_27212);
and U27566 (N_27566,N_27000,N_27044);
xor U27567 (N_27567,N_27210,N_27261);
or U27568 (N_27568,N_27242,N_27200);
nand U27569 (N_27569,N_27262,N_27293);
and U27570 (N_27570,N_27125,N_27127);
or U27571 (N_27571,N_27225,N_27060);
nand U27572 (N_27572,N_27022,N_27155);
and U27573 (N_27573,N_27236,N_27270);
xnor U27574 (N_27574,N_27124,N_27010);
nor U27575 (N_27575,N_27294,N_27211);
and U27576 (N_27576,N_27073,N_27076);
xnor U27577 (N_27577,N_27173,N_27263);
or U27578 (N_27578,N_27119,N_27288);
and U27579 (N_27579,N_27224,N_27288);
and U27580 (N_27580,N_27014,N_27174);
xnor U27581 (N_27581,N_27268,N_27096);
nor U27582 (N_27582,N_27194,N_27261);
and U27583 (N_27583,N_27239,N_27234);
and U27584 (N_27584,N_27111,N_27147);
and U27585 (N_27585,N_27012,N_27206);
nor U27586 (N_27586,N_27014,N_27080);
nor U27587 (N_27587,N_27075,N_27023);
and U27588 (N_27588,N_27212,N_27037);
nor U27589 (N_27589,N_27026,N_27119);
or U27590 (N_27590,N_27062,N_27080);
and U27591 (N_27591,N_27206,N_27246);
or U27592 (N_27592,N_27202,N_27299);
nor U27593 (N_27593,N_27209,N_27126);
nor U27594 (N_27594,N_27062,N_27209);
nor U27595 (N_27595,N_27146,N_27009);
or U27596 (N_27596,N_27003,N_27033);
nor U27597 (N_27597,N_27252,N_27054);
xnor U27598 (N_27598,N_27134,N_27063);
nor U27599 (N_27599,N_27163,N_27013);
xor U27600 (N_27600,N_27538,N_27432);
and U27601 (N_27601,N_27544,N_27341);
and U27602 (N_27602,N_27469,N_27554);
xnor U27603 (N_27603,N_27418,N_27330);
nand U27604 (N_27604,N_27334,N_27521);
nor U27605 (N_27605,N_27468,N_27381);
nand U27606 (N_27606,N_27496,N_27587);
or U27607 (N_27607,N_27446,N_27370);
or U27608 (N_27608,N_27336,N_27421);
or U27609 (N_27609,N_27519,N_27357);
xnor U27610 (N_27610,N_27505,N_27362);
nand U27611 (N_27611,N_27358,N_27593);
nand U27612 (N_27612,N_27465,N_27414);
nor U27613 (N_27613,N_27597,N_27441);
nand U27614 (N_27614,N_27562,N_27591);
and U27615 (N_27615,N_27492,N_27348);
or U27616 (N_27616,N_27328,N_27471);
or U27617 (N_27617,N_27516,N_27371);
or U27618 (N_27618,N_27360,N_27489);
nand U27619 (N_27619,N_27514,N_27327);
or U27620 (N_27620,N_27460,N_27592);
and U27621 (N_27621,N_27488,N_27555);
or U27622 (N_27622,N_27596,N_27495);
xnor U27623 (N_27623,N_27531,N_27477);
nand U27624 (N_27624,N_27551,N_27445);
and U27625 (N_27625,N_27497,N_27543);
nand U27626 (N_27626,N_27518,N_27467);
and U27627 (N_27627,N_27494,N_27504);
and U27628 (N_27628,N_27572,N_27326);
and U27629 (N_27629,N_27479,N_27352);
and U27630 (N_27630,N_27561,N_27367);
or U27631 (N_27631,N_27510,N_27399);
or U27632 (N_27632,N_27383,N_27384);
nor U27633 (N_27633,N_27584,N_27335);
nor U27634 (N_27634,N_27458,N_27324);
nand U27635 (N_27635,N_27523,N_27337);
and U27636 (N_27636,N_27579,N_27410);
and U27637 (N_27637,N_27433,N_27396);
or U27638 (N_27638,N_27322,N_27306);
nor U27639 (N_27639,N_27339,N_27319);
nand U27640 (N_27640,N_27419,N_27595);
or U27641 (N_27641,N_27570,N_27547);
xor U27642 (N_27642,N_27301,N_27478);
and U27643 (N_27643,N_27407,N_27426);
xnor U27644 (N_27644,N_27487,N_27409);
nor U27645 (N_27645,N_27552,N_27411);
xor U27646 (N_27646,N_27463,N_27388);
xnor U27647 (N_27647,N_27361,N_27585);
or U27648 (N_27648,N_27567,N_27438);
and U27649 (N_27649,N_27484,N_27316);
xor U27650 (N_27650,N_27353,N_27573);
and U27651 (N_27651,N_27393,N_27375);
and U27652 (N_27652,N_27474,N_27372);
or U27653 (N_27653,N_27449,N_27338);
nand U27654 (N_27654,N_27356,N_27507);
and U27655 (N_27655,N_27303,N_27501);
nand U27656 (N_27656,N_27333,N_27502);
and U27657 (N_27657,N_27402,N_27434);
nand U27658 (N_27658,N_27534,N_27397);
and U27659 (N_27659,N_27586,N_27448);
xor U27660 (N_27660,N_27398,N_27440);
and U27661 (N_27661,N_27363,N_27320);
xor U27662 (N_27662,N_27345,N_27424);
xor U27663 (N_27663,N_27548,N_27373);
or U27664 (N_27664,N_27347,N_27447);
and U27665 (N_27665,N_27475,N_27574);
nand U27666 (N_27666,N_27311,N_27506);
and U27667 (N_27667,N_27493,N_27359);
and U27668 (N_27668,N_27473,N_27532);
xnor U27669 (N_27669,N_27527,N_27355);
nor U27670 (N_27670,N_27412,N_27366);
or U27671 (N_27671,N_27594,N_27485);
or U27672 (N_27672,N_27408,N_27550);
xor U27673 (N_27673,N_27325,N_27450);
or U27674 (N_27674,N_27389,N_27580);
or U27675 (N_27675,N_27329,N_27403);
and U27676 (N_27676,N_27420,N_27459);
xnor U27677 (N_27677,N_27546,N_27542);
nand U27678 (N_27678,N_27342,N_27553);
nand U27679 (N_27679,N_27526,N_27391);
xnor U27680 (N_27680,N_27582,N_27490);
or U27681 (N_27681,N_27598,N_27557);
nor U27682 (N_27682,N_27332,N_27380);
nor U27683 (N_27683,N_27503,N_27590);
or U27684 (N_27684,N_27340,N_27522);
xnor U27685 (N_27685,N_27472,N_27413);
nand U27686 (N_27686,N_27315,N_27323);
or U27687 (N_27687,N_27486,N_27365);
nand U27688 (N_27688,N_27377,N_27528);
or U27689 (N_27689,N_27578,N_27382);
nor U27690 (N_27690,N_27455,N_27431);
or U27691 (N_27691,N_27453,N_27308);
xor U27692 (N_27692,N_27321,N_27310);
nor U27693 (N_27693,N_27571,N_27539);
xnor U27694 (N_27694,N_27444,N_27351);
nor U27695 (N_27695,N_27566,N_27429);
nor U27696 (N_27696,N_27378,N_27482);
and U27697 (N_27697,N_27428,N_27442);
and U27698 (N_27698,N_27464,N_27457);
and U27699 (N_27699,N_27435,N_27530);
nand U27700 (N_27700,N_27525,N_27499);
nor U27701 (N_27701,N_27524,N_27443);
xor U27702 (N_27702,N_27451,N_27309);
xnor U27703 (N_27703,N_27512,N_27563);
nand U27704 (N_27704,N_27581,N_27576);
xor U27705 (N_27705,N_27535,N_27415);
nand U27706 (N_27706,N_27500,N_27318);
and U27707 (N_27707,N_27480,N_27498);
nor U27708 (N_27708,N_27394,N_27491);
xor U27709 (N_27709,N_27588,N_27390);
xnor U27710 (N_27710,N_27589,N_27520);
nand U27711 (N_27711,N_27314,N_27583);
nor U27712 (N_27712,N_27470,N_27476);
and U27713 (N_27713,N_27511,N_27483);
nand U27714 (N_27714,N_27346,N_27466);
or U27715 (N_27715,N_27564,N_27508);
and U27716 (N_27716,N_27374,N_27385);
or U27717 (N_27717,N_27461,N_27368);
and U27718 (N_27718,N_27545,N_27577);
xor U27719 (N_27719,N_27305,N_27416);
nand U27720 (N_27720,N_27556,N_27307);
and U27721 (N_27721,N_27513,N_27331);
xor U27722 (N_27722,N_27387,N_27515);
and U27723 (N_27723,N_27529,N_27568);
nand U27724 (N_27724,N_27313,N_27427);
nand U27725 (N_27725,N_27565,N_27575);
or U27726 (N_27726,N_27452,N_27379);
or U27727 (N_27727,N_27430,N_27456);
xor U27728 (N_27728,N_27406,N_27417);
nor U27729 (N_27729,N_27439,N_27509);
and U27730 (N_27730,N_27304,N_27560);
nor U27731 (N_27731,N_27537,N_27386);
nand U27732 (N_27732,N_27569,N_27354);
nor U27733 (N_27733,N_27454,N_27481);
or U27734 (N_27734,N_27405,N_27369);
nor U27735 (N_27735,N_27558,N_27423);
and U27736 (N_27736,N_27422,N_27350);
or U27737 (N_27737,N_27400,N_27462);
nor U27738 (N_27738,N_27395,N_27392);
xor U27739 (N_27739,N_27312,N_27401);
nand U27740 (N_27740,N_27425,N_27300);
xnor U27741 (N_27741,N_27364,N_27549);
or U27742 (N_27742,N_27599,N_27541);
nor U27743 (N_27743,N_27533,N_27343);
and U27744 (N_27744,N_27349,N_27559);
nand U27745 (N_27745,N_27317,N_27404);
xor U27746 (N_27746,N_27436,N_27540);
nand U27747 (N_27747,N_27376,N_27344);
nor U27748 (N_27748,N_27437,N_27536);
nand U27749 (N_27749,N_27302,N_27517);
nor U27750 (N_27750,N_27504,N_27338);
xor U27751 (N_27751,N_27596,N_27503);
nor U27752 (N_27752,N_27389,N_27357);
and U27753 (N_27753,N_27319,N_27568);
or U27754 (N_27754,N_27326,N_27444);
nand U27755 (N_27755,N_27421,N_27419);
and U27756 (N_27756,N_27488,N_27350);
nand U27757 (N_27757,N_27325,N_27402);
nor U27758 (N_27758,N_27309,N_27371);
nor U27759 (N_27759,N_27300,N_27537);
nor U27760 (N_27760,N_27338,N_27433);
and U27761 (N_27761,N_27435,N_27590);
nor U27762 (N_27762,N_27535,N_27338);
and U27763 (N_27763,N_27337,N_27391);
nor U27764 (N_27764,N_27517,N_27492);
and U27765 (N_27765,N_27553,N_27326);
nor U27766 (N_27766,N_27571,N_27588);
nand U27767 (N_27767,N_27442,N_27564);
xor U27768 (N_27768,N_27576,N_27451);
or U27769 (N_27769,N_27337,N_27316);
nand U27770 (N_27770,N_27407,N_27566);
nor U27771 (N_27771,N_27524,N_27426);
nor U27772 (N_27772,N_27478,N_27558);
xnor U27773 (N_27773,N_27555,N_27365);
or U27774 (N_27774,N_27457,N_27479);
and U27775 (N_27775,N_27520,N_27354);
and U27776 (N_27776,N_27339,N_27560);
or U27777 (N_27777,N_27361,N_27566);
nor U27778 (N_27778,N_27421,N_27364);
and U27779 (N_27779,N_27571,N_27466);
nand U27780 (N_27780,N_27477,N_27383);
nand U27781 (N_27781,N_27392,N_27330);
or U27782 (N_27782,N_27550,N_27466);
nor U27783 (N_27783,N_27552,N_27314);
nand U27784 (N_27784,N_27580,N_27515);
xor U27785 (N_27785,N_27544,N_27462);
xnor U27786 (N_27786,N_27428,N_27542);
or U27787 (N_27787,N_27320,N_27546);
nand U27788 (N_27788,N_27596,N_27561);
and U27789 (N_27789,N_27377,N_27454);
nand U27790 (N_27790,N_27411,N_27496);
nor U27791 (N_27791,N_27301,N_27482);
or U27792 (N_27792,N_27581,N_27386);
nand U27793 (N_27793,N_27509,N_27597);
or U27794 (N_27794,N_27502,N_27584);
nor U27795 (N_27795,N_27536,N_27459);
nand U27796 (N_27796,N_27576,N_27416);
nor U27797 (N_27797,N_27587,N_27579);
or U27798 (N_27798,N_27357,N_27561);
nand U27799 (N_27799,N_27547,N_27454);
xor U27800 (N_27800,N_27338,N_27315);
and U27801 (N_27801,N_27573,N_27499);
nor U27802 (N_27802,N_27325,N_27461);
xor U27803 (N_27803,N_27552,N_27448);
and U27804 (N_27804,N_27584,N_27407);
xnor U27805 (N_27805,N_27578,N_27476);
or U27806 (N_27806,N_27309,N_27329);
nor U27807 (N_27807,N_27348,N_27501);
and U27808 (N_27808,N_27383,N_27555);
or U27809 (N_27809,N_27332,N_27383);
nor U27810 (N_27810,N_27482,N_27346);
xnor U27811 (N_27811,N_27488,N_27430);
or U27812 (N_27812,N_27385,N_27540);
or U27813 (N_27813,N_27382,N_27354);
or U27814 (N_27814,N_27521,N_27329);
or U27815 (N_27815,N_27575,N_27501);
and U27816 (N_27816,N_27593,N_27448);
and U27817 (N_27817,N_27464,N_27590);
xor U27818 (N_27818,N_27360,N_27541);
and U27819 (N_27819,N_27412,N_27405);
and U27820 (N_27820,N_27315,N_27512);
and U27821 (N_27821,N_27546,N_27553);
or U27822 (N_27822,N_27407,N_27522);
or U27823 (N_27823,N_27585,N_27416);
and U27824 (N_27824,N_27424,N_27487);
nor U27825 (N_27825,N_27368,N_27478);
nor U27826 (N_27826,N_27504,N_27444);
or U27827 (N_27827,N_27430,N_27481);
nor U27828 (N_27828,N_27592,N_27521);
and U27829 (N_27829,N_27306,N_27515);
and U27830 (N_27830,N_27316,N_27383);
nor U27831 (N_27831,N_27303,N_27399);
nand U27832 (N_27832,N_27533,N_27576);
and U27833 (N_27833,N_27546,N_27537);
or U27834 (N_27834,N_27377,N_27498);
nor U27835 (N_27835,N_27584,N_27545);
xnor U27836 (N_27836,N_27375,N_27369);
and U27837 (N_27837,N_27392,N_27317);
nor U27838 (N_27838,N_27566,N_27462);
xor U27839 (N_27839,N_27559,N_27421);
nand U27840 (N_27840,N_27384,N_27584);
and U27841 (N_27841,N_27398,N_27360);
and U27842 (N_27842,N_27569,N_27481);
nor U27843 (N_27843,N_27506,N_27586);
xnor U27844 (N_27844,N_27345,N_27352);
nor U27845 (N_27845,N_27528,N_27595);
nor U27846 (N_27846,N_27520,N_27399);
or U27847 (N_27847,N_27443,N_27514);
nand U27848 (N_27848,N_27489,N_27341);
or U27849 (N_27849,N_27342,N_27346);
and U27850 (N_27850,N_27421,N_27324);
nand U27851 (N_27851,N_27430,N_27518);
or U27852 (N_27852,N_27584,N_27423);
xor U27853 (N_27853,N_27590,N_27570);
xnor U27854 (N_27854,N_27350,N_27304);
nand U27855 (N_27855,N_27444,N_27331);
or U27856 (N_27856,N_27523,N_27322);
xor U27857 (N_27857,N_27584,N_27304);
and U27858 (N_27858,N_27563,N_27515);
xnor U27859 (N_27859,N_27428,N_27595);
or U27860 (N_27860,N_27450,N_27594);
xnor U27861 (N_27861,N_27581,N_27356);
xor U27862 (N_27862,N_27588,N_27558);
nand U27863 (N_27863,N_27394,N_27335);
or U27864 (N_27864,N_27533,N_27564);
and U27865 (N_27865,N_27473,N_27536);
nor U27866 (N_27866,N_27363,N_27415);
and U27867 (N_27867,N_27432,N_27576);
xor U27868 (N_27868,N_27387,N_27353);
and U27869 (N_27869,N_27559,N_27555);
nand U27870 (N_27870,N_27467,N_27483);
nand U27871 (N_27871,N_27389,N_27398);
or U27872 (N_27872,N_27402,N_27486);
nand U27873 (N_27873,N_27522,N_27426);
nand U27874 (N_27874,N_27508,N_27578);
and U27875 (N_27875,N_27339,N_27318);
nand U27876 (N_27876,N_27484,N_27419);
and U27877 (N_27877,N_27336,N_27320);
or U27878 (N_27878,N_27438,N_27549);
xor U27879 (N_27879,N_27351,N_27486);
or U27880 (N_27880,N_27448,N_27300);
and U27881 (N_27881,N_27488,N_27455);
and U27882 (N_27882,N_27489,N_27385);
or U27883 (N_27883,N_27315,N_27358);
xor U27884 (N_27884,N_27585,N_27512);
or U27885 (N_27885,N_27578,N_27411);
nand U27886 (N_27886,N_27567,N_27326);
nor U27887 (N_27887,N_27490,N_27502);
xor U27888 (N_27888,N_27359,N_27594);
nand U27889 (N_27889,N_27335,N_27437);
nor U27890 (N_27890,N_27542,N_27408);
and U27891 (N_27891,N_27417,N_27460);
and U27892 (N_27892,N_27582,N_27321);
nor U27893 (N_27893,N_27583,N_27462);
nor U27894 (N_27894,N_27312,N_27578);
or U27895 (N_27895,N_27419,N_27504);
xor U27896 (N_27896,N_27310,N_27383);
nand U27897 (N_27897,N_27361,N_27438);
xnor U27898 (N_27898,N_27469,N_27491);
xnor U27899 (N_27899,N_27413,N_27427);
nor U27900 (N_27900,N_27796,N_27683);
nor U27901 (N_27901,N_27729,N_27859);
or U27902 (N_27902,N_27750,N_27813);
or U27903 (N_27903,N_27670,N_27697);
and U27904 (N_27904,N_27660,N_27869);
and U27905 (N_27905,N_27814,N_27792);
nor U27906 (N_27906,N_27627,N_27806);
xor U27907 (N_27907,N_27628,N_27632);
or U27908 (N_27908,N_27654,N_27773);
nor U27909 (N_27909,N_27802,N_27789);
nand U27910 (N_27910,N_27801,N_27688);
nand U27911 (N_27911,N_27701,N_27762);
and U27912 (N_27912,N_27676,N_27879);
and U27913 (N_27913,N_27799,N_27898);
xor U27914 (N_27914,N_27848,N_27610);
and U27915 (N_27915,N_27669,N_27817);
xnor U27916 (N_27916,N_27694,N_27605);
nand U27917 (N_27917,N_27795,N_27873);
xor U27918 (N_27918,N_27893,N_27691);
nor U27919 (N_27919,N_27874,N_27744);
xor U27920 (N_27920,N_27668,N_27888);
nor U27921 (N_27921,N_27643,N_27663);
nor U27922 (N_27922,N_27680,N_27649);
or U27923 (N_27923,N_27816,N_27764);
xnor U27924 (N_27924,N_27735,N_27889);
or U27925 (N_27925,N_27661,N_27656);
and U27926 (N_27926,N_27696,N_27788);
nor U27927 (N_27927,N_27720,N_27629);
nand U27928 (N_27928,N_27650,N_27768);
nand U27929 (N_27929,N_27844,N_27864);
xnor U27930 (N_27930,N_27853,N_27836);
and U27931 (N_27931,N_27602,N_27778);
or U27932 (N_27932,N_27785,N_27835);
nand U27933 (N_27933,N_27840,N_27739);
or U27934 (N_27934,N_27711,N_27876);
nand U27935 (N_27935,N_27830,N_27726);
and U27936 (N_27936,N_27636,N_27749);
xor U27937 (N_27937,N_27713,N_27615);
nor U27938 (N_27938,N_27678,N_27884);
and U27939 (N_27939,N_27863,N_27722);
or U27940 (N_27940,N_27761,N_27639);
nand U27941 (N_27941,N_27886,N_27779);
and U27942 (N_27942,N_27803,N_27699);
nand U27943 (N_27943,N_27686,N_27815);
nand U27944 (N_27944,N_27838,N_27890);
xor U27945 (N_27945,N_27793,N_27608);
nand U27946 (N_27946,N_27673,N_27737);
xor U27947 (N_27947,N_27777,N_27883);
or U27948 (N_27948,N_27652,N_27812);
nand U27949 (N_27949,N_27727,N_27679);
nand U27950 (N_27950,N_27756,N_27700);
or U27951 (N_27951,N_27646,N_27891);
and U27952 (N_27952,N_27871,N_27621);
or U27953 (N_27953,N_27870,N_27708);
or U27954 (N_27954,N_27709,N_27872);
xor U27955 (N_27955,N_27625,N_27635);
nand U27956 (N_27956,N_27877,N_27687);
nor U27957 (N_27957,N_27748,N_27841);
or U27958 (N_27958,N_27690,N_27774);
nand U27959 (N_27959,N_27707,N_27674);
xor U27960 (N_27960,N_27682,N_27800);
nand U27961 (N_27961,N_27854,N_27622);
or U27962 (N_27962,N_27832,N_27843);
nand U27963 (N_27963,N_27767,N_27822);
xor U27964 (N_27964,N_27892,N_27633);
nand U27965 (N_27965,N_27856,N_27759);
nand U27966 (N_27966,N_27651,N_27852);
nor U27967 (N_27967,N_27725,N_27703);
nand U27968 (N_27968,N_27810,N_27825);
nor U27969 (N_27969,N_27640,N_27780);
or U27970 (N_27970,N_27881,N_27783);
or U27971 (N_27971,N_27776,N_27689);
or U27972 (N_27972,N_27693,N_27619);
nor U27973 (N_27973,N_27834,N_27710);
nor U27974 (N_27974,N_27738,N_27657);
nand U27975 (N_27975,N_27772,N_27718);
nand U27976 (N_27976,N_27752,N_27823);
xnor U27977 (N_27977,N_27775,N_27769);
nand U27978 (N_27978,N_27623,N_27751);
nand U27979 (N_27979,N_27617,N_27645);
and U27980 (N_27980,N_27704,N_27862);
xor U27981 (N_27981,N_27833,N_27787);
nor U27982 (N_27982,N_27692,N_27644);
xor U27983 (N_27983,N_27827,N_27797);
nor U27984 (N_27984,N_27601,N_27765);
xnor U27985 (N_27985,N_27857,N_27706);
and U27986 (N_27986,N_27612,N_27638);
nor U27987 (N_27987,N_27790,N_27662);
or U27988 (N_27988,N_27717,N_27613);
and U27989 (N_27989,N_27745,N_27824);
nor U27990 (N_27990,N_27819,N_27732);
nor U27991 (N_27991,N_27715,N_27741);
and U27992 (N_27992,N_27845,N_27758);
nor U27993 (N_27993,N_27743,N_27821);
nor U27994 (N_27994,N_27698,N_27653);
and U27995 (N_27995,N_27866,N_27695);
xor U27996 (N_27996,N_27641,N_27648);
and U27997 (N_27997,N_27675,N_27808);
nand U27998 (N_27998,N_27637,N_27805);
xor U27999 (N_27999,N_27728,N_27664);
or U28000 (N_28000,N_27677,N_27734);
or U28001 (N_28001,N_27747,N_27626);
and U28002 (N_28002,N_27609,N_27634);
nand U28003 (N_28003,N_27614,N_27611);
and U28004 (N_28004,N_27826,N_27798);
nor U28005 (N_28005,N_27804,N_27736);
and U28006 (N_28006,N_27642,N_27894);
nor U28007 (N_28007,N_27897,N_27868);
nand U28008 (N_28008,N_27753,N_27733);
or U28009 (N_28009,N_27731,N_27714);
nand U28010 (N_28010,N_27624,N_27899);
xnor U28011 (N_28011,N_27766,N_27672);
and U28012 (N_28012,N_27716,N_27858);
nor U28013 (N_28013,N_27702,N_27807);
nand U28014 (N_28014,N_27665,N_27620);
and U28015 (N_28015,N_27828,N_27630);
nand U28016 (N_28016,N_27885,N_27880);
nand U28017 (N_28017,N_27771,N_27604);
nand U28018 (N_28018,N_27685,N_27820);
xor U28019 (N_28019,N_27754,N_27794);
xor U28020 (N_28020,N_27846,N_27875);
nand U28021 (N_28021,N_27860,N_27684);
nand U28022 (N_28022,N_27867,N_27666);
nand U28023 (N_28023,N_27763,N_27895);
xnor U28024 (N_28024,N_27755,N_27781);
or U28025 (N_28025,N_27746,N_27851);
and U28026 (N_28026,N_27659,N_27865);
nor U28027 (N_28027,N_27606,N_27631);
nand U28028 (N_28028,N_27809,N_27842);
or U28029 (N_28029,N_27724,N_27740);
or U28030 (N_28030,N_27831,N_27647);
xor U28031 (N_28031,N_27616,N_27618);
and U28032 (N_28032,N_27658,N_27818);
nand U28033 (N_28033,N_27600,N_27791);
nor U28034 (N_28034,N_27671,N_27847);
and U28035 (N_28035,N_27784,N_27850);
or U28036 (N_28036,N_27782,N_27667);
or U28037 (N_28037,N_27730,N_27770);
or U28038 (N_28038,N_27719,N_27861);
xor U28039 (N_28039,N_27607,N_27655);
or U28040 (N_28040,N_27855,N_27882);
nor U28041 (N_28041,N_27705,N_27723);
nor U28042 (N_28042,N_27896,N_27712);
nor U28043 (N_28043,N_27849,N_27760);
or U28044 (N_28044,N_27829,N_27742);
or U28045 (N_28045,N_27721,N_27887);
or U28046 (N_28046,N_27839,N_27757);
or U28047 (N_28047,N_27681,N_27786);
nand U28048 (N_28048,N_27878,N_27837);
xor U28049 (N_28049,N_27603,N_27811);
and U28050 (N_28050,N_27877,N_27788);
nand U28051 (N_28051,N_27649,N_27836);
and U28052 (N_28052,N_27678,N_27778);
or U28053 (N_28053,N_27712,N_27897);
nand U28054 (N_28054,N_27863,N_27810);
and U28055 (N_28055,N_27734,N_27613);
xor U28056 (N_28056,N_27603,N_27711);
nor U28057 (N_28057,N_27607,N_27894);
xor U28058 (N_28058,N_27812,N_27688);
xor U28059 (N_28059,N_27727,N_27741);
or U28060 (N_28060,N_27713,N_27785);
and U28061 (N_28061,N_27833,N_27646);
xnor U28062 (N_28062,N_27798,N_27852);
and U28063 (N_28063,N_27775,N_27836);
or U28064 (N_28064,N_27704,N_27846);
nor U28065 (N_28065,N_27802,N_27731);
nor U28066 (N_28066,N_27703,N_27686);
nand U28067 (N_28067,N_27842,N_27668);
and U28068 (N_28068,N_27687,N_27771);
or U28069 (N_28069,N_27685,N_27711);
nand U28070 (N_28070,N_27899,N_27739);
and U28071 (N_28071,N_27758,N_27767);
nor U28072 (N_28072,N_27619,N_27710);
or U28073 (N_28073,N_27690,N_27647);
or U28074 (N_28074,N_27742,N_27855);
xnor U28075 (N_28075,N_27707,N_27737);
xnor U28076 (N_28076,N_27833,N_27665);
nand U28077 (N_28077,N_27890,N_27824);
nor U28078 (N_28078,N_27739,N_27857);
or U28079 (N_28079,N_27776,N_27724);
and U28080 (N_28080,N_27646,N_27855);
or U28081 (N_28081,N_27890,N_27857);
nor U28082 (N_28082,N_27612,N_27680);
nor U28083 (N_28083,N_27861,N_27850);
nand U28084 (N_28084,N_27607,N_27850);
or U28085 (N_28085,N_27651,N_27670);
nand U28086 (N_28086,N_27814,N_27604);
nand U28087 (N_28087,N_27833,N_27880);
nor U28088 (N_28088,N_27677,N_27741);
or U28089 (N_28089,N_27623,N_27629);
nor U28090 (N_28090,N_27883,N_27833);
nand U28091 (N_28091,N_27851,N_27821);
and U28092 (N_28092,N_27896,N_27784);
nand U28093 (N_28093,N_27726,N_27696);
and U28094 (N_28094,N_27744,N_27854);
and U28095 (N_28095,N_27839,N_27744);
nand U28096 (N_28096,N_27608,N_27844);
nand U28097 (N_28097,N_27728,N_27653);
xor U28098 (N_28098,N_27747,N_27682);
nor U28099 (N_28099,N_27676,N_27687);
nand U28100 (N_28100,N_27892,N_27680);
nand U28101 (N_28101,N_27610,N_27636);
nor U28102 (N_28102,N_27840,N_27639);
nor U28103 (N_28103,N_27648,N_27784);
nor U28104 (N_28104,N_27680,N_27730);
or U28105 (N_28105,N_27784,N_27671);
and U28106 (N_28106,N_27892,N_27782);
nand U28107 (N_28107,N_27723,N_27897);
nor U28108 (N_28108,N_27683,N_27605);
nor U28109 (N_28109,N_27697,N_27870);
nand U28110 (N_28110,N_27800,N_27611);
nand U28111 (N_28111,N_27612,N_27859);
xor U28112 (N_28112,N_27762,N_27647);
xnor U28113 (N_28113,N_27717,N_27751);
and U28114 (N_28114,N_27824,N_27773);
nor U28115 (N_28115,N_27736,N_27742);
nand U28116 (N_28116,N_27870,N_27630);
and U28117 (N_28117,N_27764,N_27767);
nand U28118 (N_28118,N_27839,N_27852);
xnor U28119 (N_28119,N_27735,N_27768);
nand U28120 (N_28120,N_27654,N_27709);
nand U28121 (N_28121,N_27815,N_27759);
and U28122 (N_28122,N_27784,N_27787);
and U28123 (N_28123,N_27833,N_27826);
nand U28124 (N_28124,N_27711,N_27770);
xnor U28125 (N_28125,N_27652,N_27626);
or U28126 (N_28126,N_27829,N_27667);
xnor U28127 (N_28127,N_27803,N_27733);
or U28128 (N_28128,N_27668,N_27818);
or U28129 (N_28129,N_27630,N_27806);
nor U28130 (N_28130,N_27714,N_27752);
nor U28131 (N_28131,N_27886,N_27893);
nand U28132 (N_28132,N_27813,N_27619);
nand U28133 (N_28133,N_27888,N_27847);
xor U28134 (N_28134,N_27716,N_27604);
nor U28135 (N_28135,N_27622,N_27723);
xnor U28136 (N_28136,N_27775,N_27688);
or U28137 (N_28137,N_27697,N_27780);
and U28138 (N_28138,N_27747,N_27772);
nand U28139 (N_28139,N_27820,N_27866);
nor U28140 (N_28140,N_27863,N_27624);
nand U28141 (N_28141,N_27709,N_27767);
or U28142 (N_28142,N_27836,N_27675);
nand U28143 (N_28143,N_27774,N_27747);
nor U28144 (N_28144,N_27669,N_27896);
or U28145 (N_28145,N_27670,N_27687);
xor U28146 (N_28146,N_27713,N_27823);
and U28147 (N_28147,N_27861,N_27820);
nor U28148 (N_28148,N_27652,N_27651);
xnor U28149 (N_28149,N_27759,N_27653);
xor U28150 (N_28150,N_27803,N_27805);
nor U28151 (N_28151,N_27816,N_27743);
or U28152 (N_28152,N_27890,N_27859);
or U28153 (N_28153,N_27690,N_27685);
nand U28154 (N_28154,N_27858,N_27883);
or U28155 (N_28155,N_27733,N_27712);
nor U28156 (N_28156,N_27876,N_27638);
nor U28157 (N_28157,N_27650,N_27696);
nand U28158 (N_28158,N_27713,N_27645);
or U28159 (N_28159,N_27725,N_27648);
xor U28160 (N_28160,N_27697,N_27838);
nor U28161 (N_28161,N_27694,N_27742);
or U28162 (N_28162,N_27672,N_27824);
or U28163 (N_28163,N_27776,N_27681);
xnor U28164 (N_28164,N_27883,N_27621);
nor U28165 (N_28165,N_27838,N_27886);
nor U28166 (N_28166,N_27629,N_27604);
nor U28167 (N_28167,N_27870,N_27699);
nand U28168 (N_28168,N_27600,N_27737);
and U28169 (N_28169,N_27618,N_27634);
and U28170 (N_28170,N_27648,N_27828);
nand U28171 (N_28171,N_27821,N_27868);
nand U28172 (N_28172,N_27756,N_27735);
and U28173 (N_28173,N_27770,N_27715);
nor U28174 (N_28174,N_27680,N_27767);
nand U28175 (N_28175,N_27673,N_27669);
xor U28176 (N_28176,N_27899,N_27643);
or U28177 (N_28177,N_27637,N_27750);
xor U28178 (N_28178,N_27860,N_27660);
or U28179 (N_28179,N_27706,N_27654);
and U28180 (N_28180,N_27759,N_27770);
nor U28181 (N_28181,N_27841,N_27663);
and U28182 (N_28182,N_27644,N_27854);
nand U28183 (N_28183,N_27612,N_27630);
or U28184 (N_28184,N_27770,N_27725);
or U28185 (N_28185,N_27855,N_27834);
nand U28186 (N_28186,N_27828,N_27890);
nand U28187 (N_28187,N_27815,N_27760);
nor U28188 (N_28188,N_27706,N_27840);
xnor U28189 (N_28189,N_27742,N_27767);
and U28190 (N_28190,N_27761,N_27895);
or U28191 (N_28191,N_27722,N_27890);
and U28192 (N_28192,N_27664,N_27643);
or U28193 (N_28193,N_27804,N_27775);
nor U28194 (N_28194,N_27765,N_27669);
nor U28195 (N_28195,N_27668,N_27708);
xor U28196 (N_28196,N_27777,N_27807);
or U28197 (N_28197,N_27707,N_27640);
xnor U28198 (N_28198,N_27782,N_27870);
xor U28199 (N_28199,N_27677,N_27883);
and U28200 (N_28200,N_28053,N_28005);
and U28201 (N_28201,N_27988,N_28110);
and U28202 (N_28202,N_28082,N_28193);
xor U28203 (N_28203,N_28045,N_27942);
nand U28204 (N_28204,N_27901,N_27948);
xnor U28205 (N_28205,N_27992,N_28102);
nor U28206 (N_28206,N_28140,N_28065);
nor U28207 (N_28207,N_28018,N_27940);
xnor U28208 (N_28208,N_27977,N_28146);
xor U28209 (N_28209,N_28104,N_28052);
and U28210 (N_28210,N_28056,N_28194);
or U28211 (N_28211,N_28030,N_28109);
or U28212 (N_28212,N_28176,N_28111);
nand U28213 (N_28213,N_27989,N_28195);
nor U28214 (N_28214,N_28159,N_28192);
xor U28215 (N_28215,N_28148,N_27994);
or U28216 (N_28216,N_28118,N_27906);
nand U28217 (N_28217,N_27997,N_28137);
and U28218 (N_28218,N_28022,N_28171);
or U28219 (N_28219,N_27935,N_28113);
and U28220 (N_28220,N_28071,N_28187);
xor U28221 (N_28221,N_28138,N_28196);
and U28222 (N_28222,N_27952,N_28186);
or U28223 (N_28223,N_27941,N_28069);
xor U28224 (N_28224,N_28174,N_28024);
or U28225 (N_28225,N_28054,N_28150);
nand U28226 (N_28226,N_28042,N_28015);
xor U28227 (N_28227,N_28040,N_27937);
and U28228 (N_28228,N_27964,N_27965);
nor U28229 (N_28229,N_27953,N_28084);
xnor U28230 (N_28230,N_27971,N_28136);
and U28231 (N_28231,N_28037,N_27911);
nor U28232 (N_28232,N_28026,N_28097);
nor U28233 (N_28233,N_27922,N_27913);
and U28234 (N_28234,N_28068,N_28064);
or U28235 (N_28235,N_28107,N_28017);
xor U28236 (N_28236,N_28083,N_28087);
or U28237 (N_28237,N_27934,N_28181);
nor U28238 (N_28238,N_28155,N_27925);
xor U28239 (N_28239,N_28188,N_27960);
and U28240 (N_28240,N_28143,N_28038);
or U28241 (N_28241,N_28043,N_27954);
and U28242 (N_28242,N_28013,N_28066);
nor U28243 (N_28243,N_28145,N_28166);
or U28244 (N_28244,N_28185,N_28190);
nand U28245 (N_28245,N_27903,N_28078);
nand U28246 (N_28246,N_27938,N_28074);
nor U28247 (N_28247,N_28154,N_27978);
xnor U28248 (N_28248,N_27955,N_28180);
xnor U28249 (N_28249,N_27973,N_28009);
or U28250 (N_28250,N_28008,N_28020);
and U28251 (N_28251,N_27976,N_27924);
xor U28252 (N_28252,N_28129,N_27985);
nor U28253 (N_28253,N_27968,N_28121);
nand U28254 (N_28254,N_28012,N_27939);
xor U28255 (N_28255,N_27918,N_27957);
xnor U28256 (N_28256,N_28034,N_28168);
xor U28257 (N_28257,N_27987,N_28127);
nand U28258 (N_28258,N_28170,N_28101);
nand U28259 (N_28259,N_28095,N_28062);
nand U28260 (N_28260,N_28152,N_27975);
and U28261 (N_28261,N_27963,N_28161);
nand U28262 (N_28262,N_28019,N_27919);
and U28263 (N_28263,N_28163,N_28077);
nand U28264 (N_28264,N_27995,N_28060);
and U28265 (N_28265,N_28134,N_28105);
and U28266 (N_28266,N_27972,N_27980);
and U28267 (N_28267,N_28028,N_28093);
or U28268 (N_28268,N_27909,N_28177);
or U28269 (N_28269,N_28126,N_27930);
nor U28270 (N_28270,N_28139,N_28131);
xnor U28271 (N_28271,N_28162,N_27931);
and U28272 (N_28272,N_28094,N_28001);
or U28273 (N_28273,N_27917,N_27929);
nand U28274 (N_28274,N_28165,N_28156);
xnor U28275 (N_28275,N_28090,N_28179);
or U28276 (N_28276,N_28067,N_27932);
or U28277 (N_28277,N_28182,N_27990);
nor U28278 (N_28278,N_28080,N_28075);
xor U28279 (N_28279,N_28123,N_27993);
nor U28280 (N_28280,N_27970,N_28006);
xnor U28281 (N_28281,N_28175,N_28172);
xnor U28282 (N_28282,N_27951,N_28125);
nor U28283 (N_28283,N_27907,N_27967);
and U28284 (N_28284,N_28198,N_27986);
or U28285 (N_28285,N_28128,N_27928);
xor U28286 (N_28286,N_27984,N_28096);
nand U28287 (N_28287,N_27946,N_27902);
xnor U28288 (N_28288,N_27981,N_28112);
and U28289 (N_28289,N_28091,N_27949);
or U28290 (N_28290,N_28032,N_28157);
nor U28291 (N_28291,N_28092,N_28164);
and U28292 (N_28292,N_28100,N_28035);
nor U28293 (N_28293,N_28173,N_28189);
nor U28294 (N_28294,N_28011,N_27912);
nor U28295 (N_28295,N_28081,N_28036);
and U28296 (N_28296,N_28184,N_28191);
xnor U28297 (N_28297,N_28047,N_28041);
nand U28298 (N_28298,N_28167,N_28000);
nor U28299 (N_28299,N_28151,N_27910);
nand U28300 (N_28300,N_28070,N_28079);
xnor U28301 (N_28301,N_27974,N_28160);
xnor U28302 (N_28302,N_27936,N_28169);
or U28303 (N_28303,N_28120,N_27999);
and U28304 (N_28304,N_27983,N_28025);
nor U28305 (N_28305,N_28119,N_27933);
and U28306 (N_28306,N_28144,N_27943);
nand U28307 (N_28307,N_28049,N_27998);
and U28308 (N_28308,N_28147,N_28048);
nand U28309 (N_28309,N_27950,N_27904);
or U28310 (N_28310,N_28117,N_28057);
and U28311 (N_28311,N_28004,N_28051);
and U28312 (N_28312,N_28108,N_28197);
nand U28313 (N_28313,N_28103,N_28099);
xnor U28314 (N_28314,N_28058,N_28021);
nand U28315 (N_28315,N_27956,N_27969);
nor U28316 (N_28316,N_28158,N_28141);
xnor U28317 (N_28317,N_28088,N_28014);
and U28318 (N_28318,N_28089,N_28027);
and U28319 (N_28319,N_28063,N_28133);
nor U28320 (N_28320,N_28116,N_28016);
nand U28321 (N_28321,N_27982,N_27959);
nand U28322 (N_28322,N_27914,N_28031);
and U28323 (N_28323,N_27996,N_27920);
xnor U28324 (N_28324,N_28002,N_28073);
or U28325 (N_28325,N_28106,N_28124);
nor U28326 (N_28326,N_27900,N_28199);
nor U28327 (N_28327,N_27921,N_28023);
nor U28328 (N_28328,N_28003,N_28072);
or U28329 (N_28329,N_27927,N_27966);
xnor U28330 (N_28330,N_28033,N_27991);
and U28331 (N_28331,N_27947,N_27908);
nor U28332 (N_28332,N_28076,N_27944);
and U28333 (N_28333,N_27923,N_28149);
or U28334 (N_28334,N_28061,N_28130);
nand U28335 (N_28335,N_28050,N_27916);
xor U28336 (N_28336,N_28114,N_28059);
and U28337 (N_28337,N_28039,N_27958);
and U28338 (N_28338,N_27915,N_28183);
and U28339 (N_28339,N_28115,N_28135);
nand U28340 (N_28340,N_28178,N_27979);
nand U28341 (N_28341,N_28085,N_28055);
and U28342 (N_28342,N_28046,N_27926);
xor U28343 (N_28343,N_27945,N_28132);
or U28344 (N_28344,N_28007,N_27962);
xor U28345 (N_28345,N_28044,N_28010);
nand U28346 (N_28346,N_28029,N_27905);
nand U28347 (N_28347,N_28098,N_27961);
or U28348 (N_28348,N_28142,N_28086);
nor U28349 (N_28349,N_28122,N_28153);
or U28350 (N_28350,N_28191,N_28028);
nand U28351 (N_28351,N_28060,N_28079);
and U28352 (N_28352,N_28175,N_28017);
or U28353 (N_28353,N_28144,N_27959);
or U28354 (N_28354,N_27945,N_27932);
and U28355 (N_28355,N_28047,N_28158);
or U28356 (N_28356,N_28057,N_27966);
xor U28357 (N_28357,N_28039,N_28141);
nand U28358 (N_28358,N_28001,N_27905);
xor U28359 (N_28359,N_28165,N_28093);
nand U28360 (N_28360,N_28162,N_27925);
nor U28361 (N_28361,N_28002,N_28069);
or U28362 (N_28362,N_27901,N_27986);
or U28363 (N_28363,N_27961,N_28161);
or U28364 (N_28364,N_27950,N_27961);
xor U28365 (N_28365,N_28141,N_28033);
nand U28366 (N_28366,N_28146,N_28065);
xnor U28367 (N_28367,N_28179,N_27978);
xnor U28368 (N_28368,N_28001,N_27917);
nand U28369 (N_28369,N_28010,N_28170);
xor U28370 (N_28370,N_28146,N_28087);
nor U28371 (N_28371,N_27992,N_28067);
nor U28372 (N_28372,N_27921,N_28168);
xor U28373 (N_28373,N_27907,N_28182);
nor U28374 (N_28374,N_27996,N_27989);
nand U28375 (N_28375,N_28163,N_27951);
and U28376 (N_28376,N_28017,N_28102);
nor U28377 (N_28377,N_28066,N_28102);
nor U28378 (N_28378,N_28190,N_28038);
or U28379 (N_28379,N_27901,N_27903);
and U28380 (N_28380,N_28104,N_28057);
nor U28381 (N_28381,N_28125,N_28084);
and U28382 (N_28382,N_28088,N_27905);
or U28383 (N_28383,N_27951,N_27969);
nand U28384 (N_28384,N_28095,N_27932);
and U28385 (N_28385,N_27909,N_27977);
xnor U28386 (N_28386,N_28027,N_28028);
xor U28387 (N_28387,N_28134,N_28053);
nor U28388 (N_28388,N_28018,N_27995);
xnor U28389 (N_28389,N_28029,N_28149);
nor U28390 (N_28390,N_28033,N_28087);
nand U28391 (N_28391,N_28150,N_28021);
nand U28392 (N_28392,N_27987,N_27994);
xnor U28393 (N_28393,N_28026,N_27967);
nor U28394 (N_28394,N_27968,N_28173);
nor U28395 (N_28395,N_28177,N_28063);
and U28396 (N_28396,N_28016,N_28006);
nor U28397 (N_28397,N_28097,N_28041);
nand U28398 (N_28398,N_27976,N_28191);
or U28399 (N_28399,N_28141,N_27906);
or U28400 (N_28400,N_28100,N_28186);
nand U28401 (N_28401,N_28150,N_27918);
xor U28402 (N_28402,N_28014,N_27968);
nor U28403 (N_28403,N_27928,N_27978);
and U28404 (N_28404,N_28087,N_27924);
nor U28405 (N_28405,N_27996,N_27982);
xnor U28406 (N_28406,N_28050,N_28096);
and U28407 (N_28407,N_28068,N_27939);
xnor U28408 (N_28408,N_27995,N_28175);
or U28409 (N_28409,N_28184,N_28057);
or U28410 (N_28410,N_27927,N_28117);
nor U28411 (N_28411,N_27957,N_28152);
or U28412 (N_28412,N_28103,N_27941);
xnor U28413 (N_28413,N_27987,N_28199);
and U28414 (N_28414,N_27958,N_27960);
nor U28415 (N_28415,N_28028,N_28070);
nand U28416 (N_28416,N_28133,N_27953);
xor U28417 (N_28417,N_28018,N_27936);
xor U28418 (N_28418,N_28160,N_28066);
nand U28419 (N_28419,N_28089,N_28085);
and U28420 (N_28420,N_28042,N_28023);
and U28421 (N_28421,N_27988,N_28191);
or U28422 (N_28422,N_28181,N_28174);
and U28423 (N_28423,N_28074,N_28097);
nor U28424 (N_28424,N_28077,N_28127);
xnor U28425 (N_28425,N_27930,N_28004);
xor U28426 (N_28426,N_28021,N_28166);
xnor U28427 (N_28427,N_28069,N_28186);
and U28428 (N_28428,N_28005,N_28131);
nand U28429 (N_28429,N_27921,N_28118);
xnor U28430 (N_28430,N_28011,N_28176);
or U28431 (N_28431,N_28015,N_27983);
or U28432 (N_28432,N_28088,N_28022);
nor U28433 (N_28433,N_28055,N_28186);
and U28434 (N_28434,N_28191,N_27942);
nand U28435 (N_28435,N_28076,N_28169);
nand U28436 (N_28436,N_28077,N_28011);
xnor U28437 (N_28437,N_28117,N_28192);
nor U28438 (N_28438,N_27937,N_28019);
nand U28439 (N_28439,N_28175,N_27912);
nand U28440 (N_28440,N_27919,N_28080);
nand U28441 (N_28441,N_28141,N_28008);
xor U28442 (N_28442,N_28030,N_28140);
and U28443 (N_28443,N_27912,N_28012);
nand U28444 (N_28444,N_28138,N_27908);
or U28445 (N_28445,N_28141,N_28128);
nor U28446 (N_28446,N_28046,N_27934);
nor U28447 (N_28447,N_27960,N_28192);
nor U28448 (N_28448,N_28033,N_27965);
and U28449 (N_28449,N_28134,N_28153);
nor U28450 (N_28450,N_28122,N_27969);
nor U28451 (N_28451,N_28017,N_28182);
xor U28452 (N_28452,N_28132,N_28116);
and U28453 (N_28453,N_27912,N_28129);
nand U28454 (N_28454,N_27941,N_27916);
nor U28455 (N_28455,N_27902,N_28165);
nor U28456 (N_28456,N_28079,N_28184);
or U28457 (N_28457,N_28033,N_28020);
nor U28458 (N_28458,N_27908,N_27915);
nor U28459 (N_28459,N_28198,N_28025);
xnor U28460 (N_28460,N_28182,N_28077);
and U28461 (N_28461,N_27926,N_27971);
and U28462 (N_28462,N_27951,N_27924);
and U28463 (N_28463,N_28146,N_28013);
nor U28464 (N_28464,N_28134,N_28106);
nor U28465 (N_28465,N_27953,N_27989);
nor U28466 (N_28466,N_27994,N_28190);
or U28467 (N_28467,N_27989,N_27914);
nand U28468 (N_28468,N_28125,N_27986);
nor U28469 (N_28469,N_27977,N_28075);
and U28470 (N_28470,N_28081,N_28048);
nand U28471 (N_28471,N_28064,N_28037);
nor U28472 (N_28472,N_27901,N_28155);
or U28473 (N_28473,N_28143,N_27957);
and U28474 (N_28474,N_28185,N_27928);
nand U28475 (N_28475,N_27970,N_28016);
xor U28476 (N_28476,N_27993,N_28153);
and U28477 (N_28477,N_28039,N_28144);
nor U28478 (N_28478,N_28091,N_27979);
nor U28479 (N_28479,N_28011,N_27906);
and U28480 (N_28480,N_28166,N_28006);
nor U28481 (N_28481,N_28159,N_27927);
xnor U28482 (N_28482,N_28135,N_28194);
or U28483 (N_28483,N_27964,N_28159);
xnor U28484 (N_28484,N_27958,N_28063);
or U28485 (N_28485,N_28133,N_28174);
nor U28486 (N_28486,N_27941,N_28165);
nand U28487 (N_28487,N_28192,N_28098);
and U28488 (N_28488,N_28115,N_27980);
xor U28489 (N_28489,N_27925,N_27982);
nor U28490 (N_28490,N_27979,N_27994);
nor U28491 (N_28491,N_27905,N_28058);
nor U28492 (N_28492,N_27945,N_28002);
and U28493 (N_28493,N_28186,N_28119);
or U28494 (N_28494,N_27918,N_28087);
nand U28495 (N_28495,N_28007,N_28105);
xor U28496 (N_28496,N_28054,N_28132);
nor U28497 (N_28497,N_28105,N_28015);
and U28498 (N_28498,N_27942,N_27914);
xor U28499 (N_28499,N_27977,N_27956);
nor U28500 (N_28500,N_28252,N_28202);
or U28501 (N_28501,N_28369,N_28456);
and U28502 (N_28502,N_28238,N_28404);
nor U28503 (N_28503,N_28342,N_28338);
nand U28504 (N_28504,N_28418,N_28372);
xor U28505 (N_28505,N_28472,N_28486);
nor U28506 (N_28506,N_28260,N_28207);
nor U28507 (N_28507,N_28233,N_28267);
xor U28508 (N_28508,N_28208,N_28414);
nor U28509 (N_28509,N_28446,N_28229);
xnor U28510 (N_28510,N_28381,N_28245);
nand U28511 (N_28511,N_28359,N_28259);
nor U28512 (N_28512,N_28353,N_28395);
nor U28513 (N_28513,N_28203,N_28264);
or U28514 (N_28514,N_28438,N_28488);
and U28515 (N_28515,N_28223,N_28276);
nand U28516 (N_28516,N_28289,N_28326);
or U28517 (N_28517,N_28331,N_28282);
nor U28518 (N_28518,N_28370,N_28483);
and U28519 (N_28519,N_28253,N_28270);
xor U28520 (N_28520,N_28447,N_28215);
nand U28521 (N_28521,N_28397,N_28349);
nor U28522 (N_28522,N_28330,N_28336);
xor U28523 (N_28523,N_28487,N_28494);
and U28524 (N_28524,N_28413,N_28367);
and U28525 (N_28525,N_28379,N_28204);
and U28526 (N_28526,N_28281,N_28346);
xor U28527 (N_28527,N_28429,N_28375);
nand U28528 (N_28528,N_28307,N_28268);
and U28529 (N_28529,N_28317,N_28380);
and U28530 (N_28530,N_28244,N_28328);
nand U28531 (N_28531,N_28366,N_28293);
nand U28532 (N_28532,N_28363,N_28439);
nor U28533 (N_28533,N_28361,N_28319);
or U28534 (N_28534,N_28257,N_28237);
or U28535 (N_28535,N_28426,N_28347);
and U28536 (N_28536,N_28405,N_28206);
nand U28537 (N_28537,N_28345,N_28462);
nand U28538 (N_28538,N_28211,N_28256);
or U28539 (N_28539,N_28396,N_28312);
xnor U28540 (N_28540,N_28417,N_28216);
or U28541 (N_28541,N_28287,N_28271);
or U28542 (N_28542,N_28444,N_28273);
nand U28543 (N_28543,N_28454,N_28355);
xnor U28544 (N_28544,N_28239,N_28209);
nand U28545 (N_28545,N_28343,N_28220);
xnor U28546 (N_28546,N_28224,N_28234);
xnor U28547 (N_28547,N_28467,N_28392);
nand U28548 (N_28548,N_28315,N_28272);
xor U28549 (N_28549,N_28228,N_28371);
nor U28550 (N_28550,N_28340,N_28477);
nor U28551 (N_28551,N_28401,N_28306);
nor U28552 (N_28552,N_28358,N_28246);
nand U28553 (N_28553,N_28263,N_28296);
xnor U28554 (N_28554,N_28301,N_28368);
and U28555 (N_28555,N_28266,N_28427);
and U28556 (N_28556,N_28407,N_28230);
nor U28557 (N_28557,N_28305,N_28471);
nand U28558 (N_28558,N_28295,N_28378);
or U28559 (N_28559,N_28441,N_28416);
or U28560 (N_28560,N_28394,N_28286);
nand U28561 (N_28561,N_28351,N_28464);
and U28562 (N_28562,N_28218,N_28313);
or U28563 (N_28563,N_28242,N_28217);
nand U28564 (N_28564,N_28299,N_28411);
nor U28565 (N_28565,N_28236,N_28344);
nand U28566 (N_28566,N_28466,N_28469);
or U28567 (N_28567,N_28304,N_28448);
and U28568 (N_28568,N_28322,N_28249);
or U28569 (N_28569,N_28430,N_28275);
nand U28570 (N_28570,N_28484,N_28360);
nor U28571 (N_28571,N_28357,N_28421);
nor U28572 (N_28572,N_28415,N_28496);
or U28573 (N_28573,N_28300,N_28490);
or U28574 (N_28574,N_28258,N_28442);
and U28575 (N_28575,N_28474,N_28470);
nand U28576 (N_28576,N_28314,N_28356);
xnor U28577 (N_28577,N_28241,N_28443);
xor U28578 (N_28578,N_28440,N_28388);
nor U28579 (N_28579,N_28374,N_28376);
or U28580 (N_28580,N_28311,N_28316);
nor U28581 (N_28581,N_28422,N_28320);
or U28582 (N_28582,N_28458,N_28384);
nand U28583 (N_28583,N_28221,N_28433);
nor U28584 (N_28584,N_28386,N_28200);
xor U28585 (N_28585,N_28262,N_28310);
nand U28586 (N_28586,N_28460,N_28334);
nor U28587 (N_28587,N_28461,N_28225);
nor U28588 (N_28588,N_28398,N_28435);
nor U28589 (N_28589,N_28214,N_28465);
xnor U28590 (N_28590,N_28261,N_28247);
or U28591 (N_28591,N_28431,N_28291);
nand U28592 (N_28592,N_28231,N_28478);
nand U28593 (N_28593,N_28391,N_28309);
and U28594 (N_28594,N_28341,N_28450);
xor U28595 (N_28595,N_28277,N_28284);
nor U28596 (N_28596,N_28445,N_28455);
nand U28597 (N_28597,N_28333,N_28325);
xor U28598 (N_28598,N_28213,N_28428);
xor U28599 (N_28599,N_28329,N_28393);
or U28600 (N_28600,N_28480,N_28205);
xor U28601 (N_28601,N_28294,N_28406);
xnor U28602 (N_28602,N_28482,N_28499);
nor U28603 (N_28603,N_28292,N_28308);
xnor U28604 (N_28604,N_28389,N_28385);
xor U28605 (N_28605,N_28243,N_28279);
nor U28606 (N_28606,N_28492,N_28403);
xor U28607 (N_28607,N_28410,N_28491);
xnor U28608 (N_28608,N_28409,N_28400);
xnor U28609 (N_28609,N_28383,N_28201);
and U28610 (N_28610,N_28475,N_28339);
nand U28611 (N_28611,N_28265,N_28377);
and U28612 (N_28612,N_28352,N_28297);
nand U28613 (N_28613,N_28479,N_28354);
and U28614 (N_28614,N_28432,N_28250);
nor U28615 (N_28615,N_28451,N_28278);
and U28616 (N_28616,N_28495,N_28365);
nor U28617 (N_28617,N_28280,N_28423);
and U28618 (N_28618,N_28473,N_28248);
nand U28619 (N_28619,N_28408,N_28219);
xnor U28620 (N_28620,N_28390,N_28332);
and U28621 (N_28621,N_28235,N_28274);
xnor U28622 (N_28622,N_28459,N_28437);
nor U28623 (N_28623,N_28348,N_28399);
or U28624 (N_28624,N_28425,N_28476);
and U28625 (N_28625,N_28255,N_28303);
nor U28626 (N_28626,N_28285,N_28489);
xor U28627 (N_28627,N_28321,N_28387);
and U28628 (N_28628,N_28468,N_28226);
or U28629 (N_28629,N_28222,N_28449);
and U28630 (N_28630,N_28323,N_28498);
or U28631 (N_28631,N_28335,N_28485);
nand U28632 (N_28632,N_28298,N_28463);
or U28633 (N_28633,N_28457,N_28493);
or U28634 (N_28634,N_28452,N_28327);
xor U28635 (N_28635,N_28302,N_28337);
or U28636 (N_28636,N_28210,N_28290);
xnor U28637 (N_28637,N_28350,N_28424);
and U28638 (N_28638,N_28382,N_28453);
and U28639 (N_28639,N_28254,N_28434);
xor U28640 (N_28640,N_28227,N_28419);
and U28641 (N_28641,N_28251,N_28402);
nor U28642 (N_28642,N_28318,N_28373);
or U28643 (N_28643,N_28269,N_28212);
and U28644 (N_28644,N_28232,N_28324);
nor U28645 (N_28645,N_28497,N_28283);
nand U28646 (N_28646,N_28420,N_28412);
and U28647 (N_28647,N_28288,N_28481);
and U28648 (N_28648,N_28240,N_28362);
nand U28649 (N_28649,N_28436,N_28364);
nor U28650 (N_28650,N_28285,N_28270);
nor U28651 (N_28651,N_28264,N_28339);
nor U28652 (N_28652,N_28403,N_28226);
nor U28653 (N_28653,N_28376,N_28457);
and U28654 (N_28654,N_28247,N_28307);
and U28655 (N_28655,N_28309,N_28403);
or U28656 (N_28656,N_28286,N_28360);
and U28657 (N_28657,N_28349,N_28347);
nor U28658 (N_28658,N_28338,N_28418);
nand U28659 (N_28659,N_28295,N_28466);
nor U28660 (N_28660,N_28217,N_28473);
nor U28661 (N_28661,N_28391,N_28300);
nor U28662 (N_28662,N_28272,N_28427);
nand U28663 (N_28663,N_28488,N_28274);
or U28664 (N_28664,N_28351,N_28324);
nand U28665 (N_28665,N_28265,N_28275);
nand U28666 (N_28666,N_28363,N_28488);
xor U28667 (N_28667,N_28251,N_28387);
and U28668 (N_28668,N_28202,N_28359);
xnor U28669 (N_28669,N_28479,N_28332);
nand U28670 (N_28670,N_28307,N_28478);
or U28671 (N_28671,N_28243,N_28443);
and U28672 (N_28672,N_28488,N_28427);
nor U28673 (N_28673,N_28335,N_28297);
nor U28674 (N_28674,N_28227,N_28243);
and U28675 (N_28675,N_28206,N_28278);
nor U28676 (N_28676,N_28495,N_28490);
nand U28677 (N_28677,N_28313,N_28401);
nor U28678 (N_28678,N_28245,N_28293);
or U28679 (N_28679,N_28421,N_28271);
xnor U28680 (N_28680,N_28375,N_28300);
nor U28681 (N_28681,N_28212,N_28395);
or U28682 (N_28682,N_28286,N_28287);
nand U28683 (N_28683,N_28290,N_28273);
nand U28684 (N_28684,N_28470,N_28386);
nand U28685 (N_28685,N_28477,N_28439);
or U28686 (N_28686,N_28445,N_28300);
nor U28687 (N_28687,N_28407,N_28221);
nor U28688 (N_28688,N_28484,N_28348);
nor U28689 (N_28689,N_28311,N_28309);
nand U28690 (N_28690,N_28472,N_28251);
nor U28691 (N_28691,N_28259,N_28257);
xor U28692 (N_28692,N_28433,N_28400);
and U28693 (N_28693,N_28349,N_28318);
or U28694 (N_28694,N_28371,N_28277);
or U28695 (N_28695,N_28484,N_28415);
or U28696 (N_28696,N_28435,N_28369);
or U28697 (N_28697,N_28250,N_28321);
and U28698 (N_28698,N_28308,N_28499);
xor U28699 (N_28699,N_28393,N_28234);
and U28700 (N_28700,N_28315,N_28209);
xnor U28701 (N_28701,N_28362,N_28222);
nor U28702 (N_28702,N_28467,N_28378);
nor U28703 (N_28703,N_28391,N_28372);
or U28704 (N_28704,N_28323,N_28385);
nand U28705 (N_28705,N_28321,N_28307);
or U28706 (N_28706,N_28243,N_28238);
and U28707 (N_28707,N_28285,N_28279);
nor U28708 (N_28708,N_28245,N_28489);
xor U28709 (N_28709,N_28242,N_28392);
nand U28710 (N_28710,N_28349,N_28345);
xor U28711 (N_28711,N_28274,N_28230);
or U28712 (N_28712,N_28475,N_28266);
nor U28713 (N_28713,N_28429,N_28388);
nand U28714 (N_28714,N_28340,N_28303);
xor U28715 (N_28715,N_28356,N_28413);
or U28716 (N_28716,N_28426,N_28406);
and U28717 (N_28717,N_28405,N_28319);
nor U28718 (N_28718,N_28235,N_28397);
xor U28719 (N_28719,N_28283,N_28437);
xnor U28720 (N_28720,N_28440,N_28399);
xnor U28721 (N_28721,N_28348,N_28450);
xor U28722 (N_28722,N_28343,N_28297);
nand U28723 (N_28723,N_28361,N_28347);
and U28724 (N_28724,N_28387,N_28373);
nand U28725 (N_28725,N_28497,N_28437);
nand U28726 (N_28726,N_28435,N_28475);
nand U28727 (N_28727,N_28278,N_28473);
or U28728 (N_28728,N_28218,N_28293);
nor U28729 (N_28729,N_28407,N_28282);
and U28730 (N_28730,N_28332,N_28240);
and U28731 (N_28731,N_28363,N_28461);
and U28732 (N_28732,N_28280,N_28442);
and U28733 (N_28733,N_28322,N_28247);
or U28734 (N_28734,N_28204,N_28375);
nor U28735 (N_28735,N_28270,N_28353);
or U28736 (N_28736,N_28226,N_28495);
xnor U28737 (N_28737,N_28498,N_28465);
nor U28738 (N_28738,N_28389,N_28228);
and U28739 (N_28739,N_28303,N_28230);
or U28740 (N_28740,N_28486,N_28488);
xor U28741 (N_28741,N_28232,N_28416);
xor U28742 (N_28742,N_28347,N_28449);
nand U28743 (N_28743,N_28382,N_28323);
and U28744 (N_28744,N_28203,N_28224);
and U28745 (N_28745,N_28247,N_28440);
or U28746 (N_28746,N_28359,N_28341);
nand U28747 (N_28747,N_28229,N_28204);
and U28748 (N_28748,N_28229,N_28487);
or U28749 (N_28749,N_28446,N_28230);
and U28750 (N_28750,N_28477,N_28440);
nor U28751 (N_28751,N_28254,N_28362);
or U28752 (N_28752,N_28255,N_28482);
and U28753 (N_28753,N_28220,N_28491);
and U28754 (N_28754,N_28373,N_28362);
or U28755 (N_28755,N_28261,N_28346);
or U28756 (N_28756,N_28464,N_28250);
xnor U28757 (N_28757,N_28473,N_28390);
and U28758 (N_28758,N_28232,N_28225);
or U28759 (N_28759,N_28489,N_28288);
nor U28760 (N_28760,N_28464,N_28385);
or U28761 (N_28761,N_28337,N_28303);
xnor U28762 (N_28762,N_28303,N_28247);
and U28763 (N_28763,N_28449,N_28490);
xor U28764 (N_28764,N_28392,N_28415);
nor U28765 (N_28765,N_28236,N_28224);
nor U28766 (N_28766,N_28310,N_28370);
nor U28767 (N_28767,N_28380,N_28298);
nor U28768 (N_28768,N_28361,N_28341);
nor U28769 (N_28769,N_28361,N_28464);
nor U28770 (N_28770,N_28210,N_28266);
or U28771 (N_28771,N_28332,N_28361);
xnor U28772 (N_28772,N_28325,N_28355);
xnor U28773 (N_28773,N_28228,N_28343);
or U28774 (N_28774,N_28497,N_28343);
xor U28775 (N_28775,N_28290,N_28307);
nand U28776 (N_28776,N_28357,N_28441);
xnor U28777 (N_28777,N_28362,N_28425);
and U28778 (N_28778,N_28207,N_28238);
or U28779 (N_28779,N_28315,N_28418);
xnor U28780 (N_28780,N_28327,N_28283);
nor U28781 (N_28781,N_28310,N_28392);
nor U28782 (N_28782,N_28228,N_28200);
and U28783 (N_28783,N_28425,N_28248);
and U28784 (N_28784,N_28480,N_28374);
or U28785 (N_28785,N_28328,N_28269);
and U28786 (N_28786,N_28429,N_28450);
or U28787 (N_28787,N_28377,N_28324);
nand U28788 (N_28788,N_28360,N_28410);
nor U28789 (N_28789,N_28331,N_28302);
xor U28790 (N_28790,N_28359,N_28323);
nand U28791 (N_28791,N_28376,N_28332);
xor U28792 (N_28792,N_28394,N_28353);
nand U28793 (N_28793,N_28459,N_28280);
nor U28794 (N_28794,N_28429,N_28374);
and U28795 (N_28795,N_28497,N_28262);
or U28796 (N_28796,N_28207,N_28476);
nand U28797 (N_28797,N_28274,N_28396);
nor U28798 (N_28798,N_28250,N_28496);
or U28799 (N_28799,N_28474,N_28453);
or U28800 (N_28800,N_28621,N_28706);
or U28801 (N_28801,N_28632,N_28528);
or U28802 (N_28802,N_28591,N_28618);
xnor U28803 (N_28803,N_28743,N_28588);
nand U28804 (N_28804,N_28711,N_28513);
xnor U28805 (N_28805,N_28788,N_28782);
nand U28806 (N_28806,N_28716,N_28504);
or U28807 (N_28807,N_28762,N_28587);
xor U28808 (N_28808,N_28645,N_28786);
and U28809 (N_28809,N_28506,N_28568);
xnor U28810 (N_28810,N_28644,N_28685);
or U28811 (N_28811,N_28530,N_28671);
and U28812 (N_28812,N_28534,N_28581);
nand U28813 (N_28813,N_28783,N_28520);
xnor U28814 (N_28814,N_28656,N_28714);
nand U28815 (N_28815,N_28700,N_28597);
or U28816 (N_28816,N_28546,N_28741);
nor U28817 (N_28817,N_28677,N_28503);
or U28818 (N_28818,N_28763,N_28695);
and U28819 (N_28819,N_28787,N_28679);
and U28820 (N_28820,N_28509,N_28767);
or U28821 (N_28821,N_28682,N_28798);
nor U28822 (N_28822,N_28712,N_28605);
xnor U28823 (N_28823,N_28675,N_28773);
nor U28824 (N_28824,N_28694,N_28598);
nor U28825 (N_28825,N_28541,N_28556);
nor U28826 (N_28826,N_28500,N_28639);
or U28827 (N_28827,N_28608,N_28780);
nand U28828 (N_28828,N_28594,N_28617);
nor U28829 (N_28829,N_28660,N_28651);
xor U28830 (N_28830,N_28547,N_28703);
and U28831 (N_28831,N_28582,N_28557);
nor U28832 (N_28832,N_28699,N_28579);
nor U28833 (N_28833,N_28570,N_28544);
or U28834 (N_28834,N_28664,N_28553);
nor U28835 (N_28835,N_28658,N_28585);
nor U28836 (N_28836,N_28702,N_28567);
or U28837 (N_28837,N_28564,N_28672);
nand U28838 (N_28838,N_28736,N_28758);
or U28839 (N_28839,N_28789,N_28665);
and U28840 (N_28840,N_28540,N_28596);
nor U28841 (N_28841,N_28777,N_28583);
nand U28842 (N_28842,N_28640,N_28749);
nand U28843 (N_28843,N_28523,N_28512);
and U28844 (N_28844,N_28641,N_28769);
and U28845 (N_28845,N_28717,N_28770);
nand U28846 (N_28846,N_28721,N_28696);
xnor U28847 (N_28847,N_28593,N_28750);
and U28848 (N_28848,N_28792,N_28794);
xnor U28849 (N_28849,N_28552,N_28747);
xor U28850 (N_28850,N_28616,N_28562);
and U28851 (N_28851,N_28728,N_28771);
nand U28852 (N_28852,N_28681,N_28701);
nor U28853 (N_28853,N_28555,N_28559);
xnor U28854 (N_28854,N_28691,N_28521);
or U28855 (N_28855,N_28793,N_28514);
nor U28856 (N_28856,N_28536,N_28727);
or U28857 (N_28857,N_28768,N_28775);
xnor U28858 (N_28858,N_28537,N_28667);
and U28859 (N_28859,N_28538,N_28609);
or U28860 (N_28860,N_28502,N_28508);
xor U28861 (N_28861,N_28524,N_28759);
or U28862 (N_28862,N_28566,N_28554);
or U28863 (N_28863,N_28629,N_28614);
xnor U28864 (N_28864,N_28766,N_28799);
xor U28865 (N_28865,N_28525,N_28668);
xnor U28866 (N_28866,N_28688,N_28673);
nand U28867 (N_28867,N_28742,N_28753);
xnor U28868 (N_28868,N_28560,N_28636);
xor U28869 (N_28869,N_28589,N_28516);
xnor U28870 (N_28870,N_28657,N_28628);
nor U28871 (N_28871,N_28539,N_28752);
nor U28872 (N_28872,N_28655,N_28731);
and U28873 (N_28873,N_28765,N_28590);
nand U28874 (N_28874,N_28738,N_28666);
xnor U28875 (N_28875,N_28595,N_28613);
xor U28876 (N_28876,N_28648,N_28517);
nor U28877 (N_28877,N_28729,N_28757);
nand U28878 (N_28878,N_28630,N_28584);
or U28879 (N_28879,N_28569,N_28518);
nor U28880 (N_28880,N_28548,N_28779);
or U28881 (N_28881,N_28744,N_28710);
nor U28882 (N_28882,N_28659,N_28748);
or U28883 (N_28883,N_28684,N_28674);
and U28884 (N_28884,N_28784,N_28708);
nand U28885 (N_28885,N_28693,N_28563);
and U28886 (N_28886,N_28545,N_28620);
xor U28887 (N_28887,N_28592,N_28663);
and U28888 (N_28888,N_28737,N_28709);
xor U28889 (N_28889,N_28637,N_28602);
xor U28890 (N_28890,N_28732,N_28760);
or U28891 (N_28891,N_28735,N_28661);
or U28892 (N_28892,N_28785,N_28781);
or U28893 (N_28893,N_28611,N_28751);
nor U28894 (N_28894,N_28776,N_28724);
nor U28895 (N_28895,N_28612,N_28649);
nor U28896 (N_28896,N_28745,N_28622);
nand U28897 (N_28897,N_28796,N_28551);
nor U28898 (N_28898,N_28669,N_28680);
nor U28899 (N_28899,N_28572,N_28795);
or U28900 (N_28900,N_28670,N_28533);
or U28901 (N_28901,N_28761,N_28526);
and U28902 (N_28902,N_28604,N_28790);
xor U28903 (N_28903,N_28576,N_28739);
or U28904 (N_28904,N_28558,N_28654);
and U28905 (N_28905,N_28723,N_28606);
nand U28906 (N_28906,N_28650,N_28719);
and U28907 (N_28907,N_28686,N_28510);
and U28908 (N_28908,N_28690,N_28643);
xnor U28909 (N_28909,N_28549,N_28726);
or U28910 (N_28910,N_28543,N_28638);
and U28911 (N_28911,N_28565,N_28627);
and U28912 (N_28912,N_28624,N_28619);
or U28913 (N_28913,N_28519,N_28507);
nand U28914 (N_28914,N_28704,N_28764);
or U28915 (N_28915,N_28687,N_28720);
xor U28916 (N_28916,N_28522,N_28615);
or U28917 (N_28917,N_28715,N_28550);
nand U28918 (N_28918,N_28631,N_28600);
and U28919 (N_28919,N_28705,N_28573);
nor U28920 (N_28920,N_28683,N_28713);
nor U28921 (N_28921,N_28652,N_28734);
xnor U28922 (N_28922,N_28754,N_28722);
xor U28923 (N_28923,N_28692,N_28746);
nor U28924 (N_28924,N_28797,N_28625);
or U28925 (N_28925,N_28603,N_28542);
nor U28926 (N_28926,N_28689,N_28697);
nand U28927 (N_28927,N_28755,N_28791);
and U28928 (N_28928,N_28634,N_28561);
and U28929 (N_28929,N_28535,N_28707);
xor U28930 (N_28930,N_28756,N_28642);
nor U28931 (N_28931,N_28733,N_28653);
and U28932 (N_28932,N_28740,N_28662);
nor U28933 (N_28933,N_28646,N_28599);
or U28934 (N_28934,N_28623,N_28778);
nand U28935 (N_28935,N_28580,N_28571);
xnor U28936 (N_28936,N_28718,N_28575);
nand U28937 (N_28937,N_28698,N_28505);
and U28938 (N_28938,N_28676,N_28501);
or U28939 (N_28939,N_28529,N_28678);
nor U28940 (N_28940,N_28601,N_28577);
nor U28941 (N_28941,N_28515,N_28610);
nor U28942 (N_28942,N_28531,N_28527);
and U28943 (N_28943,N_28730,N_28511);
xor U28944 (N_28944,N_28574,N_28635);
and U28945 (N_28945,N_28633,N_28774);
or U28946 (N_28946,N_28626,N_28725);
nor U28947 (N_28947,N_28586,N_28607);
or U28948 (N_28948,N_28578,N_28647);
xnor U28949 (N_28949,N_28532,N_28772);
or U28950 (N_28950,N_28609,N_28558);
xor U28951 (N_28951,N_28773,N_28732);
nand U28952 (N_28952,N_28551,N_28578);
xnor U28953 (N_28953,N_28681,N_28664);
xor U28954 (N_28954,N_28761,N_28672);
nor U28955 (N_28955,N_28789,N_28785);
nand U28956 (N_28956,N_28627,N_28548);
or U28957 (N_28957,N_28771,N_28745);
nor U28958 (N_28958,N_28668,N_28664);
or U28959 (N_28959,N_28755,N_28785);
nand U28960 (N_28960,N_28763,N_28504);
and U28961 (N_28961,N_28684,N_28622);
nor U28962 (N_28962,N_28623,N_28688);
and U28963 (N_28963,N_28645,N_28642);
nor U28964 (N_28964,N_28640,N_28723);
nand U28965 (N_28965,N_28648,N_28702);
nand U28966 (N_28966,N_28731,N_28591);
nand U28967 (N_28967,N_28501,N_28649);
and U28968 (N_28968,N_28651,N_28799);
and U28969 (N_28969,N_28713,N_28502);
and U28970 (N_28970,N_28679,N_28550);
and U28971 (N_28971,N_28594,N_28688);
xor U28972 (N_28972,N_28793,N_28682);
nand U28973 (N_28973,N_28642,N_28709);
and U28974 (N_28974,N_28566,N_28535);
xor U28975 (N_28975,N_28563,N_28598);
nand U28976 (N_28976,N_28751,N_28709);
nor U28977 (N_28977,N_28721,N_28523);
nand U28978 (N_28978,N_28583,N_28621);
xor U28979 (N_28979,N_28504,N_28721);
or U28980 (N_28980,N_28655,N_28782);
and U28981 (N_28981,N_28603,N_28595);
xor U28982 (N_28982,N_28549,N_28509);
or U28983 (N_28983,N_28749,N_28535);
nand U28984 (N_28984,N_28792,N_28578);
nor U28985 (N_28985,N_28663,N_28797);
nand U28986 (N_28986,N_28693,N_28660);
and U28987 (N_28987,N_28638,N_28636);
xnor U28988 (N_28988,N_28744,N_28501);
and U28989 (N_28989,N_28595,N_28776);
and U28990 (N_28990,N_28500,N_28593);
and U28991 (N_28991,N_28747,N_28521);
nand U28992 (N_28992,N_28642,N_28542);
or U28993 (N_28993,N_28761,N_28762);
xnor U28994 (N_28994,N_28656,N_28528);
nor U28995 (N_28995,N_28634,N_28511);
and U28996 (N_28996,N_28592,N_28526);
or U28997 (N_28997,N_28713,N_28613);
nor U28998 (N_28998,N_28656,N_28742);
and U28999 (N_28999,N_28745,N_28743);
xnor U29000 (N_29000,N_28685,N_28724);
nand U29001 (N_29001,N_28707,N_28748);
and U29002 (N_29002,N_28606,N_28638);
nor U29003 (N_29003,N_28793,N_28708);
nor U29004 (N_29004,N_28629,N_28611);
and U29005 (N_29005,N_28723,N_28761);
or U29006 (N_29006,N_28684,N_28757);
xor U29007 (N_29007,N_28522,N_28655);
nor U29008 (N_29008,N_28751,N_28503);
and U29009 (N_29009,N_28544,N_28629);
nor U29010 (N_29010,N_28600,N_28721);
nand U29011 (N_29011,N_28563,N_28793);
and U29012 (N_29012,N_28571,N_28676);
nor U29013 (N_29013,N_28722,N_28737);
and U29014 (N_29014,N_28673,N_28501);
or U29015 (N_29015,N_28569,N_28588);
xor U29016 (N_29016,N_28731,N_28626);
nand U29017 (N_29017,N_28605,N_28798);
or U29018 (N_29018,N_28561,N_28748);
nand U29019 (N_29019,N_28769,N_28602);
nand U29020 (N_29020,N_28741,N_28780);
nor U29021 (N_29021,N_28528,N_28653);
nand U29022 (N_29022,N_28657,N_28716);
xnor U29023 (N_29023,N_28509,N_28727);
or U29024 (N_29024,N_28651,N_28574);
and U29025 (N_29025,N_28718,N_28710);
nor U29026 (N_29026,N_28684,N_28784);
nor U29027 (N_29027,N_28770,N_28617);
or U29028 (N_29028,N_28739,N_28668);
nor U29029 (N_29029,N_28776,N_28530);
nor U29030 (N_29030,N_28517,N_28676);
or U29031 (N_29031,N_28611,N_28673);
xor U29032 (N_29032,N_28643,N_28688);
and U29033 (N_29033,N_28539,N_28733);
and U29034 (N_29034,N_28658,N_28616);
and U29035 (N_29035,N_28658,N_28737);
nand U29036 (N_29036,N_28566,N_28514);
nor U29037 (N_29037,N_28537,N_28768);
nand U29038 (N_29038,N_28578,N_28608);
or U29039 (N_29039,N_28729,N_28701);
xor U29040 (N_29040,N_28790,N_28775);
nand U29041 (N_29041,N_28564,N_28798);
and U29042 (N_29042,N_28547,N_28530);
or U29043 (N_29043,N_28649,N_28506);
nor U29044 (N_29044,N_28757,N_28623);
nor U29045 (N_29045,N_28554,N_28782);
xor U29046 (N_29046,N_28637,N_28644);
nand U29047 (N_29047,N_28583,N_28732);
xnor U29048 (N_29048,N_28786,N_28696);
xor U29049 (N_29049,N_28610,N_28780);
xor U29050 (N_29050,N_28766,N_28687);
nand U29051 (N_29051,N_28633,N_28707);
nand U29052 (N_29052,N_28647,N_28777);
and U29053 (N_29053,N_28702,N_28667);
nand U29054 (N_29054,N_28508,N_28570);
xor U29055 (N_29055,N_28746,N_28577);
nor U29056 (N_29056,N_28580,N_28550);
or U29057 (N_29057,N_28545,N_28716);
or U29058 (N_29058,N_28643,N_28732);
and U29059 (N_29059,N_28628,N_28608);
nand U29060 (N_29060,N_28634,N_28643);
nand U29061 (N_29061,N_28691,N_28622);
or U29062 (N_29062,N_28790,N_28503);
nor U29063 (N_29063,N_28577,N_28618);
xnor U29064 (N_29064,N_28752,N_28674);
xnor U29065 (N_29065,N_28547,N_28740);
xor U29066 (N_29066,N_28799,N_28775);
and U29067 (N_29067,N_28716,N_28783);
or U29068 (N_29068,N_28617,N_28539);
nand U29069 (N_29069,N_28767,N_28677);
nand U29070 (N_29070,N_28692,N_28794);
nand U29071 (N_29071,N_28605,N_28643);
xnor U29072 (N_29072,N_28668,N_28693);
nor U29073 (N_29073,N_28629,N_28649);
and U29074 (N_29074,N_28578,N_28582);
nand U29075 (N_29075,N_28581,N_28680);
xnor U29076 (N_29076,N_28626,N_28765);
and U29077 (N_29077,N_28682,N_28671);
nand U29078 (N_29078,N_28569,N_28551);
xnor U29079 (N_29079,N_28534,N_28604);
nor U29080 (N_29080,N_28779,N_28793);
or U29081 (N_29081,N_28661,N_28716);
and U29082 (N_29082,N_28592,N_28604);
xor U29083 (N_29083,N_28639,N_28690);
xnor U29084 (N_29084,N_28688,N_28514);
xnor U29085 (N_29085,N_28700,N_28547);
nor U29086 (N_29086,N_28668,N_28628);
xnor U29087 (N_29087,N_28792,N_28631);
nand U29088 (N_29088,N_28649,N_28739);
or U29089 (N_29089,N_28718,N_28646);
nand U29090 (N_29090,N_28517,N_28749);
nand U29091 (N_29091,N_28770,N_28758);
or U29092 (N_29092,N_28794,N_28630);
xnor U29093 (N_29093,N_28703,N_28649);
nor U29094 (N_29094,N_28503,N_28671);
or U29095 (N_29095,N_28695,N_28513);
or U29096 (N_29096,N_28720,N_28719);
xnor U29097 (N_29097,N_28680,N_28675);
xnor U29098 (N_29098,N_28716,N_28711);
nand U29099 (N_29099,N_28644,N_28600);
and U29100 (N_29100,N_29094,N_28898);
or U29101 (N_29101,N_29048,N_29072);
xnor U29102 (N_29102,N_28950,N_28859);
or U29103 (N_29103,N_28952,N_28979);
nand U29104 (N_29104,N_28995,N_28998);
or U29105 (N_29105,N_28841,N_29035);
xor U29106 (N_29106,N_29006,N_28946);
or U29107 (N_29107,N_29038,N_28965);
xor U29108 (N_29108,N_29053,N_28823);
nor U29109 (N_29109,N_29047,N_28882);
or U29110 (N_29110,N_28832,N_29069);
or U29111 (N_29111,N_28860,N_28909);
nand U29112 (N_29112,N_28991,N_29085);
and U29113 (N_29113,N_28850,N_28902);
xor U29114 (N_29114,N_28887,N_28939);
nand U29115 (N_29115,N_29095,N_29088);
xor U29116 (N_29116,N_28967,N_28918);
or U29117 (N_29117,N_28831,N_28913);
xor U29118 (N_29118,N_29022,N_28906);
nand U29119 (N_29119,N_28890,N_28808);
nand U29120 (N_29120,N_28978,N_28915);
or U29121 (N_29121,N_28815,N_28821);
nand U29122 (N_29122,N_29050,N_28805);
nor U29123 (N_29123,N_28958,N_29019);
or U29124 (N_29124,N_29054,N_28867);
and U29125 (N_29125,N_28833,N_29046);
or U29126 (N_29126,N_28857,N_28973);
nor U29127 (N_29127,N_28835,N_29049);
nand U29128 (N_29128,N_28949,N_29084);
or U29129 (N_29129,N_28907,N_28957);
xor U29130 (N_29130,N_28828,N_28986);
nand U29131 (N_29131,N_29071,N_28938);
nand U29132 (N_29132,N_28836,N_29014);
and U29133 (N_29133,N_29090,N_28800);
xnor U29134 (N_29134,N_28879,N_29075);
nand U29135 (N_29135,N_28925,N_28943);
xor U29136 (N_29136,N_28876,N_28916);
nor U29137 (N_29137,N_29067,N_29000);
nand U29138 (N_29138,N_29086,N_28845);
and U29139 (N_29139,N_28940,N_28842);
or U29140 (N_29140,N_28911,N_28944);
xor U29141 (N_29141,N_28871,N_29063);
and U29142 (N_29142,N_28947,N_29017);
nand U29143 (N_29143,N_28826,N_29015);
xnor U29144 (N_29144,N_28970,N_28830);
or U29145 (N_29145,N_28804,N_28994);
xnor U29146 (N_29146,N_28814,N_29011);
nor U29147 (N_29147,N_28825,N_28877);
nor U29148 (N_29148,N_28985,N_28863);
nand U29149 (N_29149,N_29042,N_28827);
nand U29150 (N_29150,N_29059,N_28945);
and U29151 (N_29151,N_29097,N_28977);
xnor U29152 (N_29152,N_29057,N_28921);
xor U29153 (N_29153,N_29091,N_29068);
nor U29154 (N_29154,N_28920,N_28932);
or U29155 (N_29155,N_29074,N_28904);
nand U29156 (N_29156,N_29016,N_28834);
xor U29157 (N_29157,N_29026,N_28837);
xnor U29158 (N_29158,N_28875,N_28900);
xnor U29159 (N_29159,N_28873,N_28849);
xor U29160 (N_29160,N_28839,N_28852);
xnor U29161 (N_29161,N_29009,N_28853);
and U29162 (N_29162,N_29033,N_28980);
xnor U29163 (N_29163,N_29034,N_29064);
or U29164 (N_29164,N_28865,N_28941);
nor U29165 (N_29165,N_28969,N_28844);
nor U29166 (N_29166,N_28866,N_29044);
or U29167 (N_29167,N_29020,N_29045);
nor U29168 (N_29168,N_28996,N_28955);
or U29169 (N_29169,N_28895,N_28975);
nor U29170 (N_29170,N_29013,N_28838);
nor U29171 (N_29171,N_28948,N_28822);
nand U29172 (N_29172,N_29037,N_28864);
nand U29173 (N_29173,N_29058,N_29024);
nor U29174 (N_29174,N_28893,N_29055);
nand U29175 (N_29175,N_28889,N_28884);
or U29176 (N_29176,N_28930,N_28878);
or U29177 (N_29177,N_29061,N_28910);
nand U29178 (N_29178,N_28960,N_28891);
xor U29179 (N_29179,N_28817,N_28929);
and U29180 (N_29180,N_28869,N_28966);
or U29181 (N_29181,N_29051,N_29089);
or U29182 (N_29182,N_28803,N_28820);
nor U29183 (N_29183,N_28962,N_28905);
nor U29184 (N_29184,N_28931,N_28888);
xor U29185 (N_29185,N_28984,N_28813);
and U29186 (N_29186,N_28851,N_28954);
nor U29187 (N_29187,N_28997,N_28824);
nand U29188 (N_29188,N_29021,N_29030);
or U29189 (N_29189,N_29036,N_28933);
and U29190 (N_29190,N_29066,N_28971);
and U29191 (N_29191,N_28987,N_28801);
and U29192 (N_29192,N_29065,N_29079);
nand U29193 (N_29193,N_28983,N_28829);
nor U29194 (N_29194,N_28848,N_28936);
and U29195 (N_29195,N_28976,N_28874);
nor U29196 (N_29196,N_28992,N_29082);
xor U29197 (N_29197,N_28956,N_28974);
xor U29198 (N_29198,N_29003,N_29098);
and U29199 (N_29199,N_28899,N_28858);
xnor U29200 (N_29200,N_29005,N_28892);
nand U29201 (N_29201,N_28819,N_29029);
and U29202 (N_29202,N_29018,N_28846);
nand U29203 (N_29203,N_28807,N_28885);
or U29204 (N_29204,N_28912,N_28961);
nand U29205 (N_29205,N_28968,N_29080);
xnor U29206 (N_29206,N_28880,N_28964);
nand U29207 (N_29207,N_29012,N_29060);
and U29208 (N_29208,N_28802,N_29083);
nand U29209 (N_29209,N_29078,N_28999);
xor U29210 (N_29210,N_28990,N_28855);
xnor U29211 (N_29211,N_29096,N_28816);
nor U29212 (N_29212,N_28870,N_29025);
and U29213 (N_29213,N_28982,N_28896);
nor U29214 (N_29214,N_29093,N_29087);
and U29215 (N_29215,N_28993,N_29008);
xnor U29216 (N_29216,N_28972,N_29002);
and U29217 (N_29217,N_28959,N_29062);
nand U29218 (N_29218,N_29081,N_28809);
and U29219 (N_29219,N_29077,N_29023);
xor U29220 (N_29220,N_28963,N_28810);
xnor U29221 (N_29221,N_28897,N_28812);
and U29222 (N_29222,N_29032,N_28908);
xor U29223 (N_29223,N_29092,N_29040);
nor U29224 (N_29224,N_29027,N_28942);
xor U29225 (N_29225,N_29028,N_28868);
or U29226 (N_29226,N_28923,N_28937);
and U29227 (N_29227,N_28926,N_29004);
or U29228 (N_29228,N_28924,N_29001);
or U29229 (N_29229,N_29031,N_28818);
and U29230 (N_29230,N_29073,N_28843);
xnor U29231 (N_29231,N_28894,N_29052);
nor U29232 (N_29232,N_29007,N_28981);
xor U29233 (N_29233,N_28927,N_28806);
or U29234 (N_29234,N_28886,N_28862);
or U29235 (N_29235,N_28928,N_28872);
or U29236 (N_29236,N_28935,N_28917);
xnor U29237 (N_29237,N_28901,N_29076);
nand U29238 (N_29238,N_29041,N_29099);
nand U29239 (N_29239,N_28988,N_28861);
and U29240 (N_29240,N_28953,N_28881);
and U29241 (N_29241,N_29043,N_29056);
xnor U29242 (N_29242,N_28883,N_28903);
and U29243 (N_29243,N_28914,N_28951);
xnor U29244 (N_29244,N_28919,N_28840);
or U29245 (N_29245,N_28854,N_28989);
and U29246 (N_29246,N_29010,N_28922);
and U29247 (N_29247,N_29070,N_28856);
and U29248 (N_29248,N_28811,N_28847);
or U29249 (N_29249,N_28934,N_29039);
nor U29250 (N_29250,N_29057,N_29072);
nand U29251 (N_29251,N_28821,N_28813);
nand U29252 (N_29252,N_29027,N_28975);
nor U29253 (N_29253,N_28898,N_28810);
and U29254 (N_29254,N_28976,N_29007);
nor U29255 (N_29255,N_28814,N_29017);
and U29256 (N_29256,N_29055,N_28920);
nor U29257 (N_29257,N_28881,N_29067);
xnor U29258 (N_29258,N_29001,N_29083);
nand U29259 (N_29259,N_29054,N_28986);
or U29260 (N_29260,N_28927,N_28854);
xnor U29261 (N_29261,N_28817,N_28816);
or U29262 (N_29262,N_28964,N_29051);
nor U29263 (N_29263,N_28907,N_28928);
xnor U29264 (N_29264,N_29039,N_28845);
xnor U29265 (N_29265,N_28988,N_28960);
and U29266 (N_29266,N_28908,N_28884);
nor U29267 (N_29267,N_28921,N_28886);
and U29268 (N_29268,N_28883,N_28808);
nor U29269 (N_29269,N_28960,N_28992);
nand U29270 (N_29270,N_28838,N_28958);
xnor U29271 (N_29271,N_28808,N_29090);
xnor U29272 (N_29272,N_29066,N_28855);
and U29273 (N_29273,N_29015,N_28839);
or U29274 (N_29274,N_29098,N_28876);
nor U29275 (N_29275,N_29066,N_28965);
nand U29276 (N_29276,N_28955,N_29019);
nand U29277 (N_29277,N_28803,N_28897);
nand U29278 (N_29278,N_28984,N_29038);
nor U29279 (N_29279,N_28916,N_28879);
nand U29280 (N_29280,N_28954,N_28933);
or U29281 (N_29281,N_28957,N_28976);
nor U29282 (N_29282,N_28801,N_28831);
nor U29283 (N_29283,N_28997,N_28885);
or U29284 (N_29284,N_29011,N_28801);
and U29285 (N_29285,N_28852,N_28959);
and U29286 (N_29286,N_29054,N_28851);
or U29287 (N_29287,N_29012,N_29046);
and U29288 (N_29288,N_28959,N_29009);
xnor U29289 (N_29289,N_28826,N_28863);
and U29290 (N_29290,N_28901,N_28943);
nor U29291 (N_29291,N_28905,N_29087);
and U29292 (N_29292,N_28865,N_28979);
or U29293 (N_29293,N_28866,N_29001);
and U29294 (N_29294,N_28801,N_28886);
and U29295 (N_29295,N_29035,N_29020);
nor U29296 (N_29296,N_28913,N_28919);
nor U29297 (N_29297,N_29027,N_28864);
xnor U29298 (N_29298,N_29031,N_29003);
nand U29299 (N_29299,N_28809,N_29047);
nand U29300 (N_29300,N_28958,N_28926);
nor U29301 (N_29301,N_28808,N_29062);
and U29302 (N_29302,N_29075,N_29040);
xnor U29303 (N_29303,N_28818,N_29092);
or U29304 (N_29304,N_29000,N_28885);
and U29305 (N_29305,N_28854,N_29086);
and U29306 (N_29306,N_28801,N_28955);
xnor U29307 (N_29307,N_28924,N_28815);
xnor U29308 (N_29308,N_28976,N_28803);
xor U29309 (N_29309,N_28805,N_28954);
nor U29310 (N_29310,N_29080,N_28940);
xnor U29311 (N_29311,N_28920,N_29087);
and U29312 (N_29312,N_28803,N_28986);
xor U29313 (N_29313,N_28982,N_29007);
nor U29314 (N_29314,N_29055,N_28801);
and U29315 (N_29315,N_29022,N_29024);
nor U29316 (N_29316,N_29045,N_28916);
nor U29317 (N_29317,N_28836,N_28993);
xor U29318 (N_29318,N_28805,N_28902);
xor U29319 (N_29319,N_28966,N_29047);
and U29320 (N_29320,N_28861,N_28929);
xnor U29321 (N_29321,N_29044,N_29061);
and U29322 (N_29322,N_28973,N_28866);
xnor U29323 (N_29323,N_28874,N_28850);
nor U29324 (N_29324,N_29058,N_28892);
xnor U29325 (N_29325,N_29004,N_28893);
xnor U29326 (N_29326,N_28843,N_29037);
nor U29327 (N_29327,N_28907,N_29080);
nor U29328 (N_29328,N_28907,N_28870);
nor U29329 (N_29329,N_28921,N_29087);
and U29330 (N_29330,N_28835,N_28936);
or U29331 (N_29331,N_28880,N_28888);
or U29332 (N_29332,N_28974,N_28915);
and U29333 (N_29333,N_28922,N_28890);
and U29334 (N_29334,N_28862,N_29033);
nor U29335 (N_29335,N_28828,N_28846);
nor U29336 (N_29336,N_28858,N_28847);
xor U29337 (N_29337,N_28968,N_29093);
and U29338 (N_29338,N_29046,N_28883);
nand U29339 (N_29339,N_29093,N_28815);
or U29340 (N_29340,N_29025,N_28823);
or U29341 (N_29341,N_28909,N_28865);
xnor U29342 (N_29342,N_29041,N_28863);
and U29343 (N_29343,N_29053,N_29002);
nor U29344 (N_29344,N_28919,N_28951);
or U29345 (N_29345,N_29045,N_29008);
nor U29346 (N_29346,N_29026,N_29048);
or U29347 (N_29347,N_28990,N_28934);
nor U29348 (N_29348,N_28893,N_28946);
xnor U29349 (N_29349,N_29055,N_28950);
nand U29350 (N_29350,N_28861,N_28972);
nand U29351 (N_29351,N_28990,N_28996);
and U29352 (N_29352,N_28874,N_29060);
nor U29353 (N_29353,N_29078,N_28950);
nor U29354 (N_29354,N_29013,N_28825);
nand U29355 (N_29355,N_28876,N_28812);
nand U29356 (N_29356,N_28922,N_28867);
or U29357 (N_29357,N_28850,N_28832);
and U29358 (N_29358,N_29084,N_28948);
or U29359 (N_29359,N_28843,N_28918);
xor U29360 (N_29360,N_29096,N_29070);
and U29361 (N_29361,N_29005,N_28989);
or U29362 (N_29362,N_28822,N_28888);
nor U29363 (N_29363,N_28936,N_29053);
nor U29364 (N_29364,N_28923,N_29084);
and U29365 (N_29365,N_28925,N_29027);
nand U29366 (N_29366,N_28828,N_28880);
nor U29367 (N_29367,N_28886,N_28895);
nand U29368 (N_29368,N_28972,N_28919);
and U29369 (N_29369,N_28870,N_29055);
nor U29370 (N_29370,N_28921,N_28930);
xor U29371 (N_29371,N_28866,N_29042);
and U29372 (N_29372,N_29039,N_29029);
and U29373 (N_29373,N_28878,N_28845);
xor U29374 (N_29374,N_29010,N_28824);
or U29375 (N_29375,N_28814,N_28846);
nand U29376 (N_29376,N_29070,N_28868);
nor U29377 (N_29377,N_29007,N_28859);
xnor U29378 (N_29378,N_28811,N_29028);
or U29379 (N_29379,N_28871,N_28900);
and U29380 (N_29380,N_29043,N_29021);
xor U29381 (N_29381,N_28855,N_29083);
nand U29382 (N_29382,N_28953,N_28957);
nand U29383 (N_29383,N_29051,N_28993);
or U29384 (N_29384,N_29089,N_29048);
or U29385 (N_29385,N_28821,N_28966);
xnor U29386 (N_29386,N_28955,N_28943);
and U29387 (N_29387,N_28974,N_29043);
xnor U29388 (N_29388,N_28857,N_28861);
nand U29389 (N_29389,N_28913,N_28834);
or U29390 (N_29390,N_28922,N_29062);
or U29391 (N_29391,N_29099,N_28974);
and U29392 (N_29392,N_28912,N_29037);
or U29393 (N_29393,N_28860,N_29060);
or U29394 (N_29394,N_29034,N_28853);
xnor U29395 (N_29395,N_28847,N_28913);
and U29396 (N_29396,N_28987,N_29011);
or U29397 (N_29397,N_29019,N_28855);
or U29398 (N_29398,N_28838,N_28968);
or U29399 (N_29399,N_28970,N_28998);
and U29400 (N_29400,N_29189,N_29324);
nor U29401 (N_29401,N_29336,N_29173);
and U29402 (N_29402,N_29272,N_29153);
or U29403 (N_29403,N_29318,N_29142);
and U29404 (N_29404,N_29162,N_29190);
and U29405 (N_29405,N_29184,N_29216);
and U29406 (N_29406,N_29207,N_29244);
xor U29407 (N_29407,N_29285,N_29210);
xor U29408 (N_29408,N_29140,N_29155);
or U29409 (N_29409,N_29342,N_29352);
nand U29410 (N_29410,N_29350,N_29289);
xor U29411 (N_29411,N_29167,N_29214);
nor U29412 (N_29412,N_29298,N_29398);
or U29413 (N_29413,N_29371,N_29206);
nand U29414 (N_29414,N_29123,N_29312);
nor U29415 (N_29415,N_29107,N_29311);
xnor U29416 (N_29416,N_29106,N_29361);
or U29417 (N_29417,N_29275,N_29358);
and U29418 (N_29418,N_29227,N_29302);
or U29419 (N_29419,N_29183,N_29316);
and U29420 (N_29420,N_29369,N_29322);
xor U29421 (N_29421,N_29362,N_29177);
nand U29422 (N_29422,N_29135,N_29105);
or U29423 (N_29423,N_29213,N_29327);
nand U29424 (N_29424,N_29328,N_29198);
or U29425 (N_29425,N_29228,N_29335);
nand U29426 (N_29426,N_29329,N_29175);
nor U29427 (N_29427,N_29136,N_29372);
and U29428 (N_29428,N_29197,N_29337);
xor U29429 (N_29429,N_29351,N_29345);
xor U29430 (N_29430,N_29286,N_29117);
nand U29431 (N_29431,N_29249,N_29178);
and U29432 (N_29432,N_29170,N_29268);
or U29433 (N_29433,N_29278,N_29137);
nand U29434 (N_29434,N_29396,N_29163);
xnor U29435 (N_29435,N_29200,N_29250);
xnor U29436 (N_29436,N_29113,N_29118);
or U29437 (N_29437,N_29386,N_29165);
nor U29438 (N_29438,N_29147,N_29265);
xnor U29439 (N_29439,N_29259,N_29264);
or U29440 (N_29440,N_29299,N_29271);
xor U29441 (N_29441,N_29252,N_29168);
nand U29442 (N_29442,N_29180,N_29120);
nor U29443 (N_29443,N_29330,N_29219);
nor U29444 (N_29444,N_29293,N_29157);
nor U29445 (N_29445,N_29194,N_29287);
nor U29446 (N_29446,N_29374,N_29317);
and U29447 (N_29447,N_29347,N_29122);
and U29448 (N_29448,N_29395,N_29236);
xnor U29449 (N_29449,N_29392,N_29161);
nor U29450 (N_29450,N_29338,N_29295);
or U29451 (N_29451,N_29381,N_29368);
or U29452 (N_29452,N_29232,N_29121);
or U29453 (N_29453,N_29196,N_29111);
or U29454 (N_29454,N_29367,N_29127);
or U29455 (N_29455,N_29334,N_29225);
and U29456 (N_29456,N_29388,N_29256);
xor U29457 (N_29457,N_29291,N_29365);
nand U29458 (N_29458,N_29364,N_29116);
and U29459 (N_29459,N_29212,N_29319);
and U29460 (N_29460,N_29217,N_29130);
nand U29461 (N_29461,N_29282,N_29199);
and U29462 (N_29462,N_29229,N_29174);
nor U29463 (N_29463,N_29263,N_29380);
and U29464 (N_29464,N_29208,N_29308);
nand U29465 (N_29465,N_29280,N_29304);
or U29466 (N_29466,N_29223,N_29139);
or U29467 (N_29467,N_29195,N_29211);
or U29468 (N_29468,N_29193,N_29104);
xnor U29469 (N_29469,N_29145,N_29297);
nand U29470 (N_29470,N_29235,N_29389);
and U29471 (N_29471,N_29378,N_29301);
xor U29472 (N_29472,N_29273,N_29357);
and U29473 (N_29473,N_29333,N_29240);
nor U29474 (N_29474,N_29391,N_29226);
or U29475 (N_29475,N_29377,N_29158);
or U29476 (N_29476,N_29332,N_29233);
nor U29477 (N_29477,N_29239,N_29245);
and U29478 (N_29478,N_29218,N_29313);
xnor U29479 (N_29479,N_29292,N_29128);
nor U29480 (N_29480,N_29185,N_29192);
xnor U29481 (N_29481,N_29166,N_29255);
nor U29482 (N_29482,N_29186,N_29284);
xor U29483 (N_29483,N_29363,N_29237);
and U29484 (N_29484,N_29230,N_29151);
nor U29485 (N_29485,N_29394,N_29320);
or U29486 (N_29486,N_29114,N_29187);
or U29487 (N_29487,N_29154,N_29124);
nand U29488 (N_29488,N_29254,N_29132);
or U29489 (N_29489,N_29296,N_29385);
xnor U29490 (N_29490,N_29310,N_29150);
nand U29491 (N_29491,N_29274,N_29376);
and U29492 (N_29492,N_29270,N_29182);
or U29493 (N_29493,N_29246,N_29129);
nand U29494 (N_29494,N_29305,N_29181);
nor U29495 (N_29495,N_29343,N_29300);
nand U29496 (N_29496,N_29397,N_29191);
and U29497 (N_29497,N_29146,N_29205);
or U29498 (N_29498,N_29257,N_29148);
xnor U29499 (N_29499,N_29100,N_29115);
nor U29500 (N_29500,N_29108,N_29281);
nor U29501 (N_29501,N_29138,N_29288);
or U29502 (N_29502,N_29315,N_29202);
nor U29503 (N_29503,N_29258,N_29366);
nand U29504 (N_29504,N_29248,N_29179);
xor U29505 (N_29505,N_29387,N_29125);
nor U29506 (N_29506,N_29353,N_29346);
or U29507 (N_29507,N_29399,N_29266);
nand U29508 (N_29508,N_29359,N_29110);
or U29509 (N_29509,N_29188,N_29382);
xor U29510 (N_29510,N_29215,N_29390);
and U29511 (N_29511,N_29370,N_29325);
xor U29512 (N_29512,N_29156,N_29231);
nor U29513 (N_29513,N_29109,N_29241);
or U29514 (N_29514,N_29224,N_29251);
nor U29515 (N_29515,N_29279,N_29341);
or U29516 (N_29516,N_29339,N_29326);
xor U29517 (N_29517,N_29303,N_29238);
xor U29518 (N_29518,N_29204,N_29262);
nand U29519 (N_29519,N_29373,N_29314);
and U29520 (N_29520,N_29159,N_29201);
nand U29521 (N_29521,N_29375,N_29349);
xor U29522 (N_29522,N_29383,N_29141);
nand U29523 (N_29523,N_29294,N_29393);
nor U29524 (N_29524,N_29354,N_29149);
nand U29525 (N_29525,N_29355,N_29222);
or U29526 (N_29526,N_29323,N_29176);
and U29527 (N_29527,N_29112,N_29344);
or U29528 (N_29528,N_29133,N_29253);
or U29529 (N_29529,N_29203,N_29321);
xor U29530 (N_29530,N_29277,N_29290);
or U29531 (N_29531,N_29220,N_29283);
or U29532 (N_29532,N_29243,N_29309);
xnor U29533 (N_29533,N_29209,N_29267);
xor U29534 (N_29534,N_29169,N_29160);
xor U29535 (N_29535,N_29276,N_29260);
xor U29536 (N_29536,N_29152,N_29306);
nor U29537 (N_29537,N_29103,N_29143);
and U29538 (N_29538,N_29119,N_29331);
and U29539 (N_29539,N_29384,N_29348);
or U29540 (N_29540,N_29242,N_29247);
xor U29541 (N_29541,N_29101,N_29126);
nor U29542 (N_29542,N_29171,N_29172);
and U29543 (N_29543,N_29234,N_29164);
or U29544 (N_29544,N_29340,N_29102);
and U29545 (N_29545,N_29131,N_29134);
and U29546 (N_29546,N_29360,N_29261);
nand U29547 (N_29547,N_29307,N_29221);
and U29548 (N_29548,N_29144,N_29356);
xnor U29549 (N_29549,N_29269,N_29379);
or U29550 (N_29550,N_29307,N_29277);
xor U29551 (N_29551,N_29362,N_29115);
or U29552 (N_29552,N_29204,N_29148);
or U29553 (N_29553,N_29185,N_29199);
and U29554 (N_29554,N_29274,N_29335);
nor U29555 (N_29555,N_29185,N_29176);
and U29556 (N_29556,N_29144,N_29148);
nand U29557 (N_29557,N_29149,N_29379);
nand U29558 (N_29558,N_29380,N_29180);
xnor U29559 (N_29559,N_29356,N_29243);
or U29560 (N_29560,N_29161,N_29189);
or U29561 (N_29561,N_29248,N_29261);
nand U29562 (N_29562,N_29115,N_29277);
or U29563 (N_29563,N_29337,N_29247);
and U29564 (N_29564,N_29292,N_29217);
or U29565 (N_29565,N_29226,N_29370);
xor U29566 (N_29566,N_29112,N_29374);
nor U29567 (N_29567,N_29121,N_29279);
xor U29568 (N_29568,N_29358,N_29271);
nor U29569 (N_29569,N_29148,N_29307);
or U29570 (N_29570,N_29389,N_29219);
nand U29571 (N_29571,N_29204,N_29245);
nor U29572 (N_29572,N_29395,N_29288);
nor U29573 (N_29573,N_29318,N_29181);
nand U29574 (N_29574,N_29152,N_29308);
or U29575 (N_29575,N_29372,N_29239);
nand U29576 (N_29576,N_29156,N_29216);
or U29577 (N_29577,N_29347,N_29371);
nand U29578 (N_29578,N_29229,N_29124);
xnor U29579 (N_29579,N_29102,N_29316);
or U29580 (N_29580,N_29365,N_29120);
and U29581 (N_29581,N_29315,N_29103);
nand U29582 (N_29582,N_29166,N_29189);
xor U29583 (N_29583,N_29106,N_29359);
nor U29584 (N_29584,N_29323,N_29285);
or U29585 (N_29585,N_29323,N_29105);
nand U29586 (N_29586,N_29349,N_29111);
nand U29587 (N_29587,N_29102,N_29241);
and U29588 (N_29588,N_29144,N_29339);
or U29589 (N_29589,N_29136,N_29131);
nor U29590 (N_29590,N_29145,N_29352);
xor U29591 (N_29591,N_29275,N_29360);
and U29592 (N_29592,N_29377,N_29172);
nor U29593 (N_29593,N_29263,N_29368);
nand U29594 (N_29594,N_29158,N_29200);
and U29595 (N_29595,N_29365,N_29298);
nand U29596 (N_29596,N_29243,N_29251);
or U29597 (N_29597,N_29350,N_29300);
xor U29598 (N_29598,N_29106,N_29101);
nor U29599 (N_29599,N_29388,N_29182);
nand U29600 (N_29600,N_29234,N_29392);
nor U29601 (N_29601,N_29156,N_29187);
nor U29602 (N_29602,N_29398,N_29194);
or U29603 (N_29603,N_29325,N_29380);
and U29604 (N_29604,N_29261,N_29242);
nand U29605 (N_29605,N_29178,N_29358);
and U29606 (N_29606,N_29210,N_29148);
nand U29607 (N_29607,N_29200,N_29268);
nand U29608 (N_29608,N_29276,N_29219);
or U29609 (N_29609,N_29133,N_29370);
nand U29610 (N_29610,N_29345,N_29271);
or U29611 (N_29611,N_29273,N_29227);
nand U29612 (N_29612,N_29330,N_29299);
nand U29613 (N_29613,N_29242,N_29325);
and U29614 (N_29614,N_29364,N_29375);
and U29615 (N_29615,N_29195,N_29389);
nand U29616 (N_29616,N_29107,N_29248);
and U29617 (N_29617,N_29194,N_29165);
and U29618 (N_29618,N_29344,N_29274);
nand U29619 (N_29619,N_29335,N_29299);
nor U29620 (N_29620,N_29102,N_29350);
and U29621 (N_29621,N_29210,N_29310);
and U29622 (N_29622,N_29336,N_29246);
nor U29623 (N_29623,N_29329,N_29312);
or U29624 (N_29624,N_29254,N_29117);
nor U29625 (N_29625,N_29358,N_29204);
or U29626 (N_29626,N_29264,N_29104);
or U29627 (N_29627,N_29249,N_29381);
and U29628 (N_29628,N_29366,N_29269);
nor U29629 (N_29629,N_29285,N_29172);
nor U29630 (N_29630,N_29222,N_29354);
and U29631 (N_29631,N_29286,N_29236);
xnor U29632 (N_29632,N_29109,N_29217);
and U29633 (N_29633,N_29124,N_29209);
and U29634 (N_29634,N_29380,N_29134);
xnor U29635 (N_29635,N_29390,N_29263);
xor U29636 (N_29636,N_29222,N_29147);
nor U29637 (N_29637,N_29281,N_29249);
xnor U29638 (N_29638,N_29299,N_29200);
or U29639 (N_29639,N_29271,N_29368);
nand U29640 (N_29640,N_29318,N_29396);
nand U29641 (N_29641,N_29216,N_29308);
nand U29642 (N_29642,N_29227,N_29330);
xor U29643 (N_29643,N_29376,N_29246);
or U29644 (N_29644,N_29250,N_29282);
and U29645 (N_29645,N_29124,N_29234);
and U29646 (N_29646,N_29289,N_29133);
nor U29647 (N_29647,N_29305,N_29162);
or U29648 (N_29648,N_29197,N_29221);
xnor U29649 (N_29649,N_29142,N_29121);
xnor U29650 (N_29650,N_29111,N_29124);
xnor U29651 (N_29651,N_29298,N_29380);
and U29652 (N_29652,N_29110,N_29315);
or U29653 (N_29653,N_29106,N_29399);
nor U29654 (N_29654,N_29212,N_29361);
nand U29655 (N_29655,N_29315,N_29303);
nand U29656 (N_29656,N_29202,N_29255);
or U29657 (N_29657,N_29351,N_29204);
and U29658 (N_29658,N_29152,N_29202);
or U29659 (N_29659,N_29358,N_29355);
or U29660 (N_29660,N_29356,N_29188);
nand U29661 (N_29661,N_29334,N_29182);
or U29662 (N_29662,N_29301,N_29190);
or U29663 (N_29663,N_29119,N_29297);
nand U29664 (N_29664,N_29300,N_29141);
xnor U29665 (N_29665,N_29325,N_29105);
nor U29666 (N_29666,N_29397,N_29271);
nor U29667 (N_29667,N_29334,N_29106);
or U29668 (N_29668,N_29223,N_29177);
nand U29669 (N_29669,N_29381,N_29101);
and U29670 (N_29670,N_29283,N_29278);
and U29671 (N_29671,N_29303,N_29110);
or U29672 (N_29672,N_29113,N_29194);
xor U29673 (N_29673,N_29114,N_29385);
or U29674 (N_29674,N_29200,N_29244);
nand U29675 (N_29675,N_29385,N_29390);
xnor U29676 (N_29676,N_29322,N_29149);
xnor U29677 (N_29677,N_29381,N_29110);
or U29678 (N_29678,N_29198,N_29298);
nand U29679 (N_29679,N_29167,N_29307);
nand U29680 (N_29680,N_29349,N_29225);
xor U29681 (N_29681,N_29254,N_29371);
nor U29682 (N_29682,N_29341,N_29142);
or U29683 (N_29683,N_29125,N_29100);
nor U29684 (N_29684,N_29185,N_29264);
and U29685 (N_29685,N_29175,N_29301);
nand U29686 (N_29686,N_29346,N_29242);
or U29687 (N_29687,N_29220,N_29203);
nand U29688 (N_29688,N_29344,N_29341);
xnor U29689 (N_29689,N_29336,N_29109);
or U29690 (N_29690,N_29205,N_29265);
nor U29691 (N_29691,N_29146,N_29260);
nand U29692 (N_29692,N_29328,N_29258);
or U29693 (N_29693,N_29312,N_29247);
xnor U29694 (N_29694,N_29183,N_29178);
xnor U29695 (N_29695,N_29156,N_29347);
nand U29696 (N_29696,N_29326,N_29203);
nor U29697 (N_29697,N_29184,N_29352);
and U29698 (N_29698,N_29333,N_29311);
xnor U29699 (N_29699,N_29132,N_29203);
and U29700 (N_29700,N_29454,N_29537);
nor U29701 (N_29701,N_29479,N_29651);
or U29702 (N_29702,N_29517,N_29578);
nand U29703 (N_29703,N_29459,N_29443);
or U29704 (N_29704,N_29629,N_29452);
and U29705 (N_29705,N_29694,N_29473);
and U29706 (N_29706,N_29676,N_29530);
nor U29707 (N_29707,N_29531,N_29483);
nand U29708 (N_29708,N_29668,N_29634);
or U29709 (N_29709,N_29592,N_29573);
nor U29710 (N_29710,N_29604,N_29422);
xor U29711 (N_29711,N_29491,N_29628);
nor U29712 (N_29712,N_29497,N_29420);
or U29713 (N_29713,N_29402,N_29539);
nor U29714 (N_29714,N_29632,N_29476);
xor U29715 (N_29715,N_29579,N_29412);
or U29716 (N_29716,N_29490,N_29418);
xnor U29717 (N_29717,N_29552,N_29577);
nand U29718 (N_29718,N_29563,N_29435);
nand U29719 (N_29719,N_29696,N_29515);
xnor U29720 (N_29720,N_29662,N_29607);
or U29721 (N_29721,N_29414,N_29528);
xor U29722 (N_29722,N_29511,N_29656);
nand U29723 (N_29723,N_29529,N_29618);
and U29724 (N_29724,N_29602,N_29620);
and U29725 (N_29725,N_29545,N_29465);
and U29726 (N_29726,N_29434,N_29448);
nand U29727 (N_29727,N_29400,N_29635);
or U29728 (N_29728,N_29482,N_29588);
nand U29729 (N_29729,N_29493,N_29675);
or U29730 (N_29730,N_29419,N_29468);
nand U29731 (N_29731,N_29679,N_29514);
or U29732 (N_29732,N_29432,N_29469);
or U29733 (N_29733,N_29599,N_29569);
xor U29734 (N_29734,N_29590,N_29553);
xnor U29735 (N_29735,N_29534,N_29571);
xor U29736 (N_29736,N_29484,N_29547);
and U29737 (N_29737,N_29644,N_29560);
xnor U29738 (N_29738,N_29608,N_29438);
or U29739 (N_29739,N_29688,N_29646);
xnor U29740 (N_29740,N_29404,N_29671);
or U29741 (N_29741,N_29666,N_29401);
nor U29742 (N_29742,N_29555,N_29594);
nor U29743 (N_29743,N_29472,N_29508);
and U29744 (N_29744,N_29437,N_29458);
xnor U29745 (N_29745,N_29558,N_29501);
nor U29746 (N_29746,N_29466,N_29562);
xor U29747 (N_29747,N_29664,N_29546);
nand U29748 (N_29748,N_29496,N_29647);
and U29749 (N_29749,N_29498,N_29684);
nand U29750 (N_29750,N_29587,N_29533);
nor U29751 (N_29751,N_29518,N_29663);
or U29752 (N_29752,N_29523,N_29591);
or U29753 (N_29753,N_29660,N_29674);
or U29754 (N_29754,N_29415,N_29504);
or U29755 (N_29755,N_29509,N_29446);
xor U29756 (N_29756,N_29596,N_29503);
nor U29757 (N_29757,N_29595,N_29695);
xor U29758 (N_29758,N_29642,N_29568);
and U29759 (N_29759,N_29673,N_29538);
nor U29760 (N_29760,N_29626,N_29680);
xor U29761 (N_29761,N_29630,N_29416);
xnor U29762 (N_29762,N_29460,N_29580);
or U29763 (N_29763,N_29593,N_29625);
nand U29764 (N_29764,N_29597,N_29697);
xor U29765 (N_29765,N_29510,N_29450);
nand U29766 (N_29766,N_29665,N_29502);
nand U29767 (N_29767,N_29639,N_29406);
nand U29768 (N_29768,N_29619,N_29551);
nand U29769 (N_29769,N_29512,N_29661);
xnor U29770 (N_29770,N_29451,N_29691);
nor U29771 (N_29771,N_29427,N_29506);
xnor U29772 (N_29772,N_29487,N_29544);
or U29773 (N_29773,N_29576,N_29407);
nor U29774 (N_29774,N_29658,N_29655);
or U29775 (N_29775,N_29447,N_29631);
or U29776 (N_29776,N_29669,N_29672);
nand U29777 (N_29777,N_29601,N_29456);
or U29778 (N_29778,N_29425,N_29521);
or U29779 (N_29779,N_29471,N_29535);
xnor U29780 (N_29780,N_29582,N_29565);
xnor U29781 (N_29781,N_29690,N_29621);
and U29782 (N_29782,N_29481,N_29598);
and U29783 (N_29783,N_29645,N_29572);
or U29784 (N_29784,N_29606,N_29526);
xor U29785 (N_29785,N_29623,N_29433);
xor U29786 (N_29786,N_29505,N_29648);
or U29787 (N_29787,N_29439,N_29559);
or U29788 (N_29788,N_29636,N_29603);
and U29789 (N_29789,N_29457,N_29532);
nand U29790 (N_29790,N_29683,N_29507);
xor U29791 (N_29791,N_29612,N_29605);
nor U29792 (N_29792,N_29403,N_29522);
nor U29793 (N_29793,N_29677,N_29462);
and U29794 (N_29794,N_29678,N_29453);
nand U29795 (N_29795,N_29566,N_29442);
and U29796 (N_29796,N_29583,N_29516);
nor U29797 (N_29797,N_29474,N_29567);
and U29798 (N_29798,N_29586,N_29467);
xnor U29799 (N_29799,N_29637,N_29436);
or U29800 (N_29800,N_29653,N_29525);
or U29801 (N_29801,N_29429,N_29627);
nand U29802 (N_29802,N_29652,N_29486);
and U29803 (N_29803,N_29440,N_29540);
nand U29804 (N_29804,N_29609,N_29411);
and U29805 (N_29805,N_29575,N_29692);
nand U29806 (N_29806,N_29417,N_29654);
or U29807 (N_29807,N_29622,N_29640);
nand U29808 (N_29808,N_29408,N_29681);
xor U29809 (N_29809,N_29570,N_29556);
nand U29810 (N_29810,N_29513,N_29520);
and U29811 (N_29811,N_29478,N_29423);
nor U29812 (N_29812,N_29430,N_29477);
nand U29813 (N_29813,N_29421,N_29500);
or U29814 (N_29814,N_29624,N_29686);
xor U29815 (N_29815,N_29461,N_29492);
xor U29816 (N_29816,N_29633,N_29614);
xnor U29817 (N_29817,N_29541,N_29693);
nor U29818 (N_29818,N_29689,N_29698);
nand U29819 (N_29819,N_29499,N_29641);
or U29820 (N_29820,N_29557,N_29561);
or U29821 (N_29821,N_29410,N_29613);
xor U29822 (N_29822,N_29519,N_29475);
or U29823 (N_29823,N_29649,N_29494);
nand U29824 (N_29824,N_29413,N_29616);
xnor U29825 (N_29825,N_29554,N_29550);
or U29826 (N_29826,N_29659,N_29638);
nor U29827 (N_29827,N_29480,N_29441);
and U29828 (N_29828,N_29424,N_29574);
or U29829 (N_29829,N_29488,N_29650);
nor U29830 (N_29830,N_29428,N_29464);
xor U29831 (N_29831,N_29584,N_29610);
nand U29832 (N_29832,N_29682,N_29687);
xnor U29833 (N_29833,N_29548,N_29527);
nand U29834 (N_29834,N_29485,N_29431);
and U29835 (N_29835,N_29455,N_29657);
and U29836 (N_29836,N_29536,N_29489);
nor U29837 (N_29837,N_29543,N_29405);
or U29838 (N_29838,N_29495,N_29409);
nor U29839 (N_29839,N_29564,N_29449);
or U29840 (N_29840,N_29444,N_29470);
nand U29841 (N_29841,N_29617,N_29549);
nor U29842 (N_29842,N_29585,N_29426);
and U29843 (N_29843,N_29643,N_29699);
nand U29844 (N_29844,N_29445,N_29463);
nor U29845 (N_29845,N_29615,N_29685);
nor U29846 (N_29846,N_29542,N_29524);
or U29847 (N_29847,N_29667,N_29600);
and U29848 (N_29848,N_29589,N_29611);
and U29849 (N_29849,N_29670,N_29581);
and U29850 (N_29850,N_29433,N_29506);
nand U29851 (N_29851,N_29655,N_29563);
or U29852 (N_29852,N_29678,N_29502);
xor U29853 (N_29853,N_29521,N_29593);
nand U29854 (N_29854,N_29699,N_29649);
and U29855 (N_29855,N_29628,N_29657);
and U29856 (N_29856,N_29467,N_29681);
and U29857 (N_29857,N_29518,N_29488);
or U29858 (N_29858,N_29501,N_29675);
xor U29859 (N_29859,N_29557,N_29562);
xor U29860 (N_29860,N_29495,N_29652);
xnor U29861 (N_29861,N_29563,N_29553);
nand U29862 (N_29862,N_29483,N_29667);
nor U29863 (N_29863,N_29453,N_29462);
and U29864 (N_29864,N_29404,N_29544);
nor U29865 (N_29865,N_29581,N_29640);
nor U29866 (N_29866,N_29617,N_29515);
and U29867 (N_29867,N_29571,N_29483);
xnor U29868 (N_29868,N_29404,N_29689);
nand U29869 (N_29869,N_29526,N_29637);
xor U29870 (N_29870,N_29662,N_29486);
or U29871 (N_29871,N_29607,N_29470);
and U29872 (N_29872,N_29630,N_29459);
nand U29873 (N_29873,N_29483,N_29475);
or U29874 (N_29874,N_29614,N_29685);
nand U29875 (N_29875,N_29692,N_29612);
nor U29876 (N_29876,N_29621,N_29648);
nand U29877 (N_29877,N_29689,N_29443);
nand U29878 (N_29878,N_29694,N_29406);
and U29879 (N_29879,N_29410,N_29637);
xnor U29880 (N_29880,N_29616,N_29665);
or U29881 (N_29881,N_29605,N_29637);
nor U29882 (N_29882,N_29624,N_29594);
and U29883 (N_29883,N_29589,N_29560);
and U29884 (N_29884,N_29637,N_29691);
nor U29885 (N_29885,N_29486,N_29463);
xor U29886 (N_29886,N_29437,N_29527);
xnor U29887 (N_29887,N_29615,N_29494);
nand U29888 (N_29888,N_29478,N_29660);
and U29889 (N_29889,N_29454,N_29690);
and U29890 (N_29890,N_29501,N_29534);
nor U29891 (N_29891,N_29441,N_29415);
nor U29892 (N_29892,N_29604,N_29470);
nand U29893 (N_29893,N_29657,N_29515);
nand U29894 (N_29894,N_29589,N_29535);
nor U29895 (N_29895,N_29491,N_29678);
and U29896 (N_29896,N_29687,N_29424);
nand U29897 (N_29897,N_29402,N_29612);
and U29898 (N_29898,N_29457,N_29535);
or U29899 (N_29899,N_29541,N_29588);
nand U29900 (N_29900,N_29626,N_29687);
nor U29901 (N_29901,N_29412,N_29658);
or U29902 (N_29902,N_29696,N_29650);
and U29903 (N_29903,N_29670,N_29527);
xor U29904 (N_29904,N_29592,N_29451);
nand U29905 (N_29905,N_29500,N_29435);
xnor U29906 (N_29906,N_29561,N_29506);
or U29907 (N_29907,N_29443,N_29551);
or U29908 (N_29908,N_29570,N_29523);
and U29909 (N_29909,N_29608,N_29511);
and U29910 (N_29910,N_29682,N_29405);
and U29911 (N_29911,N_29647,N_29581);
and U29912 (N_29912,N_29606,N_29582);
nor U29913 (N_29913,N_29659,N_29535);
and U29914 (N_29914,N_29590,N_29435);
nor U29915 (N_29915,N_29614,N_29649);
xnor U29916 (N_29916,N_29655,N_29562);
and U29917 (N_29917,N_29430,N_29695);
nor U29918 (N_29918,N_29483,N_29515);
nand U29919 (N_29919,N_29573,N_29486);
or U29920 (N_29920,N_29482,N_29476);
or U29921 (N_29921,N_29651,N_29507);
or U29922 (N_29922,N_29535,N_29427);
nand U29923 (N_29923,N_29694,N_29491);
xnor U29924 (N_29924,N_29458,N_29663);
nor U29925 (N_29925,N_29570,N_29455);
xor U29926 (N_29926,N_29507,N_29414);
nor U29927 (N_29927,N_29590,N_29660);
and U29928 (N_29928,N_29607,N_29474);
nor U29929 (N_29929,N_29618,N_29408);
nor U29930 (N_29930,N_29641,N_29554);
or U29931 (N_29931,N_29581,N_29464);
or U29932 (N_29932,N_29481,N_29431);
and U29933 (N_29933,N_29599,N_29461);
or U29934 (N_29934,N_29682,N_29577);
xor U29935 (N_29935,N_29485,N_29660);
nand U29936 (N_29936,N_29404,N_29556);
or U29937 (N_29937,N_29563,N_29557);
nor U29938 (N_29938,N_29482,N_29523);
nor U29939 (N_29939,N_29564,N_29571);
and U29940 (N_29940,N_29409,N_29693);
xnor U29941 (N_29941,N_29667,N_29488);
nor U29942 (N_29942,N_29402,N_29682);
and U29943 (N_29943,N_29478,N_29647);
and U29944 (N_29944,N_29686,N_29521);
nor U29945 (N_29945,N_29565,N_29640);
nand U29946 (N_29946,N_29595,N_29527);
nand U29947 (N_29947,N_29653,N_29465);
nand U29948 (N_29948,N_29699,N_29599);
nand U29949 (N_29949,N_29454,N_29678);
and U29950 (N_29950,N_29661,N_29516);
or U29951 (N_29951,N_29534,N_29402);
and U29952 (N_29952,N_29553,N_29627);
nand U29953 (N_29953,N_29502,N_29497);
xor U29954 (N_29954,N_29635,N_29448);
and U29955 (N_29955,N_29632,N_29698);
nor U29956 (N_29956,N_29446,N_29668);
nand U29957 (N_29957,N_29659,N_29542);
and U29958 (N_29958,N_29464,N_29592);
and U29959 (N_29959,N_29498,N_29419);
or U29960 (N_29960,N_29561,N_29594);
or U29961 (N_29961,N_29526,N_29648);
nand U29962 (N_29962,N_29448,N_29614);
nand U29963 (N_29963,N_29605,N_29442);
nor U29964 (N_29964,N_29455,N_29419);
and U29965 (N_29965,N_29522,N_29519);
or U29966 (N_29966,N_29537,N_29481);
and U29967 (N_29967,N_29698,N_29674);
xor U29968 (N_29968,N_29486,N_29616);
xor U29969 (N_29969,N_29524,N_29467);
or U29970 (N_29970,N_29586,N_29609);
or U29971 (N_29971,N_29560,N_29466);
nor U29972 (N_29972,N_29645,N_29578);
nand U29973 (N_29973,N_29688,N_29565);
xnor U29974 (N_29974,N_29447,N_29445);
xnor U29975 (N_29975,N_29559,N_29684);
nand U29976 (N_29976,N_29401,N_29623);
or U29977 (N_29977,N_29682,N_29416);
nand U29978 (N_29978,N_29562,N_29561);
or U29979 (N_29979,N_29685,N_29443);
nor U29980 (N_29980,N_29433,N_29477);
or U29981 (N_29981,N_29623,N_29524);
xnor U29982 (N_29982,N_29494,N_29619);
or U29983 (N_29983,N_29522,N_29551);
or U29984 (N_29984,N_29604,N_29660);
xnor U29985 (N_29985,N_29531,N_29597);
or U29986 (N_29986,N_29685,N_29525);
xor U29987 (N_29987,N_29641,N_29518);
nand U29988 (N_29988,N_29660,N_29461);
nand U29989 (N_29989,N_29591,N_29628);
and U29990 (N_29990,N_29683,N_29554);
or U29991 (N_29991,N_29574,N_29458);
or U29992 (N_29992,N_29481,N_29445);
nor U29993 (N_29993,N_29551,N_29485);
xor U29994 (N_29994,N_29509,N_29521);
nor U29995 (N_29995,N_29454,N_29484);
nor U29996 (N_29996,N_29405,N_29499);
or U29997 (N_29997,N_29411,N_29459);
and U29998 (N_29998,N_29486,N_29647);
or U29999 (N_29999,N_29597,N_29595);
nand UO_0 (O_0,N_29876,N_29709);
or UO_1 (O_1,N_29742,N_29814);
nand UO_2 (O_2,N_29800,N_29929);
nor UO_3 (O_3,N_29702,N_29995);
nor UO_4 (O_4,N_29955,N_29763);
nor UO_5 (O_5,N_29846,N_29787);
nor UO_6 (O_6,N_29915,N_29992);
nand UO_7 (O_7,N_29749,N_29966);
or UO_8 (O_8,N_29996,N_29991);
nor UO_9 (O_9,N_29808,N_29851);
nor UO_10 (O_10,N_29840,N_29874);
and UO_11 (O_11,N_29938,N_29987);
nor UO_12 (O_12,N_29954,N_29869);
nand UO_13 (O_13,N_29914,N_29871);
xnor UO_14 (O_14,N_29843,N_29827);
xor UO_15 (O_15,N_29852,N_29853);
or UO_16 (O_16,N_29792,N_29730);
or UO_17 (O_17,N_29897,N_29811);
and UO_18 (O_18,N_29816,N_29728);
xor UO_19 (O_19,N_29708,N_29879);
or UO_20 (O_20,N_29945,N_29837);
or UO_21 (O_21,N_29902,N_29986);
xor UO_22 (O_22,N_29860,N_29981);
and UO_23 (O_23,N_29822,N_29927);
or UO_24 (O_24,N_29724,N_29901);
nor UO_25 (O_25,N_29810,N_29976);
nor UO_26 (O_26,N_29799,N_29747);
xor UO_27 (O_27,N_29812,N_29834);
or UO_28 (O_28,N_29909,N_29705);
and UO_29 (O_29,N_29952,N_29790);
or UO_30 (O_30,N_29971,N_29739);
and UO_31 (O_31,N_29965,N_29823);
and UO_32 (O_32,N_29796,N_29972);
nand UO_33 (O_33,N_29795,N_29942);
xnor UO_34 (O_34,N_29782,N_29865);
or UO_35 (O_35,N_29813,N_29737);
nor UO_36 (O_36,N_29912,N_29907);
nand UO_37 (O_37,N_29890,N_29707);
xor UO_38 (O_38,N_29819,N_29752);
nor UO_39 (O_39,N_29788,N_29805);
or UO_40 (O_40,N_29974,N_29836);
or UO_41 (O_41,N_29773,N_29714);
xnor UO_42 (O_42,N_29855,N_29826);
nor UO_43 (O_43,N_29900,N_29844);
nand UO_44 (O_44,N_29839,N_29777);
or UO_45 (O_45,N_29778,N_29825);
and UO_46 (O_46,N_29875,N_29940);
and UO_47 (O_47,N_29804,N_29990);
and UO_48 (O_48,N_29740,N_29734);
xor UO_49 (O_49,N_29771,N_29960);
or UO_50 (O_50,N_29998,N_29759);
nor UO_51 (O_51,N_29849,N_29722);
and UO_52 (O_52,N_29946,N_29815);
and UO_53 (O_53,N_29729,N_29781);
and UO_54 (O_54,N_29797,N_29889);
nand UO_55 (O_55,N_29780,N_29937);
and UO_56 (O_56,N_29703,N_29906);
or UO_57 (O_57,N_29953,N_29873);
xor UO_58 (O_58,N_29726,N_29764);
or UO_59 (O_59,N_29918,N_29828);
nor UO_60 (O_60,N_29854,N_29895);
or UO_61 (O_61,N_29956,N_29924);
nor UO_62 (O_62,N_29881,N_29775);
or UO_63 (O_63,N_29923,N_29803);
nor UO_64 (O_64,N_29993,N_29717);
or UO_65 (O_65,N_29985,N_29809);
xor UO_66 (O_66,N_29761,N_29861);
nor UO_67 (O_67,N_29720,N_29975);
nand UO_68 (O_68,N_29892,N_29857);
or UO_69 (O_69,N_29922,N_29719);
xor UO_70 (O_70,N_29725,N_29829);
nor UO_71 (O_71,N_29859,N_29715);
or UO_72 (O_72,N_29982,N_29925);
nand UO_73 (O_73,N_29949,N_29967);
or UO_74 (O_74,N_29847,N_29743);
or UO_75 (O_75,N_29806,N_29753);
nand UO_76 (O_76,N_29750,N_29867);
and UO_77 (O_77,N_29833,N_29713);
and UO_78 (O_78,N_29821,N_29845);
xnor UO_79 (O_79,N_29919,N_29785);
nand UO_80 (O_80,N_29732,N_29932);
and UO_81 (O_81,N_29793,N_29983);
nand UO_82 (O_82,N_29958,N_29756);
or UO_83 (O_83,N_29898,N_29888);
and UO_84 (O_84,N_29841,N_29989);
and UO_85 (O_85,N_29911,N_29848);
and UO_86 (O_86,N_29964,N_29757);
nor UO_87 (O_87,N_29916,N_29794);
xor UO_88 (O_88,N_29904,N_29921);
nor UO_89 (O_89,N_29842,N_29899);
and UO_90 (O_90,N_29913,N_29961);
nor UO_91 (O_91,N_29935,N_29877);
nor UO_92 (O_92,N_29832,N_29870);
nor UO_93 (O_93,N_29885,N_29733);
nor UO_94 (O_94,N_29789,N_29766);
and UO_95 (O_95,N_29758,N_29887);
nor UO_96 (O_96,N_29968,N_29866);
nor UO_97 (O_97,N_29951,N_29943);
or UO_98 (O_98,N_29765,N_29762);
and UO_99 (O_99,N_29801,N_29731);
and UO_100 (O_100,N_29817,N_29882);
xnor UO_101 (O_101,N_29969,N_29858);
nor UO_102 (O_102,N_29926,N_29994);
nand UO_103 (O_103,N_29736,N_29718);
nand UO_104 (O_104,N_29872,N_29710);
xnor UO_105 (O_105,N_29770,N_29784);
nor UO_106 (O_106,N_29769,N_29893);
nand UO_107 (O_107,N_29830,N_29910);
and UO_108 (O_108,N_29807,N_29748);
or UO_109 (O_109,N_29721,N_29716);
or UO_110 (O_110,N_29891,N_29950);
nand UO_111 (O_111,N_29920,N_29959);
nand UO_112 (O_112,N_29997,N_29741);
xnor UO_113 (O_113,N_29928,N_29880);
nand UO_114 (O_114,N_29984,N_29896);
or UO_115 (O_115,N_29802,N_29835);
nor UO_116 (O_116,N_29760,N_29973);
xnor UO_117 (O_117,N_29838,N_29776);
and UO_118 (O_118,N_29936,N_29917);
nor UO_119 (O_119,N_29768,N_29820);
nand UO_120 (O_120,N_29751,N_29850);
and UO_121 (O_121,N_29783,N_29767);
nor UO_122 (O_122,N_29831,N_29856);
nor UO_123 (O_123,N_29884,N_29754);
and UO_124 (O_124,N_29934,N_29941);
or UO_125 (O_125,N_29978,N_29886);
and UO_126 (O_126,N_29939,N_29894);
nor UO_127 (O_127,N_29883,N_29711);
or UO_128 (O_128,N_29746,N_29970);
nor UO_129 (O_129,N_29977,N_29944);
xor UO_130 (O_130,N_29999,N_29947);
or UO_131 (O_131,N_29774,N_29962);
xor UO_132 (O_132,N_29744,N_29931);
and UO_133 (O_133,N_29735,N_29868);
xnor UO_134 (O_134,N_29791,N_29755);
nand UO_135 (O_135,N_29701,N_29818);
and UO_136 (O_136,N_29798,N_29988);
nand UO_137 (O_137,N_29745,N_29704);
nand UO_138 (O_138,N_29979,N_29772);
nor UO_139 (O_139,N_29862,N_29948);
or UO_140 (O_140,N_29903,N_29957);
or UO_141 (O_141,N_29738,N_29933);
xnor UO_142 (O_142,N_29864,N_29878);
nand UO_143 (O_143,N_29963,N_29727);
or UO_144 (O_144,N_29706,N_29824);
nand UO_145 (O_145,N_29779,N_29786);
and UO_146 (O_146,N_29908,N_29700);
and UO_147 (O_147,N_29980,N_29712);
nor UO_148 (O_148,N_29930,N_29723);
and UO_149 (O_149,N_29905,N_29863);
and UO_150 (O_150,N_29910,N_29864);
nand UO_151 (O_151,N_29963,N_29851);
xor UO_152 (O_152,N_29824,N_29841);
nand UO_153 (O_153,N_29864,N_29865);
nor UO_154 (O_154,N_29953,N_29964);
nand UO_155 (O_155,N_29799,N_29712);
nand UO_156 (O_156,N_29801,N_29717);
nor UO_157 (O_157,N_29982,N_29878);
xor UO_158 (O_158,N_29865,N_29702);
or UO_159 (O_159,N_29816,N_29969);
or UO_160 (O_160,N_29720,N_29737);
nand UO_161 (O_161,N_29846,N_29964);
nor UO_162 (O_162,N_29772,N_29711);
nand UO_163 (O_163,N_29703,N_29818);
xor UO_164 (O_164,N_29921,N_29877);
and UO_165 (O_165,N_29771,N_29765);
nand UO_166 (O_166,N_29996,N_29845);
nor UO_167 (O_167,N_29762,N_29747);
nand UO_168 (O_168,N_29720,N_29805);
nand UO_169 (O_169,N_29979,N_29751);
and UO_170 (O_170,N_29938,N_29720);
or UO_171 (O_171,N_29832,N_29849);
and UO_172 (O_172,N_29901,N_29811);
nor UO_173 (O_173,N_29919,N_29797);
nand UO_174 (O_174,N_29946,N_29706);
nand UO_175 (O_175,N_29855,N_29952);
and UO_176 (O_176,N_29863,N_29718);
nand UO_177 (O_177,N_29706,N_29935);
or UO_178 (O_178,N_29942,N_29811);
nand UO_179 (O_179,N_29947,N_29813);
or UO_180 (O_180,N_29706,N_29808);
xnor UO_181 (O_181,N_29881,N_29944);
nand UO_182 (O_182,N_29779,N_29971);
and UO_183 (O_183,N_29710,N_29740);
xnor UO_184 (O_184,N_29805,N_29922);
xor UO_185 (O_185,N_29991,N_29797);
and UO_186 (O_186,N_29914,N_29832);
xor UO_187 (O_187,N_29958,N_29745);
nand UO_188 (O_188,N_29790,N_29732);
and UO_189 (O_189,N_29945,N_29923);
or UO_190 (O_190,N_29867,N_29982);
and UO_191 (O_191,N_29918,N_29902);
nand UO_192 (O_192,N_29901,N_29840);
xnor UO_193 (O_193,N_29781,N_29941);
nor UO_194 (O_194,N_29835,N_29842);
nor UO_195 (O_195,N_29732,N_29838);
nand UO_196 (O_196,N_29870,N_29735);
nor UO_197 (O_197,N_29960,N_29865);
or UO_198 (O_198,N_29826,N_29836);
nand UO_199 (O_199,N_29804,N_29913);
and UO_200 (O_200,N_29808,N_29913);
nand UO_201 (O_201,N_29850,N_29917);
xor UO_202 (O_202,N_29850,N_29828);
or UO_203 (O_203,N_29956,N_29803);
and UO_204 (O_204,N_29806,N_29843);
or UO_205 (O_205,N_29960,N_29965);
xnor UO_206 (O_206,N_29969,N_29986);
and UO_207 (O_207,N_29969,N_29966);
nor UO_208 (O_208,N_29979,N_29854);
xor UO_209 (O_209,N_29848,N_29829);
nor UO_210 (O_210,N_29865,N_29915);
nor UO_211 (O_211,N_29807,N_29787);
or UO_212 (O_212,N_29938,N_29829);
and UO_213 (O_213,N_29860,N_29983);
nand UO_214 (O_214,N_29720,N_29804);
nand UO_215 (O_215,N_29748,N_29893);
nor UO_216 (O_216,N_29800,N_29829);
nor UO_217 (O_217,N_29705,N_29803);
nand UO_218 (O_218,N_29872,N_29824);
or UO_219 (O_219,N_29857,N_29776);
xor UO_220 (O_220,N_29874,N_29971);
or UO_221 (O_221,N_29897,N_29710);
nand UO_222 (O_222,N_29714,N_29754);
xnor UO_223 (O_223,N_29986,N_29817);
or UO_224 (O_224,N_29873,N_29949);
and UO_225 (O_225,N_29954,N_29962);
nor UO_226 (O_226,N_29949,N_29743);
xor UO_227 (O_227,N_29898,N_29771);
xnor UO_228 (O_228,N_29751,N_29897);
or UO_229 (O_229,N_29772,N_29798);
xnor UO_230 (O_230,N_29959,N_29799);
nor UO_231 (O_231,N_29827,N_29909);
or UO_232 (O_232,N_29702,N_29862);
xnor UO_233 (O_233,N_29959,N_29827);
nor UO_234 (O_234,N_29971,N_29907);
and UO_235 (O_235,N_29850,N_29841);
and UO_236 (O_236,N_29719,N_29800);
and UO_237 (O_237,N_29784,N_29974);
and UO_238 (O_238,N_29914,N_29757);
nor UO_239 (O_239,N_29774,N_29943);
nand UO_240 (O_240,N_29966,N_29818);
and UO_241 (O_241,N_29807,N_29898);
or UO_242 (O_242,N_29856,N_29938);
or UO_243 (O_243,N_29838,N_29837);
and UO_244 (O_244,N_29983,N_29934);
and UO_245 (O_245,N_29895,N_29909);
or UO_246 (O_246,N_29746,N_29932);
xnor UO_247 (O_247,N_29798,N_29991);
nor UO_248 (O_248,N_29771,N_29723);
nand UO_249 (O_249,N_29729,N_29964);
or UO_250 (O_250,N_29959,N_29923);
or UO_251 (O_251,N_29713,N_29944);
and UO_252 (O_252,N_29859,N_29737);
or UO_253 (O_253,N_29758,N_29946);
nor UO_254 (O_254,N_29718,N_29724);
xor UO_255 (O_255,N_29797,N_29743);
xnor UO_256 (O_256,N_29908,N_29933);
or UO_257 (O_257,N_29901,N_29822);
nor UO_258 (O_258,N_29825,N_29885);
or UO_259 (O_259,N_29742,N_29834);
or UO_260 (O_260,N_29754,N_29713);
and UO_261 (O_261,N_29843,N_29893);
or UO_262 (O_262,N_29803,N_29724);
nor UO_263 (O_263,N_29869,N_29835);
nor UO_264 (O_264,N_29712,N_29769);
or UO_265 (O_265,N_29931,N_29898);
xnor UO_266 (O_266,N_29811,N_29890);
nand UO_267 (O_267,N_29796,N_29702);
and UO_268 (O_268,N_29782,N_29847);
and UO_269 (O_269,N_29922,N_29957);
nand UO_270 (O_270,N_29938,N_29790);
nor UO_271 (O_271,N_29837,N_29908);
nand UO_272 (O_272,N_29747,N_29756);
and UO_273 (O_273,N_29909,N_29704);
or UO_274 (O_274,N_29916,N_29906);
or UO_275 (O_275,N_29727,N_29772);
and UO_276 (O_276,N_29898,N_29784);
and UO_277 (O_277,N_29936,N_29723);
and UO_278 (O_278,N_29779,N_29877);
and UO_279 (O_279,N_29799,N_29851);
nand UO_280 (O_280,N_29744,N_29846);
xnor UO_281 (O_281,N_29770,N_29911);
or UO_282 (O_282,N_29723,N_29923);
or UO_283 (O_283,N_29748,N_29931);
nor UO_284 (O_284,N_29995,N_29857);
or UO_285 (O_285,N_29836,N_29868);
nor UO_286 (O_286,N_29949,N_29963);
nor UO_287 (O_287,N_29806,N_29924);
or UO_288 (O_288,N_29880,N_29715);
and UO_289 (O_289,N_29835,N_29959);
xnor UO_290 (O_290,N_29750,N_29943);
or UO_291 (O_291,N_29871,N_29924);
xor UO_292 (O_292,N_29707,N_29706);
or UO_293 (O_293,N_29922,N_29983);
nand UO_294 (O_294,N_29915,N_29965);
xnor UO_295 (O_295,N_29954,N_29830);
xor UO_296 (O_296,N_29930,N_29901);
nand UO_297 (O_297,N_29721,N_29762);
and UO_298 (O_298,N_29714,N_29824);
or UO_299 (O_299,N_29975,N_29933);
and UO_300 (O_300,N_29983,N_29735);
or UO_301 (O_301,N_29784,N_29748);
nor UO_302 (O_302,N_29941,N_29925);
xnor UO_303 (O_303,N_29899,N_29700);
or UO_304 (O_304,N_29738,N_29767);
nor UO_305 (O_305,N_29792,N_29797);
xnor UO_306 (O_306,N_29741,N_29853);
nor UO_307 (O_307,N_29964,N_29950);
nand UO_308 (O_308,N_29887,N_29924);
nor UO_309 (O_309,N_29995,N_29741);
nand UO_310 (O_310,N_29985,N_29804);
nand UO_311 (O_311,N_29964,N_29949);
and UO_312 (O_312,N_29725,N_29904);
or UO_313 (O_313,N_29949,N_29780);
and UO_314 (O_314,N_29786,N_29794);
or UO_315 (O_315,N_29731,N_29806);
and UO_316 (O_316,N_29955,N_29760);
and UO_317 (O_317,N_29755,N_29838);
xnor UO_318 (O_318,N_29700,N_29788);
or UO_319 (O_319,N_29899,N_29949);
and UO_320 (O_320,N_29839,N_29764);
xnor UO_321 (O_321,N_29709,N_29944);
xor UO_322 (O_322,N_29742,N_29718);
xnor UO_323 (O_323,N_29888,N_29885);
or UO_324 (O_324,N_29701,N_29997);
nand UO_325 (O_325,N_29972,N_29918);
xor UO_326 (O_326,N_29899,N_29881);
nand UO_327 (O_327,N_29950,N_29795);
xnor UO_328 (O_328,N_29889,N_29814);
or UO_329 (O_329,N_29894,N_29702);
or UO_330 (O_330,N_29930,N_29987);
nand UO_331 (O_331,N_29709,N_29742);
xnor UO_332 (O_332,N_29855,N_29715);
or UO_333 (O_333,N_29748,N_29801);
nand UO_334 (O_334,N_29775,N_29742);
nand UO_335 (O_335,N_29727,N_29923);
xor UO_336 (O_336,N_29966,N_29974);
and UO_337 (O_337,N_29908,N_29731);
or UO_338 (O_338,N_29960,N_29760);
nand UO_339 (O_339,N_29743,N_29700);
and UO_340 (O_340,N_29772,N_29739);
and UO_341 (O_341,N_29876,N_29721);
nor UO_342 (O_342,N_29982,N_29938);
xnor UO_343 (O_343,N_29768,N_29862);
or UO_344 (O_344,N_29881,N_29840);
nand UO_345 (O_345,N_29808,N_29711);
and UO_346 (O_346,N_29937,N_29768);
or UO_347 (O_347,N_29844,N_29729);
and UO_348 (O_348,N_29969,N_29844);
nor UO_349 (O_349,N_29844,N_29856);
nand UO_350 (O_350,N_29773,N_29936);
and UO_351 (O_351,N_29724,N_29917);
nand UO_352 (O_352,N_29789,N_29849);
nand UO_353 (O_353,N_29916,N_29746);
nand UO_354 (O_354,N_29982,N_29798);
xnor UO_355 (O_355,N_29700,N_29749);
nor UO_356 (O_356,N_29953,N_29808);
nand UO_357 (O_357,N_29859,N_29738);
nand UO_358 (O_358,N_29850,N_29782);
nand UO_359 (O_359,N_29926,N_29752);
xor UO_360 (O_360,N_29814,N_29758);
nand UO_361 (O_361,N_29965,N_29996);
or UO_362 (O_362,N_29805,N_29738);
nor UO_363 (O_363,N_29999,N_29983);
nor UO_364 (O_364,N_29823,N_29850);
and UO_365 (O_365,N_29884,N_29928);
nand UO_366 (O_366,N_29917,N_29772);
or UO_367 (O_367,N_29799,N_29850);
xor UO_368 (O_368,N_29848,N_29826);
and UO_369 (O_369,N_29967,N_29979);
or UO_370 (O_370,N_29820,N_29981);
or UO_371 (O_371,N_29833,N_29776);
or UO_372 (O_372,N_29735,N_29816);
xor UO_373 (O_373,N_29722,N_29951);
nor UO_374 (O_374,N_29881,N_29872);
xnor UO_375 (O_375,N_29991,N_29770);
or UO_376 (O_376,N_29960,N_29851);
xnor UO_377 (O_377,N_29749,N_29927);
nand UO_378 (O_378,N_29957,N_29738);
or UO_379 (O_379,N_29886,N_29831);
xnor UO_380 (O_380,N_29725,N_29850);
or UO_381 (O_381,N_29859,N_29825);
xnor UO_382 (O_382,N_29992,N_29770);
nand UO_383 (O_383,N_29754,N_29798);
nand UO_384 (O_384,N_29862,N_29993);
or UO_385 (O_385,N_29774,N_29729);
and UO_386 (O_386,N_29891,N_29930);
and UO_387 (O_387,N_29785,N_29730);
and UO_388 (O_388,N_29851,N_29894);
and UO_389 (O_389,N_29761,N_29918);
or UO_390 (O_390,N_29970,N_29860);
and UO_391 (O_391,N_29746,N_29926);
nand UO_392 (O_392,N_29717,N_29870);
or UO_393 (O_393,N_29729,N_29745);
nand UO_394 (O_394,N_29999,N_29708);
and UO_395 (O_395,N_29920,N_29743);
nand UO_396 (O_396,N_29864,N_29950);
xor UO_397 (O_397,N_29713,N_29859);
nor UO_398 (O_398,N_29855,N_29784);
or UO_399 (O_399,N_29739,N_29849);
xnor UO_400 (O_400,N_29837,N_29975);
nor UO_401 (O_401,N_29713,N_29985);
nand UO_402 (O_402,N_29816,N_29768);
nand UO_403 (O_403,N_29868,N_29716);
xor UO_404 (O_404,N_29918,N_29963);
and UO_405 (O_405,N_29973,N_29766);
or UO_406 (O_406,N_29722,N_29982);
or UO_407 (O_407,N_29883,N_29947);
and UO_408 (O_408,N_29937,N_29853);
or UO_409 (O_409,N_29957,N_29962);
or UO_410 (O_410,N_29771,N_29984);
nor UO_411 (O_411,N_29859,N_29932);
nor UO_412 (O_412,N_29961,N_29989);
nor UO_413 (O_413,N_29725,N_29755);
or UO_414 (O_414,N_29741,N_29921);
nor UO_415 (O_415,N_29972,N_29901);
nor UO_416 (O_416,N_29751,N_29844);
xor UO_417 (O_417,N_29703,N_29964);
nand UO_418 (O_418,N_29706,N_29918);
and UO_419 (O_419,N_29863,N_29806);
nor UO_420 (O_420,N_29875,N_29787);
nor UO_421 (O_421,N_29728,N_29963);
or UO_422 (O_422,N_29879,N_29716);
xor UO_423 (O_423,N_29837,N_29771);
and UO_424 (O_424,N_29959,N_29765);
nand UO_425 (O_425,N_29721,N_29954);
xnor UO_426 (O_426,N_29922,N_29958);
xor UO_427 (O_427,N_29824,N_29910);
xor UO_428 (O_428,N_29708,N_29850);
xor UO_429 (O_429,N_29927,N_29831);
or UO_430 (O_430,N_29739,N_29993);
nand UO_431 (O_431,N_29723,N_29888);
or UO_432 (O_432,N_29965,N_29718);
or UO_433 (O_433,N_29904,N_29734);
xor UO_434 (O_434,N_29978,N_29925);
or UO_435 (O_435,N_29819,N_29905);
xor UO_436 (O_436,N_29814,N_29852);
nor UO_437 (O_437,N_29737,N_29767);
xor UO_438 (O_438,N_29876,N_29909);
nand UO_439 (O_439,N_29956,N_29985);
nand UO_440 (O_440,N_29912,N_29984);
nor UO_441 (O_441,N_29972,N_29898);
and UO_442 (O_442,N_29713,N_29903);
and UO_443 (O_443,N_29894,N_29823);
nand UO_444 (O_444,N_29755,N_29704);
nor UO_445 (O_445,N_29939,N_29742);
and UO_446 (O_446,N_29929,N_29911);
or UO_447 (O_447,N_29959,N_29728);
nand UO_448 (O_448,N_29702,N_29721);
nand UO_449 (O_449,N_29860,N_29871);
or UO_450 (O_450,N_29872,N_29985);
or UO_451 (O_451,N_29950,N_29888);
and UO_452 (O_452,N_29939,N_29778);
and UO_453 (O_453,N_29817,N_29738);
xor UO_454 (O_454,N_29780,N_29901);
nor UO_455 (O_455,N_29884,N_29828);
and UO_456 (O_456,N_29936,N_29790);
nand UO_457 (O_457,N_29854,N_29900);
nor UO_458 (O_458,N_29890,N_29846);
nand UO_459 (O_459,N_29722,N_29834);
nand UO_460 (O_460,N_29949,N_29894);
nor UO_461 (O_461,N_29784,N_29963);
and UO_462 (O_462,N_29730,N_29745);
nor UO_463 (O_463,N_29809,N_29994);
nand UO_464 (O_464,N_29751,N_29930);
or UO_465 (O_465,N_29828,N_29896);
nand UO_466 (O_466,N_29829,N_29851);
nand UO_467 (O_467,N_29843,N_29816);
and UO_468 (O_468,N_29880,N_29917);
or UO_469 (O_469,N_29902,N_29753);
xnor UO_470 (O_470,N_29995,N_29805);
nor UO_471 (O_471,N_29993,N_29723);
and UO_472 (O_472,N_29976,N_29864);
nor UO_473 (O_473,N_29935,N_29900);
nor UO_474 (O_474,N_29863,N_29931);
xor UO_475 (O_475,N_29770,N_29874);
nor UO_476 (O_476,N_29866,N_29801);
and UO_477 (O_477,N_29902,N_29946);
nor UO_478 (O_478,N_29914,N_29962);
or UO_479 (O_479,N_29815,N_29808);
nand UO_480 (O_480,N_29952,N_29787);
nor UO_481 (O_481,N_29800,N_29723);
nand UO_482 (O_482,N_29936,N_29823);
nor UO_483 (O_483,N_29767,N_29815);
nor UO_484 (O_484,N_29993,N_29972);
or UO_485 (O_485,N_29739,N_29831);
xor UO_486 (O_486,N_29731,N_29932);
nand UO_487 (O_487,N_29761,N_29981);
and UO_488 (O_488,N_29903,N_29769);
nand UO_489 (O_489,N_29910,N_29972);
and UO_490 (O_490,N_29767,N_29861);
xnor UO_491 (O_491,N_29862,N_29786);
or UO_492 (O_492,N_29845,N_29781);
and UO_493 (O_493,N_29794,N_29839);
xor UO_494 (O_494,N_29784,N_29844);
nor UO_495 (O_495,N_29856,N_29893);
nand UO_496 (O_496,N_29933,N_29767);
and UO_497 (O_497,N_29863,N_29756);
and UO_498 (O_498,N_29814,N_29753);
nor UO_499 (O_499,N_29701,N_29942);
and UO_500 (O_500,N_29776,N_29920);
or UO_501 (O_501,N_29989,N_29982);
and UO_502 (O_502,N_29796,N_29727);
and UO_503 (O_503,N_29763,N_29968);
nor UO_504 (O_504,N_29915,N_29878);
nand UO_505 (O_505,N_29786,N_29821);
and UO_506 (O_506,N_29939,N_29979);
nand UO_507 (O_507,N_29871,N_29982);
nand UO_508 (O_508,N_29899,N_29797);
xnor UO_509 (O_509,N_29790,N_29793);
nand UO_510 (O_510,N_29725,N_29713);
or UO_511 (O_511,N_29765,N_29953);
nand UO_512 (O_512,N_29926,N_29934);
nor UO_513 (O_513,N_29924,N_29991);
xor UO_514 (O_514,N_29847,N_29899);
nand UO_515 (O_515,N_29726,N_29717);
or UO_516 (O_516,N_29987,N_29746);
nand UO_517 (O_517,N_29894,N_29791);
and UO_518 (O_518,N_29961,N_29971);
xnor UO_519 (O_519,N_29824,N_29859);
nor UO_520 (O_520,N_29809,N_29946);
nor UO_521 (O_521,N_29869,N_29840);
and UO_522 (O_522,N_29736,N_29705);
and UO_523 (O_523,N_29815,N_29989);
nor UO_524 (O_524,N_29917,N_29973);
xor UO_525 (O_525,N_29882,N_29951);
and UO_526 (O_526,N_29987,N_29884);
or UO_527 (O_527,N_29890,N_29704);
and UO_528 (O_528,N_29992,N_29885);
or UO_529 (O_529,N_29922,N_29762);
or UO_530 (O_530,N_29925,N_29922);
or UO_531 (O_531,N_29722,N_29845);
nor UO_532 (O_532,N_29860,N_29945);
and UO_533 (O_533,N_29817,N_29866);
xor UO_534 (O_534,N_29918,N_29710);
and UO_535 (O_535,N_29800,N_29983);
and UO_536 (O_536,N_29814,N_29733);
xor UO_537 (O_537,N_29928,N_29904);
and UO_538 (O_538,N_29879,N_29853);
or UO_539 (O_539,N_29782,N_29895);
xor UO_540 (O_540,N_29932,N_29974);
xnor UO_541 (O_541,N_29945,N_29758);
xor UO_542 (O_542,N_29966,N_29931);
or UO_543 (O_543,N_29849,N_29761);
nor UO_544 (O_544,N_29971,N_29904);
and UO_545 (O_545,N_29936,N_29754);
xor UO_546 (O_546,N_29787,N_29763);
and UO_547 (O_547,N_29702,N_29858);
xor UO_548 (O_548,N_29709,N_29998);
and UO_549 (O_549,N_29900,N_29911);
and UO_550 (O_550,N_29966,N_29716);
xnor UO_551 (O_551,N_29992,N_29704);
nand UO_552 (O_552,N_29952,N_29926);
nand UO_553 (O_553,N_29726,N_29939);
and UO_554 (O_554,N_29911,N_29919);
and UO_555 (O_555,N_29908,N_29962);
nand UO_556 (O_556,N_29842,N_29828);
nor UO_557 (O_557,N_29870,N_29953);
and UO_558 (O_558,N_29910,N_29839);
nand UO_559 (O_559,N_29734,N_29801);
nand UO_560 (O_560,N_29824,N_29845);
or UO_561 (O_561,N_29912,N_29927);
or UO_562 (O_562,N_29852,N_29805);
xor UO_563 (O_563,N_29807,N_29703);
and UO_564 (O_564,N_29714,N_29794);
xor UO_565 (O_565,N_29941,N_29782);
nand UO_566 (O_566,N_29954,N_29750);
xnor UO_567 (O_567,N_29895,N_29808);
nand UO_568 (O_568,N_29705,N_29970);
nand UO_569 (O_569,N_29866,N_29763);
nor UO_570 (O_570,N_29709,N_29884);
and UO_571 (O_571,N_29899,N_29798);
or UO_572 (O_572,N_29796,N_29830);
nand UO_573 (O_573,N_29910,N_29846);
and UO_574 (O_574,N_29812,N_29904);
and UO_575 (O_575,N_29922,N_29888);
xnor UO_576 (O_576,N_29814,N_29887);
nor UO_577 (O_577,N_29716,N_29887);
nor UO_578 (O_578,N_29782,N_29770);
and UO_579 (O_579,N_29885,N_29828);
nor UO_580 (O_580,N_29747,N_29826);
xor UO_581 (O_581,N_29801,N_29882);
nor UO_582 (O_582,N_29768,N_29956);
nor UO_583 (O_583,N_29852,N_29794);
nor UO_584 (O_584,N_29937,N_29736);
xnor UO_585 (O_585,N_29806,N_29751);
nor UO_586 (O_586,N_29832,N_29955);
and UO_587 (O_587,N_29847,N_29823);
xor UO_588 (O_588,N_29959,N_29966);
nand UO_589 (O_589,N_29928,N_29977);
nand UO_590 (O_590,N_29841,N_29934);
xnor UO_591 (O_591,N_29842,N_29719);
nand UO_592 (O_592,N_29847,N_29962);
nand UO_593 (O_593,N_29798,N_29940);
or UO_594 (O_594,N_29744,N_29924);
and UO_595 (O_595,N_29777,N_29809);
and UO_596 (O_596,N_29991,N_29990);
and UO_597 (O_597,N_29711,N_29753);
nor UO_598 (O_598,N_29872,N_29772);
xnor UO_599 (O_599,N_29796,N_29774);
or UO_600 (O_600,N_29961,N_29856);
and UO_601 (O_601,N_29745,N_29896);
and UO_602 (O_602,N_29760,N_29941);
nor UO_603 (O_603,N_29821,N_29992);
nand UO_604 (O_604,N_29796,N_29869);
or UO_605 (O_605,N_29768,N_29866);
nor UO_606 (O_606,N_29754,N_29872);
xnor UO_607 (O_607,N_29928,N_29860);
nor UO_608 (O_608,N_29949,N_29723);
xnor UO_609 (O_609,N_29839,N_29755);
xor UO_610 (O_610,N_29732,N_29826);
or UO_611 (O_611,N_29877,N_29712);
nor UO_612 (O_612,N_29721,N_29833);
and UO_613 (O_613,N_29748,N_29958);
or UO_614 (O_614,N_29763,N_29857);
and UO_615 (O_615,N_29886,N_29945);
or UO_616 (O_616,N_29941,N_29788);
xor UO_617 (O_617,N_29960,N_29773);
xnor UO_618 (O_618,N_29810,N_29902);
nor UO_619 (O_619,N_29922,N_29809);
and UO_620 (O_620,N_29792,N_29938);
nor UO_621 (O_621,N_29713,N_29870);
xor UO_622 (O_622,N_29765,N_29750);
and UO_623 (O_623,N_29745,N_29850);
xor UO_624 (O_624,N_29829,N_29831);
xor UO_625 (O_625,N_29845,N_29815);
nor UO_626 (O_626,N_29970,N_29923);
xnor UO_627 (O_627,N_29996,N_29827);
nand UO_628 (O_628,N_29878,N_29792);
or UO_629 (O_629,N_29807,N_29969);
nor UO_630 (O_630,N_29894,N_29778);
xnor UO_631 (O_631,N_29748,N_29831);
xor UO_632 (O_632,N_29875,N_29928);
and UO_633 (O_633,N_29870,N_29879);
nor UO_634 (O_634,N_29989,N_29916);
or UO_635 (O_635,N_29975,N_29791);
and UO_636 (O_636,N_29741,N_29994);
or UO_637 (O_637,N_29932,N_29733);
and UO_638 (O_638,N_29819,N_29750);
xor UO_639 (O_639,N_29959,N_29727);
or UO_640 (O_640,N_29709,N_29948);
nand UO_641 (O_641,N_29834,N_29945);
nand UO_642 (O_642,N_29718,N_29789);
xnor UO_643 (O_643,N_29818,N_29773);
and UO_644 (O_644,N_29958,N_29927);
nor UO_645 (O_645,N_29763,N_29802);
nand UO_646 (O_646,N_29854,N_29834);
nor UO_647 (O_647,N_29750,N_29871);
xor UO_648 (O_648,N_29707,N_29888);
xor UO_649 (O_649,N_29958,N_29706);
or UO_650 (O_650,N_29843,N_29936);
nor UO_651 (O_651,N_29844,N_29749);
and UO_652 (O_652,N_29955,N_29792);
nor UO_653 (O_653,N_29891,N_29815);
and UO_654 (O_654,N_29987,N_29843);
and UO_655 (O_655,N_29740,N_29876);
nor UO_656 (O_656,N_29868,N_29911);
and UO_657 (O_657,N_29750,N_29917);
and UO_658 (O_658,N_29881,N_29852);
nand UO_659 (O_659,N_29960,N_29815);
and UO_660 (O_660,N_29847,N_29905);
nor UO_661 (O_661,N_29705,N_29913);
nand UO_662 (O_662,N_29821,N_29972);
nor UO_663 (O_663,N_29836,N_29776);
nand UO_664 (O_664,N_29988,N_29743);
nand UO_665 (O_665,N_29768,N_29738);
xnor UO_666 (O_666,N_29846,N_29860);
and UO_667 (O_667,N_29897,N_29838);
and UO_668 (O_668,N_29816,N_29886);
and UO_669 (O_669,N_29822,N_29999);
nor UO_670 (O_670,N_29729,N_29955);
and UO_671 (O_671,N_29715,N_29731);
or UO_672 (O_672,N_29919,N_29749);
or UO_673 (O_673,N_29966,N_29903);
xnor UO_674 (O_674,N_29858,N_29837);
nand UO_675 (O_675,N_29781,N_29843);
and UO_676 (O_676,N_29881,N_29968);
nor UO_677 (O_677,N_29897,N_29969);
or UO_678 (O_678,N_29841,N_29795);
xnor UO_679 (O_679,N_29805,N_29727);
and UO_680 (O_680,N_29792,N_29753);
xor UO_681 (O_681,N_29788,N_29717);
xor UO_682 (O_682,N_29853,N_29735);
xnor UO_683 (O_683,N_29807,N_29762);
nand UO_684 (O_684,N_29862,N_29765);
and UO_685 (O_685,N_29725,N_29917);
or UO_686 (O_686,N_29848,N_29822);
or UO_687 (O_687,N_29827,N_29935);
nand UO_688 (O_688,N_29774,N_29903);
and UO_689 (O_689,N_29935,N_29707);
xor UO_690 (O_690,N_29860,N_29765);
or UO_691 (O_691,N_29883,N_29792);
and UO_692 (O_692,N_29700,N_29895);
nor UO_693 (O_693,N_29962,N_29832);
or UO_694 (O_694,N_29869,N_29762);
xnor UO_695 (O_695,N_29859,N_29928);
or UO_696 (O_696,N_29930,N_29988);
or UO_697 (O_697,N_29922,N_29835);
xor UO_698 (O_698,N_29915,N_29939);
and UO_699 (O_699,N_29990,N_29904);
or UO_700 (O_700,N_29865,N_29982);
xnor UO_701 (O_701,N_29872,N_29745);
and UO_702 (O_702,N_29855,N_29866);
nand UO_703 (O_703,N_29890,N_29899);
and UO_704 (O_704,N_29705,N_29825);
nor UO_705 (O_705,N_29785,N_29953);
xor UO_706 (O_706,N_29750,N_29913);
nand UO_707 (O_707,N_29831,N_29762);
nor UO_708 (O_708,N_29746,N_29869);
xnor UO_709 (O_709,N_29826,N_29959);
and UO_710 (O_710,N_29890,N_29738);
and UO_711 (O_711,N_29840,N_29968);
or UO_712 (O_712,N_29953,N_29706);
nor UO_713 (O_713,N_29814,N_29948);
or UO_714 (O_714,N_29774,N_29776);
nand UO_715 (O_715,N_29958,N_29734);
or UO_716 (O_716,N_29884,N_29904);
nand UO_717 (O_717,N_29777,N_29733);
or UO_718 (O_718,N_29929,N_29775);
or UO_719 (O_719,N_29725,N_29825);
and UO_720 (O_720,N_29713,N_29973);
nor UO_721 (O_721,N_29884,N_29708);
nor UO_722 (O_722,N_29761,N_29915);
and UO_723 (O_723,N_29916,N_29869);
and UO_724 (O_724,N_29885,N_29796);
and UO_725 (O_725,N_29815,N_29980);
and UO_726 (O_726,N_29995,N_29860);
nand UO_727 (O_727,N_29714,N_29892);
xor UO_728 (O_728,N_29983,N_29911);
nand UO_729 (O_729,N_29828,N_29892);
and UO_730 (O_730,N_29867,N_29991);
nand UO_731 (O_731,N_29777,N_29914);
xnor UO_732 (O_732,N_29712,N_29771);
xnor UO_733 (O_733,N_29799,N_29764);
xor UO_734 (O_734,N_29944,N_29806);
nand UO_735 (O_735,N_29754,N_29779);
xor UO_736 (O_736,N_29789,N_29801);
and UO_737 (O_737,N_29866,N_29822);
xor UO_738 (O_738,N_29822,N_29833);
nand UO_739 (O_739,N_29812,N_29982);
and UO_740 (O_740,N_29926,N_29965);
nor UO_741 (O_741,N_29777,N_29845);
and UO_742 (O_742,N_29775,N_29719);
and UO_743 (O_743,N_29794,N_29806);
and UO_744 (O_744,N_29845,N_29756);
xnor UO_745 (O_745,N_29855,N_29832);
nand UO_746 (O_746,N_29878,N_29810);
nand UO_747 (O_747,N_29823,N_29726);
nor UO_748 (O_748,N_29835,N_29846);
xor UO_749 (O_749,N_29754,N_29841);
nor UO_750 (O_750,N_29883,N_29721);
nor UO_751 (O_751,N_29838,N_29745);
and UO_752 (O_752,N_29837,N_29860);
and UO_753 (O_753,N_29705,N_29725);
nand UO_754 (O_754,N_29823,N_29734);
xor UO_755 (O_755,N_29939,N_29855);
nand UO_756 (O_756,N_29904,N_29930);
and UO_757 (O_757,N_29855,N_29986);
nor UO_758 (O_758,N_29976,N_29790);
or UO_759 (O_759,N_29717,N_29909);
and UO_760 (O_760,N_29703,N_29885);
nand UO_761 (O_761,N_29884,N_29787);
nor UO_762 (O_762,N_29706,N_29919);
nand UO_763 (O_763,N_29973,N_29740);
or UO_764 (O_764,N_29982,N_29963);
nor UO_765 (O_765,N_29969,N_29843);
nor UO_766 (O_766,N_29943,N_29906);
or UO_767 (O_767,N_29705,N_29928);
or UO_768 (O_768,N_29716,N_29717);
xnor UO_769 (O_769,N_29801,N_29837);
xor UO_770 (O_770,N_29926,N_29841);
xor UO_771 (O_771,N_29939,N_29843);
xor UO_772 (O_772,N_29836,N_29739);
nand UO_773 (O_773,N_29967,N_29990);
nor UO_774 (O_774,N_29808,N_29942);
and UO_775 (O_775,N_29939,N_29715);
or UO_776 (O_776,N_29713,N_29921);
nand UO_777 (O_777,N_29956,N_29709);
and UO_778 (O_778,N_29935,N_29777);
xor UO_779 (O_779,N_29768,N_29758);
and UO_780 (O_780,N_29868,N_29753);
xnor UO_781 (O_781,N_29988,N_29896);
nor UO_782 (O_782,N_29891,N_29966);
nand UO_783 (O_783,N_29897,N_29888);
nor UO_784 (O_784,N_29939,N_29926);
or UO_785 (O_785,N_29872,N_29807);
nand UO_786 (O_786,N_29933,N_29719);
and UO_787 (O_787,N_29730,N_29894);
or UO_788 (O_788,N_29929,N_29846);
xor UO_789 (O_789,N_29710,N_29816);
xnor UO_790 (O_790,N_29835,N_29810);
or UO_791 (O_791,N_29932,N_29939);
xor UO_792 (O_792,N_29873,N_29905);
xnor UO_793 (O_793,N_29835,N_29717);
nor UO_794 (O_794,N_29790,N_29726);
or UO_795 (O_795,N_29791,N_29727);
nor UO_796 (O_796,N_29834,N_29713);
xor UO_797 (O_797,N_29856,N_29930);
and UO_798 (O_798,N_29957,N_29730);
nand UO_799 (O_799,N_29971,N_29797);
nor UO_800 (O_800,N_29864,N_29970);
and UO_801 (O_801,N_29769,N_29899);
or UO_802 (O_802,N_29907,N_29788);
nor UO_803 (O_803,N_29701,N_29965);
or UO_804 (O_804,N_29893,N_29905);
nand UO_805 (O_805,N_29856,N_29975);
xor UO_806 (O_806,N_29805,N_29854);
xor UO_807 (O_807,N_29953,N_29984);
or UO_808 (O_808,N_29869,N_29722);
and UO_809 (O_809,N_29892,N_29877);
and UO_810 (O_810,N_29973,N_29990);
xor UO_811 (O_811,N_29873,N_29886);
nor UO_812 (O_812,N_29824,N_29978);
or UO_813 (O_813,N_29988,N_29738);
or UO_814 (O_814,N_29962,N_29886);
and UO_815 (O_815,N_29887,N_29986);
xor UO_816 (O_816,N_29845,N_29710);
xor UO_817 (O_817,N_29908,N_29981);
or UO_818 (O_818,N_29943,N_29752);
nand UO_819 (O_819,N_29825,N_29903);
xnor UO_820 (O_820,N_29744,N_29768);
xnor UO_821 (O_821,N_29750,N_29961);
or UO_822 (O_822,N_29798,N_29832);
nand UO_823 (O_823,N_29973,N_29886);
nor UO_824 (O_824,N_29980,N_29764);
nor UO_825 (O_825,N_29885,N_29739);
nand UO_826 (O_826,N_29862,N_29958);
and UO_827 (O_827,N_29860,N_29783);
nand UO_828 (O_828,N_29788,N_29849);
xnor UO_829 (O_829,N_29735,N_29955);
xnor UO_830 (O_830,N_29769,N_29896);
and UO_831 (O_831,N_29908,N_29831);
nand UO_832 (O_832,N_29837,N_29722);
nand UO_833 (O_833,N_29998,N_29832);
nor UO_834 (O_834,N_29845,N_29884);
xnor UO_835 (O_835,N_29930,N_29969);
or UO_836 (O_836,N_29729,N_29986);
nand UO_837 (O_837,N_29911,N_29851);
or UO_838 (O_838,N_29956,N_29837);
xnor UO_839 (O_839,N_29941,N_29989);
xnor UO_840 (O_840,N_29881,N_29965);
nor UO_841 (O_841,N_29808,N_29874);
nor UO_842 (O_842,N_29875,N_29757);
nor UO_843 (O_843,N_29906,N_29905);
and UO_844 (O_844,N_29872,N_29808);
and UO_845 (O_845,N_29710,N_29933);
or UO_846 (O_846,N_29950,N_29765);
nand UO_847 (O_847,N_29704,N_29941);
nand UO_848 (O_848,N_29755,N_29746);
and UO_849 (O_849,N_29760,N_29842);
nand UO_850 (O_850,N_29757,N_29938);
nor UO_851 (O_851,N_29876,N_29855);
or UO_852 (O_852,N_29704,N_29702);
nand UO_853 (O_853,N_29861,N_29869);
nor UO_854 (O_854,N_29929,N_29879);
xnor UO_855 (O_855,N_29939,N_29739);
xnor UO_856 (O_856,N_29842,N_29860);
nor UO_857 (O_857,N_29801,N_29966);
or UO_858 (O_858,N_29970,N_29972);
nand UO_859 (O_859,N_29730,N_29760);
nand UO_860 (O_860,N_29749,N_29869);
nand UO_861 (O_861,N_29794,N_29886);
nor UO_862 (O_862,N_29743,N_29718);
xor UO_863 (O_863,N_29840,N_29858);
nor UO_864 (O_864,N_29883,N_29892);
or UO_865 (O_865,N_29720,N_29732);
nor UO_866 (O_866,N_29977,N_29750);
xnor UO_867 (O_867,N_29852,N_29964);
and UO_868 (O_868,N_29740,N_29893);
and UO_869 (O_869,N_29968,N_29835);
or UO_870 (O_870,N_29923,N_29754);
xor UO_871 (O_871,N_29930,N_29836);
or UO_872 (O_872,N_29706,N_29774);
xor UO_873 (O_873,N_29919,N_29732);
or UO_874 (O_874,N_29839,N_29938);
nand UO_875 (O_875,N_29772,N_29705);
xnor UO_876 (O_876,N_29984,N_29762);
or UO_877 (O_877,N_29986,N_29992);
nor UO_878 (O_878,N_29895,N_29870);
or UO_879 (O_879,N_29805,N_29740);
xnor UO_880 (O_880,N_29789,N_29954);
nand UO_881 (O_881,N_29910,N_29744);
xor UO_882 (O_882,N_29718,N_29915);
and UO_883 (O_883,N_29753,N_29828);
nand UO_884 (O_884,N_29870,N_29728);
xnor UO_885 (O_885,N_29932,N_29934);
and UO_886 (O_886,N_29986,N_29916);
xor UO_887 (O_887,N_29833,N_29795);
xnor UO_888 (O_888,N_29826,N_29738);
nor UO_889 (O_889,N_29767,N_29752);
xnor UO_890 (O_890,N_29832,N_29781);
nor UO_891 (O_891,N_29904,N_29807);
or UO_892 (O_892,N_29761,N_29945);
nand UO_893 (O_893,N_29768,N_29970);
and UO_894 (O_894,N_29787,N_29826);
nor UO_895 (O_895,N_29991,N_29756);
and UO_896 (O_896,N_29830,N_29927);
or UO_897 (O_897,N_29933,N_29712);
xnor UO_898 (O_898,N_29860,N_29888);
xnor UO_899 (O_899,N_29795,N_29943);
xnor UO_900 (O_900,N_29978,N_29703);
xor UO_901 (O_901,N_29848,N_29878);
or UO_902 (O_902,N_29868,N_29828);
and UO_903 (O_903,N_29843,N_29779);
nand UO_904 (O_904,N_29777,N_29987);
or UO_905 (O_905,N_29766,N_29787);
xnor UO_906 (O_906,N_29933,N_29941);
or UO_907 (O_907,N_29857,N_29915);
or UO_908 (O_908,N_29712,N_29792);
and UO_909 (O_909,N_29784,N_29740);
nor UO_910 (O_910,N_29835,N_29905);
xor UO_911 (O_911,N_29801,N_29957);
xnor UO_912 (O_912,N_29945,N_29741);
xnor UO_913 (O_913,N_29796,N_29823);
xnor UO_914 (O_914,N_29726,N_29852);
and UO_915 (O_915,N_29905,N_29752);
and UO_916 (O_916,N_29922,N_29967);
xnor UO_917 (O_917,N_29732,N_29727);
xnor UO_918 (O_918,N_29854,N_29947);
or UO_919 (O_919,N_29817,N_29903);
and UO_920 (O_920,N_29904,N_29979);
nand UO_921 (O_921,N_29870,N_29947);
and UO_922 (O_922,N_29971,N_29762);
nand UO_923 (O_923,N_29990,N_29844);
and UO_924 (O_924,N_29980,N_29906);
and UO_925 (O_925,N_29735,N_29884);
nand UO_926 (O_926,N_29853,N_29999);
nor UO_927 (O_927,N_29738,N_29719);
nor UO_928 (O_928,N_29847,N_29857);
xnor UO_929 (O_929,N_29927,N_29993);
nand UO_930 (O_930,N_29776,N_29932);
and UO_931 (O_931,N_29711,N_29826);
and UO_932 (O_932,N_29758,N_29782);
xnor UO_933 (O_933,N_29785,N_29946);
xor UO_934 (O_934,N_29980,N_29778);
nand UO_935 (O_935,N_29878,N_29714);
or UO_936 (O_936,N_29700,N_29764);
nor UO_937 (O_937,N_29989,N_29929);
nand UO_938 (O_938,N_29956,N_29765);
nand UO_939 (O_939,N_29728,N_29702);
and UO_940 (O_940,N_29757,N_29908);
or UO_941 (O_941,N_29702,N_29713);
and UO_942 (O_942,N_29829,N_29833);
and UO_943 (O_943,N_29795,N_29981);
nor UO_944 (O_944,N_29817,N_29849);
nor UO_945 (O_945,N_29827,N_29901);
nand UO_946 (O_946,N_29905,N_29854);
or UO_947 (O_947,N_29926,N_29724);
and UO_948 (O_948,N_29721,N_29809);
or UO_949 (O_949,N_29717,N_29744);
xor UO_950 (O_950,N_29950,N_29799);
nand UO_951 (O_951,N_29779,N_29790);
xor UO_952 (O_952,N_29914,N_29947);
nand UO_953 (O_953,N_29831,N_29809);
xor UO_954 (O_954,N_29820,N_29879);
nor UO_955 (O_955,N_29949,N_29736);
xor UO_956 (O_956,N_29759,N_29726);
and UO_957 (O_957,N_29792,N_29819);
nand UO_958 (O_958,N_29940,N_29764);
or UO_959 (O_959,N_29842,N_29804);
xnor UO_960 (O_960,N_29909,N_29812);
nor UO_961 (O_961,N_29716,N_29777);
xor UO_962 (O_962,N_29713,N_29762);
or UO_963 (O_963,N_29744,N_29913);
or UO_964 (O_964,N_29878,N_29828);
or UO_965 (O_965,N_29957,N_29782);
or UO_966 (O_966,N_29710,N_29889);
nor UO_967 (O_967,N_29890,N_29776);
nor UO_968 (O_968,N_29795,N_29848);
nor UO_969 (O_969,N_29771,N_29849);
nand UO_970 (O_970,N_29940,N_29931);
nand UO_971 (O_971,N_29806,N_29835);
and UO_972 (O_972,N_29918,N_29958);
or UO_973 (O_973,N_29851,N_29709);
xor UO_974 (O_974,N_29978,N_29997);
nor UO_975 (O_975,N_29926,N_29726);
nor UO_976 (O_976,N_29760,N_29927);
or UO_977 (O_977,N_29722,N_29880);
nor UO_978 (O_978,N_29821,N_29721);
xor UO_979 (O_979,N_29948,N_29740);
and UO_980 (O_980,N_29900,N_29951);
nand UO_981 (O_981,N_29916,N_29909);
nor UO_982 (O_982,N_29786,N_29774);
or UO_983 (O_983,N_29784,N_29700);
and UO_984 (O_984,N_29740,N_29915);
nand UO_985 (O_985,N_29950,N_29990);
nor UO_986 (O_986,N_29991,N_29747);
or UO_987 (O_987,N_29789,N_29907);
and UO_988 (O_988,N_29956,N_29976);
nand UO_989 (O_989,N_29790,N_29846);
xor UO_990 (O_990,N_29897,N_29759);
xor UO_991 (O_991,N_29930,N_29962);
xor UO_992 (O_992,N_29751,N_29767);
or UO_993 (O_993,N_29826,N_29958);
or UO_994 (O_994,N_29781,N_29809);
or UO_995 (O_995,N_29959,N_29784);
xor UO_996 (O_996,N_29801,N_29744);
and UO_997 (O_997,N_29752,N_29993);
and UO_998 (O_998,N_29949,N_29992);
xnor UO_999 (O_999,N_29708,N_29949);
nor UO_1000 (O_1000,N_29812,N_29808);
nand UO_1001 (O_1001,N_29756,N_29775);
or UO_1002 (O_1002,N_29965,N_29980);
xor UO_1003 (O_1003,N_29823,N_29769);
nor UO_1004 (O_1004,N_29735,N_29760);
or UO_1005 (O_1005,N_29723,N_29795);
nand UO_1006 (O_1006,N_29744,N_29751);
or UO_1007 (O_1007,N_29810,N_29910);
and UO_1008 (O_1008,N_29722,N_29752);
nor UO_1009 (O_1009,N_29770,N_29835);
or UO_1010 (O_1010,N_29776,N_29921);
xor UO_1011 (O_1011,N_29814,N_29924);
nand UO_1012 (O_1012,N_29763,N_29706);
and UO_1013 (O_1013,N_29870,N_29827);
nand UO_1014 (O_1014,N_29932,N_29954);
nor UO_1015 (O_1015,N_29780,N_29906);
nor UO_1016 (O_1016,N_29877,N_29747);
and UO_1017 (O_1017,N_29824,N_29940);
and UO_1018 (O_1018,N_29856,N_29715);
and UO_1019 (O_1019,N_29838,N_29885);
nor UO_1020 (O_1020,N_29753,N_29723);
nand UO_1021 (O_1021,N_29883,N_29822);
nor UO_1022 (O_1022,N_29795,N_29963);
nor UO_1023 (O_1023,N_29713,N_29847);
or UO_1024 (O_1024,N_29832,N_29980);
nand UO_1025 (O_1025,N_29746,N_29876);
or UO_1026 (O_1026,N_29827,N_29900);
nand UO_1027 (O_1027,N_29986,N_29795);
and UO_1028 (O_1028,N_29710,N_29886);
xnor UO_1029 (O_1029,N_29803,N_29908);
nand UO_1030 (O_1030,N_29803,N_29945);
xor UO_1031 (O_1031,N_29710,N_29810);
nor UO_1032 (O_1032,N_29891,N_29784);
nor UO_1033 (O_1033,N_29758,N_29875);
nand UO_1034 (O_1034,N_29972,N_29743);
nor UO_1035 (O_1035,N_29885,N_29715);
nand UO_1036 (O_1036,N_29824,N_29790);
nand UO_1037 (O_1037,N_29724,N_29774);
or UO_1038 (O_1038,N_29714,N_29817);
nand UO_1039 (O_1039,N_29824,N_29948);
or UO_1040 (O_1040,N_29814,N_29941);
nand UO_1041 (O_1041,N_29956,N_29907);
nand UO_1042 (O_1042,N_29730,N_29821);
xnor UO_1043 (O_1043,N_29722,N_29769);
nor UO_1044 (O_1044,N_29731,N_29736);
and UO_1045 (O_1045,N_29713,N_29818);
xnor UO_1046 (O_1046,N_29894,N_29743);
nand UO_1047 (O_1047,N_29816,N_29864);
and UO_1048 (O_1048,N_29935,N_29800);
and UO_1049 (O_1049,N_29789,N_29717);
nor UO_1050 (O_1050,N_29711,N_29888);
or UO_1051 (O_1051,N_29968,N_29806);
nand UO_1052 (O_1052,N_29954,N_29924);
nand UO_1053 (O_1053,N_29884,N_29714);
nor UO_1054 (O_1054,N_29831,N_29721);
nor UO_1055 (O_1055,N_29747,N_29786);
nand UO_1056 (O_1056,N_29702,N_29785);
nor UO_1057 (O_1057,N_29769,N_29819);
nor UO_1058 (O_1058,N_29936,N_29866);
nand UO_1059 (O_1059,N_29878,N_29782);
nor UO_1060 (O_1060,N_29914,N_29831);
nand UO_1061 (O_1061,N_29970,N_29926);
xor UO_1062 (O_1062,N_29965,N_29826);
or UO_1063 (O_1063,N_29740,N_29939);
nor UO_1064 (O_1064,N_29940,N_29956);
xnor UO_1065 (O_1065,N_29820,N_29730);
nor UO_1066 (O_1066,N_29748,N_29701);
xor UO_1067 (O_1067,N_29878,N_29818);
nor UO_1068 (O_1068,N_29711,N_29897);
nor UO_1069 (O_1069,N_29805,N_29840);
nand UO_1070 (O_1070,N_29838,N_29955);
or UO_1071 (O_1071,N_29748,N_29981);
or UO_1072 (O_1072,N_29781,N_29769);
nor UO_1073 (O_1073,N_29992,N_29909);
nand UO_1074 (O_1074,N_29922,N_29952);
nor UO_1075 (O_1075,N_29836,N_29900);
nand UO_1076 (O_1076,N_29747,N_29764);
and UO_1077 (O_1077,N_29884,N_29806);
nand UO_1078 (O_1078,N_29735,N_29728);
and UO_1079 (O_1079,N_29831,N_29862);
xnor UO_1080 (O_1080,N_29795,N_29956);
or UO_1081 (O_1081,N_29848,N_29714);
nor UO_1082 (O_1082,N_29793,N_29714);
nand UO_1083 (O_1083,N_29930,N_29833);
or UO_1084 (O_1084,N_29713,N_29963);
or UO_1085 (O_1085,N_29757,N_29904);
nand UO_1086 (O_1086,N_29983,N_29994);
and UO_1087 (O_1087,N_29728,N_29824);
nand UO_1088 (O_1088,N_29956,N_29743);
nor UO_1089 (O_1089,N_29766,N_29925);
nor UO_1090 (O_1090,N_29926,N_29705);
or UO_1091 (O_1091,N_29992,N_29787);
nand UO_1092 (O_1092,N_29948,N_29920);
nand UO_1093 (O_1093,N_29727,N_29974);
or UO_1094 (O_1094,N_29734,N_29708);
and UO_1095 (O_1095,N_29996,N_29734);
and UO_1096 (O_1096,N_29891,N_29976);
nand UO_1097 (O_1097,N_29819,N_29749);
and UO_1098 (O_1098,N_29798,N_29781);
xor UO_1099 (O_1099,N_29961,N_29776);
or UO_1100 (O_1100,N_29770,N_29790);
xor UO_1101 (O_1101,N_29925,N_29995);
or UO_1102 (O_1102,N_29868,N_29783);
and UO_1103 (O_1103,N_29990,N_29715);
and UO_1104 (O_1104,N_29740,N_29824);
nor UO_1105 (O_1105,N_29857,N_29709);
nand UO_1106 (O_1106,N_29951,N_29779);
and UO_1107 (O_1107,N_29763,N_29790);
and UO_1108 (O_1108,N_29783,N_29740);
or UO_1109 (O_1109,N_29826,N_29942);
and UO_1110 (O_1110,N_29871,N_29915);
nor UO_1111 (O_1111,N_29873,N_29740);
xor UO_1112 (O_1112,N_29773,N_29783);
and UO_1113 (O_1113,N_29720,N_29807);
or UO_1114 (O_1114,N_29991,N_29914);
nor UO_1115 (O_1115,N_29941,N_29995);
nor UO_1116 (O_1116,N_29943,N_29825);
xor UO_1117 (O_1117,N_29884,N_29717);
nand UO_1118 (O_1118,N_29770,N_29780);
or UO_1119 (O_1119,N_29913,N_29713);
nand UO_1120 (O_1120,N_29741,N_29935);
nand UO_1121 (O_1121,N_29751,N_29706);
nor UO_1122 (O_1122,N_29758,N_29965);
and UO_1123 (O_1123,N_29970,N_29736);
and UO_1124 (O_1124,N_29968,N_29838);
xor UO_1125 (O_1125,N_29968,N_29780);
xor UO_1126 (O_1126,N_29849,N_29823);
or UO_1127 (O_1127,N_29949,N_29719);
or UO_1128 (O_1128,N_29769,N_29705);
nor UO_1129 (O_1129,N_29945,N_29878);
and UO_1130 (O_1130,N_29899,N_29863);
nor UO_1131 (O_1131,N_29944,N_29757);
and UO_1132 (O_1132,N_29718,N_29706);
nor UO_1133 (O_1133,N_29743,N_29940);
nor UO_1134 (O_1134,N_29734,N_29851);
nand UO_1135 (O_1135,N_29705,N_29711);
xor UO_1136 (O_1136,N_29754,N_29956);
or UO_1137 (O_1137,N_29870,N_29719);
nor UO_1138 (O_1138,N_29940,N_29983);
or UO_1139 (O_1139,N_29841,N_29767);
and UO_1140 (O_1140,N_29806,N_29986);
nor UO_1141 (O_1141,N_29807,N_29881);
xnor UO_1142 (O_1142,N_29933,N_29724);
nand UO_1143 (O_1143,N_29977,N_29844);
nand UO_1144 (O_1144,N_29727,N_29891);
and UO_1145 (O_1145,N_29836,N_29856);
nor UO_1146 (O_1146,N_29821,N_29963);
and UO_1147 (O_1147,N_29841,N_29966);
or UO_1148 (O_1148,N_29785,N_29990);
nand UO_1149 (O_1149,N_29760,N_29995);
xor UO_1150 (O_1150,N_29998,N_29725);
and UO_1151 (O_1151,N_29988,N_29828);
nand UO_1152 (O_1152,N_29882,N_29986);
nor UO_1153 (O_1153,N_29861,N_29800);
nor UO_1154 (O_1154,N_29951,N_29851);
nor UO_1155 (O_1155,N_29936,N_29709);
xor UO_1156 (O_1156,N_29885,N_29868);
nand UO_1157 (O_1157,N_29794,N_29796);
nand UO_1158 (O_1158,N_29773,N_29839);
nor UO_1159 (O_1159,N_29728,N_29792);
nor UO_1160 (O_1160,N_29810,N_29879);
nand UO_1161 (O_1161,N_29946,N_29949);
xor UO_1162 (O_1162,N_29911,N_29877);
and UO_1163 (O_1163,N_29932,N_29737);
or UO_1164 (O_1164,N_29765,N_29889);
nand UO_1165 (O_1165,N_29869,N_29704);
nand UO_1166 (O_1166,N_29802,N_29920);
xor UO_1167 (O_1167,N_29842,N_29870);
or UO_1168 (O_1168,N_29951,N_29794);
or UO_1169 (O_1169,N_29846,N_29947);
nand UO_1170 (O_1170,N_29904,N_29941);
and UO_1171 (O_1171,N_29888,N_29790);
and UO_1172 (O_1172,N_29917,N_29798);
nor UO_1173 (O_1173,N_29999,N_29820);
nand UO_1174 (O_1174,N_29701,N_29988);
nand UO_1175 (O_1175,N_29924,N_29874);
or UO_1176 (O_1176,N_29709,N_29976);
nand UO_1177 (O_1177,N_29958,N_29995);
nor UO_1178 (O_1178,N_29701,N_29919);
nor UO_1179 (O_1179,N_29891,N_29802);
nand UO_1180 (O_1180,N_29777,N_29782);
nor UO_1181 (O_1181,N_29813,N_29931);
or UO_1182 (O_1182,N_29870,N_29709);
nand UO_1183 (O_1183,N_29946,N_29867);
nor UO_1184 (O_1184,N_29777,N_29979);
and UO_1185 (O_1185,N_29742,N_29723);
nor UO_1186 (O_1186,N_29774,N_29787);
or UO_1187 (O_1187,N_29786,N_29925);
xnor UO_1188 (O_1188,N_29741,N_29887);
nor UO_1189 (O_1189,N_29902,N_29988);
and UO_1190 (O_1190,N_29817,N_29700);
xnor UO_1191 (O_1191,N_29711,N_29780);
and UO_1192 (O_1192,N_29971,N_29836);
and UO_1193 (O_1193,N_29734,N_29713);
xnor UO_1194 (O_1194,N_29770,N_29904);
nand UO_1195 (O_1195,N_29773,N_29897);
nor UO_1196 (O_1196,N_29861,N_29741);
nor UO_1197 (O_1197,N_29752,N_29725);
nor UO_1198 (O_1198,N_29946,N_29910);
nand UO_1199 (O_1199,N_29968,N_29872);
or UO_1200 (O_1200,N_29739,N_29890);
xnor UO_1201 (O_1201,N_29760,N_29732);
or UO_1202 (O_1202,N_29830,N_29709);
and UO_1203 (O_1203,N_29975,N_29981);
xor UO_1204 (O_1204,N_29898,N_29956);
and UO_1205 (O_1205,N_29960,N_29727);
nand UO_1206 (O_1206,N_29896,N_29857);
nand UO_1207 (O_1207,N_29950,N_29921);
and UO_1208 (O_1208,N_29886,N_29756);
or UO_1209 (O_1209,N_29818,N_29731);
nand UO_1210 (O_1210,N_29733,N_29739);
xnor UO_1211 (O_1211,N_29790,N_29787);
xor UO_1212 (O_1212,N_29984,N_29729);
nand UO_1213 (O_1213,N_29815,N_29786);
or UO_1214 (O_1214,N_29892,N_29784);
nor UO_1215 (O_1215,N_29851,N_29849);
nand UO_1216 (O_1216,N_29938,N_29732);
or UO_1217 (O_1217,N_29713,N_29748);
or UO_1218 (O_1218,N_29737,N_29880);
xor UO_1219 (O_1219,N_29884,N_29901);
nor UO_1220 (O_1220,N_29768,N_29881);
or UO_1221 (O_1221,N_29861,N_29877);
nor UO_1222 (O_1222,N_29894,N_29776);
and UO_1223 (O_1223,N_29881,N_29827);
nand UO_1224 (O_1224,N_29902,N_29862);
nor UO_1225 (O_1225,N_29741,N_29850);
or UO_1226 (O_1226,N_29769,N_29996);
or UO_1227 (O_1227,N_29771,N_29817);
and UO_1228 (O_1228,N_29770,N_29916);
and UO_1229 (O_1229,N_29851,N_29731);
and UO_1230 (O_1230,N_29757,N_29747);
nand UO_1231 (O_1231,N_29796,N_29933);
nor UO_1232 (O_1232,N_29968,N_29722);
nor UO_1233 (O_1233,N_29873,N_29728);
or UO_1234 (O_1234,N_29829,N_29715);
nand UO_1235 (O_1235,N_29830,N_29969);
nor UO_1236 (O_1236,N_29868,N_29898);
and UO_1237 (O_1237,N_29793,N_29892);
or UO_1238 (O_1238,N_29770,N_29986);
nand UO_1239 (O_1239,N_29860,N_29857);
nand UO_1240 (O_1240,N_29908,N_29946);
nor UO_1241 (O_1241,N_29786,N_29716);
nor UO_1242 (O_1242,N_29758,N_29730);
and UO_1243 (O_1243,N_29826,N_29860);
or UO_1244 (O_1244,N_29752,N_29768);
nand UO_1245 (O_1245,N_29782,N_29837);
nand UO_1246 (O_1246,N_29964,N_29716);
nand UO_1247 (O_1247,N_29866,N_29760);
nor UO_1248 (O_1248,N_29756,N_29772);
nand UO_1249 (O_1249,N_29801,N_29701);
nor UO_1250 (O_1250,N_29836,N_29767);
xnor UO_1251 (O_1251,N_29896,N_29778);
xnor UO_1252 (O_1252,N_29725,N_29800);
and UO_1253 (O_1253,N_29791,N_29986);
or UO_1254 (O_1254,N_29763,N_29874);
and UO_1255 (O_1255,N_29817,N_29780);
nand UO_1256 (O_1256,N_29999,N_29810);
or UO_1257 (O_1257,N_29945,N_29929);
xor UO_1258 (O_1258,N_29756,N_29732);
nor UO_1259 (O_1259,N_29822,N_29903);
or UO_1260 (O_1260,N_29909,N_29901);
and UO_1261 (O_1261,N_29935,N_29978);
and UO_1262 (O_1262,N_29918,N_29876);
and UO_1263 (O_1263,N_29762,N_29708);
xor UO_1264 (O_1264,N_29823,N_29968);
nor UO_1265 (O_1265,N_29749,N_29909);
nor UO_1266 (O_1266,N_29700,N_29969);
xnor UO_1267 (O_1267,N_29763,N_29986);
or UO_1268 (O_1268,N_29876,N_29765);
xnor UO_1269 (O_1269,N_29903,N_29782);
and UO_1270 (O_1270,N_29913,N_29747);
xnor UO_1271 (O_1271,N_29986,N_29836);
nor UO_1272 (O_1272,N_29930,N_29765);
or UO_1273 (O_1273,N_29895,N_29715);
nand UO_1274 (O_1274,N_29877,N_29808);
nor UO_1275 (O_1275,N_29783,N_29746);
nand UO_1276 (O_1276,N_29940,N_29820);
xor UO_1277 (O_1277,N_29933,N_29952);
and UO_1278 (O_1278,N_29837,N_29856);
and UO_1279 (O_1279,N_29740,N_29874);
and UO_1280 (O_1280,N_29720,N_29772);
nor UO_1281 (O_1281,N_29825,N_29842);
nor UO_1282 (O_1282,N_29927,N_29872);
xnor UO_1283 (O_1283,N_29899,N_29818);
xnor UO_1284 (O_1284,N_29923,N_29763);
nand UO_1285 (O_1285,N_29702,N_29746);
nor UO_1286 (O_1286,N_29709,N_29972);
xor UO_1287 (O_1287,N_29913,N_29959);
and UO_1288 (O_1288,N_29722,N_29956);
xnor UO_1289 (O_1289,N_29753,N_29705);
and UO_1290 (O_1290,N_29853,N_29839);
nand UO_1291 (O_1291,N_29842,N_29993);
or UO_1292 (O_1292,N_29971,N_29716);
xnor UO_1293 (O_1293,N_29859,N_29754);
xor UO_1294 (O_1294,N_29756,N_29921);
or UO_1295 (O_1295,N_29891,N_29805);
xor UO_1296 (O_1296,N_29735,N_29716);
xor UO_1297 (O_1297,N_29745,N_29786);
or UO_1298 (O_1298,N_29706,N_29800);
or UO_1299 (O_1299,N_29877,N_29780);
nor UO_1300 (O_1300,N_29950,N_29968);
nor UO_1301 (O_1301,N_29905,N_29946);
xor UO_1302 (O_1302,N_29868,N_29889);
and UO_1303 (O_1303,N_29764,N_29786);
and UO_1304 (O_1304,N_29880,N_29794);
or UO_1305 (O_1305,N_29752,N_29927);
and UO_1306 (O_1306,N_29916,N_29947);
nor UO_1307 (O_1307,N_29963,N_29735);
xnor UO_1308 (O_1308,N_29822,N_29892);
nor UO_1309 (O_1309,N_29882,N_29878);
and UO_1310 (O_1310,N_29763,N_29735);
nand UO_1311 (O_1311,N_29757,N_29826);
xnor UO_1312 (O_1312,N_29830,N_29730);
and UO_1313 (O_1313,N_29700,N_29761);
and UO_1314 (O_1314,N_29993,N_29857);
xnor UO_1315 (O_1315,N_29924,N_29873);
and UO_1316 (O_1316,N_29952,N_29917);
and UO_1317 (O_1317,N_29749,N_29722);
or UO_1318 (O_1318,N_29963,N_29995);
or UO_1319 (O_1319,N_29951,N_29889);
and UO_1320 (O_1320,N_29775,N_29846);
xnor UO_1321 (O_1321,N_29706,N_29813);
and UO_1322 (O_1322,N_29931,N_29916);
xor UO_1323 (O_1323,N_29991,N_29846);
and UO_1324 (O_1324,N_29962,N_29880);
and UO_1325 (O_1325,N_29775,N_29816);
or UO_1326 (O_1326,N_29968,N_29815);
or UO_1327 (O_1327,N_29939,N_29866);
nor UO_1328 (O_1328,N_29915,N_29826);
or UO_1329 (O_1329,N_29834,N_29928);
xor UO_1330 (O_1330,N_29743,N_29980);
or UO_1331 (O_1331,N_29769,N_29876);
or UO_1332 (O_1332,N_29860,N_29940);
xnor UO_1333 (O_1333,N_29979,N_29722);
nand UO_1334 (O_1334,N_29813,N_29879);
or UO_1335 (O_1335,N_29839,N_29856);
nor UO_1336 (O_1336,N_29977,N_29918);
nor UO_1337 (O_1337,N_29772,N_29839);
or UO_1338 (O_1338,N_29933,N_29939);
and UO_1339 (O_1339,N_29826,N_29872);
nor UO_1340 (O_1340,N_29702,N_29827);
or UO_1341 (O_1341,N_29795,N_29869);
and UO_1342 (O_1342,N_29922,N_29866);
or UO_1343 (O_1343,N_29906,N_29850);
and UO_1344 (O_1344,N_29768,N_29869);
nand UO_1345 (O_1345,N_29759,N_29994);
and UO_1346 (O_1346,N_29989,N_29773);
xor UO_1347 (O_1347,N_29932,N_29729);
and UO_1348 (O_1348,N_29849,N_29806);
nor UO_1349 (O_1349,N_29973,N_29893);
or UO_1350 (O_1350,N_29959,N_29770);
xor UO_1351 (O_1351,N_29875,N_29975);
or UO_1352 (O_1352,N_29827,N_29719);
or UO_1353 (O_1353,N_29993,N_29848);
nor UO_1354 (O_1354,N_29891,N_29956);
or UO_1355 (O_1355,N_29947,N_29811);
or UO_1356 (O_1356,N_29825,N_29837);
xor UO_1357 (O_1357,N_29928,N_29732);
nand UO_1358 (O_1358,N_29728,N_29919);
and UO_1359 (O_1359,N_29923,N_29905);
nor UO_1360 (O_1360,N_29979,N_29819);
and UO_1361 (O_1361,N_29798,N_29826);
nor UO_1362 (O_1362,N_29843,N_29913);
nand UO_1363 (O_1363,N_29991,N_29746);
nand UO_1364 (O_1364,N_29825,N_29756);
and UO_1365 (O_1365,N_29795,N_29719);
nand UO_1366 (O_1366,N_29814,N_29918);
xnor UO_1367 (O_1367,N_29885,N_29723);
nor UO_1368 (O_1368,N_29991,N_29862);
and UO_1369 (O_1369,N_29864,N_29943);
or UO_1370 (O_1370,N_29979,N_29902);
and UO_1371 (O_1371,N_29889,N_29914);
xnor UO_1372 (O_1372,N_29983,N_29736);
xor UO_1373 (O_1373,N_29848,N_29895);
nand UO_1374 (O_1374,N_29760,N_29867);
nor UO_1375 (O_1375,N_29705,N_29981);
xor UO_1376 (O_1376,N_29709,N_29719);
or UO_1377 (O_1377,N_29731,N_29897);
nor UO_1378 (O_1378,N_29736,N_29809);
nand UO_1379 (O_1379,N_29964,N_29764);
and UO_1380 (O_1380,N_29975,N_29832);
nand UO_1381 (O_1381,N_29762,N_29888);
xnor UO_1382 (O_1382,N_29818,N_29748);
or UO_1383 (O_1383,N_29886,N_29728);
nand UO_1384 (O_1384,N_29971,N_29841);
nand UO_1385 (O_1385,N_29921,N_29801);
xnor UO_1386 (O_1386,N_29911,N_29880);
and UO_1387 (O_1387,N_29987,N_29762);
and UO_1388 (O_1388,N_29859,N_29794);
nor UO_1389 (O_1389,N_29981,N_29879);
or UO_1390 (O_1390,N_29842,N_29906);
nor UO_1391 (O_1391,N_29824,N_29801);
nand UO_1392 (O_1392,N_29843,N_29865);
or UO_1393 (O_1393,N_29787,N_29854);
and UO_1394 (O_1394,N_29816,N_29797);
nor UO_1395 (O_1395,N_29786,N_29884);
nand UO_1396 (O_1396,N_29795,N_29749);
nand UO_1397 (O_1397,N_29864,N_29703);
or UO_1398 (O_1398,N_29977,N_29921);
nor UO_1399 (O_1399,N_29750,N_29805);
or UO_1400 (O_1400,N_29749,N_29777);
and UO_1401 (O_1401,N_29790,N_29948);
nor UO_1402 (O_1402,N_29824,N_29704);
nor UO_1403 (O_1403,N_29746,N_29824);
xor UO_1404 (O_1404,N_29813,N_29848);
or UO_1405 (O_1405,N_29759,N_29968);
or UO_1406 (O_1406,N_29936,N_29910);
xor UO_1407 (O_1407,N_29704,N_29746);
nand UO_1408 (O_1408,N_29792,N_29864);
and UO_1409 (O_1409,N_29926,N_29825);
nor UO_1410 (O_1410,N_29745,N_29837);
or UO_1411 (O_1411,N_29719,N_29930);
and UO_1412 (O_1412,N_29901,N_29967);
and UO_1413 (O_1413,N_29708,N_29806);
xor UO_1414 (O_1414,N_29880,N_29977);
and UO_1415 (O_1415,N_29714,N_29917);
xnor UO_1416 (O_1416,N_29766,N_29790);
nand UO_1417 (O_1417,N_29994,N_29800);
xor UO_1418 (O_1418,N_29968,N_29909);
nor UO_1419 (O_1419,N_29793,N_29913);
or UO_1420 (O_1420,N_29780,N_29904);
xnor UO_1421 (O_1421,N_29796,N_29732);
xor UO_1422 (O_1422,N_29831,N_29965);
and UO_1423 (O_1423,N_29864,N_29769);
and UO_1424 (O_1424,N_29762,N_29749);
and UO_1425 (O_1425,N_29851,N_29830);
nand UO_1426 (O_1426,N_29883,N_29835);
nor UO_1427 (O_1427,N_29758,N_29901);
and UO_1428 (O_1428,N_29766,N_29823);
nand UO_1429 (O_1429,N_29909,N_29728);
xor UO_1430 (O_1430,N_29831,N_29868);
or UO_1431 (O_1431,N_29708,N_29902);
xor UO_1432 (O_1432,N_29809,N_29755);
and UO_1433 (O_1433,N_29827,N_29837);
xor UO_1434 (O_1434,N_29914,N_29934);
and UO_1435 (O_1435,N_29749,N_29908);
xor UO_1436 (O_1436,N_29905,N_29953);
nor UO_1437 (O_1437,N_29979,N_29708);
nor UO_1438 (O_1438,N_29974,N_29701);
or UO_1439 (O_1439,N_29828,N_29879);
or UO_1440 (O_1440,N_29846,N_29968);
nand UO_1441 (O_1441,N_29915,N_29936);
nand UO_1442 (O_1442,N_29990,N_29908);
or UO_1443 (O_1443,N_29721,N_29863);
and UO_1444 (O_1444,N_29842,N_29994);
nor UO_1445 (O_1445,N_29714,N_29888);
xor UO_1446 (O_1446,N_29866,N_29907);
nor UO_1447 (O_1447,N_29723,N_29754);
nor UO_1448 (O_1448,N_29744,N_29878);
and UO_1449 (O_1449,N_29837,N_29971);
nand UO_1450 (O_1450,N_29794,N_29910);
nor UO_1451 (O_1451,N_29776,N_29949);
nand UO_1452 (O_1452,N_29718,N_29770);
and UO_1453 (O_1453,N_29721,N_29705);
nand UO_1454 (O_1454,N_29770,N_29909);
or UO_1455 (O_1455,N_29762,N_29808);
and UO_1456 (O_1456,N_29846,N_29831);
and UO_1457 (O_1457,N_29999,N_29881);
nor UO_1458 (O_1458,N_29963,N_29793);
nor UO_1459 (O_1459,N_29788,N_29766);
or UO_1460 (O_1460,N_29738,N_29797);
xnor UO_1461 (O_1461,N_29876,N_29947);
nor UO_1462 (O_1462,N_29722,N_29893);
or UO_1463 (O_1463,N_29784,N_29929);
nand UO_1464 (O_1464,N_29890,N_29877);
or UO_1465 (O_1465,N_29975,N_29799);
and UO_1466 (O_1466,N_29978,N_29733);
nand UO_1467 (O_1467,N_29899,N_29768);
and UO_1468 (O_1468,N_29803,N_29957);
nor UO_1469 (O_1469,N_29737,N_29875);
or UO_1470 (O_1470,N_29775,N_29798);
nand UO_1471 (O_1471,N_29723,N_29935);
or UO_1472 (O_1472,N_29984,N_29872);
or UO_1473 (O_1473,N_29704,N_29881);
xor UO_1474 (O_1474,N_29889,N_29907);
nand UO_1475 (O_1475,N_29816,N_29936);
nand UO_1476 (O_1476,N_29986,N_29957);
and UO_1477 (O_1477,N_29827,N_29942);
xnor UO_1478 (O_1478,N_29846,N_29782);
or UO_1479 (O_1479,N_29840,N_29712);
and UO_1480 (O_1480,N_29753,N_29858);
and UO_1481 (O_1481,N_29752,N_29729);
and UO_1482 (O_1482,N_29810,N_29829);
or UO_1483 (O_1483,N_29862,N_29912);
or UO_1484 (O_1484,N_29954,N_29831);
nand UO_1485 (O_1485,N_29820,N_29714);
or UO_1486 (O_1486,N_29977,N_29812);
nand UO_1487 (O_1487,N_29916,N_29994);
nor UO_1488 (O_1488,N_29912,N_29932);
and UO_1489 (O_1489,N_29926,N_29992);
nand UO_1490 (O_1490,N_29830,N_29722);
xnor UO_1491 (O_1491,N_29991,N_29865);
and UO_1492 (O_1492,N_29799,N_29730);
nand UO_1493 (O_1493,N_29988,N_29816);
nand UO_1494 (O_1494,N_29939,N_29948);
xor UO_1495 (O_1495,N_29848,N_29734);
xor UO_1496 (O_1496,N_29757,N_29729);
xor UO_1497 (O_1497,N_29745,N_29816);
nand UO_1498 (O_1498,N_29706,N_29756);
or UO_1499 (O_1499,N_29831,N_29756);
and UO_1500 (O_1500,N_29978,N_29714);
nand UO_1501 (O_1501,N_29899,N_29988);
nor UO_1502 (O_1502,N_29841,N_29838);
and UO_1503 (O_1503,N_29903,N_29792);
nand UO_1504 (O_1504,N_29801,N_29912);
nand UO_1505 (O_1505,N_29849,N_29784);
nor UO_1506 (O_1506,N_29823,N_29783);
and UO_1507 (O_1507,N_29873,N_29917);
nand UO_1508 (O_1508,N_29751,N_29869);
nor UO_1509 (O_1509,N_29917,N_29747);
nor UO_1510 (O_1510,N_29825,N_29784);
nor UO_1511 (O_1511,N_29791,N_29729);
or UO_1512 (O_1512,N_29720,N_29878);
and UO_1513 (O_1513,N_29875,N_29723);
nor UO_1514 (O_1514,N_29935,N_29791);
and UO_1515 (O_1515,N_29749,N_29813);
and UO_1516 (O_1516,N_29737,N_29804);
xor UO_1517 (O_1517,N_29983,N_29924);
nor UO_1518 (O_1518,N_29949,N_29969);
and UO_1519 (O_1519,N_29947,N_29759);
or UO_1520 (O_1520,N_29981,N_29922);
or UO_1521 (O_1521,N_29705,N_29785);
or UO_1522 (O_1522,N_29954,N_29868);
xor UO_1523 (O_1523,N_29718,N_29925);
nor UO_1524 (O_1524,N_29760,N_29833);
xnor UO_1525 (O_1525,N_29825,N_29940);
nand UO_1526 (O_1526,N_29905,N_29840);
nor UO_1527 (O_1527,N_29858,N_29730);
and UO_1528 (O_1528,N_29925,N_29737);
nor UO_1529 (O_1529,N_29733,N_29951);
nand UO_1530 (O_1530,N_29889,N_29815);
nor UO_1531 (O_1531,N_29934,N_29985);
or UO_1532 (O_1532,N_29727,N_29953);
and UO_1533 (O_1533,N_29770,N_29994);
xnor UO_1534 (O_1534,N_29847,N_29863);
and UO_1535 (O_1535,N_29915,N_29963);
nor UO_1536 (O_1536,N_29796,N_29767);
xnor UO_1537 (O_1537,N_29807,N_29951);
nor UO_1538 (O_1538,N_29793,N_29857);
nor UO_1539 (O_1539,N_29931,N_29743);
xnor UO_1540 (O_1540,N_29950,N_29725);
or UO_1541 (O_1541,N_29819,N_29975);
or UO_1542 (O_1542,N_29774,N_29895);
and UO_1543 (O_1543,N_29991,N_29912);
or UO_1544 (O_1544,N_29716,N_29943);
nand UO_1545 (O_1545,N_29905,N_29848);
xor UO_1546 (O_1546,N_29826,N_29782);
nor UO_1547 (O_1547,N_29909,N_29711);
nor UO_1548 (O_1548,N_29849,N_29868);
or UO_1549 (O_1549,N_29860,N_29911);
nor UO_1550 (O_1550,N_29869,N_29744);
nor UO_1551 (O_1551,N_29778,N_29987);
or UO_1552 (O_1552,N_29855,N_29738);
or UO_1553 (O_1553,N_29786,N_29890);
and UO_1554 (O_1554,N_29915,N_29913);
nand UO_1555 (O_1555,N_29868,N_29764);
and UO_1556 (O_1556,N_29850,N_29960);
nand UO_1557 (O_1557,N_29741,N_29928);
and UO_1558 (O_1558,N_29914,N_29764);
nor UO_1559 (O_1559,N_29981,N_29735);
or UO_1560 (O_1560,N_29720,N_29783);
nor UO_1561 (O_1561,N_29833,N_29887);
nand UO_1562 (O_1562,N_29745,N_29794);
or UO_1563 (O_1563,N_29898,N_29985);
and UO_1564 (O_1564,N_29701,N_29761);
nor UO_1565 (O_1565,N_29877,N_29939);
nor UO_1566 (O_1566,N_29732,N_29782);
and UO_1567 (O_1567,N_29722,N_29744);
or UO_1568 (O_1568,N_29706,N_29817);
nand UO_1569 (O_1569,N_29936,N_29733);
or UO_1570 (O_1570,N_29954,N_29956);
xnor UO_1571 (O_1571,N_29984,N_29925);
and UO_1572 (O_1572,N_29984,N_29930);
or UO_1573 (O_1573,N_29709,N_29765);
and UO_1574 (O_1574,N_29795,N_29765);
nand UO_1575 (O_1575,N_29838,N_29864);
nor UO_1576 (O_1576,N_29716,N_29795);
and UO_1577 (O_1577,N_29828,N_29748);
xor UO_1578 (O_1578,N_29811,N_29728);
nand UO_1579 (O_1579,N_29986,N_29914);
xor UO_1580 (O_1580,N_29724,N_29934);
and UO_1581 (O_1581,N_29831,N_29951);
nor UO_1582 (O_1582,N_29798,N_29812);
nand UO_1583 (O_1583,N_29720,N_29779);
or UO_1584 (O_1584,N_29741,N_29871);
xor UO_1585 (O_1585,N_29824,N_29938);
or UO_1586 (O_1586,N_29872,N_29875);
xnor UO_1587 (O_1587,N_29889,N_29711);
and UO_1588 (O_1588,N_29970,N_29912);
or UO_1589 (O_1589,N_29869,N_29872);
nor UO_1590 (O_1590,N_29960,N_29882);
and UO_1591 (O_1591,N_29888,N_29960);
nand UO_1592 (O_1592,N_29952,N_29887);
and UO_1593 (O_1593,N_29907,N_29880);
xor UO_1594 (O_1594,N_29978,N_29838);
xnor UO_1595 (O_1595,N_29978,N_29949);
xnor UO_1596 (O_1596,N_29710,N_29795);
and UO_1597 (O_1597,N_29794,N_29749);
or UO_1598 (O_1598,N_29778,N_29820);
nor UO_1599 (O_1599,N_29816,N_29742);
nor UO_1600 (O_1600,N_29907,N_29834);
or UO_1601 (O_1601,N_29891,N_29935);
nand UO_1602 (O_1602,N_29803,N_29873);
nand UO_1603 (O_1603,N_29864,N_29780);
or UO_1604 (O_1604,N_29759,N_29922);
and UO_1605 (O_1605,N_29704,N_29862);
and UO_1606 (O_1606,N_29988,N_29954);
or UO_1607 (O_1607,N_29906,N_29939);
and UO_1608 (O_1608,N_29716,N_29862);
nor UO_1609 (O_1609,N_29972,N_29766);
xor UO_1610 (O_1610,N_29739,N_29727);
nand UO_1611 (O_1611,N_29968,N_29764);
and UO_1612 (O_1612,N_29739,N_29933);
nor UO_1613 (O_1613,N_29802,N_29822);
and UO_1614 (O_1614,N_29736,N_29914);
and UO_1615 (O_1615,N_29972,N_29855);
nor UO_1616 (O_1616,N_29858,N_29866);
xnor UO_1617 (O_1617,N_29840,N_29801);
or UO_1618 (O_1618,N_29798,N_29744);
xor UO_1619 (O_1619,N_29775,N_29866);
xnor UO_1620 (O_1620,N_29719,N_29872);
and UO_1621 (O_1621,N_29770,N_29807);
xor UO_1622 (O_1622,N_29774,N_29794);
xor UO_1623 (O_1623,N_29956,N_29969);
or UO_1624 (O_1624,N_29738,N_29735);
xnor UO_1625 (O_1625,N_29732,N_29952);
nand UO_1626 (O_1626,N_29958,N_29866);
xnor UO_1627 (O_1627,N_29823,N_29782);
nor UO_1628 (O_1628,N_29854,N_29723);
nor UO_1629 (O_1629,N_29937,N_29808);
xor UO_1630 (O_1630,N_29747,N_29892);
nor UO_1631 (O_1631,N_29734,N_29742);
nand UO_1632 (O_1632,N_29801,N_29983);
or UO_1633 (O_1633,N_29843,N_29772);
or UO_1634 (O_1634,N_29989,N_29968);
or UO_1635 (O_1635,N_29903,N_29725);
or UO_1636 (O_1636,N_29730,N_29736);
xnor UO_1637 (O_1637,N_29757,N_29949);
or UO_1638 (O_1638,N_29979,N_29957);
nand UO_1639 (O_1639,N_29933,N_29763);
and UO_1640 (O_1640,N_29806,N_29727);
xor UO_1641 (O_1641,N_29876,N_29938);
nand UO_1642 (O_1642,N_29928,N_29751);
xor UO_1643 (O_1643,N_29842,N_29758);
nor UO_1644 (O_1644,N_29919,N_29891);
or UO_1645 (O_1645,N_29886,N_29842);
nand UO_1646 (O_1646,N_29962,N_29995);
or UO_1647 (O_1647,N_29841,N_29945);
nand UO_1648 (O_1648,N_29804,N_29862);
nand UO_1649 (O_1649,N_29851,N_29768);
xnor UO_1650 (O_1650,N_29868,N_29793);
nor UO_1651 (O_1651,N_29739,N_29899);
and UO_1652 (O_1652,N_29972,N_29820);
and UO_1653 (O_1653,N_29854,N_29876);
xnor UO_1654 (O_1654,N_29999,N_29925);
xor UO_1655 (O_1655,N_29761,N_29938);
xor UO_1656 (O_1656,N_29732,N_29989);
and UO_1657 (O_1657,N_29985,N_29792);
nor UO_1658 (O_1658,N_29745,N_29922);
xor UO_1659 (O_1659,N_29702,N_29912);
or UO_1660 (O_1660,N_29856,N_29898);
nand UO_1661 (O_1661,N_29899,N_29874);
nor UO_1662 (O_1662,N_29885,N_29747);
and UO_1663 (O_1663,N_29931,N_29983);
nand UO_1664 (O_1664,N_29807,N_29908);
and UO_1665 (O_1665,N_29755,N_29737);
and UO_1666 (O_1666,N_29702,N_29736);
nand UO_1667 (O_1667,N_29777,N_29789);
nand UO_1668 (O_1668,N_29932,N_29727);
nor UO_1669 (O_1669,N_29913,N_29857);
and UO_1670 (O_1670,N_29987,N_29890);
nor UO_1671 (O_1671,N_29880,N_29780);
xnor UO_1672 (O_1672,N_29872,N_29954);
or UO_1673 (O_1673,N_29879,N_29885);
and UO_1674 (O_1674,N_29852,N_29916);
and UO_1675 (O_1675,N_29941,N_29863);
nor UO_1676 (O_1676,N_29947,N_29969);
nand UO_1677 (O_1677,N_29903,N_29991);
nand UO_1678 (O_1678,N_29977,N_29749);
xnor UO_1679 (O_1679,N_29916,N_29963);
nor UO_1680 (O_1680,N_29800,N_29961);
or UO_1681 (O_1681,N_29943,N_29996);
and UO_1682 (O_1682,N_29738,N_29799);
and UO_1683 (O_1683,N_29946,N_29843);
xnor UO_1684 (O_1684,N_29789,N_29997);
xor UO_1685 (O_1685,N_29713,N_29718);
and UO_1686 (O_1686,N_29858,N_29786);
nand UO_1687 (O_1687,N_29831,N_29755);
and UO_1688 (O_1688,N_29774,N_29956);
xor UO_1689 (O_1689,N_29755,N_29703);
nand UO_1690 (O_1690,N_29965,N_29798);
nor UO_1691 (O_1691,N_29883,N_29997);
nand UO_1692 (O_1692,N_29788,N_29784);
xor UO_1693 (O_1693,N_29791,N_29720);
and UO_1694 (O_1694,N_29750,N_29712);
xnor UO_1695 (O_1695,N_29801,N_29965);
nand UO_1696 (O_1696,N_29990,N_29940);
xor UO_1697 (O_1697,N_29766,N_29826);
or UO_1698 (O_1698,N_29756,N_29720);
and UO_1699 (O_1699,N_29792,N_29769);
xnor UO_1700 (O_1700,N_29900,N_29711);
and UO_1701 (O_1701,N_29829,N_29855);
nor UO_1702 (O_1702,N_29949,N_29818);
and UO_1703 (O_1703,N_29714,N_29719);
nor UO_1704 (O_1704,N_29745,N_29889);
nand UO_1705 (O_1705,N_29844,N_29704);
and UO_1706 (O_1706,N_29744,N_29782);
or UO_1707 (O_1707,N_29745,N_29774);
or UO_1708 (O_1708,N_29742,N_29820);
or UO_1709 (O_1709,N_29875,N_29870);
and UO_1710 (O_1710,N_29994,N_29968);
nor UO_1711 (O_1711,N_29927,N_29773);
xor UO_1712 (O_1712,N_29974,N_29753);
nand UO_1713 (O_1713,N_29917,N_29943);
and UO_1714 (O_1714,N_29866,N_29810);
or UO_1715 (O_1715,N_29738,N_29833);
and UO_1716 (O_1716,N_29882,N_29937);
and UO_1717 (O_1717,N_29708,N_29872);
and UO_1718 (O_1718,N_29923,N_29841);
nor UO_1719 (O_1719,N_29950,N_29989);
nor UO_1720 (O_1720,N_29796,N_29894);
or UO_1721 (O_1721,N_29852,N_29908);
and UO_1722 (O_1722,N_29722,N_29945);
nand UO_1723 (O_1723,N_29912,N_29831);
nand UO_1724 (O_1724,N_29840,N_29843);
xor UO_1725 (O_1725,N_29927,N_29915);
and UO_1726 (O_1726,N_29984,N_29718);
nor UO_1727 (O_1727,N_29945,N_29869);
xor UO_1728 (O_1728,N_29879,N_29771);
and UO_1729 (O_1729,N_29811,N_29914);
xnor UO_1730 (O_1730,N_29862,N_29969);
nor UO_1731 (O_1731,N_29851,N_29726);
nor UO_1732 (O_1732,N_29907,N_29900);
and UO_1733 (O_1733,N_29994,N_29756);
nor UO_1734 (O_1734,N_29950,N_29792);
nor UO_1735 (O_1735,N_29835,N_29897);
xor UO_1736 (O_1736,N_29765,N_29912);
nor UO_1737 (O_1737,N_29856,N_29990);
and UO_1738 (O_1738,N_29842,N_29704);
xor UO_1739 (O_1739,N_29875,N_29770);
xor UO_1740 (O_1740,N_29714,N_29787);
and UO_1741 (O_1741,N_29994,N_29862);
xor UO_1742 (O_1742,N_29866,N_29800);
and UO_1743 (O_1743,N_29892,N_29913);
and UO_1744 (O_1744,N_29798,N_29897);
or UO_1745 (O_1745,N_29888,N_29739);
nand UO_1746 (O_1746,N_29902,N_29746);
or UO_1747 (O_1747,N_29724,N_29898);
and UO_1748 (O_1748,N_29775,N_29998);
nand UO_1749 (O_1749,N_29830,N_29839);
and UO_1750 (O_1750,N_29925,N_29907);
nand UO_1751 (O_1751,N_29981,N_29828);
nand UO_1752 (O_1752,N_29890,N_29752);
nor UO_1753 (O_1753,N_29929,N_29764);
or UO_1754 (O_1754,N_29778,N_29938);
nor UO_1755 (O_1755,N_29832,N_29905);
nand UO_1756 (O_1756,N_29780,N_29874);
and UO_1757 (O_1757,N_29882,N_29908);
nor UO_1758 (O_1758,N_29881,N_29831);
nand UO_1759 (O_1759,N_29801,N_29896);
and UO_1760 (O_1760,N_29874,N_29932);
and UO_1761 (O_1761,N_29770,N_29825);
nand UO_1762 (O_1762,N_29729,N_29894);
nor UO_1763 (O_1763,N_29840,N_29903);
nor UO_1764 (O_1764,N_29988,N_29711);
and UO_1765 (O_1765,N_29883,N_29918);
and UO_1766 (O_1766,N_29951,N_29866);
or UO_1767 (O_1767,N_29741,N_29882);
nand UO_1768 (O_1768,N_29856,N_29716);
nand UO_1769 (O_1769,N_29839,N_29852);
and UO_1770 (O_1770,N_29895,N_29897);
nand UO_1771 (O_1771,N_29774,N_29993);
or UO_1772 (O_1772,N_29705,N_29965);
nor UO_1773 (O_1773,N_29998,N_29824);
nand UO_1774 (O_1774,N_29736,N_29985);
nand UO_1775 (O_1775,N_29865,N_29996);
nor UO_1776 (O_1776,N_29815,N_29706);
and UO_1777 (O_1777,N_29772,N_29903);
nor UO_1778 (O_1778,N_29871,N_29732);
nand UO_1779 (O_1779,N_29702,N_29970);
nor UO_1780 (O_1780,N_29877,N_29912);
and UO_1781 (O_1781,N_29748,N_29922);
or UO_1782 (O_1782,N_29785,N_29948);
or UO_1783 (O_1783,N_29955,N_29883);
nand UO_1784 (O_1784,N_29787,N_29946);
nor UO_1785 (O_1785,N_29884,N_29784);
nand UO_1786 (O_1786,N_29898,N_29917);
nand UO_1787 (O_1787,N_29878,N_29789);
xor UO_1788 (O_1788,N_29914,N_29854);
nand UO_1789 (O_1789,N_29907,N_29817);
or UO_1790 (O_1790,N_29972,N_29877);
or UO_1791 (O_1791,N_29710,N_29911);
and UO_1792 (O_1792,N_29801,N_29761);
xor UO_1793 (O_1793,N_29991,N_29799);
or UO_1794 (O_1794,N_29703,N_29719);
xor UO_1795 (O_1795,N_29957,N_29796);
xnor UO_1796 (O_1796,N_29860,N_29759);
xor UO_1797 (O_1797,N_29972,N_29782);
xnor UO_1798 (O_1798,N_29875,N_29726);
nor UO_1799 (O_1799,N_29839,N_29992);
xor UO_1800 (O_1800,N_29971,N_29734);
nand UO_1801 (O_1801,N_29721,N_29910);
or UO_1802 (O_1802,N_29928,N_29842);
xnor UO_1803 (O_1803,N_29734,N_29982);
or UO_1804 (O_1804,N_29785,N_29742);
nand UO_1805 (O_1805,N_29907,N_29941);
nor UO_1806 (O_1806,N_29725,N_29791);
xnor UO_1807 (O_1807,N_29920,N_29758);
nand UO_1808 (O_1808,N_29886,N_29898);
or UO_1809 (O_1809,N_29933,N_29954);
nand UO_1810 (O_1810,N_29857,N_29851);
xor UO_1811 (O_1811,N_29734,N_29799);
xor UO_1812 (O_1812,N_29822,N_29825);
nor UO_1813 (O_1813,N_29756,N_29919);
and UO_1814 (O_1814,N_29977,N_29837);
nand UO_1815 (O_1815,N_29788,N_29995);
nor UO_1816 (O_1816,N_29807,N_29734);
nand UO_1817 (O_1817,N_29944,N_29742);
nor UO_1818 (O_1818,N_29765,N_29982);
xor UO_1819 (O_1819,N_29957,N_29996);
and UO_1820 (O_1820,N_29763,N_29734);
nand UO_1821 (O_1821,N_29915,N_29754);
nand UO_1822 (O_1822,N_29706,N_29963);
and UO_1823 (O_1823,N_29954,N_29819);
or UO_1824 (O_1824,N_29929,N_29798);
nor UO_1825 (O_1825,N_29750,N_29922);
or UO_1826 (O_1826,N_29945,N_29940);
and UO_1827 (O_1827,N_29848,N_29808);
and UO_1828 (O_1828,N_29898,N_29914);
nor UO_1829 (O_1829,N_29893,N_29854);
xnor UO_1830 (O_1830,N_29841,N_29736);
nand UO_1831 (O_1831,N_29972,N_29996);
nand UO_1832 (O_1832,N_29992,N_29841);
nor UO_1833 (O_1833,N_29970,N_29895);
nor UO_1834 (O_1834,N_29864,N_29975);
or UO_1835 (O_1835,N_29951,N_29782);
nand UO_1836 (O_1836,N_29798,N_29913);
or UO_1837 (O_1837,N_29712,N_29899);
or UO_1838 (O_1838,N_29755,N_29947);
nand UO_1839 (O_1839,N_29759,N_29775);
nor UO_1840 (O_1840,N_29744,N_29898);
or UO_1841 (O_1841,N_29747,N_29817);
or UO_1842 (O_1842,N_29980,N_29772);
nand UO_1843 (O_1843,N_29745,N_29755);
nand UO_1844 (O_1844,N_29840,N_29930);
nor UO_1845 (O_1845,N_29833,N_29913);
or UO_1846 (O_1846,N_29951,N_29727);
and UO_1847 (O_1847,N_29926,N_29937);
nor UO_1848 (O_1848,N_29901,N_29958);
or UO_1849 (O_1849,N_29923,N_29977);
and UO_1850 (O_1850,N_29803,N_29777);
or UO_1851 (O_1851,N_29760,N_29793);
xnor UO_1852 (O_1852,N_29932,N_29951);
and UO_1853 (O_1853,N_29910,N_29812);
xnor UO_1854 (O_1854,N_29773,N_29998);
xor UO_1855 (O_1855,N_29923,N_29881);
and UO_1856 (O_1856,N_29841,N_29993);
nand UO_1857 (O_1857,N_29779,N_29865);
and UO_1858 (O_1858,N_29854,N_29920);
or UO_1859 (O_1859,N_29795,N_29750);
xnor UO_1860 (O_1860,N_29798,N_29880);
xnor UO_1861 (O_1861,N_29711,N_29879);
or UO_1862 (O_1862,N_29739,N_29927);
or UO_1863 (O_1863,N_29730,N_29968);
nor UO_1864 (O_1864,N_29936,N_29960);
nand UO_1865 (O_1865,N_29769,N_29843);
nor UO_1866 (O_1866,N_29734,N_29923);
and UO_1867 (O_1867,N_29930,N_29800);
and UO_1868 (O_1868,N_29965,N_29929);
or UO_1869 (O_1869,N_29968,N_29990);
nor UO_1870 (O_1870,N_29877,N_29760);
and UO_1871 (O_1871,N_29802,N_29989);
nor UO_1872 (O_1872,N_29967,N_29966);
or UO_1873 (O_1873,N_29960,N_29800);
nand UO_1874 (O_1874,N_29925,N_29913);
xnor UO_1875 (O_1875,N_29764,N_29854);
xnor UO_1876 (O_1876,N_29725,N_29706);
or UO_1877 (O_1877,N_29770,N_29761);
xor UO_1878 (O_1878,N_29882,N_29748);
or UO_1879 (O_1879,N_29833,N_29993);
nor UO_1880 (O_1880,N_29937,N_29803);
nor UO_1881 (O_1881,N_29773,N_29894);
nand UO_1882 (O_1882,N_29904,N_29842);
and UO_1883 (O_1883,N_29931,N_29794);
or UO_1884 (O_1884,N_29862,N_29735);
or UO_1885 (O_1885,N_29788,N_29781);
and UO_1886 (O_1886,N_29739,N_29821);
nand UO_1887 (O_1887,N_29930,N_29873);
nor UO_1888 (O_1888,N_29704,N_29808);
or UO_1889 (O_1889,N_29859,N_29988);
nor UO_1890 (O_1890,N_29730,N_29981);
and UO_1891 (O_1891,N_29768,N_29894);
nor UO_1892 (O_1892,N_29753,N_29837);
nor UO_1893 (O_1893,N_29705,N_29977);
nand UO_1894 (O_1894,N_29918,N_29843);
nand UO_1895 (O_1895,N_29733,N_29904);
nand UO_1896 (O_1896,N_29746,N_29945);
and UO_1897 (O_1897,N_29903,N_29980);
xnor UO_1898 (O_1898,N_29956,N_29753);
nor UO_1899 (O_1899,N_29747,N_29883);
xor UO_1900 (O_1900,N_29927,N_29753);
or UO_1901 (O_1901,N_29992,N_29846);
nand UO_1902 (O_1902,N_29757,N_29868);
nor UO_1903 (O_1903,N_29940,N_29797);
and UO_1904 (O_1904,N_29976,N_29850);
and UO_1905 (O_1905,N_29748,N_29948);
or UO_1906 (O_1906,N_29897,N_29959);
nor UO_1907 (O_1907,N_29760,N_29773);
nor UO_1908 (O_1908,N_29787,N_29998);
nand UO_1909 (O_1909,N_29804,N_29777);
xor UO_1910 (O_1910,N_29754,N_29724);
nand UO_1911 (O_1911,N_29733,N_29956);
or UO_1912 (O_1912,N_29954,N_29947);
and UO_1913 (O_1913,N_29854,N_29777);
nor UO_1914 (O_1914,N_29979,N_29706);
nor UO_1915 (O_1915,N_29957,N_29712);
nor UO_1916 (O_1916,N_29855,N_29923);
or UO_1917 (O_1917,N_29897,N_29702);
and UO_1918 (O_1918,N_29818,N_29760);
or UO_1919 (O_1919,N_29798,N_29951);
nand UO_1920 (O_1920,N_29729,N_29957);
nor UO_1921 (O_1921,N_29899,N_29785);
nand UO_1922 (O_1922,N_29895,N_29723);
and UO_1923 (O_1923,N_29828,N_29984);
nand UO_1924 (O_1924,N_29870,N_29744);
nand UO_1925 (O_1925,N_29795,N_29863);
or UO_1926 (O_1926,N_29786,N_29860);
nor UO_1927 (O_1927,N_29795,N_29947);
nor UO_1928 (O_1928,N_29839,N_29939);
and UO_1929 (O_1929,N_29901,N_29937);
nor UO_1930 (O_1930,N_29842,N_29986);
and UO_1931 (O_1931,N_29801,N_29827);
and UO_1932 (O_1932,N_29737,N_29919);
nor UO_1933 (O_1933,N_29988,N_29846);
nor UO_1934 (O_1934,N_29844,N_29864);
or UO_1935 (O_1935,N_29796,N_29961);
xor UO_1936 (O_1936,N_29871,N_29797);
nand UO_1937 (O_1937,N_29791,N_29985);
nor UO_1938 (O_1938,N_29746,N_29717);
and UO_1939 (O_1939,N_29831,N_29853);
or UO_1940 (O_1940,N_29839,N_29768);
and UO_1941 (O_1941,N_29967,N_29718);
xnor UO_1942 (O_1942,N_29776,N_29850);
xor UO_1943 (O_1943,N_29844,N_29916);
nand UO_1944 (O_1944,N_29934,N_29859);
nor UO_1945 (O_1945,N_29967,N_29847);
nand UO_1946 (O_1946,N_29760,N_29803);
or UO_1947 (O_1947,N_29875,N_29837);
or UO_1948 (O_1948,N_29983,N_29847);
and UO_1949 (O_1949,N_29797,N_29866);
and UO_1950 (O_1950,N_29737,N_29797);
or UO_1951 (O_1951,N_29977,N_29974);
nand UO_1952 (O_1952,N_29727,N_29926);
and UO_1953 (O_1953,N_29703,N_29945);
nor UO_1954 (O_1954,N_29845,N_29947);
xor UO_1955 (O_1955,N_29819,N_29876);
nor UO_1956 (O_1956,N_29757,N_29834);
and UO_1957 (O_1957,N_29772,N_29899);
and UO_1958 (O_1958,N_29934,N_29817);
xnor UO_1959 (O_1959,N_29741,N_29790);
nand UO_1960 (O_1960,N_29858,N_29908);
nand UO_1961 (O_1961,N_29959,N_29870);
nand UO_1962 (O_1962,N_29721,N_29937);
nor UO_1963 (O_1963,N_29861,N_29895);
nor UO_1964 (O_1964,N_29816,N_29871);
or UO_1965 (O_1965,N_29714,N_29748);
or UO_1966 (O_1966,N_29790,N_29848);
xnor UO_1967 (O_1967,N_29835,N_29748);
nor UO_1968 (O_1968,N_29866,N_29887);
nor UO_1969 (O_1969,N_29880,N_29954);
nand UO_1970 (O_1970,N_29903,N_29893);
xor UO_1971 (O_1971,N_29834,N_29822);
or UO_1972 (O_1972,N_29823,N_29817);
or UO_1973 (O_1973,N_29813,N_29863);
nand UO_1974 (O_1974,N_29972,N_29713);
xor UO_1975 (O_1975,N_29717,N_29948);
and UO_1976 (O_1976,N_29786,N_29953);
and UO_1977 (O_1977,N_29809,N_29868);
xor UO_1978 (O_1978,N_29941,N_29717);
or UO_1979 (O_1979,N_29732,N_29705);
nor UO_1980 (O_1980,N_29849,N_29908);
xor UO_1981 (O_1981,N_29816,N_29741);
and UO_1982 (O_1982,N_29755,N_29769);
and UO_1983 (O_1983,N_29718,N_29747);
nor UO_1984 (O_1984,N_29989,N_29770);
xor UO_1985 (O_1985,N_29908,N_29876);
nor UO_1986 (O_1986,N_29881,N_29771);
or UO_1987 (O_1987,N_29858,N_29997);
xor UO_1988 (O_1988,N_29836,N_29785);
xnor UO_1989 (O_1989,N_29742,N_29717);
nand UO_1990 (O_1990,N_29818,N_29805);
and UO_1991 (O_1991,N_29962,N_29706);
nor UO_1992 (O_1992,N_29937,N_29841);
xor UO_1993 (O_1993,N_29830,N_29785);
nor UO_1994 (O_1994,N_29888,N_29850);
and UO_1995 (O_1995,N_29963,N_29734);
xnor UO_1996 (O_1996,N_29744,N_29716);
xor UO_1997 (O_1997,N_29923,N_29740);
or UO_1998 (O_1998,N_29917,N_29907);
and UO_1999 (O_1999,N_29801,N_29820);
or UO_2000 (O_2000,N_29859,N_29783);
nand UO_2001 (O_2001,N_29909,N_29802);
nor UO_2002 (O_2002,N_29996,N_29817);
and UO_2003 (O_2003,N_29747,N_29989);
xor UO_2004 (O_2004,N_29704,N_29962);
nor UO_2005 (O_2005,N_29815,N_29899);
xor UO_2006 (O_2006,N_29980,N_29848);
xnor UO_2007 (O_2007,N_29851,N_29776);
or UO_2008 (O_2008,N_29966,N_29867);
or UO_2009 (O_2009,N_29862,N_29844);
nor UO_2010 (O_2010,N_29900,N_29875);
or UO_2011 (O_2011,N_29894,N_29882);
and UO_2012 (O_2012,N_29707,N_29744);
xor UO_2013 (O_2013,N_29971,N_29773);
nand UO_2014 (O_2014,N_29905,N_29822);
and UO_2015 (O_2015,N_29946,N_29731);
and UO_2016 (O_2016,N_29740,N_29841);
xor UO_2017 (O_2017,N_29957,N_29904);
xnor UO_2018 (O_2018,N_29740,N_29742);
xnor UO_2019 (O_2019,N_29942,N_29913);
xor UO_2020 (O_2020,N_29794,N_29998);
nor UO_2021 (O_2021,N_29709,N_29988);
nand UO_2022 (O_2022,N_29830,N_29780);
xor UO_2023 (O_2023,N_29912,N_29908);
nor UO_2024 (O_2024,N_29836,N_29781);
nand UO_2025 (O_2025,N_29927,N_29725);
and UO_2026 (O_2026,N_29774,N_29735);
nor UO_2027 (O_2027,N_29979,N_29848);
nor UO_2028 (O_2028,N_29993,N_29824);
nand UO_2029 (O_2029,N_29851,N_29787);
nor UO_2030 (O_2030,N_29744,N_29796);
nor UO_2031 (O_2031,N_29794,N_29861);
nand UO_2032 (O_2032,N_29803,N_29917);
nand UO_2033 (O_2033,N_29778,N_29802);
or UO_2034 (O_2034,N_29946,N_29945);
nand UO_2035 (O_2035,N_29900,N_29873);
nand UO_2036 (O_2036,N_29877,N_29996);
and UO_2037 (O_2037,N_29961,N_29757);
and UO_2038 (O_2038,N_29906,N_29896);
and UO_2039 (O_2039,N_29741,N_29789);
or UO_2040 (O_2040,N_29933,N_29998);
nand UO_2041 (O_2041,N_29848,N_29792);
xnor UO_2042 (O_2042,N_29903,N_29794);
xnor UO_2043 (O_2043,N_29760,N_29814);
xnor UO_2044 (O_2044,N_29890,N_29981);
nand UO_2045 (O_2045,N_29762,N_29715);
nor UO_2046 (O_2046,N_29754,N_29823);
or UO_2047 (O_2047,N_29812,N_29802);
or UO_2048 (O_2048,N_29920,N_29879);
and UO_2049 (O_2049,N_29980,N_29841);
nand UO_2050 (O_2050,N_29848,N_29946);
nand UO_2051 (O_2051,N_29808,N_29842);
xnor UO_2052 (O_2052,N_29730,N_29935);
or UO_2053 (O_2053,N_29843,N_29954);
nor UO_2054 (O_2054,N_29798,N_29959);
xnor UO_2055 (O_2055,N_29720,N_29846);
nand UO_2056 (O_2056,N_29753,N_29769);
or UO_2057 (O_2057,N_29779,N_29700);
or UO_2058 (O_2058,N_29772,N_29712);
nand UO_2059 (O_2059,N_29815,N_29763);
nand UO_2060 (O_2060,N_29836,N_29749);
nor UO_2061 (O_2061,N_29877,N_29869);
and UO_2062 (O_2062,N_29885,N_29746);
xor UO_2063 (O_2063,N_29941,N_29869);
xor UO_2064 (O_2064,N_29802,N_29938);
or UO_2065 (O_2065,N_29917,N_29984);
and UO_2066 (O_2066,N_29885,N_29977);
nor UO_2067 (O_2067,N_29803,N_29886);
xnor UO_2068 (O_2068,N_29749,N_29948);
xor UO_2069 (O_2069,N_29707,N_29779);
nor UO_2070 (O_2070,N_29917,N_29997);
or UO_2071 (O_2071,N_29924,N_29816);
nand UO_2072 (O_2072,N_29945,N_29855);
xor UO_2073 (O_2073,N_29978,N_29932);
and UO_2074 (O_2074,N_29784,N_29858);
nor UO_2075 (O_2075,N_29726,N_29800);
nor UO_2076 (O_2076,N_29896,N_29951);
nor UO_2077 (O_2077,N_29785,N_29904);
xnor UO_2078 (O_2078,N_29858,N_29844);
and UO_2079 (O_2079,N_29818,N_29907);
nor UO_2080 (O_2080,N_29755,N_29869);
nor UO_2081 (O_2081,N_29867,N_29960);
nand UO_2082 (O_2082,N_29914,N_29845);
xnor UO_2083 (O_2083,N_29833,N_29827);
or UO_2084 (O_2084,N_29710,N_29916);
xnor UO_2085 (O_2085,N_29988,N_29760);
xor UO_2086 (O_2086,N_29908,N_29861);
nand UO_2087 (O_2087,N_29927,N_29736);
and UO_2088 (O_2088,N_29904,N_29881);
nor UO_2089 (O_2089,N_29901,N_29897);
or UO_2090 (O_2090,N_29760,N_29729);
xnor UO_2091 (O_2091,N_29729,N_29724);
xor UO_2092 (O_2092,N_29974,N_29704);
or UO_2093 (O_2093,N_29894,N_29805);
nand UO_2094 (O_2094,N_29950,N_29881);
nand UO_2095 (O_2095,N_29921,N_29763);
xor UO_2096 (O_2096,N_29752,N_29885);
nor UO_2097 (O_2097,N_29711,N_29899);
xnor UO_2098 (O_2098,N_29911,N_29789);
xor UO_2099 (O_2099,N_29806,N_29900);
xor UO_2100 (O_2100,N_29701,N_29861);
or UO_2101 (O_2101,N_29784,N_29707);
xnor UO_2102 (O_2102,N_29866,N_29991);
xnor UO_2103 (O_2103,N_29959,N_29999);
nor UO_2104 (O_2104,N_29828,N_29905);
or UO_2105 (O_2105,N_29772,N_29815);
and UO_2106 (O_2106,N_29764,N_29757);
and UO_2107 (O_2107,N_29816,N_29739);
or UO_2108 (O_2108,N_29929,N_29955);
nor UO_2109 (O_2109,N_29802,N_29988);
or UO_2110 (O_2110,N_29800,N_29773);
nand UO_2111 (O_2111,N_29980,N_29746);
or UO_2112 (O_2112,N_29701,N_29767);
or UO_2113 (O_2113,N_29702,N_29892);
xnor UO_2114 (O_2114,N_29984,N_29948);
nand UO_2115 (O_2115,N_29846,N_29994);
or UO_2116 (O_2116,N_29882,N_29856);
nand UO_2117 (O_2117,N_29986,N_29933);
and UO_2118 (O_2118,N_29923,N_29838);
or UO_2119 (O_2119,N_29757,N_29716);
xnor UO_2120 (O_2120,N_29751,N_29892);
or UO_2121 (O_2121,N_29835,N_29933);
or UO_2122 (O_2122,N_29779,N_29736);
or UO_2123 (O_2123,N_29992,N_29758);
nand UO_2124 (O_2124,N_29957,N_29905);
nor UO_2125 (O_2125,N_29947,N_29980);
or UO_2126 (O_2126,N_29925,N_29971);
xnor UO_2127 (O_2127,N_29992,N_29802);
nor UO_2128 (O_2128,N_29806,N_29848);
or UO_2129 (O_2129,N_29724,N_29955);
nor UO_2130 (O_2130,N_29819,N_29883);
or UO_2131 (O_2131,N_29828,N_29722);
xor UO_2132 (O_2132,N_29867,N_29925);
nor UO_2133 (O_2133,N_29800,N_29850);
xor UO_2134 (O_2134,N_29933,N_29964);
nor UO_2135 (O_2135,N_29861,N_29760);
or UO_2136 (O_2136,N_29979,N_29741);
or UO_2137 (O_2137,N_29892,N_29871);
and UO_2138 (O_2138,N_29937,N_29786);
and UO_2139 (O_2139,N_29849,N_29873);
or UO_2140 (O_2140,N_29800,N_29820);
nor UO_2141 (O_2141,N_29729,N_29795);
nand UO_2142 (O_2142,N_29995,N_29834);
nor UO_2143 (O_2143,N_29832,N_29989);
nor UO_2144 (O_2144,N_29720,N_29889);
nand UO_2145 (O_2145,N_29888,N_29991);
nor UO_2146 (O_2146,N_29815,N_29922);
nor UO_2147 (O_2147,N_29983,N_29840);
or UO_2148 (O_2148,N_29975,N_29823);
nand UO_2149 (O_2149,N_29878,N_29956);
xor UO_2150 (O_2150,N_29976,N_29746);
or UO_2151 (O_2151,N_29875,N_29816);
nor UO_2152 (O_2152,N_29766,N_29768);
nor UO_2153 (O_2153,N_29713,N_29915);
xor UO_2154 (O_2154,N_29741,N_29781);
nor UO_2155 (O_2155,N_29721,N_29785);
xor UO_2156 (O_2156,N_29962,N_29863);
and UO_2157 (O_2157,N_29985,N_29876);
or UO_2158 (O_2158,N_29752,N_29835);
or UO_2159 (O_2159,N_29848,N_29758);
or UO_2160 (O_2160,N_29848,N_29919);
or UO_2161 (O_2161,N_29817,N_29820);
nand UO_2162 (O_2162,N_29860,N_29976);
or UO_2163 (O_2163,N_29839,N_29981);
nor UO_2164 (O_2164,N_29765,N_29985);
or UO_2165 (O_2165,N_29740,N_29772);
nor UO_2166 (O_2166,N_29896,N_29710);
nand UO_2167 (O_2167,N_29985,N_29738);
and UO_2168 (O_2168,N_29707,N_29979);
and UO_2169 (O_2169,N_29882,N_29805);
or UO_2170 (O_2170,N_29856,N_29752);
nand UO_2171 (O_2171,N_29750,N_29829);
nand UO_2172 (O_2172,N_29725,N_29711);
nor UO_2173 (O_2173,N_29855,N_29887);
xor UO_2174 (O_2174,N_29843,N_29994);
nor UO_2175 (O_2175,N_29837,N_29711);
xnor UO_2176 (O_2176,N_29744,N_29936);
and UO_2177 (O_2177,N_29993,N_29860);
xnor UO_2178 (O_2178,N_29921,N_29897);
nor UO_2179 (O_2179,N_29924,N_29964);
nor UO_2180 (O_2180,N_29829,N_29731);
nand UO_2181 (O_2181,N_29982,N_29771);
and UO_2182 (O_2182,N_29947,N_29972);
or UO_2183 (O_2183,N_29712,N_29945);
or UO_2184 (O_2184,N_29946,N_29863);
or UO_2185 (O_2185,N_29838,N_29765);
nor UO_2186 (O_2186,N_29852,N_29815);
nand UO_2187 (O_2187,N_29830,N_29882);
nand UO_2188 (O_2188,N_29842,N_29912);
nor UO_2189 (O_2189,N_29905,N_29780);
or UO_2190 (O_2190,N_29742,N_29877);
nand UO_2191 (O_2191,N_29785,N_29957);
xor UO_2192 (O_2192,N_29700,N_29907);
and UO_2193 (O_2193,N_29888,N_29930);
or UO_2194 (O_2194,N_29824,N_29757);
xor UO_2195 (O_2195,N_29835,N_29916);
and UO_2196 (O_2196,N_29881,N_29894);
and UO_2197 (O_2197,N_29925,N_29821);
nor UO_2198 (O_2198,N_29884,N_29971);
nand UO_2199 (O_2199,N_29785,N_29975);
nor UO_2200 (O_2200,N_29904,N_29987);
and UO_2201 (O_2201,N_29840,N_29964);
nor UO_2202 (O_2202,N_29817,N_29779);
xor UO_2203 (O_2203,N_29894,N_29830);
nand UO_2204 (O_2204,N_29852,N_29725);
and UO_2205 (O_2205,N_29930,N_29730);
or UO_2206 (O_2206,N_29981,N_29793);
nor UO_2207 (O_2207,N_29793,N_29896);
nand UO_2208 (O_2208,N_29806,N_29916);
and UO_2209 (O_2209,N_29973,N_29931);
and UO_2210 (O_2210,N_29844,N_29987);
xnor UO_2211 (O_2211,N_29897,N_29814);
and UO_2212 (O_2212,N_29919,N_29746);
xor UO_2213 (O_2213,N_29768,N_29995);
nand UO_2214 (O_2214,N_29775,N_29729);
or UO_2215 (O_2215,N_29773,N_29990);
or UO_2216 (O_2216,N_29778,N_29844);
nor UO_2217 (O_2217,N_29858,N_29952);
nor UO_2218 (O_2218,N_29874,N_29841);
nand UO_2219 (O_2219,N_29893,N_29942);
and UO_2220 (O_2220,N_29940,N_29863);
nor UO_2221 (O_2221,N_29730,N_29924);
and UO_2222 (O_2222,N_29755,N_29773);
and UO_2223 (O_2223,N_29736,N_29967);
xnor UO_2224 (O_2224,N_29973,N_29881);
nor UO_2225 (O_2225,N_29930,N_29993);
nand UO_2226 (O_2226,N_29754,N_29751);
nor UO_2227 (O_2227,N_29980,N_29898);
or UO_2228 (O_2228,N_29731,N_29802);
and UO_2229 (O_2229,N_29724,N_29881);
and UO_2230 (O_2230,N_29829,N_29895);
nor UO_2231 (O_2231,N_29913,N_29779);
and UO_2232 (O_2232,N_29966,N_29756);
nand UO_2233 (O_2233,N_29850,N_29919);
or UO_2234 (O_2234,N_29970,N_29744);
nand UO_2235 (O_2235,N_29756,N_29901);
or UO_2236 (O_2236,N_29915,N_29907);
nand UO_2237 (O_2237,N_29747,N_29940);
xnor UO_2238 (O_2238,N_29984,N_29918);
xor UO_2239 (O_2239,N_29802,N_29961);
or UO_2240 (O_2240,N_29870,N_29811);
and UO_2241 (O_2241,N_29891,N_29893);
and UO_2242 (O_2242,N_29741,N_29967);
nor UO_2243 (O_2243,N_29932,N_29922);
and UO_2244 (O_2244,N_29991,N_29881);
nor UO_2245 (O_2245,N_29892,N_29713);
and UO_2246 (O_2246,N_29914,N_29979);
nor UO_2247 (O_2247,N_29824,N_29747);
and UO_2248 (O_2248,N_29868,N_29758);
nor UO_2249 (O_2249,N_29968,N_29927);
xnor UO_2250 (O_2250,N_29905,N_29914);
and UO_2251 (O_2251,N_29771,N_29746);
nor UO_2252 (O_2252,N_29868,N_29937);
or UO_2253 (O_2253,N_29982,N_29795);
xor UO_2254 (O_2254,N_29977,N_29859);
or UO_2255 (O_2255,N_29788,N_29855);
nand UO_2256 (O_2256,N_29783,N_29763);
nand UO_2257 (O_2257,N_29721,N_29994);
or UO_2258 (O_2258,N_29864,N_29814);
and UO_2259 (O_2259,N_29926,N_29838);
or UO_2260 (O_2260,N_29815,N_29871);
or UO_2261 (O_2261,N_29822,N_29914);
xor UO_2262 (O_2262,N_29764,N_29819);
nand UO_2263 (O_2263,N_29783,N_29952);
and UO_2264 (O_2264,N_29772,N_29921);
nand UO_2265 (O_2265,N_29808,N_29878);
or UO_2266 (O_2266,N_29925,N_29770);
xnor UO_2267 (O_2267,N_29718,N_29919);
nand UO_2268 (O_2268,N_29911,N_29787);
xor UO_2269 (O_2269,N_29788,N_29977);
or UO_2270 (O_2270,N_29879,N_29812);
nand UO_2271 (O_2271,N_29965,N_29720);
nand UO_2272 (O_2272,N_29883,N_29785);
or UO_2273 (O_2273,N_29957,N_29799);
nor UO_2274 (O_2274,N_29847,N_29884);
nand UO_2275 (O_2275,N_29971,N_29761);
nor UO_2276 (O_2276,N_29864,N_29945);
nor UO_2277 (O_2277,N_29800,N_29776);
xnor UO_2278 (O_2278,N_29869,N_29901);
or UO_2279 (O_2279,N_29756,N_29849);
or UO_2280 (O_2280,N_29883,N_29708);
nor UO_2281 (O_2281,N_29850,N_29983);
or UO_2282 (O_2282,N_29965,N_29916);
or UO_2283 (O_2283,N_29990,N_29887);
and UO_2284 (O_2284,N_29886,N_29726);
or UO_2285 (O_2285,N_29703,N_29901);
nor UO_2286 (O_2286,N_29869,N_29772);
xnor UO_2287 (O_2287,N_29816,N_29983);
nor UO_2288 (O_2288,N_29844,N_29736);
and UO_2289 (O_2289,N_29835,N_29917);
and UO_2290 (O_2290,N_29719,N_29780);
xor UO_2291 (O_2291,N_29852,N_29925);
xnor UO_2292 (O_2292,N_29932,N_29748);
nand UO_2293 (O_2293,N_29843,N_29749);
nand UO_2294 (O_2294,N_29983,N_29888);
and UO_2295 (O_2295,N_29758,N_29863);
xnor UO_2296 (O_2296,N_29947,N_29701);
xor UO_2297 (O_2297,N_29772,N_29707);
or UO_2298 (O_2298,N_29717,N_29900);
nand UO_2299 (O_2299,N_29705,N_29712);
xor UO_2300 (O_2300,N_29848,N_29867);
or UO_2301 (O_2301,N_29960,N_29769);
nand UO_2302 (O_2302,N_29862,N_29711);
xnor UO_2303 (O_2303,N_29702,N_29846);
nor UO_2304 (O_2304,N_29798,N_29720);
and UO_2305 (O_2305,N_29820,N_29825);
nand UO_2306 (O_2306,N_29938,N_29920);
and UO_2307 (O_2307,N_29943,N_29873);
nor UO_2308 (O_2308,N_29705,N_29770);
or UO_2309 (O_2309,N_29788,N_29921);
and UO_2310 (O_2310,N_29947,N_29869);
or UO_2311 (O_2311,N_29785,N_29893);
nor UO_2312 (O_2312,N_29961,N_29995);
xor UO_2313 (O_2313,N_29990,N_29732);
nor UO_2314 (O_2314,N_29726,N_29841);
or UO_2315 (O_2315,N_29781,N_29700);
nor UO_2316 (O_2316,N_29842,N_29792);
or UO_2317 (O_2317,N_29933,N_29997);
or UO_2318 (O_2318,N_29878,N_29861);
and UO_2319 (O_2319,N_29725,N_29965);
nor UO_2320 (O_2320,N_29839,N_29746);
or UO_2321 (O_2321,N_29870,N_29897);
nor UO_2322 (O_2322,N_29999,N_29972);
nor UO_2323 (O_2323,N_29926,N_29811);
and UO_2324 (O_2324,N_29817,N_29734);
and UO_2325 (O_2325,N_29711,N_29978);
nor UO_2326 (O_2326,N_29755,N_29968);
nor UO_2327 (O_2327,N_29827,N_29985);
and UO_2328 (O_2328,N_29869,N_29903);
nand UO_2329 (O_2329,N_29731,N_29790);
or UO_2330 (O_2330,N_29799,N_29816);
nor UO_2331 (O_2331,N_29728,N_29788);
and UO_2332 (O_2332,N_29791,N_29754);
xor UO_2333 (O_2333,N_29986,N_29832);
nor UO_2334 (O_2334,N_29890,N_29874);
nor UO_2335 (O_2335,N_29788,N_29743);
nand UO_2336 (O_2336,N_29753,N_29701);
or UO_2337 (O_2337,N_29704,N_29767);
xor UO_2338 (O_2338,N_29727,N_29735);
xnor UO_2339 (O_2339,N_29866,N_29909);
nand UO_2340 (O_2340,N_29746,N_29940);
or UO_2341 (O_2341,N_29793,N_29903);
nand UO_2342 (O_2342,N_29961,N_29994);
nor UO_2343 (O_2343,N_29836,N_29912);
nand UO_2344 (O_2344,N_29731,N_29779);
or UO_2345 (O_2345,N_29722,N_29781);
or UO_2346 (O_2346,N_29890,N_29860);
nor UO_2347 (O_2347,N_29815,N_29736);
nor UO_2348 (O_2348,N_29953,N_29992);
and UO_2349 (O_2349,N_29798,N_29734);
or UO_2350 (O_2350,N_29729,N_29822);
or UO_2351 (O_2351,N_29786,N_29853);
nand UO_2352 (O_2352,N_29729,N_29750);
nand UO_2353 (O_2353,N_29915,N_29921);
and UO_2354 (O_2354,N_29968,N_29896);
and UO_2355 (O_2355,N_29743,N_29924);
or UO_2356 (O_2356,N_29932,N_29810);
nand UO_2357 (O_2357,N_29972,N_29927);
and UO_2358 (O_2358,N_29835,N_29732);
nand UO_2359 (O_2359,N_29895,N_29957);
nor UO_2360 (O_2360,N_29749,N_29982);
nand UO_2361 (O_2361,N_29803,N_29906);
or UO_2362 (O_2362,N_29973,N_29726);
xor UO_2363 (O_2363,N_29861,N_29955);
and UO_2364 (O_2364,N_29757,N_29711);
or UO_2365 (O_2365,N_29773,N_29930);
nor UO_2366 (O_2366,N_29892,N_29943);
and UO_2367 (O_2367,N_29847,N_29821);
nand UO_2368 (O_2368,N_29995,N_29886);
nor UO_2369 (O_2369,N_29927,N_29726);
nor UO_2370 (O_2370,N_29958,N_29786);
and UO_2371 (O_2371,N_29895,N_29781);
and UO_2372 (O_2372,N_29788,N_29703);
and UO_2373 (O_2373,N_29955,N_29766);
nor UO_2374 (O_2374,N_29751,N_29716);
xor UO_2375 (O_2375,N_29983,N_29886);
nand UO_2376 (O_2376,N_29899,N_29976);
nand UO_2377 (O_2377,N_29798,N_29876);
nor UO_2378 (O_2378,N_29896,N_29843);
nand UO_2379 (O_2379,N_29915,N_29987);
xor UO_2380 (O_2380,N_29880,N_29752);
or UO_2381 (O_2381,N_29966,N_29744);
or UO_2382 (O_2382,N_29934,N_29708);
nor UO_2383 (O_2383,N_29945,N_29964);
nor UO_2384 (O_2384,N_29949,N_29900);
nor UO_2385 (O_2385,N_29714,N_29844);
nand UO_2386 (O_2386,N_29793,N_29886);
nand UO_2387 (O_2387,N_29834,N_29728);
and UO_2388 (O_2388,N_29942,N_29726);
xnor UO_2389 (O_2389,N_29949,N_29823);
and UO_2390 (O_2390,N_29983,N_29949);
nand UO_2391 (O_2391,N_29774,N_29954);
nor UO_2392 (O_2392,N_29818,N_29940);
and UO_2393 (O_2393,N_29800,N_29934);
or UO_2394 (O_2394,N_29807,N_29702);
and UO_2395 (O_2395,N_29811,N_29766);
nor UO_2396 (O_2396,N_29901,N_29750);
or UO_2397 (O_2397,N_29761,N_29759);
nand UO_2398 (O_2398,N_29868,N_29935);
xor UO_2399 (O_2399,N_29742,N_29738);
or UO_2400 (O_2400,N_29966,N_29816);
nor UO_2401 (O_2401,N_29866,N_29917);
or UO_2402 (O_2402,N_29815,N_29878);
nand UO_2403 (O_2403,N_29726,N_29838);
and UO_2404 (O_2404,N_29709,N_29903);
xnor UO_2405 (O_2405,N_29996,N_29851);
nor UO_2406 (O_2406,N_29901,N_29844);
nor UO_2407 (O_2407,N_29796,N_29890);
nor UO_2408 (O_2408,N_29801,N_29960);
nand UO_2409 (O_2409,N_29733,N_29828);
or UO_2410 (O_2410,N_29974,N_29757);
nor UO_2411 (O_2411,N_29810,N_29799);
xor UO_2412 (O_2412,N_29840,N_29811);
nand UO_2413 (O_2413,N_29882,N_29810);
xor UO_2414 (O_2414,N_29881,N_29802);
nand UO_2415 (O_2415,N_29812,N_29991);
or UO_2416 (O_2416,N_29982,N_29823);
or UO_2417 (O_2417,N_29950,N_29764);
nand UO_2418 (O_2418,N_29913,N_29718);
and UO_2419 (O_2419,N_29744,N_29754);
xor UO_2420 (O_2420,N_29839,N_29931);
nand UO_2421 (O_2421,N_29789,N_29850);
or UO_2422 (O_2422,N_29701,N_29752);
and UO_2423 (O_2423,N_29856,N_29899);
nor UO_2424 (O_2424,N_29802,N_29785);
nor UO_2425 (O_2425,N_29705,N_29937);
and UO_2426 (O_2426,N_29737,N_29931);
nor UO_2427 (O_2427,N_29874,N_29782);
or UO_2428 (O_2428,N_29798,N_29952);
nor UO_2429 (O_2429,N_29958,N_29987);
nand UO_2430 (O_2430,N_29791,N_29962);
nand UO_2431 (O_2431,N_29920,N_29794);
nor UO_2432 (O_2432,N_29925,N_29710);
nand UO_2433 (O_2433,N_29955,N_29757);
nand UO_2434 (O_2434,N_29867,N_29945);
xnor UO_2435 (O_2435,N_29812,N_29800);
or UO_2436 (O_2436,N_29932,N_29923);
or UO_2437 (O_2437,N_29720,N_29817);
and UO_2438 (O_2438,N_29996,N_29755);
nor UO_2439 (O_2439,N_29777,N_29791);
and UO_2440 (O_2440,N_29929,N_29891);
xnor UO_2441 (O_2441,N_29748,N_29880);
nand UO_2442 (O_2442,N_29954,N_29802);
nor UO_2443 (O_2443,N_29810,N_29990);
nand UO_2444 (O_2444,N_29818,N_29711);
and UO_2445 (O_2445,N_29976,N_29839);
nor UO_2446 (O_2446,N_29982,N_29858);
and UO_2447 (O_2447,N_29887,N_29922);
or UO_2448 (O_2448,N_29881,N_29859);
nor UO_2449 (O_2449,N_29740,N_29978);
xnor UO_2450 (O_2450,N_29887,N_29778);
xnor UO_2451 (O_2451,N_29823,N_29860);
or UO_2452 (O_2452,N_29746,N_29969);
nor UO_2453 (O_2453,N_29748,N_29724);
nor UO_2454 (O_2454,N_29739,N_29720);
nand UO_2455 (O_2455,N_29883,N_29789);
and UO_2456 (O_2456,N_29762,N_29825);
or UO_2457 (O_2457,N_29902,N_29815);
and UO_2458 (O_2458,N_29818,N_29767);
xor UO_2459 (O_2459,N_29708,N_29771);
xnor UO_2460 (O_2460,N_29732,N_29985);
nor UO_2461 (O_2461,N_29817,N_29808);
xor UO_2462 (O_2462,N_29930,N_29831);
nand UO_2463 (O_2463,N_29996,N_29881);
xnor UO_2464 (O_2464,N_29853,N_29779);
nor UO_2465 (O_2465,N_29889,N_29923);
xnor UO_2466 (O_2466,N_29901,N_29705);
xor UO_2467 (O_2467,N_29934,N_29987);
xor UO_2468 (O_2468,N_29868,N_29899);
nor UO_2469 (O_2469,N_29831,N_29911);
nand UO_2470 (O_2470,N_29735,N_29882);
or UO_2471 (O_2471,N_29709,N_29710);
xnor UO_2472 (O_2472,N_29884,N_29915);
nand UO_2473 (O_2473,N_29929,N_29799);
nor UO_2474 (O_2474,N_29805,N_29724);
and UO_2475 (O_2475,N_29803,N_29763);
nor UO_2476 (O_2476,N_29701,N_29729);
nand UO_2477 (O_2477,N_29927,N_29826);
xor UO_2478 (O_2478,N_29705,N_29878);
nor UO_2479 (O_2479,N_29946,N_29928);
nand UO_2480 (O_2480,N_29714,N_29863);
or UO_2481 (O_2481,N_29800,N_29845);
and UO_2482 (O_2482,N_29956,N_29957);
or UO_2483 (O_2483,N_29973,N_29930);
xor UO_2484 (O_2484,N_29879,N_29938);
nor UO_2485 (O_2485,N_29907,N_29878);
and UO_2486 (O_2486,N_29995,N_29738);
or UO_2487 (O_2487,N_29846,N_29792);
nand UO_2488 (O_2488,N_29990,N_29704);
nor UO_2489 (O_2489,N_29773,N_29717);
or UO_2490 (O_2490,N_29969,N_29996);
nor UO_2491 (O_2491,N_29928,N_29981);
xor UO_2492 (O_2492,N_29741,N_29898);
or UO_2493 (O_2493,N_29846,N_29877);
nand UO_2494 (O_2494,N_29854,N_29864);
xor UO_2495 (O_2495,N_29882,N_29924);
or UO_2496 (O_2496,N_29886,N_29771);
nand UO_2497 (O_2497,N_29970,N_29745);
nand UO_2498 (O_2498,N_29769,N_29811);
nand UO_2499 (O_2499,N_29845,N_29863);
or UO_2500 (O_2500,N_29790,N_29879);
nand UO_2501 (O_2501,N_29969,N_29757);
or UO_2502 (O_2502,N_29764,N_29993);
xor UO_2503 (O_2503,N_29705,N_29992);
xnor UO_2504 (O_2504,N_29813,N_29767);
and UO_2505 (O_2505,N_29825,N_29715);
and UO_2506 (O_2506,N_29946,N_29991);
xor UO_2507 (O_2507,N_29730,N_29925);
xnor UO_2508 (O_2508,N_29736,N_29895);
xnor UO_2509 (O_2509,N_29914,N_29865);
nor UO_2510 (O_2510,N_29959,N_29911);
nor UO_2511 (O_2511,N_29921,N_29940);
nor UO_2512 (O_2512,N_29999,N_29860);
xor UO_2513 (O_2513,N_29865,N_29945);
nor UO_2514 (O_2514,N_29720,N_29884);
nand UO_2515 (O_2515,N_29984,N_29885);
xor UO_2516 (O_2516,N_29998,N_29899);
nand UO_2517 (O_2517,N_29740,N_29838);
nand UO_2518 (O_2518,N_29858,N_29708);
nor UO_2519 (O_2519,N_29772,N_29701);
or UO_2520 (O_2520,N_29811,N_29907);
nand UO_2521 (O_2521,N_29734,N_29773);
nand UO_2522 (O_2522,N_29835,N_29997);
or UO_2523 (O_2523,N_29771,N_29714);
or UO_2524 (O_2524,N_29767,N_29852);
xor UO_2525 (O_2525,N_29982,N_29748);
xor UO_2526 (O_2526,N_29767,N_29800);
nand UO_2527 (O_2527,N_29733,N_29962);
nor UO_2528 (O_2528,N_29792,N_29911);
or UO_2529 (O_2529,N_29890,N_29741);
and UO_2530 (O_2530,N_29783,N_29994);
nand UO_2531 (O_2531,N_29882,N_29816);
xnor UO_2532 (O_2532,N_29939,N_29974);
and UO_2533 (O_2533,N_29758,N_29725);
xor UO_2534 (O_2534,N_29932,N_29807);
nor UO_2535 (O_2535,N_29925,N_29998);
xor UO_2536 (O_2536,N_29749,N_29766);
nor UO_2537 (O_2537,N_29833,N_29775);
nor UO_2538 (O_2538,N_29965,N_29982);
nor UO_2539 (O_2539,N_29928,N_29899);
and UO_2540 (O_2540,N_29859,N_29728);
nand UO_2541 (O_2541,N_29934,N_29797);
nor UO_2542 (O_2542,N_29754,N_29705);
nand UO_2543 (O_2543,N_29934,N_29779);
nor UO_2544 (O_2544,N_29727,N_29828);
or UO_2545 (O_2545,N_29768,N_29846);
xor UO_2546 (O_2546,N_29801,N_29728);
xor UO_2547 (O_2547,N_29755,N_29953);
and UO_2548 (O_2548,N_29796,N_29713);
nor UO_2549 (O_2549,N_29707,N_29747);
nor UO_2550 (O_2550,N_29967,N_29992);
nor UO_2551 (O_2551,N_29713,N_29980);
nor UO_2552 (O_2552,N_29957,N_29978);
xnor UO_2553 (O_2553,N_29768,N_29944);
xor UO_2554 (O_2554,N_29808,N_29875);
nor UO_2555 (O_2555,N_29728,N_29931);
nor UO_2556 (O_2556,N_29943,N_29969);
xor UO_2557 (O_2557,N_29872,N_29736);
xor UO_2558 (O_2558,N_29841,N_29866);
xnor UO_2559 (O_2559,N_29709,N_29865);
nand UO_2560 (O_2560,N_29906,N_29965);
nor UO_2561 (O_2561,N_29976,N_29816);
or UO_2562 (O_2562,N_29995,N_29917);
and UO_2563 (O_2563,N_29821,N_29752);
or UO_2564 (O_2564,N_29818,N_29998);
or UO_2565 (O_2565,N_29935,N_29973);
nand UO_2566 (O_2566,N_29905,N_29735);
nand UO_2567 (O_2567,N_29963,N_29711);
and UO_2568 (O_2568,N_29937,N_29776);
nor UO_2569 (O_2569,N_29810,N_29851);
nand UO_2570 (O_2570,N_29931,N_29857);
xnor UO_2571 (O_2571,N_29856,N_29918);
and UO_2572 (O_2572,N_29926,N_29896);
nand UO_2573 (O_2573,N_29755,N_29969);
xor UO_2574 (O_2574,N_29885,N_29841);
and UO_2575 (O_2575,N_29923,N_29993);
and UO_2576 (O_2576,N_29850,N_29845);
and UO_2577 (O_2577,N_29875,N_29754);
or UO_2578 (O_2578,N_29916,N_29731);
and UO_2579 (O_2579,N_29950,N_29999);
xnor UO_2580 (O_2580,N_29833,N_29982);
nor UO_2581 (O_2581,N_29723,N_29744);
xnor UO_2582 (O_2582,N_29809,N_29877);
and UO_2583 (O_2583,N_29834,N_29934);
nor UO_2584 (O_2584,N_29791,N_29931);
or UO_2585 (O_2585,N_29917,N_29926);
and UO_2586 (O_2586,N_29795,N_29724);
nor UO_2587 (O_2587,N_29877,N_29828);
nor UO_2588 (O_2588,N_29938,N_29960);
nand UO_2589 (O_2589,N_29938,N_29810);
or UO_2590 (O_2590,N_29748,N_29954);
nand UO_2591 (O_2591,N_29911,N_29963);
or UO_2592 (O_2592,N_29907,N_29875);
nand UO_2593 (O_2593,N_29785,N_29921);
and UO_2594 (O_2594,N_29718,N_29916);
xor UO_2595 (O_2595,N_29947,N_29833);
and UO_2596 (O_2596,N_29802,N_29898);
and UO_2597 (O_2597,N_29739,N_29967);
and UO_2598 (O_2598,N_29890,N_29957);
nand UO_2599 (O_2599,N_29933,N_29770);
nor UO_2600 (O_2600,N_29868,N_29993);
nor UO_2601 (O_2601,N_29992,N_29763);
and UO_2602 (O_2602,N_29809,N_29876);
nand UO_2603 (O_2603,N_29853,N_29709);
nand UO_2604 (O_2604,N_29943,N_29764);
nor UO_2605 (O_2605,N_29809,N_29957);
nand UO_2606 (O_2606,N_29925,N_29817);
nand UO_2607 (O_2607,N_29910,N_29828);
or UO_2608 (O_2608,N_29704,N_29713);
xnor UO_2609 (O_2609,N_29964,N_29825);
or UO_2610 (O_2610,N_29946,N_29982);
nor UO_2611 (O_2611,N_29717,N_29885);
or UO_2612 (O_2612,N_29752,N_29761);
and UO_2613 (O_2613,N_29901,N_29731);
xor UO_2614 (O_2614,N_29861,N_29907);
nand UO_2615 (O_2615,N_29906,N_29822);
and UO_2616 (O_2616,N_29976,N_29975);
and UO_2617 (O_2617,N_29746,N_29882);
xnor UO_2618 (O_2618,N_29959,N_29886);
and UO_2619 (O_2619,N_29849,N_29847);
nor UO_2620 (O_2620,N_29854,N_29925);
xnor UO_2621 (O_2621,N_29710,N_29989);
and UO_2622 (O_2622,N_29980,N_29704);
and UO_2623 (O_2623,N_29724,N_29944);
and UO_2624 (O_2624,N_29737,N_29869);
nor UO_2625 (O_2625,N_29767,N_29887);
or UO_2626 (O_2626,N_29946,N_29729);
nand UO_2627 (O_2627,N_29920,N_29748);
nor UO_2628 (O_2628,N_29976,N_29895);
and UO_2629 (O_2629,N_29784,N_29859);
nand UO_2630 (O_2630,N_29909,N_29794);
nand UO_2631 (O_2631,N_29924,N_29837);
or UO_2632 (O_2632,N_29770,N_29915);
and UO_2633 (O_2633,N_29780,N_29927);
and UO_2634 (O_2634,N_29716,N_29831);
and UO_2635 (O_2635,N_29997,N_29865);
nand UO_2636 (O_2636,N_29772,N_29754);
or UO_2637 (O_2637,N_29817,N_29752);
xor UO_2638 (O_2638,N_29755,N_29747);
and UO_2639 (O_2639,N_29733,N_29916);
and UO_2640 (O_2640,N_29758,N_29844);
nor UO_2641 (O_2641,N_29897,N_29839);
nor UO_2642 (O_2642,N_29734,N_29777);
and UO_2643 (O_2643,N_29974,N_29824);
and UO_2644 (O_2644,N_29759,N_29890);
nand UO_2645 (O_2645,N_29803,N_29847);
nor UO_2646 (O_2646,N_29892,N_29991);
xnor UO_2647 (O_2647,N_29813,N_29787);
nand UO_2648 (O_2648,N_29751,N_29935);
xor UO_2649 (O_2649,N_29974,N_29852);
nor UO_2650 (O_2650,N_29730,N_29807);
xnor UO_2651 (O_2651,N_29868,N_29751);
nand UO_2652 (O_2652,N_29782,N_29700);
and UO_2653 (O_2653,N_29737,N_29867);
nand UO_2654 (O_2654,N_29917,N_29732);
nor UO_2655 (O_2655,N_29843,N_29929);
nand UO_2656 (O_2656,N_29728,N_29905);
nor UO_2657 (O_2657,N_29793,N_29792);
and UO_2658 (O_2658,N_29802,N_29716);
nor UO_2659 (O_2659,N_29758,N_29726);
or UO_2660 (O_2660,N_29835,N_29876);
or UO_2661 (O_2661,N_29937,N_29980);
nand UO_2662 (O_2662,N_29775,N_29912);
nor UO_2663 (O_2663,N_29857,N_29882);
xnor UO_2664 (O_2664,N_29792,N_29908);
nand UO_2665 (O_2665,N_29814,N_29967);
and UO_2666 (O_2666,N_29743,N_29919);
and UO_2667 (O_2667,N_29996,N_29933);
xnor UO_2668 (O_2668,N_29783,N_29796);
nand UO_2669 (O_2669,N_29999,N_29877);
nand UO_2670 (O_2670,N_29735,N_29813);
nand UO_2671 (O_2671,N_29914,N_29993);
nand UO_2672 (O_2672,N_29934,N_29828);
or UO_2673 (O_2673,N_29905,N_29746);
nand UO_2674 (O_2674,N_29901,N_29722);
nand UO_2675 (O_2675,N_29754,N_29813);
nor UO_2676 (O_2676,N_29717,N_29722);
and UO_2677 (O_2677,N_29805,N_29940);
nand UO_2678 (O_2678,N_29700,N_29737);
xor UO_2679 (O_2679,N_29789,N_29726);
or UO_2680 (O_2680,N_29797,N_29823);
xnor UO_2681 (O_2681,N_29772,N_29863);
nand UO_2682 (O_2682,N_29798,N_29845);
or UO_2683 (O_2683,N_29914,N_29833);
nand UO_2684 (O_2684,N_29794,N_29887);
or UO_2685 (O_2685,N_29718,N_29784);
nor UO_2686 (O_2686,N_29803,N_29969);
xnor UO_2687 (O_2687,N_29721,N_29775);
or UO_2688 (O_2688,N_29770,N_29775);
or UO_2689 (O_2689,N_29911,N_29749);
or UO_2690 (O_2690,N_29999,N_29994);
xnor UO_2691 (O_2691,N_29804,N_29993);
nand UO_2692 (O_2692,N_29715,N_29899);
and UO_2693 (O_2693,N_29846,N_29911);
and UO_2694 (O_2694,N_29866,N_29879);
or UO_2695 (O_2695,N_29918,N_29939);
nand UO_2696 (O_2696,N_29966,N_29878);
nor UO_2697 (O_2697,N_29726,N_29925);
or UO_2698 (O_2698,N_29976,N_29855);
nand UO_2699 (O_2699,N_29985,N_29794);
nand UO_2700 (O_2700,N_29846,N_29887);
nand UO_2701 (O_2701,N_29837,N_29811);
nor UO_2702 (O_2702,N_29831,N_29708);
or UO_2703 (O_2703,N_29736,N_29912);
or UO_2704 (O_2704,N_29873,N_29852);
or UO_2705 (O_2705,N_29776,N_29819);
and UO_2706 (O_2706,N_29873,N_29989);
nor UO_2707 (O_2707,N_29885,N_29945);
nand UO_2708 (O_2708,N_29950,N_29979);
and UO_2709 (O_2709,N_29934,N_29911);
nor UO_2710 (O_2710,N_29803,N_29715);
nand UO_2711 (O_2711,N_29734,N_29787);
nand UO_2712 (O_2712,N_29875,N_29788);
xor UO_2713 (O_2713,N_29870,N_29849);
nor UO_2714 (O_2714,N_29758,N_29976);
nor UO_2715 (O_2715,N_29881,N_29700);
xor UO_2716 (O_2716,N_29791,N_29971);
nor UO_2717 (O_2717,N_29989,N_29958);
and UO_2718 (O_2718,N_29795,N_29887);
and UO_2719 (O_2719,N_29793,N_29706);
nor UO_2720 (O_2720,N_29744,N_29742);
xnor UO_2721 (O_2721,N_29952,N_29721);
nand UO_2722 (O_2722,N_29960,N_29889);
or UO_2723 (O_2723,N_29744,N_29855);
nor UO_2724 (O_2724,N_29886,N_29929);
nor UO_2725 (O_2725,N_29955,N_29720);
or UO_2726 (O_2726,N_29738,N_29764);
nor UO_2727 (O_2727,N_29980,N_29925);
and UO_2728 (O_2728,N_29832,N_29750);
nor UO_2729 (O_2729,N_29839,N_29790);
and UO_2730 (O_2730,N_29910,N_29905);
xnor UO_2731 (O_2731,N_29711,N_29764);
nand UO_2732 (O_2732,N_29787,N_29731);
or UO_2733 (O_2733,N_29868,N_29785);
xnor UO_2734 (O_2734,N_29892,N_29819);
or UO_2735 (O_2735,N_29958,N_29722);
nand UO_2736 (O_2736,N_29829,N_29993);
or UO_2737 (O_2737,N_29880,N_29870);
nor UO_2738 (O_2738,N_29886,N_29885);
or UO_2739 (O_2739,N_29749,N_29838);
or UO_2740 (O_2740,N_29998,N_29922);
nand UO_2741 (O_2741,N_29790,N_29823);
xnor UO_2742 (O_2742,N_29946,N_29820);
or UO_2743 (O_2743,N_29766,N_29930);
xnor UO_2744 (O_2744,N_29916,N_29820);
xor UO_2745 (O_2745,N_29948,N_29943);
nor UO_2746 (O_2746,N_29937,N_29907);
or UO_2747 (O_2747,N_29907,N_29730);
nor UO_2748 (O_2748,N_29794,N_29928);
or UO_2749 (O_2749,N_29853,N_29885);
and UO_2750 (O_2750,N_29722,N_29863);
and UO_2751 (O_2751,N_29742,N_29795);
nor UO_2752 (O_2752,N_29730,N_29859);
xnor UO_2753 (O_2753,N_29948,N_29759);
nand UO_2754 (O_2754,N_29759,N_29799);
xnor UO_2755 (O_2755,N_29708,N_29878);
nand UO_2756 (O_2756,N_29912,N_29738);
or UO_2757 (O_2757,N_29954,N_29826);
and UO_2758 (O_2758,N_29781,N_29980);
xnor UO_2759 (O_2759,N_29729,N_29967);
or UO_2760 (O_2760,N_29800,N_29974);
and UO_2761 (O_2761,N_29856,N_29905);
nor UO_2762 (O_2762,N_29986,N_29854);
and UO_2763 (O_2763,N_29815,N_29832);
nor UO_2764 (O_2764,N_29748,N_29730);
xor UO_2765 (O_2765,N_29780,N_29782);
xnor UO_2766 (O_2766,N_29843,N_29739);
and UO_2767 (O_2767,N_29993,N_29831);
or UO_2768 (O_2768,N_29871,N_29949);
xor UO_2769 (O_2769,N_29853,N_29989);
xnor UO_2770 (O_2770,N_29720,N_29873);
nand UO_2771 (O_2771,N_29894,N_29973);
or UO_2772 (O_2772,N_29845,N_29740);
nand UO_2773 (O_2773,N_29969,N_29831);
and UO_2774 (O_2774,N_29911,N_29756);
xnor UO_2775 (O_2775,N_29993,N_29793);
nor UO_2776 (O_2776,N_29904,N_29781);
xor UO_2777 (O_2777,N_29746,N_29809);
xor UO_2778 (O_2778,N_29928,N_29995);
nor UO_2779 (O_2779,N_29860,N_29939);
nand UO_2780 (O_2780,N_29879,N_29785);
nor UO_2781 (O_2781,N_29916,N_29875);
xnor UO_2782 (O_2782,N_29791,N_29976);
or UO_2783 (O_2783,N_29742,N_29905);
xor UO_2784 (O_2784,N_29941,N_29714);
nand UO_2785 (O_2785,N_29863,N_29834);
nand UO_2786 (O_2786,N_29996,N_29810);
nor UO_2787 (O_2787,N_29981,N_29835);
xnor UO_2788 (O_2788,N_29756,N_29913);
or UO_2789 (O_2789,N_29804,N_29829);
or UO_2790 (O_2790,N_29746,N_29764);
nor UO_2791 (O_2791,N_29891,N_29768);
and UO_2792 (O_2792,N_29914,N_29983);
xnor UO_2793 (O_2793,N_29770,N_29981);
or UO_2794 (O_2794,N_29736,N_29744);
and UO_2795 (O_2795,N_29713,N_29901);
nand UO_2796 (O_2796,N_29830,N_29717);
and UO_2797 (O_2797,N_29785,N_29732);
nor UO_2798 (O_2798,N_29906,N_29828);
and UO_2799 (O_2799,N_29733,N_29881);
xnor UO_2800 (O_2800,N_29833,N_29799);
and UO_2801 (O_2801,N_29722,N_29846);
or UO_2802 (O_2802,N_29788,N_29742);
or UO_2803 (O_2803,N_29765,N_29812);
or UO_2804 (O_2804,N_29737,N_29842);
or UO_2805 (O_2805,N_29707,N_29999);
nand UO_2806 (O_2806,N_29801,N_29792);
and UO_2807 (O_2807,N_29982,N_29974);
xnor UO_2808 (O_2808,N_29974,N_29742);
nand UO_2809 (O_2809,N_29872,N_29799);
nand UO_2810 (O_2810,N_29892,N_29839);
nor UO_2811 (O_2811,N_29816,N_29974);
or UO_2812 (O_2812,N_29797,N_29775);
and UO_2813 (O_2813,N_29971,N_29835);
nand UO_2814 (O_2814,N_29996,N_29731);
nand UO_2815 (O_2815,N_29847,N_29808);
nand UO_2816 (O_2816,N_29858,N_29965);
or UO_2817 (O_2817,N_29913,N_29815);
or UO_2818 (O_2818,N_29724,N_29767);
or UO_2819 (O_2819,N_29825,N_29888);
and UO_2820 (O_2820,N_29868,N_29978);
or UO_2821 (O_2821,N_29753,N_29712);
and UO_2822 (O_2822,N_29728,N_29838);
nand UO_2823 (O_2823,N_29777,N_29957);
and UO_2824 (O_2824,N_29933,N_29716);
nand UO_2825 (O_2825,N_29861,N_29989);
xnor UO_2826 (O_2826,N_29975,N_29880);
or UO_2827 (O_2827,N_29862,N_29797);
nand UO_2828 (O_2828,N_29981,N_29767);
nand UO_2829 (O_2829,N_29997,N_29984);
xnor UO_2830 (O_2830,N_29826,N_29980);
nand UO_2831 (O_2831,N_29978,N_29830);
xor UO_2832 (O_2832,N_29864,N_29774);
nand UO_2833 (O_2833,N_29903,N_29917);
nand UO_2834 (O_2834,N_29821,N_29882);
or UO_2835 (O_2835,N_29800,N_29780);
or UO_2836 (O_2836,N_29807,N_29856);
xor UO_2837 (O_2837,N_29939,N_29890);
xor UO_2838 (O_2838,N_29929,N_29810);
nor UO_2839 (O_2839,N_29853,N_29758);
xnor UO_2840 (O_2840,N_29737,N_29858);
or UO_2841 (O_2841,N_29735,N_29861);
or UO_2842 (O_2842,N_29716,N_29818);
nand UO_2843 (O_2843,N_29909,N_29977);
nor UO_2844 (O_2844,N_29804,N_29714);
nand UO_2845 (O_2845,N_29812,N_29835);
nand UO_2846 (O_2846,N_29776,N_29744);
nor UO_2847 (O_2847,N_29908,N_29919);
xor UO_2848 (O_2848,N_29996,N_29980);
and UO_2849 (O_2849,N_29937,N_29963);
and UO_2850 (O_2850,N_29884,N_29706);
nand UO_2851 (O_2851,N_29937,N_29749);
nand UO_2852 (O_2852,N_29834,N_29844);
nand UO_2853 (O_2853,N_29865,N_29966);
or UO_2854 (O_2854,N_29700,N_29942);
nand UO_2855 (O_2855,N_29935,N_29945);
xor UO_2856 (O_2856,N_29751,N_29987);
or UO_2857 (O_2857,N_29710,N_29790);
or UO_2858 (O_2858,N_29933,N_29965);
xor UO_2859 (O_2859,N_29967,N_29708);
nor UO_2860 (O_2860,N_29708,N_29844);
nand UO_2861 (O_2861,N_29971,N_29910);
and UO_2862 (O_2862,N_29973,N_29960);
and UO_2863 (O_2863,N_29767,N_29872);
and UO_2864 (O_2864,N_29848,N_29929);
xor UO_2865 (O_2865,N_29971,N_29770);
nand UO_2866 (O_2866,N_29747,N_29872);
xor UO_2867 (O_2867,N_29937,N_29754);
xnor UO_2868 (O_2868,N_29712,N_29883);
or UO_2869 (O_2869,N_29826,N_29922);
nand UO_2870 (O_2870,N_29977,N_29811);
and UO_2871 (O_2871,N_29976,N_29903);
nor UO_2872 (O_2872,N_29994,N_29706);
or UO_2873 (O_2873,N_29700,N_29924);
and UO_2874 (O_2874,N_29826,N_29953);
and UO_2875 (O_2875,N_29915,N_29755);
nor UO_2876 (O_2876,N_29724,N_29830);
nor UO_2877 (O_2877,N_29841,N_29784);
nand UO_2878 (O_2878,N_29928,N_29921);
or UO_2879 (O_2879,N_29963,N_29842);
and UO_2880 (O_2880,N_29813,N_29803);
and UO_2881 (O_2881,N_29849,N_29734);
nand UO_2882 (O_2882,N_29806,N_29931);
xnor UO_2883 (O_2883,N_29779,N_29816);
nor UO_2884 (O_2884,N_29753,N_29907);
or UO_2885 (O_2885,N_29931,N_29902);
nand UO_2886 (O_2886,N_29848,N_29704);
and UO_2887 (O_2887,N_29808,N_29932);
nand UO_2888 (O_2888,N_29835,N_29907);
and UO_2889 (O_2889,N_29936,N_29961);
and UO_2890 (O_2890,N_29961,N_29756);
or UO_2891 (O_2891,N_29915,N_29709);
nand UO_2892 (O_2892,N_29947,N_29979);
and UO_2893 (O_2893,N_29742,N_29972);
nor UO_2894 (O_2894,N_29779,N_29872);
xnor UO_2895 (O_2895,N_29849,N_29772);
nand UO_2896 (O_2896,N_29857,N_29955);
xor UO_2897 (O_2897,N_29946,N_29781);
or UO_2898 (O_2898,N_29859,N_29925);
and UO_2899 (O_2899,N_29843,N_29908);
and UO_2900 (O_2900,N_29998,N_29931);
nand UO_2901 (O_2901,N_29870,N_29861);
nand UO_2902 (O_2902,N_29939,N_29781);
xor UO_2903 (O_2903,N_29880,N_29926);
nor UO_2904 (O_2904,N_29894,N_29852);
nand UO_2905 (O_2905,N_29721,N_29895);
nor UO_2906 (O_2906,N_29912,N_29755);
nand UO_2907 (O_2907,N_29953,N_29945);
and UO_2908 (O_2908,N_29786,N_29798);
nor UO_2909 (O_2909,N_29815,N_29972);
or UO_2910 (O_2910,N_29734,N_29739);
nor UO_2911 (O_2911,N_29960,N_29892);
nand UO_2912 (O_2912,N_29791,N_29797);
nand UO_2913 (O_2913,N_29788,N_29988);
xnor UO_2914 (O_2914,N_29713,N_29817);
nor UO_2915 (O_2915,N_29884,N_29751);
xnor UO_2916 (O_2916,N_29829,N_29950);
nor UO_2917 (O_2917,N_29776,N_29781);
or UO_2918 (O_2918,N_29777,N_29771);
nand UO_2919 (O_2919,N_29985,N_29991);
or UO_2920 (O_2920,N_29846,N_29996);
and UO_2921 (O_2921,N_29914,N_29786);
nor UO_2922 (O_2922,N_29704,N_29855);
nor UO_2923 (O_2923,N_29922,N_29731);
xor UO_2924 (O_2924,N_29901,N_29708);
and UO_2925 (O_2925,N_29997,N_29906);
xor UO_2926 (O_2926,N_29750,N_29773);
xnor UO_2927 (O_2927,N_29985,N_29712);
or UO_2928 (O_2928,N_29889,N_29996);
nor UO_2929 (O_2929,N_29960,N_29828);
xnor UO_2930 (O_2930,N_29857,N_29879);
nor UO_2931 (O_2931,N_29920,N_29710);
xor UO_2932 (O_2932,N_29729,N_29876);
nor UO_2933 (O_2933,N_29918,N_29766);
nor UO_2934 (O_2934,N_29703,N_29837);
and UO_2935 (O_2935,N_29790,N_29792);
or UO_2936 (O_2936,N_29927,N_29944);
nor UO_2937 (O_2937,N_29854,N_29726);
nand UO_2938 (O_2938,N_29757,N_29986);
or UO_2939 (O_2939,N_29726,N_29822);
or UO_2940 (O_2940,N_29981,N_29756);
or UO_2941 (O_2941,N_29707,N_29894);
xor UO_2942 (O_2942,N_29805,N_29711);
nand UO_2943 (O_2943,N_29845,N_29883);
or UO_2944 (O_2944,N_29968,N_29782);
nor UO_2945 (O_2945,N_29906,N_29879);
nand UO_2946 (O_2946,N_29765,N_29712);
and UO_2947 (O_2947,N_29791,N_29927);
nand UO_2948 (O_2948,N_29765,N_29856);
nor UO_2949 (O_2949,N_29918,N_29805);
nor UO_2950 (O_2950,N_29737,N_29777);
nor UO_2951 (O_2951,N_29744,N_29946);
nor UO_2952 (O_2952,N_29987,N_29721);
and UO_2953 (O_2953,N_29827,N_29823);
nand UO_2954 (O_2954,N_29774,N_29916);
or UO_2955 (O_2955,N_29725,N_29848);
or UO_2956 (O_2956,N_29929,N_29760);
xor UO_2957 (O_2957,N_29957,N_29892);
and UO_2958 (O_2958,N_29855,N_29850);
xnor UO_2959 (O_2959,N_29985,N_29950);
nand UO_2960 (O_2960,N_29929,N_29905);
or UO_2961 (O_2961,N_29702,N_29966);
nor UO_2962 (O_2962,N_29914,N_29957);
nor UO_2963 (O_2963,N_29917,N_29833);
xor UO_2964 (O_2964,N_29895,N_29838);
or UO_2965 (O_2965,N_29727,N_29978);
and UO_2966 (O_2966,N_29870,N_29902);
nand UO_2967 (O_2967,N_29910,N_29923);
or UO_2968 (O_2968,N_29700,N_29973);
xor UO_2969 (O_2969,N_29742,N_29913);
or UO_2970 (O_2970,N_29994,N_29749);
nand UO_2971 (O_2971,N_29750,N_29715);
xor UO_2972 (O_2972,N_29719,N_29815);
and UO_2973 (O_2973,N_29766,N_29828);
nand UO_2974 (O_2974,N_29710,N_29958);
and UO_2975 (O_2975,N_29960,N_29749);
nor UO_2976 (O_2976,N_29861,N_29812);
or UO_2977 (O_2977,N_29846,N_29753);
xor UO_2978 (O_2978,N_29734,N_29934);
nand UO_2979 (O_2979,N_29839,N_29933);
and UO_2980 (O_2980,N_29789,N_29893);
nand UO_2981 (O_2981,N_29861,N_29992);
or UO_2982 (O_2982,N_29763,N_29719);
nand UO_2983 (O_2983,N_29964,N_29977);
and UO_2984 (O_2984,N_29794,N_29719);
nand UO_2985 (O_2985,N_29849,N_29941);
or UO_2986 (O_2986,N_29772,N_29926);
and UO_2987 (O_2987,N_29845,N_29937);
and UO_2988 (O_2988,N_29947,N_29993);
xor UO_2989 (O_2989,N_29743,N_29963);
xor UO_2990 (O_2990,N_29984,N_29846);
xor UO_2991 (O_2991,N_29851,N_29884);
xnor UO_2992 (O_2992,N_29965,N_29950);
nand UO_2993 (O_2993,N_29937,N_29855);
nand UO_2994 (O_2994,N_29740,N_29757);
and UO_2995 (O_2995,N_29842,N_29837);
or UO_2996 (O_2996,N_29848,N_29777);
nand UO_2997 (O_2997,N_29969,N_29985);
or UO_2998 (O_2998,N_29993,N_29964);
nand UO_2999 (O_2999,N_29753,N_29876);
nand UO_3000 (O_3000,N_29973,N_29849);
and UO_3001 (O_3001,N_29798,N_29828);
xor UO_3002 (O_3002,N_29963,N_29791);
or UO_3003 (O_3003,N_29976,N_29972);
nor UO_3004 (O_3004,N_29954,N_29796);
nor UO_3005 (O_3005,N_29873,N_29871);
xnor UO_3006 (O_3006,N_29798,N_29849);
or UO_3007 (O_3007,N_29782,N_29871);
nand UO_3008 (O_3008,N_29926,N_29868);
or UO_3009 (O_3009,N_29710,N_29723);
nand UO_3010 (O_3010,N_29791,N_29775);
xnor UO_3011 (O_3011,N_29944,N_29721);
nor UO_3012 (O_3012,N_29855,N_29767);
xnor UO_3013 (O_3013,N_29722,N_29857);
or UO_3014 (O_3014,N_29795,N_29876);
nand UO_3015 (O_3015,N_29900,N_29862);
and UO_3016 (O_3016,N_29726,N_29830);
xnor UO_3017 (O_3017,N_29756,N_29998);
or UO_3018 (O_3018,N_29852,N_29848);
and UO_3019 (O_3019,N_29922,N_29901);
nor UO_3020 (O_3020,N_29841,N_29984);
or UO_3021 (O_3021,N_29891,N_29731);
xnor UO_3022 (O_3022,N_29858,N_29981);
and UO_3023 (O_3023,N_29738,N_29982);
and UO_3024 (O_3024,N_29708,N_29738);
nand UO_3025 (O_3025,N_29708,N_29907);
or UO_3026 (O_3026,N_29971,N_29749);
and UO_3027 (O_3027,N_29714,N_29867);
nor UO_3028 (O_3028,N_29795,N_29763);
nand UO_3029 (O_3029,N_29869,N_29852);
xnor UO_3030 (O_3030,N_29929,N_29984);
and UO_3031 (O_3031,N_29878,N_29811);
or UO_3032 (O_3032,N_29749,N_29713);
or UO_3033 (O_3033,N_29810,N_29937);
and UO_3034 (O_3034,N_29819,N_29903);
or UO_3035 (O_3035,N_29929,N_29931);
xnor UO_3036 (O_3036,N_29837,N_29830);
and UO_3037 (O_3037,N_29859,N_29973);
xnor UO_3038 (O_3038,N_29774,N_29939);
and UO_3039 (O_3039,N_29829,N_29940);
or UO_3040 (O_3040,N_29709,N_29896);
nand UO_3041 (O_3041,N_29999,N_29926);
and UO_3042 (O_3042,N_29742,N_29801);
nor UO_3043 (O_3043,N_29925,N_29785);
nand UO_3044 (O_3044,N_29733,N_29785);
or UO_3045 (O_3045,N_29906,N_29733);
nor UO_3046 (O_3046,N_29995,N_29785);
nand UO_3047 (O_3047,N_29955,N_29938);
or UO_3048 (O_3048,N_29828,N_29712);
nor UO_3049 (O_3049,N_29949,N_29773);
xor UO_3050 (O_3050,N_29963,N_29778);
and UO_3051 (O_3051,N_29771,N_29719);
and UO_3052 (O_3052,N_29964,N_29992);
nand UO_3053 (O_3053,N_29940,N_29830);
xor UO_3054 (O_3054,N_29909,N_29808);
or UO_3055 (O_3055,N_29829,N_29702);
nor UO_3056 (O_3056,N_29919,N_29925);
xor UO_3057 (O_3057,N_29959,N_29969);
xor UO_3058 (O_3058,N_29807,N_29966);
xnor UO_3059 (O_3059,N_29774,N_29980);
xor UO_3060 (O_3060,N_29706,N_29925);
nor UO_3061 (O_3061,N_29726,N_29842);
xor UO_3062 (O_3062,N_29911,N_29981);
or UO_3063 (O_3063,N_29892,N_29949);
nand UO_3064 (O_3064,N_29902,N_29968);
and UO_3065 (O_3065,N_29926,N_29912);
and UO_3066 (O_3066,N_29830,N_29805);
nand UO_3067 (O_3067,N_29825,N_29907);
and UO_3068 (O_3068,N_29735,N_29781);
and UO_3069 (O_3069,N_29986,N_29892);
or UO_3070 (O_3070,N_29941,N_29801);
and UO_3071 (O_3071,N_29818,N_29842);
or UO_3072 (O_3072,N_29806,N_29959);
xnor UO_3073 (O_3073,N_29986,N_29816);
and UO_3074 (O_3074,N_29984,N_29765);
and UO_3075 (O_3075,N_29829,N_29746);
xnor UO_3076 (O_3076,N_29733,N_29942);
nand UO_3077 (O_3077,N_29762,N_29939);
xnor UO_3078 (O_3078,N_29945,N_29794);
or UO_3079 (O_3079,N_29843,N_29815);
xnor UO_3080 (O_3080,N_29973,N_29720);
nand UO_3081 (O_3081,N_29894,N_29947);
and UO_3082 (O_3082,N_29951,N_29952);
and UO_3083 (O_3083,N_29824,N_29962);
xor UO_3084 (O_3084,N_29808,N_29726);
nand UO_3085 (O_3085,N_29929,N_29889);
nand UO_3086 (O_3086,N_29930,N_29974);
or UO_3087 (O_3087,N_29926,N_29930);
or UO_3088 (O_3088,N_29840,N_29828);
or UO_3089 (O_3089,N_29920,N_29984);
nor UO_3090 (O_3090,N_29743,N_29734);
nand UO_3091 (O_3091,N_29871,N_29906);
xnor UO_3092 (O_3092,N_29920,N_29852);
nor UO_3093 (O_3093,N_29732,N_29843);
nand UO_3094 (O_3094,N_29795,N_29991);
nor UO_3095 (O_3095,N_29885,N_29874);
xor UO_3096 (O_3096,N_29813,N_29926);
nand UO_3097 (O_3097,N_29900,N_29980);
or UO_3098 (O_3098,N_29983,N_29896);
xor UO_3099 (O_3099,N_29867,N_29882);
nand UO_3100 (O_3100,N_29896,N_29734);
and UO_3101 (O_3101,N_29984,N_29837);
nand UO_3102 (O_3102,N_29913,N_29935);
or UO_3103 (O_3103,N_29792,N_29963);
or UO_3104 (O_3104,N_29712,N_29960);
or UO_3105 (O_3105,N_29776,N_29729);
nor UO_3106 (O_3106,N_29718,N_29755);
xor UO_3107 (O_3107,N_29947,N_29803);
nor UO_3108 (O_3108,N_29980,N_29982);
nand UO_3109 (O_3109,N_29758,N_29738);
nand UO_3110 (O_3110,N_29884,N_29883);
nand UO_3111 (O_3111,N_29979,N_29956);
or UO_3112 (O_3112,N_29943,N_29995);
and UO_3113 (O_3113,N_29701,N_29791);
xnor UO_3114 (O_3114,N_29986,N_29884);
nor UO_3115 (O_3115,N_29794,N_29818);
and UO_3116 (O_3116,N_29768,N_29838);
or UO_3117 (O_3117,N_29939,N_29883);
nand UO_3118 (O_3118,N_29784,N_29710);
nand UO_3119 (O_3119,N_29848,N_29809);
xnor UO_3120 (O_3120,N_29758,N_29989);
nand UO_3121 (O_3121,N_29760,N_29825);
and UO_3122 (O_3122,N_29777,N_29864);
xor UO_3123 (O_3123,N_29967,N_29752);
nor UO_3124 (O_3124,N_29910,N_29919);
nand UO_3125 (O_3125,N_29796,N_29822);
nor UO_3126 (O_3126,N_29914,N_29925);
or UO_3127 (O_3127,N_29751,N_29775);
nand UO_3128 (O_3128,N_29939,N_29745);
nand UO_3129 (O_3129,N_29772,N_29968);
xor UO_3130 (O_3130,N_29742,N_29833);
nand UO_3131 (O_3131,N_29897,N_29830);
and UO_3132 (O_3132,N_29946,N_29901);
nor UO_3133 (O_3133,N_29810,N_29876);
nand UO_3134 (O_3134,N_29925,N_29814);
or UO_3135 (O_3135,N_29705,N_29715);
xor UO_3136 (O_3136,N_29708,N_29981);
or UO_3137 (O_3137,N_29865,N_29943);
and UO_3138 (O_3138,N_29826,N_29718);
or UO_3139 (O_3139,N_29805,N_29997);
nand UO_3140 (O_3140,N_29780,N_29762);
and UO_3141 (O_3141,N_29798,N_29909);
nand UO_3142 (O_3142,N_29733,N_29989);
xnor UO_3143 (O_3143,N_29782,N_29961);
or UO_3144 (O_3144,N_29867,N_29775);
nor UO_3145 (O_3145,N_29863,N_29830);
xnor UO_3146 (O_3146,N_29731,N_29894);
and UO_3147 (O_3147,N_29702,N_29980);
or UO_3148 (O_3148,N_29923,N_29720);
and UO_3149 (O_3149,N_29811,N_29934);
nand UO_3150 (O_3150,N_29728,N_29966);
or UO_3151 (O_3151,N_29749,N_29921);
and UO_3152 (O_3152,N_29795,N_29818);
nor UO_3153 (O_3153,N_29978,N_29754);
nor UO_3154 (O_3154,N_29905,N_29924);
or UO_3155 (O_3155,N_29953,N_29741);
xor UO_3156 (O_3156,N_29985,N_29702);
nor UO_3157 (O_3157,N_29749,N_29796);
xnor UO_3158 (O_3158,N_29766,N_29717);
nor UO_3159 (O_3159,N_29735,N_29749);
nand UO_3160 (O_3160,N_29953,N_29986);
or UO_3161 (O_3161,N_29969,N_29728);
or UO_3162 (O_3162,N_29893,N_29970);
or UO_3163 (O_3163,N_29751,N_29770);
and UO_3164 (O_3164,N_29833,N_29970);
nor UO_3165 (O_3165,N_29761,N_29773);
xnor UO_3166 (O_3166,N_29916,N_29745);
nand UO_3167 (O_3167,N_29777,N_29720);
and UO_3168 (O_3168,N_29941,N_29737);
nand UO_3169 (O_3169,N_29822,N_29968);
xor UO_3170 (O_3170,N_29964,N_29922);
xnor UO_3171 (O_3171,N_29967,N_29954);
nor UO_3172 (O_3172,N_29924,N_29935);
xnor UO_3173 (O_3173,N_29720,N_29879);
or UO_3174 (O_3174,N_29888,N_29757);
xnor UO_3175 (O_3175,N_29719,N_29897);
nor UO_3176 (O_3176,N_29729,N_29906);
xnor UO_3177 (O_3177,N_29903,N_29896);
xnor UO_3178 (O_3178,N_29897,N_29994);
and UO_3179 (O_3179,N_29856,N_29834);
nand UO_3180 (O_3180,N_29761,N_29751);
nand UO_3181 (O_3181,N_29937,N_29894);
and UO_3182 (O_3182,N_29750,N_29771);
nand UO_3183 (O_3183,N_29756,N_29748);
nor UO_3184 (O_3184,N_29807,N_29939);
nor UO_3185 (O_3185,N_29969,N_29715);
nor UO_3186 (O_3186,N_29737,N_29953);
or UO_3187 (O_3187,N_29833,N_29806);
nand UO_3188 (O_3188,N_29787,N_29964);
or UO_3189 (O_3189,N_29730,N_29806);
nand UO_3190 (O_3190,N_29724,N_29703);
xor UO_3191 (O_3191,N_29722,N_29777);
or UO_3192 (O_3192,N_29755,N_29851);
or UO_3193 (O_3193,N_29809,N_29941);
and UO_3194 (O_3194,N_29825,N_29928);
xnor UO_3195 (O_3195,N_29915,N_29830);
nor UO_3196 (O_3196,N_29945,N_29833);
xnor UO_3197 (O_3197,N_29958,N_29870);
xnor UO_3198 (O_3198,N_29940,N_29753);
or UO_3199 (O_3199,N_29791,N_29852);
xnor UO_3200 (O_3200,N_29701,N_29706);
nor UO_3201 (O_3201,N_29969,N_29875);
and UO_3202 (O_3202,N_29962,N_29973);
nand UO_3203 (O_3203,N_29887,N_29951);
xnor UO_3204 (O_3204,N_29971,N_29851);
xor UO_3205 (O_3205,N_29907,N_29786);
xnor UO_3206 (O_3206,N_29895,N_29709);
nor UO_3207 (O_3207,N_29914,N_29873);
or UO_3208 (O_3208,N_29979,N_29909);
and UO_3209 (O_3209,N_29965,N_29865);
nor UO_3210 (O_3210,N_29898,N_29786);
and UO_3211 (O_3211,N_29726,N_29922);
or UO_3212 (O_3212,N_29810,N_29956);
or UO_3213 (O_3213,N_29861,N_29985);
nand UO_3214 (O_3214,N_29803,N_29936);
nand UO_3215 (O_3215,N_29959,N_29937);
or UO_3216 (O_3216,N_29986,N_29702);
xnor UO_3217 (O_3217,N_29763,N_29869);
and UO_3218 (O_3218,N_29940,N_29991);
nand UO_3219 (O_3219,N_29845,N_29974);
nor UO_3220 (O_3220,N_29880,N_29753);
and UO_3221 (O_3221,N_29890,N_29937);
and UO_3222 (O_3222,N_29918,N_29974);
nor UO_3223 (O_3223,N_29870,N_29988);
or UO_3224 (O_3224,N_29942,N_29717);
nand UO_3225 (O_3225,N_29964,N_29872);
and UO_3226 (O_3226,N_29914,N_29820);
nor UO_3227 (O_3227,N_29924,N_29769);
nor UO_3228 (O_3228,N_29773,N_29913);
and UO_3229 (O_3229,N_29734,N_29994);
or UO_3230 (O_3230,N_29885,N_29863);
xor UO_3231 (O_3231,N_29953,N_29811);
nand UO_3232 (O_3232,N_29815,N_29879);
nor UO_3233 (O_3233,N_29928,N_29947);
and UO_3234 (O_3234,N_29849,N_29741);
or UO_3235 (O_3235,N_29905,N_29932);
nand UO_3236 (O_3236,N_29811,N_29924);
xor UO_3237 (O_3237,N_29800,N_29729);
and UO_3238 (O_3238,N_29904,N_29791);
nor UO_3239 (O_3239,N_29818,N_29810);
nand UO_3240 (O_3240,N_29821,N_29991);
and UO_3241 (O_3241,N_29875,N_29943);
and UO_3242 (O_3242,N_29971,N_29820);
nand UO_3243 (O_3243,N_29781,N_29707);
nand UO_3244 (O_3244,N_29960,N_29899);
nor UO_3245 (O_3245,N_29833,N_29906);
nand UO_3246 (O_3246,N_29962,N_29926);
and UO_3247 (O_3247,N_29813,N_29817);
nor UO_3248 (O_3248,N_29841,N_29930);
and UO_3249 (O_3249,N_29733,N_29792);
nand UO_3250 (O_3250,N_29834,N_29749);
xor UO_3251 (O_3251,N_29809,N_29970);
or UO_3252 (O_3252,N_29701,N_29883);
nand UO_3253 (O_3253,N_29906,N_29990);
or UO_3254 (O_3254,N_29820,N_29958);
nand UO_3255 (O_3255,N_29997,N_29857);
or UO_3256 (O_3256,N_29820,N_29889);
xor UO_3257 (O_3257,N_29972,N_29780);
or UO_3258 (O_3258,N_29999,N_29785);
xor UO_3259 (O_3259,N_29733,N_29779);
or UO_3260 (O_3260,N_29899,N_29759);
and UO_3261 (O_3261,N_29920,N_29947);
and UO_3262 (O_3262,N_29769,N_29751);
xor UO_3263 (O_3263,N_29864,N_29735);
nand UO_3264 (O_3264,N_29760,N_29791);
nand UO_3265 (O_3265,N_29780,N_29986);
xor UO_3266 (O_3266,N_29763,N_29804);
nor UO_3267 (O_3267,N_29982,N_29832);
and UO_3268 (O_3268,N_29799,N_29825);
or UO_3269 (O_3269,N_29751,N_29822);
xor UO_3270 (O_3270,N_29960,N_29822);
nor UO_3271 (O_3271,N_29911,N_29888);
and UO_3272 (O_3272,N_29816,N_29788);
xor UO_3273 (O_3273,N_29967,N_29734);
or UO_3274 (O_3274,N_29981,N_29927);
nand UO_3275 (O_3275,N_29989,N_29991);
and UO_3276 (O_3276,N_29796,N_29984);
nor UO_3277 (O_3277,N_29965,N_29850);
xor UO_3278 (O_3278,N_29810,N_29703);
nor UO_3279 (O_3279,N_29707,N_29808);
and UO_3280 (O_3280,N_29851,N_29908);
and UO_3281 (O_3281,N_29991,N_29810);
xnor UO_3282 (O_3282,N_29984,N_29945);
xnor UO_3283 (O_3283,N_29864,N_29914);
xnor UO_3284 (O_3284,N_29949,N_29766);
xnor UO_3285 (O_3285,N_29951,N_29850);
xor UO_3286 (O_3286,N_29902,N_29849);
nand UO_3287 (O_3287,N_29875,N_29744);
nor UO_3288 (O_3288,N_29944,N_29917);
nand UO_3289 (O_3289,N_29801,N_29739);
nand UO_3290 (O_3290,N_29734,N_29728);
nand UO_3291 (O_3291,N_29875,N_29803);
nand UO_3292 (O_3292,N_29713,N_29800);
xor UO_3293 (O_3293,N_29794,N_29850);
xnor UO_3294 (O_3294,N_29712,N_29723);
nand UO_3295 (O_3295,N_29898,N_29889);
xnor UO_3296 (O_3296,N_29855,N_29904);
xnor UO_3297 (O_3297,N_29927,N_29740);
nor UO_3298 (O_3298,N_29965,N_29857);
and UO_3299 (O_3299,N_29734,N_29815);
nand UO_3300 (O_3300,N_29891,N_29983);
nand UO_3301 (O_3301,N_29739,N_29986);
and UO_3302 (O_3302,N_29829,N_29898);
nor UO_3303 (O_3303,N_29707,N_29716);
nor UO_3304 (O_3304,N_29901,N_29843);
nor UO_3305 (O_3305,N_29894,N_29927);
xnor UO_3306 (O_3306,N_29984,N_29715);
xnor UO_3307 (O_3307,N_29757,N_29753);
or UO_3308 (O_3308,N_29865,N_29974);
nor UO_3309 (O_3309,N_29889,N_29830);
nand UO_3310 (O_3310,N_29747,N_29897);
nor UO_3311 (O_3311,N_29700,N_29902);
xor UO_3312 (O_3312,N_29789,N_29842);
and UO_3313 (O_3313,N_29888,N_29972);
or UO_3314 (O_3314,N_29860,N_29950);
or UO_3315 (O_3315,N_29907,N_29882);
or UO_3316 (O_3316,N_29995,N_29986);
nand UO_3317 (O_3317,N_29998,N_29867);
or UO_3318 (O_3318,N_29985,N_29932);
nand UO_3319 (O_3319,N_29976,N_29929);
nor UO_3320 (O_3320,N_29746,N_29874);
nor UO_3321 (O_3321,N_29987,N_29979);
or UO_3322 (O_3322,N_29884,N_29899);
xnor UO_3323 (O_3323,N_29741,N_29910);
nor UO_3324 (O_3324,N_29961,N_29984);
or UO_3325 (O_3325,N_29948,N_29786);
nor UO_3326 (O_3326,N_29981,N_29870);
nand UO_3327 (O_3327,N_29781,N_29872);
and UO_3328 (O_3328,N_29968,N_29771);
or UO_3329 (O_3329,N_29940,N_29915);
nand UO_3330 (O_3330,N_29987,N_29894);
xor UO_3331 (O_3331,N_29806,N_29814);
nand UO_3332 (O_3332,N_29810,N_29843);
and UO_3333 (O_3333,N_29724,N_29960);
and UO_3334 (O_3334,N_29788,N_29822);
nand UO_3335 (O_3335,N_29810,N_29827);
nor UO_3336 (O_3336,N_29798,N_29983);
nor UO_3337 (O_3337,N_29991,N_29987);
xor UO_3338 (O_3338,N_29802,N_29913);
nor UO_3339 (O_3339,N_29756,N_29778);
or UO_3340 (O_3340,N_29709,N_29721);
or UO_3341 (O_3341,N_29806,N_29940);
nand UO_3342 (O_3342,N_29770,N_29944);
xnor UO_3343 (O_3343,N_29759,N_29735);
or UO_3344 (O_3344,N_29918,N_29917);
xnor UO_3345 (O_3345,N_29966,N_29720);
and UO_3346 (O_3346,N_29793,N_29810);
nand UO_3347 (O_3347,N_29777,N_29902);
nand UO_3348 (O_3348,N_29733,N_29968);
xnor UO_3349 (O_3349,N_29856,N_29988);
or UO_3350 (O_3350,N_29846,N_29736);
xor UO_3351 (O_3351,N_29709,N_29850);
nor UO_3352 (O_3352,N_29803,N_29979);
and UO_3353 (O_3353,N_29788,N_29800);
or UO_3354 (O_3354,N_29961,N_29860);
nor UO_3355 (O_3355,N_29736,N_29801);
nor UO_3356 (O_3356,N_29931,N_29825);
and UO_3357 (O_3357,N_29932,N_29973);
or UO_3358 (O_3358,N_29776,N_29854);
nor UO_3359 (O_3359,N_29996,N_29701);
xnor UO_3360 (O_3360,N_29843,N_29912);
nor UO_3361 (O_3361,N_29920,N_29925);
and UO_3362 (O_3362,N_29927,N_29926);
nor UO_3363 (O_3363,N_29919,N_29820);
nor UO_3364 (O_3364,N_29935,N_29970);
or UO_3365 (O_3365,N_29813,N_29724);
or UO_3366 (O_3366,N_29910,N_29820);
nand UO_3367 (O_3367,N_29774,N_29930);
and UO_3368 (O_3368,N_29999,N_29761);
nand UO_3369 (O_3369,N_29993,N_29910);
nand UO_3370 (O_3370,N_29936,N_29970);
nand UO_3371 (O_3371,N_29706,N_29731);
or UO_3372 (O_3372,N_29804,N_29835);
nand UO_3373 (O_3373,N_29720,N_29860);
nand UO_3374 (O_3374,N_29706,N_29834);
xnor UO_3375 (O_3375,N_29799,N_29818);
or UO_3376 (O_3376,N_29927,N_29918);
nor UO_3377 (O_3377,N_29703,N_29793);
xor UO_3378 (O_3378,N_29705,N_29822);
and UO_3379 (O_3379,N_29938,N_29915);
or UO_3380 (O_3380,N_29837,N_29938);
xor UO_3381 (O_3381,N_29776,N_29804);
nor UO_3382 (O_3382,N_29941,N_29868);
or UO_3383 (O_3383,N_29885,N_29754);
xnor UO_3384 (O_3384,N_29926,N_29914);
and UO_3385 (O_3385,N_29805,N_29883);
nor UO_3386 (O_3386,N_29844,N_29880);
nor UO_3387 (O_3387,N_29924,N_29750);
and UO_3388 (O_3388,N_29927,N_29841);
nor UO_3389 (O_3389,N_29930,N_29747);
or UO_3390 (O_3390,N_29885,N_29871);
and UO_3391 (O_3391,N_29969,N_29802);
nor UO_3392 (O_3392,N_29940,N_29767);
or UO_3393 (O_3393,N_29989,N_29945);
xor UO_3394 (O_3394,N_29936,N_29840);
nor UO_3395 (O_3395,N_29789,N_29868);
or UO_3396 (O_3396,N_29864,N_29790);
nor UO_3397 (O_3397,N_29883,N_29935);
and UO_3398 (O_3398,N_29758,N_29749);
nand UO_3399 (O_3399,N_29784,N_29714);
nand UO_3400 (O_3400,N_29739,N_29775);
nor UO_3401 (O_3401,N_29960,N_29946);
xnor UO_3402 (O_3402,N_29892,N_29882);
or UO_3403 (O_3403,N_29909,N_29786);
nor UO_3404 (O_3404,N_29749,N_29902);
or UO_3405 (O_3405,N_29743,N_29823);
xnor UO_3406 (O_3406,N_29924,N_29791);
xor UO_3407 (O_3407,N_29729,N_29851);
and UO_3408 (O_3408,N_29891,N_29834);
xor UO_3409 (O_3409,N_29865,N_29756);
nand UO_3410 (O_3410,N_29718,N_29797);
nor UO_3411 (O_3411,N_29771,N_29979);
nand UO_3412 (O_3412,N_29959,N_29857);
xnor UO_3413 (O_3413,N_29854,N_29962);
nand UO_3414 (O_3414,N_29977,N_29726);
and UO_3415 (O_3415,N_29714,N_29981);
nand UO_3416 (O_3416,N_29708,N_29920);
nand UO_3417 (O_3417,N_29812,N_29789);
nand UO_3418 (O_3418,N_29863,N_29890);
xor UO_3419 (O_3419,N_29855,N_29723);
xnor UO_3420 (O_3420,N_29718,N_29938);
nor UO_3421 (O_3421,N_29982,N_29844);
xor UO_3422 (O_3422,N_29787,N_29917);
or UO_3423 (O_3423,N_29741,N_29918);
nor UO_3424 (O_3424,N_29749,N_29787);
xor UO_3425 (O_3425,N_29951,N_29818);
and UO_3426 (O_3426,N_29801,N_29815);
xnor UO_3427 (O_3427,N_29750,N_29874);
xor UO_3428 (O_3428,N_29707,N_29955);
nor UO_3429 (O_3429,N_29839,N_29757);
nor UO_3430 (O_3430,N_29913,N_29727);
and UO_3431 (O_3431,N_29809,N_29974);
nor UO_3432 (O_3432,N_29848,N_29898);
xnor UO_3433 (O_3433,N_29957,N_29797);
nor UO_3434 (O_3434,N_29966,N_29753);
nor UO_3435 (O_3435,N_29813,N_29856);
or UO_3436 (O_3436,N_29938,N_29827);
and UO_3437 (O_3437,N_29991,N_29870);
xnor UO_3438 (O_3438,N_29839,N_29715);
nor UO_3439 (O_3439,N_29834,N_29929);
xnor UO_3440 (O_3440,N_29931,N_29734);
xor UO_3441 (O_3441,N_29807,N_29853);
and UO_3442 (O_3442,N_29917,N_29746);
and UO_3443 (O_3443,N_29727,N_29722);
xor UO_3444 (O_3444,N_29728,N_29872);
and UO_3445 (O_3445,N_29805,N_29851);
or UO_3446 (O_3446,N_29870,N_29844);
nor UO_3447 (O_3447,N_29976,N_29732);
xnor UO_3448 (O_3448,N_29865,N_29703);
nand UO_3449 (O_3449,N_29856,N_29993);
xor UO_3450 (O_3450,N_29897,N_29862);
or UO_3451 (O_3451,N_29799,N_29944);
nand UO_3452 (O_3452,N_29871,N_29738);
nor UO_3453 (O_3453,N_29893,N_29774);
nor UO_3454 (O_3454,N_29911,N_29833);
nor UO_3455 (O_3455,N_29979,N_29776);
xnor UO_3456 (O_3456,N_29710,N_29939);
or UO_3457 (O_3457,N_29802,N_29797);
and UO_3458 (O_3458,N_29717,N_29754);
xor UO_3459 (O_3459,N_29951,N_29839);
xor UO_3460 (O_3460,N_29853,N_29816);
xnor UO_3461 (O_3461,N_29878,N_29827);
or UO_3462 (O_3462,N_29844,N_29772);
nor UO_3463 (O_3463,N_29896,N_29758);
nand UO_3464 (O_3464,N_29943,N_29869);
nand UO_3465 (O_3465,N_29949,N_29721);
xor UO_3466 (O_3466,N_29714,N_29946);
nor UO_3467 (O_3467,N_29952,N_29820);
nand UO_3468 (O_3468,N_29714,N_29758);
nand UO_3469 (O_3469,N_29904,N_29709);
nor UO_3470 (O_3470,N_29932,N_29979);
or UO_3471 (O_3471,N_29800,N_29728);
xor UO_3472 (O_3472,N_29896,N_29775);
nand UO_3473 (O_3473,N_29911,N_29775);
or UO_3474 (O_3474,N_29999,N_29910);
nor UO_3475 (O_3475,N_29743,N_29777);
and UO_3476 (O_3476,N_29855,N_29988);
nor UO_3477 (O_3477,N_29975,N_29902);
xnor UO_3478 (O_3478,N_29977,N_29725);
and UO_3479 (O_3479,N_29705,N_29728);
or UO_3480 (O_3480,N_29985,N_29884);
and UO_3481 (O_3481,N_29835,N_29927);
and UO_3482 (O_3482,N_29703,N_29732);
nand UO_3483 (O_3483,N_29941,N_29840);
nand UO_3484 (O_3484,N_29738,N_29918);
and UO_3485 (O_3485,N_29882,N_29981);
nor UO_3486 (O_3486,N_29702,N_29929);
xor UO_3487 (O_3487,N_29791,N_29936);
or UO_3488 (O_3488,N_29924,N_29894);
and UO_3489 (O_3489,N_29815,N_29931);
nor UO_3490 (O_3490,N_29793,N_29867);
xor UO_3491 (O_3491,N_29795,N_29980);
nor UO_3492 (O_3492,N_29997,N_29710);
nand UO_3493 (O_3493,N_29786,N_29918);
xnor UO_3494 (O_3494,N_29769,N_29732);
or UO_3495 (O_3495,N_29915,N_29731);
and UO_3496 (O_3496,N_29865,N_29799);
and UO_3497 (O_3497,N_29727,N_29972);
or UO_3498 (O_3498,N_29747,N_29955);
xor UO_3499 (O_3499,N_29763,N_29754);
endmodule