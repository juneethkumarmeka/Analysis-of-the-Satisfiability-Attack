module basic_500_3000_500_6_levels_1xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_409,In_69);
xor U1 (N_1,In_263,In_481);
and U2 (N_2,In_279,In_261);
nand U3 (N_3,In_337,In_239);
and U4 (N_4,In_389,In_424);
and U5 (N_5,In_15,In_336);
and U6 (N_6,In_485,In_117);
nor U7 (N_7,In_451,In_235);
or U8 (N_8,In_57,In_269);
nor U9 (N_9,In_222,In_56);
or U10 (N_10,In_1,In_355);
or U11 (N_11,In_305,In_496);
or U12 (N_12,In_349,In_465);
nand U13 (N_13,In_47,In_456);
nand U14 (N_14,In_65,In_4);
and U15 (N_15,In_135,In_414);
nand U16 (N_16,In_123,In_229);
or U17 (N_17,In_7,In_205);
or U18 (N_18,In_29,In_433);
and U19 (N_19,In_395,In_266);
nor U20 (N_20,In_233,In_126);
or U21 (N_21,In_248,In_498);
or U22 (N_22,In_330,In_323);
and U23 (N_23,In_25,In_209);
nor U24 (N_24,In_489,In_163);
and U25 (N_25,In_371,In_367);
and U26 (N_26,In_119,In_92);
or U27 (N_27,In_315,In_84);
nor U28 (N_28,In_335,In_272);
or U29 (N_29,In_404,In_434);
and U30 (N_30,In_36,In_6);
or U31 (N_31,In_76,In_319);
or U32 (N_32,In_444,In_197);
and U33 (N_33,In_386,In_368);
or U34 (N_34,In_215,In_180);
or U35 (N_35,In_447,In_394);
or U36 (N_36,In_254,In_11);
nor U37 (N_37,In_361,In_155);
nor U38 (N_38,In_369,In_353);
nor U39 (N_39,In_463,In_24);
and U40 (N_40,In_396,In_78);
nor U41 (N_41,In_12,In_283);
nand U42 (N_42,In_291,In_352);
or U43 (N_43,In_246,In_177);
nor U44 (N_44,In_2,In_364);
or U45 (N_45,In_50,In_164);
and U46 (N_46,In_322,In_129);
nor U47 (N_47,In_74,In_412);
nand U48 (N_48,In_111,In_179);
and U49 (N_49,In_347,In_309);
nand U50 (N_50,In_181,In_213);
and U51 (N_51,In_268,In_243);
or U52 (N_52,In_391,In_267);
nand U53 (N_53,In_462,In_423);
nand U54 (N_54,In_170,In_143);
nor U55 (N_55,In_372,In_341);
nand U56 (N_56,In_468,In_41);
or U57 (N_57,In_431,In_362);
and U58 (N_58,In_326,In_61);
or U59 (N_59,In_294,In_342);
xnor U60 (N_60,In_86,In_473);
and U61 (N_61,In_317,In_397);
or U62 (N_62,In_174,In_38);
nand U63 (N_63,In_26,In_259);
and U64 (N_64,In_437,In_488);
and U65 (N_65,In_441,In_120);
nand U66 (N_66,In_313,In_172);
and U67 (N_67,In_30,In_82);
nor U68 (N_68,In_125,In_350);
nand U69 (N_69,In_381,In_124);
nor U70 (N_70,In_234,In_471);
or U71 (N_71,In_399,In_188);
and U72 (N_72,In_478,In_348);
or U73 (N_73,In_48,In_118);
nand U74 (N_74,In_405,In_208);
nand U75 (N_75,In_320,In_192);
or U76 (N_76,In_311,In_55);
nand U77 (N_77,In_327,In_277);
or U78 (N_78,In_303,In_392);
nand U79 (N_79,In_220,In_278);
or U80 (N_80,In_210,In_23);
nor U81 (N_81,In_101,In_310);
or U82 (N_82,In_132,In_285);
nand U83 (N_83,In_257,In_71);
or U84 (N_84,In_255,In_206);
and U85 (N_85,In_344,In_5);
and U86 (N_86,In_284,In_228);
xor U87 (N_87,In_9,In_318);
or U88 (N_88,In_122,In_448);
or U89 (N_89,In_75,In_469);
nand U90 (N_90,In_19,In_144);
nand U91 (N_91,In_443,In_385);
or U92 (N_92,In_44,In_432);
or U93 (N_93,In_33,In_360);
or U94 (N_94,In_383,In_288);
or U95 (N_95,In_316,In_499);
nor U96 (N_96,In_491,In_88);
nor U97 (N_97,In_312,In_321);
or U98 (N_98,In_147,In_438);
nand U99 (N_99,In_31,In_487);
and U100 (N_100,In_64,In_128);
or U101 (N_101,In_449,In_230);
nor U102 (N_102,In_380,In_271);
nor U103 (N_103,In_133,In_152);
and U104 (N_104,In_116,In_426);
nand U105 (N_105,In_354,In_211);
nand U106 (N_106,In_238,In_241);
or U107 (N_107,In_453,In_388);
or U108 (N_108,In_258,In_202);
and U109 (N_109,In_393,In_265);
nand U110 (N_110,In_160,In_379);
or U111 (N_111,In_137,In_52);
nor U112 (N_112,In_338,In_474);
and U113 (N_113,In_419,In_136);
or U114 (N_114,In_8,In_45);
and U115 (N_115,In_13,In_356);
and U116 (N_116,In_245,In_95);
and U117 (N_117,In_231,In_176);
or U118 (N_118,In_182,In_89);
or U119 (N_119,In_332,In_292);
nand U120 (N_120,In_403,In_457);
nor U121 (N_121,In_363,In_195);
nand U122 (N_122,In_400,In_186);
nand U123 (N_123,In_264,In_401);
nor U124 (N_124,In_333,In_35);
and U125 (N_125,In_459,In_314);
or U126 (N_126,In_227,In_113);
nor U127 (N_127,In_430,In_154);
and U128 (N_128,In_280,In_276);
nor U129 (N_129,In_219,In_439);
nand U130 (N_130,In_328,In_304);
and U131 (N_131,In_273,In_112);
and U132 (N_132,In_458,In_308);
nor U133 (N_133,In_121,In_18);
and U134 (N_134,In_413,In_454);
nor U135 (N_135,In_387,In_274);
and U136 (N_136,In_198,In_40);
nand U137 (N_137,In_27,In_460);
nand U138 (N_138,In_226,In_58);
nor U139 (N_139,In_183,In_452);
nand U140 (N_140,In_260,In_106);
or U141 (N_141,In_196,In_166);
and U142 (N_142,In_168,In_79);
nor U143 (N_143,In_169,In_300);
and U144 (N_144,In_237,In_3);
or U145 (N_145,In_203,In_67);
and U146 (N_146,In_60,In_435);
nor U147 (N_147,In_420,In_306);
nor U148 (N_148,In_217,In_297);
nand U149 (N_149,In_96,In_127);
or U150 (N_150,In_140,In_91);
nor U151 (N_151,In_429,In_83);
nor U152 (N_152,In_49,In_214);
or U153 (N_153,In_94,In_224);
nor U154 (N_154,In_290,In_493);
nand U155 (N_155,In_99,In_199);
or U156 (N_156,In_244,In_109);
and U157 (N_157,In_175,In_43);
or U158 (N_158,In_376,In_110);
or U159 (N_159,In_296,In_194);
and U160 (N_160,In_77,In_105);
and U161 (N_161,In_289,In_373);
nand U162 (N_162,In_165,In_374);
and U163 (N_163,In_398,In_455);
and U164 (N_164,In_256,In_242);
nor U165 (N_165,In_150,In_85);
and U166 (N_166,In_384,In_0);
or U167 (N_167,In_422,In_73);
or U168 (N_168,In_80,In_286);
nand U169 (N_169,In_200,In_21);
nand U170 (N_170,In_87,In_149);
and U171 (N_171,In_20,In_446);
or U172 (N_172,In_477,In_358);
nand U173 (N_173,In_416,In_161);
or U174 (N_174,In_62,In_93);
and U175 (N_175,In_467,In_298);
nor U176 (N_176,In_247,In_299);
and U177 (N_177,In_301,In_334);
nand U178 (N_178,In_325,In_32);
nand U179 (N_179,In_159,In_167);
or U180 (N_180,In_494,In_351);
and U181 (N_181,In_148,In_39);
nand U182 (N_182,In_107,In_331);
nor U183 (N_183,In_377,In_72);
and U184 (N_184,In_100,In_406);
nand U185 (N_185,In_53,In_486);
and U186 (N_186,In_470,In_492);
or U187 (N_187,In_440,In_483);
nor U188 (N_188,In_216,In_157);
or U189 (N_189,In_131,In_10);
and U190 (N_190,In_282,In_402);
nor U191 (N_191,In_14,In_357);
or U192 (N_192,In_340,In_218);
and U193 (N_193,In_153,In_90);
or U194 (N_194,In_54,In_421);
or U195 (N_195,In_145,In_345);
nand U196 (N_196,In_189,In_302);
and U197 (N_197,In_343,In_251);
nand U198 (N_198,In_466,In_130);
and U199 (N_199,In_418,In_28);
or U200 (N_200,In_225,In_221);
nor U201 (N_201,In_68,In_171);
nand U202 (N_202,In_97,In_425);
nor U203 (N_203,In_472,In_461);
or U204 (N_204,In_275,In_464);
and U205 (N_205,In_223,In_442);
nor U206 (N_206,In_490,In_115);
nor U207 (N_207,In_295,In_34);
or U208 (N_208,In_370,In_249);
nand U209 (N_209,In_495,In_236);
or U210 (N_210,In_427,In_187);
nor U211 (N_211,In_193,In_270);
nor U212 (N_212,In_339,In_212);
nor U213 (N_213,In_151,In_103);
and U214 (N_214,In_410,In_436);
or U215 (N_215,In_42,In_365);
nand U216 (N_216,In_146,In_232);
or U217 (N_217,In_476,In_46);
and U218 (N_218,In_59,In_480);
nor U219 (N_219,In_324,In_204);
or U220 (N_220,In_415,In_191);
nor U221 (N_221,In_417,In_482);
nor U222 (N_222,In_190,In_329);
and U223 (N_223,In_382,In_70);
nor U224 (N_224,In_185,In_479);
nand U225 (N_225,In_158,In_63);
nor U226 (N_226,In_287,In_37);
or U227 (N_227,In_240,In_102);
nor U228 (N_228,In_281,In_262);
or U229 (N_229,In_114,In_184);
nor U230 (N_230,In_66,In_250);
or U231 (N_231,In_141,In_178);
nand U232 (N_232,In_378,In_207);
nand U233 (N_233,In_445,In_138);
nor U234 (N_234,In_134,In_98);
nand U235 (N_235,In_293,In_484);
and U236 (N_236,In_162,In_252);
or U237 (N_237,In_497,In_142);
or U238 (N_238,In_253,In_201);
and U239 (N_239,In_51,In_104);
or U240 (N_240,In_359,In_411);
or U241 (N_241,In_408,In_16);
and U242 (N_242,In_139,In_390);
or U243 (N_243,In_346,In_375);
or U244 (N_244,In_17,In_173);
or U245 (N_245,In_366,In_407);
nor U246 (N_246,In_475,In_428);
and U247 (N_247,In_156,In_22);
and U248 (N_248,In_450,In_108);
nand U249 (N_249,In_81,In_307);
xnor U250 (N_250,In_124,In_198);
or U251 (N_251,In_367,In_92);
nand U252 (N_252,In_343,In_374);
and U253 (N_253,In_456,In_25);
nor U254 (N_254,In_499,In_305);
nor U255 (N_255,In_329,In_191);
nand U256 (N_256,In_338,In_277);
nor U257 (N_257,In_220,In_9);
nor U258 (N_258,In_247,In_467);
nor U259 (N_259,In_294,In_457);
nand U260 (N_260,In_228,In_103);
and U261 (N_261,In_187,In_297);
nand U262 (N_262,In_250,In_385);
or U263 (N_263,In_447,In_86);
nor U264 (N_264,In_61,In_70);
nand U265 (N_265,In_331,In_452);
and U266 (N_266,In_434,In_340);
nor U267 (N_267,In_127,In_17);
and U268 (N_268,In_292,In_126);
or U269 (N_269,In_468,In_112);
and U270 (N_270,In_2,In_112);
nand U271 (N_271,In_283,In_27);
and U272 (N_272,In_145,In_394);
nor U273 (N_273,In_336,In_61);
nor U274 (N_274,In_321,In_126);
nor U275 (N_275,In_299,In_377);
or U276 (N_276,In_116,In_384);
nand U277 (N_277,In_146,In_282);
nand U278 (N_278,In_499,In_227);
and U279 (N_279,In_161,In_28);
nand U280 (N_280,In_359,In_185);
nor U281 (N_281,In_108,In_306);
or U282 (N_282,In_229,In_271);
and U283 (N_283,In_127,In_158);
or U284 (N_284,In_315,In_338);
and U285 (N_285,In_223,In_371);
nor U286 (N_286,In_52,In_257);
and U287 (N_287,In_411,In_495);
nand U288 (N_288,In_401,In_90);
nor U289 (N_289,In_10,In_463);
nand U290 (N_290,In_356,In_404);
and U291 (N_291,In_132,In_106);
or U292 (N_292,In_440,In_153);
nor U293 (N_293,In_353,In_107);
and U294 (N_294,In_268,In_57);
nand U295 (N_295,In_179,In_391);
nor U296 (N_296,In_315,In_211);
or U297 (N_297,In_437,In_98);
nor U298 (N_298,In_72,In_224);
nor U299 (N_299,In_479,In_233);
nand U300 (N_300,In_294,In_285);
and U301 (N_301,In_221,In_260);
nor U302 (N_302,In_286,In_65);
nor U303 (N_303,In_204,In_23);
nand U304 (N_304,In_485,In_314);
nand U305 (N_305,In_403,In_48);
nand U306 (N_306,In_17,In_211);
and U307 (N_307,In_207,In_52);
xnor U308 (N_308,In_447,In_330);
nand U309 (N_309,In_407,In_180);
or U310 (N_310,In_313,In_275);
and U311 (N_311,In_313,In_393);
nand U312 (N_312,In_20,In_255);
or U313 (N_313,In_230,In_199);
nor U314 (N_314,In_255,In_391);
nor U315 (N_315,In_181,In_176);
nand U316 (N_316,In_477,In_264);
and U317 (N_317,In_463,In_401);
and U318 (N_318,In_269,In_495);
or U319 (N_319,In_206,In_80);
and U320 (N_320,In_384,In_433);
or U321 (N_321,In_484,In_307);
nand U322 (N_322,In_480,In_184);
nor U323 (N_323,In_234,In_35);
or U324 (N_324,In_103,In_342);
nand U325 (N_325,In_92,In_185);
xor U326 (N_326,In_205,In_262);
nand U327 (N_327,In_484,In_103);
nor U328 (N_328,In_193,In_179);
nor U329 (N_329,In_432,In_23);
nand U330 (N_330,In_328,In_106);
or U331 (N_331,In_264,In_4);
and U332 (N_332,In_303,In_363);
or U333 (N_333,In_393,In_140);
nand U334 (N_334,In_428,In_297);
or U335 (N_335,In_402,In_129);
nand U336 (N_336,In_381,In_196);
or U337 (N_337,In_319,In_323);
or U338 (N_338,In_279,In_401);
or U339 (N_339,In_161,In_199);
or U340 (N_340,In_216,In_27);
nor U341 (N_341,In_57,In_19);
or U342 (N_342,In_266,In_48);
and U343 (N_343,In_377,In_194);
and U344 (N_344,In_398,In_437);
nor U345 (N_345,In_251,In_344);
and U346 (N_346,In_247,In_85);
nand U347 (N_347,In_482,In_305);
nor U348 (N_348,In_448,In_312);
nor U349 (N_349,In_313,In_76);
nor U350 (N_350,In_460,In_15);
and U351 (N_351,In_478,In_340);
nor U352 (N_352,In_440,In_148);
and U353 (N_353,In_134,In_188);
or U354 (N_354,In_369,In_348);
nor U355 (N_355,In_353,In_429);
or U356 (N_356,In_92,In_198);
nand U357 (N_357,In_437,In_304);
nand U358 (N_358,In_86,In_293);
nor U359 (N_359,In_371,In_366);
nand U360 (N_360,In_447,In_238);
or U361 (N_361,In_209,In_358);
or U362 (N_362,In_1,In_476);
nand U363 (N_363,In_293,In_470);
and U364 (N_364,In_268,In_185);
or U365 (N_365,In_96,In_298);
nand U366 (N_366,In_285,In_168);
nand U367 (N_367,In_443,In_361);
nor U368 (N_368,In_417,In_356);
nor U369 (N_369,In_249,In_151);
nor U370 (N_370,In_481,In_208);
nand U371 (N_371,In_210,In_313);
and U372 (N_372,In_351,In_139);
nand U373 (N_373,In_472,In_283);
nor U374 (N_374,In_206,In_230);
nor U375 (N_375,In_224,In_489);
and U376 (N_376,In_58,In_439);
or U377 (N_377,In_279,In_27);
and U378 (N_378,In_299,In_439);
or U379 (N_379,In_252,In_463);
nand U380 (N_380,In_306,In_381);
nand U381 (N_381,In_339,In_14);
nor U382 (N_382,In_430,In_389);
nand U383 (N_383,In_490,In_415);
nor U384 (N_384,In_397,In_285);
and U385 (N_385,In_279,In_204);
or U386 (N_386,In_146,In_105);
nor U387 (N_387,In_179,In_357);
xnor U388 (N_388,In_122,In_112);
nor U389 (N_389,In_73,In_484);
and U390 (N_390,In_282,In_141);
and U391 (N_391,In_51,In_496);
and U392 (N_392,In_193,In_392);
nand U393 (N_393,In_312,In_74);
nand U394 (N_394,In_479,In_1);
nand U395 (N_395,In_401,In_229);
nand U396 (N_396,In_44,In_91);
nor U397 (N_397,In_26,In_12);
nand U398 (N_398,In_75,In_113);
and U399 (N_399,In_194,In_40);
and U400 (N_400,In_458,In_211);
nand U401 (N_401,In_371,In_340);
nand U402 (N_402,In_148,In_373);
nor U403 (N_403,In_123,In_228);
nor U404 (N_404,In_394,In_32);
nor U405 (N_405,In_111,In_152);
and U406 (N_406,In_74,In_47);
nor U407 (N_407,In_200,In_124);
or U408 (N_408,In_455,In_380);
nand U409 (N_409,In_152,In_387);
nand U410 (N_410,In_311,In_492);
and U411 (N_411,In_304,In_255);
or U412 (N_412,In_183,In_361);
and U413 (N_413,In_353,In_304);
or U414 (N_414,In_476,In_180);
or U415 (N_415,In_492,In_478);
nor U416 (N_416,In_428,In_87);
nand U417 (N_417,In_290,In_367);
nor U418 (N_418,In_130,In_304);
nand U419 (N_419,In_39,In_274);
or U420 (N_420,In_17,In_281);
or U421 (N_421,In_110,In_481);
xor U422 (N_422,In_302,In_312);
nor U423 (N_423,In_105,In_469);
and U424 (N_424,In_147,In_218);
nor U425 (N_425,In_167,In_497);
nor U426 (N_426,In_459,In_60);
nand U427 (N_427,In_238,In_338);
nand U428 (N_428,In_40,In_313);
or U429 (N_429,In_396,In_400);
nor U430 (N_430,In_128,In_495);
or U431 (N_431,In_276,In_301);
and U432 (N_432,In_29,In_482);
nand U433 (N_433,In_466,In_417);
and U434 (N_434,In_208,In_494);
and U435 (N_435,In_497,In_481);
or U436 (N_436,In_302,In_108);
nand U437 (N_437,In_333,In_166);
and U438 (N_438,In_254,In_365);
or U439 (N_439,In_305,In_150);
nand U440 (N_440,In_303,In_33);
or U441 (N_441,In_99,In_14);
and U442 (N_442,In_317,In_182);
nand U443 (N_443,In_4,In_23);
or U444 (N_444,In_201,In_259);
and U445 (N_445,In_367,In_489);
nand U446 (N_446,In_256,In_282);
nand U447 (N_447,In_305,In_85);
or U448 (N_448,In_75,In_89);
nor U449 (N_449,In_393,In_341);
nand U450 (N_450,In_198,In_59);
nand U451 (N_451,In_45,In_421);
and U452 (N_452,In_110,In_377);
and U453 (N_453,In_170,In_383);
or U454 (N_454,In_51,In_477);
nand U455 (N_455,In_246,In_70);
and U456 (N_456,In_81,In_8);
and U457 (N_457,In_382,In_246);
nor U458 (N_458,In_294,In_97);
and U459 (N_459,In_10,In_336);
or U460 (N_460,In_193,In_291);
nor U461 (N_461,In_125,In_342);
nor U462 (N_462,In_13,In_469);
nor U463 (N_463,In_429,In_484);
nor U464 (N_464,In_439,In_454);
nor U465 (N_465,In_277,In_56);
nor U466 (N_466,In_459,In_139);
and U467 (N_467,In_448,In_206);
and U468 (N_468,In_261,In_348);
nand U469 (N_469,In_439,In_217);
and U470 (N_470,In_370,In_207);
nand U471 (N_471,In_343,In_400);
or U472 (N_472,In_239,In_12);
nand U473 (N_473,In_412,In_233);
nand U474 (N_474,In_80,In_112);
nor U475 (N_475,In_119,In_276);
and U476 (N_476,In_7,In_462);
nand U477 (N_477,In_187,In_235);
or U478 (N_478,In_337,In_427);
and U479 (N_479,In_38,In_51);
nand U480 (N_480,In_37,In_229);
nor U481 (N_481,In_498,In_265);
or U482 (N_482,In_407,In_490);
nand U483 (N_483,In_332,In_438);
nor U484 (N_484,In_284,In_446);
nor U485 (N_485,In_491,In_166);
or U486 (N_486,In_230,In_293);
nor U487 (N_487,In_161,In_224);
nand U488 (N_488,In_151,In_478);
nand U489 (N_489,In_216,In_191);
nand U490 (N_490,In_349,In_47);
or U491 (N_491,In_370,In_492);
or U492 (N_492,In_244,In_384);
and U493 (N_493,In_39,In_212);
and U494 (N_494,In_88,In_304);
or U495 (N_495,In_462,In_97);
nand U496 (N_496,In_476,In_113);
nand U497 (N_497,In_55,In_348);
nor U498 (N_498,In_359,In_402);
and U499 (N_499,In_198,In_217);
and U500 (N_500,N_209,N_118);
nor U501 (N_501,N_103,N_473);
nor U502 (N_502,N_408,N_309);
or U503 (N_503,N_87,N_183);
nand U504 (N_504,N_300,N_353);
nand U505 (N_505,N_66,N_215);
and U506 (N_506,N_438,N_277);
and U507 (N_507,N_211,N_255);
nand U508 (N_508,N_371,N_53);
nor U509 (N_509,N_433,N_282);
or U510 (N_510,N_377,N_30);
and U511 (N_511,N_264,N_281);
nor U512 (N_512,N_100,N_315);
nand U513 (N_513,N_329,N_499);
and U514 (N_514,N_213,N_405);
nor U515 (N_515,N_461,N_401);
or U516 (N_516,N_276,N_271);
nor U517 (N_517,N_81,N_137);
and U518 (N_518,N_252,N_71);
nand U519 (N_519,N_304,N_67);
nand U520 (N_520,N_159,N_373);
nand U521 (N_521,N_131,N_201);
or U522 (N_522,N_170,N_241);
and U523 (N_523,N_199,N_345);
and U524 (N_524,N_322,N_3);
nand U525 (N_525,N_99,N_341);
nand U526 (N_526,N_95,N_4);
and U527 (N_527,N_383,N_111);
and U528 (N_528,N_143,N_495);
xor U529 (N_529,N_75,N_445);
or U530 (N_530,N_244,N_45);
or U531 (N_531,N_279,N_348);
and U532 (N_532,N_226,N_289);
nor U533 (N_533,N_290,N_372);
or U534 (N_534,N_306,N_80);
nand U535 (N_535,N_466,N_181);
and U536 (N_536,N_272,N_479);
nand U537 (N_537,N_367,N_478);
and U538 (N_538,N_34,N_370);
nor U539 (N_539,N_64,N_157);
nand U540 (N_540,N_196,N_337);
nand U541 (N_541,N_173,N_317);
nand U542 (N_542,N_406,N_292);
or U543 (N_543,N_327,N_312);
or U544 (N_544,N_263,N_121);
nand U545 (N_545,N_19,N_480);
nor U546 (N_546,N_485,N_114);
and U547 (N_547,N_26,N_357);
nor U548 (N_548,N_283,N_227);
and U549 (N_549,N_85,N_325);
and U550 (N_550,N_220,N_351);
and U551 (N_551,N_409,N_313);
nor U552 (N_552,N_65,N_236);
nor U553 (N_553,N_490,N_278);
or U554 (N_554,N_413,N_331);
nand U555 (N_555,N_303,N_462);
and U556 (N_556,N_140,N_135);
or U557 (N_557,N_185,N_486);
and U558 (N_558,N_402,N_294);
and U559 (N_559,N_422,N_41);
or U560 (N_560,N_37,N_437);
and U561 (N_561,N_22,N_350);
nor U562 (N_562,N_334,N_54);
nor U563 (N_563,N_129,N_84);
xnor U564 (N_564,N_295,N_18);
or U565 (N_565,N_78,N_247);
nand U566 (N_566,N_117,N_262);
or U567 (N_567,N_430,N_460);
nand U568 (N_568,N_1,N_464);
nor U569 (N_569,N_275,N_219);
nand U570 (N_570,N_128,N_191);
and U571 (N_571,N_69,N_122);
nor U572 (N_572,N_17,N_239);
nand U573 (N_573,N_61,N_43);
nor U574 (N_574,N_369,N_342);
nand U575 (N_575,N_432,N_182);
or U576 (N_576,N_447,N_204);
nor U577 (N_577,N_228,N_355);
and U578 (N_578,N_8,N_206);
or U579 (N_579,N_200,N_119);
nand U580 (N_580,N_392,N_302);
xnor U581 (N_581,N_179,N_444);
and U582 (N_582,N_463,N_29);
or U583 (N_583,N_127,N_494);
nand U584 (N_584,N_165,N_364);
and U585 (N_585,N_393,N_47);
or U586 (N_586,N_15,N_189);
nand U587 (N_587,N_139,N_5);
nor U588 (N_588,N_256,N_352);
nor U589 (N_589,N_60,N_101);
and U590 (N_590,N_484,N_316);
or U591 (N_591,N_375,N_391);
nor U592 (N_592,N_188,N_431);
nand U593 (N_593,N_55,N_208);
or U594 (N_594,N_266,N_172);
nand U595 (N_595,N_166,N_234);
nand U596 (N_596,N_218,N_399);
nor U597 (N_597,N_138,N_359);
or U598 (N_598,N_471,N_270);
and U599 (N_599,N_378,N_48);
or U600 (N_600,N_92,N_50);
and U601 (N_601,N_472,N_374);
nor U602 (N_602,N_324,N_420);
nor U603 (N_603,N_68,N_365);
nand U604 (N_604,N_31,N_416);
and U605 (N_605,N_269,N_88);
or U606 (N_606,N_160,N_449);
and U607 (N_607,N_492,N_382);
nand U608 (N_608,N_97,N_202);
or U609 (N_609,N_70,N_496);
and U610 (N_610,N_418,N_27);
nor U611 (N_611,N_89,N_308);
or U612 (N_612,N_453,N_424);
and U613 (N_613,N_57,N_323);
and U614 (N_614,N_212,N_328);
nor U615 (N_615,N_305,N_104);
nand U616 (N_616,N_198,N_301);
nor U617 (N_617,N_77,N_91);
and U618 (N_618,N_169,N_176);
or U619 (N_619,N_38,N_242);
nand U620 (N_620,N_126,N_116);
nor U621 (N_621,N_123,N_343);
nor U622 (N_622,N_307,N_253);
nand U623 (N_623,N_6,N_321);
nand U624 (N_624,N_178,N_389);
and U625 (N_625,N_245,N_224);
and U626 (N_626,N_132,N_476);
and U627 (N_627,N_440,N_40);
nor U628 (N_628,N_25,N_425);
or U629 (N_629,N_207,N_28);
nor U630 (N_630,N_297,N_368);
nor U631 (N_631,N_474,N_35);
or U632 (N_632,N_238,N_388);
nand U633 (N_633,N_380,N_381);
nor U634 (N_634,N_42,N_216);
or U635 (N_635,N_194,N_435);
xnor U636 (N_636,N_39,N_59);
nand U637 (N_637,N_141,N_153);
nand U638 (N_638,N_452,N_360);
or U639 (N_639,N_442,N_481);
nand U640 (N_640,N_470,N_190);
nor U641 (N_641,N_318,N_20);
nand U642 (N_642,N_51,N_36);
or U643 (N_643,N_347,N_164);
nand U644 (N_644,N_175,N_232);
and U645 (N_645,N_150,N_287);
nor U646 (N_646,N_109,N_274);
nor U647 (N_647,N_299,N_465);
or U648 (N_648,N_161,N_477);
and U649 (N_649,N_248,N_125);
or U650 (N_650,N_148,N_497);
nand U651 (N_651,N_407,N_163);
or U652 (N_652,N_32,N_94);
nand U653 (N_653,N_82,N_291);
or U654 (N_654,N_330,N_251);
xor U655 (N_655,N_286,N_62);
and U656 (N_656,N_133,N_423);
and U657 (N_657,N_362,N_63);
or U658 (N_658,N_427,N_249);
nor U659 (N_659,N_469,N_144);
or U660 (N_660,N_214,N_33);
and U661 (N_661,N_311,N_180);
nor U662 (N_662,N_98,N_197);
or U663 (N_663,N_468,N_396);
and U664 (N_664,N_387,N_298);
or U665 (N_665,N_483,N_108);
nor U666 (N_666,N_326,N_265);
and U667 (N_667,N_237,N_412);
nand U668 (N_668,N_205,N_105);
or U669 (N_669,N_443,N_124);
and U670 (N_670,N_152,N_439);
and U671 (N_671,N_296,N_456);
nand U672 (N_672,N_366,N_428);
nand U673 (N_673,N_254,N_338);
or U674 (N_674,N_13,N_250);
nand U675 (N_675,N_349,N_386);
nor U676 (N_676,N_49,N_448);
nor U677 (N_677,N_261,N_426);
nor U678 (N_678,N_421,N_268);
nor U679 (N_679,N_14,N_488);
or U680 (N_680,N_340,N_414);
or U681 (N_681,N_21,N_96);
or U682 (N_682,N_403,N_390);
and U683 (N_683,N_361,N_146);
nor U684 (N_684,N_155,N_451);
and U685 (N_685,N_79,N_243);
nand U686 (N_686,N_230,N_293);
nand U687 (N_687,N_107,N_400);
nand U688 (N_688,N_72,N_106);
or U689 (N_689,N_225,N_333);
nor U690 (N_690,N_384,N_142);
nand U691 (N_691,N_454,N_222);
or U692 (N_692,N_455,N_115);
nand U693 (N_693,N_491,N_9);
and U694 (N_694,N_235,N_260);
or U695 (N_695,N_288,N_217);
or U696 (N_696,N_149,N_436);
and U697 (N_697,N_184,N_192);
or U698 (N_698,N_0,N_446);
or U699 (N_699,N_154,N_177);
nor U700 (N_700,N_24,N_459);
and U701 (N_701,N_487,N_354);
nor U702 (N_702,N_467,N_498);
or U703 (N_703,N_457,N_221);
or U704 (N_704,N_332,N_167);
or U705 (N_705,N_319,N_7);
nor U706 (N_706,N_93,N_46);
and U707 (N_707,N_397,N_147);
nand U708 (N_708,N_120,N_168);
and U709 (N_709,N_489,N_90);
and U710 (N_710,N_356,N_240);
xor U711 (N_711,N_344,N_379);
nor U712 (N_712,N_23,N_73);
and U713 (N_713,N_493,N_410);
and U714 (N_714,N_130,N_102);
and U715 (N_715,N_223,N_231);
nor U716 (N_716,N_257,N_56);
and U717 (N_717,N_44,N_16);
nor U718 (N_718,N_156,N_52);
and U719 (N_719,N_113,N_419);
nand U720 (N_720,N_12,N_187);
and U721 (N_721,N_310,N_385);
nand U722 (N_722,N_174,N_363);
nor U723 (N_723,N_482,N_285);
and U724 (N_724,N_76,N_171);
and U725 (N_725,N_314,N_404);
nor U726 (N_726,N_335,N_394);
nand U727 (N_727,N_193,N_417);
nor U728 (N_728,N_339,N_267);
nor U729 (N_729,N_429,N_258);
or U730 (N_730,N_441,N_450);
nand U731 (N_731,N_151,N_398);
or U732 (N_732,N_415,N_259);
nor U733 (N_733,N_229,N_320);
and U734 (N_734,N_475,N_336);
or U735 (N_735,N_110,N_280);
or U736 (N_736,N_358,N_10);
nor U737 (N_737,N_145,N_2);
or U738 (N_738,N_434,N_246);
and U739 (N_739,N_86,N_395);
nand U740 (N_740,N_83,N_136);
nor U741 (N_741,N_346,N_112);
and U742 (N_742,N_411,N_11);
nand U743 (N_743,N_458,N_195);
nand U744 (N_744,N_158,N_376);
nor U745 (N_745,N_58,N_233);
nor U746 (N_746,N_203,N_210);
or U747 (N_747,N_134,N_186);
nand U748 (N_748,N_74,N_284);
nor U749 (N_749,N_273,N_162);
nand U750 (N_750,N_220,N_284);
nand U751 (N_751,N_19,N_34);
or U752 (N_752,N_336,N_224);
and U753 (N_753,N_77,N_120);
nand U754 (N_754,N_343,N_13);
or U755 (N_755,N_332,N_66);
nand U756 (N_756,N_62,N_3);
or U757 (N_757,N_345,N_235);
and U758 (N_758,N_497,N_291);
and U759 (N_759,N_153,N_26);
or U760 (N_760,N_304,N_277);
nor U761 (N_761,N_448,N_116);
or U762 (N_762,N_259,N_369);
and U763 (N_763,N_91,N_6);
and U764 (N_764,N_393,N_212);
and U765 (N_765,N_29,N_281);
nor U766 (N_766,N_320,N_353);
and U767 (N_767,N_408,N_162);
or U768 (N_768,N_28,N_188);
nand U769 (N_769,N_101,N_220);
nand U770 (N_770,N_111,N_83);
nor U771 (N_771,N_333,N_475);
nor U772 (N_772,N_280,N_201);
nor U773 (N_773,N_263,N_191);
or U774 (N_774,N_25,N_73);
or U775 (N_775,N_474,N_12);
and U776 (N_776,N_409,N_254);
or U777 (N_777,N_78,N_295);
or U778 (N_778,N_100,N_99);
nor U779 (N_779,N_22,N_103);
nor U780 (N_780,N_282,N_97);
or U781 (N_781,N_174,N_38);
nor U782 (N_782,N_293,N_486);
or U783 (N_783,N_292,N_497);
and U784 (N_784,N_347,N_379);
and U785 (N_785,N_492,N_304);
or U786 (N_786,N_125,N_81);
nand U787 (N_787,N_23,N_131);
nor U788 (N_788,N_25,N_483);
or U789 (N_789,N_238,N_315);
nor U790 (N_790,N_84,N_312);
nor U791 (N_791,N_198,N_154);
and U792 (N_792,N_354,N_271);
and U793 (N_793,N_211,N_128);
nor U794 (N_794,N_86,N_189);
or U795 (N_795,N_104,N_236);
nor U796 (N_796,N_468,N_84);
or U797 (N_797,N_77,N_342);
nor U798 (N_798,N_232,N_438);
or U799 (N_799,N_374,N_156);
nand U800 (N_800,N_169,N_276);
xor U801 (N_801,N_53,N_431);
or U802 (N_802,N_472,N_256);
nand U803 (N_803,N_80,N_451);
nor U804 (N_804,N_7,N_325);
or U805 (N_805,N_179,N_79);
nand U806 (N_806,N_250,N_424);
and U807 (N_807,N_162,N_202);
and U808 (N_808,N_43,N_34);
and U809 (N_809,N_270,N_229);
and U810 (N_810,N_237,N_376);
and U811 (N_811,N_385,N_438);
and U812 (N_812,N_391,N_271);
and U813 (N_813,N_421,N_214);
and U814 (N_814,N_474,N_139);
and U815 (N_815,N_131,N_341);
nor U816 (N_816,N_412,N_486);
nor U817 (N_817,N_1,N_81);
nand U818 (N_818,N_390,N_282);
or U819 (N_819,N_440,N_136);
or U820 (N_820,N_431,N_107);
nand U821 (N_821,N_93,N_363);
or U822 (N_822,N_324,N_368);
and U823 (N_823,N_93,N_324);
and U824 (N_824,N_255,N_445);
nand U825 (N_825,N_179,N_316);
or U826 (N_826,N_236,N_370);
and U827 (N_827,N_274,N_185);
or U828 (N_828,N_479,N_210);
nor U829 (N_829,N_313,N_435);
and U830 (N_830,N_295,N_395);
nand U831 (N_831,N_228,N_67);
or U832 (N_832,N_209,N_22);
nor U833 (N_833,N_300,N_483);
or U834 (N_834,N_76,N_424);
nand U835 (N_835,N_186,N_275);
nor U836 (N_836,N_382,N_0);
and U837 (N_837,N_365,N_332);
nor U838 (N_838,N_66,N_206);
nor U839 (N_839,N_319,N_223);
and U840 (N_840,N_225,N_134);
and U841 (N_841,N_334,N_397);
or U842 (N_842,N_73,N_424);
nand U843 (N_843,N_27,N_37);
nand U844 (N_844,N_474,N_178);
or U845 (N_845,N_357,N_399);
or U846 (N_846,N_327,N_347);
nor U847 (N_847,N_251,N_448);
nor U848 (N_848,N_217,N_495);
nand U849 (N_849,N_250,N_325);
or U850 (N_850,N_193,N_106);
and U851 (N_851,N_164,N_469);
nor U852 (N_852,N_310,N_27);
xor U853 (N_853,N_295,N_105);
nand U854 (N_854,N_73,N_318);
or U855 (N_855,N_281,N_380);
nand U856 (N_856,N_304,N_409);
nand U857 (N_857,N_386,N_339);
or U858 (N_858,N_62,N_11);
or U859 (N_859,N_122,N_297);
and U860 (N_860,N_241,N_491);
nand U861 (N_861,N_492,N_347);
and U862 (N_862,N_340,N_184);
nand U863 (N_863,N_376,N_483);
nand U864 (N_864,N_471,N_428);
and U865 (N_865,N_60,N_102);
or U866 (N_866,N_489,N_285);
and U867 (N_867,N_314,N_499);
or U868 (N_868,N_252,N_193);
or U869 (N_869,N_317,N_86);
nand U870 (N_870,N_275,N_36);
nor U871 (N_871,N_252,N_473);
nor U872 (N_872,N_160,N_150);
or U873 (N_873,N_198,N_426);
nand U874 (N_874,N_351,N_276);
nor U875 (N_875,N_150,N_9);
nand U876 (N_876,N_446,N_42);
nand U877 (N_877,N_487,N_463);
and U878 (N_878,N_486,N_479);
nor U879 (N_879,N_146,N_459);
nor U880 (N_880,N_413,N_273);
and U881 (N_881,N_196,N_294);
nand U882 (N_882,N_398,N_259);
nor U883 (N_883,N_97,N_207);
or U884 (N_884,N_439,N_389);
nor U885 (N_885,N_478,N_328);
or U886 (N_886,N_262,N_449);
nor U887 (N_887,N_163,N_383);
or U888 (N_888,N_486,N_419);
nand U889 (N_889,N_119,N_337);
or U890 (N_890,N_369,N_10);
nand U891 (N_891,N_485,N_199);
nor U892 (N_892,N_129,N_334);
nand U893 (N_893,N_460,N_251);
nor U894 (N_894,N_407,N_470);
and U895 (N_895,N_424,N_10);
nand U896 (N_896,N_414,N_298);
nand U897 (N_897,N_448,N_132);
and U898 (N_898,N_353,N_464);
nor U899 (N_899,N_89,N_232);
nand U900 (N_900,N_323,N_403);
nor U901 (N_901,N_191,N_241);
or U902 (N_902,N_52,N_274);
nand U903 (N_903,N_189,N_410);
nor U904 (N_904,N_31,N_99);
and U905 (N_905,N_310,N_267);
nand U906 (N_906,N_168,N_239);
nand U907 (N_907,N_462,N_319);
and U908 (N_908,N_179,N_322);
nor U909 (N_909,N_79,N_248);
nor U910 (N_910,N_141,N_144);
or U911 (N_911,N_316,N_114);
nand U912 (N_912,N_157,N_60);
and U913 (N_913,N_161,N_285);
or U914 (N_914,N_172,N_328);
and U915 (N_915,N_307,N_80);
or U916 (N_916,N_246,N_107);
or U917 (N_917,N_161,N_24);
nand U918 (N_918,N_365,N_323);
or U919 (N_919,N_208,N_306);
and U920 (N_920,N_410,N_110);
nor U921 (N_921,N_154,N_328);
and U922 (N_922,N_425,N_338);
nor U923 (N_923,N_111,N_488);
and U924 (N_924,N_395,N_232);
nand U925 (N_925,N_418,N_60);
or U926 (N_926,N_454,N_168);
nor U927 (N_927,N_256,N_307);
or U928 (N_928,N_273,N_42);
nor U929 (N_929,N_407,N_477);
nand U930 (N_930,N_24,N_56);
or U931 (N_931,N_312,N_165);
or U932 (N_932,N_480,N_427);
or U933 (N_933,N_267,N_271);
and U934 (N_934,N_0,N_331);
and U935 (N_935,N_387,N_198);
or U936 (N_936,N_118,N_227);
and U937 (N_937,N_80,N_275);
or U938 (N_938,N_453,N_268);
nor U939 (N_939,N_263,N_133);
nand U940 (N_940,N_140,N_36);
nor U941 (N_941,N_295,N_400);
and U942 (N_942,N_284,N_58);
nor U943 (N_943,N_432,N_49);
or U944 (N_944,N_54,N_476);
nand U945 (N_945,N_308,N_433);
nand U946 (N_946,N_357,N_488);
nand U947 (N_947,N_416,N_404);
nor U948 (N_948,N_436,N_3);
and U949 (N_949,N_176,N_227);
or U950 (N_950,N_206,N_54);
nand U951 (N_951,N_78,N_494);
nor U952 (N_952,N_306,N_370);
or U953 (N_953,N_22,N_123);
nand U954 (N_954,N_30,N_23);
and U955 (N_955,N_130,N_254);
nor U956 (N_956,N_490,N_322);
and U957 (N_957,N_6,N_22);
or U958 (N_958,N_326,N_257);
nand U959 (N_959,N_496,N_348);
nand U960 (N_960,N_43,N_190);
and U961 (N_961,N_18,N_289);
or U962 (N_962,N_90,N_144);
or U963 (N_963,N_410,N_32);
nand U964 (N_964,N_348,N_293);
and U965 (N_965,N_122,N_229);
xnor U966 (N_966,N_430,N_433);
nand U967 (N_967,N_230,N_265);
and U968 (N_968,N_62,N_260);
nand U969 (N_969,N_77,N_246);
nand U970 (N_970,N_338,N_272);
or U971 (N_971,N_93,N_193);
or U972 (N_972,N_1,N_84);
and U973 (N_973,N_360,N_139);
nand U974 (N_974,N_230,N_87);
nor U975 (N_975,N_133,N_86);
or U976 (N_976,N_84,N_266);
and U977 (N_977,N_134,N_337);
or U978 (N_978,N_477,N_224);
and U979 (N_979,N_497,N_9);
nor U980 (N_980,N_13,N_84);
and U981 (N_981,N_176,N_287);
nor U982 (N_982,N_490,N_438);
nand U983 (N_983,N_25,N_476);
and U984 (N_984,N_369,N_7);
and U985 (N_985,N_330,N_369);
and U986 (N_986,N_453,N_405);
nor U987 (N_987,N_371,N_177);
nand U988 (N_988,N_135,N_98);
and U989 (N_989,N_340,N_63);
xnor U990 (N_990,N_32,N_374);
and U991 (N_991,N_492,N_56);
nand U992 (N_992,N_399,N_0);
and U993 (N_993,N_103,N_459);
or U994 (N_994,N_81,N_91);
nor U995 (N_995,N_189,N_310);
nor U996 (N_996,N_219,N_337);
nand U997 (N_997,N_378,N_253);
nor U998 (N_998,N_335,N_441);
or U999 (N_999,N_456,N_279);
nor U1000 (N_1000,N_782,N_841);
and U1001 (N_1001,N_962,N_503);
nor U1002 (N_1002,N_644,N_664);
or U1003 (N_1003,N_853,N_734);
nand U1004 (N_1004,N_639,N_974);
and U1005 (N_1005,N_945,N_653);
nor U1006 (N_1006,N_711,N_788);
nand U1007 (N_1007,N_537,N_846);
or U1008 (N_1008,N_880,N_547);
and U1009 (N_1009,N_719,N_886);
and U1010 (N_1010,N_614,N_616);
and U1011 (N_1011,N_992,N_756);
and U1012 (N_1012,N_958,N_910);
or U1013 (N_1013,N_933,N_567);
nand U1014 (N_1014,N_512,N_743);
nor U1015 (N_1015,N_517,N_584);
and U1016 (N_1016,N_666,N_918);
nand U1017 (N_1017,N_595,N_559);
nand U1018 (N_1018,N_990,N_767);
nor U1019 (N_1019,N_583,N_833);
nor U1020 (N_1020,N_681,N_835);
or U1021 (N_1021,N_546,N_942);
nor U1022 (N_1022,N_713,N_613);
nor U1023 (N_1023,N_976,N_899);
or U1024 (N_1024,N_715,N_580);
nor U1025 (N_1025,N_949,N_760);
and U1026 (N_1026,N_954,N_898);
nor U1027 (N_1027,N_520,N_722);
xnor U1028 (N_1028,N_508,N_981);
xnor U1029 (N_1029,N_998,N_912);
and U1030 (N_1030,N_634,N_564);
and U1031 (N_1031,N_731,N_971);
or U1032 (N_1032,N_861,N_550);
nor U1033 (N_1033,N_618,N_553);
and U1034 (N_1034,N_577,N_862);
and U1035 (N_1035,N_730,N_591);
nor U1036 (N_1036,N_592,N_852);
nor U1037 (N_1037,N_600,N_645);
nand U1038 (N_1038,N_891,N_959);
nand U1039 (N_1039,N_643,N_611);
nand U1040 (N_1040,N_540,N_854);
nor U1041 (N_1041,N_604,N_972);
nand U1042 (N_1042,N_935,N_778);
nand U1043 (N_1043,N_516,N_802);
or U1044 (N_1044,N_948,N_624);
or U1045 (N_1045,N_951,N_510);
nand U1046 (N_1046,N_904,N_741);
nand U1047 (N_1047,N_915,N_527);
and U1048 (N_1048,N_876,N_863);
or U1049 (N_1049,N_578,N_628);
and U1050 (N_1050,N_661,N_947);
nor U1051 (N_1051,N_548,N_748);
or U1052 (N_1052,N_896,N_800);
nor U1053 (N_1053,N_562,N_890);
nor U1054 (N_1054,N_685,N_809);
and U1055 (N_1055,N_968,N_997);
or U1056 (N_1056,N_630,N_593);
nor U1057 (N_1057,N_795,N_502);
or U1058 (N_1058,N_830,N_667);
or U1059 (N_1059,N_554,N_594);
and U1060 (N_1060,N_928,N_957);
or U1061 (N_1061,N_786,N_813);
nor U1062 (N_1062,N_768,N_825);
or U1063 (N_1063,N_921,N_569);
xnor U1064 (N_1064,N_894,N_943);
and U1065 (N_1065,N_574,N_626);
or U1066 (N_1066,N_859,N_827);
nand U1067 (N_1067,N_588,N_521);
and U1068 (N_1068,N_680,N_615);
nor U1069 (N_1069,N_934,N_999);
and U1070 (N_1070,N_961,N_944);
and U1071 (N_1071,N_761,N_893);
and U1072 (N_1072,N_837,N_638);
nor U1073 (N_1073,N_905,N_586);
and U1074 (N_1074,N_621,N_987);
nand U1075 (N_1075,N_845,N_532);
and U1076 (N_1076,N_623,N_581);
nand U1077 (N_1077,N_609,N_602);
nor U1078 (N_1078,N_919,N_705);
or U1079 (N_1079,N_884,N_885);
and U1080 (N_1080,N_975,N_729);
nand U1081 (N_1081,N_668,N_513);
nand U1082 (N_1082,N_920,N_526);
nand U1083 (N_1083,N_946,N_892);
or U1084 (N_1084,N_849,N_829);
nor U1085 (N_1085,N_690,N_907);
nand U1086 (N_1086,N_950,N_763);
nor U1087 (N_1087,N_608,N_599);
and U1088 (N_1088,N_978,N_828);
and U1089 (N_1089,N_877,N_582);
nor U1090 (N_1090,N_575,N_983);
or U1091 (N_1091,N_710,N_777);
xnor U1092 (N_1092,N_989,N_860);
nor U1093 (N_1093,N_847,N_814);
nor U1094 (N_1094,N_585,N_775);
or U1095 (N_1095,N_881,N_673);
nand U1096 (N_1096,N_511,N_789);
nand U1097 (N_1097,N_816,N_901);
and U1098 (N_1098,N_798,N_683);
nand U1099 (N_1099,N_679,N_738);
nand U1100 (N_1100,N_771,N_820);
and U1101 (N_1101,N_783,N_514);
nor U1102 (N_1102,N_790,N_796);
or U1103 (N_1103,N_808,N_631);
and U1104 (N_1104,N_721,N_652);
nor U1105 (N_1105,N_751,N_530);
or U1106 (N_1106,N_888,N_801);
or U1107 (N_1107,N_823,N_563);
and U1108 (N_1108,N_762,N_501);
nand U1109 (N_1109,N_541,N_504);
and U1110 (N_1110,N_807,N_507);
and U1111 (N_1111,N_878,N_804);
nand U1112 (N_1112,N_793,N_803);
nand U1113 (N_1113,N_648,N_923);
xnor U1114 (N_1114,N_936,N_686);
or U1115 (N_1115,N_701,N_691);
xor U1116 (N_1116,N_996,N_766);
or U1117 (N_1117,N_579,N_826);
nand U1118 (N_1118,N_662,N_576);
nor U1119 (N_1119,N_620,N_839);
or U1120 (N_1120,N_857,N_965);
nor U1121 (N_1121,N_744,N_682);
or U1122 (N_1122,N_650,N_570);
nor U1123 (N_1123,N_696,N_925);
and U1124 (N_1124,N_676,N_769);
nor U1125 (N_1125,N_779,N_855);
or U1126 (N_1126,N_560,N_797);
or U1127 (N_1127,N_703,N_746);
or U1128 (N_1128,N_688,N_674);
nor U1129 (N_1129,N_873,N_874);
or U1130 (N_1130,N_566,N_720);
or U1131 (N_1131,N_843,N_952);
nor U1132 (N_1132,N_557,N_969);
or U1133 (N_1133,N_571,N_597);
nor U1134 (N_1134,N_723,N_817);
nand U1135 (N_1135,N_812,N_709);
nand U1136 (N_1136,N_538,N_655);
nor U1137 (N_1137,N_757,N_551);
or U1138 (N_1138,N_818,N_635);
nor U1139 (N_1139,N_770,N_519);
nor U1140 (N_1140,N_887,N_754);
nor U1141 (N_1141,N_821,N_840);
nand U1142 (N_1142,N_544,N_642);
nand U1143 (N_1143,N_646,N_908);
nand U1144 (N_1144,N_883,N_824);
and U1145 (N_1145,N_932,N_742);
nand U1146 (N_1146,N_543,N_970);
nand U1147 (N_1147,N_692,N_780);
and U1148 (N_1148,N_900,N_589);
nand U1149 (N_1149,N_749,N_733);
or U1150 (N_1150,N_759,N_601);
or U1151 (N_1151,N_930,N_700);
and U1152 (N_1152,N_806,N_776);
nor U1153 (N_1153,N_953,N_606);
nand U1154 (N_1154,N_714,N_500);
and U1155 (N_1155,N_663,N_509);
nor U1156 (N_1156,N_963,N_895);
nor U1157 (N_1157,N_993,N_922);
and U1158 (N_1158,N_549,N_607);
and U1159 (N_1159,N_505,N_805);
and U1160 (N_1160,N_791,N_697);
nor U1161 (N_1161,N_740,N_794);
and U1162 (N_1162,N_656,N_792);
nor U1163 (N_1163,N_964,N_529);
or U1164 (N_1164,N_637,N_672);
nor U1165 (N_1165,N_707,N_758);
or U1166 (N_1166,N_747,N_590);
nand U1167 (N_1167,N_955,N_931);
nand U1168 (N_1168,N_605,N_651);
nand U1169 (N_1169,N_725,N_670);
or U1170 (N_1170,N_773,N_870);
nor U1171 (N_1171,N_534,N_524);
or U1172 (N_1172,N_882,N_665);
nor U1173 (N_1173,N_702,N_572);
and U1174 (N_1174,N_764,N_938);
nand U1175 (N_1175,N_610,N_675);
nor U1176 (N_1176,N_629,N_909);
and U1177 (N_1177,N_871,N_832);
nor U1178 (N_1178,N_525,N_752);
nor U1179 (N_1179,N_985,N_924);
nand U1180 (N_1180,N_716,N_596);
or U1181 (N_1181,N_755,N_658);
or U1182 (N_1182,N_929,N_869);
nand U1183 (N_1183,N_506,N_879);
nor U1184 (N_1184,N_864,N_772);
nor U1185 (N_1185,N_659,N_850);
nand U1186 (N_1186,N_657,N_939);
and U1187 (N_1187,N_875,N_556);
nand U1188 (N_1188,N_906,N_718);
and U1189 (N_1189,N_535,N_649);
and U1190 (N_1190,N_986,N_897);
nand U1191 (N_1191,N_889,N_539);
nor U1192 (N_1192,N_982,N_784);
or U1193 (N_1193,N_868,N_984);
or U1194 (N_1194,N_858,N_712);
nor U1195 (N_1195,N_937,N_727);
nand U1196 (N_1196,N_917,N_979);
nor U1197 (N_1197,N_926,N_515);
or U1198 (N_1198,N_552,N_956);
nand U1199 (N_1199,N_617,N_724);
nor U1200 (N_1200,N_636,N_811);
nor U1201 (N_1201,N_647,N_916);
and U1202 (N_1202,N_528,N_531);
nand U1203 (N_1203,N_695,N_678);
or U1204 (N_1204,N_732,N_834);
or U1205 (N_1205,N_573,N_684);
nand U1206 (N_1206,N_641,N_911);
or U1207 (N_1207,N_977,N_603);
nor U1208 (N_1208,N_848,N_598);
nor U1209 (N_1209,N_633,N_851);
nand U1210 (N_1210,N_698,N_866);
and U1211 (N_1211,N_903,N_810);
or U1212 (N_1212,N_536,N_728);
and U1213 (N_1213,N_842,N_980);
and U1214 (N_1214,N_902,N_941);
or U1215 (N_1215,N_708,N_872);
or U1216 (N_1216,N_522,N_736);
nand U1217 (N_1217,N_561,N_838);
and U1218 (N_1218,N_991,N_960);
xor U1219 (N_1219,N_787,N_627);
nand U1220 (N_1220,N_671,N_545);
or U1221 (N_1221,N_967,N_587);
nand U1222 (N_1222,N_704,N_677);
nand U1223 (N_1223,N_815,N_927);
nor U1224 (N_1224,N_785,N_774);
and U1225 (N_1225,N_753,N_717);
or U1226 (N_1226,N_737,N_669);
nor U1227 (N_1227,N_632,N_856);
nand U1228 (N_1228,N_568,N_619);
nand U1229 (N_1229,N_867,N_660);
nand U1230 (N_1230,N_558,N_625);
or U1231 (N_1231,N_523,N_654);
nor U1232 (N_1232,N_865,N_687);
nor U1233 (N_1233,N_699,N_799);
nand U1234 (N_1234,N_542,N_706);
nor U1235 (N_1235,N_940,N_994);
nand U1236 (N_1236,N_913,N_735);
nor U1237 (N_1237,N_844,N_819);
nor U1238 (N_1238,N_966,N_822);
nand U1239 (N_1239,N_518,N_689);
nor U1240 (N_1240,N_693,N_533);
or U1241 (N_1241,N_622,N_914);
or U1242 (N_1242,N_694,N_565);
or U1243 (N_1243,N_739,N_831);
and U1244 (N_1244,N_988,N_726);
and U1245 (N_1245,N_555,N_612);
xor U1246 (N_1246,N_995,N_765);
or U1247 (N_1247,N_781,N_745);
or U1248 (N_1248,N_640,N_750);
and U1249 (N_1249,N_973,N_836);
or U1250 (N_1250,N_868,N_927);
or U1251 (N_1251,N_749,N_934);
nand U1252 (N_1252,N_537,N_941);
and U1253 (N_1253,N_912,N_583);
nor U1254 (N_1254,N_620,N_920);
nand U1255 (N_1255,N_899,N_658);
and U1256 (N_1256,N_819,N_700);
nor U1257 (N_1257,N_745,N_839);
nor U1258 (N_1258,N_816,N_561);
and U1259 (N_1259,N_951,N_976);
or U1260 (N_1260,N_526,N_820);
and U1261 (N_1261,N_501,N_933);
nand U1262 (N_1262,N_901,N_652);
and U1263 (N_1263,N_503,N_935);
or U1264 (N_1264,N_542,N_525);
nand U1265 (N_1265,N_862,N_799);
nand U1266 (N_1266,N_899,N_794);
or U1267 (N_1267,N_905,N_757);
and U1268 (N_1268,N_549,N_975);
or U1269 (N_1269,N_850,N_800);
nor U1270 (N_1270,N_680,N_965);
nand U1271 (N_1271,N_946,N_548);
or U1272 (N_1272,N_981,N_916);
or U1273 (N_1273,N_951,N_842);
nor U1274 (N_1274,N_790,N_918);
nor U1275 (N_1275,N_773,N_679);
nor U1276 (N_1276,N_715,N_567);
or U1277 (N_1277,N_758,N_588);
or U1278 (N_1278,N_765,N_759);
and U1279 (N_1279,N_952,N_769);
or U1280 (N_1280,N_596,N_768);
nand U1281 (N_1281,N_534,N_543);
xnor U1282 (N_1282,N_619,N_873);
and U1283 (N_1283,N_679,N_889);
or U1284 (N_1284,N_882,N_744);
and U1285 (N_1285,N_891,N_545);
or U1286 (N_1286,N_862,N_863);
and U1287 (N_1287,N_751,N_705);
nand U1288 (N_1288,N_734,N_711);
or U1289 (N_1289,N_910,N_705);
or U1290 (N_1290,N_904,N_962);
or U1291 (N_1291,N_923,N_590);
and U1292 (N_1292,N_861,N_507);
or U1293 (N_1293,N_724,N_501);
nor U1294 (N_1294,N_709,N_623);
and U1295 (N_1295,N_859,N_948);
or U1296 (N_1296,N_735,N_742);
nor U1297 (N_1297,N_809,N_915);
nor U1298 (N_1298,N_584,N_925);
or U1299 (N_1299,N_520,N_915);
nor U1300 (N_1300,N_763,N_854);
nor U1301 (N_1301,N_799,N_882);
nand U1302 (N_1302,N_966,N_983);
and U1303 (N_1303,N_711,N_816);
or U1304 (N_1304,N_740,N_532);
or U1305 (N_1305,N_773,N_536);
or U1306 (N_1306,N_953,N_652);
or U1307 (N_1307,N_519,N_504);
nor U1308 (N_1308,N_521,N_991);
nand U1309 (N_1309,N_540,N_861);
nor U1310 (N_1310,N_728,N_724);
or U1311 (N_1311,N_587,N_934);
nor U1312 (N_1312,N_815,N_882);
and U1313 (N_1313,N_922,N_750);
nor U1314 (N_1314,N_507,N_872);
nand U1315 (N_1315,N_880,N_613);
or U1316 (N_1316,N_730,N_986);
or U1317 (N_1317,N_531,N_917);
xor U1318 (N_1318,N_806,N_975);
and U1319 (N_1319,N_608,N_561);
nor U1320 (N_1320,N_607,N_852);
or U1321 (N_1321,N_817,N_505);
nor U1322 (N_1322,N_824,N_884);
nor U1323 (N_1323,N_584,N_519);
or U1324 (N_1324,N_592,N_907);
nor U1325 (N_1325,N_854,N_920);
and U1326 (N_1326,N_557,N_517);
and U1327 (N_1327,N_833,N_993);
nand U1328 (N_1328,N_562,N_788);
or U1329 (N_1329,N_606,N_923);
or U1330 (N_1330,N_877,N_967);
nand U1331 (N_1331,N_917,N_816);
nor U1332 (N_1332,N_600,N_899);
nor U1333 (N_1333,N_992,N_582);
nand U1334 (N_1334,N_863,N_534);
and U1335 (N_1335,N_828,N_561);
nor U1336 (N_1336,N_910,N_819);
and U1337 (N_1337,N_548,N_966);
nor U1338 (N_1338,N_913,N_739);
and U1339 (N_1339,N_712,N_949);
nand U1340 (N_1340,N_643,N_699);
and U1341 (N_1341,N_826,N_985);
nor U1342 (N_1342,N_686,N_839);
nor U1343 (N_1343,N_817,N_708);
nand U1344 (N_1344,N_919,N_620);
nor U1345 (N_1345,N_629,N_925);
nand U1346 (N_1346,N_666,N_682);
nand U1347 (N_1347,N_813,N_821);
or U1348 (N_1348,N_765,N_571);
and U1349 (N_1349,N_725,N_863);
or U1350 (N_1350,N_984,N_816);
and U1351 (N_1351,N_627,N_749);
or U1352 (N_1352,N_636,N_909);
nand U1353 (N_1353,N_876,N_773);
nor U1354 (N_1354,N_843,N_901);
or U1355 (N_1355,N_871,N_712);
nand U1356 (N_1356,N_848,N_504);
or U1357 (N_1357,N_741,N_685);
and U1358 (N_1358,N_829,N_554);
and U1359 (N_1359,N_995,N_855);
nor U1360 (N_1360,N_965,N_837);
nor U1361 (N_1361,N_749,N_806);
nor U1362 (N_1362,N_883,N_600);
nand U1363 (N_1363,N_761,N_869);
nand U1364 (N_1364,N_980,N_840);
nand U1365 (N_1365,N_976,N_658);
and U1366 (N_1366,N_631,N_682);
nor U1367 (N_1367,N_625,N_631);
nor U1368 (N_1368,N_614,N_722);
or U1369 (N_1369,N_966,N_529);
and U1370 (N_1370,N_864,N_611);
nor U1371 (N_1371,N_637,N_775);
or U1372 (N_1372,N_552,N_682);
nor U1373 (N_1373,N_940,N_698);
nor U1374 (N_1374,N_707,N_922);
or U1375 (N_1375,N_570,N_751);
nor U1376 (N_1376,N_604,N_869);
or U1377 (N_1377,N_740,N_664);
and U1378 (N_1378,N_794,N_606);
or U1379 (N_1379,N_683,N_862);
or U1380 (N_1380,N_537,N_956);
and U1381 (N_1381,N_876,N_662);
nand U1382 (N_1382,N_745,N_732);
or U1383 (N_1383,N_567,N_562);
nand U1384 (N_1384,N_867,N_862);
and U1385 (N_1385,N_906,N_994);
and U1386 (N_1386,N_654,N_741);
or U1387 (N_1387,N_534,N_619);
and U1388 (N_1388,N_828,N_527);
nand U1389 (N_1389,N_574,N_760);
or U1390 (N_1390,N_831,N_864);
nand U1391 (N_1391,N_720,N_808);
nor U1392 (N_1392,N_736,N_533);
nand U1393 (N_1393,N_599,N_832);
or U1394 (N_1394,N_928,N_672);
nor U1395 (N_1395,N_951,N_697);
or U1396 (N_1396,N_612,N_959);
nand U1397 (N_1397,N_911,N_763);
or U1398 (N_1398,N_760,N_634);
and U1399 (N_1399,N_691,N_930);
nor U1400 (N_1400,N_527,N_726);
nand U1401 (N_1401,N_883,N_548);
nand U1402 (N_1402,N_835,N_778);
or U1403 (N_1403,N_620,N_661);
nand U1404 (N_1404,N_590,N_518);
nand U1405 (N_1405,N_855,N_694);
nor U1406 (N_1406,N_723,N_527);
nor U1407 (N_1407,N_579,N_628);
nor U1408 (N_1408,N_586,N_984);
or U1409 (N_1409,N_828,N_649);
nor U1410 (N_1410,N_786,N_826);
nand U1411 (N_1411,N_854,N_771);
or U1412 (N_1412,N_671,N_836);
nor U1413 (N_1413,N_916,N_955);
nand U1414 (N_1414,N_608,N_713);
and U1415 (N_1415,N_574,N_754);
or U1416 (N_1416,N_548,N_817);
and U1417 (N_1417,N_599,N_621);
and U1418 (N_1418,N_625,N_766);
and U1419 (N_1419,N_713,N_575);
and U1420 (N_1420,N_782,N_673);
and U1421 (N_1421,N_767,N_936);
or U1422 (N_1422,N_826,N_967);
nor U1423 (N_1423,N_563,N_874);
or U1424 (N_1424,N_623,N_626);
nor U1425 (N_1425,N_578,N_664);
or U1426 (N_1426,N_532,N_536);
nand U1427 (N_1427,N_551,N_556);
or U1428 (N_1428,N_674,N_696);
nand U1429 (N_1429,N_864,N_539);
and U1430 (N_1430,N_796,N_649);
nand U1431 (N_1431,N_797,N_782);
and U1432 (N_1432,N_600,N_830);
nand U1433 (N_1433,N_732,N_726);
and U1434 (N_1434,N_978,N_850);
nand U1435 (N_1435,N_829,N_621);
nor U1436 (N_1436,N_670,N_625);
and U1437 (N_1437,N_993,N_733);
nand U1438 (N_1438,N_809,N_528);
or U1439 (N_1439,N_812,N_813);
and U1440 (N_1440,N_754,N_685);
or U1441 (N_1441,N_651,N_568);
nand U1442 (N_1442,N_534,N_563);
or U1443 (N_1443,N_946,N_722);
nand U1444 (N_1444,N_570,N_913);
or U1445 (N_1445,N_621,N_514);
xor U1446 (N_1446,N_577,N_852);
nand U1447 (N_1447,N_564,N_984);
nor U1448 (N_1448,N_929,N_611);
nand U1449 (N_1449,N_818,N_629);
or U1450 (N_1450,N_881,N_716);
and U1451 (N_1451,N_811,N_884);
nand U1452 (N_1452,N_707,N_611);
and U1453 (N_1453,N_589,N_871);
and U1454 (N_1454,N_921,N_641);
nand U1455 (N_1455,N_926,N_599);
or U1456 (N_1456,N_634,N_622);
nand U1457 (N_1457,N_640,N_718);
nand U1458 (N_1458,N_811,N_539);
nand U1459 (N_1459,N_794,N_502);
or U1460 (N_1460,N_546,N_964);
nand U1461 (N_1461,N_907,N_633);
nor U1462 (N_1462,N_789,N_890);
nand U1463 (N_1463,N_519,N_680);
and U1464 (N_1464,N_686,N_707);
nand U1465 (N_1465,N_928,N_516);
nand U1466 (N_1466,N_569,N_919);
nor U1467 (N_1467,N_562,N_605);
or U1468 (N_1468,N_567,N_665);
or U1469 (N_1469,N_632,N_868);
and U1470 (N_1470,N_611,N_924);
and U1471 (N_1471,N_967,N_595);
or U1472 (N_1472,N_877,N_884);
and U1473 (N_1473,N_561,N_525);
and U1474 (N_1474,N_647,N_558);
or U1475 (N_1475,N_767,N_620);
nor U1476 (N_1476,N_570,N_707);
nand U1477 (N_1477,N_629,N_567);
nand U1478 (N_1478,N_717,N_822);
and U1479 (N_1479,N_553,N_749);
nor U1480 (N_1480,N_538,N_615);
nand U1481 (N_1481,N_792,N_902);
and U1482 (N_1482,N_994,N_791);
or U1483 (N_1483,N_609,N_775);
or U1484 (N_1484,N_695,N_921);
nor U1485 (N_1485,N_578,N_799);
or U1486 (N_1486,N_752,N_697);
or U1487 (N_1487,N_507,N_547);
nor U1488 (N_1488,N_671,N_957);
nand U1489 (N_1489,N_844,N_681);
nor U1490 (N_1490,N_703,N_529);
and U1491 (N_1491,N_864,N_558);
nand U1492 (N_1492,N_865,N_835);
nand U1493 (N_1493,N_558,N_666);
or U1494 (N_1494,N_765,N_808);
nand U1495 (N_1495,N_816,N_518);
nand U1496 (N_1496,N_964,N_592);
and U1497 (N_1497,N_649,N_978);
or U1498 (N_1498,N_697,N_997);
or U1499 (N_1499,N_864,N_970);
nand U1500 (N_1500,N_1393,N_1196);
and U1501 (N_1501,N_1285,N_1403);
nand U1502 (N_1502,N_1370,N_1060);
and U1503 (N_1503,N_1088,N_1014);
nor U1504 (N_1504,N_1408,N_1070);
nor U1505 (N_1505,N_1349,N_1449);
nor U1506 (N_1506,N_1202,N_1025);
nand U1507 (N_1507,N_1033,N_1359);
and U1508 (N_1508,N_1276,N_1032);
nor U1509 (N_1509,N_1068,N_1290);
and U1510 (N_1510,N_1004,N_1081);
nor U1511 (N_1511,N_1394,N_1007);
nand U1512 (N_1512,N_1227,N_1369);
nor U1513 (N_1513,N_1392,N_1065);
or U1514 (N_1514,N_1079,N_1071);
or U1515 (N_1515,N_1429,N_1288);
or U1516 (N_1516,N_1256,N_1150);
and U1517 (N_1517,N_1265,N_1261);
nand U1518 (N_1518,N_1303,N_1248);
nor U1519 (N_1519,N_1054,N_1270);
or U1520 (N_1520,N_1472,N_1491);
nand U1521 (N_1521,N_1199,N_1286);
and U1522 (N_1522,N_1277,N_1149);
nor U1523 (N_1523,N_1192,N_1105);
or U1524 (N_1524,N_1010,N_1380);
or U1525 (N_1525,N_1053,N_1419);
and U1526 (N_1526,N_1425,N_1254);
nand U1527 (N_1527,N_1201,N_1047);
or U1528 (N_1528,N_1271,N_1113);
nor U1529 (N_1529,N_1005,N_1336);
or U1530 (N_1530,N_1385,N_1367);
or U1531 (N_1531,N_1397,N_1405);
nor U1532 (N_1532,N_1305,N_1095);
and U1533 (N_1533,N_1215,N_1282);
and U1534 (N_1534,N_1445,N_1440);
nor U1535 (N_1535,N_1019,N_1387);
nand U1536 (N_1536,N_1187,N_1330);
or U1537 (N_1537,N_1211,N_1224);
or U1538 (N_1538,N_1326,N_1153);
nand U1539 (N_1539,N_1448,N_1465);
nand U1540 (N_1540,N_1024,N_1441);
and U1541 (N_1541,N_1361,N_1300);
nand U1542 (N_1542,N_1189,N_1168);
and U1543 (N_1543,N_1239,N_1173);
nor U1544 (N_1544,N_1076,N_1127);
nor U1545 (N_1545,N_1297,N_1116);
nor U1546 (N_1546,N_1100,N_1308);
and U1547 (N_1547,N_1052,N_1471);
nand U1548 (N_1548,N_1075,N_1186);
nor U1549 (N_1549,N_1135,N_1030);
nand U1550 (N_1550,N_1073,N_1041);
nor U1551 (N_1551,N_1158,N_1258);
and U1552 (N_1552,N_1238,N_1147);
nand U1553 (N_1553,N_1077,N_1456);
or U1554 (N_1554,N_1118,N_1307);
or U1555 (N_1555,N_1123,N_1094);
and U1556 (N_1556,N_1103,N_1119);
nor U1557 (N_1557,N_1412,N_1063);
nor U1558 (N_1558,N_1083,N_1011);
nor U1559 (N_1559,N_1344,N_1437);
nor U1560 (N_1560,N_1411,N_1244);
and U1561 (N_1561,N_1241,N_1329);
or U1562 (N_1562,N_1365,N_1036);
nand U1563 (N_1563,N_1314,N_1049);
and U1564 (N_1564,N_1249,N_1318);
nand U1565 (N_1565,N_1353,N_1000);
nand U1566 (N_1566,N_1454,N_1266);
or U1567 (N_1567,N_1001,N_1120);
and U1568 (N_1568,N_1428,N_1480);
and U1569 (N_1569,N_1096,N_1252);
nand U1570 (N_1570,N_1421,N_1031);
nand U1571 (N_1571,N_1023,N_1046);
nor U1572 (N_1572,N_1486,N_1287);
and U1573 (N_1573,N_1058,N_1346);
or U1574 (N_1574,N_1184,N_1133);
or U1575 (N_1575,N_1231,N_1461);
and U1576 (N_1576,N_1163,N_1279);
and U1577 (N_1577,N_1495,N_1057);
and U1578 (N_1578,N_1061,N_1274);
nor U1579 (N_1579,N_1229,N_1435);
and U1580 (N_1580,N_1432,N_1386);
nor U1581 (N_1581,N_1328,N_1460);
nand U1582 (N_1582,N_1175,N_1354);
nor U1583 (N_1583,N_1193,N_1458);
nor U1584 (N_1584,N_1391,N_1414);
or U1585 (N_1585,N_1423,N_1453);
nand U1586 (N_1586,N_1469,N_1131);
nor U1587 (N_1587,N_1475,N_1015);
or U1588 (N_1588,N_1051,N_1289);
nand U1589 (N_1589,N_1212,N_1137);
or U1590 (N_1590,N_1398,N_1451);
and U1591 (N_1591,N_1371,N_1124);
and U1592 (N_1592,N_1132,N_1037);
nor U1593 (N_1593,N_1101,N_1395);
nand U1594 (N_1594,N_1228,N_1223);
xnor U1595 (N_1595,N_1402,N_1415);
nor U1596 (N_1596,N_1216,N_1204);
nor U1597 (N_1597,N_1427,N_1008);
and U1598 (N_1598,N_1375,N_1164);
and U1599 (N_1599,N_1165,N_1358);
nand U1600 (N_1600,N_1012,N_1337);
and U1601 (N_1601,N_1309,N_1170);
nand U1602 (N_1602,N_1172,N_1038);
and U1603 (N_1603,N_1160,N_1488);
nor U1604 (N_1604,N_1301,N_1139);
or U1605 (N_1605,N_1409,N_1484);
nor U1606 (N_1606,N_1479,N_1293);
and U1607 (N_1607,N_1413,N_1436);
or U1608 (N_1608,N_1138,N_1457);
and U1609 (N_1609,N_1197,N_1226);
nor U1610 (N_1610,N_1478,N_1292);
nand U1611 (N_1611,N_1040,N_1462);
and U1612 (N_1612,N_1322,N_1169);
and U1613 (N_1613,N_1230,N_1264);
nor U1614 (N_1614,N_1373,N_1157);
or U1615 (N_1615,N_1129,N_1232);
nor U1616 (N_1616,N_1390,N_1207);
or U1617 (N_1617,N_1340,N_1098);
nor U1618 (N_1618,N_1464,N_1039);
nand U1619 (N_1619,N_1306,N_1243);
or U1620 (N_1620,N_1166,N_1059);
nand U1621 (N_1621,N_1210,N_1066);
or U1622 (N_1622,N_1018,N_1179);
nand U1623 (N_1623,N_1302,N_1283);
nor U1624 (N_1624,N_1209,N_1284);
nand U1625 (N_1625,N_1259,N_1388);
or U1626 (N_1626,N_1143,N_1316);
or U1627 (N_1627,N_1152,N_1363);
and U1628 (N_1628,N_1177,N_1273);
and U1629 (N_1629,N_1242,N_1443);
or U1630 (N_1630,N_1108,N_1250);
nor U1631 (N_1631,N_1022,N_1222);
nor U1632 (N_1632,N_1320,N_1317);
nor U1633 (N_1633,N_1325,N_1418);
nand U1634 (N_1634,N_1122,N_1217);
nor U1635 (N_1635,N_1017,N_1466);
nor U1636 (N_1636,N_1121,N_1278);
and U1637 (N_1637,N_1183,N_1102);
nor U1638 (N_1638,N_1218,N_1442);
and U1639 (N_1639,N_1013,N_1020);
xnor U1640 (N_1640,N_1396,N_1235);
nand U1641 (N_1641,N_1294,N_1378);
nand U1642 (N_1642,N_1364,N_1195);
or U1643 (N_1643,N_1404,N_1474);
and U1644 (N_1644,N_1112,N_1490);
and U1645 (N_1645,N_1281,N_1084);
nand U1646 (N_1646,N_1482,N_1110);
nor U1647 (N_1647,N_1009,N_1422);
and U1648 (N_1648,N_1027,N_1089);
and U1649 (N_1649,N_1029,N_1191);
and U1650 (N_1650,N_1247,N_1452);
and U1651 (N_1651,N_1481,N_1406);
and U1652 (N_1652,N_1087,N_1144);
and U1653 (N_1653,N_1091,N_1269);
nand U1654 (N_1654,N_1450,N_1497);
xnor U1655 (N_1655,N_1171,N_1140);
nor U1656 (N_1656,N_1323,N_1048);
xnor U1657 (N_1657,N_1026,N_1220);
and U1658 (N_1658,N_1080,N_1006);
and U1659 (N_1659,N_1181,N_1180);
or U1660 (N_1660,N_1214,N_1174);
or U1661 (N_1661,N_1221,N_1485);
and U1662 (N_1662,N_1352,N_1494);
and U1663 (N_1663,N_1348,N_1304);
nor U1664 (N_1664,N_1275,N_1003);
nor U1665 (N_1665,N_1034,N_1377);
or U1666 (N_1666,N_1342,N_1257);
nor U1667 (N_1667,N_1155,N_1470);
or U1668 (N_1668,N_1324,N_1280);
or U1669 (N_1669,N_1489,N_1115);
and U1670 (N_1670,N_1295,N_1416);
and U1671 (N_1671,N_1381,N_1355);
and U1672 (N_1672,N_1267,N_1447);
nand U1673 (N_1673,N_1296,N_1347);
nand U1674 (N_1674,N_1374,N_1114);
and U1675 (N_1675,N_1107,N_1345);
nor U1676 (N_1676,N_1128,N_1360);
or U1677 (N_1677,N_1233,N_1044);
nor U1678 (N_1678,N_1251,N_1142);
or U1679 (N_1679,N_1148,N_1321);
nand U1680 (N_1680,N_1298,N_1439);
and U1681 (N_1681,N_1327,N_1104);
nand U1682 (N_1682,N_1069,N_1382);
and U1683 (N_1683,N_1263,N_1126);
or U1684 (N_1684,N_1255,N_1268);
xnor U1685 (N_1685,N_1473,N_1332);
or U1686 (N_1686,N_1424,N_1438);
or U1687 (N_1687,N_1028,N_1161);
nor U1688 (N_1688,N_1198,N_1384);
and U1689 (N_1689,N_1400,N_1072);
or U1690 (N_1690,N_1136,N_1185);
and U1691 (N_1691,N_1097,N_1067);
and U1692 (N_1692,N_1130,N_1182);
and U1693 (N_1693,N_1343,N_1426);
or U1694 (N_1694,N_1085,N_1372);
and U1695 (N_1695,N_1357,N_1433);
nand U1696 (N_1696,N_1246,N_1154);
or U1697 (N_1697,N_1141,N_1056);
nand U1698 (N_1698,N_1237,N_1236);
nor U1699 (N_1699,N_1351,N_1253);
nand U1700 (N_1700,N_1078,N_1090);
and U1701 (N_1701,N_1335,N_1167);
or U1702 (N_1702,N_1042,N_1319);
or U1703 (N_1703,N_1002,N_1106);
or U1704 (N_1704,N_1206,N_1176);
and U1705 (N_1705,N_1455,N_1313);
or U1706 (N_1706,N_1134,N_1109);
nor U1707 (N_1707,N_1219,N_1366);
nor U1708 (N_1708,N_1299,N_1315);
and U1709 (N_1709,N_1389,N_1074);
xnor U1710 (N_1710,N_1272,N_1499);
nand U1711 (N_1711,N_1356,N_1213);
nor U1712 (N_1712,N_1021,N_1434);
or U1713 (N_1713,N_1368,N_1468);
nor U1714 (N_1714,N_1162,N_1062);
and U1715 (N_1715,N_1092,N_1420);
or U1716 (N_1716,N_1341,N_1417);
nor U1717 (N_1717,N_1483,N_1093);
nand U1718 (N_1718,N_1099,N_1159);
or U1719 (N_1719,N_1498,N_1446);
nor U1720 (N_1720,N_1262,N_1496);
or U1721 (N_1721,N_1260,N_1151);
nor U1722 (N_1722,N_1203,N_1043);
xor U1723 (N_1723,N_1476,N_1156);
nor U1724 (N_1724,N_1362,N_1125);
nor U1725 (N_1725,N_1379,N_1050);
nor U1726 (N_1726,N_1410,N_1376);
and U1727 (N_1727,N_1055,N_1016);
nand U1728 (N_1728,N_1111,N_1492);
nand U1729 (N_1729,N_1045,N_1401);
and U1730 (N_1730,N_1086,N_1178);
and U1731 (N_1731,N_1487,N_1117);
or U1732 (N_1732,N_1208,N_1467);
and U1733 (N_1733,N_1245,N_1240);
or U1734 (N_1734,N_1311,N_1225);
nand U1735 (N_1735,N_1035,N_1064);
nor U1736 (N_1736,N_1334,N_1459);
nand U1737 (N_1737,N_1145,N_1399);
nor U1738 (N_1738,N_1310,N_1444);
xnor U1739 (N_1739,N_1146,N_1188);
nor U1740 (N_1740,N_1200,N_1190);
and U1741 (N_1741,N_1333,N_1430);
and U1742 (N_1742,N_1338,N_1082);
nand U1743 (N_1743,N_1493,N_1291);
nand U1744 (N_1744,N_1194,N_1331);
or U1745 (N_1745,N_1205,N_1431);
and U1746 (N_1746,N_1312,N_1350);
or U1747 (N_1747,N_1463,N_1339);
nor U1748 (N_1748,N_1383,N_1234);
nor U1749 (N_1749,N_1477,N_1407);
and U1750 (N_1750,N_1197,N_1010);
nand U1751 (N_1751,N_1056,N_1360);
and U1752 (N_1752,N_1304,N_1104);
nand U1753 (N_1753,N_1450,N_1266);
nand U1754 (N_1754,N_1178,N_1367);
and U1755 (N_1755,N_1238,N_1381);
nand U1756 (N_1756,N_1101,N_1115);
nand U1757 (N_1757,N_1098,N_1026);
and U1758 (N_1758,N_1296,N_1205);
nor U1759 (N_1759,N_1294,N_1470);
and U1760 (N_1760,N_1264,N_1496);
nor U1761 (N_1761,N_1135,N_1184);
or U1762 (N_1762,N_1184,N_1405);
or U1763 (N_1763,N_1380,N_1134);
nor U1764 (N_1764,N_1113,N_1489);
and U1765 (N_1765,N_1199,N_1035);
nor U1766 (N_1766,N_1302,N_1295);
and U1767 (N_1767,N_1028,N_1265);
nand U1768 (N_1768,N_1442,N_1103);
or U1769 (N_1769,N_1220,N_1335);
or U1770 (N_1770,N_1317,N_1291);
or U1771 (N_1771,N_1012,N_1300);
nand U1772 (N_1772,N_1073,N_1301);
nor U1773 (N_1773,N_1183,N_1073);
and U1774 (N_1774,N_1376,N_1497);
nor U1775 (N_1775,N_1144,N_1461);
nand U1776 (N_1776,N_1352,N_1010);
nor U1777 (N_1777,N_1470,N_1392);
nor U1778 (N_1778,N_1485,N_1120);
nand U1779 (N_1779,N_1352,N_1218);
nand U1780 (N_1780,N_1419,N_1073);
or U1781 (N_1781,N_1232,N_1235);
or U1782 (N_1782,N_1382,N_1275);
or U1783 (N_1783,N_1089,N_1250);
or U1784 (N_1784,N_1101,N_1157);
nor U1785 (N_1785,N_1130,N_1368);
nand U1786 (N_1786,N_1299,N_1163);
nor U1787 (N_1787,N_1321,N_1465);
nor U1788 (N_1788,N_1332,N_1253);
or U1789 (N_1789,N_1291,N_1352);
or U1790 (N_1790,N_1077,N_1233);
nand U1791 (N_1791,N_1119,N_1310);
or U1792 (N_1792,N_1096,N_1188);
or U1793 (N_1793,N_1364,N_1421);
nor U1794 (N_1794,N_1296,N_1218);
and U1795 (N_1795,N_1380,N_1093);
and U1796 (N_1796,N_1055,N_1496);
nand U1797 (N_1797,N_1004,N_1222);
nor U1798 (N_1798,N_1075,N_1145);
nor U1799 (N_1799,N_1477,N_1358);
nand U1800 (N_1800,N_1380,N_1074);
nor U1801 (N_1801,N_1414,N_1269);
or U1802 (N_1802,N_1491,N_1050);
nand U1803 (N_1803,N_1072,N_1034);
and U1804 (N_1804,N_1114,N_1275);
or U1805 (N_1805,N_1178,N_1172);
nor U1806 (N_1806,N_1159,N_1237);
or U1807 (N_1807,N_1383,N_1351);
nor U1808 (N_1808,N_1118,N_1201);
nand U1809 (N_1809,N_1119,N_1262);
and U1810 (N_1810,N_1062,N_1401);
and U1811 (N_1811,N_1021,N_1028);
xor U1812 (N_1812,N_1462,N_1398);
nor U1813 (N_1813,N_1307,N_1071);
and U1814 (N_1814,N_1174,N_1185);
and U1815 (N_1815,N_1290,N_1329);
nand U1816 (N_1816,N_1102,N_1038);
nand U1817 (N_1817,N_1488,N_1270);
nand U1818 (N_1818,N_1382,N_1057);
nand U1819 (N_1819,N_1072,N_1478);
nand U1820 (N_1820,N_1426,N_1177);
nand U1821 (N_1821,N_1201,N_1293);
nand U1822 (N_1822,N_1443,N_1445);
nand U1823 (N_1823,N_1015,N_1404);
nor U1824 (N_1824,N_1022,N_1471);
nor U1825 (N_1825,N_1240,N_1185);
or U1826 (N_1826,N_1296,N_1190);
nor U1827 (N_1827,N_1266,N_1317);
nand U1828 (N_1828,N_1005,N_1085);
nand U1829 (N_1829,N_1114,N_1211);
and U1830 (N_1830,N_1490,N_1020);
and U1831 (N_1831,N_1436,N_1265);
nand U1832 (N_1832,N_1442,N_1067);
or U1833 (N_1833,N_1334,N_1017);
and U1834 (N_1834,N_1221,N_1253);
and U1835 (N_1835,N_1056,N_1237);
nand U1836 (N_1836,N_1165,N_1010);
and U1837 (N_1837,N_1168,N_1103);
nor U1838 (N_1838,N_1412,N_1478);
nand U1839 (N_1839,N_1236,N_1332);
or U1840 (N_1840,N_1143,N_1339);
nor U1841 (N_1841,N_1158,N_1367);
nor U1842 (N_1842,N_1103,N_1087);
nor U1843 (N_1843,N_1452,N_1050);
nand U1844 (N_1844,N_1116,N_1382);
nand U1845 (N_1845,N_1055,N_1088);
nand U1846 (N_1846,N_1057,N_1128);
nand U1847 (N_1847,N_1457,N_1348);
and U1848 (N_1848,N_1459,N_1100);
and U1849 (N_1849,N_1486,N_1144);
nand U1850 (N_1850,N_1065,N_1317);
nor U1851 (N_1851,N_1020,N_1192);
nand U1852 (N_1852,N_1306,N_1380);
or U1853 (N_1853,N_1481,N_1254);
nand U1854 (N_1854,N_1474,N_1087);
xor U1855 (N_1855,N_1377,N_1068);
or U1856 (N_1856,N_1384,N_1278);
nand U1857 (N_1857,N_1471,N_1153);
nor U1858 (N_1858,N_1329,N_1101);
and U1859 (N_1859,N_1434,N_1373);
and U1860 (N_1860,N_1494,N_1139);
or U1861 (N_1861,N_1338,N_1044);
nor U1862 (N_1862,N_1184,N_1092);
nand U1863 (N_1863,N_1177,N_1494);
nor U1864 (N_1864,N_1281,N_1059);
and U1865 (N_1865,N_1439,N_1128);
or U1866 (N_1866,N_1049,N_1083);
xnor U1867 (N_1867,N_1186,N_1313);
nor U1868 (N_1868,N_1037,N_1005);
nor U1869 (N_1869,N_1274,N_1459);
and U1870 (N_1870,N_1346,N_1101);
nor U1871 (N_1871,N_1466,N_1355);
nand U1872 (N_1872,N_1367,N_1332);
nand U1873 (N_1873,N_1478,N_1311);
and U1874 (N_1874,N_1266,N_1320);
and U1875 (N_1875,N_1474,N_1157);
nand U1876 (N_1876,N_1135,N_1070);
nand U1877 (N_1877,N_1000,N_1233);
nor U1878 (N_1878,N_1302,N_1176);
and U1879 (N_1879,N_1080,N_1342);
nand U1880 (N_1880,N_1056,N_1343);
nand U1881 (N_1881,N_1201,N_1448);
and U1882 (N_1882,N_1431,N_1120);
or U1883 (N_1883,N_1189,N_1353);
or U1884 (N_1884,N_1027,N_1366);
nor U1885 (N_1885,N_1488,N_1284);
and U1886 (N_1886,N_1478,N_1402);
nor U1887 (N_1887,N_1195,N_1258);
and U1888 (N_1888,N_1430,N_1402);
nand U1889 (N_1889,N_1421,N_1132);
nand U1890 (N_1890,N_1008,N_1246);
nand U1891 (N_1891,N_1006,N_1458);
or U1892 (N_1892,N_1417,N_1395);
nor U1893 (N_1893,N_1164,N_1271);
and U1894 (N_1894,N_1383,N_1238);
or U1895 (N_1895,N_1211,N_1448);
nand U1896 (N_1896,N_1292,N_1338);
nand U1897 (N_1897,N_1193,N_1135);
and U1898 (N_1898,N_1304,N_1200);
nand U1899 (N_1899,N_1451,N_1457);
nand U1900 (N_1900,N_1248,N_1428);
nor U1901 (N_1901,N_1416,N_1182);
nand U1902 (N_1902,N_1330,N_1429);
or U1903 (N_1903,N_1195,N_1062);
nand U1904 (N_1904,N_1291,N_1470);
nor U1905 (N_1905,N_1158,N_1161);
and U1906 (N_1906,N_1081,N_1114);
nand U1907 (N_1907,N_1306,N_1163);
and U1908 (N_1908,N_1111,N_1480);
or U1909 (N_1909,N_1052,N_1212);
and U1910 (N_1910,N_1344,N_1066);
nor U1911 (N_1911,N_1297,N_1005);
nand U1912 (N_1912,N_1453,N_1164);
nand U1913 (N_1913,N_1165,N_1298);
nand U1914 (N_1914,N_1330,N_1102);
nor U1915 (N_1915,N_1053,N_1172);
nand U1916 (N_1916,N_1217,N_1419);
and U1917 (N_1917,N_1112,N_1393);
or U1918 (N_1918,N_1439,N_1249);
nor U1919 (N_1919,N_1365,N_1059);
nor U1920 (N_1920,N_1098,N_1011);
or U1921 (N_1921,N_1324,N_1234);
and U1922 (N_1922,N_1369,N_1226);
nor U1923 (N_1923,N_1255,N_1242);
or U1924 (N_1924,N_1395,N_1232);
nor U1925 (N_1925,N_1023,N_1102);
and U1926 (N_1926,N_1293,N_1137);
or U1927 (N_1927,N_1170,N_1002);
nand U1928 (N_1928,N_1283,N_1039);
nand U1929 (N_1929,N_1127,N_1155);
nor U1930 (N_1930,N_1219,N_1100);
and U1931 (N_1931,N_1077,N_1482);
or U1932 (N_1932,N_1130,N_1003);
and U1933 (N_1933,N_1321,N_1053);
nand U1934 (N_1934,N_1481,N_1388);
or U1935 (N_1935,N_1299,N_1108);
nand U1936 (N_1936,N_1231,N_1438);
and U1937 (N_1937,N_1356,N_1171);
or U1938 (N_1938,N_1482,N_1479);
or U1939 (N_1939,N_1022,N_1008);
nand U1940 (N_1940,N_1005,N_1281);
nand U1941 (N_1941,N_1107,N_1480);
nor U1942 (N_1942,N_1491,N_1446);
and U1943 (N_1943,N_1033,N_1078);
nor U1944 (N_1944,N_1120,N_1177);
nand U1945 (N_1945,N_1216,N_1205);
nor U1946 (N_1946,N_1123,N_1083);
or U1947 (N_1947,N_1110,N_1424);
nand U1948 (N_1948,N_1220,N_1239);
and U1949 (N_1949,N_1350,N_1089);
or U1950 (N_1950,N_1354,N_1295);
and U1951 (N_1951,N_1160,N_1112);
and U1952 (N_1952,N_1420,N_1256);
or U1953 (N_1953,N_1469,N_1140);
or U1954 (N_1954,N_1451,N_1189);
nand U1955 (N_1955,N_1121,N_1186);
and U1956 (N_1956,N_1305,N_1372);
or U1957 (N_1957,N_1420,N_1238);
or U1958 (N_1958,N_1228,N_1328);
and U1959 (N_1959,N_1052,N_1193);
or U1960 (N_1960,N_1201,N_1457);
nor U1961 (N_1961,N_1385,N_1323);
and U1962 (N_1962,N_1413,N_1202);
nor U1963 (N_1963,N_1005,N_1305);
and U1964 (N_1964,N_1009,N_1374);
nor U1965 (N_1965,N_1216,N_1156);
or U1966 (N_1966,N_1467,N_1287);
nor U1967 (N_1967,N_1305,N_1176);
nand U1968 (N_1968,N_1149,N_1475);
nor U1969 (N_1969,N_1454,N_1469);
nand U1970 (N_1970,N_1171,N_1007);
and U1971 (N_1971,N_1190,N_1220);
nor U1972 (N_1972,N_1050,N_1004);
nand U1973 (N_1973,N_1063,N_1327);
xnor U1974 (N_1974,N_1456,N_1139);
or U1975 (N_1975,N_1204,N_1105);
nand U1976 (N_1976,N_1444,N_1482);
nor U1977 (N_1977,N_1262,N_1276);
nand U1978 (N_1978,N_1046,N_1177);
and U1979 (N_1979,N_1068,N_1381);
and U1980 (N_1980,N_1081,N_1086);
and U1981 (N_1981,N_1259,N_1270);
and U1982 (N_1982,N_1168,N_1151);
or U1983 (N_1983,N_1383,N_1337);
and U1984 (N_1984,N_1433,N_1403);
nor U1985 (N_1985,N_1106,N_1080);
nor U1986 (N_1986,N_1219,N_1382);
nor U1987 (N_1987,N_1164,N_1071);
and U1988 (N_1988,N_1021,N_1367);
or U1989 (N_1989,N_1411,N_1366);
or U1990 (N_1990,N_1435,N_1462);
nor U1991 (N_1991,N_1066,N_1463);
and U1992 (N_1992,N_1495,N_1265);
nand U1993 (N_1993,N_1227,N_1485);
and U1994 (N_1994,N_1389,N_1328);
and U1995 (N_1995,N_1092,N_1040);
nor U1996 (N_1996,N_1217,N_1463);
nand U1997 (N_1997,N_1478,N_1474);
or U1998 (N_1998,N_1037,N_1326);
or U1999 (N_1999,N_1114,N_1360);
and U2000 (N_2000,N_1501,N_1688);
nand U2001 (N_2001,N_1809,N_1507);
and U2002 (N_2002,N_1813,N_1830);
or U2003 (N_2003,N_1767,N_1974);
or U2004 (N_2004,N_1758,N_1981);
or U2005 (N_2005,N_1804,N_1722);
nor U2006 (N_2006,N_1972,N_1627);
nand U2007 (N_2007,N_1651,N_1669);
or U2008 (N_2008,N_1951,N_1628);
and U2009 (N_2009,N_1694,N_1984);
nand U2010 (N_2010,N_1662,N_1761);
or U2011 (N_2011,N_1668,N_1573);
or U2012 (N_2012,N_1900,N_1744);
xor U2013 (N_2013,N_1901,N_1533);
nand U2014 (N_2014,N_1535,N_1559);
or U2015 (N_2015,N_1759,N_1942);
or U2016 (N_2016,N_1864,N_1913);
and U2017 (N_2017,N_1964,N_1608);
nor U2018 (N_2018,N_1868,N_1824);
nor U2019 (N_2019,N_1701,N_1750);
and U2020 (N_2020,N_1873,N_1992);
and U2021 (N_2021,N_1703,N_1998);
or U2022 (N_2022,N_1505,N_1816);
or U2023 (N_2023,N_1966,N_1756);
or U2024 (N_2024,N_1817,N_1725);
nor U2025 (N_2025,N_1677,N_1819);
and U2026 (N_2026,N_1866,N_1939);
xor U2027 (N_2027,N_1692,N_1825);
nand U2028 (N_2028,N_1990,N_1956);
nand U2029 (N_2029,N_1684,N_1869);
and U2030 (N_2030,N_1745,N_1516);
nor U2031 (N_2031,N_1615,N_1691);
nand U2032 (N_2032,N_1739,N_1567);
or U2033 (N_2033,N_1920,N_1892);
nor U2034 (N_2034,N_1777,N_1571);
nand U2035 (N_2035,N_1714,N_1988);
nor U2036 (N_2036,N_1967,N_1637);
nor U2037 (N_2037,N_1704,N_1860);
and U2038 (N_2038,N_1896,N_1619);
nor U2039 (N_2039,N_1757,N_1959);
or U2040 (N_2040,N_1524,N_1909);
and U2041 (N_2041,N_1854,N_1898);
nor U2042 (N_2042,N_1975,N_1616);
nor U2043 (N_2043,N_1924,N_1595);
and U2044 (N_2044,N_1560,N_1877);
nor U2045 (N_2045,N_1729,N_1514);
or U2046 (N_2046,N_1926,N_1686);
nand U2047 (N_2047,N_1857,N_1855);
nor U2048 (N_2048,N_1636,N_1609);
or U2049 (N_2049,N_1927,N_1800);
and U2050 (N_2050,N_1790,N_1952);
or U2051 (N_2051,N_1706,N_1755);
and U2052 (N_2052,N_1922,N_1598);
nor U2053 (N_2053,N_1837,N_1808);
nand U2054 (N_2054,N_1687,N_1544);
nor U2055 (N_2055,N_1566,N_1579);
or U2056 (N_2056,N_1787,N_1995);
or U2057 (N_2057,N_1944,N_1648);
and U2058 (N_2058,N_1614,N_1957);
or U2059 (N_2059,N_1679,N_1580);
or U2060 (N_2060,N_1699,N_1563);
or U2061 (N_2061,N_1806,N_1530);
or U2062 (N_2062,N_1764,N_1589);
and U2063 (N_2063,N_1862,N_1564);
nor U2064 (N_2064,N_1638,N_1958);
nor U2065 (N_2065,N_1879,N_1941);
nor U2066 (N_2066,N_1548,N_1517);
nor U2067 (N_2067,N_1602,N_1712);
and U2068 (N_2068,N_1891,N_1557);
or U2069 (N_2069,N_1680,N_1789);
nand U2070 (N_2070,N_1858,N_1778);
and U2071 (N_2071,N_1751,N_1834);
or U2072 (N_2072,N_1805,N_1907);
nor U2073 (N_2073,N_1618,N_1730);
and U2074 (N_2074,N_1653,N_1949);
nand U2075 (N_2075,N_1885,N_1803);
or U2076 (N_2076,N_1818,N_1705);
nand U2077 (N_2077,N_1523,N_1591);
nand U2078 (N_2078,N_1979,N_1675);
or U2079 (N_2079,N_1953,N_1856);
nand U2080 (N_2080,N_1810,N_1536);
and U2081 (N_2081,N_1748,N_1781);
and U2082 (N_2082,N_1645,N_1776);
or U2083 (N_2083,N_1508,N_1693);
or U2084 (N_2084,N_1768,N_1503);
or U2085 (N_2085,N_1689,N_1644);
nand U2086 (N_2086,N_1683,N_1925);
or U2087 (N_2087,N_1801,N_1793);
or U2088 (N_2088,N_1574,N_1812);
nand U2089 (N_2089,N_1547,N_1795);
or U2090 (N_2090,N_1720,N_1664);
nor U2091 (N_2091,N_1785,N_1918);
and U2092 (N_2092,N_1632,N_1921);
or U2093 (N_2093,N_1641,N_1954);
or U2094 (N_2094,N_1534,N_1696);
and U2095 (N_2095,N_1655,N_1791);
or U2096 (N_2096,N_1500,N_1843);
nand U2097 (N_2097,N_1786,N_1635);
nor U2098 (N_2098,N_1707,N_1577);
nand U2099 (N_2099,N_1605,N_1999);
nand U2100 (N_2100,N_1780,N_1875);
nand U2101 (N_2101,N_1646,N_1831);
nor U2102 (N_2102,N_1702,N_1889);
or U2103 (N_2103,N_1697,N_1634);
nor U2104 (N_2104,N_1977,N_1665);
nand U2105 (N_2105,N_1586,N_1842);
nand U2106 (N_2106,N_1610,N_1626);
and U2107 (N_2107,N_1642,N_1948);
and U2108 (N_2108,N_1597,N_1839);
or U2109 (N_2109,N_1711,N_1894);
and U2110 (N_2110,N_1844,N_1727);
nor U2111 (N_2111,N_1512,N_1732);
and U2112 (N_2112,N_1775,N_1719);
nand U2113 (N_2113,N_1742,N_1823);
nor U2114 (N_2114,N_1519,N_1763);
or U2115 (N_2115,N_1596,N_1731);
or U2116 (N_2116,N_1960,N_1915);
nor U2117 (N_2117,N_1562,N_1674);
nor U2118 (N_2118,N_1695,N_1936);
nor U2119 (N_2119,N_1603,N_1565);
and U2120 (N_2120,N_1661,N_1685);
nand U2121 (N_2121,N_1623,N_1724);
or U2122 (N_2122,N_1518,N_1876);
nand U2123 (N_2123,N_1903,N_1982);
nand U2124 (N_2124,N_1989,N_1550);
nand U2125 (N_2125,N_1652,N_1887);
or U2126 (N_2126,N_1600,N_1584);
or U2127 (N_2127,N_1511,N_1983);
and U2128 (N_2128,N_1772,N_1766);
or U2129 (N_2129,N_1765,N_1513);
nor U2130 (N_2130,N_1723,N_1576);
and U2131 (N_2131,N_1993,N_1746);
nor U2132 (N_2132,N_1538,N_1607);
and U2133 (N_2133,N_1760,N_1715);
and U2134 (N_2134,N_1553,N_1752);
nand U2135 (N_2135,N_1708,N_1713);
and U2136 (N_2136,N_1561,N_1946);
and U2137 (N_2137,N_1933,N_1542);
or U2138 (N_2138,N_1911,N_1672);
or U2139 (N_2139,N_1671,N_1852);
or U2140 (N_2140,N_1601,N_1572);
or U2141 (N_2141,N_1643,N_1734);
nand U2142 (N_2142,N_1845,N_1867);
and U2143 (N_2143,N_1718,N_1840);
and U2144 (N_2144,N_1794,N_1882);
and U2145 (N_2145,N_1888,N_1740);
nor U2146 (N_2146,N_1802,N_1822);
and U2147 (N_2147,N_1916,N_1502);
nor U2148 (N_2148,N_1541,N_1861);
and U2149 (N_2149,N_1509,N_1784);
or U2150 (N_2150,N_1878,N_1811);
and U2151 (N_2151,N_1821,N_1893);
and U2152 (N_2152,N_1910,N_1994);
nor U2153 (N_2153,N_1543,N_1950);
or U2154 (N_2154,N_1594,N_1585);
or U2155 (N_2155,N_1678,N_1826);
nor U2156 (N_2156,N_1897,N_1884);
nor U2157 (N_2157,N_1558,N_1996);
nor U2158 (N_2158,N_1851,N_1621);
nor U2159 (N_2159,N_1531,N_1880);
nor U2160 (N_2160,N_1955,N_1629);
nand U2161 (N_2161,N_1575,N_1710);
nor U2162 (N_2162,N_1779,N_1552);
nor U2163 (N_2163,N_1522,N_1792);
and U2164 (N_2164,N_1770,N_1836);
and U2165 (N_2165,N_1895,N_1622);
nor U2166 (N_2166,N_1647,N_1798);
nor U2167 (N_2167,N_1700,N_1871);
or U2168 (N_2168,N_1617,N_1846);
or U2169 (N_2169,N_1991,N_1886);
or U2170 (N_2170,N_1947,N_1904);
and U2171 (N_2171,N_1578,N_1797);
nand U2172 (N_2172,N_1735,N_1630);
nor U2173 (N_2173,N_1961,N_1506);
nand U2174 (N_2174,N_1666,N_1539);
nor U2175 (N_2175,N_1935,N_1733);
or U2176 (N_2176,N_1737,N_1849);
nand U2177 (N_2177,N_1673,N_1592);
or U2178 (N_2178,N_1520,N_1970);
nand U2179 (N_2179,N_1774,N_1504);
and U2180 (N_2180,N_1848,N_1537);
nand U2181 (N_2181,N_1938,N_1555);
or U2182 (N_2182,N_1660,N_1976);
nor U2183 (N_2183,N_1649,N_1963);
and U2184 (N_2184,N_1593,N_1783);
and U2185 (N_2185,N_1741,N_1659);
nor U2186 (N_2186,N_1569,N_1968);
and U2187 (N_2187,N_1676,N_1625);
or U2188 (N_2188,N_1604,N_1997);
nor U2189 (N_2189,N_1870,N_1527);
or U2190 (N_2190,N_1650,N_1510);
nor U2191 (N_2191,N_1859,N_1639);
and U2192 (N_2192,N_1515,N_1670);
and U2193 (N_2193,N_1987,N_1754);
nand U2194 (N_2194,N_1624,N_1929);
or U2195 (N_2195,N_1850,N_1820);
and U2196 (N_2196,N_1890,N_1881);
and U2197 (N_2197,N_1698,N_1853);
nor U2198 (N_2198,N_1528,N_1769);
nand U2199 (N_2199,N_1716,N_1654);
nor U2200 (N_2200,N_1841,N_1726);
and U2201 (N_2201,N_1788,N_1545);
or U2202 (N_2202,N_1633,N_1606);
nand U2203 (N_2203,N_1923,N_1681);
and U2204 (N_2204,N_1908,N_1932);
nor U2205 (N_2205,N_1832,N_1930);
nand U2206 (N_2206,N_1863,N_1613);
or U2207 (N_2207,N_1581,N_1717);
and U2208 (N_2208,N_1838,N_1728);
nand U2209 (N_2209,N_1874,N_1658);
nor U2210 (N_2210,N_1978,N_1599);
nand U2211 (N_2211,N_1928,N_1835);
nor U2212 (N_2212,N_1872,N_1914);
and U2213 (N_2213,N_1943,N_1883);
or U2214 (N_2214,N_1753,N_1521);
nand U2215 (N_2215,N_1847,N_1546);
or U2216 (N_2216,N_1556,N_1771);
nor U2217 (N_2217,N_1934,N_1568);
nor U2218 (N_2218,N_1940,N_1899);
and U2219 (N_2219,N_1833,N_1931);
and U2220 (N_2220,N_1551,N_1554);
and U2221 (N_2221,N_1640,N_1986);
or U2222 (N_2222,N_1905,N_1762);
nor U2223 (N_2223,N_1540,N_1865);
or U2224 (N_2224,N_1663,N_1969);
and U2225 (N_2225,N_1980,N_1782);
nand U2226 (N_2226,N_1814,N_1973);
or U2227 (N_2227,N_1612,N_1749);
nor U2228 (N_2228,N_1631,N_1709);
or U2229 (N_2229,N_1587,N_1799);
nand U2230 (N_2230,N_1912,N_1917);
nand U2231 (N_2231,N_1965,N_1529);
nand U2232 (N_2232,N_1583,N_1588);
xor U2233 (N_2233,N_1682,N_1937);
and U2234 (N_2234,N_1828,N_1743);
and U2235 (N_2235,N_1829,N_1919);
or U2236 (N_2236,N_1815,N_1590);
nor U2237 (N_2237,N_1902,N_1985);
or U2238 (N_2238,N_1945,N_1525);
and U2239 (N_2239,N_1736,N_1657);
nand U2240 (N_2240,N_1667,N_1532);
nor U2241 (N_2241,N_1620,N_1962);
nor U2242 (N_2242,N_1738,N_1971);
nand U2243 (N_2243,N_1773,N_1526);
or U2244 (N_2244,N_1747,N_1549);
and U2245 (N_2245,N_1827,N_1906);
nor U2246 (N_2246,N_1656,N_1611);
or U2247 (N_2247,N_1807,N_1570);
nand U2248 (N_2248,N_1796,N_1721);
nand U2249 (N_2249,N_1690,N_1582);
nor U2250 (N_2250,N_1521,N_1717);
or U2251 (N_2251,N_1998,N_1944);
and U2252 (N_2252,N_1879,N_1947);
nor U2253 (N_2253,N_1506,N_1904);
or U2254 (N_2254,N_1963,N_1519);
or U2255 (N_2255,N_1852,N_1614);
and U2256 (N_2256,N_1936,N_1583);
or U2257 (N_2257,N_1878,N_1698);
and U2258 (N_2258,N_1618,N_1674);
or U2259 (N_2259,N_1685,N_1652);
and U2260 (N_2260,N_1924,N_1965);
or U2261 (N_2261,N_1504,N_1827);
or U2262 (N_2262,N_1712,N_1865);
nand U2263 (N_2263,N_1736,N_1952);
or U2264 (N_2264,N_1529,N_1897);
and U2265 (N_2265,N_1556,N_1842);
nor U2266 (N_2266,N_1740,N_1561);
nor U2267 (N_2267,N_1898,N_1779);
or U2268 (N_2268,N_1753,N_1944);
or U2269 (N_2269,N_1904,N_1976);
nand U2270 (N_2270,N_1843,N_1817);
or U2271 (N_2271,N_1739,N_1949);
or U2272 (N_2272,N_1642,N_1741);
and U2273 (N_2273,N_1999,N_1627);
nand U2274 (N_2274,N_1977,N_1826);
or U2275 (N_2275,N_1578,N_1945);
or U2276 (N_2276,N_1726,N_1886);
or U2277 (N_2277,N_1722,N_1753);
nor U2278 (N_2278,N_1679,N_1802);
nor U2279 (N_2279,N_1920,N_1953);
and U2280 (N_2280,N_1723,N_1685);
and U2281 (N_2281,N_1649,N_1951);
or U2282 (N_2282,N_1932,N_1584);
nor U2283 (N_2283,N_1637,N_1602);
nand U2284 (N_2284,N_1526,N_1965);
or U2285 (N_2285,N_1547,N_1989);
nand U2286 (N_2286,N_1509,N_1807);
or U2287 (N_2287,N_1565,N_1686);
or U2288 (N_2288,N_1648,N_1589);
nand U2289 (N_2289,N_1604,N_1684);
nand U2290 (N_2290,N_1633,N_1729);
or U2291 (N_2291,N_1708,N_1998);
nand U2292 (N_2292,N_1910,N_1572);
or U2293 (N_2293,N_1829,N_1718);
nand U2294 (N_2294,N_1818,N_1567);
nor U2295 (N_2295,N_1869,N_1924);
or U2296 (N_2296,N_1685,N_1837);
nand U2297 (N_2297,N_1932,N_1655);
nand U2298 (N_2298,N_1502,N_1510);
nand U2299 (N_2299,N_1730,N_1595);
nor U2300 (N_2300,N_1839,N_1890);
nor U2301 (N_2301,N_1889,N_1888);
and U2302 (N_2302,N_1948,N_1774);
nor U2303 (N_2303,N_1594,N_1746);
and U2304 (N_2304,N_1741,N_1513);
and U2305 (N_2305,N_1722,N_1960);
or U2306 (N_2306,N_1626,N_1756);
and U2307 (N_2307,N_1856,N_1693);
and U2308 (N_2308,N_1981,N_1957);
and U2309 (N_2309,N_1730,N_1949);
or U2310 (N_2310,N_1607,N_1853);
and U2311 (N_2311,N_1910,N_1969);
nand U2312 (N_2312,N_1690,N_1506);
and U2313 (N_2313,N_1592,N_1581);
or U2314 (N_2314,N_1665,N_1917);
and U2315 (N_2315,N_1922,N_1901);
or U2316 (N_2316,N_1616,N_1802);
nor U2317 (N_2317,N_1743,N_1554);
or U2318 (N_2318,N_1690,N_1605);
and U2319 (N_2319,N_1779,N_1589);
nand U2320 (N_2320,N_1553,N_1744);
or U2321 (N_2321,N_1871,N_1756);
and U2322 (N_2322,N_1947,N_1624);
or U2323 (N_2323,N_1870,N_1658);
and U2324 (N_2324,N_1508,N_1710);
nor U2325 (N_2325,N_1810,N_1575);
nor U2326 (N_2326,N_1834,N_1894);
nor U2327 (N_2327,N_1830,N_1987);
nand U2328 (N_2328,N_1809,N_1833);
nand U2329 (N_2329,N_1501,N_1710);
and U2330 (N_2330,N_1513,N_1898);
or U2331 (N_2331,N_1752,N_1986);
and U2332 (N_2332,N_1956,N_1730);
nor U2333 (N_2333,N_1802,N_1749);
nor U2334 (N_2334,N_1671,N_1805);
and U2335 (N_2335,N_1843,N_1688);
nor U2336 (N_2336,N_1650,N_1935);
nor U2337 (N_2337,N_1524,N_1685);
or U2338 (N_2338,N_1534,N_1749);
nor U2339 (N_2339,N_1709,N_1828);
nor U2340 (N_2340,N_1507,N_1859);
or U2341 (N_2341,N_1548,N_1988);
nor U2342 (N_2342,N_1711,N_1989);
nor U2343 (N_2343,N_1605,N_1570);
or U2344 (N_2344,N_1509,N_1583);
nor U2345 (N_2345,N_1501,N_1615);
nand U2346 (N_2346,N_1687,N_1525);
nand U2347 (N_2347,N_1823,N_1749);
and U2348 (N_2348,N_1981,N_1953);
and U2349 (N_2349,N_1682,N_1702);
and U2350 (N_2350,N_1570,N_1712);
nand U2351 (N_2351,N_1858,N_1918);
or U2352 (N_2352,N_1855,N_1726);
and U2353 (N_2353,N_1871,N_1714);
and U2354 (N_2354,N_1628,N_1939);
and U2355 (N_2355,N_1685,N_1912);
and U2356 (N_2356,N_1756,N_1613);
or U2357 (N_2357,N_1949,N_1688);
nand U2358 (N_2358,N_1839,N_1537);
nor U2359 (N_2359,N_1696,N_1799);
nor U2360 (N_2360,N_1669,N_1890);
and U2361 (N_2361,N_1843,N_1700);
and U2362 (N_2362,N_1749,N_1766);
and U2363 (N_2363,N_1883,N_1523);
nand U2364 (N_2364,N_1573,N_1936);
nand U2365 (N_2365,N_1931,N_1641);
nand U2366 (N_2366,N_1573,N_1740);
nand U2367 (N_2367,N_1995,N_1500);
nand U2368 (N_2368,N_1677,N_1543);
nand U2369 (N_2369,N_1826,N_1604);
or U2370 (N_2370,N_1665,N_1806);
nand U2371 (N_2371,N_1944,N_1623);
nand U2372 (N_2372,N_1958,N_1721);
and U2373 (N_2373,N_1645,N_1727);
nor U2374 (N_2374,N_1539,N_1651);
and U2375 (N_2375,N_1924,N_1758);
or U2376 (N_2376,N_1829,N_1688);
or U2377 (N_2377,N_1690,N_1999);
nor U2378 (N_2378,N_1607,N_1521);
nand U2379 (N_2379,N_1572,N_1936);
and U2380 (N_2380,N_1640,N_1670);
and U2381 (N_2381,N_1745,N_1732);
nor U2382 (N_2382,N_1993,N_1910);
nor U2383 (N_2383,N_1906,N_1931);
nor U2384 (N_2384,N_1912,N_1592);
nand U2385 (N_2385,N_1749,N_1714);
or U2386 (N_2386,N_1994,N_1769);
and U2387 (N_2387,N_1715,N_1652);
or U2388 (N_2388,N_1665,N_1877);
nand U2389 (N_2389,N_1879,N_1902);
and U2390 (N_2390,N_1960,N_1919);
or U2391 (N_2391,N_1983,N_1564);
and U2392 (N_2392,N_1519,N_1528);
or U2393 (N_2393,N_1844,N_1951);
nor U2394 (N_2394,N_1787,N_1508);
and U2395 (N_2395,N_1815,N_1783);
nor U2396 (N_2396,N_1945,N_1826);
nor U2397 (N_2397,N_1552,N_1725);
or U2398 (N_2398,N_1649,N_1936);
or U2399 (N_2399,N_1608,N_1806);
or U2400 (N_2400,N_1588,N_1512);
or U2401 (N_2401,N_1623,N_1620);
and U2402 (N_2402,N_1666,N_1993);
nor U2403 (N_2403,N_1872,N_1907);
and U2404 (N_2404,N_1707,N_1832);
and U2405 (N_2405,N_1836,N_1708);
nor U2406 (N_2406,N_1696,N_1819);
and U2407 (N_2407,N_1695,N_1719);
nand U2408 (N_2408,N_1566,N_1898);
or U2409 (N_2409,N_1579,N_1655);
nor U2410 (N_2410,N_1982,N_1977);
and U2411 (N_2411,N_1851,N_1871);
and U2412 (N_2412,N_1578,N_1633);
xnor U2413 (N_2413,N_1845,N_1629);
nor U2414 (N_2414,N_1769,N_1718);
nor U2415 (N_2415,N_1621,N_1756);
or U2416 (N_2416,N_1794,N_1798);
and U2417 (N_2417,N_1550,N_1764);
nor U2418 (N_2418,N_1720,N_1976);
nand U2419 (N_2419,N_1603,N_1932);
nand U2420 (N_2420,N_1564,N_1964);
and U2421 (N_2421,N_1895,N_1620);
xor U2422 (N_2422,N_1895,N_1723);
or U2423 (N_2423,N_1974,N_1798);
nor U2424 (N_2424,N_1911,N_1866);
or U2425 (N_2425,N_1920,N_1527);
or U2426 (N_2426,N_1531,N_1937);
and U2427 (N_2427,N_1969,N_1988);
nor U2428 (N_2428,N_1627,N_1807);
or U2429 (N_2429,N_1891,N_1665);
nor U2430 (N_2430,N_1914,N_1610);
nand U2431 (N_2431,N_1798,N_1770);
or U2432 (N_2432,N_1663,N_1709);
and U2433 (N_2433,N_1543,N_1949);
and U2434 (N_2434,N_1777,N_1832);
or U2435 (N_2435,N_1942,N_1845);
xnor U2436 (N_2436,N_1604,N_1967);
nor U2437 (N_2437,N_1560,N_1643);
and U2438 (N_2438,N_1890,N_1767);
nand U2439 (N_2439,N_1736,N_1821);
nand U2440 (N_2440,N_1966,N_1512);
nand U2441 (N_2441,N_1908,N_1582);
nor U2442 (N_2442,N_1636,N_1895);
or U2443 (N_2443,N_1993,N_1924);
nor U2444 (N_2444,N_1971,N_1525);
nand U2445 (N_2445,N_1750,N_1649);
or U2446 (N_2446,N_1815,N_1987);
and U2447 (N_2447,N_1557,N_1647);
or U2448 (N_2448,N_1649,N_1632);
or U2449 (N_2449,N_1570,N_1903);
and U2450 (N_2450,N_1749,N_1815);
nand U2451 (N_2451,N_1708,N_1826);
nor U2452 (N_2452,N_1691,N_1720);
or U2453 (N_2453,N_1729,N_1821);
nor U2454 (N_2454,N_1704,N_1515);
nand U2455 (N_2455,N_1679,N_1561);
or U2456 (N_2456,N_1688,N_1990);
nor U2457 (N_2457,N_1892,N_1842);
or U2458 (N_2458,N_1996,N_1898);
or U2459 (N_2459,N_1631,N_1507);
nand U2460 (N_2460,N_1852,N_1907);
or U2461 (N_2461,N_1886,N_1875);
or U2462 (N_2462,N_1639,N_1767);
nor U2463 (N_2463,N_1999,N_1581);
nor U2464 (N_2464,N_1686,N_1952);
and U2465 (N_2465,N_1936,N_1995);
nand U2466 (N_2466,N_1760,N_1772);
nand U2467 (N_2467,N_1837,N_1761);
and U2468 (N_2468,N_1540,N_1536);
nand U2469 (N_2469,N_1795,N_1572);
and U2470 (N_2470,N_1548,N_1899);
or U2471 (N_2471,N_1704,N_1764);
nand U2472 (N_2472,N_1689,N_1608);
nand U2473 (N_2473,N_1788,N_1668);
and U2474 (N_2474,N_1801,N_1938);
and U2475 (N_2475,N_1557,N_1752);
nand U2476 (N_2476,N_1765,N_1600);
or U2477 (N_2477,N_1845,N_1535);
and U2478 (N_2478,N_1977,N_1580);
nand U2479 (N_2479,N_1837,N_1642);
or U2480 (N_2480,N_1569,N_1749);
or U2481 (N_2481,N_1964,N_1775);
nand U2482 (N_2482,N_1756,N_1851);
and U2483 (N_2483,N_1859,N_1575);
and U2484 (N_2484,N_1945,N_1519);
and U2485 (N_2485,N_1677,N_1768);
or U2486 (N_2486,N_1949,N_1942);
nor U2487 (N_2487,N_1799,N_1651);
nand U2488 (N_2488,N_1859,N_1954);
nand U2489 (N_2489,N_1636,N_1922);
nor U2490 (N_2490,N_1918,N_1772);
or U2491 (N_2491,N_1913,N_1859);
nand U2492 (N_2492,N_1785,N_1731);
or U2493 (N_2493,N_1772,N_1916);
nor U2494 (N_2494,N_1685,N_1840);
nand U2495 (N_2495,N_1999,N_1733);
and U2496 (N_2496,N_1626,N_1545);
or U2497 (N_2497,N_1558,N_1572);
nor U2498 (N_2498,N_1898,N_1981);
or U2499 (N_2499,N_1909,N_1599);
nor U2500 (N_2500,N_2001,N_2188);
and U2501 (N_2501,N_2359,N_2080);
nand U2502 (N_2502,N_2217,N_2118);
nand U2503 (N_2503,N_2027,N_2132);
and U2504 (N_2504,N_2067,N_2427);
and U2505 (N_2505,N_2232,N_2452);
or U2506 (N_2506,N_2225,N_2270);
and U2507 (N_2507,N_2262,N_2363);
and U2508 (N_2508,N_2407,N_2162);
nand U2509 (N_2509,N_2249,N_2177);
nor U2510 (N_2510,N_2248,N_2304);
nor U2511 (N_2511,N_2441,N_2137);
nand U2512 (N_2512,N_2488,N_2199);
and U2513 (N_2513,N_2043,N_2054);
and U2514 (N_2514,N_2064,N_2330);
nand U2515 (N_2515,N_2050,N_2448);
nor U2516 (N_2516,N_2444,N_2034);
xnor U2517 (N_2517,N_2108,N_2372);
or U2518 (N_2518,N_2336,N_2158);
nor U2519 (N_2519,N_2065,N_2429);
nor U2520 (N_2520,N_2038,N_2149);
and U2521 (N_2521,N_2391,N_2288);
nor U2522 (N_2522,N_2128,N_2409);
nor U2523 (N_2523,N_2022,N_2004);
or U2524 (N_2524,N_2339,N_2364);
and U2525 (N_2525,N_2436,N_2115);
or U2526 (N_2526,N_2279,N_2224);
nand U2527 (N_2527,N_2009,N_2209);
and U2528 (N_2528,N_2099,N_2286);
and U2529 (N_2529,N_2333,N_2066);
nor U2530 (N_2530,N_2013,N_2063);
and U2531 (N_2531,N_2155,N_2349);
nor U2532 (N_2532,N_2335,N_2218);
nand U2533 (N_2533,N_2052,N_2216);
nor U2534 (N_2534,N_2134,N_2252);
or U2535 (N_2535,N_2474,N_2408);
nand U2536 (N_2536,N_2173,N_2097);
and U2537 (N_2537,N_2422,N_2076);
and U2538 (N_2538,N_2111,N_2200);
nor U2539 (N_2539,N_2397,N_2018);
nand U2540 (N_2540,N_2344,N_2451);
nand U2541 (N_2541,N_2124,N_2040);
or U2542 (N_2542,N_2074,N_2443);
nor U2543 (N_2543,N_2498,N_2142);
nand U2544 (N_2544,N_2306,N_2398);
or U2545 (N_2545,N_2459,N_2011);
nor U2546 (N_2546,N_2073,N_2401);
nor U2547 (N_2547,N_2166,N_2123);
and U2548 (N_2548,N_2144,N_2223);
and U2549 (N_2549,N_2490,N_2057);
nand U2550 (N_2550,N_2323,N_2376);
or U2551 (N_2551,N_2193,N_2412);
nor U2552 (N_2552,N_2228,N_2293);
or U2553 (N_2553,N_2187,N_2321);
nor U2554 (N_2554,N_2470,N_2240);
or U2555 (N_2555,N_2070,N_2127);
or U2556 (N_2556,N_2475,N_2319);
or U2557 (N_2557,N_2480,N_2437);
or U2558 (N_2558,N_2112,N_2312);
nor U2559 (N_2559,N_2213,N_2423);
and U2560 (N_2560,N_2077,N_2210);
nor U2561 (N_2561,N_2375,N_2109);
nor U2562 (N_2562,N_2150,N_2289);
nor U2563 (N_2563,N_2296,N_2340);
nand U2564 (N_2564,N_2211,N_2017);
xor U2565 (N_2565,N_2447,N_2492);
and U2566 (N_2566,N_2325,N_2455);
and U2567 (N_2567,N_2174,N_2131);
or U2568 (N_2568,N_2117,N_2085);
nand U2569 (N_2569,N_2389,N_2396);
or U2570 (N_2570,N_2386,N_2291);
nor U2571 (N_2571,N_2495,N_2160);
and U2572 (N_2572,N_2007,N_2461);
nor U2573 (N_2573,N_2192,N_2159);
nand U2574 (N_2574,N_2251,N_2136);
nand U2575 (N_2575,N_2230,N_2308);
nor U2576 (N_2576,N_2247,N_2298);
nand U2577 (N_2577,N_2404,N_2014);
and U2578 (N_2578,N_2190,N_2163);
or U2579 (N_2579,N_2345,N_2287);
nand U2580 (N_2580,N_2322,N_2318);
nand U2581 (N_2581,N_2047,N_2453);
nand U2582 (N_2582,N_2121,N_2028);
and U2583 (N_2583,N_2395,N_2140);
nand U2584 (N_2584,N_2183,N_2012);
nor U2585 (N_2585,N_2393,N_2305);
and U2586 (N_2586,N_2297,N_2171);
nand U2587 (N_2587,N_2487,N_2244);
or U2588 (N_2588,N_2433,N_2354);
and U2589 (N_2589,N_2428,N_2167);
nor U2590 (N_2590,N_2438,N_2479);
nor U2591 (N_2591,N_2403,N_2311);
and U2592 (N_2592,N_2129,N_2434);
nor U2593 (N_2593,N_2332,N_2069);
or U2594 (N_2594,N_2044,N_2464);
nand U2595 (N_2595,N_2274,N_2029);
or U2596 (N_2596,N_2058,N_2161);
or U2597 (N_2597,N_2237,N_2031);
or U2598 (N_2598,N_2267,N_2178);
or U2599 (N_2599,N_2374,N_2046);
or U2600 (N_2600,N_2116,N_2263);
nor U2601 (N_2601,N_2275,N_2035);
nor U2602 (N_2602,N_2493,N_2019);
nand U2603 (N_2603,N_2104,N_2169);
and U2604 (N_2604,N_2334,N_2320);
and U2605 (N_2605,N_2186,N_2039);
and U2606 (N_2606,N_2426,N_2098);
or U2607 (N_2607,N_2338,N_2465);
or U2608 (N_2608,N_2093,N_2457);
nand U2609 (N_2609,N_2421,N_2059);
or U2610 (N_2610,N_2281,N_2399);
or U2611 (N_2611,N_2241,N_2156);
nand U2612 (N_2612,N_2273,N_2350);
nand U2613 (N_2613,N_2154,N_2435);
nor U2614 (N_2614,N_2406,N_2316);
nand U2615 (N_2615,N_2125,N_2486);
or U2616 (N_2616,N_2265,N_2016);
and U2617 (N_2617,N_2416,N_2152);
or U2618 (N_2618,N_2260,N_2103);
or U2619 (N_2619,N_2382,N_2424);
nand U2620 (N_2620,N_2201,N_2072);
or U2621 (N_2621,N_2147,N_2204);
and U2622 (N_2622,N_2413,N_2003);
and U2623 (N_2623,N_2477,N_2483);
or U2624 (N_2624,N_2258,N_2256);
nor U2625 (N_2625,N_2170,N_2010);
and U2626 (N_2626,N_2324,N_2353);
and U2627 (N_2627,N_2439,N_2410);
nor U2628 (N_2628,N_2292,N_2417);
and U2629 (N_2629,N_2207,N_2377);
or U2630 (N_2630,N_2277,N_2235);
nand U2631 (N_2631,N_2294,N_2078);
or U2632 (N_2632,N_2153,N_2450);
and U2633 (N_2633,N_2092,N_2264);
nor U2634 (N_2634,N_2105,N_2405);
or U2635 (N_2635,N_2212,N_2357);
nand U2636 (N_2636,N_2238,N_2411);
and U2637 (N_2637,N_2049,N_2485);
and U2638 (N_2638,N_2387,N_2491);
nand U2639 (N_2639,N_2346,N_2361);
and U2640 (N_2640,N_2494,N_2060);
nor U2641 (N_2641,N_2303,N_2185);
and U2642 (N_2642,N_2309,N_2055);
or U2643 (N_2643,N_2276,N_2091);
nor U2644 (N_2644,N_2499,N_2400);
nor U2645 (N_2645,N_2000,N_2290);
nand U2646 (N_2646,N_2195,N_2478);
and U2647 (N_2647,N_2284,N_2037);
nand U2648 (N_2648,N_2165,N_2432);
nor U2649 (N_2649,N_2243,N_2214);
or U2650 (N_2650,N_2024,N_2100);
nand U2651 (N_2651,N_2233,N_2176);
or U2652 (N_2652,N_2094,N_2369);
nor U2653 (N_2653,N_2075,N_2222);
or U2654 (N_2654,N_2126,N_2315);
and U2655 (N_2655,N_2084,N_2088);
nand U2656 (N_2656,N_2371,N_2056);
nor U2657 (N_2657,N_2083,N_2471);
or U2658 (N_2658,N_2197,N_2221);
or U2659 (N_2659,N_2328,N_2096);
nor U2660 (N_2660,N_2138,N_2326);
or U2661 (N_2661,N_2048,N_2442);
nand U2662 (N_2662,N_2145,N_2025);
and U2663 (N_2663,N_2236,N_2229);
or U2664 (N_2664,N_2420,N_2133);
and U2665 (N_2665,N_2191,N_2157);
nor U2666 (N_2666,N_2071,N_2419);
and U2667 (N_2667,N_2164,N_2068);
nand U2668 (N_2668,N_2440,N_2226);
and U2669 (N_2669,N_2380,N_2005);
nor U2670 (N_2670,N_2268,N_2239);
nor U2671 (N_2671,N_2388,N_2042);
and U2672 (N_2672,N_2384,N_2307);
or U2673 (N_2673,N_2476,N_2402);
nand U2674 (N_2674,N_2082,N_2272);
and U2675 (N_2675,N_2081,N_2469);
or U2676 (N_2676,N_2266,N_2041);
or U2677 (N_2677,N_2310,N_2087);
nor U2678 (N_2678,N_2458,N_2194);
and U2679 (N_2679,N_2030,N_2352);
nand U2680 (N_2680,N_2143,N_2381);
and U2681 (N_2681,N_2489,N_2379);
or U2682 (N_2682,N_2472,N_2360);
or U2683 (N_2683,N_2367,N_2181);
nand U2684 (N_2684,N_2445,N_2370);
and U2685 (N_2685,N_2351,N_2415);
nand U2686 (N_2686,N_2107,N_2365);
or U2687 (N_2687,N_2497,N_2378);
nand U2688 (N_2688,N_2473,N_2114);
or U2689 (N_2689,N_2189,N_2449);
nand U2690 (N_2690,N_2255,N_2430);
xnor U2691 (N_2691,N_2203,N_2313);
and U2692 (N_2692,N_2175,N_2215);
nor U2693 (N_2693,N_2120,N_2261);
nand U2694 (N_2694,N_2342,N_2278);
nor U2695 (N_2695,N_2337,N_2021);
or U2696 (N_2696,N_2141,N_2246);
nor U2697 (N_2697,N_2356,N_2366);
and U2698 (N_2698,N_2341,N_2250);
or U2699 (N_2699,N_2347,N_2295);
and U2700 (N_2700,N_2285,N_2245);
or U2701 (N_2701,N_2026,N_2023);
or U2702 (N_2702,N_2184,N_2205);
and U2703 (N_2703,N_2394,N_2089);
and U2704 (N_2704,N_2385,N_2033);
nand U2705 (N_2705,N_2045,N_2198);
and U2706 (N_2706,N_2456,N_2343);
or U2707 (N_2707,N_2102,N_2182);
and U2708 (N_2708,N_2468,N_2269);
or U2709 (N_2709,N_2146,N_2355);
nand U2710 (N_2710,N_2135,N_2463);
or U2711 (N_2711,N_2172,N_2119);
and U2712 (N_2712,N_2302,N_2348);
nor U2713 (N_2713,N_2418,N_2101);
and U2714 (N_2714,N_2257,N_2300);
and U2715 (N_2715,N_2208,N_2095);
and U2716 (N_2716,N_2425,N_2227);
or U2717 (N_2717,N_2231,N_2299);
nand U2718 (N_2718,N_2496,N_2368);
nor U2719 (N_2719,N_2280,N_2148);
or U2720 (N_2720,N_2110,N_2446);
and U2721 (N_2721,N_2482,N_2202);
or U2722 (N_2722,N_2106,N_2020);
or U2723 (N_2723,N_2151,N_2253);
nand U2724 (N_2724,N_2168,N_2414);
xor U2725 (N_2725,N_2079,N_2206);
or U2726 (N_2726,N_2219,N_2327);
xnor U2727 (N_2727,N_2484,N_2271);
nor U2728 (N_2728,N_2220,N_2466);
nand U2729 (N_2729,N_2032,N_2454);
nor U2730 (N_2730,N_2282,N_2006);
nand U2731 (N_2731,N_2392,N_2283);
nor U2732 (N_2732,N_2301,N_2460);
nor U2733 (N_2733,N_2062,N_2362);
nor U2734 (N_2734,N_2053,N_2329);
nor U2735 (N_2735,N_2113,N_2317);
nor U2736 (N_2736,N_2234,N_2090);
or U2737 (N_2737,N_2036,N_2008);
xor U2738 (N_2738,N_2051,N_2254);
or U2739 (N_2739,N_2061,N_2358);
and U2740 (N_2740,N_2139,N_2467);
and U2741 (N_2741,N_2196,N_2331);
or U2742 (N_2742,N_2015,N_2462);
nor U2743 (N_2743,N_2122,N_2481);
nor U2744 (N_2744,N_2373,N_2002);
xor U2745 (N_2745,N_2242,N_2314);
or U2746 (N_2746,N_2390,N_2383);
nand U2747 (N_2747,N_2130,N_2086);
nor U2748 (N_2748,N_2259,N_2179);
or U2749 (N_2749,N_2180,N_2431);
nor U2750 (N_2750,N_2204,N_2323);
or U2751 (N_2751,N_2415,N_2263);
nor U2752 (N_2752,N_2494,N_2147);
and U2753 (N_2753,N_2290,N_2118);
nor U2754 (N_2754,N_2467,N_2373);
nor U2755 (N_2755,N_2319,N_2165);
nor U2756 (N_2756,N_2358,N_2210);
nand U2757 (N_2757,N_2085,N_2108);
nor U2758 (N_2758,N_2209,N_2221);
nand U2759 (N_2759,N_2078,N_2221);
nor U2760 (N_2760,N_2053,N_2312);
and U2761 (N_2761,N_2224,N_2056);
and U2762 (N_2762,N_2349,N_2091);
nor U2763 (N_2763,N_2287,N_2462);
nor U2764 (N_2764,N_2228,N_2204);
nand U2765 (N_2765,N_2256,N_2040);
nand U2766 (N_2766,N_2232,N_2091);
or U2767 (N_2767,N_2345,N_2035);
nand U2768 (N_2768,N_2223,N_2305);
nand U2769 (N_2769,N_2364,N_2099);
nand U2770 (N_2770,N_2484,N_2175);
and U2771 (N_2771,N_2422,N_2486);
nor U2772 (N_2772,N_2301,N_2310);
xor U2773 (N_2773,N_2060,N_2463);
and U2774 (N_2774,N_2008,N_2280);
nand U2775 (N_2775,N_2109,N_2411);
nor U2776 (N_2776,N_2151,N_2057);
nor U2777 (N_2777,N_2100,N_2486);
and U2778 (N_2778,N_2483,N_2316);
nand U2779 (N_2779,N_2472,N_2274);
nor U2780 (N_2780,N_2180,N_2086);
nor U2781 (N_2781,N_2465,N_2146);
nand U2782 (N_2782,N_2165,N_2188);
nor U2783 (N_2783,N_2450,N_2276);
nand U2784 (N_2784,N_2258,N_2040);
nand U2785 (N_2785,N_2320,N_2367);
nor U2786 (N_2786,N_2114,N_2176);
nor U2787 (N_2787,N_2270,N_2066);
nand U2788 (N_2788,N_2068,N_2321);
nor U2789 (N_2789,N_2166,N_2281);
and U2790 (N_2790,N_2153,N_2373);
xnor U2791 (N_2791,N_2193,N_2005);
nor U2792 (N_2792,N_2413,N_2174);
nor U2793 (N_2793,N_2132,N_2015);
and U2794 (N_2794,N_2028,N_2290);
or U2795 (N_2795,N_2343,N_2470);
and U2796 (N_2796,N_2418,N_2298);
nor U2797 (N_2797,N_2490,N_2079);
nor U2798 (N_2798,N_2268,N_2180);
and U2799 (N_2799,N_2048,N_2192);
nor U2800 (N_2800,N_2414,N_2182);
and U2801 (N_2801,N_2187,N_2390);
nor U2802 (N_2802,N_2168,N_2357);
or U2803 (N_2803,N_2078,N_2073);
nand U2804 (N_2804,N_2136,N_2275);
or U2805 (N_2805,N_2483,N_2117);
or U2806 (N_2806,N_2204,N_2258);
or U2807 (N_2807,N_2281,N_2394);
and U2808 (N_2808,N_2029,N_2108);
nor U2809 (N_2809,N_2091,N_2495);
nor U2810 (N_2810,N_2428,N_2287);
nand U2811 (N_2811,N_2362,N_2002);
nand U2812 (N_2812,N_2317,N_2254);
or U2813 (N_2813,N_2064,N_2208);
and U2814 (N_2814,N_2089,N_2132);
and U2815 (N_2815,N_2185,N_2462);
or U2816 (N_2816,N_2466,N_2245);
nor U2817 (N_2817,N_2067,N_2232);
nor U2818 (N_2818,N_2241,N_2300);
or U2819 (N_2819,N_2434,N_2160);
or U2820 (N_2820,N_2226,N_2118);
nor U2821 (N_2821,N_2374,N_2182);
xor U2822 (N_2822,N_2009,N_2114);
nor U2823 (N_2823,N_2084,N_2095);
nand U2824 (N_2824,N_2133,N_2124);
xnor U2825 (N_2825,N_2492,N_2072);
nor U2826 (N_2826,N_2389,N_2226);
or U2827 (N_2827,N_2496,N_2112);
and U2828 (N_2828,N_2213,N_2404);
nor U2829 (N_2829,N_2405,N_2267);
nand U2830 (N_2830,N_2275,N_2092);
and U2831 (N_2831,N_2062,N_2057);
nor U2832 (N_2832,N_2092,N_2004);
nor U2833 (N_2833,N_2311,N_2389);
nand U2834 (N_2834,N_2176,N_2074);
xor U2835 (N_2835,N_2265,N_2047);
nor U2836 (N_2836,N_2326,N_2130);
nand U2837 (N_2837,N_2474,N_2413);
and U2838 (N_2838,N_2180,N_2251);
and U2839 (N_2839,N_2027,N_2361);
nor U2840 (N_2840,N_2494,N_2032);
nor U2841 (N_2841,N_2290,N_2289);
nor U2842 (N_2842,N_2336,N_2436);
nor U2843 (N_2843,N_2178,N_2404);
nand U2844 (N_2844,N_2068,N_2276);
nand U2845 (N_2845,N_2471,N_2106);
nand U2846 (N_2846,N_2490,N_2477);
nor U2847 (N_2847,N_2107,N_2451);
nor U2848 (N_2848,N_2096,N_2082);
or U2849 (N_2849,N_2317,N_2363);
and U2850 (N_2850,N_2333,N_2254);
or U2851 (N_2851,N_2434,N_2483);
or U2852 (N_2852,N_2328,N_2117);
xor U2853 (N_2853,N_2495,N_2122);
nand U2854 (N_2854,N_2412,N_2470);
and U2855 (N_2855,N_2422,N_2021);
nand U2856 (N_2856,N_2383,N_2208);
nand U2857 (N_2857,N_2304,N_2032);
nand U2858 (N_2858,N_2056,N_2395);
nand U2859 (N_2859,N_2413,N_2046);
nor U2860 (N_2860,N_2142,N_2246);
nor U2861 (N_2861,N_2141,N_2283);
or U2862 (N_2862,N_2155,N_2325);
nand U2863 (N_2863,N_2007,N_2115);
nor U2864 (N_2864,N_2279,N_2235);
and U2865 (N_2865,N_2470,N_2429);
nand U2866 (N_2866,N_2342,N_2416);
or U2867 (N_2867,N_2307,N_2357);
xnor U2868 (N_2868,N_2232,N_2267);
and U2869 (N_2869,N_2443,N_2350);
nor U2870 (N_2870,N_2466,N_2155);
nor U2871 (N_2871,N_2363,N_2007);
nand U2872 (N_2872,N_2393,N_2349);
and U2873 (N_2873,N_2119,N_2438);
nor U2874 (N_2874,N_2330,N_2323);
nor U2875 (N_2875,N_2247,N_2475);
and U2876 (N_2876,N_2222,N_2195);
nor U2877 (N_2877,N_2188,N_2242);
nor U2878 (N_2878,N_2301,N_2290);
and U2879 (N_2879,N_2173,N_2219);
or U2880 (N_2880,N_2356,N_2309);
and U2881 (N_2881,N_2229,N_2135);
and U2882 (N_2882,N_2449,N_2161);
nor U2883 (N_2883,N_2050,N_2490);
or U2884 (N_2884,N_2137,N_2341);
nand U2885 (N_2885,N_2373,N_2205);
xor U2886 (N_2886,N_2464,N_2449);
or U2887 (N_2887,N_2180,N_2214);
or U2888 (N_2888,N_2164,N_2427);
and U2889 (N_2889,N_2001,N_2227);
nand U2890 (N_2890,N_2311,N_2373);
nor U2891 (N_2891,N_2359,N_2440);
nand U2892 (N_2892,N_2302,N_2299);
and U2893 (N_2893,N_2415,N_2131);
and U2894 (N_2894,N_2358,N_2399);
nor U2895 (N_2895,N_2376,N_2009);
nor U2896 (N_2896,N_2335,N_2481);
nor U2897 (N_2897,N_2390,N_2136);
nor U2898 (N_2898,N_2019,N_2378);
nor U2899 (N_2899,N_2304,N_2178);
and U2900 (N_2900,N_2175,N_2310);
nand U2901 (N_2901,N_2136,N_2364);
nand U2902 (N_2902,N_2147,N_2412);
and U2903 (N_2903,N_2016,N_2013);
or U2904 (N_2904,N_2248,N_2025);
and U2905 (N_2905,N_2238,N_2415);
nand U2906 (N_2906,N_2060,N_2135);
nor U2907 (N_2907,N_2088,N_2303);
and U2908 (N_2908,N_2292,N_2277);
or U2909 (N_2909,N_2243,N_2036);
or U2910 (N_2910,N_2303,N_2443);
nand U2911 (N_2911,N_2454,N_2110);
and U2912 (N_2912,N_2365,N_2192);
and U2913 (N_2913,N_2224,N_2041);
and U2914 (N_2914,N_2452,N_2405);
nand U2915 (N_2915,N_2280,N_2189);
or U2916 (N_2916,N_2214,N_2342);
nand U2917 (N_2917,N_2128,N_2182);
nand U2918 (N_2918,N_2346,N_2037);
nand U2919 (N_2919,N_2260,N_2351);
and U2920 (N_2920,N_2292,N_2471);
and U2921 (N_2921,N_2124,N_2077);
nand U2922 (N_2922,N_2061,N_2486);
nor U2923 (N_2923,N_2431,N_2194);
or U2924 (N_2924,N_2167,N_2283);
and U2925 (N_2925,N_2195,N_2026);
xor U2926 (N_2926,N_2260,N_2043);
nor U2927 (N_2927,N_2137,N_2451);
and U2928 (N_2928,N_2029,N_2291);
and U2929 (N_2929,N_2366,N_2059);
nor U2930 (N_2930,N_2359,N_2219);
and U2931 (N_2931,N_2160,N_2228);
or U2932 (N_2932,N_2213,N_2196);
or U2933 (N_2933,N_2493,N_2002);
or U2934 (N_2934,N_2113,N_2417);
nand U2935 (N_2935,N_2020,N_2118);
nand U2936 (N_2936,N_2309,N_2070);
nor U2937 (N_2937,N_2270,N_2085);
and U2938 (N_2938,N_2044,N_2043);
nand U2939 (N_2939,N_2354,N_2420);
or U2940 (N_2940,N_2092,N_2060);
nand U2941 (N_2941,N_2226,N_2314);
nand U2942 (N_2942,N_2202,N_2358);
and U2943 (N_2943,N_2470,N_2007);
nor U2944 (N_2944,N_2410,N_2074);
nand U2945 (N_2945,N_2419,N_2342);
or U2946 (N_2946,N_2014,N_2299);
and U2947 (N_2947,N_2061,N_2343);
nor U2948 (N_2948,N_2271,N_2137);
or U2949 (N_2949,N_2402,N_2396);
or U2950 (N_2950,N_2131,N_2411);
xnor U2951 (N_2951,N_2488,N_2274);
nand U2952 (N_2952,N_2361,N_2006);
and U2953 (N_2953,N_2207,N_2401);
nor U2954 (N_2954,N_2223,N_2052);
nand U2955 (N_2955,N_2352,N_2355);
and U2956 (N_2956,N_2251,N_2012);
or U2957 (N_2957,N_2371,N_2422);
or U2958 (N_2958,N_2058,N_2063);
or U2959 (N_2959,N_2395,N_2012);
or U2960 (N_2960,N_2109,N_2353);
and U2961 (N_2961,N_2028,N_2466);
nor U2962 (N_2962,N_2254,N_2128);
nand U2963 (N_2963,N_2444,N_2344);
nor U2964 (N_2964,N_2305,N_2356);
nor U2965 (N_2965,N_2497,N_2395);
nand U2966 (N_2966,N_2053,N_2073);
and U2967 (N_2967,N_2307,N_2239);
or U2968 (N_2968,N_2153,N_2203);
or U2969 (N_2969,N_2094,N_2467);
and U2970 (N_2970,N_2108,N_2232);
and U2971 (N_2971,N_2102,N_2400);
and U2972 (N_2972,N_2024,N_2485);
and U2973 (N_2973,N_2446,N_2062);
and U2974 (N_2974,N_2258,N_2468);
nand U2975 (N_2975,N_2324,N_2029);
nand U2976 (N_2976,N_2054,N_2075);
nand U2977 (N_2977,N_2409,N_2145);
and U2978 (N_2978,N_2476,N_2293);
and U2979 (N_2979,N_2472,N_2272);
and U2980 (N_2980,N_2080,N_2454);
or U2981 (N_2981,N_2165,N_2284);
or U2982 (N_2982,N_2076,N_2258);
or U2983 (N_2983,N_2112,N_2129);
nand U2984 (N_2984,N_2309,N_2093);
nor U2985 (N_2985,N_2177,N_2080);
nand U2986 (N_2986,N_2309,N_2473);
nand U2987 (N_2987,N_2210,N_2303);
nand U2988 (N_2988,N_2270,N_2274);
nand U2989 (N_2989,N_2262,N_2123);
nor U2990 (N_2990,N_2185,N_2271);
nand U2991 (N_2991,N_2441,N_2496);
or U2992 (N_2992,N_2399,N_2364);
nor U2993 (N_2993,N_2417,N_2496);
or U2994 (N_2994,N_2036,N_2162);
and U2995 (N_2995,N_2414,N_2326);
and U2996 (N_2996,N_2395,N_2061);
nand U2997 (N_2997,N_2212,N_2029);
and U2998 (N_2998,N_2074,N_2262);
or U2999 (N_2999,N_2449,N_2286);
nor UO_0 (O_0,N_2960,N_2730);
or UO_1 (O_1,N_2878,N_2552);
and UO_2 (O_2,N_2614,N_2754);
nor UO_3 (O_3,N_2737,N_2965);
nor UO_4 (O_4,N_2873,N_2992);
and UO_5 (O_5,N_2951,N_2809);
nand UO_6 (O_6,N_2793,N_2736);
nor UO_7 (O_7,N_2521,N_2905);
or UO_8 (O_8,N_2771,N_2944);
or UO_9 (O_9,N_2916,N_2645);
nor UO_10 (O_10,N_2704,N_2915);
or UO_11 (O_11,N_2538,N_2648);
nor UO_12 (O_12,N_2909,N_2987);
and UO_13 (O_13,N_2925,N_2627);
and UO_14 (O_14,N_2658,N_2655);
nor UO_15 (O_15,N_2852,N_2796);
nor UO_16 (O_16,N_2841,N_2966);
nand UO_17 (O_17,N_2826,N_2632);
xor UO_18 (O_18,N_2767,N_2742);
nor UO_19 (O_19,N_2980,N_2622);
or UO_20 (O_20,N_2586,N_2681);
nand UO_21 (O_21,N_2813,N_2642);
and UO_22 (O_22,N_2696,N_2939);
nor UO_23 (O_23,N_2685,N_2733);
nand UO_24 (O_24,N_2777,N_2518);
nand UO_25 (O_25,N_2663,N_2972);
or UO_26 (O_26,N_2662,N_2956);
nor UO_27 (O_27,N_2723,N_2840);
and UO_28 (O_28,N_2590,N_2759);
nor UO_29 (O_29,N_2516,N_2668);
and UO_30 (O_30,N_2933,N_2805);
and UO_31 (O_31,N_2949,N_2863);
nor UO_32 (O_32,N_2866,N_2531);
and UO_33 (O_33,N_2931,N_2678);
nor UO_34 (O_34,N_2529,N_2541);
or UO_35 (O_35,N_2650,N_2862);
nand UO_36 (O_36,N_2515,N_2692);
and UO_37 (O_37,N_2667,N_2785);
and UO_38 (O_38,N_2691,N_2790);
nand UO_39 (O_39,N_2546,N_2810);
or UO_40 (O_40,N_2540,N_2877);
nor UO_41 (O_41,N_2881,N_2760);
or UO_42 (O_42,N_2528,N_2643);
or UO_43 (O_43,N_2526,N_2930);
and UO_44 (O_44,N_2867,N_2714);
or UO_45 (O_45,N_2695,N_2902);
nor UO_46 (O_46,N_2795,N_2556);
and UO_47 (O_47,N_2783,N_2636);
nor UO_48 (O_48,N_2860,N_2784);
nand UO_49 (O_49,N_2948,N_2698);
or UO_50 (O_50,N_2917,N_2782);
and UO_51 (O_51,N_2690,N_2808);
and UO_52 (O_52,N_2981,N_2578);
or UO_53 (O_53,N_2660,N_2659);
and UO_54 (O_54,N_2848,N_2907);
nand UO_55 (O_55,N_2654,N_2854);
xor UO_56 (O_56,N_2613,N_2510);
and UO_57 (O_57,N_2594,N_2740);
or UO_58 (O_58,N_2670,N_2687);
and UO_59 (O_59,N_2601,N_2787);
or UO_60 (O_60,N_2936,N_2845);
and UO_61 (O_61,N_2514,N_2804);
and UO_62 (O_62,N_2582,N_2911);
and UO_63 (O_63,N_2884,N_2994);
nor UO_64 (O_64,N_2971,N_2503);
or UO_65 (O_65,N_2797,N_2707);
and UO_66 (O_66,N_2729,N_2522);
nand UO_67 (O_67,N_2686,N_2588);
nor UO_68 (O_68,N_2550,N_2768);
nand UO_69 (O_69,N_2587,N_2741);
and UO_70 (O_70,N_2722,N_2638);
nor UO_71 (O_71,N_2975,N_2505);
and UO_72 (O_72,N_2816,N_2812);
nor UO_73 (O_73,N_2637,N_2547);
nor UO_74 (O_74,N_2802,N_2527);
nor UO_75 (O_75,N_2589,N_2864);
nor UO_76 (O_76,N_2605,N_2834);
nor UO_77 (O_77,N_2904,N_2523);
nand UO_78 (O_78,N_2828,N_2525);
nand UO_79 (O_79,N_2892,N_2776);
and UO_80 (O_80,N_2652,N_2616);
and UO_81 (O_81,N_2819,N_2947);
or UO_82 (O_82,N_2563,N_2886);
nand UO_83 (O_83,N_2673,N_2575);
and UO_84 (O_84,N_2815,N_2679);
or UO_85 (O_85,N_2524,N_2548);
nand UO_86 (O_86,N_2739,N_2568);
and UO_87 (O_87,N_2592,N_2702);
and UO_88 (O_88,N_2851,N_2982);
nor UO_89 (O_89,N_2898,N_2830);
nand UO_90 (O_90,N_2928,N_2676);
nand UO_91 (O_91,N_2762,N_2891);
nand UO_92 (O_92,N_2532,N_2969);
and UO_93 (O_93,N_2609,N_2724);
and UO_94 (O_94,N_2718,N_2943);
nor UO_95 (O_95,N_2604,N_2520);
or UO_96 (O_96,N_2836,N_2932);
or UO_97 (O_97,N_2758,N_2500);
and UO_98 (O_98,N_2926,N_2629);
or UO_99 (O_99,N_2850,N_2952);
or UO_100 (O_100,N_2634,N_2572);
nor UO_101 (O_101,N_2746,N_2693);
or UO_102 (O_102,N_2964,N_2842);
nor UO_103 (O_103,N_2619,N_2986);
and UO_104 (O_104,N_2769,N_2856);
nand UO_105 (O_105,N_2651,N_2688);
and UO_106 (O_106,N_2537,N_2913);
and UO_107 (O_107,N_2921,N_2709);
nor UO_108 (O_108,N_2557,N_2630);
or UO_109 (O_109,N_2606,N_2923);
nand UO_110 (O_110,N_2788,N_2720);
nor UO_111 (O_111,N_2879,N_2621);
and UO_112 (O_112,N_2827,N_2983);
nor UO_113 (O_113,N_2791,N_2875);
and UO_114 (O_114,N_2938,N_2779);
or UO_115 (O_115,N_2927,N_2753);
and UO_116 (O_116,N_2677,N_2935);
nor UO_117 (O_117,N_2833,N_2874);
and UO_118 (O_118,N_2897,N_2990);
and UO_119 (O_119,N_2647,N_2978);
and UO_120 (O_120,N_2504,N_2998);
and UO_121 (O_121,N_2910,N_2901);
nor UO_122 (O_122,N_2542,N_2774);
nor UO_123 (O_123,N_2764,N_2896);
nand UO_124 (O_124,N_2789,N_2993);
nor UO_125 (O_125,N_2567,N_2708);
nor UO_126 (O_126,N_2562,N_2991);
or UO_127 (O_127,N_2888,N_2639);
or UO_128 (O_128,N_2700,N_2817);
nor UO_129 (O_129,N_2626,N_2835);
nor UO_130 (O_130,N_2801,N_2940);
nand UO_131 (O_131,N_2745,N_2735);
nand UO_132 (O_132,N_2871,N_2853);
and UO_133 (O_133,N_2988,N_2876);
nand UO_134 (O_134,N_2569,N_2780);
nand UO_135 (O_135,N_2807,N_2974);
or UO_136 (O_136,N_2599,N_2880);
nor UO_137 (O_137,N_2766,N_2890);
or UO_138 (O_138,N_2560,N_2608);
nor UO_139 (O_139,N_2544,N_2914);
or UO_140 (O_140,N_2976,N_2640);
or UO_141 (O_141,N_2749,N_2501);
and UO_142 (O_142,N_2765,N_2574);
or UO_143 (O_143,N_2946,N_2732);
or UO_144 (O_144,N_2712,N_2600);
nand UO_145 (O_145,N_2653,N_2832);
nor UO_146 (O_146,N_2738,N_2573);
nand UO_147 (O_147,N_2674,N_2953);
or UO_148 (O_148,N_2744,N_2962);
nor UO_149 (O_149,N_2803,N_2664);
nand UO_150 (O_150,N_2752,N_2814);
nand UO_151 (O_151,N_2607,N_2644);
and UO_152 (O_152,N_2502,N_2584);
nand UO_153 (O_153,N_2872,N_2699);
and UO_154 (O_154,N_2822,N_2612);
and UO_155 (O_155,N_2564,N_2773);
or UO_156 (O_156,N_2716,N_2671);
nor UO_157 (O_157,N_2770,N_2615);
nor UO_158 (O_158,N_2549,N_2628);
or UO_159 (O_159,N_2519,N_2581);
nand UO_160 (O_160,N_2649,N_2508);
or UO_161 (O_161,N_2530,N_2535);
nand UO_162 (O_162,N_2979,N_2750);
and UO_163 (O_163,N_2989,N_2610);
nor UO_164 (O_164,N_2543,N_2843);
nor UO_165 (O_165,N_2908,N_2625);
nand UO_166 (O_166,N_2798,N_2967);
nand UO_167 (O_167,N_2893,N_2846);
nor UO_168 (O_168,N_2726,N_2997);
nand UO_169 (O_169,N_2857,N_2887);
or UO_170 (O_170,N_2585,N_2763);
and UO_171 (O_171,N_2799,N_2961);
or UO_172 (O_172,N_2558,N_2995);
and UO_173 (O_173,N_2984,N_2900);
or UO_174 (O_174,N_2977,N_2715);
nor UO_175 (O_175,N_2641,N_2885);
and UO_176 (O_176,N_2684,N_2838);
nand UO_177 (O_177,N_2823,N_2682);
nand UO_178 (O_178,N_2924,N_2985);
or UO_179 (O_179,N_2706,N_2761);
and UO_180 (O_180,N_2533,N_2861);
nor UO_181 (O_181,N_2577,N_2849);
nor UO_182 (O_182,N_2595,N_2565);
nor UO_183 (O_183,N_2618,N_2747);
nor UO_184 (O_184,N_2922,N_2603);
nand UO_185 (O_185,N_2945,N_2539);
nor UO_186 (O_186,N_2869,N_2839);
or UO_187 (O_187,N_2999,N_2680);
nor UO_188 (O_188,N_2536,N_2689);
and UO_189 (O_189,N_2666,N_2781);
nand UO_190 (O_190,N_2882,N_2942);
and UO_191 (O_191,N_2868,N_2786);
xor UO_192 (O_192,N_2870,N_2545);
or UO_193 (O_193,N_2576,N_2919);
nor UO_194 (O_194,N_2847,N_2561);
or UO_195 (O_195,N_2955,N_2566);
nor UO_196 (O_196,N_2617,N_2941);
and UO_197 (O_197,N_2865,N_2748);
or UO_198 (O_198,N_2937,N_2683);
and UO_199 (O_199,N_2705,N_2623);
and UO_200 (O_200,N_2509,N_2855);
nand UO_201 (O_201,N_2602,N_2710);
nor UO_202 (O_202,N_2656,N_2513);
and UO_203 (O_203,N_2958,N_2811);
nand UO_204 (O_204,N_2772,N_2713);
nand UO_205 (O_205,N_2725,N_2775);
and UO_206 (O_206,N_2968,N_2721);
nand UO_207 (O_207,N_2507,N_2829);
nor UO_208 (O_208,N_2511,N_2889);
nand UO_209 (O_209,N_2934,N_2593);
or UO_210 (O_210,N_2597,N_2818);
nand UO_211 (O_211,N_2611,N_2895);
nor UO_212 (O_212,N_2957,N_2734);
nand UO_213 (O_213,N_2727,N_2570);
and UO_214 (O_214,N_2824,N_2620);
nor UO_215 (O_215,N_2583,N_2920);
and UO_216 (O_216,N_2963,N_2598);
nand UO_217 (O_217,N_2675,N_2728);
nor UO_218 (O_218,N_2596,N_2792);
xor UO_219 (O_219,N_2929,N_2717);
and UO_220 (O_220,N_2657,N_2669);
nor UO_221 (O_221,N_2954,N_2756);
and UO_222 (O_222,N_2755,N_2731);
and UO_223 (O_223,N_2778,N_2665);
and UO_224 (O_224,N_2554,N_2831);
nor UO_225 (O_225,N_2899,N_2571);
and UO_226 (O_226,N_2794,N_2631);
or UO_227 (O_227,N_2661,N_2883);
nor UO_228 (O_228,N_2672,N_2743);
nand UO_229 (O_229,N_2806,N_2697);
nand UO_230 (O_230,N_2551,N_2633);
nor UO_231 (O_231,N_2821,N_2973);
and UO_232 (O_232,N_2800,N_2757);
nand UO_233 (O_233,N_2906,N_2959);
nand UO_234 (O_234,N_2559,N_2970);
nor UO_235 (O_235,N_2646,N_2694);
nor UO_236 (O_236,N_2703,N_2579);
nor UO_237 (O_237,N_2837,N_2517);
nor UO_238 (O_238,N_2751,N_2553);
nand UO_239 (O_239,N_2894,N_2506);
nand UO_240 (O_240,N_2918,N_2950);
or UO_241 (O_241,N_2512,N_2858);
or UO_242 (O_242,N_2534,N_2719);
and UO_243 (O_243,N_2820,N_2701);
or UO_244 (O_244,N_2825,N_2555);
and UO_245 (O_245,N_2903,N_2711);
nand UO_246 (O_246,N_2580,N_2912);
nand UO_247 (O_247,N_2859,N_2591);
and UO_248 (O_248,N_2624,N_2996);
and UO_249 (O_249,N_2635,N_2844);
and UO_250 (O_250,N_2610,N_2744);
nor UO_251 (O_251,N_2530,N_2856);
nand UO_252 (O_252,N_2799,N_2891);
nand UO_253 (O_253,N_2957,N_2850);
nand UO_254 (O_254,N_2794,N_2739);
nand UO_255 (O_255,N_2887,N_2847);
and UO_256 (O_256,N_2975,N_2717);
nand UO_257 (O_257,N_2590,N_2540);
and UO_258 (O_258,N_2821,N_2810);
and UO_259 (O_259,N_2652,N_2788);
or UO_260 (O_260,N_2690,N_2978);
and UO_261 (O_261,N_2698,N_2783);
or UO_262 (O_262,N_2613,N_2889);
nand UO_263 (O_263,N_2607,N_2748);
and UO_264 (O_264,N_2537,N_2926);
and UO_265 (O_265,N_2551,N_2776);
or UO_266 (O_266,N_2721,N_2578);
nand UO_267 (O_267,N_2821,N_2705);
nor UO_268 (O_268,N_2932,N_2635);
or UO_269 (O_269,N_2878,N_2621);
nor UO_270 (O_270,N_2625,N_2984);
nor UO_271 (O_271,N_2834,N_2753);
and UO_272 (O_272,N_2727,N_2819);
or UO_273 (O_273,N_2762,N_2950);
and UO_274 (O_274,N_2634,N_2538);
nor UO_275 (O_275,N_2540,N_2896);
and UO_276 (O_276,N_2924,N_2563);
nand UO_277 (O_277,N_2516,N_2750);
or UO_278 (O_278,N_2734,N_2864);
or UO_279 (O_279,N_2882,N_2807);
nor UO_280 (O_280,N_2544,N_2991);
nor UO_281 (O_281,N_2640,N_2589);
or UO_282 (O_282,N_2930,N_2821);
nand UO_283 (O_283,N_2589,N_2754);
nand UO_284 (O_284,N_2725,N_2822);
nand UO_285 (O_285,N_2598,N_2765);
or UO_286 (O_286,N_2850,N_2894);
nand UO_287 (O_287,N_2955,N_2905);
nor UO_288 (O_288,N_2827,N_2882);
nand UO_289 (O_289,N_2948,N_2759);
xor UO_290 (O_290,N_2577,N_2687);
and UO_291 (O_291,N_2787,N_2547);
nor UO_292 (O_292,N_2791,N_2922);
or UO_293 (O_293,N_2893,N_2850);
and UO_294 (O_294,N_2849,N_2843);
and UO_295 (O_295,N_2697,N_2660);
or UO_296 (O_296,N_2976,N_2895);
nor UO_297 (O_297,N_2626,N_2554);
and UO_298 (O_298,N_2507,N_2855);
nor UO_299 (O_299,N_2815,N_2556);
nor UO_300 (O_300,N_2787,N_2956);
and UO_301 (O_301,N_2849,N_2719);
and UO_302 (O_302,N_2863,N_2914);
or UO_303 (O_303,N_2806,N_2746);
nand UO_304 (O_304,N_2586,N_2817);
and UO_305 (O_305,N_2668,N_2917);
and UO_306 (O_306,N_2587,N_2813);
nand UO_307 (O_307,N_2896,N_2633);
nor UO_308 (O_308,N_2969,N_2894);
nor UO_309 (O_309,N_2933,N_2702);
and UO_310 (O_310,N_2536,N_2613);
nand UO_311 (O_311,N_2877,N_2860);
and UO_312 (O_312,N_2719,N_2552);
or UO_313 (O_313,N_2735,N_2937);
nand UO_314 (O_314,N_2771,N_2836);
and UO_315 (O_315,N_2589,N_2975);
nor UO_316 (O_316,N_2662,N_2743);
nor UO_317 (O_317,N_2689,N_2711);
or UO_318 (O_318,N_2983,N_2830);
or UO_319 (O_319,N_2965,N_2695);
nand UO_320 (O_320,N_2866,N_2523);
nor UO_321 (O_321,N_2921,N_2928);
and UO_322 (O_322,N_2689,N_2903);
nand UO_323 (O_323,N_2939,N_2683);
nand UO_324 (O_324,N_2634,N_2516);
and UO_325 (O_325,N_2878,N_2681);
nor UO_326 (O_326,N_2500,N_2963);
and UO_327 (O_327,N_2753,N_2998);
nand UO_328 (O_328,N_2726,N_2999);
or UO_329 (O_329,N_2620,N_2633);
nand UO_330 (O_330,N_2806,N_2506);
nand UO_331 (O_331,N_2917,N_2532);
nor UO_332 (O_332,N_2673,N_2587);
nand UO_333 (O_333,N_2896,N_2614);
nor UO_334 (O_334,N_2915,N_2787);
and UO_335 (O_335,N_2724,N_2925);
nor UO_336 (O_336,N_2729,N_2712);
or UO_337 (O_337,N_2838,N_2630);
and UO_338 (O_338,N_2937,N_2553);
nand UO_339 (O_339,N_2581,N_2655);
nor UO_340 (O_340,N_2717,N_2772);
nor UO_341 (O_341,N_2617,N_2549);
or UO_342 (O_342,N_2841,N_2520);
nand UO_343 (O_343,N_2522,N_2545);
nor UO_344 (O_344,N_2992,N_2849);
or UO_345 (O_345,N_2654,N_2716);
or UO_346 (O_346,N_2636,N_2694);
nand UO_347 (O_347,N_2978,N_2747);
nand UO_348 (O_348,N_2969,N_2881);
or UO_349 (O_349,N_2518,N_2551);
and UO_350 (O_350,N_2537,N_2627);
nand UO_351 (O_351,N_2530,N_2729);
or UO_352 (O_352,N_2975,N_2721);
nand UO_353 (O_353,N_2609,N_2818);
nor UO_354 (O_354,N_2799,N_2596);
nand UO_355 (O_355,N_2923,N_2509);
nand UO_356 (O_356,N_2674,N_2976);
or UO_357 (O_357,N_2948,N_2592);
and UO_358 (O_358,N_2664,N_2907);
nand UO_359 (O_359,N_2941,N_2769);
or UO_360 (O_360,N_2983,N_2631);
nor UO_361 (O_361,N_2821,N_2591);
nor UO_362 (O_362,N_2548,N_2813);
nand UO_363 (O_363,N_2993,N_2503);
and UO_364 (O_364,N_2569,N_2598);
nand UO_365 (O_365,N_2504,N_2548);
nand UO_366 (O_366,N_2974,N_2541);
nand UO_367 (O_367,N_2857,N_2504);
and UO_368 (O_368,N_2840,N_2692);
and UO_369 (O_369,N_2559,N_2551);
nor UO_370 (O_370,N_2752,N_2899);
and UO_371 (O_371,N_2702,N_2701);
and UO_372 (O_372,N_2958,N_2980);
and UO_373 (O_373,N_2892,N_2844);
nand UO_374 (O_374,N_2782,N_2575);
and UO_375 (O_375,N_2920,N_2650);
and UO_376 (O_376,N_2847,N_2705);
nor UO_377 (O_377,N_2733,N_2705);
and UO_378 (O_378,N_2956,N_2901);
or UO_379 (O_379,N_2890,N_2822);
nand UO_380 (O_380,N_2590,N_2747);
nor UO_381 (O_381,N_2742,N_2917);
or UO_382 (O_382,N_2670,N_2785);
or UO_383 (O_383,N_2541,N_2565);
and UO_384 (O_384,N_2791,N_2723);
nor UO_385 (O_385,N_2972,N_2782);
and UO_386 (O_386,N_2551,N_2770);
nor UO_387 (O_387,N_2980,N_2950);
or UO_388 (O_388,N_2969,N_2932);
or UO_389 (O_389,N_2970,N_2673);
nor UO_390 (O_390,N_2856,N_2605);
nor UO_391 (O_391,N_2780,N_2652);
nand UO_392 (O_392,N_2968,N_2793);
or UO_393 (O_393,N_2738,N_2845);
and UO_394 (O_394,N_2654,N_2657);
nand UO_395 (O_395,N_2756,N_2702);
nor UO_396 (O_396,N_2658,N_2886);
nand UO_397 (O_397,N_2714,N_2724);
and UO_398 (O_398,N_2746,N_2807);
xor UO_399 (O_399,N_2893,N_2797);
nor UO_400 (O_400,N_2515,N_2566);
and UO_401 (O_401,N_2838,N_2834);
nor UO_402 (O_402,N_2823,N_2929);
and UO_403 (O_403,N_2631,N_2614);
nand UO_404 (O_404,N_2536,N_2998);
nand UO_405 (O_405,N_2638,N_2941);
nand UO_406 (O_406,N_2569,N_2918);
and UO_407 (O_407,N_2789,N_2927);
nor UO_408 (O_408,N_2978,N_2708);
nor UO_409 (O_409,N_2916,N_2860);
or UO_410 (O_410,N_2783,N_2992);
and UO_411 (O_411,N_2510,N_2789);
nor UO_412 (O_412,N_2516,N_2951);
nor UO_413 (O_413,N_2823,N_2956);
or UO_414 (O_414,N_2643,N_2704);
nand UO_415 (O_415,N_2898,N_2779);
nor UO_416 (O_416,N_2892,N_2624);
or UO_417 (O_417,N_2654,N_2955);
nor UO_418 (O_418,N_2770,N_2794);
nand UO_419 (O_419,N_2534,N_2742);
and UO_420 (O_420,N_2520,N_2661);
and UO_421 (O_421,N_2829,N_2979);
or UO_422 (O_422,N_2599,N_2972);
nor UO_423 (O_423,N_2971,N_2865);
or UO_424 (O_424,N_2796,N_2840);
nand UO_425 (O_425,N_2713,N_2892);
nor UO_426 (O_426,N_2772,N_2641);
xnor UO_427 (O_427,N_2849,N_2628);
nand UO_428 (O_428,N_2509,N_2578);
and UO_429 (O_429,N_2970,N_2960);
nor UO_430 (O_430,N_2600,N_2729);
nor UO_431 (O_431,N_2968,N_2637);
nand UO_432 (O_432,N_2839,N_2614);
nand UO_433 (O_433,N_2907,N_2924);
nand UO_434 (O_434,N_2786,N_2908);
nand UO_435 (O_435,N_2594,N_2986);
or UO_436 (O_436,N_2858,N_2738);
nor UO_437 (O_437,N_2745,N_2556);
and UO_438 (O_438,N_2684,N_2712);
or UO_439 (O_439,N_2967,N_2896);
nand UO_440 (O_440,N_2596,N_2726);
or UO_441 (O_441,N_2875,N_2956);
or UO_442 (O_442,N_2583,N_2953);
nand UO_443 (O_443,N_2711,N_2503);
or UO_444 (O_444,N_2845,N_2519);
nor UO_445 (O_445,N_2517,N_2627);
nor UO_446 (O_446,N_2663,N_2804);
nand UO_447 (O_447,N_2638,N_2748);
and UO_448 (O_448,N_2711,N_2597);
or UO_449 (O_449,N_2575,N_2879);
nand UO_450 (O_450,N_2871,N_2664);
and UO_451 (O_451,N_2935,N_2986);
nor UO_452 (O_452,N_2667,N_2583);
nand UO_453 (O_453,N_2658,N_2510);
or UO_454 (O_454,N_2781,N_2687);
nand UO_455 (O_455,N_2744,N_2959);
xor UO_456 (O_456,N_2706,N_2835);
and UO_457 (O_457,N_2687,N_2753);
and UO_458 (O_458,N_2582,N_2822);
nand UO_459 (O_459,N_2953,N_2581);
nand UO_460 (O_460,N_2504,N_2572);
nor UO_461 (O_461,N_2773,N_2559);
nand UO_462 (O_462,N_2628,N_2993);
nand UO_463 (O_463,N_2552,N_2718);
and UO_464 (O_464,N_2614,N_2630);
nand UO_465 (O_465,N_2663,N_2836);
nand UO_466 (O_466,N_2734,N_2974);
nand UO_467 (O_467,N_2761,N_2518);
nor UO_468 (O_468,N_2792,N_2525);
or UO_469 (O_469,N_2840,N_2968);
and UO_470 (O_470,N_2882,N_2522);
nand UO_471 (O_471,N_2887,N_2910);
or UO_472 (O_472,N_2958,N_2678);
nand UO_473 (O_473,N_2994,N_2685);
and UO_474 (O_474,N_2580,N_2831);
and UO_475 (O_475,N_2583,N_2566);
nand UO_476 (O_476,N_2781,N_2857);
nand UO_477 (O_477,N_2839,N_2824);
nand UO_478 (O_478,N_2702,N_2777);
nor UO_479 (O_479,N_2784,N_2917);
nand UO_480 (O_480,N_2946,N_2857);
nor UO_481 (O_481,N_2843,N_2654);
nor UO_482 (O_482,N_2710,N_2664);
or UO_483 (O_483,N_2787,N_2620);
and UO_484 (O_484,N_2528,N_2586);
nand UO_485 (O_485,N_2993,N_2510);
or UO_486 (O_486,N_2905,N_2694);
nor UO_487 (O_487,N_2930,N_2947);
nor UO_488 (O_488,N_2997,N_2792);
and UO_489 (O_489,N_2635,N_2732);
and UO_490 (O_490,N_2681,N_2838);
nor UO_491 (O_491,N_2841,N_2921);
or UO_492 (O_492,N_2645,N_2724);
nand UO_493 (O_493,N_2886,N_2909);
or UO_494 (O_494,N_2944,N_2934);
or UO_495 (O_495,N_2770,N_2844);
nor UO_496 (O_496,N_2947,N_2666);
or UO_497 (O_497,N_2919,N_2623);
nor UO_498 (O_498,N_2862,N_2918);
nor UO_499 (O_499,N_2611,N_2985);
endmodule