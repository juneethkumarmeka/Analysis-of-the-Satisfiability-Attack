module basic_2000_20000_2500_5_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nand U0 (N_0,In_1691,In_1925);
nor U1 (N_1,In_47,In_1744);
xnor U2 (N_2,In_724,In_747);
nor U3 (N_3,In_391,In_265);
nor U4 (N_4,In_165,In_1884);
nor U5 (N_5,In_1880,In_1549);
nand U6 (N_6,In_822,In_667);
nand U7 (N_7,In_1604,In_609);
nor U8 (N_8,In_138,In_1947);
xor U9 (N_9,In_1521,In_1311);
and U10 (N_10,In_1444,In_741);
nor U11 (N_11,In_1229,In_1175);
and U12 (N_12,In_1700,In_1321);
xnor U13 (N_13,In_34,In_1010);
and U14 (N_14,In_1781,In_1776);
and U15 (N_15,In_72,In_607);
xor U16 (N_16,In_1245,In_517);
and U17 (N_17,In_1657,In_1217);
nand U18 (N_18,In_1663,In_309);
nand U19 (N_19,In_1921,In_1091);
nor U20 (N_20,In_1392,In_826);
nand U21 (N_21,In_136,In_407);
nor U22 (N_22,In_1507,In_1165);
nor U23 (N_23,In_405,In_214);
nor U24 (N_24,In_1149,In_529);
nor U25 (N_25,In_595,In_468);
nand U26 (N_26,In_751,In_1067);
nand U27 (N_27,In_1068,In_1591);
nor U28 (N_28,In_1757,In_1096);
or U29 (N_29,In_764,In_1435);
nand U30 (N_30,In_1734,In_455);
xnor U31 (N_31,In_24,In_1991);
and U32 (N_32,In_1942,In_660);
nor U33 (N_33,In_1467,In_1395);
nand U34 (N_34,In_1054,In_723);
nor U35 (N_35,In_1473,In_1794);
or U36 (N_36,In_27,In_750);
and U37 (N_37,In_1178,In_1851);
or U38 (N_38,In_549,In_645);
or U39 (N_39,In_838,In_1584);
nand U40 (N_40,In_426,In_1737);
or U41 (N_41,In_1348,In_132);
or U42 (N_42,In_489,In_900);
nand U43 (N_43,In_1650,In_1709);
xnor U44 (N_44,In_1556,In_185);
xor U45 (N_45,In_1423,In_762);
and U46 (N_46,In_913,In_627);
or U47 (N_47,In_1483,In_1579);
nor U48 (N_48,In_1014,In_1544);
or U49 (N_49,In_1751,In_1920);
and U50 (N_50,In_226,In_1222);
nor U51 (N_51,In_1249,In_883);
and U52 (N_52,In_401,In_1971);
nand U53 (N_53,In_470,In_654);
nand U54 (N_54,In_1258,In_1923);
or U55 (N_55,In_1858,In_87);
and U56 (N_56,In_1466,In_676);
nor U57 (N_57,In_61,In_453);
xor U58 (N_58,In_230,In_753);
and U59 (N_59,In_933,In_780);
nand U60 (N_60,In_596,In_1257);
xor U61 (N_61,In_1793,In_1083);
or U62 (N_62,In_263,In_222);
nor U63 (N_63,In_1824,In_504);
or U64 (N_64,In_111,In_1397);
and U65 (N_65,In_224,In_1902);
or U66 (N_66,In_1020,In_431);
xor U67 (N_67,In_618,In_1834);
or U68 (N_68,In_178,In_1883);
xnor U69 (N_69,In_606,In_1255);
and U70 (N_70,In_1652,In_40);
nand U71 (N_71,In_819,In_1580);
nand U72 (N_72,In_1050,In_1280);
and U73 (N_73,In_243,In_802);
or U74 (N_74,In_610,In_1551);
and U75 (N_75,In_1537,In_691);
and U76 (N_76,In_887,In_63);
xor U77 (N_77,In_1957,In_1189);
or U78 (N_78,In_76,In_663);
xnor U79 (N_79,In_408,In_698);
nor U80 (N_80,In_1148,In_1132);
nand U81 (N_81,In_1837,In_1973);
xnor U82 (N_82,In_97,In_1845);
xnor U83 (N_83,In_1384,In_1898);
xnor U84 (N_84,In_1320,In_1689);
nor U85 (N_85,In_443,In_1351);
and U86 (N_86,In_264,In_1574);
nand U87 (N_87,In_460,In_1388);
xor U88 (N_88,In_808,In_54);
or U89 (N_89,In_1586,In_1156);
nand U90 (N_90,In_604,In_1241);
xnor U91 (N_91,In_535,In_1716);
and U92 (N_92,In_1200,In_1823);
and U93 (N_93,In_1949,In_547);
nor U94 (N_94,In_1021,In_938);
and U95 (N_95,In_492,In_684);
nand U96 (N_96,In_129,In_1036);
and U97 (N_97,In_769,In_458);
nand U98 (N_98,In_1643,In_1405);
xnor U99 (N_99,In_1198,In_1266);
xnor U100 (N_100,In_1345,In_1938);
or U101 (N_101,In_304,In_857);
nor U102 (N_102,In_1540,In_153);
xor U103 (N_103,In_176,In_1300);
xor U104 (N_104,In_646,In_540);
xor U105 (N_105,In_745,In_1380);
nor U106 (N_106,In_1896,In_472);
nor U107 (N_107,In_1235,In_78);
and U108 (N_108,In_385,In_1450);
and U109 (N_109,In_56,In_668);
and U110 (N_110,In_314,In_791);
xnor U111 (N_111,In_1188,In_858);
xor U112 (N_112,In_1412,In_1952);
and U113 (N_113,In_400,In_1511);
nand U114 (N_114,In_1099,In_13);
and U115 (N_115,In_150,In_671);
xor U116 (N_116,In_1489,In_479);
nand U117 (N_117,In_21,In_772);
and U118 (N_118,In_60,In_149);
nor U119 (N_119,In_1022,In_898);
nand U120 (N_120,In_1012,In_1806);
or U121 (N_121,In_1937,In_801);
or U122 (N_122,In_1057,In_1370);
nor U123 (N_123,In_485,In_1975);
xnor U124 (N_124,In_905,In_636);
or U125 (N_125,In_907,In_152);
nor U126 (N_126,In_1157,In_313);
and U127 (N_127,In_1956,In_137);
and U128 (N_128,In_1576,In_1950);
xnor U129 (N_129,In_1869,In_296);
nand U130 (N_130,In_1843,In_510);
xnor U131 (N_131,In_1798,In_1379);
nand U132 (N_132,In_934,In_903);
xnor U133 (N_133,In_522,In_79);
nor U134 (N_134,In_1356,In_269);
xnor U135 (N_135,In_711,In_568);
xnor U136 (N_136,In_979,In_1026);
xnor U137 (N_137,In_1998,In_1908);
and U138 (N_138,In_716,In_1581);
xor U139 (N_139,In_93,In_327);
or U140 (N_140,In_1494,In_10);
nand U141 (N_141,In_651,In_1621);
and U142 (N_142,In_1897,In_1597);
nand U143 (N_143,In_1485,In_1163);
and U144 (N_144,In_1327,In_1019);
or U145 (N_145,In_975,In_1176);
nand U146 (N_146,In_930,In_1210);
nor U147 (N_147,In_208,In_1982);
and U148 (N_148,In_1475,In_451);
xor U149 (N_149,In_733,In_554);
nor U150 (N_150,In_1808,In_1676);
or U151 (N_151,In_1917,In_953);
and U152 (N_152,In_1290,In_478);
and U153 (N_153,In_1878,In_1219);
nor U154 (N_154,In_167,In_1109);
xor U155 (N_155,In_65,In_1134);
nand U156 (N_156,In_1717,In_133);
or U157 (N_157,In_1608,In_1005);
or U158 (N_158,In_1654,In_970);
xnor U159 (N_159,In_1941,In_614);
xor U160 (N_160,In_1342,In_1498);
nor U161 (N_161,In_1616,In_1394);
or U162 (N_162,In_379,In_1894);
or U163 (N_163,In_1243,In_1764);
or U164 (N_164,In_306,In_1545);
and U165 (N_165,In_899,In_1140);
nor U166 (N_166,In_871,In_843);
xor U167 (N_167,In_1725,In_559);
nand U168 (N_168,In_1501,In_1461);
or U169 (N_169,In_523,In_592);
xnor U170 (N_170,In_1490,In_447);
or U171 (N_171,In_565,In_186);
nor U172 (N_172,In_25,In_556);
and U173 (N_173,In_323,In_1864);
nor U174 (N_174,In_641,In_18);
nor U175 (N_175,In_1840,In_1382);
xnor U176 (N_176,In_1557,In_1192);
nand U177 (N_177,In_864,In_1914);
xnor U178 (N_178,In_874,In_1530);
nor U179 (N_179,In_581,In_6);
nor U180 (N_180,In_188,In_276);
xor U181 (N_181,In_625,In_1775);
xor U182 (N_182,In_1063,In_156);
or U183 (N_183,In_1733,In_1431);
and U184 (N_184,In_1754,In_834);
or U185 (N_185,In_1034,In_561);
xor U186 (N_186,In_1990,In_1680);
and U187 (N_187,In_960,In_748);
xnor U188 (N_188,In_1968,In_1169);
or U189 (N_189,In_812,In_359);
nand U190 (N_190,In_807,In_1100);
and U191 (N_191,In_1297,In_823);
nand U192 (N_192,In_928,In_1527);
or U193 (N_193,In_344,In_1730);
and U194 (N_194,In_612,In_294);
nand U195 (N_195,In_760,In_825);
xor U196 (N_196,In_55,In_1193);
or U197 (N_197,In_1008,In_566);
xnor U198 (N_198,In_289,In_1442);
xor U199 (N_199,In_301,In_1197);
nor U200 (N_200,In_1055,In_36);
and U201 (N_201,In_818,In_1276);
xor U202 (N_202,In_1948,In_1391);
nor U203 (N_203,In_544,In_1122);
xnor U204 (N_204,In_1301,In_1578);
xor U205 (N_205,In_1889,In_1999);
nor U206 (N_206,In_244,In_1575);
xor U207 (N_207,In_971,In_525);
xnor U208 (N_208,In_520,In_1518);
or U209 (N_209,In_530,In_15);
xor U210 (N_210,In_12,In_873);
nor U211 (N_211,In_1129,In_1570);
or U212 (N_212,In_58,In_991);
xnor U213 (N_213,In_225,In_1905);
xnor U214 (N_214,In_312,In_282);
or U215 (N_215,In_1334,In_1859);
nand U216 (N_216,In_1600,In_1164);
xnor U217 (N_217,In_981,In_141);
nand U218 (N_218,In_914,In_1305);
and U219 (N_219,In_1086,In_923);
xor U220 (N_220,In_318,In_120);
nor U221 (N_221,In_703,In_1462);
nor U222 (N_222,In_742,In_175);
xor U223 (N_223,In_594,In_1996);
or U224 (N_224,In_1907,In_1051);
nand U225 (N_225,In_1115,In_1316);
xor U226 (N_226,In_774,In_115);
or U227 (N_227,In_666,In_257);
nor U228 (N_228,In_66,In_701);
xor U229 (N_229,In_285,In_1747);
and U230 (N_230,In_1162,In_1625);
nor U231 (N_231,In_280,In_386);
xor U232 (N_232,In_528,In_669);
nor U233 (N_233,In_1817,In_1871);
nor U234 (N_234,In_1313,In_1963);
xor U235 (N_235,In_1230,In_1773);
nor U236 (N_236,In_14,In_1136);
or U237 (N_237,In_1403,In_255);
xnor U238 (N_238,In_1337,In_964);
nand U239 (N_239,In_396,In_597);
nand U240 (N_240,In_1944,In_1220);
nand U241 (N_241,In_219,In_1278);
nor U242 (N_242,In_246,In_1419);
nor U243 (N_243,In_810,In_1088);
or U244 (N_244,In_155,In_575);
nand U245 (N_245,In_1283,In_466);
nor U246 (N_246,In_1992,In_1205);
xnor U247 (N_247,In_746,In_200);
and U248 (N_248,In_75,In_1719);
or U249 (N_249,In_574,In_531);
nor U250 (N_250,In_1770,In_1177);
nor U251 (N_251,In_1378,In_1343);
nand U252 (N_252,In_849,In_1786);
nand U253 (N_253,In_869,In_1989);
and U254 (N_254,In_241,In_1383);
nand U255 (N_255,In_1879,In_853);
and U256 (N_256,In_1868,In_1656);
nand U257 (N_257,In_1174,In_1653);
and U258 (N_258,In_1911,In_1066);
nor U259 (N_259,In_394,In_613);
and U260 (N_260,In_1906,In_330);
nand U261 (N_261,In_495,In_793);
nor U262 (N_262,In_1801,In_602);
and U263 (N_263,In_171,In_128);
and U264 (N_264,In_117,In_1553);
or U265 (N_265,In_1799,In_982);
nand U266 (N_266,In_821,In_194);
and U267 (N_267,In_560,In_783);
or U268 (N_268,In_537,In_1712);
nor U269 (N_269,In_254,In_1111);
and U270 (N_270,In_1244,In_974);
or U271 (N_271,In_707,In_1354);
nor U272 (N_272,In_1838,In_1682);
nand U273 (N_273,In_1504,In_1274);
and U274 (N_274,In_1438,In_82);
nor U275 (N_275,In_183,In_62);
nor U276 (N_276,In_692,In_570);
nor U277 (N_277,In_406,In_1705);
xor U278 (N_278,In_8,In_190);
and U279 (N_279,In_139,In_1614);
nand U280 (N_280,In_513,In_392);
xor U281 (N_281,In_778,In_218);
nand U282 (N_282,In_1797,In_300);
nand U283 (N_283,In_1454,In_1409);
nor U284 (N_284,In_697,In_939);
or U285 (N_285,In_177,In_1374);
nor U286 (N_286,In_1264,In_918);
or U287 (N_287,In_1726,In_1030);
xnor U288 (N_288,In_259,In_1510);
and U289 (N_289,In_233,In_1254);
xnor U290 (N_290,In_123,In_28);
nor U291 (N_291,In_99,In_474);
nand U292 (N_292,In_937,In_1202);
nor U293 (N_293,In_395,In_1662);
and U294 (N_294,In_1738,In_1500);
or U295 (N_295,In_1832,In_740);
and U296 (N_296,In_1548,In_885);
xor U297 (N_297,In_500,In_1913);
nand U298 (N_298,In_985,In_1784);
and U299 (N_299,In_1150,In_681);
or U300 (N_300,In_929,In_172);
and U301 (N_301,In_865,In_146);
nor U302 (N_302,In_722,In_345);
nand U303 (N_303,In_680,In_1155);
nor U304 (N_304,In_1247,In_74);
nor U305 (N_305,In_1685,In_720);
nor U306 (N_306,In_1547,In_1401);
or U307 (N_307,In_1541,In_1520);
nor U308 (N_308,In_567,In_1605);
xnor U309 (N_309,In_1459,In_1309);
or U310 (N_310,In_499,In_1833);
or U311 (N_311,In_1571,In_1821);
nor U312 (N_312,In_256,In_603);
nand U313 (N_313,In_794,In_1138);
nor U314 (N_314,In_1127,In_332);
nand U315 (N_315,In_1018,In_1287);
xor U316 (N_316,In_1302,In_1335);
nand U317 (N_317,In_1167,In_940);
nand U318 (N_318,In_1376,In_890);
and U319 (N_319,In_1116,In_508);
nor U320 (N_320,In_855,In_1281);
nand U321 (N_321,In_1723,In_1559);
and U322 (N_322,In_1550,In_377);
nor U323 (N_323,In_1208,In_1488);
xor U324 (N_324,In_1315,In_712);
or U325 (N_325,In_585,In_768);
nand U326 (N_326,In_295,In_1890);
xor U327 (N_327,In_1692,In_1103);
and U328 (N_328,In_992,In_168);
nor U329 (N_329,In_1620,In_755);
xnor U330 (N_330,In_1729,In_1273);
xor U331 (N_331,In_211,In_1361);
xor U332 (N_332,In_1629,In_1895);
nand U333 (N_333,In_983,In_192);
and U334 (N_334,In_1828,In_328);
nand U335 (N_335,In_493,In_1007);
nand U336 (N_336,In_1515,In_416);
or U337 (N_337,In_162,In_767);
nor U338 (N_338,In_496,In_990);
nor U339 (N_339,In_846,In_1152);
and U340 (N_340,In_270,In_752);
xnor U341 (N_341,In_1533,In_904);
nor U342 (N_342,In_376,In_968);
and U343 (N_343,In_840,In_112);
xor U344 (N_344,In_677,In_1736);
and U345 (N_345,In_1678,In_580);
nand U346 (N_346,In_1299,In_632);
nand U347 (N_347,In_418,In_770);
nand U348 (N_348,In_1118,In_1027);
nand U349 (N_349,In_1146,In_1420);
or U350 (N_350,In_688,In_999);
or U351 (N_351,In_665,In_57);
nand U352 (N_352,In_1032,In_107);
nand U353 (N_353,In_1695,In_1710);
nand U354 (N_354,In_1104,In_7);
and U355 (N_355,In_956,In_324);
nor U356 (N_356,In_1194,In_1318);
or U357 (N_357,In_587,In_494);
and U358 (N_358,In_310,In_100);
xor U359 (N_359,In_886,In_1933);
or U360 (N_360,In_1482,In_702);
nand U361 (N_361,In_1644,In_1661);
nand U362 (N_362,In_976,In_813);
or U363 (N_363,In_773,In_110);
and U364 (N_364,In_1953,In_1265);
or U365 (N_365,In_1870,In_98);
nor U366 (N_366,In_1922,In_221);
nor U367 (N_367,In_611,In_1977);
and U368 (N_368,In_1788,In_1250);
or U369 (N_369,In_445,In_338);
nand U370 (N_370,In_88,In_430);
nor U371 (N_371,In_1528,In_1204);
nor U372 (N_372,In_572,In_1269);
nand U373 (N_373,In_1002,In_776);
nand U374 (N_374,In_1958,In_1633);
nand U375 (N_375,In_884,In_817);
xor U376 (N_376,In_122,In_1093);
xnor U377 (N_377,In_1288,In_1985);
xor U378 (N_378,In_467,In_215);
or U379 (N_379,In_827,In_1160);
or U380 (N_380,In_1826,In_739);
nor U381 (N_381,In_1293,In_1915);
nor U382 (N_382,In_624,In_1964);
nand U383 (N_383,In_135,In_1955);
or U384 (N_384,In_42,In_1844);
xor U385 (N_385,In_213,In_558);
nand U386 (N_386,In_471,In_440);
nand U387 (N_387,In_1505,In_675);
nor U388 (N_388,In_1009,In_1767);
xnor U389 (N_389,In_1499,In_19);
xor U390 (N_390,In_1829,In_199);
xor U391 (N_391,In_815,In_1404);
and U392 (N_392,In_286,In_958);
nand U393 (N_393,In_1873,In_1037);
nand U394 (N_394,In_1039,In_238);
and U395 (N_395,In_831,In_1753);
or U396 (N_396,In_650,In_1159);
nor U397 (N_397,In_1624,In_719);
nand U398 (N_398,In_1769,In_1408);
nand U399 (N_399,In_879,In_240);
nand U400 (N_400,In_329,In_920);
and U401 (N_401,In_1227,In_456);
and U402 (N_402,In_1465,In_571);
nand U403 (N_403,In_652,In_388);
nor U404 (N_404,In_657,In_868);
and U405 (N_405,In_973,In_1024);
or U406 (N_406,In_134,In_357);
or U407 (N_407,In_548,In_1761);
nand U408 (N_408,In_114,In_737);
xnor U409 (N_409,In_1735,In_833);
and U410 (N_410,In_891,In_163);
and U411 (N_411,In_1367,In_105);
xor U412 (N_412,In_1886,In_1232);
and U413 (N_413,In_1790,In_1961);
xor U414 (N_414,In_505,In_766);
or U415 (N_415,In_919,In_1377);
and U416 (N_416,In_399,In_1183);
or U417 (N_417,In_1195,In_197);
and U418 (N_418,In_488,In_1453);
nand U419 (N_419,In_448,In_526);
or U420 (N_420,In_434,In_1285);
nor U421 (N_421,In_1529,In_631);
and U422 (N_422,In_1071,In_1349);
or U423 (N_423,In_1268,In_1481);
xnor U424 (N_424,In_380,In_1017);
or U425 (N_425,In_1166,In_1517);
nor U426 (N_426,In_1704,In_308);
or U427 (N_427,In_384,In_901);
and U428 (N_428,In_387,In_1415);
xor U429 (N_429,In_1237,In_305);
and U430 (N_430,In_459,In_1090);
and U431 (N_431,In_1672,In_1813);
xor U432 (N_432,In_84,In_1901);
nor U433 (N_433,In_354,In_693);
xor U434 (N_434,In_848,In_109);
nor U435 (N_435,In_909,In_1267);
xor U436 (N_436,In_1410,In_1406);
nand U437 (N_437,In_427,In_311);
nor U438 (N_438,In_785,In_1561);
xor U439 (N_439,In_1569,In_368);
nand U440 (N_440,In_161,In_1011);
or U441 (N_441,In_1231,In_1411);
or U442 (N_442,In_1749,In_1674);
nor U443 (N_443,In_1314,In_203);
nor U444 (N_444,In_1807,In_1688);
nand U445 (N_445,In_1523,In_1471);
nand U446 (N_446,In_220,In_1647);
or U447 (N_447,In_1137,In_779);
nand U448 (N_448,In_235,In_1279);
xor U449 (N_449,In_337,In_31);
nand U450 (N_450,In_1945,In_428);
nand U451 (N_451,In_867,In_1135);
nand U452 (N_452,In_1659,In_46);
nand U453 (N_453,In_1242,In_293);
nand U454 (N_454,In_789,In_464);
xor U455 (N_455,In_1147,In_924);
and U456 (N_456,In_127,In_482);
nor U457 (N_457,In_598,In_364);
and U458 (N_458,In_452,In_1655);
xnor U459 (N_459,In_378,In_617);
xor U460 (N_460,In_1815,In_423);
and U461 (N_461,In_1509,In_360);
and U462 (N_462,In_619,In_373);
or U463 (N_463,In_1699,In_1339);
or U464 (N_464,In_1585,In_1493);
xor U465 (N_465,In_935,In_227);
nor U466 (N_466,In_1675,In_1721);
and U467 (N_467,In_965,In_616);
xnor U468 (N_468,In_851,In_621);
or U469 (N_469,In_145,In_577);
or U470 (N_470,In_1046,In_1839);
nor U471 (N_471,In_1827,In_1209);
nand U472 (N_472,In_81,In_1782);
and U473 (N_473,In_1363,In_1497);
nand U474 (N_474,In_95,In_638);
nor U475 (N_475,In_591,In_1246);
nor U476 (N_476,In_350,In_1308);
xor U477 (N_477,In_1218,In_1632);
and U478 (N_478,In_1087,In_144);
nor U479 (N_479,In_1123,In_1084);
and U480 (N_480,In_1765,In_894);
or U481 (N_481,In_1919,In_759);
and U482 (N_482,In_1151,In_1755);
xnor U483 (N_483,In_435,In_389);
xnor U484 (N_484,In_1325,In_229);
or U485 (N_485,In_714,In_1669);
nor U486 (N_486,In_1618,In_1702);
and U487 (N_487,In_1094,In_1731);
nor U488 (N_488,In_158,In_734);
nor U489 (N_489,In_1664,In_1590);
nand U490 (N_490,In_1554,In_1207);
nor U491 (N_491,In_397,In_541);
nor U492 (N_492,In_866,In_361);
or U493 (N_493,In_989,In_268);
and U494 (N_494,In_841,In_1718);
or U495 (N_495,In_1000,In_1263);
or U496 (N_496,In_1607,In_1417);
and U497 (N_497,In_1872,In_191);
or U498 (N_498,In_1543,In_842);
nor U499 (N_499,In_555,In_1366);
xnor U500 (N_500,In_835,In_1638);
and U501 (N_501,In_1074,In_316);
xnor U502 (N_502,In_491,In_538);
or U503 (N_503,In_800,In_1424);
nand U504 (N_504,In_444,In_729);
nand U505 (N_505,In_358,In_398);
nor U506 (N_506,In_1965,In_1693);
or U507 (N_507,In_1038,In_212);
nor U508 (N_508,In_1789,In_271);
and U509 (N_509,In_1877,In_623);
and U510 (N_510,In_601,In_1577);
and U511 (N_511,In_1903,In_1631);
and U512 (N_512,In_1847,In_23);
nand U513 (N_513,In_1525,In_888);
or U514 (N_514,In_1270,In_805);
or U515 (N_515,In_1830,In_828);
or U516 (N_516,In_1289,In_932);
xor U517 (N_517,In_1317,In_1058);
nor U518 (N_518,In_20,In_994);
xor U519 (N_519,In_1874,In_696);
xor U520 (N_520,In_189,In_1035);
or U521 (N_521,In_1800,In_1082);
nor U522 (N_522,In_374,In_507);
nor U523 (N_523,In_980,In_381);
nor U524 (N_524,In_86,In_708);
and U525 (N_525,In_1259,In_454);
nor U526 (N_526,In_947,In_1935);
or U527 (N_527,In_551,In_519);
xor U528 (N_528,In_988,In_160);
xnor U529 (N_529,In_948,In_1443);
xor U530 (N_530,In_1199,In_727);
or U531 (N_531,In_169,In_1114);
nand U532 (N_532,In_1402,In_1856);
and U533 (N_533,In_942,In_881);
and U534 (N_534,In_1651,In_1592);
nand U535 (N_535,In_249,In_274);
and U536 (N_536,In_1572,In_1951);
nor U537 (N_537,In_690,In_620);
and U538 (N_538,In_775,In_736);
or U539 (N_539,In_1857,In_1783);
xor U540 (N_540,In_1696,In_809);
nand U541 (N_541,In_1003,In_1924);
and U542 (N_542,In_512,In_1564);
nor U543 (N_543,In_1816,In_73);
or U544 (N_544,In_1286,In_1061);
or U545 (N_545,In_781,In_685);
nand U546 (N_546,In_1480,In_1330);
nand U547 (N_547,In_844,In_1056);
nand U548 (N_548,In_615,In_670);
nand U549 (N_549,In_422,In_824);
nor U550 (N_550,In_1429,In_1203);
or U551 (N_551,In_1414,In_1640);
and U552 (N_552,In_382,In_383);
xor U553 (N_553,In_1430,In_1421);
or U554 (N_554,In_1526,In_725);
xor U555 (N_555,In_546,In_1125);
xor U556 (N_556,In_1671,In_353);
nor U557 (N_557,In_1850,In_411);
or U558 (N_558,In_322,In_298);
nand U559 (N_559,In_1449,In_761);
and U560 (N_560,In_210,In_292);
and U561 (N_561,In_1762,In_1389);
and U562 (N_562,In_1092,In_1029);
nor U563 (N_563,In_465,In_1954);
or U564 (N_564,In_626,In_1170);
xnor U565 (N_565,In_1440,In_967);
and U566 (N_566,In_369,In_1399);
nor U567 (N_567,In_1930,In_1187);
or U568 (N_568,In_1455,In_237);
nor U569 (N_569,In_576,In_1984);
nor U570 (N_570,In_1739,In_438);
nor U571 (N_571,In_302,In_563);
xor U572 (N_572,In_80,In_39);
nor U573 (N_573,In_877,In_103);
or U574 (N_574,In_1552,In_706);
nand U575 (N_575,In_777,In_1364);
xor U576 (N_576,In_1225,In_130);
nor U577 (N_577,In_1885,In_1168);
nand U578 (N_578,In_814,In_1179);
and U579 (N_579,In_366,In_198);
nand U580 (N_580,In_600,In_33);
or U581 (N_581,In_1425,In_1447);
and U582 (N_582,In_490,In_957);
xor U583 (N_583,In_291,In_1025);
nor U584 (N_584,In_441,In_1771);
nand U585 (N_585,In_288,In_250);
or U586 (N_586,In_1967,In_1534);
and U587 (N_587,In_22,In_524);
nand U588 (N_588,In_346,In_393);
or U589 (N_589,In_1373,In_1387);
nor U590 (N_590,In_686,In_1974);
nand U591 (N_591,In_365,In_763);
nor U592 (N_592,In_1506,In_258);
nor U593 (N_593,In_1422,In_232);
or U594 (N_594,In_253,In_1503);
xnor U595 (N_595,In_1627,In_209);
nor U596 (N_596,In_1213,In_1602);
nor U597 (N_597,In_1139,In_1929);
xor U598 (N_598,In_687,In_1196);
or U599 (N_599,In_202,In_1298);
nor U600 (N_600,In_412,In_1665);
xnor U601 (N_601,In_806,In_367);
nor U602 (N_602,In_889,In_1740);
nand U603 (N_603,In_1102,In_439);
nand U604 (N_604,In_506,In_977);
xor U605 (N_605,In_1745,In_90);
xnor U606 (N_606,In_1001,In_532);
nand U607 (N_607,In_966,In_897);
or U608 (N_608,In_1787,In_1040);
and U609 (N_609,In_267,In_281);
or U610 (N_610,In_1120,In_829);
xnor U611 (N_611,In_1312,In_1161);
or U612 (N_612,In_1812,In_786);
or U613 (N_613,In_234,In_1398);
or U614 (N_614,In_1158,In_820);
and U615 (N_615,In_870,In_1);
xnor U616 (N_616,In_1333,In_343);
or U617 (N_617,In_754,In_1531);
xor U618 (N_618,In_511,In_1226);
xor U619 (N_619,In_1720,In_1727);
or U620 (N_620,In_1825,In_1479);
nand U621 (N_621,In_1329,In_151);
and U622 (N_622,In_193,In_96);
nor U623 (N_623,In_315,In_502);
nand U624 (N_624,In_1310,In_1648);
xnor U625 (N_625,In_1772,In_1081);
nor U626 (N_626,In_303,In_462);
xor U627 (N_627,In_1460,In_1660);
xor U628 (N_628,In_1882,In_11);
xnor U629 (N_629,In_266,In_1458);
xnor U630 (N_630,In_351,In_573);
or U631 (N_631,In_863,In_1900);
or U632 (N_632,In_278,In_658);
and U633 (N_633,In_339,In_475);
nor U634 (N_634,In_424,In_340);
or U635 (N_635,In_290,In_916);
or U636 (N_636,In_1960,In_1666);
nor U637 (N_637,In_993,In_880);
nor U638 (N_638,In_644,In_5);
or U639 (N_639,In_16,In_1080);
nor U640 (N_640,In_1400,In_1248);
xor U641 (N_641,In_1048,In_950);
nor U642 (N_642,In_749,In_1697);
nor U643 (N_643,In_705,In_432);
or U644 (N_644,In_1606,In_893);
or U645 (N_645,In_1623,In_1491);
xnor U646 (N_646,In_1583,In_1062);
and U647 (N_647,In_1617,In_181);
xor U648 (N_648,In_371,In_1677);
or U649 (N_649,In_32,In_148);
or U650 (N_650,In_1171,In_902);
nand U651 (N_651,In_896,In_963);
nand U652 (N_652,In_195,In_1645);
nand U653 (N_653,In_593,In_765);
or U654 (N_654,In_347,In_1637);
xnor U655 (N_655,In_1514,In_1639);
or U656 (N_656,In_1441,In_457);
or U657 (N_657,In_1369,In_514);
and U658 (N_658,In_217,In_1047);
xnor U659 (N_659,In_297,In_1707);
or U660 (N_660,In_1658,In_584);
or U661 (N_661,In_1836,In_1888);
and U662 (N_662,In_1698,In_390);
nand U663 (N_663,In_1760,In_449);
xor U664 (N_664,In_978,In_1701);
and U665 (N_665,In_1743,In_1918);
or U666 (N_666,In_299,In_1296);
or U667 (N_667,In_355,In_1184);
nor U668 (N_668,In_179,In_1180);
xnor U669 (N_669,In_1538,In_926);
nor U670 (N_670,In_1588,In_375);
xor U671 (N_671,In_1272,In_732);
nand U672 (N_672,In_70,In_1646);
nand U673 (N_673,In_104,In_1595);
nor U674 (N_674,In_1206,In_1307);
nor U675 (N_675,In_1741,In_1126);
nand U676 (N_676,In_622,In_1340);
nor U677 (N_677,In_1635,In_317);
xnor U678 (N_678,In_1256,In_1835);
or U679 (N_679,In_1439,In_943);
or U680 (N_680,In_672,In_1464);
nand U681 (N_681,In_216,In_1634);
xor U682 (N_682,In_341,In_1041);
or U683 (N_683,In_159,In_521);
xnor U684 (N_684,In_1642,In_1448);
nand U685 (N_685,In_463,In_944);
or U686 (N_686,In_1346,In_1033);
xor U687 (N_687,In_995,In_1778);
nor U688 (N_688,In_437,In_319);
or U689 (N_689,In_187,In_875);
nand U690 (N_690,In_436,In_882);
nand U691 (N_691,In_1796,In_1463);
nor U692 (N_692,In_92,In_539);
and U693 (N_693,In_1072,In_1758);
xor U694 (N_694,In_503,In_1436);
or U695 (N_695,In_1524,In_1802);
and U696 (N_696,In_683,In_588);
nand U697 (N_697,In_1622,In_30);
nor U698 (N_698,In_1323,In_44);
and U699 (N_699,In_1536,In_583);
or U700 (N_700,In_1611,In_1587);
nand U701 (N_701,In_1854,In_140);
or U702 (N_702,In_1015,In_1819);
nand U703 (N_703,In_1820,In_1486);
nand U704 (N_704,In_1936,In_1516);
nor U705 (N_705,In_1916,In_450);
nor U706 (N_706,In_1028,In_1910);
nor U707 (N_707,In_275,In_872);
xor U708 (N_708,In_1234,In_1943);
xnor U709 (N_709,In_231,In_1252);
xor U710 (N_710,In_1306,In_402);
or U711 (N_711,In_1236,In_628);
or U712 (N_712,In_1108,In_921);
xnor U713 (N_713,In_895,In_1089);
or U714 (N_714,In_845,In_1070);
or U715 (N_715,In_649,In_878);
nand U716 (N_716,In_372,In_1703);
xnor U717 (N_717,In_718,In_483);
and U718 (N_718,In_184,In_77);
and U719 (N_719,In_799,In_1013);
xor U720 (N_720,In_1714,In_124);
nor U721 (N_721,In_207,In_1995);
xnor U722 (N_722,In_1931,In_1049);
and U723 (N_723,In_166,In_413);
and U724 (N_724,In_1484,In_1940);
nor U725 (N_725,In_1386,In_1861);
nor U726 (N_726,In_961,In_656);
and U727 (N_727,In_1434,In_1076);
or U728 (N_728,In_1154,In_910);
xnor U729 (N_729,In_1221,In_721);
and U730 (N_730,In_425,In_1841);
nand U731 (N_731,In_1393,In_157);
nand U732 (N_732,In_1932,In_629);
or U733 (N_733,In_1432,In_71);
xor U734 (N_734,In_1988,In_582);
or U735 (N_735,In_91,In_1347);
xor U736 (N_736,In_1451,In_1119);
xnor U737 (N_737,In_1978,In_1887);
and U738 (N_738,In_1846,In_1487);
or U739 (N_739,In_1078,In_1909);
or U740 (N_740,In_1130,In_1980);
xnor U741 (N_741,In_860,In_1238);
and U742 (N_742,In_247,In_480);
nor U743 (N_743,In_1470,In_142);
or U744 (N_744,In_1322,In_1331);
nor U745 (N_745,In_1344,In_1779);
and U746 (N_746,In_461,In_1502);
or U747 (N_747,In_1113,In_433);
or U748 (N_748,In_484,In_1742);
nand U749 (N_749,In_1694,In_1277);
or U750 (N_750,In_1805,In_1558);
xnor U751 (N_751,In_797,In_1275);
nand U752 (N_752,In_1997,In_49);
or U753 (N_753,In_273,In_1756);
nor U754 (N_754,In_1862,In_1469);
nor U755 (N_755,In_501,In_67);
or U756 (N_756,In_1876,In_803);
or U757 (N_757,In_1891,In_41);
nor U758 (N_758,In_1368,In_415);
nor U759 (N_759,In_1437,In_1512);
and U760 (N_760,In_1513,In_1390);
nand U761 (N_761,In_633,In_1809);
or U762 (N_762,In_986,In_1939);
nand U763 (N_763,In_782,In_1075);
or U764 (N_764,In_1681,In_1928);
or U765 (N_765,In_1239,In_946);
and U766 (N_766,In_642,In_1045);
or U767 (N_767,In_536,In_1172);
nand U768 (N_768,In_1365,In_726);
xnor U769 (N_769,In_262,In_1468);
xor U770 (N_770,In_557,In_1261);
xnor U771 (N_771,In_709,In_699);
or U772 (N_772,In_1649,In_792);
nor U773 (N_773,In_2,In_579);
nor U774 (N_774,In_1190,In_941);
or U775 (N_775,In_1567,In_277);
xnor U776 (N_776,In_1145,In_756);
and U777 (N_777,In_1708,In_1352);
nand U778 (N_778,In_1141,In_1212);
xnor U779 (N_779,In_272,In_1085);
and U780 (N_780,In_1792,In_476);
nand U781 (N_781,In_998,In_1295);
xnor U782 (N_782,In_409,In_1811);
or U783 (N_783,In_1927,In_1892);
nor U784 (N_784,In_854,In_728);
xnor U785 (N_785,In_839,In_356);
and U786 (N_786,In_43,In_1686);
nor U787 (N_787,In_1211,In_917);
nand U788 (N_788,In_1044,In_911);
xnor U789 (N_789,In_1628,In_469);
and U790 (N_790,In_125,In_1251);
nand U791 (N_791,In_1589,In_659);
xor U792 (N_792,In_682,In_1381);
or U793 (N_793,In_119,In_248);
or U794 (N_794,In_53,In_429);
nand U795 (N_795,In_1630,In_710);
and U796 (N_796,In_1546,In_1875);
and U797 (N_797,In_1848,In_1328);
or U798 (N_798,In_674,In_850);
xnor U799 (N_799,In_1986,In_29);
nor U800 (N_800,In_1360,In_1069);
nor U801 (N_801,In_599,In_348);
nand U802 (N_802,In_922,In_1496);
and U803 (N_803,In_121,In_590);
nor U804 (N_804,In_1031,In_927);
xnor U805 (N_805,In_730,In_116);
nor U806 (N_806,In_1668,In_552);
xnor U807 (N_807,In_1966,In_333);
or U808 (N_808,In_1215,In_180);
nand U809 (N_809,In_1724,In_1427);
xor U810 (N_810,In_1396,In_1542);
and U811 (N_811,In_1474,In_1987);
xnor U812 (N_812,In_1535,In_473);
and U813 (N_813,In_704,In_1385);
nor U814 (N_814,In_859,In_1748);
nor U815 (N_815,In_50,In_1191);
or U816 (N_816,In_569,In_861);
xnor U817 (N_817,In_68,In_758);
xor U818 (N_818,In_1372,In_118);
and U819 (N_819,In_915,In_334);
xor U820 (N_820,In_89,In_798);
nand U821 (N_821,In_1182,In_201);
or U822 (N_822,In_101,In_1214);
xor U823 (N_823,In_326,In_251);
or U824 (N_824,In_640,In_1353);
nor U825 (N_825,In_223,In_1979);
xnor U826 (N_826,In_790,In_1562);
xor U827 (N_827,In_477,In_1101);
or U828 (N_828,In_1609,In_1713);
nand U829 (N_829,In_1319,In_245);
nand U830 (N_830,In_486,In_48);
nor U831 (N_831,In_1912,In_1582);
xor U832 (N_832,In_1338,In_1476);
nand U833 (N_833,In_996,In_1687);
nor U834 (N_834,In_795,In_533);
and U835 (N_835,In_1842,In_1359);
nand U836 (N_836,In_284,In_936);
and U837 (N_837,In_647,In_1294);
and U838 (N_838,In_205,In_527);
and U839 (N_839,In_1133,In_349);
or U840 (N_840,In_1228,In_1641);
nand U841 (N_841,In_59,In_1357);
or U842 (N_842,In_403,In_1407);
and U843 (N_843,In_771,In_1994);
or U844 (N_844,In_1073,In_38);
and U845 (N_845,In_419,In_1418);
or U846 (N_846,In_635,In_1457);
xor U847 (N_847,In_634,In_1477);
nand U848 (N_848,In_1690,In_414);
and U849 (N_849,In_206,In_69);
nand U850 (N_850,In_1594,In_1934);
and U851 (N_851,In_335,In_1573);
and U852 (N_852,In_1216,In_1768);
and U853 (N_853,In_1433,In_1706);
nor U854 (N_854,In_637,In_1110);
nand U855 (N_855,In_1128,In_1124);
or U856 (N_856,In_331,In_283);
nand U857 (N_857,In_252,In_1131);
xor U858 (N_858,In_242,In_446);
xnor U859 (N_859,In_1253,In_1106);
or U860 (N_860,In_287,In_1926);
nor U861 (N_861,In_955,In_673);
nand U862 (N_862,In_1893,In_1117);
and U863 (N_863,In_352,In_892);
xor U864 (N_864,In_1711,In_1853);
nand U865 (N_865,In_1043,In_1804);
nor U866 (N_866,In_1532,In_487);
and U867 (N_867,In_856,In_1962);
nand U868 (N_868,In_417,In_1810);
xnor U869 (N_869,In_481,In_1774);
or U870 (N_870,In_578,In_497);
xnor U871 (N_871,In_1763,In_951);
and U872 (N_872,In_228,In_1636);
nand U873 (N_873,In_1185,In_816);
xnor U874 (N_874,In_1291,In_1059);
nand U875 (N_875,In_1780,In_648);
xnor U876 (N_876,In_662,In_1112);
nor U877 (N_877,In_236,In_106);
or U878 (N_878,In_847,In_9);
nand U879 (N_879,In_678,In_170);
xnor U880 (N_880,In_410,In_1603);
xnor U881 (N_881,In_962,In_3);
nor U882 (N_882,In_925,In_1593);
nor U883 (N_883,In_1042,In_362);
nand U884 (N_884,In_1746,In_239);
and U885 (N_885,In_1904,In_630);
or U886 (N_886,In_876,In_1292);
xnor U887 (N_887,In_1599,In_1004);
or U888 (N_888,In_1006,In_550);
and U889 (N_889,In_1852,In_321);
xnor U890 (N_890,In_912,In_174);
or U891 (N_891,In_1282,In_987);
nand U892 (N_892,In_1060,In_836);
nor U893 (N_893,In_515,In_1855);
nand U894 (N_894,In_1981,In_1508);
nor U895 (N_895,In_131,In_126);
and U896 (N_896,In_1679,In_908);
xor U897 (N_897,In_731,In_1777);
nor U898 (N_898,In_717,In_1750);
xor U899 (N_899,In_738,In_1667);
xor U900 (N_900,In_743,In_1023);
xor U901 (N_901,In_1959,In_1223);
xor U902 (N_902,In_518,In_1284);
or U903 (N_903,In_173,In_1426);
and U904 (N_904,In_26,In_837);
nor U905 (N_905,In_608,In_1814);
and U906 (N_906,In_1849,In_1271);
or U907 (N_907,In_906,In_1445);
nand U908 (N_908,In_154,In_1053);
xor U909 (N_909,In_404,In_342);
nand U910 (N_910,In_1375,In_1673);
nand U911 (N_911,In_1759,In_1728);
xnor U912 (N_912,In_1324,In_1240);
xor U913 (N_913,In_442,In_1863);
or U914 (N_914,In_498,In_811);
and U915 (N_915,In_984,In_862);
or U916 (N_916,In_1670,In_261);
or U917 (N_917,In_586,In_972);
and U918 (N_918,In_1976,In_1568);
nor U919 (N_919,In_1016,In_1303);
nor U920 (N_920,In_1860,In_1052);
and U921 (N_921,In_1899,In_1079);
and U922 (N_922,In_1260,In_113);
and U923 (N_923,In_516,In_735);
nand U924 (N_924,In_1142,In_1626);
or U925 (N_925,In_1866,In_1881);
or U926 (N_926,In_1803,In_1865);
or U927 (N_927,In_1350,In_164);
xnor U928 (N_928,In_1121,In_102);
nor U929 (N_929,In_1098,In_320);
nor U930 (N_930,In_260,In_1596);
nand U931 (N_931,In_0,In_1341);
nor U932 (N_932,In_969,In_700);
and U933 (N_933,In_1867,In_661);
nor U934 (N_934,In_1732,In_605);
xor U935 (N_935,In_1358,In_1565);
and U936 (N_936,In_85,In_1153);
and U937 (N_937,In_182,In_45);
and U938 (N_938,In_784,In_1831);
nor U939 (N_939,In_94,In_1612);
and U940 (N_940,In_52,In_1791);
nand U941 (N_941,In_796,In_1818);
nor U942 (N_942,In_4,In_1143);
nor U943 (N_943,In_788,In_1064);
nand U944 (N_944,In_1566,In_997);
nand U945 (N_945,In_1683,In_325);
nor U946 (N_946,In_787,In_655);
xnor U947 (N_947,In_1095,In_949);
nor U948 (N_948,In_664,In_83);
xor U949 (N_949,In_1413,In_1613);
nor U950 (N_950,In_1598,In_1601);
xnor U951 (N_951,In_370,In_1224);
nand U952 (N_952,In_1262,In_1946);
xor U953 (N_953,In_1619,In_954);
or U954 (N_954,In_564,In_1610);
nor U955 (N_955,In_643,In_757);
nor U956 (N_956,In_1355,In_1495);
xnor U957 (N_957,In_1555,In_1233);
or U958 (N_958,In_1615,In_279);
and U959 (N_959,In_1560,In_852);
and U960 (N_960,In_695,In_689);
or U961 (N_961,In_509,In_1065);
nor U962 (N_962,In_1304,In_1452);
and U963 (N_963,In_1715,In_51);
nor U964 (N_964,In_1326,In_204);
or U965 (N_965,In_589,In_1722);
and U966 (N_966,In_744,In_952);
nor U967 (N_967,In_1983,In_639);
nand U968 (N_968,In_553,In_1173);
nor U969 (N_969,In_1539,In_1492);
nor U970 (N_970,In_715,In_336);
and U971 (N_971,In_1362,In_945);
xnor U972 (N_972,In_363,In_653);
nand U973 (N_973,In_713,In_1993);
or U974 (N_974,In_1766,In_1472);
or U975 (N_975,In_147,In_830);
and U976 (N_976,In_1201,In_37);
nor U977 (N_977,In_694,In_542);
nand U978 (N_978,In_64,In_562);
nand U979 (N_979,In_35,In_1563);
nand U980 (N_980,In_1969,In_1107);
nand U981 (N_981,In_307,In_543);
xnor U982 (N_982,In_1428,In_1416);
xnor U983 (N_983,In_1144,In_534);
xor U984 (N_984,In_1752,In_196);
and U985 (N_985,In_1478,In_1970);
and U986 (N_986,In_1097,In_1795);
nand U987 (N_987,In_832,In_1522);
nand U988 (N_988,In_545,In_1972);
nand U989 (N_989,In_1684,In_1446);
and U990 (N_990,In_959,In_1077);
or U991 (N_991,In_143,In_679);
nand U992 (N_992,In_17,In_931);
nand U993 (N_993,In_1181,In_1105);
or U994 (N_994,In_1456,In_1822);
and U995 (N_995,In_108,In_1336);
xor U996 (N_996,In_804,In_421);
or U997 (N_997,In_1519,In_1371);
and U998 (N_998,In_1785,In_1332);
nand U999 (N_999,In_1186,In_420);
nand U1000 (N_1000,In_347,In_1575);
nor U1001 (N_1001,In_1655,In_1261);
nor U1002 (N_1002,In_8,In_501);
nor U1003 (N_1003,In_962,In_1871);
nor U1004 (N_1004,In_575,In_296);
nand U1005 (N_1005,In_13,In_1678);
nor U1006 (N_1006,In_147,In_1116);
xnor U1007 (N_1007,In_1860,In_1182);
and U1008 (N_1008,In_55,In_840);
nand U1009 (N_1009,In_1458,In_537);
nor U1010 (N_1010,In_703,In_1408);
and U1011 (N_1011,In_633,In_517);
and U1012 (N_1012,In_1973,In_154);
xor U1013 (N_1013,In_745,In_1234);
xnor U1014 (N_1014,In_1694,In_1196);
xnor U1015 (N_1015,In_1745,In_1270);
and U1016 (N_1016,In_1853,In_1790);
nand U1017 (N_1017,In_1912,In_1619);
xnor U1018 (N_1018,In_1041,In_611);
or U1019 (N_1019,In_246,In_461);
and U1020 (N_1020,In_1681,In_1002);
or U1021 (N_1021,In_459,In_1439);
nor U1022 (N_1022,In_178,In_326);
nor U1023 (N_1023,In_749,In_848);
xnor U1024 (N_1024,In_860,In_1808);
and U1025 (N_1025,In_886,In_268);
nor U1026 (N_1026,In_125,In_828);
and U1027 (N_1027,In_1346,In_745);
nand U1028 (N_1028,In_753,In_1624);
and U1029 (N_1029,In_574,In_1379);
xor U1030 (N_1030,In_722,In_1442);
or U1031 (N_1031,In_1457,In_744);
nor U1032 (N_1032,In_1876,In_2);
xnor U1033 (N_1033,In_923,In_841);
xnor U1034 (N_1034,In_991,In_114);
nor U1035 (N_1035,In_1852,In_1729);
and U1036 (N_1036,In_1195,In_1840);
nand U1037 (N_1037,In_1865,In_455);
or U1038 (N_1038,In_1187,In_493);
nand U1039 (N_1039,In_1137,In_1523);
nand U1040 (N_1040,In_1979,In_1928);
xor U1041 (N_1041,In_711,In_1452);
and U1042 (N_1042,In_1065,In_1716);
nor U1043 (N_1043,In_885,In_386);
or U1044 (N_1044,In_574,In_1360);
and U1045 (N_1045,In_1928,In_1698);
and U1046 (N_1046,In_883,In_288);
nand U1047 (N_1047,In_7,In_822);
xnor U1048 (N_1048,In_1185,In_711);
and U1049 (N_1049,In_47,In_1823);
and U1050 (N_1050,In_1921,In_1822);
xnor U1051 (N_1051,In_1608,In_1211);
nor U1052 (N_1052,In_1271,In_483);
nor U1053 (N_1053,In_57,In_1982);
nand U1054 (N_1054,In_423,In_677);
nand U1055 (N_1055,In_888,In_1403);
nor U1056 (N_1056,In_829,In_1594);
nand U1057 (N_1057,In_492,In_1531);
xnor U1058 (N_1058,In_46,In_188);
xnor U1059 (N_1059,In_1414,In_1396);
xnor U1060 (N_1060,In_1334,In_420);
and U1061 (N_1061,In_1068,In_1282);
and U1062 (N_1062,In_764,In_61);
nand U1063 (N_1063,In_1160,In_210);
nand U1064 (N_1064,In_836,In_1178);
nor U1065 (N_1065,In_1160,In_720);
and U1066 (N_1066,In_669,In_732);
nor U1067 (N_1067,In_1918,In_1670);
and U1068 (N_1068,In_1118,In_156);
and U1069 (N_1069,In_1494,In_377);
nor U1070 (N_1070,In_519,In_1193);
nand U1071 (N_1071,In_1828,In_1187);
nand U1072 (N_1072,In_350,In_828);
xnor U1073 (N_1073,In_1401,In_1202);
xnor U1074 (N_1074,In_906,In_398);
xor U1075 (N_1075,In_1617,In_1538);
nand U1076 (N_1076,In_1114,In_1017);
xnor U1077 (N_1077,In_915,In_1783);
or U1078 (N_1078,In_257,In_1375);
nor U1079 (N_1079,In_692,In_825);
nand U1080 (N_1080,In_745,In_1758);
xor U1081 (N_1081,In_1210,In_1017);
and U1082 (N_1082,In_669,In_1653);
nand U1083 (N_1083,In_308,In_1284);
xnor U1084 (N_1084,In_704,In_1420);
nor U1085 (N_1085,In_205,In_145);
nor U1086 (N_1086,In_1798,In_236);
and U1087 (N_1087,In_391,In_78);
or U1088 (N_1088,In_1631,In_1940);
nor U1089 (N_1089,In_1775,In_246);
nand U1090 (N_1090,In_264,In_205);
or U1091 (N_1091,In_1834,In_1227);
and U1092 (N_1092,In_1524,In_775);
nor U1093 (N_1093,In_1086,In_100);
nand U1094 (N_1094,In_1027,In_426);
xor U1095 (N_1095,In_248,In_1174);
and U1096 (N_1096,In_1943,In_1810);
nand U1097 (N_1097,In_1350,In_170);
xor U1098 (N_1098,In_1205,In_1183);
nand U1099 (N_1099,In_1914,In_184);
xnor U1100 (N_1100,In_1720,In_1402);
and U1101 (N_1101,In_506,In_1256);
or U1102 (N_1102,In_1266,In_1860);
xor U1103 (N_1103,In_1165,In_1952);
or U1104 (N_1104,In_974,In_1000);
and U1105 (N_1105,In_80,In_1201);
and U1106 (N_1106,In_1700,In_42);
xor U1107 (N_1107,In_1410,In_1799);
or U1108 (N_1108,In_1114,In_1649);
nand U1109 (N_1109,In_539,In_1660);
or U1110 (N_1110,In_1075,In_1232);
nor U1111 (N_1111,In_178,In_855);
and U1112 (N_1112,In_1939,In_819);
xor U1113 (N_1113,In_443,In_1538);
xor U1114 (N_1114,In_308,In_1598);
and U1115 (N_1115,In_369,In_1392);
or U1116 (N_1116,In_1946,In_1589);
and U1117 (N_1117,In_1479,In_1183);
xor U1118 (N_1118,In_1969,In_951);
nor U1119 (N_1119,In_142,In_294);
nor U1120 (N_1120,In_821,In_1062);
nor U1121 (N_1121,In_445,In_736);
or U1122 (N_1122,In_1904,In_1306);
and U1123 (N_1123,In_907,In_1581);
or U1124 (N_1124,In_673,In_507);
nor U1125 (N_1125,In_72,In_552);
xnor U1126 (N_1126,In_1538,In_1912);
nor U1127 (N_1127,In_1811,In_1920);
or U1128 (N_1128,In_1857,In_1135);
and U1129 (N_1129,In_788,In_1884);
xor U1130 (N_1130,In_719,In_1534);
xnor U1131 (N_1131,In_768,In_249);
xor U1132 (N_1132,In_293,In_1448);
or U1133 (N_1133,In_689,In_1164);
nor U1134 (N_1134,In_1201,In_1842);
and U1135 (N_1135,In_247,In_253);
and U1136 (N_1136,In_593,In_539);
nand U1137 (N_1137,In_1386,In_387);
nor U1138 (N_1138,In_1170,In_230);
xnor U1139 (N_1139,In_1845,In_597);
or U1140 (N_1140,In_1590,In_1841);
nor U1141 (N_1141,In_1399,In_1531);
nand U1142 (N_1142,In_227,In_1748);
xor U1143 (N_1143,In_1708,In_230);
and U1144 (N_1144,In_1162,In_609);
xnor U1145 (N_1145,In_920,In_572);
and U1146 (N_1146,In_638,In_196);
and U1147 (N_1147,In_1063,In_134);
xnor U1148 (N_1148,In_1858,In_1696);
or U1149 (N_1149,In_116,In_1959);
or U1150 (N_1150,In_1737,In_1908);
xnor U1151 (N_1151,In_375,In_978);
nand U1152 (N_1152,In_837,In_1107);
and U1153 (N_1153,In_535,In_1930);
or U1154 (N_1154,In_1034,In_289);
or U1155 (N_1155,In_228,In_1550);
nand U1156 (N_1156,In_1650,In_672);
xnor U1157 (N_1157,In_1323,In_1778);
or U1158 (N_1158,In_1802,In_1610);
or U1159 (N_1159,In_1044,In_1791);
nor U1160 (N_1160,In_1641,In_1032);
nor U1161 (N_1161,In_604,In_1099);
nand U1162 (N_1162,In_303,In_43);
nand U1163 (N_1163,In_363,In_618);
and U1164 (N_1164,In_1947,In_617);
xor U1165 (N_1165,In_485,In_1255);
and U1166 (N_1166,In_623,In_834);
or U1167 (N_1167,In_51,In_592);
xnor U1168 (N_1168,In_450,In_389);
and U1169 (N_1169,In_561,In_1640);
or U1170 (N_1170,In_1251,In_105);
nand U1171 (N_1171,In_897,In_1084);
nand U1172 (N_1172,In_448,In_168);
xnor U1173 (N_1173,In_1296,In_456);
nor U1174 (N_1174,In_151,In_920);
nand U1175 (N_1175,In_1886,In_1733);
or U1176 (N_1176,In_464,In_935);
and U1177 (N_1177,In_52,In_1929);
nand U1178 (N_1178,In_271,In_231);
nand U1179 (N_1179,In_1168,In_1016);
nor U1180 (N_1180,In_1147,In_1023);
or U1181 (N_1181,In_861,In_755);
and U1182 (N_1182,In_1591,In_886);
and U1183 (N_1183,In_743,In_534);
xnor U1184 (N_1184,In_34,In_702);
and U1185 (N_1185,In_1313,In_1549);
and U1186 (N_1186,In_802,In_1510);
or U1187 (N_1187,In_216,In_1820);
xor U1188 (N_1188,In_1015,In_1814);
nor U1189 (N_1189,In_959,In_538);
nand U1190 (N_1190,In_458,In_121);
nor U1191 (N_1191,In_377,In_1863);
xnor U1192 (N_1192,In_1921,In_1384);
xnor U1193 (N_1193,In_1525,In_965);
xnor U1194 (N_1194,In_878,In_1285);
xor U1195 (N_1195,In_1907,In_1706);
or U1196 (N_1196,In_1074,In_1226);
and U1197 (N_1197,In_773,In_174);
nand U1198 (N_1198,In_462,In_132);
xnor U1199 (N_1199,In_63,In_449);
nor U1200 (N_1200,In_839,In_1557);
or U1201 (N_1201,In_820,In_457);
xor U1202 (N_1202,In_203,In_877);
or U1203 (N_1203,In_969,In_1091);
xor U1204 (N_1204,In_308,In_124);
xnor U1205 (N_1205,In_1645,In_901);
nand U1206 (N_1206,In_81,In_1007);
and U1207 (N_1207,In_1394,In_626);
and U1208 (N_1208,In_821,In_1623);
xor U1209 (N_1209,In_278,In_1702);
nand U1210 (N_1210,In_1353,In_189);
or U1211 (N_1211,In_1063,In_405);
xor U1212 (N_1212,In_1875,In_1956);
nand U1213 (N_1213,In_135,In_648);
xnor U1214 (N_1214,In_779,In_689);
nand U1215 (N_1215,In_1249,In_445);
and U1216 (N_1216,In_1303,In_921);
xnor U1217 (N_1217,In_1974,In_1742);
nand U1218 (N_1218,In_1473,In_1735);
xor U1219 (N_1219,In_1069,In_1538);
nand U1220 (N_1220,In_205,In_688);
xor U1221 (N_1221,In_94,In_877);
or U1222 (N_1222,In_694,In_1034);
xnor U1223 (N_1223,In_1081,In_712);
and U1224 (N_1224,In_594,In_683);
xnor U1225 (N_1225,In_1832,In_778);
nor U1226 (N_1226,In_1657,In_542);
nor U1227 (N_1227,In_1245,In_84);
nand U1228 (N_1228,In_689,In_547);
nor U1229 (N_1229,In_1712,In_1954);
xor U1230 (N_1230,In_1618,In_747);
xnor U1231 (N_1231,In_1969,In_1176);
nand U1232 (N_1232,In_1477,In_916);
or U1233 (N_1233,In_361,In_760);
xor U1234 (N_1234,In_1123,In_1598);
or U1235 (N_1235,In_1619,In_345);
or U1236 (N_1236,In_1999,In_1225);
and U1237 (N_1237,In_1080,In_414);
xnor U1238 (N_1238,In_61,In_1048);
nand U1239 (N_1239,In_547,In_1119);
nand U1240 (N_1240,In_1052,In_930);
and U1241 (N_1241,In_257,In_1706);
nand U1242 (N_1242,In_1920,In_363);
or U1243 (N_1243,In_1625,In_178);
nor U1244 (N_1244,In_487,In_605);
nand U1245 (N_1245,In_143,In_1284);
nor U1246 (N_1246,In_202,In_609);
nor U1247 (N_1247,In_1508,In_914);
nand U1248 (N_1248,In_398,In_1533);
nand U1249 (N_1249,In_1651,In_221);
nand U1250 (N_1250,In_1361,In_1140);
nand U1251 (N_1251,In_1870,In_239);
xor U1252 (N_1252,In_1439,In_159);
and U1253 (N_1253,In_1529,In_1115);
and U1254 (N_1254,In_698,In_307);
nor U1255 (N_1255,In_165,In_623);
nor U1256 (N_1256,In_1258,In_1823);
nand U1257 (N_1257,In_467,In_1753);
nor U1258 (N_1258,In_849,In_1976);
nor U1259 (N_1259,In_1354,In_352);
or U1260 (N_1260,In_1634,In_1011);
nand U1261 (N_1261,In_963,In_539);
nand U1262 (N_1262,In_1324,In_748);
nor U1263 (N_1263,In_68,In_415);
xnor U1264 (N_1264,In_545,In_1351);
and U1265 (N_1265,In_1785,In_1669);
and U1266 (N_1266,In_457,In_475);
or U1267 (N_1267,In_1805,In_1438);
nor U1268 (N_1268,In_1520,In_1472);
or U1269 (N_1269,In_1508,In_1464);
nand U1270 (N_1270,In_261,In_697);
nor U1271 (N_1271,In_836,In_1461);
or U1272 (N_1272,In_373,In_778);
and U1273 (N_1273,In_51,In_1633);
nor U1274 (N_1274,In_450,In_828);
nand U1275 (N_1275,In_978,In_1289);
nand U1276 (N_1276,In_1857,In_1220);
nor U1277 (N_1277,In_1517,In_1079);
nor U1278 (N_1278,In_1634,In_1690);
nor U1279 (N_1279,In_25,In_1547);
or U1280 (N_1280,In_64,In_8);
xnor U1281 (N_1281,In_1226,In_175);
nor U1282 (N_1282,In_1417,In_1581);
and U1283 (N_1283,In_1694,In_829);
xnor U1284 (N_1284,In_1119,In_915);
and U1285 (N_1285,In_1877,In_846);
and U1286 (N_1286,In_1878,In_1458);
xor U1287 (N_1287,In_1114,In_258);
xor U1288 (N_1288,In_1724,In_355);
nand U1289 (N_1289,In_155,In_1307);
or U1290 (N_1290,In_1042,In_1808);
nand U1291 (N_1291,In_53,In_749);
xor U1292 (N_1292,In_1943,In_317);
or U1293 (N_1293,In_1155,In_431);
nor U1294 (N_1294,In_1699,In_1441);
nor U1295 (N_1295,In_332,In_692);
and U1296 (N_1296,In_1192,In_902);
and U1297 (N_1297,In_1351,In_547);
or U1298 (N_1298,In_123,In_696);
nand U1299 (N_1299,In_23,In_1313);
nor U1300 (N_1300,In_1085,In_492);
nor U1301 (N_1301,In_1486,In_155);
nor U1302 (N_1302,In_865,In_472);
xnor U1303 (N_1303,In_268,In_269);
nand U1304 (N_1304,In_740,In_325);
nor U1305 (N_1305,In_993,In_1174);
or U1306 (N_1306,In_20,In_878);
nor U1307 (N_1307,In_1374,In_653);
or U1308 (N_1308,In_648,In_196);
and U1309 (N_1309,In_189,In_95);
or U1310 (N_1310,In_1788,In_1733);
and U1311 (N_1311,In_1423,In_979);
xor U1312 (N_1312,In_1545,In_501);
nor U1313 (N_1313,In_1242,In_1486);
or U1314 (N_1314,In_1118,In_1995);
nor U1315 (N_1315,In_1674,In_1856);
and U1316 (N_1316,In_507,In_1200);
or U1317 (N_1317,In_1010,In_1808);
and U1318 (N_1318,In_424,In_1303);
or U1319 (N_1319,In_1788,In_539);
and U1320 (N_1320,In_1091,In_1919);
xor U1321 (N_1321,In_774,In_675);
or U1322 (N_1322,In_1426,In_258);
and U1323 (N_1323,In_1987,In_828);
and U1324 (N_1324,In_1511,In_1761);
and U1325 (N_1325,In_773,In_1454);
and U1326 (N_1326,In_761,In_975);
or U1327 (N_1327,In_823,In_1843);
and U1328 (N_1328,In_1640,In_240);
or U1329 (N_1329,In_1907,In_733);
or U1330 (N_1330,In_1274,In_524);
nor U1331 (N_1331,In_75,In_1993);
nand U1332 (N_1332,In_1984,In_107);
nor U1333 (N_1333,In_573,In_916);
xnor U1334 (N_1334,In_585,In_334);
and U1335 (N_1335,In_23,In_1164);
xnor U1336 (N_1336,In_1320,In_1917);
xor U1337 (N_1337,In_836,In_1695);
nor U1338 (N_1338,In_1530,In_1093);
xor U1339 (N_1339,In_613,In_36);
nor U1340 (N_1340,In_1358,In_37);
or U1341 (N_1341,In_296,In_479);
and U1342 (N_1342,In_1086,In_1941);
nand U1343 (N_1343,In_1394,In_1533);
or U1344 (N_1344,In_1572,In_1553);
xor U1345 (N_1345,In_1200,In_1489);
or U1346 (N_1346,In_1384,In_890);
xor U1347 (N_1347,In_1983,In_1625);
or U1348 (N_1348,In_4,In_734);
nand U1349 (N_1349,In_1174,In_1425);
and U1350 (N_1350,In_971,In_60);
and U1351 (N_1351,In_810,In_805);
nor U1352 (N_1352,In_123,In_1957);
or U1353 (N_1353,In_1098,In_319);
nor U1354 (N_1354,In_1901,In_1067);
or U1355 (N_1355,In_366,In_433);
nand U1356 (N_1356,In_128,In_184);
nor U1357 (N_1357,In_803,In_295);
xor U1358 (N_1358,In_1471,In_1711);
xor U1359 (N_1359,In_387,In_856);
xnor U1360 (N_1360,In_47,In_435);
nand U1361 (N_1361,In_1991,In_1258);
and U1362 (N_1362,In_1495,In_110);
nor U1363 (N_1363,In_1041,In_28);
nor U1364 (N_1364,In_1487,In_335);
nand U1365 (N_1365,In_1635,In_643);
or U1366 (N_1366,In_376,In_1855);
nand U1367 (N_1367,In_1418,In_1595);
and U1368 (N_1368,In_1548,In_1935);
xnor U1369 (N_1369,In_1092,In_420);
xor U1370 (N_1370,In_1151,In_773);
nand U1371 (N_1371,In_513,In_1953);
xnor U1372 (N_1372,In_1536,In_23);
xor U1373 (N_1373,In_373,In_1332);
nor U1374 (N_1374,In_1082,In_1628);
or U1375 (N_1375,In_1109,In_1897);
nand U1376 (N_1376,In_1706,In_1009);
or U1377 (N_1377,In_559,In_909);
nor U1378 (N_1378,In_1569,In_1927);
nand U1379 (N_1379,In_265,In_617);
and U1380 (N_1380,In_1004,In_1069);
or U1381 (N_1381,In_1617,In_1855);
xor U1382 (N_1382,In_556,In_13);
nor U1383 (N_1383,In_875,In_302);
and U1384 (N_1384,In_369,In_1227);
nor U1385 (N_1385,In_1563,In_573);
or U1386 (N_1386,In_1220,In_1794);
nor U1387 (N_1387,In_69,In_258);
or U1388 (N_1388,In_1279,In_1101);
or U1389 (N_1389,In_373,In_1471);
nand U1390 (N_1390,In_0,In_107);
xor U1391 (N_1391,In_961,In_1168);
or U1392 (N_1392,In_1677,In_1013);
and U1393 (N_1393,In_865,In_341);
and U1394 (N_1394,In_279,In_1712);
xor U1395 (N_1395,In_1991,In_1753);
or U1396 (N_1396,In_1777,In_1912);
xor U1397 (N_1397,In_1515,In_1291);
nor U1398 (N_1398,In_1836,In_1084);
nand U1399 (N_1399,In_999,In_459);
nor U1400 (N_1400,In_1351,In_1722);
or U1401 (N_1401,In_1439,In_1522);
or U1402 (N_1402,In_374,In_890);
nand U1403 (N_1403,In_1442,In_1119);
xnor U1404 (N_1404,In_466,In_1884);
and U1405 (N_1405,In_1030,In_1225);
nand U1406 (N_1406,In_478,In_1300);
and U1407 (N_1407,In_1497,In_1611);
nand U1408 (N_1408,In_1366,In_994);
and U1409 (N_1409,In_486,In_575);
and U1410 (N_1410,In_1654,In_1244);
and U1411 (N_1411,In_1192,In_999);
nor U1412 (N_1412,In_926,In_916);
xnor U1413 (N_1413,In_130,In_714);
and U1414 (N_1414,In_423,In_1492);
nand U1415 (N_1415,In_1637,In_57);
nand U1416 (N_1416,In_904,In_983);
and U1417 (N_1417,In_1998,In_1323);
or U1418 (N_1418,In_90,In_45);
xnor U1419 (N_1419,In_1133,In_242);
nand U1420 (N_1420,In_1131,In_1982);
nor U1421 (N_1421,In_58,In_1259);
and U1422 (N_1422,In_1809,In_825);
nor U1423 (N_1423,In_1646,In_1963);
and U1424 (N_1424,In_1339,In_289);
xnor U1425 (N_1425,In_218,In_1939);
nor U1426 (N_1426,In_906,In_66);
nand U1427 (N_1427,In_658,In_655);
xnor U1428 (N_1428,In_461,In_519);
or U1429 (N_1429,In_1218,In_410);
or U1430 (N_1430,In_1506,In_1374);
and U1431 (N_1431,In_869,In_187);
and U1432 (N_1432,In_946,In_271);
nor U1433 (N_1433,In_807,In_1835);
nand U1434 (N_1434,In_669,In_1107);
nand U1435 (N_1435,In_1745,In_1594);
xor U1436 (N_1436,In_1160,In_1324);
nor U1437 (N_1437,In_1612,In_383);
and U1438 (N_1438,In_896,In_553);
xor U1439 (N_1439,In_304,In_1121);
xor U1440 (N_1440,In_243,In_1959);
or U1441 (N_1441,In_1322,In_250);
nand U1442 (N_1442,In_709,In_467);
or U1443 (N_1443,In_1461,In_574);
nor U1444 (N_1444,In_270,In_1220);
nand U1445 (N_1445,In_1814,In_1123);
xor U1446 (N_1446,In_1677,In_583);
nand U1447 (N_1447,In_203,In_943);
xor U1448 (N_1448,In_1842,In_76);
nand U1449 (N_1449,In_887,In_1185);
nand U1450 (N_1450,In_836,In_856);
xor U1451 (N_1451,In_531,In_1741);
and U1452 (N_1452,In_1766,In_1756);
nand U1453 (N_1453,In_930,In_1622);
nand U1454 (N_1454,In_435,In_597);
nor U1455 (N_1455,In_618,In_1886);
nor U1456 (N_1456,In_1152,In_1386);
or U1457 (N_1457,In_1419,In_228);
xor U1458 (N_1458,In_620,In_1530);
xnor U1459 (N_1459,In_197,In_1556);
nor U1460 (N_1460,In_1023,In_1241);
and U1461 (N_1461,In_38,In_242);
xnor U1462 (N_1462,In_1212,In_489);
or U1463 (N_1463,In_1670,In_325);
xnor U1464 (N_1464,In_1940,In_1438);
nand U1465 (N_1465,In_1233,In_1246);
nand U1466 (N_1466,In_880,In_469);
and U1467 (N_1467,In_1506,In_440);
and U1468 (N_1468,In_1164,In_1182);
nand U1469 (N_1469,In_153,In_1657);
xnor U1470 (N_1470,In_729,In_18);
nand U1471 (N_1471,In_1740,In_297);
or U1472 (N_1472,In_1245,In_981);
xnor U1473 (N_1473,In_22,In_94);
xor U1474 (N_1474,In_1838,In_656);
xnor U1475 (N_1475,In_1963,In_826);
nor U1476 (N_1476,In_1061,In_1770);
or U1477 (N_1477,In_1541,In_1307);
nand U1478 (N_1478,In_1890,In_180);
nor U1479 (N_1479,In_1630,In_1315);
or U1480 (N_1480,In_1800,In_159);
nand U1481 (N_1481,In_1702,In_920);
and U1482 (N_1482,In_663,In_1702);
nand U1483 (N_1483,In_1553,In_1007);
xnor U1484 (N_1484,In_983,In_211);
nand U1485 (N_1485,In_89,In_733);
or U1486 (N_1486,In_931,In_1161);
nor U1487 (N_1487,In_1258,In_1117);
nor U1488 (N_1488,In_1522,In_1343);
and U1489 (N_1489,In_842,In_463);
and U1490 (N_1490,In_195,In_1815);
nand U1491 (N_1491,In_380,In_992);
xor U1492 (N_1492,In_1979,In_1218);
or U1493 (N_1493,In_571,In_391);
and U1494 (N_1494,In_1448,In_76);
xnor U1495 (N_1495,In_134,In_1841);
xor U1496 (N_1496,In_1169,In_656);
and U1497 (N_1497,In_604,In_1274);
nor U1498 (N_1498,In_853,In_1328);
or U1499 (N_1499,In_1379,In_1580);
and U1500 (N_1500,In_217,In_1482);
nor U1501 (N_1501,In_161,In_1210);
or U1502 (N_1502,In_321,In_1126);
xnor U1503 (N_1503,In_1444,In_1151);
or U1504 (N_1504,In_1386,In_569);
and U1505 (N_1505,In_70,In_1481);
and U1506 (N_1506,In_1505,In_515);
or U1507 (N_1507,In_466,In_1804);
xor U1508 (N_1508,In_1708,In_1821);
and U1509 (N_1509,In_1077,In_1839);
nand U1510 (N_1510,In_57,In_1163);
xnor U1511 (N_1511,In_1626,In_1023);
or U1512 (N_1512,In_1931,In_1189);
or U1513 (N_1513,In_1598,In_1104);
xnor U1514 (N_1514,In_1767,In_591);
xnor U1515 (N_1515,In_1635,In_237);
and U1516 (N_1516,In_519,In_1518);
nor U1517 (N_1517,In_494,In_64);
xor U1518 (N_1518,In_829,In_1004);
nand U1519 (N_1519,In_1207,In_777);
or U1520 (N_1520,In_84,In_1222);
nand U1521 (N_1521,In_508,In_1314);
nand U1522 (N_1522,In_743,In_1217);
and U1523 (N_1523,In_1882,In_935);
and U1524 (N_1524,In_1755,In_1490);
nand U1525 (N_1525,In_1727,In_647);
nand U1526 (N_1526,In_1854,In_1447);
nor U1527 (N_1527,In_1374,In_1735);
nand U1528 (N_1528,In_1401,In_97);
xnor U1529 (N_1529,In_46,In_1461);
and U1530 (N_1530,In_1661,In_445);
or U1531 (N_1531,In_663,In_447);
or U1532 (N_1532,In_572,In_1010);
or U1533 (N_1533,In_187,In_1817);
and U1534 (N_1534,In_1130,In_1366);
xor U1535 (N_1535,In_766,In_1683);
nand U1536 (N_1536,In_48,In_358);
nor U1537 (N_1537,In_213,In_1185);
nand U1538 (N_1538,In_1784,In_131);
nor U1539 (N_1539,In_1916,In_868);
and U1540 (N_1540,In_642,In_469);
or U1541 (N_1541,In_587,In_609);
nand U1542 (N_1542,In_1624,In_1150);
nand U1543 (N_1543,In_1534,In_1210);
and U1544 (N_1544,In_111,In_987);
and U1545 (N_1545,In_1185,In_1578);
or U1546 (N_1546,In_990,In_1267);
or U1547 (N_1547,In_563,In_1317);
and U1548 (N_1548,In_179,In_755);
xor U1549 (N_1549,In_1287,In_1711);
and U1550 (N_1550,In_905,In_32);
nor U1551 (N_1551,In_608,In_13);
xor U1552 (N_1552,In_1141,In_948);
and U1553 (N_1553,In_197,In_1180);
nand U1554 (N_1554,In_1270,In_669);
xor U1555 (N_1555,In_935,In_1346);
and U1556 (N_1556,In_879,In_198);
nand U1557 (N_1557,In_1398,In_1178);
and U1558 (N_1558,In_812,In_694);
xor U1559 (N_1559,In_1400,In_629);
xor U1560 (N_1560,In_1232,In_596);
xor U1561 (N_1561,In_779,In_1915);
and U1562 (N_1562,In_1592,In_717);
and U1563 (N_1563,In_518,In_1615);
or U1564 (N_1564,In_651,In_1718);
and U1565 (N_1565,In_1878,In_1283);
nand U1566 (N_1566,In_241,In_931);
nand U1567 (N_1567,In_1287,In_685);
or U1568 (N_1568,In_1923,In_1135);
or U1569 (N_1569,In_1408,In_1844);
nor U1570 (N_1570,In_1570,In_1207);
nor U1571 (N_1571,In_772,In_539);
and U1572 (N_1572,In_81,In_423);
xnor U1573 (N_1573,In_675,In_1392);
nand U1574 (N_1574,In_881,In_138);
and U1575 (N_1575,In_1512,In_1399);
xor U1576 (N_1576,In_1520,In_161);
and U1577 (N_1577,In_142,In_1164);
nor U1578 (N_1578,In_665,In_211);
and U1579 (N_1579,In_1953,In_900);
and U1580 (N_1580,In_1680,In_936);
and U1581 (N_1581,In_592,In_762);
or U1582 (N_1582,In_1904,In_1641);
nor U1583 (N_1583,In_1082,In_459);
xor U1584 (N_1584,In_1195,In_1382);
and U1585 (N_1585,In_1806,In_595);
xor U1586 (N_1586,In_1266,In_594);
or U1587 (N_1587,In_524,In_1814);
nand U1588 (N_1588,In_288,In_1147);
nand U1589 (N_1589,In_1801,In_251);
xor U1590 (N_1590,In_498,In_914);
nand U1591 (N_1591,In_537,In_1860);
or U1592 (N_1592,In_446,In_1540);
xor U1593 (N_1593,In_16,In_1939);
nand U1594 (N_1594,In_398,In_644);
nand U1595 (N_1595,In_1972,In_269);
and U1596 (N_1596,In_1585,In_60);
and U1597 (N_1597,In_536,In_1237);
xnor U1598 (N_1598,In_948,In_1444);
xnor U1599 (N_1599,In_1731,In_1368);
or U1600 (N_1600,In_1572,In_894);
nor U1601 (N_1601,In_363,In_1421);
or U1602 (N_1602,In_637,In_1718);
or U1603 (N_1603,In_1655,In_890);
or U1604 (N_1604,In_819,In_1847);
nor U1605 (N_1605,In_1092,In_1912);
or U1606 (N_1606,In_1718,In_631);
xnor U1607 (N_1607,In_681,In_1788);
or U1608 (N_1608,In_842,In_1994);
nand U1609 (N_1609,In_18,In_367);
and U1610 (N_1610,In_762,In_1952);
xor U1611 (N_1611,In_302,In_1480);
xnor U1612 (N_1612,In_1216,In_1370);
xor U1613 (N_1613,In_445,In_1055);
nor U1614 (N_1614,In_1461,In_882);
nor U1615 (N_1615,In_1608,In_895);
or U1616 (N_1616,In_120,In_576);
or U1617 (N_1617,In_1088,In_1825);
nand U1618 (N_1618,In_1866,In_1513);
or U1619 (N_1619,In_1810,In_457);
and U1620 (N_1620,In_1473,In_1910);
or U1621 (N_1621,In_657,In_1248);
or U1622 (N_1622,In_741,In_362);
nand U1623 (N_1623,In_1634,In_1941);
and U1624 (N_1624,In_1613,In_721);
nor U1625 (N_1625,In_225,In_29);
nor U1626 (N_1626,In_1736,In_221);
xor U1627 (N_1627,In_736,In_209);
nor U1628 (N_1628,In_1233,In_1623);
nand U1629 (N_1629,In_540,In_644);
nor U1630 (N_1630,In_122,In_724);
nor U1631 (N_1631,In_1961,In_1573);
nand U1632 (N_1632,In_690,In_405);
nand U1633 (N_1633,In_1564,In_491);
nor U1634 (N_1634,In_1110,In_1044);
nand U1635 (N_1635,In_1591,In_1224);
nor U1636 (N_1636,In_1921,In_413);
and U1637 (N_1637,In_1541,In_1682);
or U1638 (N_1638,In_657,In_1892);
and U1639 (N_1639,In_1721,In_884);
nand U1640 (N_1640,In_7,In_467);
xor U1641 (N_1641,In_604,In_1518);
xor U1642 (N_1642,In_688,In_110);
and U1643 (N_1643,In_1340,In_460);
xor U1644 (N_1644,In_1932,In_568);
and U1645 (N_1645,In_230,In_163);
and U1646 (N_1646,In_879,In_1053);
and U1647 (N_1647,In_272,In_994);
nor U1648 (N_1648,In_1838,In_1115);
nand U1649 (N_1649,In_345,In_1505);
nand U1650 (N_1650,In_1450,In_1094);
and U1651 (N_1651,In_1057,In_1367);
and U1652 (N_1652,In_183,In_642);
xnor U1653 (N_1653,In_683,In_383);
xnor U1654 (N_1654,In_1539,In_1005);
xnor U1655 (N_1655,In_1411,In_1988);
xor U1656 (N_1656,In_332,In_568);
xnor U1657 (N_1657,In_308,In_39);
nor U1658 (N_1658,In_1393,In_1796);
nor U1659 (N_1659,In_1670,In_499);
nor U1660 (N_1660,In_439,In_1721);
nand U1661 (N_1661,In_408,In_1758);
and U1662 (N_1662,In_550,In_1034);
nor U1663 (N_1663,In_1295,In_1129);
nand U1664 (N_1664,In_276,In_1794);
nor U1665 (N_1665,In_1224,In_9);
nor U1666 (N_1666,In_1826,In_338);
or U1667 (N_1667,In_1413,In_745);
nor U1668 (N_1668,In_568,In_448);
or U1669 (N_1669,In_404,In_173);
nor U1670 (N_1670,In_943,In_436);
and U1671 (N_1671,In_153,In_248);
and U1672 (N_1672,In_905,In_1369);
nand U1673 (N_1673,In_262,In_1668);
or U1674 (N_1674,In_1843,In_488);
xor U1675 (N_1675,In_672,In_306);
or U1676 (N_1676,In_634,In_1401);
or U1677 (N_1677,In_828,In_146);
nand U1678 (N_1678,In_1679,In_787);
or U1679 (N_1679,In_1292,In_710);
xnor U1680 (N_1680,In_576,In_1543);
or U1681 (N_1681,In_1715,In_387);
nand U1682 (N_1682,In_763,In_1186);
nor U1683 (N_1683,In_861,In_1724);
nor U1684 (N_1684,In_1930,In_1694);
nand U1685 (N_1685,In_1249,In_1963);
xor U1686 (N_1686,In_233,In_862);
xor U1687 (N_1687,In_60,In_3);
and U1688 (N_1688,In_1087,In_1035);
nor U1689 (N_1689,In_1679,In_1009);
nand U1690 (N_1690,In_566,In_794);
nor U1691 (N_1691,In_801,In_869);
xnor U1692 (N_1692,In_431,In_1279);
xor U1693 (N_1693,In_26,In_1988);
nand U1694 (N_1694,In_405,In_1269);
nand U1695 (N_1695,In_521,In_1847);
nand U1696 (N_1696,In_83,In_237);
nor U1697 (N_1697,In_931,In_124);
or U1698 (N_1698,In_1845,In_814);
and U1699 (N_1699,In_499,In_1933);
nand U1700 (N_1700,In_216,In_1308);
and U1701 (N_1701,In_1815,In_393);
xnor U1702 (N_1702,In_612,In_969);
nand U1703 (N_1703,In_494,In_1341);
xor U1704 (N_1704,In_156,In_685);
and U1705 (N_1705,In_1212,In_938);
nand U1706 (N_1706,In_456,In_1340);
nor U1707 (N_1707,In_1511,In_320);
nand U1708 (N_1708,In_787,In_1991);
or U1709 (N_1709,In_226,In_656);
nor U1710 (N_1710,In_1619,In_1005);
nor U1711 (N_1711,In_1601,In_611);
xor U1712 (N_1712,In_803,In_1794);
or U1713 (N_1713,In_1499,In_598);
xnor U1714 (N_1714,In_1792,In_833);
xnor U1715 (N_1715,In_886,In_1161);
nand U1716 (N_1716,In_683,In_1391);
nand U1717 (N_1717,In_127,In_202);
nand U1718 (N_1718,In_95,In_1673);
nand U1719 (N_1719,In_1172,In_1135);
or U1720 (N_1720,In_600,In_1139);
or U1721 (N_1721,In_473,In_177);
xnor U1722 (N_1722,In_954,In_1632);
or U1723 (N_1723,In_1046,In_189);
nand U1724 (N_1724,In_1872,In_907);
or U1725 (N_1725,In_483,In_663);
and U1726 (N_1726,In_688,In_513);
xor U1727 (N_1727,In_989,In_1705);
or U1728 (N_1728,In_870,In_1795);
xor U1729 (N_1729,In_1553,In_1327);
and U1730 (N_1730,In_1308,In_940);
xor U1731 (N_1731,In_788,In_1261);
and U1732 (N_1732,In_1857,In_745);
nor U1733 (N_1733,In_520,In_1941);
nand U1734 (N_1734,In_296,In_189);
and U1735 (N_1735,In_1348,In_316);
nor U1736 (N_1736,In_510,In_441);
xor U1737 (N_1737,In_1380,In_892);
or U1738 (N_1738,In_1239,In_361);
xnor U1739 (N_1739,In_167,In_73);
xor U1740 (N_1740,In_527,In_947);
nor U1741 (N_1741,In_1447,In_872);
xor U1742 (N_1742,In_1721,In_164);
nand U1743 (N_1743,In_1429,In_1988);
xor U1744 (N_1744,In_1393,In_42);
and U1745 (N_1745,In_1757,In_1971);
nand U1746 (N_1746,In_54,In_1212);
nand U1747 (N_1747,In_580,In_1228);
and U1748 (N_1748,In_1455,In_527);
or U1749 (N_1749,In_1664,In_1606);
nand U1750 (N_1750,In_145,In_1135);
nor U1751 (N_1751,In_1964,In_1379);
or U1752 (N_1752,In_1978,In_1122);
xor U1753 (N_1753,In_299,In_1480);
and U1754 (N_1754,In_1667,In_872);
and U1755 (N_1755,In_1628,In_169);
xor U1756 (N_1756,In_1015,In_1981);
or U1757 (N_1757,In_199,In_1010);
or U1758 (N_1758,In_1652,In_744);
or U1759 (N_1759,In_1531,In_314);
nand U1760 (N_1760,In_161,In_1162);
and U1761 (N_1761,In_1848,In_1978);
or U1762 (N_1762,In_654,In_818);
nor U1763 (N_1763,In_391,In_1044);
or U1764 (N_1764,In_1703,In_885);
nor U1765 (N_1765,In_1278,In_1234);
or U1766 (N_1766,In_1825,In_191);
nor U1767 (N_1767,In_1696,In_1066);
or U1768 (N_1768,In_153,In_780);
nand U1769 (N_1769,In_1811,In_267);
nand U1770 (N_1770,In_862,In_1393);
or U1771 (N_1771,In_869,In_1814);
and U1772 (N_1772,In_1223,In_154);
xor U1773 (N_1773,In_440,In_276);
xor U1774 (N_1774,In_391,In_513);
and U1775 (N_1775,In_1372,In_1546);
nor U1776 (N_1776,In_1182,In_885);
nand U1777 (N_1777,In_232,In_278);
nand U1778 (N_1778,In_661,In_732);
xor U1779 (N_1779,In_1741,In_271);
nand U1780 (N_1780,In_1772,In_1527);
xnor U1781 (N_1781,In_510,In_667);
and U1782 (N_1782,In_1040,In_26);
or U1783 (N_1783,In_10,In_385);
or U1784 (N_1784,In_1942,In_1433);
or U1785 (N_1785,In_892,In_733);
nand U1786 (N_1786,In_1197,In_1800);
xnor U1787 (N_1787,In_211,In_1117);
and U1788 (N_1788,In_1222,In_667);
or U1789 (N_1789,In_1720,In_1366);
xnor U1790 (N_1790,In_482,In_1408);
nor U1791 (N_1791,In_1442,In_231);
and U1792 (N_1792,In_1563,In_272);
or U1793 (N_1793,In_276,In_1686);
xor U1794 (N_1794,In_411,In_325);
and U1795 (N_1795,In_702,In_482);
xor U1796 (N_1796,In_824,In_1512);
or U1797 (N_1797,In_1606,In_1056);
or U1798 (N_1798,In_67,In_92);
xnor U1799 (N_1799,In_1032,In_869);
nand U1800 (N_1800,In_291,In_1984);
xor U1801 (N_1801,In_1276,In_1960);
nand U1802 (N_1802,In_126,In_1270);
and U1803 (N_1803,In_967,In_1842);
nand U1804 (N_1804,In_1751,In_1873);
and U1805 (N_1805,In_160,In_1149);
nor U1806 (N_1806,In_330,In_192);
or U1807 (N_1807,In_1425,In_789);
nand U1808 (N_1808,In_311,In_700);
nand U1809 (N_1809,In_413,In_204);
or U1810 (N_1810,In_156,In_1731);
nand U1811 (N_1811,In_1396,In_131);
nor U1812 (N_1812,In_1976,In_410);
and U1813 (N_1813,In_770,In_1700);
nand U1814 (N_1814,In_1964,In_1088);
nand U1815 (N_1815,In_1393,In_1487);
or U1816 (N_1816,In_568,In_185);
nor U1817 (N_1817,In_318,In_901);
nor U1818 (N_1818,In_584,In_1041);
nand U1819 (N_1819,In_309,In_1119);
nand U1820 (N_1820,In_336,In_1488);
or U1821 (N_1821,In_1305,In_522);
nor U1822 (N_1822,In_1119,In_1660);
and U1823 (N_1823,In_511,In_1542);
xor U1824 (N_1824,In_1665,In_80);
xor U1825 (N_1825,In_1221,In_1430);
nor U1826 (N_1826,In_39,In_973);
nand U1827 (N_1827,In_86,In_1711);
and U1828 (N_1828,In_1259,In_1761);
and U1829 (N_1829,In_1807,In_1682);
xor U1830 (N_1830,In_306,In_1742);
nor U1831 (N_1831,In_1166,In_551);
and U1832 (N_1832,In_12,In_1223);
nor U1833 (N_1833,In_1806,In_1612);
xnor U1834 (N_1834,In_63,In_313);
nor U1835 (N_1835,In_217,In_616);
nand U1836 (N_1836,In_1015,In_139);
or U1837 (N_1837,In_150,In_1468);
xor U1838 (N_1838,In_770,In_1794);
xor U1839 (N_1839,In_1530,In_1397);
xor U1840 (N_1840,In_783,In_1916);
or U1841 (N_1841,In_1426,In_509);
and U1842 (N_1842,In_1539,In_141);
nand U1843 (N_1843,In_822,In_1356);
or U1844 (N_1844,In_400,In_1329);
xnor U1845 (N_1845,In_1894,In_384);
and U1846 (N_1846,In_996,In_1350);
nand U1847 (N_1847,In_958,In_855);
or U1848 (N_1848,In_1224,In_1205);
nor U1849 (N_1849,In_377,In_701);
xnor U1850 (N_1850,In_1866,In_468);
xor U1851 (N_1851,In_64,In_644);
or U1852 (N_1852,In_934,In_191);
and U1853 (N_1853,In_1375,In_693);
nand U1854 (N_1854,In_1099,In_487);
or U1855 (N_1855,In_1405,In_234);
nand U1856 (N_1856,In_556,In_1873);
or U1857 (N_1857,In_1388,In_1090);
xnor U1858 (N_1858,In_1805,In_643);
or U1859 (N_1859,In_862,In_346);
xor U1860 (N_1860,In_1168,In_1661);
nand U1861 (N_1861,In_1861,In_870);
and U1862 (N_1862,In_1893,In_1792);
nand U1863 (N_1863,In_1504,In_578);
xnor U1864 (N_1864,In_284,In_243);
xnor U1865 (N_1865,In_767,In_779);
and U1866 (N_1866,In_1471,In_1448);
xnor U1867 (N_1867,In_655,In_1954);
and U1868 (N_1868,In_1725,In_1271);
nand U1869 (N_1869,In_36,In_638);
xnor U1870 (N_1870,In_1800,In_1263);
xnor U1871 (N_1871,In_1230,In_494);
nand U1872 (N_1872,In_1952,In_1560);
xor U1873 (N_1873,In_1370,In_1118);
or U1874 (N_1874,In_1212,In_1762);
or U1875 (N_1875,In_225,In_1744);
and U1876 (N_1876,In_941,In_1721);
or U1877 (N_1877,In_769,In_589);
or U1878 (N_1878,In_447,In_851);
nand U1879 (N_1879,In_84,In_1704);
nor U1880 (N_1880,In_1651,In_1150);
or U1881 (N_1881,In_1660,In_787);
nand U1882 (N_1882,In_50,In_1777);
nor U1883 (N_1883,In_800,In_881);
and U1884 (N_1884,In_1658,In_579);
nand U1885 (N_1885,In_1046,In_806);
nand U1886 (N_1886,In_144,In_1494);
xnor U1887 (N_1887,In_1980,In_1314);
nand U1888 (N_1888,In_1727,In_429);
xor U1889 (N_1889,In_25,In_366);
nand U1890 (N_1890,In_984,In_1255);
or U1891 (N_1891,In_285,In_755);
and U1892 (N_1892,In_1753,In_1117);
nand U1893 (N_1893,In_697,In_998);
nand U1894 (N_1894,In_201,In_62);
nand U1895 (N_1895,In_893,In_232);
xor U1896 (N_1896,In_181,In_114);
or U1897 (N_1897,In_35,In_118);
nor U1898 (N_1898,In_1975,In_1852);
nand U1899 (N_1899,In_1193,In_1434);
xor U1900 (N_1900,In_261,In_1416);
and U1901 (N_1901,In_1333,In_362);
xor U1902 (N_1902,In_1507,In_1894);
nand U1903 (N_1903,In_777,In_715);
and U1904 (N_1904,In_1653,In_421);
nor U1905 (N_1905,In_765,In_1599);
and U1906 (N_1906,In_57,In_839);
nand U1907 (N_1907,In_1032,In_852);
nor U1908 (N_1908,In_1391,In_611);
and U1909 (N_1909,In_1417,In_55);
and U1910 (N_1910,In_70,In_1955);
nand U1911 (N_1911,In_128,In_444);
and U1912 (N_1912,In_1083,In_929);
nand U1913 (N_1913,In_1650,In_1001);
nand U1914 (N_1914,In_1079,In_524);
and U1915 (N_1915,In_1547,In_769);
or U1916 (N_1916,In_589,In_1496);
nand U1917 (N_1917,In_39,In_1159);
nand U1918 (N_1918,In_1952,In_840);
nand U1919 (N_1919,In_1763,In_1319);
nand U1920 (N_1920,In_1172,In_1688);
and U1921 (N_1921,In_1027,In_1401);
nor U1922 (N_1922,In_1077,In_1166);
or U1923 (N_1923,In_1513,In_94);
nor U1924 (N_1924,In_1988,In_1884);
and U1925 (N_1925,In_1660,In_1570);
or U1926 (N_1926,In_1735,In_320);
nor U1927 (N_1927,In_48,In_264);
nand U1928 (N_1928,In_483,In_1785);
and U1929 (N_1929,In_1770,In_977);
or U1930 (N_1930,In_285,In_869);
or U1931 (N_1931,In_261,In_85);
nand U1932 (N_1932,In_35,In_1929);
or U1933 (N_1933,In_540,In_1103);
nor U1934 (N_1934,In_296,In_1639);
and U1935 (N_1935,In_249,In_931);
and U1936 (N_1936,In_287,In_1521);
and U1937 (N_1937,In_924,In_1764);
and U1938 (N_1938,In_959,In_8);
nor U1939 (N_1939,In_1263,In_1680);
and U1940 (N_1940,In_230,In_1126);
and U1941 (N_1941,In_57,In_106);
nor U1942 (N_1942,In_1866,In_6);
nor U1943 (N_1943,In_479,In_1817);
xnor U1944 (N_1944,In_1756,In_1781);
or U1945 (N_1945,In_349,In_1353);
xor U1946 (N_1946,In_514,In_944);
nor U1947 (N_1947,In_1935,In_1541);
nand U1948 (N_1948,In_45,In_1076);
xor U1949 (N_1949,In_1631,In_1433);
nand U1950 (N_1950,In_1730,In_1815);
nand U1951 (N_1951,In_215,In_1025);
nand U1952 (N_1952,In_885,In_1345);
and U1953 (N_1953,In_1643,In_1181);
xnor U1954 (N_1954,In_1147,In_1164);
nand U1955 (N_1955,In_953,In_1173);
xnor U1956 (N_1956,In_864,In_352);
and U1957 (N_1957,In_36,In_627);
nor U1958 (N_1958,In_836,In_894);
xnor U1959 (N_1959,In_1039,In_1575);
and U1960 (N_1960,In_322,In_534);
and U1961 (N_1961,In_1311,In_546);
nand U1962 (N_1962,In_576,In_967);
and U1963 (N_1963,In_954,In_723);
or U1964 (N_1964,In_213,In_282);
nand U1965 (N_1965,In_1962,In_1632);
nand U1966 (N_1966,In_1834,In_461);
and U1967 (N_1967,In_1707,In_500);
and U1968 (N_1968,In_1773,In_562);
and U1969 (N_1969,In_1918,In_1050);
xnor U1970 (N_1970,In_227,In_1333);
xor U1971 (N_1971,In_1643,In_460);
nand U1972 (N_1972,In_1837,In_1215);
xor U1973 (N_1973,In_687,In_1586);
nand U1974 (N_1974,In_1650,In_1367);
nand U1975 (N_1975,In_853,In_402);
or U1976 (N_1976,In_855,In_1050);
nand U1977 (N_1977,In_1422,In_1027);
nor U1978 (N_1978,In_1862,In_1385);
nor U1979 (N_1979,In_384,In_1760);
nor U1980 (N_1980,In_367,In_1492);
xnor U1981 (N_1981,In_661,In_1171);
nor U1982 (N_1982,In_1028,In_1118);
or U1983 (N_1983,In_116,In_329);
or U1984 (N_1984,In_210,In_747);
and U1985 (N_1985,In_1263,In_524);
or U1986 (N_1986,In_556,In_1695);
and U1987 (N_1987,In_1658,In_684);
nor U1988 (N_1988,In_322,In_1512);
and U1989 (N_1989,In_1342,In_91);
nor U1990 (N_1990,In_1289,In_1587);
nor U1991 (N_1991,In_975,In_505);
xnor U1992 (N_1992,In_286,In_440);
or U1993 (N_1993,In_1319,In_67);
or U1994 (N_1994,In_172,In_1332);
nor U1995 (N_1995,In_392,In_1108);
xor U1996 (N_1996,In_987,In_1592);
xor U1997 (N_1997,In_1683,In_1225);
and U1998 (N_1998,In_708,In_798);
nor U1999 (N_1999,In_480,In_532);
xnor U2000 (N_2000,In_183,In_1254);
xnor U2001 (N_2001,In_1391,In_823);
nand U2002 (N_2002,In_497,In_59);
nor U2003 (N_2003,In_1216,In_1123);
nor U2004 (N_2004,In_1042,In_1621);
and U2005 (N_2005,In_559,In_1822);
xor U2006 (N_2006,In_1399,In_166);
xor U2007 (N_2007,In_1227,In_1235);
xnor U2008 (N_2008,In_1365,In_1944);
and U2009 (N_2009,In_1265,In_745);
xnor U2010 (N_2010,In_588,In_1038);
or U2011 (N_2011,In_1359,In_485);
xnor U2012 (N_2012,In_599,In_204);
nand U2013 (N_2013,In_1950,In_238);
nor U2014 (N_2014,In_1070,In_674);
nor U2015 (N_2015,In_1464,In_420);
or U2016 (N_2016,In_1010,In_565);
xor U2017 (N_2017,In_1867,In_256);
or U2018 (N_2018,In_1114,In_434);
nand U2019 (N_2019,In_201,In_497);
or U2020 (N_2020,In_573,In_1674);
nor U2021 (N_2021,In_1597,In_1301);
nor U2022 (N_2022,In_662,In_1715);
nand U2023 (N_2023,In_272,In_1047);
or U2024 (N_2024,In_1922,In_204);
nor U2025 (N_2025,In_913,In_269);
nand U2026 (N_2026,In_1861,In_566);
and U2027 (N_2027,In_1078,In_689);
and U2028 (N_2028,In_997,In_204);
nor U2029 (N_2029,In_1577,In_81);
nor U2030 (N_2030,In_1235,In_1087);
nand U2031 (N_2031,In_1583,In_1592);
and U2032 (N_2032,In_878,In_547);
xor U2033 (N_2033,In_1733,In_1885);
or U2034 (N_2034,In_403,In_300);
or U2035 (N_2035,In_249,In_80);
nand U2036 (N_2036,In_1296,In_1786);
xor U2037 (N_2037,In_398,In_1309);
or U2038 (N_2038,In_1145,In_775);
and U2039 (N_2039,In_1472,In_1294);
xor U2040 (N_2040,In_1306,In_1565);
or U2041 (N_2041,In_1525,In_1062);
xnor U2042 (N_2042,In_330,In_237);
or U2043 (N_2043,In_1067,In_853);
and U2044 (N_2044,In_1868,In_802);
nand U2045 (N_2045,In_1113,In_395);
xor U2046 (N_2046,In_1120,In_128);
or U2047 (N_2047,In_1032,In_1918);
and U2048 (N_2048,In_1641,In_1957);
xor U2049 (N_2049,In_1153,In_366);
nand U2050 (N_2050,In_98,In_330);
nand U2051 (N_2051,In_681,In_1211);
or U2052 (N_2052,In_1966,In_88);
nand U2053 (N_2053,In_1970,In_323);
xnor U2054 (N_2054,In_887,In_1686);
nor U2055 (N_2055,In_1751,In_1024);
xor U2056 (N_2056,In_702,In_929);
or U2057 (N_2057,In_36,In_1225);
xor U2058 (N_2058,In_1441,In_1698);
or U2059 (N_2059,In_1480,In_974);
or U2060 (N_2060,In_1372,In_680);
xor U2061 (N_2061,In_335,In_414);
nor U2062 (N_2062,In_354,In_1431);
nand U2063 (N_2063,In_1080,In_931);
nand U2064 (N_2064,In_777,In_129);
nand U2065 (N_2065,In_765,In_1067);
or U2066 (N_2066,In_1521,In_1351);
nor U2067 (N_2067,In_1652,In_704);
and U2068 (N_2068,In_445,In_960);
or U2069 (N_2069,In_1397,In_689);
or U2070 (N_2070,In_1829,In_1233);
xor U2071 (N_2071,In_1949,In_1003);
and U2072 (N_2072,In_1317,In_956);
or U2073 (N_2073,In_1911,In_1880);
or U2074 (N_2074,In_188,In_1137);
and U2075 (N_2075,In_574,In_1352);
xor U2076 (N_2076,In_1828,In_61);
nor U2077 (N_2077,In_922,In_1862);
xnor U2078 (N_2078,In_921,In_1298);
or U2079 (N_2079,In_716,In_728);
and U2080 (N_2080,In_966,In_1517);
or U2081 (N_2081,In_989,In_280);
nand U2082 (N_2082,In_402,In_785);
or U2083 (N_2083,In_1256,In_1062);
or U2084 (N_2084,In_190,In_1102);
and U2085 (N_2085,In_684,In_1001);
nand U2086 (N_2086,In_582,In_734);
nor U2087 (N_2087,In_899,In_1594);
nor U2088 (N_2088,In_1616,In_1551);
xnor U2089 (N_2089,In_1142,In_1905);
nor U2090 (N_2090,In_704,In_1235);
and U2091 (N_2091,In_1460,In_1760);
or U2092 (N_2092,In_15,In_257);
nand U2093 (N_2093,In_1579,In_1032);
or U2094 (N_2094,In_1472,In_961);
or U2095 (N_2095,In_1832,In_505);
nand U2096 (N_2096,In_1810,In_717);
or U2097 (N_2097,In_396,In_439);
nor U2098 (N_2098,In_1298,In_1000);
or U2099 (N_2099,In_95,In_1514);
nor U2100 (N_2100,In_1683,In_412);
nor U2101 (N_2101,In_318,In_56);
or U2102 (N_2102,In_1012,In_1691);
nor U2103 (N_2103,In_926,In_1043);
and U2104 (N_2104,In_310,In_67);
nand U2105 (N_2105,In_1306,In_379);
and U2106 (N_2106,In_750,In_1953);
nand U2107 (N_2107,In_1880,In_1424);
nor U2108 (N_2108,In_27,In_548);
nor U2109 (N_2109,In_1292,In_778);
xor U2110 (N_2110,In_840,In_547);
or U2111 (N_2111,In_1219,In_98);
or U2112 (N_2112,In_297,In_1538);
nand U2113 (N_2113,In_1498,In_219);
nand U2114 (N_2114,In_184,In_455);
nor U2115 (N_2115,In_406,In_242);
nand U2116 (N_2116,In_1772,In_503);
and U2117 (N_2117,In_1169,In_519);
or U2118 (N_2118,In_12,In_400);
nor U2119 (N_2119,In_1810,In_1112);
nor U2120 (N_2120,In_727,In_1439);
and U2121 (N_2121,In_1397,In_399);
xor U2122 (N_2122,In_1280,In_1187);
nor U2123 (N_2123,In_1325,In_676);
or U2124 (N_2124,In_734,In_1178);
nand U2125 (N_2125,In_1632,In_1652);
nand U2126 (N_2126,In_585,In_1500);
and U2127 (N_2127,In_762,In_210);
xnor U2128 (N_2128,In_1052,In_1927);
xor U2129 (N_2129,In_1507,In_1324);
or U2130 (N_2130,In_1411,In_1117);
xnor U2131 (N_2131,In_1917,In_1089);
and U2132 (N_2132,In_548,In_1261);
nor U2133 (N_2133,In_510,In_866);
xnor U2134 (N_2134,In_1938,In_1326);
nand U2135 (N_2135,In_340,In_1657);
nand U2136 (N_2136,In_1695,In_1664);
xor U2137 (N_2137,In_637,In_1958);
and U2138 (N_2138,In_792,In_503);
nor U2139 (N_2139,In_1014,In_364);
nor U2140 (N_2140,In_128,In_751);
nand U2141 (N_2141,In_1573,In_1291);
nand U2142 (N_2142,In_455,In_1840);
nor U2143 (N_2143,In_1469,In_273);
xnor U2144 (N_2144,In_397,In_942);
xor U2145 (N_2145,In_617,In_1281);
nor U2146 (N_2146,In_301,In_1584);
nand U2147 (N_2147,In_208,In_1019);
and U2148 (N_2148,In_437,In_252);
nor U2149 (N_2149,In_1948,In_840);
nand U2150 (N_2150,In_953,In_148);
xnor U2151 (N_2151,In_1694,In_150);
and U2152 (N_2152,In_197,In_1786);
nor U2153 (N_2153,In_4,In_282);
and U2154 (N_2154,In_1704,In_1738);
xnor U2155 (N_2155,In_740,In_878);
nor U2156 (N_2156,In_133,In_1914);
xor U2157 (N_2157,In_232,In_657);
and U2158 (N_2158,In_1076,In_1935);
or U2159 (N_2159,In_1957,In_1169);
xnor U2160 (N_2160,In_1658,In_239);
and U2161 (N_2161,In_504,In_1400);
nand U2162 (N_2162,In_550,In_1675);
nor U2163 (N_2163,In_13,In_40);
nand U2164 (N_2164,In_145,In_235);
xnor U2165 (N_2165,In_62,In_411);
nand U2166 (N_2166,In_1640,In_413);
nor U2167 (N_2167,In_1716,In_1200);
nor U2168 (N_2168,In_1813,In_649);
xor U2169 (N_2169,In_807,In_361);
nand U2170 (N_2170,In_1130,In_816);
nand U2171 (N_2171,In_1314,In_1237);
nor U2172 (N_2172,In_1907,In_1691);
xor U2173 (N_2173,In_61,In_1688);
nand U2174 (N_2174,In_1053,In_1227);
and U2175 (N_2175,In_1357,In_1293);
or U2176 (N_2176,In_941,In_997);
nand U2177 (N_2177,In_1442,In_1860);
nor U2178 (N_2178,In_957,In_454);
nand U2179 (N_2179,In_1355,In_52);
nor U2180 (N_2180,In_616,In_868);
xnor U2181 (N_2181,In_1148,In_750);
nand U2182 (N_2182,In_1192,In_1999);
nand U2183 (N_2183,In_10,In_198);
xor U2184 (N_2184,In_695,In_1886);
xnor U2185 (N_2185,In_1798,In_1234);
nor U2186 (N_2186,In_1931,In_434);
nor U2187 (N_2187,In_787,In_1487);
nor U2188 (N_2188,In_1534,In_1167);
or U2189 (N_2189,In_822,In_1919);
nor U2190 (N_2190,In_436,In_102);
xor U2191 (N_2191,In_467,In_1380);
nor U2192 (N_2192,In_422,In_78);
and U2193 (N_2193,In_1445,In_454);
or U2194 (N_2194,In_176,In_1604);
or U2195 (N_2195,In_1829,In_722);
nor U2196 (N_2196,In_802,In_491);
nor U2197 (N_2197,In_870,In_251);
xnor U2198 (N_2198,In_639,In_756);
nor U2199 (N_2199,In_693,In_1207);
and U2200 (N_2200,In_680,In_1426);
xor U2201 (N_2201,In_1641,In_1865);
nand U2202 (N_2202,In_1191,In_372);
nor U2203 (N_2203,In_341,In_784);
and U2204 (N_2204,In_598,In_1906);
nor U2205 (N_2205,In_1977,In_608);
or U2206 (N_2206,In_1956,In_1164);
and U2207 (N_2207,In_1235,In_437);
nor U2208 (N_2208,In_1200,In_669);
xnor U2209 (N_2209,In_1052,In_1424);
and U2210 (N_2210,In_1257,In_480);
nor U2211 (N_2211,In_445,In_1831);
xnor U2212 (N_2212,In_253,In_1977);
nand U2213 (N_2213,In_53,In_968);
nor U2214 (N_2214,In_615,In_444);
and U2215 (N_2215,In_1918,In_41);
nand U2216 (N_2216,In_36,In_1977);
nor U2217 (N_2217,In_226,In_1944);
nand U2218 (N_2218,In_1474,In_579);
or U2219 (N_2219,In_559,In_1170);
and U2220 (N_2220,In_80,In_460);
and U2221 (N_2221,In_1464,In_235);
nor U2222 (N_2222,In_1919,In_746);
nand U2223 (N_2223,In_1956,In_470);
or U2224 (N_2224,In_1067,In_469);
and U2225 (N_2225,In_1170,In_1849);
and U2226 (N_2226,In_760,In_1765);
nor U2227 (N_2227,In_781,In_1153);
or U2228 (N_2228,In_270,In_1312);
nand U2229 (N_2229,In_1171,In_421);
or U2230 (N_2230,In_1977,In_1611);
xor U2231 (N_2231,In_257,In_417);
and U2232 (N_2232,In_365,In_113);
xnor U2233 (N_2233,In_530,In_1458);
nor U2234 (N_2234,In_1664,In_1650);
nor U2235 (N_2235,In_1631,In_68);
nand U2236 (N_2236,In_1275,In_417);
xnor U2237 (N_2237,In_487,In_127);
and U2238 (N_2238,In_1588,In_848);
or U2239 (N_2239,In_1169,In_514);
and U2240 (N_2240,In_1071,In_404);
nor U2241 (N_2241,In_1880,In_1098);
nand U2242 (N_2242,In_913,In_1743);
nor U2243 (N_2243,In_1984,In_1543);
or U2244 (N_2244,In_901,In_1323);
nor U2245 (N_2245,In_576,In_1721);
nand U2246 (N_2246,In_172,In_1891);
or U2247 (N_2247,In_1563,In_1438);
nand U2248 (N_2248,In_787,In_1125);
and U2249 (N_2249,In_934,In_913);
nor U2250 (N_2250,In_5,In_821);
or U2251 (N_2251,In_1547,In_1856);
or U2252 (N_2252,In_1704,In_402);
or U2253 (N_2253,In_753,In_1325);
nor U2254 (N_2254,In_1631,In_194);
and U2255 (N_2255,In_1289,In_1457);
and U2256 (N_2256,In_549,In_882);
nand U2257 (N_2257,In_1536,In_1917);
xnor U2258 (N_2258,In_748,In_429);
or U2259 (N_2259,In_1081,In_1783);
nand U2260 (N_2260,In_507,In_477);
and U2261 (N_2261,In_952,In_136);
nand U2262 (N_2262,In_1392,In_385);
nor U2263 (N_2263,In_112,In_1768);
xnor U2264 (N_2264,In_1556,In_1408);
or U2265 (N_2265,In_851,In_635);
nand U2266 (N_2266,In_627,In_1948);
and U2267 (N_2267,In_311,In_1457);
or U2268 (N_2268,In_1267,In_20);
or U2269 (N_2269,In_1750,In_763);
xnor U2270 (N_2270,In_1439,In_1953);
or U2271 (N_2271,In_56,In_1171);
nand U2272 (N_2272,In_755,In_237);
nand U2273 (N_2273,In_1197,In_1041);
and U2274 (N_2274,In_1861,In_1361);
nor U2275 (N_2275,In_1517,In_1816);
xnor U2276 (N_2276,In_688,In_560);
or U2277 (N_2277,In_930,In_1227);
and U2278 (N_2278,In_1328,In_1055);
or U2279 (N_2279,In_210,In_269);
nor U2280 (N_2280,In_1064,In_130);
xnor U2281 (N_2281,In_104,In_380);
or U2282 (N_2282,In_551,In_20);
xor U2283 (N_2283,In_657,In_775);
and U2284 (N_2284,In_882,In_1717);
and U2285 (N_2285,In_284,In_1010);
or U2286 (N_2286,In_1453,In_1436);
xnor U2287 (N_2287,In_1565,In_1018);
xnor U2288 (N_2288,In_823,In_380);
nand U2289 (N_2289,In_169,In_496);
or U2290 (N_2290,In_494,In_558);
and U2291 (N_2291,In_368,In_1436);
or U2292 (N_2292,In_1008,In_1984);
and U2293 (N_2293,In_1132,In_1316);
and U2294 (N_2294,In_263,In_711);
nand U2295 (N_2295,In_114,In_996);
xor U2296 (N_2296,In_130,In_1006);
nor U2297 (N_2297,In_468,In_1921);
or U2298 (N_2298,In_281,In_1507);
nor U2299 (N_2299,In_827,In_630);
or U2300 (N_2300,In_1079,In_726);
xor U2301 (N_2301,In_1359,In_1954);
xor U2302 (N_2302,In_1410,In_379);
nor U2303 (N_2303,In_689,In_1599);
nand U2304 (N_2304,In_864,In_868);
and U2305 (N_2305,In_701,In_1323);
or U2306 (N_2306,In_1855,In_979);
nor U2307 (N_2307,In_1571,In_1280);
and U2308 (N_2308,In_1284,In_390);
nor U2309 (N_2309,In_100,In_453);
nor U2310 (N_2310,In_96,In_1314);
nand U2311 (N_2311,In_1578,In_316);
and U2312 (N_2312,In_1075,In_1938);
nand U2313 (N_2313,In_1221,In_1147);
nor U2314 (N_2314,In_28,In_1233);
xor U2315 (N_2315,In_1921,In_1086);
xnor U2316 (N_2316,In_1854,In_16);
nor U2317 (N_2317,In_1194,In_1595);
and U2318 (N_2318,In_591,In_1607);
or U2319 (N_2319,In_420,In_1578);
nor U2320 (N_2320,In_1552,In_533);
or U2321 (N_2321,In_1888,In_806);
xor U2322 (N_2322,In_1946,In_1157);
nand U2323 (N_2323,In_1862,In_1334);
or U2324 (N_2324,In_382,In_363);
xor U2325 (N_2325,In_1952,In_907);
nor U2326 (N_2326,In_1498,In_1321);
nor U2327 (N_2327,In_1706,In_1479);
xnor U2328 (N_2328,In_1246,In_858);
nand U2329 (N_2329,In_1047,In_910);
or U2330 (N_2330,In_1820,In_1574);
and U2331 (N_2331,In_506,In_1763);
nor U2332 (N_2332,In_1242,In_1510);
xnor U2333 (N_2333,In_1243,In_986);
nor U2334 (N_2334,In_1244,In_1610);
or U2335 (N_2335,In_227,In_1911);
nor U2336 (N_2336,In_373,In_1643);
nor U2337 (N_2337,In_622,In_1379);
xor U2338 (N_2338,In_849,In_171);
nor U2339 (N_2339,In_659,In_260);
or U2340 (N_2340,In_723,In_151);
or U2341 (N_2341,In_1312,In_801);
nand U2342 (N_2342,In_1081,In_721);
or U2343 (N_2343,In_1751,In_1632);
or U2344 (N_2344,In_1996,In_367);
xnor U2345 (N_2345,In_812,In_595);
or U2346 (N_2346,In_140,In_369);
xnor U2347 (N_2347,In_1028,In_1399);
xnor U2348 (N_2348,In_1655,In_951);
or U2349 (N_2349,In_1252,In_352);
nor U2350 (N_2350,In_1697,In_1488);
xnor U2351 (N_2351,In_1830,In_1505);
nand U2352 (N_2352,In_498,In_1208);
or U2353 (N_2353,In_905,In_1551);
or U2354 (N_2354,In_1411,In_114);
xnor U2355 (N_2355,In_386,In_570);
and U2356 (N_2356,In_748,In_191);
xnor U2357 (N_2357,In_198,In_1307);
or U2358 (N_2358,In_1723,In_1091);
or U2359 (N_2359,In_1347,In_1135);
nor U2360 (N_2360,In_85,In_520);
and U2361 (N_2361,In_83,In_856);
xor U2362 (N_2362,In_1739,In_1052);
nor U2363 (N_2363,In_659,In_794);
or U2364 (N_2364,In_1771,In_1215);
xnor U2365 (N_2365,In_124,In_1223);
and U2366 (N_2366,In_252,In_45);
nor U2367 (N_2367,In_599,In_462);
and U2368 (N_2368,In_1329,In_791);
and U2369 (N_2369,In_1452,In_524);
and U2370 (N_2370,In_1875,In_252);
or U2371 (N_2371,In_1128,In_1107);
xnor U2372 (N_2372,In_1811,In_780);
or U2373 (N_2373,In_1611,In_915);
and U2374 (N_2374,In_1538,In_133);
and U2375 (N_2375,In_1968,In_11);
nor U2376 (N_2376,In_1905,In_1445);
or U2377 (N_2377,In_567,In_800);
or U2378 (N_2378,In_1509,In_1141);
nor U2379 (N_2379,In_565,In_1963);
and U2380 (N_2380,In_104,In_539);
and U2381 (N_2381,In_232,In_499);
and U2382 (N_2382,In_1381,In_864);
xor U2383 (N_2383,In_1429,In_601);
nand U2384 (N_2384,In_227,In_992);
and U2385 (N_2385,In_1791,In_833);
nand U2386 (N_2386,In_1067,In_1428);
and U2387 (N_2387,In_622,In_1615);
nand U2388 (N_2388,In_1980,In_722);
or U2389 (N_2389,In_1643,In_31);
nor U2390 (N_2390,In_101,In_1568);
and U2391 (N_2391,In_1331,In_481);
and U2392 (N_2392,In_842,In_1871);
nor U2393 (N_2393,In_524,In_1642);
xor U2394 (N_2394,In_1011,In_810);
xnor U2395 (N_2395,In_1901,In_1699);
xor U2396 (N_2396,In_1834,In_146);
xor U2397 (N_2397,In_239,In_1727);
nor U2398 (N_2398,In_1410,In_1906);
or U2399 (N_2399,In_1249,In_114);
or U2400 (N_2400,In_1283,In_1931);
or U2401 (N_2401,In_1488,In_1113);
or U2402 (N_2402,In_81,In_1925);
xor U2403 (N_2403,In_1544,In_1983);
or U2404 (N_2404,In_1921,In_1911);
nor U2405 (N_2405,In_935,In_58);
nor U2406 (N_2406,In_1378,In_1698);
xnor U2407 (N_2407,In_1277,In_1362);
xnor U2408 (N_2408,In_1360,In_1377);
nor U2409 (N_2409,In_430,In_790);
and U2410 (N_2410,In_822,In_798);
nand U2411 (N_2411,In_182,In_1332);
nand U2412 (N_2412,In_1005,In_1684);
nor U2413 (N_2413,In_59,In_1205);
nor U2414 (N_2414,In_919,In_1192);
xor U2415 (N_2415,In_1019,In_800);
nand U2416 (N_2416,In_1524,In_9);
xnor U2417 (N_2417,In_594,In_868);
xnor U2418 (N_2418,In_1532,In_1133);
xnor U2419 (N_2419,In_1065,In_860);
or U2420 (N_2420,In_1872,In_1954);
nor U2421 (N_2421,In_33,In_762);
and U2422 (N_2422,In_785,In_1142);
or U2423 (N_2423,In_1110,In_480);
nand U2424 (N_2424,In_1539,In_1991);
and U2425 (N_2425,In_1591,In_1741);
and U2426 (N_2426,In_337,In_677);
nand U2427 (N_2427,In_676,In_374);
xor U2428 (N_2428,In_824,In_764);
nand U2429 (N_2429,In_1894,In_207);
xnor U2430 (N_2430,In_1138,In_384);
or U2431 (N_2431,In_327,In_1962);
nor U2432 (N_2432,In_1653,In_540);
or U2433 (N_2433,In_1084,In_1677);
and U2434 (N_2434,In_104,In_1665);
and U2435 (N_2435,In_60,In_1194);
nor U2436 (N_2436,In_444,In_1736);
nor U2437 (N_2437,In_770,In_1092);
or U2438 (N_2438,In_1937,In_325);
xnor U2439 (N_2439,In_1646,In_1787);
or U2440 (N_2440,In_24,In_198);
nor U2441 (N_2441,In_1391,In_1109);
nor U2442 (N_2442,In_192,In_1554);
nor U2443 (N_2443,In_1300,In_1426);
xnor U2444 (N_2444,In_193,In_352);
or U2445 (N_2445,In_524,In_923);
nor U2446 (N_2446,In_1734,In_1670);
xnor U2447 (N_2447,In_1865,In_1165);
or U2448 (N_2448,In_369,In_1655);
xnor U2449 (N_2449,In_1682,In_1022);
or U2450 (N_2450,In_1564,In_892);
xor U2451 (N_2451,In_1691,In_415);
and U2452 (N_2452,In_1658,In_1562);
nand U2453 (N_2453,In_48,In_1200);
or U2454 (N_2454,In_321,In_1946);
and U2455 (N_2455,In_3,In_1627);
or U2456 (N_2456,In_1062,In_217);
and U2457 (N_2457,In_396,In_683);
nor U2458 (N_2458,In_500,In_317);
and U2459 (N_2459,In_1795,In_805);
nor U2460 (N_2460,In_428,In_340);
or U2461 (N_2461,In_1949,In_103);
nor U2462 (N_2462,In_1212,In_35);
xor U2463 (N_2463,In_567,In_1207);
and U2464 (N_2464,In_975,In_1015);
or U2465 (N_2465,In_222,In_498);
nor U2466 (N_2466,In_1250,In_1987);
or U2467 (N_2467,In_370,In_203);
or U2468 (N_2468,In_790,In_540);
nand U2469 (N_2469,In_1951,In_1286);
nand U2470 (N_2470,In_1184,In_1104);
xor U2471 (N_2471,In_119,In_1016);
nor U2472 (N_2472,In_42,In_1993);
nor U2473 (N_2473,In_1140,In_679);
nand U2474 (N_2474,In_585,In_1893);
xor U2475 (N_2475,In_135,In_1330);
or U2476 (N_2476,In_1899,In_823);
nand U2477 (N_2477,In_911,In_99);
and U2478 (N_2478,In_1240,In_1934);
nand U2479 (N_2479,In_1409,In_1369);
nor U2480 (N_2480,In_379,In_1463);
or U2481 (N_2481,In_1098,In_757);
or U2482 (N_2482,In_33,In_1994);
or U2483 (N_2483,In_859,In_665);
xnor U2484 (N_2484,In_1079,In_278);
and U2485 (N_2485,In_42,In_1802);
xor U2486 (N_2486,In_1742,In_1203);
and U2487 (N_2487,In_1006,In_1978);
nor U2488 (N_2488,In_829,In_520);
nor U2489 (N_2489,In_949,In_108);
nor U2490 (N_2490,In_55,In_509);
nor U2491 (N_2491,In_66,In_1066);
nand U2492 (N_2492,In_394,In_1900);
nand U2493 (N_2493,In_172,In_1934);
and U2494 (N_2494,In_1263,In_1775);
nand U2495 (N_2495,In_1581,In_41);
or U2496 (N_2496,In_665,In_949);
nand U2497 (N_2497,In_1998,In_1089);
or U2498 (N_2498,In_455,In_779);
or U2499 (N_2499,In_1364,In_475);
nand U2500 (N_2500,In_1758,In_1165);
and U2501 (N_2501,In_83,In_1639);
nand U2502 (N_2502,In_661,In_1365);
xnor U2503 (N_2503,In_737,In_684);
xor U2504 (N_2504,In_1865,In_1596);
or U2505 (N_2505,In_369,In_1057);
nor U2506 (N_2506,In_1168,In_688);
xnor U2507 (N_2507,In_937,In_316);
nor U2508 (N_2508,In_1478,In_245);
xor U2509 (N_2509,In_1719,In_612);
nand U2510 (N_2510,In_1010,In_761);
nor U2511 (N_2511,In_910,In_226);
xor U2512 (N_2512,In_429,In_1640);
and U2513 (N_2513,In_1699,In_1312);
and U2514 (N_2514,In_1019,In_1532);
or U2515 (N_2515,In_712,In_809);
and U2516 (N_2516,In_1570,In_624);
and U2517 (N_2517,In_1519,In_198);
xnor U2518 (N_2518,In_881,In_677);
nor U2519 (N_2519,In_483,In_1312);
and U2520 (N_2520,In_1236,In_463);
and U2521 (N_2521,In_1030,In_1270);
nand U2522 (N_2522,In_66,In_1363);
and U2523 (N_2523,In_528,In_1780);
nor U2524 (N_2524,In_1876,In_146);
nor U2525 (N_2525,In_447,In_889);
xnor U2526 (N_2526,In_1774,In_1067);
nor U2527 (N_2527,In_559,In_746);
nand U2528 (N_2528,In_1018,In_462);
nor U2529 (N_2529,In_245,In_1989);
nand U2530 (N_2530,In_428,In_1356);
nand U2531 (N_2531,In_1473,In_417);
or U2532 (N_2532,In_1692,In_1025);
and U2533 (N_2533,In_1873,In_1937);
or U2534 (N_2534,In_1420,In_1990);
xor U2535 (N_2535,In_777,In_844);
nand U2536 (N_2536,In_1906,In_536);
xor U2537 (N_2537,In_738,In_1585);
and U2538 (N_2538,In_338,In_1732);
or U2539 (N_2539,In_1742,In_1262);
nand U2540 (N_2540,In_1493,In_1027);
or U2541 (N_2541,In_907,In_1419);
nand U2542 (N_2542,In_431,In_1940);
or U2543 (N_2543,In_163,In_1552);
xnor U2544 (N_2544,In_1209,In_517);
xnor U2545 (N_2545,In_1738,In_50);
and U2546 (N_2546,In_1048,In_715);
xnor U2547 (N_2547,In_555,In_1619);
xor U2548 (N_2548,In_1461,In_1583);
or U2549 (N_2549,In_662,In_1348);
and U2550 (N_2550,In_633,In_835);
or U2551 (N_2551,In_785,In_1856);
nand U2552 (N_2552,In_520,In_739);
or U2553 (N_2553,In_550,In_291);
xnor U2554 (N_2554,In_28,In_1417);
nand U2555 (N_2555,In_74,In_948);
nand U2556 (N_2556,In_16,In_944);
or U2557 (N_2557,In_1308,In_1564);
and U2558 (N_2558,In_1403,In_1540);
and U2559 (N_2559,In_1461,In_1233);
and U2560 (N_2560,In_1439,In_1191);
or U2561 (N_2561,In_512,In_576);
nor U2562 (N_2562,In_1594,In_947);
xnor U2563 (N_2563,In_1686,In_244);
nand U2564 (N_2564,In_252,In_1424);
nor U2565 (N_2565,In_667,In_1421);
nor U2566 (N_2566,In_1530,In_359);
xor U2567 (N_2567,In_788,In_465);
xor U2568 (N_2568,In_1009,In_1236);
nand U2569 (N_2569,In_690,In_1798);
xor U2570 (N_2570,In_1096,In_1011);
xor U2571 (N_2571,In_1229,In_1801);
nand U2572 (N_2572,In_1323,In_1545);
nor U2573 (N_2573,In_578,In_724);
nor U2574 (N_2574,In_1374,In_1678);
nor U2575 (N_2575,In_1355,In_257);
or U2576 (N_2576,In_1744,In_1456);
and U2577 (N_2577,In_311,In_845);
or U2578 (N_2578,In_418,In_1332);
nand U2579 (N_2579,In_1891,In_1401);
nor U2580 (N_2580,In_973,In_1675);
or U2581 (N_2581,In_169,In_129);
nor U2582 (N_2582,In_919,In_1345);
nor U2583 (N_2583,In_35,In_1885);
nand U2584 (N_2584,In_286,In_954);
nor U2585 (N_2585,In_479,In_592);
or U2586 (N_2586,In_1108,In_1526);
nand U2587 (N_2587,In_1105,In_306);
nand U2588 (N_2588,In_945,In_673);
xnor U2589 (N_2589,In_1571,In_59);
nor U2590 (N_2590,In_784,In_794);
nor U2591 (N_2591,In_923,In_1464);
xnor U2592 (N_2592,In_691,In_283);
nand U2593 (N_2593,In_1815,In_1534);
or U2594 (N_2594,In_122,In_1929);
and U2595 (N_2595,In_146,In_214);
nor U2596 (N_2596,In_378,In_7);
xor U2597 (N_2597,In_56,In_1700);
xor U2598 (N_2598,In_1532,In_1804);
or U2599 (N_2599,In_715,In_183);
or U2600 (N_2600,In_1414,In_388);
xor U2601 (N_2601,In_6,In_1535);
or U2602 (N_2602,In_774,In_890);
and U2603 (N_2603,In_1891,In_576);
and U2604 (N_2604,In_1696,In_1204);
xor U2605 (N_2605,In_402,In_11);
xnor U2606 (N_2606,In_124,In_56);
xor U2607 (N_2607,In_1336,In_446);
or U2608 (N_2608,In_810,In_1603);
or U2609 (N_2609,In_175,In_1654);
nand U2610 (N_2610,In_877,In_725);
and U2611 (N_2611,In_1073,In_55);
xor U2612 (N_2612,In_1377,In_1412);
nor U2613 (N_2613,In_1660,In_495);
and U2614 (N_2614,In_1082,In_1782);
xor U2615 (N_2615,In_1677,In_1188);
nand U2616 (N_2616,In_1575,In_7);
or U2617 (N_2617,In_1640,In_46);
and U2618 (N_2618,In_1695,In_1388);
nor U2619 (N_2619,In_878,In_978);
and U2620 (N_2620,In_1834,In_962);
or U2621 (N_2621,In_658,In_481);
nor U2622 (N_2622,In_857,In_337);
and U2623 (N_2623,In_1083,In_964);
xor U2624 (N_2624,In_984,In_1439);
or U2625 (N_2625,In_1958,In_1809);
or U2626 (N_2626,In_1876,In_719);
nor U2627 (N_2627,In_207,In_1493);
nor U2628 (N_2628,In_18,In_516);
or U2629 (N_2629,In_1210,In_1697);
or U2630 (N_2630,In_1805,In_923);
nor U2631 (N_2631,In_875,In_1224);
nor U2632 (N_2632,In_1400,In_755);
or U2633 (N_2633,In_793,In_631);
nor U2634 (N_2634,In_1308,In_1715);
and U2635 (N_2635,In_192,In_203);
nor U2636 (N_2636,In_160,In_789);
nand U2637 (N_2637,In_293,In_1957);
and U2638 (N_2638,In_1060,In_1154);
nor U2639 (N_2639,In_1176,In_1855);
xor U2640 (N_2640,In_819,In_155);
and U2641 (N_2641,In_377,In_841);
xnor U2642 (N_2642,In_1407,In_1931);
or U2643 (N_2643,In_1031,In_1993);
or U2644 (N_2644,In_29,In_711);
nand U2645 (N_2645,In_1445,In_1051);
and U2646 (N_2646,In_984,In_1571);
nand U2647 (N_2647,In_47,In_272);
and U2648 (N_2648,In_1691,In_425);
nor U2649 (N_2649,In_438,In_1384);
nor U2650 (N_2650,In_403,In_1350);
nor U2651 (N_2651,In_67,In_1457);
nor U2652 (N_2652,In_273,In_1704);
and U2653 (N_2653,In_1211,In_1251);
nor U2654 (N_2654,In_1484,In_1784);
xnor U2655 (N_2655,In_1009,In_247);
and U2656 (N_2656,In_733,In_1800);
and U2657 (N_2657,In_356,In_1447);
and U2658 (N_2658,In_1852,In_1643);
or U2659 (N_2659,In_1770,In_1897);
xor U2660 (N_2660,In_1530,In_808);
nand U2661 (N_2661,In_844,In_1106);
nor U2662 (N_2662,In_898,In_782);
or U2663 (N_2663,In_1187,In_1197);
xor U2664 (N_2664,In_1927,In_280);
or U2665 (N_2665,In_1658,In_296);
nand U2666 (N_2666,In_441,In_1673);
or U2667 (N_2667,In_1100,In_1826);
and U2668 (N_2668,In_1365,In_1919);
and U2669 (N_2669,In_1192,In_734);
nor U2670 (N_2670,In_1500,In_21);
nor U2671 (N_2671,In_667,In_829);
nor U2672 (N_2672,In_380,In_582);
and U2673 (N_2673,In_492,In_581);
xor U2674 (N_2674,In_138,In_470);
or U2675 (N_2675,In_474,In_891);
nor U2676 (N_2676,In_244,In_1863);
nand U2677 (N_2677,In_260,In_918);
or U2678 (N_2678,In_1371,In_1937);
nand U2679 (N_2679,In_1286,In_1877);
nand U2680 (N_2680,In_35,In_1011);
and U2681 (N_2681,In_380,In_1353);
xnor U2682 (N_2682,In_953,In_1777);
and U2683 (N_2683,In_576,In_495);
xnor U2684 (N_2684,In_1686,In_558);
or U2685 (N_2685,In_969,In_110);
and U2686 (N_2686,In_823,In_638);
nor U2687 (N_2687,In_551,In_1777);
nor U2688 (N_2688,In_1024,In_917);
or U2689 (N_2689,In_85,In_113);
or U2690 (N_2690,In_1624,In_1243);
nand U2691 (N_2691,In_496,In_1240);
or U2692 (N_2692,In_1854,In_809);
nor U2693 (N_2693,In_382,In_1255);
nand U2694 (N_2694,In_1486,In_668);
and U2695 (N_2695,In_220,In_1680);
nand U2696 (N_2696,In_625,In_1303);
or U2697 (N_2697,In_1888,In_355);
nand U2698 (N_2698,In_1294,In_1991);
nor U2699 (N_2699,In_876,In_912);
nor U2700 (N_2700,In_1956,In_920);
nor U2701 (N_2701,In_885,In_185);
nor U2702 (N_2702,In_1007,In_1785);
and U2703 (N_2703,In_706,In_877);
nand U2704 (N_2704,In_1667,In_647);
or U2705 (N_2705,In_329,In_1819);
xor U2706 (N_2706,In_970,In_295);
nand U2707 (N_2707,In_342,In_887);
and U2708 (N_2708,In_10,In_1734);
and U2709 (N_2709,In_471,In_1573);
nor U2710 (N_2710,In_1972,In_1234);
and U2711 (N_2711,In_1639,In_1703);
nand U2712 (N_2712,In_1468,In_406);
nor U2713 (N_2713,In_239,In_645);
nor U2714 (N_2714,In_1199,In_599);
nor U2715 (N_2715,In_508,In_1281);
or U2716 (N_2716,In_1855,In_1090);
and U2717 (N_2717,In_1853,In_1605);
nor U2718 (N_2718,In_529,In_1297);
or U2719 (N_2719,In_1460,In_1822);
nor U2720 (N_2720,In_1882,In_428);
or U2721 (N_2721,In_1245,In_1095);
nand U2722 (N_2722,In_59,In_1775);
nor U2723 (N_2723,In_1305,In_1469);
nor U2724 (N_2724,In_983,In_807);
nand U2725 (N_2725,In_1199,In_576);
nor U2726 (N_2726,In_81,In_628);
nor U2727 (N_2727,In_1550,In_1326);
and U2728 (N_2728,In_1033,In_574);
nand U2729 (N_2729,In_1109,In_89);
nand U2730 (N_2730,In_372,In_1325);
or U2731 (N_2731,In_729,In_947);
nor U2732 (N_2732,In_683,In_1508);
nor U2733 (N_2733,In_1136,In_1780);
or U2734 (N_2734,In_1247,In_1487);
nor U2735 (N_2735,In_1775,In_79);
xnor U2736 (N_2736,In_436,In_659);
nand U2737 (N_2737,In_1108,In_971);
xor U2738 (N_2738,In_590,In_105);
nand U2739 (N_2739,In_1138,In_797);
xnor U2740 (N_2740,In_228,In_1873);
or U2741 (N_2741,In_953,In_104);
xor U2742 (N_2742,In_1436,In_672);
nor U2743 (N_2743,In_697,In_1177);
xnor U2744 (N_2744,In_282,In_580);
or U2745 (N_2745,In_1978,In_714);
and U2746 (N_2746,In_262,In_1987);
nor U2747 (N_2747,In_36,In_41);
nand U2748 (N_2748,In_345,In_1743);
nand U2749 (N_2749,In_642,In_507);
nor U2750 (N_2750,In_208,In_1679);
and U2751 (N_2751,In_449,In_532);
or U2752 (N_2752,In_152,In_931);
nand U2753 (N_2753,In_306,In_1951);
or U2754 (N_2754,In_557,In_1537);
nor U2755 (N_2755,In_1803,In_209);
or U2756 (N_2756,In_1223,In_19);
xor U2757 (N_2757,In_313,In_162);
nand U2758 (N_2758,In_1734,In_435);
or U2759 (N_2759,In_1721,In_335);
and U2760 (N_2760,In_1955,In_353);
or U2761 (N_2761,In_796,In_722);
nand U2762 (N_2762,In_1518,In_1106);
and U2763 (N_2763,In_1705,In_61);
xor U2764 (N_2764,In_1181,In_1040);
nor U2765 (N_2765,In_743,In_171);
nor U2766 (N_2766,In_303,In_2);
nand U2767 (N_2767,In_716,In_1457);
nand U2768 (N_2768,In_1433,In_758);
and U2769 (N_2769,In_1770,In_1939);
nand U2770 (N_2770,In_552,In_1967);
or U2771 (N_2771,In_512,In_1267);
nor U2772 (N_2772,In_1727,In_512);
nand U2773 (N_2773,In_1228,In_1343);
xnor U2774 (N_2774,In_222,In_1939);
xor U2775 (N_2775,In_772,In_521);
xnor U2776 (N_2776,In_1526,In_1762);
xor U2777 (N_2777,In_843,In_1193);
nand U2778 (N_2778,In_620,In_625);
or U2779 (N_2779,In_1956,In_1037);
nand U2780 (N_2780,In_1483,In_941);
nor U2781 (N_2781,In_964,In_1216);
and U2782 (N_2782,In_1641,In_1625);
nor U2783 (N_2783,In_327,In_1321);
nor U2784 (N_2784,In_970,In_844);
xor U2785 (N_2785,In_1523,In_1503);
or U2786 (N_2786,In_979,In_1534);
and U2787 (N_2787,In_828,In_1094);
nor U2788 (N_2788,In_1891,In_1369);
or U2789 (N_2789,In_617,In_1284);
or U2790 (N_2790,In_215,In_807);
and U2791 (N_2791,In_632,In_1205);
xor U2792 (N_2792,In_1797,In_1465);
or U2793 (N_2793,In_1489,In_1822);
or U2794 (N_2794,In_43,In_428);
xnor U2795 (N_2795,In_1758,In_1414);
or U2796 (N_2796,In_1248,In_1941);
xnor U2797 (N_2797,In_459,In_1119);
nand U2798 (N_2798,In_13,In_1229);
nand U2799 (N_2799,In_1860,In_1536);
or U2800 (N_2800,In_1297,In_140);
nand U2801 (N_2801,In_1382,In_839);
and U2802 (N_2802,In_1143,In_1379);
and U2803 (N_2803,In_1282,In_328);
nor U2804 (N_2804,In_976,In_1927);
xor U2805 (N_2805,In_659,In_625);
or U2806 (N_2806,In_987,In_15);
nand U2807 (N_2807,In_1957,In_989);
nand U2808 (N_2808,In_948,In_525);
and U2809 (N_2809,In_1385,In_1066);
or U2810 (N_2810,In_456,In_861);
nor U2811 (N_2811,In_914,In_540);
nor U2812 (N_2812,In_779,In_1996);
xor U2813 (N_2813,In_312,In_1518);
and U2814 (N_2814,In_1925,In_334);
or U2815 (N_2815,In_318,In_1446);
or U2816 (N_2816,In_1357,In_692);
nor U2817 (N_2817,In_1978,In_1971);
xor U2818 (N_2818,In_451,In_591);
nand U2819 (N_2819,In_840,In_1396);
nand U2820 (N_2820,In_1389,In_575);
xor U2821 (N_2821,In_1820,In_685);
xor U2822 (N_2822,In_1301,In_1069);
xnor U2823 (N_2823,In_1539,In_1505);
nor U2824 (N_2824,In_577,In_7);
and U2825 (N_2825,In_155,In_502);
nor U2826 (N_2826,In_1448,In_1703);
xnor U2827 (N_2827,In_713,In_1090);
nor U2828 (N_2828,In_289,In_617);
nor U2829 (N_2829,In_841,In_1595);
xor U2830 (N_2830,In_1221,In_211);
nor U2831 (N_2831,In_1281,In_832);
xor U2832 (N_2832,In_682,In_988);
nor U2833 (N_2833,In_1932,In_59);
xnor U2834 (N_2834,In_1592,In_1466);
or U2835 (N_2835,In_1325,In_1032);
or U2836 (N_2836,In_938,In_992);
or U2837 (N_2837,In_1179,In_1334);
nor U2838 (N_2838,In_1541,In_1743);
and U2839 (N_2839,In_1207,In_785);
or U2840 (N_2840,In_500,In_543);
nor U2841 (N_2841,In_1491,In_994);
nand U2842 (N_2842,In_1831,In_103);
and U2843 (N_2843,In_1365,In_807);
and U2844 (N_2844,In_1641,In_569);
xor U2845 (N_2845,In_1047,In_241);
xor U2846 (N_2846,In_431,In_837);
xnor U2847 (N_2847,In_1341,In_419);
or U2848 (N_2848,In_1697,In_1782);
nand U2849 (N_2849,In_1226,In_518);
and U2850 (N_2850,In_1401,In_175);
or U2851 (N_2851,In_206,In_1362);
or U2852 (N_2852,In_1172,In_1343);
nor U2853 (N_2853,In_1683,In_1524);
nand U2854 (N_2854,In_1473,In_1405);
xnor U2855 (N_2855,In_551,In_1417);
or U2856 (N_2856,In_235,In_1095);
or U2857 (N_2857,In_942,In_237);
xor U2858 (N_2858,In_370,In_1303);
xor U2859 (N_2859,In_455,In_220);
and U2860 (N_2860,In_446,In_228);
nor U2861 (N_2861,In_212,In_1920);
nand U2862 (N_2862,In_58,In_1112);
and U2863 (N_2863,In_1348,In_873);
or U2864 (N_2864,In_404,In_1483);
xnor U2865 (N_2865,In_313,In_1587);
nor U2866 (N_2866,In_706,In_1973);
nand U2867 (N_2867,In_90,In_337);
xnor U2868 (N_2868,In_595,In_938);
and U2869 (N_2869,In_211,In_108);
nor U2870 (N_2870,In_394,In_1107);
nand U2871 (N_2871,In_841,In_1525);
and U2872 (N_2872,In_1481,In_217);
and U2873 (N_2873,In_687,In_1979);
xor U2874 (N_2874,In_966,In_898);
xor U2875 (N_2875,In_310,In_105);
xor U2876 (N_2876,In_401,In_1370);
or U2877 (N_2877,In_590,In_892);
nand U2878 (N_2878,In_1328,In_336);
nand U2879 (N_2879,In_1615,In_1923);
or U2880 (N_2880,In_756,In_518);
nand U2881 (N_2881,In_702,In_1439);
nand U2882 (N_2882,In_579,In_1375);
or U2883 (N_2883,In_525,In_622);
nor U2884 (N_2884,In_787,In_85);
or U2885 (N_2885,In_1707,In_1225);
and U2886 (N_2886,In_412,In_803);
nor U2887 (N_2887,In_107,In_166);
nand U2888 (N_2888,In_1698,In_1260);
xnor U2889 (N_2889,In_567,In_1238);
nand U2890 (N_2890,In_422,In_807);
and U2891 (N_2891,In_231,In_946);
nand U2892 (N_2892,In_456,In_1019);
nor U2893 (N_2893,In_149,In_866);
or U2894 (N_2894,In_1855,In_1519);
and U2895 (N_2895,In_1877,In_1946);
and U2896 (N_2896,In_1434,In_1288);
xor U2897 (N_2897,In_1550,In_1467);
and U2898 (N_2898,In_1557,In_16);
nand U2899 (N_2899,In_1794,In_158);
xnor U2900 (N_2900,In_1988,In_935);
nor U2901 (N_2901,In_279,In_295);
nand U2902 (N_2902,In_215,In_1772);
nand U2903 (N_2903,In_392,In_790);
and U2904 (N_2904,In_284,In_1699);
and U2905 (N_2905,In_691,In_1384);
nor U2906 (N_2906,In_1849,In_1106);
xnor U2907 (N_2907,In_144,In_1342);
xnor U2908 (N_2908,In_482,In_908);
nand U2909 (N_2909,In_166,In_1031);
or U2910 (N_2910,In_1235,In_451);
xor U2911 (N_2911,In_624,In_902);
nor U2912 (N_2912,In_1453,In_1841);
nor U2913 (N_2913,In_1130,In_1811);
xor U2914 (N_2914,In_286,In_327);
nand U2915 (N_2915,In_285,In_1834);
nor U2916 (N_2916,In_1467,In_1792);
nor U2917 (N_2917,In_1170,In_1356);
xor U2918 (N_2918,In_1991,In_1096);
or U2919 (N_2919,In_552,In_1586);
nor U2920 (N_2920,In_491,In_452);
and U2921 (N_2921,In_1049,In_1973);
or U2922 (N_2922,In_117,In_603);
xor U2923 (N_2923,In_442,In_1281);
nand U2924 (N_2924,In_456,In_33);
xnor U2925 (N_2925,In_1956,In_142);
and U2926 (N_2926,In_283,In_897);
xnor U2927 (N_2927,In_628,In_1730);
nor U2928 (N_2928,In_435,In_70);
or U2929 (N_2929,In_1138,In_1652);
and U2930 (N_2930,In_1731,In_1919);
xnor U2931 (N_2931,In_328,In_1550);
nand U2932 (N_2932,In_1935,In_305);
xnor U2933 (N_2933,In_1207,In_263);
nor U2934 (N_2934,In_833,In_1851);
nand U2935 (N_2935,In_329,In_1129);
and U2936 (N_2936,In_594,In_436);
nand U2937 (N_2937,In_571,In_930);
nand U2938 (N_2938,In_1148,In_510);
nand U2939 (N_2939,In_1129,In_1429);
nand U2940 (N_2940,In_421,In_1173);
and U2941 (N_2941,In_633,In_296);
or U2942 (N_2942,In_331,In_1971);
nor U2943 (N_2943,In_775,In_1749);
and U2944 (N_2944,In_1638,In_818);
nand U2945 (N_2945,In_1722,In_1327);
nor U2946 (N_2946,In_1225,In_1537);
nand U2947 (N_2947,In_1070,In_1822);
nor U2948 (N_2948,In_1025,In_1157);
nor U2949 (N_2949,In_1534,In_1464);
and U2950 (N_2950,In_37,In_499);
nand U2951 (N_2951,In_148,In_1019);
and U2952 (N_2952,In_735,In_1151);
nand U2953 (N_2953,In_281,In_778);
nor U2954 (N_2954,In_1796,In_796);
or U2955 (N_2955,In_1662,In_1044);
or U2956 (N_2956,In_1285,In_1703);
nor U2957 (N_2957,In_1470,In_1571);
or U2958 (N_2958,In_1192,In_1382);
or U2959 (N_2959,In_1159,In_1336);
or U2960 (N_2960,In_1304,In_26);
xnor U2961 (N_2961,In_1182,In_1947);
or U2962 (N_2962,In_707,In_548);
or U2963 (N_2963,In_191,In_103);
xor U2964 (N_2964,In_1665,In_1427);
nand U2965 (N_2965,In_510,In_402);
or U2966 (N_2966,In_813,In_1076);
and U2967 (N_2967,In_1981,In_1206);
nor U2968 (N_2968,In_1392,In_1379);
and U2969 (N_2969,In_1841,In_591);
and U2970 (N_2970,In_752,In_1030);
and U2971 (N_2971,In_997,In_686);
xor U2972 (N_2972,In_91,In_1148);
and U2973 (N_2973,In_461,In_689);
nand U2974 (N_2974,In_560,In_1413);
xnor U2975 (N_2975,In_411,In_354);
xor U2976 (N_2976,In_942,In_895);
nor U2977 (N_2977,In_1706,In_1485);
xor U2978 (N_2978,In_1463,In_880);
and U2979 (N_2979,In_72,In_146);
xor U2980 (N_2980,In_717,In_1351);
or U2981 (N_2981,In_1667,In_1207);
xor U2982 (N_2982,In_1956,In_739);
xnor U2983 (N_2983,In_895,In_698);
nand U2984 (N_2984,In_685,In_1362);
or U2985 (N_2985,In_1906,In_99);
nand U2986 (N_2986,In_586,In_1290);
nor U2987 (N_2987,In_1568,In_1280);
and U2988 (N_2988,In_414,In_1878);
nand U2989 (N_2989,In_176,In_1674);
or U2990 (N_2990,In_565,In_1153);
xnor U2991 (N_2991,In_1137,In_1836);
or U2992 (N_2992,In_1720,In_630);
nor U2993 (N_2993,In_1566,In_256);
or U2994 (N_2994,In_241,In_1316);
nor U2995 (N_2995,In_1622,In_1770);
xnor U2996 (N_2996,In_99,In_1264);
or U2997 (N_2997,In_855,In_949);
xnor U2998 (N_2998,In_470,In_1171);
nor U2999 (N_2999,In_306,In_1709);
xnor U3000 (N_3000,In_553,In_1494);
and U3001 (N_3001,In_1752,In_1002);
nand U3002 (N_3002,In_873,In_1945);
nand U3003 (N_3003,In_305,In_691);
nand U3004 (N_3004,In_1409,In_1865);
xor U3005 (N_3005,In_566,In_1307);
and U3006 (N_3006,In_1212,In_441);
and U3007 (N_3007,In_390,In_1413);
or U3008 (N_3008,In_335,In_1705);
nand U3009 (N_3009,In_1048,In_678);
nand U3010 (N_3010,In_545,In_1323);
or U3011 (N_3011,In_272,In_7);
xor U3012 (N_3012,In_1277,In_182);
nor U3013 (N_3013,In_141,In_1428);
or U3014 (N_3014,In_374,In_1079);
or U3015 (N_3015,In_924,In_442);
and U3016 (N_3016,In_261,In_1846);
nor U3017 (N_3017,In_854,In_1677);
or U3018 (N_3018,In_590,In_1127);
and U3019 (N_3019,In_752,In_1193);
and U3020 (N_3020,In_458,In_420);
and U3021 (N_3021,In_445,In_1527);
and U3022 (N_3022,In_350,In_1664);
or U3023 (N_3023,In_1257,In_1739);
nor U3024 (N_3024,In_174,In_439);
nor U3025 (N_3025,In_36,In_1616);
and U3026 (N_3026,In_827,In_801);
or U3027 (N_3027,In_387,In_1295);
nand U3028 (N_3028,In_1362,In_1742);
nor U3029 (N_3029,In_1114,In_595);
xor U3030 (N_3030,In_556,In_226);
and U3031 (N_3031,In_628,In_892);
xnor U3032 (N_3032,In_1841,In_1715);
or U3033 (N_3033,In_391,In_1960);
xnor U3034 (N_3034,In_1945,In_836);
or U3035 (N_3035,In_1254,In_515);
and U3036 (N_3036,In_40,In_121);
xor U3037 (N_3037,In_1455,In_1029);
and U3038 (N_3038,In_358,In_1953);
nor U3039 (N_3039,In_473,In_1432);
xor U3040 (N_3040,In_1855,In_277);
nand U3041 (N_3041,In_1920,In_1372);
xnor U3042 (N_3042,In_601,In_711);
or U3043 (N_3043,In_835,In_615);
xor U3044 (N_3044,In_178,In_1231);
and U3045 (N_3045,In_1362,In_212);
nand U3046 (N_3046,In_903,In_155);
xnor U3047 (N_3047,In_1254,In_128);
nand U3048 (N_3048,In_395,In_1425);
nor U3049 (N_3049,In_992,In_670);
or U3050 (N_3050,In_621,In_549);
nand U3051 (N_3051,In_881,In_874);
nor U3052 (N_3052,In_469,In_69);
nor U3053 (N_3053,In_1847,In_1810);
and U3054 (N_3054,In_1913,In_268);
and U3055 (N_3055,In_330,In_1635);
xnor U3056 (N_3056,In_1666,In_1560);
xor U3057 (N_3057,In_1519,In_385);
and U3058 (N_3058,In_1933,In_1847);
xnor U3059 (N_3059,In_587,In_1208);
nand U3060 (N_3060,In_1214,In_1076);
nand U3061 (N_3061,In_1551,In_749);
and U3062 (N_3062,In_19,In_1650);
or U3063 (N_3063,In_1877,In_904);
or U3064 (N_3064,In_1712,In_443);
or U3065 (N_3065,In_1846,In_1937);
nor U3066 (N_3066,In_1731,In_62);
and U3067 (N_3067,In_638,In_1837);
xnor U3068 (N_3068,In_1594,In_1997);
nor U3069 (N_3069,In_321,In_1107);
xor U3070 (N_3070,In_1811,In_608);
xnor U3071 (N_3071,In_85,In_651);
nor U3072 (N_3072,In_927,In_81);
or U3073 (N_3073,In_399,In_800);
nor U3074 (N_3074,In_1237,In_410);
xnor U3075 (N_3075,In_376,In_1099);
xor U3076 (N_3076,In_919,In_1656);
nand U3077 (N_3077,In_948,In_1194);
nor U3078 (N_3078,In_1516,In_1067);
and U3079 (N_3079,In_1690,In_744);
nor U3080 (N_3080,In_94,In_1081);
nor U3081 (N_3081,In_962,In_1030);
xor U3082 (N_3082,In_571,In_558);
or U3083 (N_3083,In_155,In_1306);
or U3084 (N_3084,In_426,In_14);
and U3085 (N_3085,In_1271,In_82);
nor U3086 (N_3086,In_1033,In_1948);
and U3087 (N_3087,In_462,In_1116);
and U3088 (N_3088,In_1942,In_673);
xor U3089 (N_3089,In_497,In_1094);
nand U3090 (N_3090,In_959,In_1255);
xor U3091 (N_3091,In_1461,In_988);
nor U3092 (N_3092,In_650,In_120);
nor U3093 (N_3093,In_172,In_7);
or U3094 (N_3094,In_417,In_609);
nand U3095 (N_3095,In_1601,In_930);
or U3096 (N_3096,In_1065,In_1241);
or U3097 (N_3097,In_134,In_1944);
nor U3098 (N_3098,In_981,In_1862);
nand U3099 (N_3099,In_1626,In_776);
nor U3100 (N_3100,In_1183,In_266);
nor U3101 (N_3101,In_1241,In_1389);
nand U3102 (N_3102,In_220,In_792);
nor U3103 (N_3103,In_1211,In_590);
and U3104 (N_3104,In_461,In_1353);
and U3105 (N_3105,In_750,In_1613);
and U3106 (N_3106,In_826,In_289);
and U3107 (N_3107,In_17,In_611);
or U3108 (N_3108,In_882,In_1075);
nand U3109 (N_3109,In_663,In_1778);
or U3110 (N_3110,In_526,In_1657);
xnor U3111 (N_3111,In_813,In_936);
or U3112 (N_3112,In_831,In_583);
xor U3113 (N_3113,In_1388,In_1327);
nand U3114 (N_3114,In_1174,In_409);
and U3115 (N_3115,In_283,In_567);
and U3116 (N_3116,In_850,In_129);
nor U3117 (N_3117,In_438,In_447);
and U3118 (N_3118,In_1696,In_1972);
and U3119 (N_3119,In_214,In_170);
nand U3120 (N_3120,In_798,In_679);
nor U3121 (N_3121,In_1470,In_1691);
xnor U3122 (N_3122,In_1539,In_1009);
nand U3123 (N_3123,In_159,In_1389);
or U3124 (N_3124,In_1109,In_554);
or U3125 (N_3125,In_1028,In_1476);
nand U3126 (N_3126,In_1246,In_1719);
nand U3127 (N_3127,In_1483,In_178);
or U3128 (N_3128,In_1004,In_1677);
xnor U3129 (N_3129,In_1232,In_1387);
xnor U3130 (N_3130,In_362,In_221);
nor U3131 (N_3131,In_214,In_1147);
xor U3132 (N_3132,In_1642,In_627);
xnor U3133 (N_3133,In_1335,In_89);
nor U3134 (N_3134,In_214,In_1048);
and U3135 (N_3135,In_124,In_422);
and U3136 (N_3136,In_1899,In_520);
or U3137 (N_3137,In_1416,In_1116);
nor U3138 (N_3138,In_491,In_1788);
or U3139 (N_3139,In_456,In_1413);
nand U3140 (N_3140,In_1885,In_644);
nand U3141 (N_3141,In_1362,In_1714);
xnor U3142 (N_3142,In_956,In_1090);
xnor U3143 (N_3143,In_1014,In_65);
nand U3144 (N_3144,In_954,In_912);
and U3145 (N_3145,In_57,In_257);
nand U3146 (N_3146,In_1867,In_1219);
or U3147 (N_3147,In_383,In_787);
or U3148 (N_3148,In_660,In_285);
nand U3149 (N_3149,In_437,In_812);
xor U3150 (N_3150,In_273,In_1502);
nand U3151 (N_3151,In_1810,In_1364);
nand U3152 (N_3152,In_1835,In_654);
xnor U3153 (N_3153,In_1139,In_252);
and U3154 (N_3154,In_1174,In_1205);
and U3155 (N_3155,In_262,In_1276);
nand U3156 (N_3156,In_807,In_1988);
xor U3157 (N_3157,In_1540,In_1622);
nand U3158 (N_3158,In_644,In_1300);
xnor U3159 (N_3159,In_344,In_114);
nand U3160 (N_3160,In_1515,In_485);
xor U3161 (N_3161,In_1783,In_1254);
nor U3162 (N_3162,In_869,In_1879);
xnor U3163 (N_3163,In_1199,In_366);
xor U3164 (N_3164,In_1869,In_456);
or U3165 (N_3165,In_677,In_1952);
xnor U3166 (N_3166,In_143,In_338);
and U3167 (N_3167,In_432,In_1345);
nand U3168 (N_3168,In_493,In_791);
nor U3169 (N_3169,In_660,In_246);
nor U3170 (N_3170,In_813,In_448);
or U3171 (N_3171,In_885,In_689);
nor U3172 (N_3172,In_1846,In_1220);
nand U3173 (N_3173,In_427,In_104);
nor U3174 (N_3174,In_557,In_291);
or U3175 (N_3175,In_267,In_1755);
nand U3176 (N_3176,In_397,In_1809);
nand U3177 (N_3177,In_1916,In_1597);
or U3178 (N_3178,In_1349,In_715);
and U3179 (N_3179,In_141,In_1445);
nor U3180 (N_3180,In_1365,In_300);
xnor U3181 (N_3181,In_1137,In_1049);
nand U3182 (N_3182,In_430,In_1409);
xnor U3183 (N_3183,In_765,In_1260);
xnor U3184 (N_3184,In_1791,In_974);
and U3185 (N_3185,In_559,In_1532);
and U3186 (N_3186,In_1647,In_1964);
nor U3187 (N_3187,In_1208,In_333);
xnor U3188 (N_3188,In_1899,In_1038);
nor U3189 (N_3189,In_356,In_1681);
nor U3190 (N_3190,In_1735,In_1693);
and U3191 (N_3191,In_608,In_1547);
nand U3192 (N_3192,In_1655,In_119);
and U3193 (N_3193,In_599,In_669);
and U3194 (N_3194,In_191,In_458);
xnor U3195 (N_3195,In_979,In_1138);
xnor U3196 (N_3196,In_267,In_431);
and U3197 (N_3197,In_674,In_1588);
and U3198 (N_3198,In_251,In_947);
and U3199 (N_3199,In_407,In_1272);
nand U3200 (N_3200,In_404,In_1905);
xor U3201 (N_3201,In_1089,In_491);
nand U3202 (N_3202,In_902,In_674);
nor U3203 (N_3203,In_1165,In_785);
nor U3204 (N_3204,In_1290,In_986);
nor U3205 (N_3205,In_1275,In_1523);
nor U3206 (N_3206,In_1853,In_1925);
nor U3207 (N_3207,In_1094,In_1287);
nor U3208 (N_3208,In_449,In_113);
nor U3209 (N_3209,In_1736,In_1215);
xnor U3210 (N_3210,In_1938,In_1812);
or U3211 (N_3211,In_400,In_1580);
nand U3212 (N_3212,In_1067,In_1540);
xnor U3213 (N_3213,In_580,In_1298);
or U3214 (N_3214,In_172,In_307);
or U3215 (N_3215,In_1900,In_65);
nor U3216 (N_3216,In_1725,In_445);
xor U3217 (N_3217,In_1813,In_1189);
nor U3218 (N_3218,In_82,In_1852);
nand U3219 (N_3219,In_1395,In_1434);
or U3220 (N_3220,In_44,In_1582);
nor U3221 (N_3221,In_132,In_1011);
xor U3222 (N_3222,In_119,In_1493);
nand U3223 (N_3223,In_273,In_1779);
nor U3224 (N_3224,In_516,In_129);
and U3225 (N_3225,In_1965,In_460);
and U3226 (N_3226,In_861,In_995);
or U3227 (N_3227,In_465,In_681);
nor U3228 (N_3228,In_1202,In_1252);
nor U3229 (N_3229,In_1740,In_101);
nand U3230 (N_3230,In_948,In_173);
nor U3231 (N_3231,In_1005,In_1771);
and U3232 (N_3232,In_1374,In_605);
and U3233 (N_3233,In_453,In_358);
xor U3234 (N_3234,In_974,In_352);
xnor U3235 (N_3235,In_1625,In_62);
or U3236 (N_3236,In_1746,In_1445);
nor U3237 (N_3237,In_440,In_336);
nor U3238 (N_3238,In_286,In_704);
xor U3239 (N_3239,In_843,In_616);
xor U3240 (N_3240,In_1754,In_1286);
nor U3241 (N_3241,In_828,In_1553);
nand U3242 (N_3242,In_1332,In_579);
nand U3243 (N_3243,In_1720,In_492);
or U3244 (N_3244,In_817,In_418);
and U3245 (N_3245,In_1006,In_1591);
nand U3246 (N_3246,In_1190,In_206);
nand U3247 (N_3247,In_1181,In_1313);
and U3248 (N_3248,In_1924,In_1926);
nor U3249 (N_3249,In_861,In_1267);
nor U3250 (N_3250,In_1294,In_227);
or U3251 (N_3251,In_1130,In_1665);
or U3252 (N_3252,In_936,In_462);
nand U3253 (N_3253,In_881,In_444);
or U3254 (N_3254,In_776,In_281);
or U3255 (N_3255,In_1970,In_888);
nor U3256 (N_3256,In_66,In_255);
and U3257 (N_3257,In_1024,In_325);
xor U3258 (N_3258,In_1258,In_342);
nand U3259 (N_3259,In_444,In_1340);
nor U3260 (N_3260,In_1386,In_38);
and U3261 (N_3261,In_481,In_1626);
or U3262 (N_3262,In_1222,In_589);
and U3263 (N_3263,In_1381,In_48);
or U3264 (N_3264,In_1275,In_1199);
or U3265 (N_3265,In_672,In_1856);
and U3266 (N_3266,In_806,In_1296);
or U3267 (N_3267,In_1247,In_446);
nand U3268 (N_3268,In_688,In_346);
xor U3269 (N_3269,In_1368,In_68);
or U3270 (N_3270,In_439,In_1457);
or U3271 (N_3271,In_214,In_1987);
nand U3272 (N_3272,In_1013,In_924);
nor U3273 (N_3273,In_1112,In_1486);
or U3274 (N_3274,In_513,In_413);
xnor U3275 (N_3275,In_1687,In_1090);
or U3276 (N_3276,In_1362,In_1095);
and U3277 (N_3277,In_635,In_1925);
nor U3278 (N_3278,In_1390,In_1194);
or U3279 (N_3279,In_1138,In_1048);
nor U3280 (N_3280,In_619,In_1528);
nand U3281 (N_3281,In_229,In_987);
and U3282 (N_3282,In_1411,In_17);
xnor U3283 (N_3283,In_1372,In_1773);
xor U3284 (N_3284,In_1974,In_579);
or U3285 (N_3285,In_1036,In_1687);
nand U3286 (N_3286,In_1119,In_1580);
or U3287 (N_3287,In_1352,In_736);
and U3288 (N_3288,In_1767,In_755);
nor U3289 (N_3289,In_69,In_1902);
xor U3290 (N_3290,In_1058,In_1250);
nand U3291 (N_3291,In_1687,In_188);
and U3292 (N_3292,In_304,In_1448);
nand U3293 (N_3293,In_279,In_740);
nand U3294 (N_3294,In_555,In_1508);
xor U3295 (N_3295,In_677,In_1143);
or U3296 (N_3296,In_1413,In_458);
or U3297 (N_3297,In_269,In_669);
or U3298 (N_3298,In_143,In_1943);
or U3299 (N_3299,In_143,In_810);
and U3300 (N_3300,In_1938,In_1398);
nor U3301 (N_3301,In_1556,In_637);
nor U3302 (N_3302,In_1582,In_815);
and U3303 (N_3303,In_605,In_1488);
nor U3304 (N_3304,In_1628,In_21);
and U3305 (N_3305,In_523,In_1648);
and U3306 (N_3306,In_569,In_233);
nor U3307 (N_3307,In_713,In_226);
nor U3308 (N_3308,In_1641,In_1777);
xor U3309 (N_3309,In_192,In_1391);
and U3310 (N_3310,In_165,In_486);
or U3311 (N_3311,In_678,In_191);
xnor U3312 (N_3312,In_623,In_546);
nand U3313 (N_3313,In_161,In_422);
or U3314 (N_3314,In_255,In_553);
nand U3315 (N_3315,In_110,In_226);
xnor U3316 (N_3316,In_327,In_1685);
or U3317 (N_3317,In_1597,In_1659);
nand U3318 (N_3318,In_1773,In_318);
nand U3319 (N_3319,In_780,In_1029);
and U3320 (N_3320,In_1457,In_73);
nand U3321 (N_3321,In_990,In_423);
xor U3322 (N_3322,In_793,In_1912);
and U3323 (N_3323,In_1621,In_815);
and U3324 (N_3324,In_1549,In_884);
and U3325 (N_3325,In_310,In_991);
nand U3326 (N_3326,In_1214,In_213);
nor U3327 (N_3327,In_1304,In_252);
and U3328 (N_3328,In_1101,In_472);
and U3329 (N_3329,In_1387,In_254);
and U3330 (N_3330,In_1824,In_1939);
or U3331 (N_3331,In_309,In_570);
xnor U3332 (N_3332,In_181,In_388);
and U3333 (N_3333,In_675,In_1946);
xor U3334 (N_3334,In_660,In_1565);
nor U3335 (N_3335,In_61,In_1944);
or U3336 (N_3336,In_266,In_255);
or U3337 (N_3337,In_1567,In_1209);
nand U3338 (N_3338,In_1499,In_1135);
and U3339 (N_3339,In_1398,In_1027);
nor U3340 (N_3340,In_1821,In_197);
nor U3341 (N_3341,In_658,In_706);
nor U3342 (N_3342,In_1480,In_1842);
xnor U3343 (N_3343,In_1574,In_1414);
nor U3344 (N_3344,In_1054,In_1326);
nand U3345 (N_3345,In_1342,In_368);
and U3346 (N_3346,In_304,In_1050);
or U3347 (N_3347,In_297,In_592);
nand U3348 (N_3348,In_1588,In_1775);
and U3349 (N_3349,In_1824,In_102);
nor U3350 (N_3350,In_1427,In_494);
nor U3351 (N_3351,In_367,In_941);
nor U3352 (N_3352,In_1005,In_446);
xor U3353 (N_3353,In_637,In_327);
or U3354 (N_3354,In_1585,In_720);
xor U3355 (N_3355,In_1688,In_1963);
or U3356 (N_3356,In_1837,In_1322);
and U3357 (N_3357,In_101,In_330);
nand U3358 (N_3358,In_677,In_710);
nor U3359 (N_3359,In_123,In_1231);
and U3360 (N_3360,In_1650,In_593);
nor U3361 (N_3361,In_1896,In_622);
nor U3362 (N_3362,In_944,In_932);
nor U3363 (N_3363,In_467,In_173);
xnor U3364 (N_3364,In_1033,In_1113);
nand U3365 (N_3365,In_1787,In_588);
or U3366 (N_3366,In_1949,In_1841);
or U3367 (N_3367,In_951,In_25);
nor U3368 (N_3368,In_1717,In_58);
nand U3369 (N_3369,In_1709,In_677);
xor U3370 (N_3370,In_1675,In_1374);
nand U3371 (N_3371,In_843,In_1641);
nand U3372 (N_3372,In_1395,In_812);
and U3373 (N_3373,In_403,In_637);
and U3374 (N_3374,In_1968,In_267);
and U3375 (N_3375,In_1077,In_1541);
or U3376 (N_3376,In_921,In_1687);
or U3377 (N_3377,In_216,In_1991);
nand U3378 (N_3378,In_822,In_1727);
nor U3379 (N_3379,In_726,In_8);
or U3380 (N_3380,In_342,In_1320);
xor U3381 (N_3381,In_1706,In_686);
nor U3382 (N_3382,In_1044,In_1210);
xnor U3383 (N_3383,In_816,In_991);
or U3384 (N_3384,In_821,In_29);
and U3385 (N_3385,In_167,In_209);
xnor U3386 (N_3386,In_1460,In_940);
xor U3387 (N_3387,In_658,In_1312);
nand U3388 (N_3388,In_1618,In_1879);
nand U3389 (N_3389,In_803,In_884);
xnor U3390 (N_3390,In_1755,In_192);
nor U3391 (N_3391,In_358,In_637);
and U3392 (N_3392,In_898,In_1977);
xnor U3393 (N_3393,In_1730,In_1114);
xor U3394 (N_3394,In_414,In_1281);
nand U3395 (N_3395,In_1000,In_1537);
nor U3396 (N_3396,In_1715,In_347);
and U3397 (N_3397,In_105,In_1538);
nand U3398 (N_3398,In_727,In_1673);
and U3399 (N_3399,In_536,In_49);
and U3400 (N_3400,In_481,In_479);
or U3401 (N_3401,In_759,In_247);
or U3402 (N_3402,In_1663,In_1984);
nand U3403 (N_3403,In_712,In_1921);
or U3404 (N_3404,In_1615,In_1399);
xor U3405 (N_3405,In_235,In_871);
or U3406 (N_3406,In_1203,In_916);
xnor U3407 (N_3407,In_1727,In_1802);
xor U3408 (N_3408,In_861,In_160);
nor U3409 (N_3409,In_1700,In_1131);
and U3410 (N_3410,In_1188,In_1160);
xnor U3411 (N_3411,In_911,In_760);
or U3412 (N_3412,In_389,In_1280);
nand U3413 (N_3413,In_375,In_351);
and U3414 (N_3414,In_356,In_92);
xnor U3415 (N_3415,In_1851,In_462);
xor U3416 (N_3416,In_812,In_1267);
and U3417 (N_3417,In_74,In_329);
xnor U3418 (N_3418,In_225,In_1997);
xnor U3419 (N_3419,In_796,In_579);
nor U3420 (N_3420,In_1699,In_562);
and U3421 (N_3421,In_208,In_1735);
nor U3422 (N_3422,In_233,In_224);
nor U3423 (N_3423,In_1753,In_443);
and U3424 (N_3424,In_1041,In_1283);
nand U3425 (N_3425,In_331,In_1556);
nand U3426 (N_3426,In_800,In_1444);
or U3427 (N_3427,In_1177,In_1621);
and U3428 (N_3428,In_758,In_1599);
xnor U3429 (N_3429,In_1593,In_1227);
nor U3430 (N_3430,In_750,In_1001);
nor U3431 (N_3431,In_1475,In_1713);
and U3432 (N_3432,In_367,In_1265);
nand U3433 (N_3433,In_569,In_676);
nand U3434 (N_3434,In_521,In_779);
nand U3435 (N_3435,In_1076,In_1849);
xor U3436 (N_3436,In_1512,In_1970);
xor U3437 (N_3437,In_62,In_1698);
nand U3438 (N_3438,In_194,In_435);
or U3439 (N_3439,In_1705,In_68);
nor U3440 (N_3440,In_1309,In_457);
or U3441 (N_3441,In_1438,In_929);
nor U3442 (N_3442,In_1254,In_1662);
or U3443 (N_3443,In_988,In_1554);
or U3444 (N_3444,In_1542,In_1855);
nand U3445 (N_3445,In_1604,In_544);
nand U3446 (N_3446,In_462,In_1842);
and U3447 (N_3447,In_895,In_1400);
nand U3448 (N_3448,In_1983,In_961);
nand U3449 (N_3449,In_1176,In_564);
and U3450 (N_3450,In_913,In_1596);
xor U3451 (N_3451,In_1512,In_1947);
nand U3452 (N_3452,In_1220,In_1380);
nand U3453 (N_3453,In_1813,In_1645);
and U3454 (N_3454,In_1198,In_1373);
nand U3455 (N_3455,In_596,In_1374);
or U3456 (N_3456,In_1574,In_1949);
or U3457 (N_3457,In_1000,In_806);
xnor U3458 (N_3458,In_628,In_1936);
nor U3459 (N_3459,In_792,In_1530);
xnor U3460 (N_3460,In_1411,In_862);
xnor U3461 (N_3461,In_1391,In_1493);
xor U3462 (N_3462,In_791,In_1139);
nor U3463 (N_3463,In_1451,In_1306);
xnor U3464 (N_3464,In_597,In_1810);
or U3465 (N_3465,In_1104,In_1147);
and U3466 (N_3466,In_421,In_658);
and U3467 (N_3467,In_963,In_1043);
xor U3468 (N_3468,In_1087,In_1040);
and U3469 (N_3469,In_671,In_727);
or U3470 (N_3470,In_1922,In_1781);
nand U3471 (N_3471,In_1023,In_1623);
and U3472 (N_3472,In_785,In_378);
nand U3473 (N_3473,In_215,In_838);
nor U3474 (N_3474,In_129,In_246);
nor U3475 (N_3475,In_1654,In_241);
nor U3476 (N_3476,In_1378,In_1993);
and U3477 (N_3477,In_1659,In_1774);
xnor U3478 (N_3478,In_412,In_925);
or U3479 (N_3479,In_739,In_1623);
xnor U3480 (N_3480,In_167,In_1746);
nand U3481 (N_3481,In_1383,In_946);
or U3482 (N_3482,In_44,In_1683);
or U3483 (N_3483,In_1457,In_155);
and U3484 (N_3484,In_1626,In_1878);
nand U3485 (N_3485,In_214,In_1435);
nor U3486 (N_3486,In_1,In_1236);
xor U3487 (N_3487,In_987,In_1633);
and U3488 (N_3488,In_1692,In_701);
or U3489 (N_3489,In_1739,In_1379);
nand U3490 (N_3490,In_732,In_1992);
nand U3491 (N_3491,In_1483,In_330);
or U3492 (N_3492,In_661,In_256);
xor U3493 (N_3493,In_853,In_1177);
nor U3494 (N_3494,In_1174,In_1048);
or U3495 (N_3495,In_752,In_1756);
and U3496 (N_3496,In_667,In_631);
nor U3497 (N_3497,In_637,In_1565);
xor U3498 (N_3498,In_1739,In_1541);
nor U3499 (N_3499,In_1862,In_1590);
and U3500 (N_3500,In_1140,In_1853);
nand U3501 (N_3501,In_1655,In_448);
nand U3502 (N_3502,In_1576,In_129);
nand U3503 (N_3503,In_1841,In_110);
nor U3504 (N_3504,In_1702,In_672);
nand U3505 (N_3505,In_1430,In_139);
nor U3506 (N_3506,In_1010,In_1077);
and U3507 (N_3507,In_1010,In_483);
nor U3508 (N_3508,In_380,In_598);
and U3509 (N_3509,In_1525,In_1640);
nand U3510 (N_3510,In_1922,In_1929);
nand U3511 (N_3511,In_1886,In_1025);
and U3512 (N_3512,In_1076,In_35);
or U3513 (N_3513,In_1049,In_952);
nand U3514 (N_3514,In_1681,In_1848);
and U3515 (N_3515,In_933,In_1322);
xor U3516 (N_3516,In_1610,In_424);
or U3517 (N_3517,In_760,In_1972);
xor U3518 (N_3518,In_1174,In_1148);
nand U3519 (N_3519,In_1224,In_652);
nor U3520 (N_3520,In_1403,In_1577);
nor U3521 (N_3521,In_1063,In_904);
or U3522 (N_3522,In_1433,In_1869);
nor U3523 (N_3523,In_1035,In_1864);
nand U3524 (N_3524,In_821,In_652);
and U3525 (N_3525,In_1587,In_930);
or U3526 (N_3526,In_1551,In_1350);
xor U3527 (N_3527,In_1832,In_464);
xor U3528 (N_3528,In_819,In_1007);
and U3529 (N_3529,In_566,In_312);
nand U3530 (N_3530,In_1326,In_798);
or U3531 (N_3531,In_1757,In_429);
xor U3532 (N_3532,In_1563,In_1336);
and U3533 (N_3533,In_229,In_344);
nand U3534 (N_3534,In_550,In_1072);
xnor U3535 (N_3535,In_441,In_634);
xor U3536 (N_3536,In_1501,In_1284);
and U3537 (N_3537,In_912,In_1883);
or U3538 (N_3538,In_37,In_1899);
xor U3539 (N_3539,In_1800,In_1915);
nand U3540 (N_3540,In_1242,In_671);
nor U3541 (N_3541,In_1663,In_1307);
or U3542 (N_3542,In_569,In_935);
and U3543 (N_3543,In_1856,In_1081);
or U3544 (N_3544,In_913,In_1516);
nor U3545 (N_3545,In_1720,In_384);
nand U3546 (N_3546,In_1497,In_331);
or U3547 (N_3547,In_501,In_404);
nand U3548 (N_3548,In_1516,In_1686);
or U3549 (N_3549,In_4,In_808);
nand U3550 (N_3550,In_620,In_1795);
nand U3551 (N_3551,In_897,In_1237);
or U3552 (N_3552,In_458,In_1627);
nor U3553 (N_3553,In_1915,In_850);
xnor U3554 (N_3554,In_1131,In_648);
nor U3555 (N_3555,In_248,In_1863);
nor U3556 (N_3556,In_152,In_300);
nor U3557 (N_3557,In_920,In_543);
nor U3558 (N_3558,In_1135,In_596);
nor U3559 (N_3559,In_393,In_384);
xnor U3560 (N_3560,In_1015,In_182);
nor U3561 (N_3561,In_1618,In_1440);
nand U3562 (N_3562,In_714,In_1787);
nand U3563 (N_3563,In_178,In_16);
nand U3564 (N_3564,In_484,In_607);
or U3565 (N_3565,In_477,In_697);
or U3566 (N_3566,In_807,In_1044);
nand U3567 (N_3567,In_1806,In_878);
and U3568 (N_3568,In_191,In_330);
nand U3569 (N_3569,In_981,In_278);
xor U3570 (N_3570,In_282,In_1521);
xnor U3571 (N_3571,In_1077,In_590);
or U3572 (N_3572,In_993,In_1217);
xor U3573 (N_3573,In_94,In_680);
and U3574 (N_3574,In_1037,In_225);
and U3575 (N_3575,In_972,In_1474);
nand U3576 (N_3576,In_428,In_921);
nand U3577 (N_3577,In_443,In_484);
nand U3578 (N_3578,In_783,In_1904);
or U3579 (N_3579,In_1010,In_751);
nor U3580 (N_3580,In_1139,In_1390);
nor U3581 (N_3581,In_1813,In_1952);
or U3582 (N_3582,In_1814,In_269);
and U3583 (N_3583,In_1068,In_1467);
nor U3584 (N_3584,In_1538,In_1992);
nor U3585 (N_3585,In_689,In_1559);
nor U3586 (N_3586,In_1657,In_324);
nand U3587 (N_3587,In_1747,In_1607);
nor U3588 (N_3588,In_1289,In_760);
and U3589 (N_3589,In_1514,In_1467);
and U3590 (N_3590,In_1312,In_1448);
nor U3591 (N_3591,In_802,In_1124);
nor U3592 (N_3592,In_1077,In_101);
nand U3593 (N_3593,In_1612,In_1495);
xnor U3594 (N_3594,In_1098,In_1705);
and U3595 (N_3595,In_291,In_602);
and U3596 (N_3596,In_878,In_1789);
xnor U3597 (N_3597,In_344,In_1972);
nor U3598 (N_3598,In_1458,In_1352);
xnor U3599 (N_3599,In_1471,In_1890);
nor U3600 (N_3600,In_955,In_1483);
xor U3601 (N_3601,In_1059,In_1241);
or U3602 (N_3602,In_84,In_16);
and U3603 (N_3603,In_1073,In_1257);
nor U3604 (N_3604,In_432,In_1789);
or U3605 (N_3605,In_1270,In_1701);
nor U3606 (N_3606,In_1680,In_381);
nand U3607 (N_3607,In_1714,In_990);
nand U3608 (N_3608,In_975,In_64);
nand U3609 (N_3609,In_243,In_1319);
or U3610 (N_3610,In_1511,In_1572);
or U3611 (N_3611,In_1478,In_1013);
nor U3612 (N_3612,In_34,In_855);
or U3613 (N_3613,In_1876,In_1097);
nor U3614 (N_3614,In_648,In_545);
xnor U3615 (N_3615,In_1655,In_1454);
nand U3616 (N_3616,In_1315,In_1189);
nand U3617 (N_3617,In_130,In_154);
and U3618 (N_3618,In_1556,In_592);
nand U3619 (N_3619,In_1406,In_1679);
nor U3620 (N_3620,In_45,In_1361);
or U3621 (N_3621,In_876,In_69);
nand U3622 (N_3622,In_1219,In_540);
nor U3623 (N_3623,In_1472,In_52);
and U3624 (N_3624,In_736,In_1694);
nor U3625 (N_3625,In_438,In_1189);
xnor U3626 (N_3626,In_1421,In_515);
nand U3627 (N_3627,In_503,In_1419);
or U3628 (N_3628,In_1325,In_1566);
and U3629 (N_3629,In_787,In_1163);
nor U3630 (N_3630,In_527,In_207);
xnor U3631 (N_3631,In_250,In_797);
and U3632 (N_3632,In_580,In_768);
and U3633 (N_3633,In_237,In_1608);
nor U3634 (N_3634,In_1936,In_1610);
nor U3635 (N_3635,In_1551,In_864);
or U3636 (N_3636,In_1301,In_1587);
nor U3637 (N_3637,In_32,In_1037);
or U3638 (N_3638,In_1745,In_1680);
nor U3639 (N_3639,In_1314,In_276);
and U3640 (N_3640,In_1738,In_1276);
and U3641 (N_3641,In_982,In_399);
nand U3642 (N_3642,In_898,In_690);
nor U3643 (N_3643,In_1303,In_460);
and U3644 (N_3644,In_444,In_138);
and U3645 (N_3645,In_562,In_1681);
nor U3646 (N_3646,In_1635,In_654);
nand U3647 (N_3647,In_1001,In_939);
nand U3648 (N_3648,In_1631,In_1319);
xnor U3649 (N_3649,In_634,In_1537);
xnor U3650 (N_3650,In_617,In_782);
and U3651 (N_3651,In_1710,In_619);
nor U3652 (N_3652,In_1702,In_893);
xor U3653 (N_3653,In_388,In_1068);
xnor U3654 (N_3654,In_8,In_398);
or U3655 (N_3655,In_1595,In_1525);
nand U3656 (N_3656,In_192,In_1465);
or U3657 (N_3657,In_1397,In_1713);
xor U3658 (N_3658,In_741,In_1297);
xor U3659 (N_3659,In_1655,In_133);
or U3660 (N_3660,In_1604,In_402);
nor U3661 (N_3661,In_1940,In_1623);
and U3662 (N_3662,In_769,In_1922);
nand U3663 (N_3663,In_1495,In_1868);
xor U3664 (N_3664,In_98,In_1363);
xnor U3665 (N_3665,In_1449,In_1839);
and U3666 (N_3666,In_1075,In_1540);
nor U3667 (N_3667,In_1868,In_1786);
nor U3668 (N_3668,In_199,In_1260);
xor U3669 (N_3669,In_1034,In_728);
nor U3670 (N_3670,In_1312,In_417);
nand U3671 (N_3671,In_1057,In_583);
xor U3672 (N_3672,In_711,In_1524);
and U3673 (N_3673,In_1560,In_1921);
nand U3674 (N_3674,In_164,In_320);
or U3675 (N_3675,In_1803,In_1914);
and U3676 (N_3676,In_1339,In_1855);
xnor U3677 (N_3677,In_285,In_512);
nor U3678 (N_3678,In_1949,In_1620);
or U3679 (N_3679,In_1758,In_691);
nand U3680 (N_3680,In_1214,In_1516);
xor U3681 (N_3681,In_1165,In_891);
and U3682 (N_3682,In_934,In_573);
nor U3683 (N_3683,In_1708,In_601);
or U3684 (N_3684,In_1118,In_283);
nor U3685 (N_3685,In_1253,In_476);
and U3686 (N_3686,In_1093,In_446);
and U3687 (N_3687,In_706,In_176);
nand U3688 (N_3688,In_1194,In_1324);
nor U3689 (N_3689,In_607,In_1110);
or U3690 (N_3690,In_1531,In_123);
and U3691 (N_3691,In_597,In_70);
nand U3692 (N_3692,In_880,In_1949);
and U3693 (N_3693,In_724,In_1430);
or U3694 (N_3694,In_1597,In_1);
nand U3695 (N_3695,In_1527,In_489);
nand U3696 (N_3696,In_1815,In_52);
or U3697 (N_3697,In_677,In_642);
or U3698 (N_3698,In_613,In_1601);
xor U3699 (N_3699,In_1113,In_1449);
xnor U3700 (N_3700,In_394,In_336);
nor U3701 (N_3701,In_778,In_1297);
and U3702 (N_3702,In_1703,In_1618);
xnor U3703 (N_3703,In_110,In_1662);
nand U3704 (N_3704,In_1290,In_78);
or U3705 (N_3705,In_1171,In_1474);
or U3706 (N_3706,In_1719,In_1546);
nand U3707 (N_3707,In_1767,In_131);
xor U3708 (N_3708,In_996,In_305);
nor U3709 (N_3709,In_774,In_1180);
xor U3710 (N_3710,In_1695,In_1166);
or U3711 (N_3711,In_1568,In_1309);
nor U3712 (N_3712,In_60,In_1380);
and U3713 (N_3713,In_1429,In_682);
and U3714 (N_3714,In_1718,In_1812);
and U3715 (N_3715,In_1662,In_1108);
xnor U3716 (N_3716,In_838,In_962);
xor U3717 (N_3717,In_492,In_1609);
and U3718 (N_3718,In_1158,In_430);
nor U3719 (N_3719,In_1635,In_1751);
xnor U3720 (N_3720,In_1856,In_779);
or U3721 (N_3721,In_305,In_143);
and U3722 (N_3722,In_1162,In_469);
or U3723 (N_3723,In_398,In_835);
nand U3724 (N_3724,In_1533,In_143);
and U3725 (N_3725,In_124,In_296);
or U3726 (N_3726,In_1294,In_1913);
xnor U3727 (N_3727,In_778,In_1000);
nand U3728 (N_3728,In_499,In_648);
nand U3729 (N_3729,In_1792,In_3);
nor U3730 (N_3730,In_1330,In_494);
xor U3731 (N_3731,In_233,In_1846);
or U3732 (N_3732,In_1630,In_1743);
or U3733 (N_3733,In_1461,In_747);
nor U3734 (N_3734,In_1976,In_538);
or U3735 (N_3735,In_1274,In_1938);
xor U3736 (N_3736,In_1737,In_1140);
and U3737 (N_3737,In_1522,In_795);
nor U3738 (N_3738,In_1724,In_1807);
nor U3739 (N_3739,In_473,In_1189);
nor U3740 (N_3740,In_1468,In_1298);
or U3741 (N_3741,In_125,In_1723);
or U3742 (N_3742,In_897,In_1395);
nor U3743 (N_3743,In_450,In_1996);
nor U3744 (N_3744,In_822,In_1746);
and U3745 (N_3745,In_273,In_1001);
nor U3746 (N_3746,In_367,In_354);
nand U3747 (N_3747,In_1464,In_1780);
xor U3748 (N_3748,In_395,In_1166);
nor U3749 (N_3749,In_670,In_912);
xor U3750 (N_3750,In_54,In_472);
xnor U3751 (N_3751,In_898,In_184);
nor U3752 (N_3752,In_1457,In_1985);
xor U3753 (N_3753,In_1565,In_529);
nand U3754 (N_3754,In_274,In_105);
and U3755 (N_3755,In_738,In_484);
and U3756 (N_3756,In_369,In_1879);
nand U3757 (N_3757,In_637,In_1866);
nand U3758 (N_3758,In_1960,In_1940);
xnor U3759 (N_3759,In_513,In_153);
nand U3760 (N_3760,In_414,In_509);
nor U3761 (N_3761,In_952,In_798);
or U3762 (N_3762,In_1504,In_1599);
nand U3763 (N_3763,In_251,In_1650);
nor U3764 (N_3764,In_616,In_1927);
and U3765 (N_3765,In_1785,In_1881);
xnor U3766 (N_3766,In_1543,In_1246);
or U3767 (N_3767,In_1264,In_230);
xnor U3768 (N_3768,In_1773,In_681);
nand U3769 (N_3769,In_322,In_621);
and U3770 (N_3770,In_1579,In_1758);
xnor U3771 (N_3771,In_230,In_356);
and U3772 (N_3772,In_11,In_83);
or U3773 (N_3773,In_478,In_700);
nor U3774 (N_3774,In_1349,In_1430);
nand U3775 (N_3775,In_1383,In_134);
and U3776 (N_3776,In_635,In_414);
or U3777 (N_3777,In_1076,In_494);
or U3778 (N_3778,In_1856,In_831);
and U3779 (N_3779,In_595,In_1308);
nand U3780 (N_3780,In_1988,In_776);
nor U3781 (N_3781,In_588,In_1457);
or U3782 (N_3782,In_1019,In_161);
and U3783 (N_3783,In_87,In_1000);
nor U3784 (N_3784,In_713,In_349);
xor U3785 (N_3785,In_1638,In_259);
nand U3786 (N_3786,In_1177,In_1160);
and U3787 (N_3787,In_150,In_133);
or U3788 (N_3788,In_1743,In_1573);
or U3789 (N_3789,In_1826,In_1331);
nor U3790 (N_3790,In_1799,In_201);
and U3791 (N_3791,In_997,In_203);
nor U3792 (N_3792,In_1381,In_1944);
and U3793 (N_3793,In_1981,In_761);
nor U3794 (N_3794,In_766,In_1244);
nor U3795 (N_3795,In_1187,In_151);
or U3796 (N_3796,In_540,In_1569);
or U3797 (N_3797,In_241,In_61);
or U3798 (N_3798,In_1473,In_1291);
or U3799 (N_3799,In_227,In_575);
nand U3800 (N_3800,In_1536,In_695);
or U3801 (N_3801,In_82,In_850);
or U3802 (N_3802,In_175,In_600);
xnor U3803 (N_3803,In_1106,In_1311);
nor U3804 (N_3804,In_1308,In_346);
and U3805 (N_3805,In_41,In_1170);
nor U3806 (N_3806,In_1994,In_624);
nand U3807 (N_3807,In_356,In_795);
xor U3808 (N_3808,In_118,In_1589);
and U3809 (N_3809,In_446,In_896);
nor U3810 (N_3810,In_1596,In_431);
xnor U3811 (N_3811,In_1681,In_158);
and U3812 (N_3812,In_904,In_571);
xor U3813 (N_3813,In_832,In_1339);
and U3814 (N_3814,In_924,In_802);
xor U3815 (N_3815,In_541,In_1778);
and U3816 (N_3816,In_645,In_1070);
nand U3817 (N_3817,In_1531,In_1039);
nor U3818 (N_3818,In_589,In_663);
xor U3819 (N_3819,In_1959,In_564);
and U3820 (N_3820,In_590,In_106);
nand U3821 (N_3821,In_1149,In_1601);
or U3822 (N_3822,In_1270,In_651);
nand U3823 (N_3823,In_1837,In_1153);
xnor U3824 (N_3824,In_422,In_1685);
or U3825 (N_3825,In_441,In_826);
and U3826 (N_3826,In_390,In_375);
nand U3827 (N_3827,In_1714,In_535);
xor U3828 (N_3828,In_786,In_1254);
and U3829 (N_3829,In_470,In_877);
xor U3830 (N_3830,In_786,In_1640);
nor U3831 (N_3831,In_1802,In_1134);
nand U3832 (N_3832,In_64,In_891);
xnor U3833 (N_3833,In_1021,In_993);
nand U3834 (N_3834,In_1500,In_175);
nor U3835 (N_3835,In_70,In_1040);
or U3836 (N_3836,In_1127,In_508);
xnor U3837 (N_3837,In_641,In_743);
nand U3838 (N_3838,In_1727,In_183);
nand U3839 (N_3839,In_832,In_1445);
and U3840 (N_3840,In_907,In_579);
or U3841 (N_3841,In_267,In_1043);
or U3842 (N_3842,In_709,In_1165);
nor U3843 (N_3843,In_1856,In_904);
xnor U3844 (N_3844,In_365,In_1211);
xor U3845 (N_3845,In_1648,In_1517);
xnor U3846 (N_3846,In_569,In_992);
nor U3847 (N_3847,In_818,In_313);
and U3848 (N_3848,In_121,In_638);
and U3849 (N_3849,In_496,In_1113);
nand U3850 (N_3850,In_1665,In_831);
nor U3851 (N_3851,In_935,In_1722);
nor U3852 (N_3852,In_727,In_703);
xnor U3853 (N_3853,In_978,In_734);
and U3854 (N_3854,In_21,In_1659);
nand U3855 (N_3855,In_192,In_861);
xor U3856 (N_3856,In_956,In_968);
and U3857 (N_3857,In_770,In_606);
or U3858 (N_3858,In_294,In_1958);
nor U3859 (N_3859,In_84,In_916);
nor U3860 (N_3860,In_1945,In_862);
and U3861 (N_3861,In_1940,In_87);
nand U3862 (N_3862,In_267,In_9);
or U3863 (N_3863,In_1089,In_1922);
xor U3864 (N_3864,In_1920,In_1932);
and U3865 (N_3865,In_1040,In_1093);
or U3866 (N_3866,In_585,In_1935);
xor U3867 (N_3867,In_1217,In_83);
nor U3868 (N_3868,In_525,In_613);
nand U3869 (N_3869,In_427,In_991);
xnor U3870 (N_3870,In_813,In_1914);
nand U3871 (N_3871,In_1780,In_1417);
and U3872 (N_3872,In_1715,In_1578);
or U3873 (N_3873,In_1979,In_364);
nor U3874 (N_3874,In_1344,In_195);
and U3875 (N_3875,In_1658,In_1495);
nand U3876 (N_3876,In_757,In_149);
xor U3877 (N_3877,In_463,In_434);
and U3878 (N_3878,In_1304,In_1009);
or U3879 (N_3879,In_1154,In_1987);
and U3880 (N_3880,In_1741,In_1535);
nor U3881 (N_3881,In_1973,In_1461);
nand U3882 (N_3882,In_730,In_1900);
nor U3883 (N_3883,In_500,In_226);
xor U3884 (N_3884,In_263,In_1803);
or U3885 (N_3885,In_1502,In_563);
xnor U3886 (N_3886,In_594,In_233);
and U3887 (N_3887,In_1765,In_721);
or U3888 (N_3888,In_200,In_549);
nand U3889 (N_3889,In_1762,In_1618);
xnor U3890 (N_3890,In_573,In_276);
nand U3891 (N_3891,In_1260,In_928);
nor U3892 (N_3892,In_1190,In_819);
nor U3893 (N_3893,In_1929,In_575);
nor U3894 (N_3894,In_184,In_662);
and U3895 (N_3895,In_57,In_1504);
nor U3896 (N_3896,In_425,In_586);
nand U3897 (N_3897,In_1954,In_1868);
xor U3898 (N_3898,In_1575,In_1720);
and U3899 (N_3899,In_408,In_544);
nand U3900 (N_3900,In_1806,In_1588);
or U3901 (N_3901,In_1654,In_1205);
xnor U3902 (N_3902,In_129,In_1919);
and U3903 (N_3903,In_488,In_1526);
nand U3904 (N_3904,In_902,In_1836);
and U3905 (N_3905,In_777,In_743);
xnor U3906 (N_3906,In_1245,In_1558);
and U3907 (N_3907,In_921,In_1145);
and U3908 (N_3908,In_499,In_425);
nand U3909 (N_3909,In_1668,In_1509);
nand U3910 (N_3910,In_1481,In_1463);
xnor U3911 (N_3911,In_1402,In_834);
and U3912 (N_3912,In_884,In_700);
nand U3913 (N_3913,In_571,In_1992);
xnor U3914 (N_3914,In_239,In_491);
xnor U3915 (N_3915,In_643,In_1515);
and U3916 (N_3916,In_1588,In_1402);
and U3917 (N_3917,In_735,In_454);
xor U3918 (N_3918,In_1371,In_1360);
xnor U3919 (N_3919,In_1272,In_269);
nor U3920 (N_3920,In_1663,In_1310);
nor U3921 (N_3921,In_1179,In_415);
xor U3922 (N_3922,In_1856,In_1888);
xnor U3923 (N_3923,In_1203,In_1439);
nand U3924 (N_3924,In_1010,In_1605);
nor U3925 (N_3925,In_174,In_831);
nor U3926 (N_3926,In_232,In_1090);
xor U3927 (N_3927,In_1963,In_1204);
xnor U3928 (N_3928,In_310,In_881);
nand U3929 (N_3929,In_387,In_1964);
and U3930 (N_3930,In_1010,In_1744);
or U3931 (N_3931,In_1829,In_1613);
and U3932 (N_3932,In_22,In_1587);
nand U3933 (N_3933,In_1955,In_1430);
xnor U3934 (N_3934,In_778,In_1733);
or U3935 (N_3935,In_661,In_1348);
or U3936 (N_3936,In_535,In_487);
and U3937 (N_3937,In_1518,In_335);
nor U3938 (N_3938,In_1070,In_1259);
or U3939 (N_3939,In_538,In_1099);
or U3940 (N_3940,In_446,In_724);
nor U3941 (N_3941,In_1041,In_1976);
nor U3942 (N_3942,In_1413,In_921);
xor U3943 (N_3943,In_619,In_1383);
xor U3944 (N_3944,In_1217,In_943);
xnor U3945 (N_3945,In_689,In_756);
and U3946 (N_3946,In_1778,In_709);
nand U3947 (N_3947,In_1914,In_913);
nand U3948 (N_3948,In_886,In_260);
and U3949 (N_3949,In_1971,In_1286);
and U3950 (N_3950,In_1553,In_948);
and U3951 (N_3951,In_825,In_768);
or U3952 (N_3952,In_460,In_1652);
or U3953 (N_3953,In_694,In_710);
or U3954 (N_3954,In_593,In_34);
nand U3955 (N_3955,In_971,In_841);
nand U3956 (N_3956,In_1679,In_425);
nor U3957 (N_3957,In_470,In_174);
or U3958 (N_3958,In_1201,In_63);
and U3959 (N_3959,In_805,In_969);
nand U3960 (N_3960,In_303,In_161);
or U3961 (N_3961,In_1692,In_1292);
nor U3962 (N_3962,In_1274,In_1109);
or U3963 (N_3963,In_1198,In_122);
nand U3964 (N_3964,In_834,In_1766);
nor U3965 (N_3965,In_1827,In_104);
xor U3966 (N_3966,In_1393,In_1542);
and U3967 (N_3967,In_1147,In_506);
nand U3968 (N_3968,In_760,In_1808);
and U3969 (N_3969,In_1931,In_195);
xor U3970 (N_3970,In_1515,In_1199);
or U3971 (N_3971,In_94,In_178);
nand U3972 (N_3972,In_880,In_1683);
and U3973 (N_3973,In_1546,In_873);
nand U3974 (N_3974,In_876,In_1336);
nand U3975 (N_3975,In_847,In_1200);
and U3976 (N_3976,In_198,In_104);
nor U3977 (N_3977,In_1889,In_962);
nand U3978 (N_3978,In_171,In_1453);
nor U3979 (N_3979,In_1407,In_528);
or U3980 (N_3980,In_1783,In_1430);
and U3981 (N_3981,In_474,In_715);
xor U3982 (N_3982,In_395,In_1290);
nand U3983 (N_3983,In_1920,In_1057);
xnor U3984 (N_3984,In_1129,In_1055);
and U3985 (N_3985,In_1389,In_1242);
nand U3986 (N_3986,In_1921,In_1300);
or U3987 (N_3987,In_1140,In_475);
xor U3988 (N_3988,In_1457,In_539);
nor U3989 (N_3989,In_1674,In_1613);
xor U3990 (N_3990,In_658,In_1519);
nor U3991 (N_3991,In_1905,In_1981);
xnor U3992 (N_3992,In_1015,In_428);
nor U3993 (N_3993,In_12,In_909);
and U3994 (N_3994,In_1604,In_1460);
or U3995 (N_3995,In_340,In_515);
xor U3996 (N_3996,In_1842,In_1844);
and U3997 (N_3997,In_1116,In_314);
nand U3998 (N_3998,In_1423,In_235);
xor U3999 (N_3999,In_914,In_1509);
xnor U4000 (N_4000,N_2438,N_427);
nor U4001 (N_4001,N_640,N_1041);
or U4002 (N_4002,N_1498,N_503);
xnor U4003 (N_4003,N_746,N_3297);
and U4004 (N_4004,N_465,N_1791);
or U4005 (N_4005,N_882,N_1625);
or U4006 (N_4006,N_3059,N_1114);
xnor U4007 (N_4007,N_2801,N_560);
and U4008 (N_4008,N_3236,N_2540);
nor U4009 (N_4009,N_647,N_2319);
xor U4010 (N_4010,N_1429,N_2283);
xor U4011 (N_4011,N_592,N_1242);
nand U4012 (N_4012,N_1239,N_1997);
nand U4013 (N_4013,N_2790,N_1620);
and U4014 (N_4014,N_3791,N_2094);
nor U4015 (N_4015,N_2033,N_275);
xor U4016 (N_4016,N_3692,N_2683);
nor U4017 (N_4017,N_1749,N_3591);
or U4018 (N_4018,N_3495,N_1070);
and U4019 (N_4019,N_167,N_1612);
nor U4020 (N_4020,N_998,N_970);
or U4021 (N_4021,N_2224,N_2492);
or U4022 (N_4022,N_2884,N_1712);
xor U4023 (N_4023,N_3090,N_3725);
and U4024 (N_4024,N_3604,N_729);
xnor U4025 (N_4025,N_3994,N_758);
and U4026 (N_4026,N_1998,N_3746);
or U4027 (N_4027,N_392,N_2309);
or U4028 (N_4028,N_3575,N_2610);
or U4029 (N_4029,N_1533,N_3909);
nand U4030 (N_4030,N_1435,N_691);
nor U4031 (N_4031,N_1300,N_1019);
or U4032 (N_4032,N_656,N_1484);
nor U4033 (N_4033,N_19,N_1021);
and U4034 (N_4034,N_1848,N_1146);
and U4035 (N_4035,N_1343,N_3112);
and U4036 (N_4036,N_303,N_1619);
xor U4037 (N_4037,N_1942,N_3846);
nand U4038 (N_4038,N_2418,N_1911);
or U4039 (N_4039,N_2975,N_122);
nor U4040 (N_4040,N_3427,N_1601);
or U4041 (N_4041,N_1390,N_3709);
nor U4042 (N_4042,N_3043,N_1076);
xor U4043 (N_4043,N_1072,N_3167);
nor U4044 (N_4044,N_3176,N_1787);
and U4045 (N_4045,N_80,N_788);
and U4046 (N_4046,N_3232,N_3129);
nand U4047 (N_4047,N_1876,N_3186);
nor U4048 (N_4048,N_2839,N_2205);
or U4049 (N_4049,N_147,N_519);
xnor U4050 (N_4050,N_2534,N_651);
or U4051 (N_4051,N_3408,N_1093);
xnor U4052 (N_4052,N_1884,N_938);
nand U4053 (N_4053,N_3126,N_3927);
or U4054 (N_4054,N_48,N_3060);
nor U4055 (N_4055,N_1843,N_2793);
and U4056 (N_4056,N_3263,N_1560);
nand U4057 (N_4057,N_3844,N_1388);
and U4058 (N_4058,N_1531,N_2302);
xor U4059 (N_4059,N_505,N_3109);
xor U4060 (N_4060,N_1077,N_1550);
or U4061 (N_4061,N_1565,N_3895);
nor U4062 (N_4062,N_452,N_3979);
and U4063 (N_4063,N_2417,N_1258);
nand U4064 (N_4064,N_2850,N_845);
nand U4065 (N_4065,N_2660,N_1815);
nor U4066 (N_4066,N_3985,N_2897);
nand U4067 (N_4067,N_856,N_1134);
and U4068 (N_4068,N_272,N_1264);
nand U4069 (N_4069,N_3269,N_2246);
xnor U4070 (N_4070,N_2297,N_1187);
nor U4071 (N_4071,N_2789,N_3945);
nand U4072 (N_4072,N_3758,N_1737);
nor U4073 (N_4073,N_289,N_3188);
or U4074 (N_4074,N_3726,N_634);
or U4075 (N_4075,N_1013,N_1663);
or U4076 (N_4076,N_2741,N_1925);
nand U4077 (N_4077,N_51,N_2366);
xor U4078 (N_4078,N_3564,N_3107);
nand U4079 (N_4079,N_388,N_1411);
nand U4080 (N_4080,N_1478,N_3634);
nand U4081 (N_4081,N_545,N_1744);
and U4082 (N_4082,N_3539,N_3125);
and U4083 (N_4083,N_3140,N_368);
and U4084 (N_4084,N_1852,N_2862);
and U4085 (N_4085,N_3192,N_2076);
or U4086 (N_4086,N_2405,N_2103);
xor U4087 (N_4087,N_2933,N_2112);
xnor U4088 (N_4088,N_688,N_237);
nor U4089 (N_4089,N_2983,N_2774);
nor U4090 (N_4090,N_1144,N_468);
or U4091 (N_4091,N_2653,N_3958);
xor U4092 (N_4092,N_2248,N_792);
or U4093 (N_4093,N_3750,N_2835);
or U4094 (N_4094,N_3077,N_3982);
or U4095 (N_4095,N_444,N_2035);
or U4096 (N_4096,N_236,N_1539);
xnor U4097 (N_4097,N_2692,N_3132);
nand U4098 (N_4098,N_294,N_512);
nor U4099 (N_4099,N_3893,N_1816);
and U4100 (N_4100,N_3199,N_1594);
nand U4101 (N_4101,N_3016,N_3870);
and U4102 (N_4102,N_2488,N_914);
nand U4103 (N_4103,N_736,N_508);
and U4104 (N_4104,N_937,N_3524);
or U4105 (N_4105,N_3550,N_3648);
nor U4106 (N_4106,N_2077,N_3926);
and U4107 (N_4107,N_1856,N_1129);
nand U4108 (N_4108,N_3312,N_457);
nand U4109 (N_4109,N_2649,N_3930);
nor U4110 (N_4110,N_105,N_2592);
and U4111 (N_4111,N_2082,N_1564);
xnor U4112 (N_4112,N_1424,N_2133);
and U4113 (N_4113,N_499,N_259);
nand U4114 (N_4114,N_2874,N_2397);
and U4115 (N_4115,N_2898,N_1222);
xor U4116 (N_4116,N_669,N_1382);
nand U4117 (N_4117,N_3617,N_2894);
and U4118 (N_4118,N_2546,N_2219);
and U4119 (N_4119,N_3589,N_386);
or U4120 (N_4120,N_1698,N_2819);
xor U4121 (N_4121,N_3385,N_3600);
nor U4122 (N_4122,N_3456,N_787);
xor U4123 (N_4123,N_3659,N_2731);
nand U4124 (N_4124,N_1004,N_1951);
nor U4125 (N_4125,N_1024,N_365);
xnor U4126 (N_4126,N_1198,N_2760);
nor U4127 (N_4127,N_2006,N_3625);
or U4128 (N_4128,N_293,N_836);
nand U4129 (N_4129,N_3742,N_438);
nand U4130 (N_4130,N_888,N_1631);
nor U4131 (N_4131,N_3511,N_2645);
xor U4132 (N_4132,N_3546,N_2221);
nand U4133 (N_4133,N_1888,N_1794);
and U4134 (N_4134,N_3688,N_2615);
and U4135 (N_4135,N_3466,N_1027);
nand U4136 (N_4136,N_2617,N_2415);
nor U4137 (N_4137,N_1551,N_606);
nand U4138 (N_4138,N_3204,N_65);
xnor U4139 (N_4139,N_20,N_751);
and U4140 (N_4140,N_3992,N_2034);
or U4141 (N_4141,N_927,N_3367);
xnor U4142 (N_4142,N_3538,N_3912);
xnor U4143 (N_4143,N_2114,N_1806);
and U4144 (N_4144,N_1895,N_672);
and U4145 (N_4145,N_2041,N_1523);
nor U4146 (N_4146,N_2486,N_2334);
nand U4147 (N_4147,N_1923,N_3485);
nand U4148 (N_4148,N_2730,N_614);
nand U4149 (N_4149,N_701,N_859);
nor U4150 (N_4150,N_1307,N_2456);
xor U4151 (N_4151,N_3697,N_1509);
nand U4152 (N_4152,N_1866,N_2644);
and U4153 (N_4153,N_153,N_715);
nand U4154 (N_4154,N_494,N_2202);
nor U4155 (N_4155,N_1012,N_1005);
and U4156 (N_4156,N_607,N_430);
and U4157 (N_4157,N_316,N_1814);
nor U4158 (N_4158,N_233,N_2542);
or U4159 (N_4159,N_1432,N_3028);
and U4160 (N_4160,N_87,N_3437);
nand U4161 (N_4161,N_1212,N_354);
nor U4162 (N_4162,N_1984,N_3464);
nand U4163 (N_4163,N_1172,N_1053);
or U4164 (N_4164,N_994,N_2588);
xor U4165 (N_4165,N_1635,N_1659);
xnor U4166 (N_4166,N_3598,N_111);
nand U4167 (N_4167,N_3151,N_3970);
or U4168 (N_4168,N_1955,N_2608);
nand U4169 (N_4169,N_1701,N_1147);
and U4170 (N_4170,N_2820,N_2066);
nand U4171 (N_4171,N_849,N_627);
xnor U4172 (N_4172,N_1930,N_1769);
nor U4173 (N_4173,N_3214,N_3250);
and U4174 (N_4174,N_3031,N_322);
nor U4175 (N_4175,N_234,N_3139);
and U4176 (N_4176,N_1610,N_690);
and U4177 (N_4177,N_828,N_2576);
xnor U4178 (N_4178,N_2565,N_570);
xnor U4179 (N_4179,N_2485,N_2721);
xnor U4180 (N_4180,N_3121,N_3620);
and U4181 (N_4181,N_3444,N_2704);
xnor U4182 (N_4182,N_3910,N_473);
and U4183 (N_4183,N_1628,N_247);
xnor U4184 (N_4184,N_3476,N_2938);
nor U4185 (N_4185,N_2152,N_1330);
nand U4186 (N_4186,N_1237,N_83);
and U4187 (N_4187,N_2264,N_2996);
nand U4188 (N_4188,N_969,N_1779);
and U4189 (N_4189,N_2009,N_3369);
or U4190 (N_4190,N_2395,N_2708);
and U4191 (N_4191,N_3148,N_588);
nand U4192 (N_4192,N_295,N_2869);
or U4193 (N_4193,N_2022,N_1125);
nor U4194 (N_4194,N_549,N_2362);
xor U4195 (N_4195,N_3002,N_38);
nand U4196 (N_4196,N_1753,N_1151);
nand U4197 (N_4197,N_531,N_3622);
xnor U4198 (N_4198,N_1195,N_674);
xnor U4199 (N_4199,N_3631,N_1571);
and U4200 (N_4200,N_3197,N_3790);
xnor U4201 (N_4201,N_3379,N_2055);
nand U4202 (N_4202,N_2904,N_3441);
or U4203 (N_4203,N_1099,N_243);
nand U4204 (N_4204,N_3527,N_3587);
or U4205 (N_4205,N_2343,N_2265);
and U4206 (N_4206,N_2437,N_3956);
nand U4207 (N_4207,N_1873,N_2177);
xor U4208 (N_4208,N_3545,N_2229);
nand U4209 (N_4209,N_2602,N_3265);
xor U4210 (N_4210,N_2183,N_2738);
nor U4211 (N_4211,N_2383,N_2075);
or U4212 (N_4212,N_1149,N_534);
and U4213 (N_4213,N_1243,N_3768);
or U4214 (N_4214,N_3718,N_3123);
and U4215 (N_4215,N_32,N_3235);
and U4216 (N_4216,N_2080,N_2315);
nor U4217 (N_4217,N_1689,N_1036);
or U4218 (N_4218,N_1494,N_3084);
xor U4219 (N_4219,N_741,N_802);
xor U4220 (N_4220,N_2794,N_2454);
xor U4221 (N_4221,N_832,N_2761);
and U4222 (N_4222,N_2915,N_2384);
xnor U4223 (N_4223,N_3057,N_2880);
nand U4224 (N_4224,N_2681,N_2155);
xnor U4225 (N_4225,N_2108,N_1621);
or U4226 (N_4226,N_328,N_3789);
and U4227 (N_4227,N_3405,N_5);
nor U4228 (N_4228,N_3158,N_271);
xor U4229 (N_4229,N_3997,N_3779);
and U4230 (N_4230,N_601,N_1169);
and U4231 (N_4231,N_3892,N_3344);
or U4232 (N_4232,N_2690,N_2331);
xor U4233 (N_4233,N_1765,N_2044);
nand U4234 (N_4234,N_267,N_3076);
nor U4235 (N_4235,N_3258,N_1685);
or U4236 (N_4236,N_694,N_2313);
nand U4237 (N_4237,N_2652,N_3515);
and U4238 (N_4238,N_2392,N_1810);
nand U4239 (N_4239,N_2266,N_3479);
and U4240 (N_4240,N_2157,N_3323);
or U4241 (N_4241,N_1600,N_3406);
or U4242 (N_4242,N_2040,N_1991);
nand U4243 (N_4243,N_3691,N_95);
and U4244 (N_4244,N_319,N_3829);
nor U4245 (N_4245,N_2491,N_2857);
nand U4246 (N_4246,N_2051,N_223);
nor U4247 (N_4247,N_2348,N_76);
or U4248 (N_4248,N_1104,N_873);
nand U4249 (N_4249,N_3488,N_460);
xnor U4250 (N_4250,N_266,N_3403);
nand U4251 (N_4251,N_3968,N_2256);
nor U4252 (N_4252,N_1812,N_2671);
and U4253 (N_4253,N_1965,N_1451);
xor U4254 (N_4254,N_3737,N_1073);
xnor U4255 (N_4255,N_3723,N_1651);
or U4256 (N_4256,N_1761,N_2502);
nor U4257 (N_4257,N_2647,N_2749);
xor U4258 (N_4258,N_171,N_769);
or U4259 (N_4259,N_2156,N_706);
or U4260 (N_4260,N_1842,N_3651);
and U4261 (N_4261,N_1361,N_3666);
xor U4262 (N_4262,N_1363,N_1047);
or U4263 (N_4263,N_2512,N_2840);
nand U4264 (N_4264,N_3954,N_1200);
xor U4265 (N_4265,N_2093,N_2633);
nor U4266 (N_4266,N_3357,N_2679);
or U4267 (N_4267,N_96,N_2030);
nand U4268 (N_4268,N_2352,N_1064);
xor U4269 (N_4269,N_113,N_799);
nand U4270 (N_4270,N_3509,N_0);
or U4271 (N_4271,N_3283,N_3044);
xor U4272 (N_4272,N_2797,N_1106);
xor U4273 (N_4273,N_3729,N_3243);
nand U4274 (N_4274,N_2402,N_2587);
and U4275 (N_4275,N_990,N_2198);
and U4276 (N_4276,N_1890,N_2976);
or U4277 (N_4277,N_1966,N_3594);
or U4278 (N_4278,N_14,N_834);
nor U4279 (N_4279,N_3834,N_3719);
and U4280 (N_4280,N_119,N_1287);
nor U4281 (N_4281,N_2187,N_1786);
xor U4282 (N_4282,N_3241,N_184);
nand U4283 (N_4283,N_1861,N_3608);
and U4284 (N_4284,N_3461,N_1249);
and U4285 (N_4285,N_2128,N_2665);
xnor U4286 (N_4286,N_1978,N_913);
xnor U4287 (N_4287,N_1098,N_3070);
xor U4288 (N_4288,N_2175,N_1720);
xor U4289 (N_4289,N_2934,N_399);
and U4290 (N_4290,N_3519,N_323);
xor U4291 (N_4291,N_2543,N_1774);
or U4292 (N_4292,N_16,N_1598);
xnor U4293 (N_4293,N_1975,N_3819);
nor U4294 (N_4294,N_3683,N_447);
or U4295 (N_4295,N_900,N_3096);
and U4296 (N_4296,N_2470,N_823);
nand U4297 (N_4297,N_1375,N_1870);
nor U4298 (N_4298,N_1556,N_2410);
nand U4299 (N_4299,N_126,N_2670);
nand U4300 (N_4300,N_3097,N_2712);
nand U4301 (N_4301,N_3083,N_2257);
nand U4302 (N_4302,N_2477,N_1480);
or U4303 (N_4303,N_860,N_3337);
xnor U4304 (N_4304,N_1583,N_3771);
nor U4305 (N_4305,N_455,N_2635);
nor U4306 (N_4306,N_3548,N_23);
nand U4307 (N_4307,N_890,N_976);
and U4308 (N_4308,N_3135,N_1026);
xnor U4309 (N_4309,N_3316,N_3430);
nand U4310 (N_4310,N_2432,N_2270);
nor U4311 (N_4311,N_3940,N_692);
nor U4312 (N_4312,N_1409,N_2784);
nor U4313 (N_4313,N_3439,N_3404);
nand U4314 (N_4314,N_719,N_2631);
or U4315 (N_4315,N_3510,N_2640);
nor U4316 (N_4316,N_619,N_2893);
and U4317 (N_4317,N_667,N_712);
or U4318 (N_4318,N_3517,N_22);
xnor U4319 (N_4319,N_3803,N_2988);
or U4320 (N_4320,N_2100,N_577);
and U4321 (N_4321,N_3676,N_3671);
xnor U4322 (N_4322,N_775,N_1949);
xnor U4323 (N_4323,N_3008,N_3917);
or U4324 (N_4324,N_2688,N_3003);
nand U4325 (N_4325,N_1735,N_624);
or U4326 (N_4326,N_1121,N_2012);
nand U4327 (N_4327,N_1183,N_3347);
xor U4328 (N_4328,N_2151,N_1223);
and U4329 (N_4329,N_1356,N_3629);
xor U4330 (N_4330,N_3303,N_3300);
nor U4331 (N_4331,N_2909,N_2255);
nor U4332 (N_4332,N_3313,N_3293);
or U4333 (N_4333,N_1437,N_894);
or U4334 (N_4334,N_1028,N_3583);
nor U4335 (N_4335,N_768,N_3436);
and U4336 (N_4336,N_2958,N_1405);
and U4337 (N_4337,N_1225,N_2249);
or U4338 (N_4338,N_2355,N_3766);
and U4339 (N_4339,N_1881,N_488);
nand U4340 (N_4340,N_1711,N_1383);
nand U4341 (N_4341,N_464,N_3655);
nand U4342 (N_4342,N_2911,N_1344);
xor U4343 (N_4343,N_2042,N_3396);
nand U4344 (N_4344,N_8,N_3784);
and U4345 (N_4345,N_1699,N_644);
and U4346 (N_4346,N_387,N_3939);
nor U4347 (N_4347,N_2131,N_1384);
xor U4348 (N_4348,N_2173,N_909);
nor U4349 (N_4349,N_2657,N_3864);
nor U4350 (N_4350,N_2337,N_2537);
nand U4351 (N_4351,N_1,N_1917);
or U4352 (N_4352,N_1700,N_3500);
or U4353 (N_4353,N_637,N_1760);
and U4354 (N_4354,N_2474,N_230);
or U4355 (N_4355,N_2772,N_2825);
xor U4356 (N_4356,N_2001,N_131);
and U4357 (N_4357,N_2335,N_2572);
nor U4358 (N_4358,N_1992,N_2902);
nor U4359 (N_4359,N_1194,N_540);
and U4360 (N_4360,N_3327,N_1033);
and U4361 (N_4361,N_1900,N_912);
or U4362 (N_4362,N_3134,N_1286);
nand U4363 (N_4363,N_60,N_2028);
or U4364 (N_4364,N_3179,N_3949);
nor U4365 (N_4365,N_1387,N_1639);
and U4366 (N_4366,N_824,N_3826);
or U4367 (N_4367,N_381,N_557);
nor U4368 (N_4368,N_2917,N_1416);
xor U4369 (N_4369,N_1441,N_889);
nor U4370 (N_4370,N_1426,N_2578);
nand U4371 (N_4371,N_1703,N_1574);
xnor U4372 (N_4372,N_1482,N_3908);
nor U4373 (N_4373,N_3266,N_2773);
and U4374 (N_4374,N_3682,N_1825);
nand U4375 (N_4375,N_684,N_1839);
nand U4376 (N_4376,N_3435,N_521);
nand U4377 (N_4377,N_2750,N_3628);
or U4378 (N_4378,N_1952,N_75);
nand U4379 (N_4379,N_3896,N_206);
or U4380 (N_4380,N_3644,N_1553);
and U4381 (N_4381,N_2725,N_1165);
xor U4382 (N_4382,N_853,N_2509);
nor U4383 (N_4383,N_64,N_917);
or U4384 (N_4384,N_1868,N_918);
nor U4385 (N_4385,N_3665,N_150);
xnor U4386 (N_4386,N_1575,N_825);
nor U4387 (N_4387,N_1788,N_86);
nor U4388 (N_4388,N_2827,N_925);
nand U4389 (N_4389,N_599,N_819);
nand U4390 (N_4390,N_2382,N_1609);
and U4391 (N_4391,N_309,N_377);
xnor U4392 (N_4392,N_2843,N_1479);
nand U4393 (N_4393,N_3547,N_2079);
nand U4394 (N_4394,N_1377,N_160);
and U4395 (N_4395,N_3014,N_1926);
nand U4396 (N_4396,N_1717,N_304);
and U4397 (N_4397,N_443,N_2398);
and U4398 (N_4398,N_161,N_2247);
and U4399 (N_4399,N_1813,N_1898);
nor U4400 (N_4400,N_3965,N_3049);
nand U4401 (N_4401,N_1702,N_821);
and U4402 (N_4402,N_3983,N_391);
or U4403 (N_4403,N_500,N_2826);
or U4404 (N_4404,N_2710,N_3760);
or U4405 (N_4405,N_3823,N_590);
or U4406 (N_4406,N_2928,N_1299);
and U4407 (N_4407,N_2081,N_3781);
nand U4408 (N_4408,N_3966,N_2083);
nand U4409 (N_4409,N_595,N_1419);
nand U4410 (N_4410,N_3695,N_1821);
nor U4411 (N_4411,N_2320,N_2465);
or U4412 (N_4412,N_1557,N_2788);
xnor U4413 (N_4413,N_3365,N_1905);
or U4414 (N_4414,N_3795,N_3732);
xnor U4415 (N_4415,N_1964,N_820);
nor U4416 (N_4416,N_1563,N_1323);
xnor U4417 (N_4417,N_612,N_1097);
xnor U4418 (N_4418,N_1181,N_3525);
or U4419 (N_4419,N_1935,N_1269);
and U4420 (N_4420,N_2955,N_1590);
xor U4421 (N_4421,N_1562,N_2207);
xnor U4422 (N_4422,N_2394,N_1453);
or U4423 (N_4423,N_3833,N_3001);
xnor U4424 (N_4424,N_1408,N_1155);
nand U4425 (N_4425,N_989,N_872);
xnor U4426 (N_4426,N_1246,N_2468);
and U4427 (N_4427,N_3880,N_489);
or U4428 (N_4428,N_831,N_1279);
or U4429 (N_4429,N_2853,N_3428);
nor U4430 (N_4430,N_1003,N_3041);
nand U4431 (N_4431,N_3331,N_2192);
and U4432 (N_4432,N_3005,N_2220);
or U4433 (N_4433,N_2935,N_1887);
xor U4434 (N_4434,N_2161,N_3413);
nand U4435 (N_4435,N_1337,N_2551);
nor U4436 (N_4436,N_1558,N_3017);
and U4437 (N_4437,N_2011,N_643);
nor U4438 (N_4438,N_1078,N_3552);
nand U4439 (N_4439,N_1745,N_2482);
and U4440 (N_4440,N_435,N_3494);
or U4441 (N_4441,N_1800,N_2686);
or U4442 (N_4442,N_2450,N_3046);
xnor U4443 (N_4443,N_3161,N_2966);
xor U4444 (N_4444,N_2144,N_3812);
xnor U4445 (N_4445,N_881,N_1948);
and U4446 (N_4446,N_2048,N_613);
xor U4447 (N_4447,N_1710,N_636);
xor U4448 (N_4448,N_2120,N_2185);
nor U4449 (N_4449,N_728,N_2792);
nor U4450 (N_4450,N_2882,N_1985);
xor U4451 (N_4451,N_255,N_3149);
nand U4452 (N_4452,N_527,N_1049);
nand U4453 (N_4453,N_1804,N_202);
or U4454 (N_4454,N_626,N_169);
nor U4455 (N_4455,N_2726,N_1986);
and U4456 (N_4456,N_2194,N_2550);
and U4457 (N_4457,N_79,N_176);
or U4458 (N_4458,N_3392,N_3577);
nand U4459 (N_4459,N_2707,N_3840);
nor U4460 (N_4460,N_2101,N_953);
and U4461 (N_4461,N_3556,N_52);
and U4462 (N_4462,N_1950,N_3424);
nand U4463 (N_4463,N_2324,N_1614);
and U4464 (N_4464,N_3409,N_1224);
and U4465 (N_4465,N_1874,N_2559);
and U4466 (N_4466,N_1537,N_3499);
nand U4467 (N_4467,N_164,N_3281);
nor U4468 (N_4468,N_1555,N_477);
and U4469 (N_4469,N_3287,N_311);
or U4470 (N_4470,N_300,N_1840);
nor U4471 (N_4471,N_2190,N_3289);
or U4472 (N_4472,N_2049,N_1213);
nand U4473 (N_4473,N_3417,N_3401);
xnor U4474 (N_4474,N_1379,N_697);
or U4475 (N_4475,N_3085,N_253);
xor U4476 (N_4476,N_3138,N_2733);
and U4477 (N_4477,N_911,N_562);
nand U4478 (N_4478,N_472,N_1595);
nand U4479 (N_4479,N_1492,N_988);
nand U4480 (N_4480,N_2922,N_3630);
xnor U4481 (N_4481,N_2732,N_497);
or U4482 (N_4482,N_1235,N_3662);
xnor U4483 (N_4483,N_3749,N_2282);
nor U4484 (N_4484,N_81,N_2703);
or U4485 (N_4485,N_1543,N_3118);
and U4486 (N_4486,N_2369,N_2879);
nor U4487 (N_4487,N_1807,N_1240);
nand U4488 (N_4488,N_2332,N_3035);
nand U4489 (N_4489,N_3251,N_179);
and U4490 (N_4490,N_458,N_3609);
or U4491 (N_4491,N_739,N_3573);
and U4492 (N_4492,N_916,N_3884);
nor U4493 (N_4493,N_550,N_3821);
xnor U4494 (N_4494,N_2664,N_1075);
and U4495 (N_4495,N_1878,N_2304);
xor U4496 (N_4496,N_2024,N_921);
and U4497 (N_4497,N_3114,N_2895);
or U4498 (N_4498,N_2498,N_3831);
and U4499 (N_4499,N_2627,N_783);
or U4500 (N_4500,N_1400,N_3980);
nor U4501 (N_4501,N_301,N_1939);
or U4502 (N_4502,N_593,N_3669);
nor U4503 (N_4503,N_1713,N_3861);
or U4504 (N_4504,N_2281,N_946);
nand U4505 (N_4505,N_2429,N_2501);
xor U4506 (N_4506,N_3291,N_3894);
or U4507 (N_4507,N_2518,N_718);
and U4508 (N_4508,N_2393,N_1420);
or U4509 (N_4509,N_2497,N_635);
and U4510 (N_4510,N_1116,N_31);
nand U4511 (N_4511,N_2691,N_454);
or U4512 (N_4512,N_1573,N_992);
nor U4513 (N_4513,N_3601,N_3371);
nor U4514 (N_4514,N_1896,N_3911);
nor U4515 (N_4515,N_2872,N_2696);
nand U4516 (N_4516,N_104,N_2629);
and U4517 (N_4517,N_1029,N_2778);
nand U4518 (N_4518,N_722,N_2193);
xor U4519 (N_4519,N_2052,N_1485);
xnor U4520 (N_4520,N_683,N_25);
and U4521 (N_4521,N_2122,N_1718);
nand U4522 (N_4522,N_3394,N_2566);
xor U4523 (N_4523,N_2804,N_2002);
and U4524 (N_4524,N_3411,N_603);
xnor U4525 (N_4525,N_2208,N_3168);
xnor U4526 (N_4526,N_547,N_3678);
or U4527 (N_4527,N_3730,N_663);
nor U4528 (N_4528,N_491,N_1746);
or U4529 (N_4529,N_1945,N_2541);
or U4530 (N_4530,N_2956,N_1273);
xnor U4531 (N_4531,N_3721,N_1616);
or U4532 (N_4532,N_2245,N_2285);
nor U4533 (N_4533,N_854,N_1291);
nand U4534 (N_4534,N_1002,N_1345);
and U4535 (N_4535,N_1389,N_1637);
nor U4536 (N_4536,N_1977,N_140);
xnor U4537 (N_4537,N_1739,N_3216);
nor U4538 (N_4538,N_954,N_2713);
and U4539 (N_4539,N_170,N_1442);
nand U4540 (N_4540,N_1646,N_187);
nor U4541 (N_4541,N_359,N_308);
nor U4542 (N_4542,N_2775,N_421);
or U4543 (N_4543,N_310,N_3777);
and U4544 (N_4544,N_241,N_70);
nor U4545 (N_4545,N_2702,N_1695);
nor U4546 (N_4546,N_1960,N_2735);
nand U4547 (N_4547,N_3815,N_1559);
xnor U4548 (N_4548,N_3217,N_210);
nand U4549 (N_4549,N_2206,N_717);
nor U4550 (N_4550,N_1381,N_3818);
and U4551 (N_4551,N_2025,N_3146);
nand U4552 (N_4552,N_1440,N_1906);
nand U4553 (N_4553,N_1270,N_3613);
and U4554 (N_4554,N_2036,N_2547);
nand U4555 (N_4555,N_1855,N_677);
nor U4556 (N_4556,N_2469,N_3885);
xor U4557 (N_4557,N_960,N_3866);
nor U4558 (N_4558,N_2848,N_3901);
nand U4559 (N_4559,N_496,N_3639);
and U4560 (N_4560,N_1582,N_2496);
and U4561 (N_4561,N_1056,N_1404);
nand U4562 (N_4562,N_671,N_3322);
nor U4563 (N_4563,N_3991,N_515);
xnor U4564 (N_4564,N_2717,N_878);
nor U4565 (N_4565,N_2411,N_1359);
or U4566 (N_4566,N_2182,N_895);
or U4567 (N_4567,N_1253,N_3969);
and U4568 (N_4568,N_476,N_933);
nand U4569 (N_4569,N_3673,N_1202);
nor U4570 (N_4570,N_3173,N_1941);
nand U4571 (N_4571,N_196,N_3822);
and U4572 (N_4572,N_2087,N_2701);
and U4573 (N_4573,N_3505,N_2597);
or U4574 (N_4574,N_811,N_395);
xnor U4575 (N_4575,N_567,N_3883);
xor U4576 (N_4576,N_2176,N_173);
or U4577 (N_4577,N_1785,N_3452);
nor U4578 (N_4578,N_3213,N_867);
xnor U4579 (N_4579,N_797,N_317);
nor U4580 (N_4580,N_3948,N_1422);
nand U4581 (N_4581,N_805,N_1386);
and U4582 (N_4582,N_257,N_1841);
nand U4583 (N_4583,N_3025,N_1305);
xnor U4584 (N_4584,N_3256,N_416);
or U4585 (N_4585,N_1694,N_632);
xnor U4586 (N_4586,N_2489,N_2997);
nor U4587 (N_4587,N_3030,N_3332);
nor U4588 (N_4588,N_2923,N_2232);
and U4589 (N_4589,N_3015,N_2507);
xor U4590 (N_4590,N_1122,N_945);
nand U4591 (N_4591,N_3414,N_276);
and U4592 (N_4592,N_268,N_2471);
nand U4593 (N_4593,N_3679,N_436);
nor U4594 (N_4594,N_2737,N_3722);
xnor U4595 (N_4595,N_1524,N_2329);
or U4596 (N_4596,N_1642,N_3951);
nand U4597 (N_4597,N_629,N_361);
nor U4598 (N_4598,N_1335,N_1062);
or U4599 (N_4599,N_848,N_2296);
or U4600 (N_4600,N_3599,N_1820);
nand U4601 (N_4601,N_3649,N_3817);
nand U4602 (N_4602,N_3947,N_535);
xor U4603 (N_4603,N_1090,N_3443);
xor U4604 (N_4604,N_958,N_2333);
nor U4605 (N_4605,N_190,N_1088);
nand U4606 (N_4606,N_2699,N_3971);
xnor U4607 (N_4607,N_3504,N_3879);
or U4608 (N_4608,N_3806,N_3916);
nor U4609 (N_4609,N_2783,N_1293);
xor U4610 (N_4610,N_2057,N_3486);
and U4611 (N_4611,N_941,N_2650);
nor U4612 (N_4612,N_1133,N_2399);
nor U4613 (N_4613,N_935,N_551);
nor U4614 (N_4614,N_984,N_2231);
and U4615 (N_4615,N_2341,N_2213);
nor U4616 (N_4616,N_733,N_2912);
nand U4617 (N_4617,N_2866,N_3194);
nand U4618 (N_4618,N_1452,N_49);
nor U4619 (N_4619,N_1466,N_1350);
xnor U4620 (N_4620,N_1446,N_2388);
nand U4621 (N_4621,N_520,N_481);
or U4622 (N_4622,N_659,N_940);
or U4623 (N_4623,N_3259,N_3626);
nand U4624 (N_4624,N_2865,N_808);
and U4625 (N_4625,N_760,N_302);
nand U4626 (N_4626,N_2045,N_863);
nand U4627 (N_4627,N_763,N_333);
nand U4628 (N_4628,N_2724,N_681);
xnor U4629 (N_4629,N_286,N_2558);
nor U4630 (N_4630,N_3101,N_1636);
and U4631 (N_4631,N_1140,N_68);
or U4632 (N_4632,N_1436,N_2969);
and U4633 (N_4633,N_199,N_1901);
nor U4634 (N_4634,N_2799,N_1781);
and U4635 (N_4635,N_696,N_1245);
and U4636 (N_4636,N_3851,N_3660);
and U4637 (N_4637,N_2505,N_389);
nand U4638 (N_4638,N_3147,N_415);
nand U4639 (N_4639,N_3307,N_2770);
nor U4640 (N_4640,N_509,N_2624);
xnor U4641 (N_4641,N_2163,N_3953);
xor U4642 (N_4642,N_2407,N_3257);
xor U4643 (N_4643,N_3382,N_923);
nand U4644 (N_4644,N_3531,N_1506);
and U4645 (N_4645,N_1561,N_1265);
xor U4646 (N_4646,N_2330,N_291);
xor U4647 (N_4647,N_1988,N_3207);
nand U4648 (N_4648,N_2225,N_380);
or U4649 (N_4649,N_2169,N_133);
nor U4650 (N_4650,N_3597,N_695);
xor U4651 (N_4651,N_3612,N_581);
nand U4652 (N_4652,N_2073,N_1758);
xnor U4653 (N_4653,N_1068,N_2714);
xor U4654 (N_4654,N_1398,N_1417);
nand U4655 (N_4655,N_1283,N_922);
nand U4656 (N_4656,N_327,N_1185);
nor U4657 (N_4657,N_3280,N_2885);
nand U4658 (N_4658,N_579,N_752);
and U4659 (N_4659,N_2963,N_822);
or U4660 (N_4660,N_2029,N_2287);
nand U4661 (N_4661,N_88,N_2435);
and U4662 (N_4662,N_2729,N_2557);
or U4663 (N_4663,N_2372,N_1714);
and U4664 (N_4664,N_3352,N_3145);
nand U4665 (N_4665,N_1357,N_3735);
nor U4666 (N_4666,N_3963,N_3934);
nand U4667 (N_4667,N_1678,N_1725);
and U4668 (N_4668,N_62,N_724);
xnor U4669 (N_4669,N_633,N_1011);
and U4670 (N_4670,N_3560,N_2416);
xor U4671 (N_4671,N_2971,N_1038);
or U4672 (N_4672,N_1863,N_3462);
nor U4673 (N_4673,N_3715,N_2360);
nand U4674 (N_4674,N_229,N_2476);
or U4675 (N_4675,N_3453,N_138);
xnor U4676 (N_4676,N_564,N_1880);
and U4677 (N_4677,N_3984,N_628);
xnor U4678 (N_4678,N_1000,N_1633);
and U4679 (N_4679,N_1394,N_1458);
nor U4680 (N_4680,N_245,N_1274);
xor U4681 (N_4681,N_1414,N_3032);
nand U4682 (N_4682,N_1535,N_1728);
xor U4683 (N_4683,N_2046,N_1660);
and U4684 (N_4684,N_1163,N_1094);
or U4685 (N_4685,N_3026,N_798);
nor U4686 (N_4686,N_639,N_2449);
nor U4687 (N_4687,N_950,N_866);
and U4688 (N_4688,N_3778,N_2186);
nand U4689 (N_4689,N_1693,N_1358);
and U4690 (N_4690,N_2237,N_2223);
nand U4691 (N_4691,N_865,N_1092);
and U4692 (N_4692,N_2727,N_3596);
or U4693 (N_4693,N_3751,N_2965);
and U4694 (N_4694,N_1792,N_11);
or U4695 (N_4695,N_2995,N_1707);
xor U4696 (N_4696,N_3239,N_2196);
xor U4697 (N_4697,N_1516,N_3136);
nand U4698 (N_4698,N_215,N_3324);
or U4699 (N_4699,N_1160,N_2104);
nand U4700 (N_4700,N_1327,N_216);
xor U4701 (N_4701,N_3553,N_375);
and U4702 (N_4702,N_3460,N_1921);
nor U4703 (N_4703,N_98,N_1467);
or U4704 (N_4704,N_55,N_3388);
or U4705 (N_4705,N_2986,N_1643);
nand U4706 (N_4706,N_279,N_971);
or U4707 (N_4707,N_2178,N_1204);
nand U4708 (N_4708,N_123,N_3182);
or U4709 (N_4709,N_3633,N_782);
nor U4710 (N_4710,N_2243,N_3481);
nand U4711 (N_4711,N_1290,N_2317);
nor U4712 (N_4712,N_3584,N_3640);
xor U4713 (N_4713,N_2503,N_2630);
or U4714 (N_4714,N_326,N_1503);
nand U4715 (N_4715,N_3804,N_3876);
nor U4716 (N_4716,N_3807,N_871);
or U4717 (N_4717,N_2216,N_3811);
or U4718 (N_4718,N_2621,N_3995);
xor U4719 (N_4719,N_966,N_1970);
nor U4720 (N_4720,N_3580,N_2236);
nor U4721 (N_4721,N_2562,N_470);
nor U4722 (N_4722,N_3459,N_2387);
nand U4723 (N_4723,N_1406,N_641);
and U4724 (N_4724,N_1837,N_3616);
and U4725 (N_4725,N_679,N_1830);
and U4726 (N_4726,N_2188,N_919);
nor U4727 (N_4727,N_1241,N_1741);
and U4728 (N_4728,N_3386,N_3295);
nor U4729 (N_4729,N_1250,N_1464);
xor U4730 (N_4730,N_565,N_3402);
or U4731 (N_4731,N_2278,N_397);
or U4732 (N_4732,N_1339,N_3929);
xor U4733 (N_4733,N_3802,N_41);
and U4734 (N_4734,N_1757,N_3105);
and U4735 (N_4735,N_2117,N_163);
xor U4736 (N_4736,N_3931,N_1111);
nand U4737 (N_4737,N_1180,N_351);
xor U4738 (N_4738,N_1534,N_3117);
and U4739 (N_4739,N_2127,N_1943);
nor U4740 (N_4740,N_3825,N_1139);
and U4741 (N_4741,N_2831,N_115);
xor U4742 (N_4742,N_1336,N_2697);
and U4743 (N_4743,N_1278,N_2504);
or U4744 (N_4744,N_2179,N_3805);
and U4745 (N_4745,N_1261,N_3272);
nor U4746 (N_4746,N_1538,N_1459);
nor U4747 (N_4747,N_1704,N_2089);
and U4748 (N_4748,N_1010,N_2218);
or U4749 (N_4749,N_3429,N_1851);
xnor U4750 (N_4750,N_412,N_1530);
and U4751 (N_4751,N_985,N_46);
and U4752 (N_4752,N_3753,N_2636);
nand U4753 (N_4753,N_3890,N_2531);
and U4754 (N_4754,N_1510,N_1367);
or U4755 (N_4755,N_3063,N_256);
xor U4756 (N_4756,N_3492,N_3317);
or U4757 (N_4757,N_2942,N_3950);
or U4758 (N_4758,N_2068,N_2782);
xnor U4759 (N_4759,N_2740,N_2426);
nor U4760 (N_4760,N_2159,N_3582);
nor U4761 (N_4761,N_3023,N_217);
nor U4762 (N_4762,N_2460,N_3776);
and U4763 (N_4763,N_2555,N_621);
and U4764 (N_4764,N_2300,N_56);
nor U4765 (N_4765,N_670,N_522);
nand U4766 (N_4766,N_3624,N_2069);
nand U4767 (N_4767,N_1117,N_2619);
nand U4768 (N_4768,N_2867,N_44);
nor U4769 (N_4769,N_3038,N_432);
xnor U4770 (N_4770,N_2462,N_1309);
and U4771 (N_4771,N_1673,N_574);
and U4772 (N_4772,N_3702,N_1476);
and U4773 (N_4773,N_623,N_2200);
nor U4774 (N_4774,N_1924,N_942);
and U4775 (N_4775,N_3184,N_1681);
and U4776 (N_4776,N_1006,N_3863);
nor U4777 (N_4777,N_2181,N_558);
xnor U4778 (N_4778,N_439,N_1128);
or U4779 (N_4779,N_3716,N_3978);
nand U4780 (N_4780,N_977,N_2845);
nor U4781 (N_4781,N_2342,N_1764);
nand U4782 (N_4782,N_1871,N_2085);
or U4783 (N_4783,N_2201,N_765);
nor U4784 (N_4784,N_148,N_2716);
nand U4785 (N_4785,N_149,N_47);
xor U4786 (N_4786,N_1326,N_1465);
xor U4787 (N_4787,N_582,N_142);
nor U4788 (N_4788,N_3021,N_1412);
xnor U4789 (N_4789,N_382,N_1944);
nor U4790 (N_4790,N_1392,N_3690);
and U4791 (N_4791,N_2595,N_2318);
nor U4792 (N_4792,N_778,N_3793);
nor U4793 (N_4793,N_3254,N_1802);
nor U4794 (N_4794,N_3473,N_2091);
and U4795 (N_4795,N_1922,N_1691);
and U4796 (N_4796,N_2259,N_2058);
and U4797 (N_4797,N_1447,N_3588);
nor U4798 (N_4798,N_1164,N_118);
nand U4799 (N_4799,N_3451,N_3530);
or U4800 (N_4800,N_1074,N_3391);
and U4801 (N_4801,N_3273,N_906);
nor U4802 (N_4802,N_466,N_3286);
nor U4803 (N_4803,N_1497,N_110);
or U4804 (N_4804,N_3062,N_3472);
or U4805 (N_4805,N_2916,N_3302);
or U4806 (N_4806,N_3503,N_693);
and U4807 (N_4807,N_1910,N_2147);
or U4808 (N_4808,N_510,N_703);
or U4809 (N_4809,N_883,N_1971);
nor U4810 (N_4810,N_3946,N_2768);
or U4811 (N_4811,N_598,N_2135);
nor U4812 (N_4812,N_3048,N_2389);
nand U4813 (N_4813,N_1057,N_1366);
nand U4814 (N_4814,N_1566,N_968);
and U4815 (N_4815,N_930,N_1322);
and U4816 (N_4816,N_3706,N_1415);
or U4817 (N_4817,N_467,N_3421);
nand U4818 (N_4818,N_2808,N_3009);
nor U4819 (N_4819,N_2623,N_373);
nor U4820 (N_4820,N_2682,N_1238);
xor U4821 (N_4821,N_3474,N_2153);
nor U4822 (N_4822,N_2575,N_2875);
nand U4823 (N_4823,N_885,N_3657);
nor U4824 (N_4824,N_1502,N_1203);
nor U4825 (N_4825,N_1762,N_3229);
nor U4826 (N_4826,N_3534,N_3832);
or U4827 (N_4827,N_195,N_3252);
or U4828 (N_4828,N_1969,N_1067);
xnor U4829 (N_4829,N_3398,N_3094);
or U4830 (N_4830,N_1589,N_2585);
or U4831 (N_4831,N_3809,N_3618);
nand U4832 (N_4832,N_666,N_1836);
xnor U4833 (N_4833,N_615,N_3296);
or U4834 (N_4834,N_2299,N_3423);
nand U4835 (N_4835,N_3319,N_144);
or U4836 (N_4836,N_15,N_1471);
xor U4837 (N_4837,N_2288,N_3786);
xor U4838 (N_4838,N_3738,N_242);
and U4839 (N_4839,N_1544,N_2763);
nor U4840 (N_4840,N_1674,N_3990);
or U4841 (N_4841,N_2579,N_1919);
xor U4842 (N_4842,N_3810,N_1044);
xnor U4843 (N_4843,N_936,N_742);
and U4844 (N_4844,N_2800,N_2124);
nor U4845 (N_4845,N_1727,N_109);
and U4846 (N_4846,N_1191,N_967);
nor U4847 (N_4847,N_3103,N_2620);
or U4848 (N_4848,N_3087,N_3073);
nand U4849 (N_4849,N_2071,N_2940);
nand U4850 (N_4850,N_1031,N_1570);
nand U4851 (N_4851,N_3837,N_2110);
nor U4852 (N_4852,N_1995,N_1529);
nor U4853 (N_4853,N_3568,N_3128);
nand U4854 (N_4854,N_2158,N_720);
xor U4855 (N_4855,N_1679,N_3852);
nor U4856 (N_4856,N_2227,N_2115);
nor U4857 (N_4857,N_2292,N_1161);
nand U4858 (N_4858,N_1540,N_1607);
xnor U4859 (N_4859,N_471,N_2828);
nand U4860 (N_4860,N_3514,N_1522);
nand U4861 (N_4861,N_107,N_2849);
nor U4862 (N_4862,N_886,N_2648);
nor U4863 (N_4863,N_2746,N_2212);
nand U4864 (N_4864,N_2,N_61);
or U4865 (N_4865,N_89,N_1796);
nor U4866 (N_4866,N_3838,N_3675);
nor U4867 (N_4867,N_3349,N_2053);
nand U4868 (N_4868,N_846,N_2408);
and U4869 (N_4869,N_1159,N_3362);
or U4870 (N_4870,N_2817,N_1298);
and U4871 (N_4871,N_2346,N_1899);
nand U4872 (N_4872,N_273,N_3871);
and U4873 (N_4873,N_1495,N_2753);
or U4874 (N_4874,N_1719,N_3308);
nor U4875 (N_4875,N_1940,N_2569);
nand U4876 (N_4876,N_2172,N_3000);
or U4877 (N_4877,N_575,N_563);
nor U4878 (N_4878,N_3080,N_3981);
nor U4879 (N_4879,N_2998,N_1023);
or U4880 (N_4880,N_1214,N_2695);
and U4881 (N_4881,N_194,N_3226);
nand U4882 (N_4882,N_2291,N_3033);
and U4883 (N_4883,N_3843,N_3468);
xor U4884 (N_4884,N_1578,N_71);
nand U4885 (N_4885,N_3928,N_665);
and U4886 (N_4886,N_710,N_112);
and U4887 (N_4887,N_1664,N_3841);
xor U4888 (N_4888,N_999,N_1552);
nor U4889 (N_4889,N_1216,N_3882);
xnor U4890 (N_4890,N_2589,N_3449);
nor U4891 (N_4891,N_1475,N_2254);
nor U4892 (N_4892,N_239,N_2890);
xnor U4893 (N_4893,N_3165,N_1108);
and U4894 (N_4894,N_2038,N_3152);
and U4895 (N_4895,N_2994,N_3193);
nand U4896 (N_4896,N_3366,N_1082);
and U4897 (N_4897,N_837,N_3794);
nand U4898 (N_4898,N_1050,N_36);
or U4899 (N_4899,N_3915,N_1188);
nand U4900 (N_4900,N_3681,N_2345);
nor U4901 (N_4901,N_2628,N_2279);
or U4902 (N_4902,N_1095,N_2891);
nand U4903 (N_4903,N_1897,N_3333);
or U4904 (N_4904,N_2240,N_905);
nand U4905 (N_4905,N_784,N_2706);
xor U4906 (N_4906,N_2074,N_374);
nand U4907 (N_4907,N_541,N_1834);
or U4908 (N_4908,N_2021,N_222);
xnor U4909 (N_4909,N_1795,N_1507);
nor U4910 (N_4910,N_3471,N_3482);
or U4911 (N_4911,N_858,N_934);
or U4912 (N_4912,N_1775,N_287);
or U4913 (N_4913,N_2832,N_1624);
and U4914 (N_4914,N_986,N_248);
or U4915 (N_4915,N_2349,N_225);
nand U4916 (N_4916,N_1933,N_2339);
nand U4917 (N_4917,N_2250,N_812);
and U4918 (N_4918,N_2480,N_2930);
nand U4919 (N_4919,N_2719,N_3318);
xor U4920 (N_4920,N_1962,N_662);
nor U4921 (N_4921,N_3074,N_1931);
xor U4922 (N_4922,N_2374,N_3743);
or U4923 (N_4923,N_995,N_1915);
and U4924 (N_4924,N_341,N_1665);
nor U4925 (N_4925,N_2642,N_983);
xor U4926 (N_4926,N_3434,N_972);
xnor U4927 (N_4927,N_2211,N_2413);
nor U4928 (N_4928,N_422,N_2043);
and U4929 (N_4929,N_2228,N_2209);
or U4930 (N_4930,N_2892,N_2581);
or U4931 (N_4931,N_3244,N_2371);
nand U4932 (N_4932,N_28,N_2422);
xnor U4933 (N_4933,N_3972,N_1773);
or U4934 (N_4934,N_1182,N_771);
nor U4935 (N_4935,N_3763,N_3565);
xor U4936 (N_4936,N_3065,N_610);
xnor U4937 (N_4937,N_1680,N_502);
xor U4938 (N_4938,N_1135,N_495);
nor U4939 (N_4939,N_3516,N_9);
xnor U4940 (N_4940,N_2412,N_789);
or U4941 (N_4941,N_2325,N_1512);
and U4942 (N_4942,N_3467,N_3656);
nor U4943 (N_4943,N_1219,N_2638);
and U4944 (N_4944,N_77,N_1981);
xnor U4945 (N_4945,N_3942,N_3395);
nor U4946 (N_4946,N_1101,N_3341);
nand U4947 (N_4947,N_3034,N_3569);
xnor U4948 (N_4948,N_1109,N_2752);
or U4949 (N_4949,N_91,N_1173);
nand U4950 (N_4950,N_3373,N_3567);
nand U4951 (N_4951,N_2105,N_973);
xor U4952 (N_4952,N_532,N_2459);
xor U4953 (N_4953,N_2390,N_2600);
xnor U4954 (N_4954,N_2959,N_2481);
nor U4955 (N_4955,N_2166,N_862);
nor U4956 (N_4956,N_673,N_794);
nand U4957 (N_4957,N_3667,N_3571);
nor U4958 (N_4958,N_810,N_3198);
nor U4959 (N_4959,N_616,N_3309);
xor U4960 (N_4960,N_1771,N_2618);
or U4961 (N_4961,N_332,N_364);
and U4962 (N_4962,N_2979,N_3240);
xnor U4963 (N_4963,N_2858,N_2092);
nor U4964 (N_4964,N_3202,N_2072);
xor U4965 (N_4965,N_2993,N_1328);
and U4966 (N_4966,N_285,N_1016);
nand U4967 (N_4967,N_1818,N_3739);
and U4968 (N_4968,N_3636,N_699);
and U4969 (N_4969,N_2563,N_3542);
or U4970 (N_4970,N_2170,N_738);
or U4971 (N_4971,N_137,N_2810);
nand U4972 (N_4972,N_2625,N_490);
xor U4973 (N_4973,N_3705,N_2098);
or U4974 (N_4974,N_3611,N_1127);
or U4975 (N_4975,N_2121,N_136);
xnor U4976 (N_4976,N_1145,N_431);
nand U4977 (N_4977,N_1083,N_1190);
or U4978 (N_4978,N_2373,N_868);
nand U4979 (N_4979,N_1425,N_504);
nand U4980 (N_4980,N_2180,N_2655);
or U4981 (N_4981,N_337,N_749);
nor U4982 (N_4982,N_42,N_1706);
xnor U4983 (N_4983,N_3171,N_631);
xor U4984 (N_4984,N_3680,N_2948);
or U4985 (N_4985,N_1979,N_2567);
and U4986 (N_4986,N_2943,N_3433);
and U4987 (N_4987,N_731,N_2500);
xor U4988 (N_4988,N_1845,N_1644);
and U4989 (N_4989,N_2146,N_3210);
and U4990 (N_4990,N_660,N_3508);
or U4991 (N_4991,N_209,N_3875);
nand U4992 (N_4992,N_1341,N_3974);
or U4993 (N_4993,N_3554,N_1705);
nor U4994 (N_4994,N_1894,N_826);
nand U4995 (N_4995,N_3234,N_3551);
or U4996 (N_4996,N_3201,N_1864);
xor U4997 (N_4997,N_2574,N_1811);
nand U4998 (N_4998,N_2791,N_1107);
xnor U4999 (N_4999,N_3342,N_344);
xnor U5000 (N_5000,N_143,N_1913);
nor U5001 (N_5001,N_604,N_2375);
or U5002 (N_5002,N_3338,N_2409);
xnor U5003 (N_5003,N_3220,N_2980);
nand U5004 (N_5004,N_2129,N_1597);
nand U5005 (N_5005,N_518,N_325);
nor U5006 (N_5006,N_3724,N_2675);
or U5007 (N_5007,N_1937,N_1311);
and U5008 (N_5008,N_246,N_2945);
or U5009 (N_5009,N_1572,N_1835);
or U5010 (N_5010,N_843,N_1100);
and U5011 (N_5011,N_3976,N_2106);
and U5012 (N_5012,N_2705,N_2967);
and U5013 (N_5013,N_372,N_1872);
and U5014 (N_5014,N_3769,N_3627);
nor U5015 (N_5015,N_2593,N_1677);
and U5016 (N_5016,N_1008,N_3796);
nor U5017 (N_5017,N_1670,N_192);
nand U5018 (N_5018,N_3491,N_2992);
nand U5019 (N_5019,N_1176,N_1687);
nor U5020 (N_5020,N_3445,N_1039);
or U5021 (N_5021,N_2367,N_2549);
nor U5022 (N_5022,N_1828,N_1374);
nand U5023 (N_5023,N_1653,N_90);
nand U5024 (N_5024,N_406,N_770);
nand U5025 (N_5025,N_191,N_3187);
and U5026 (N_5026,N_646,N_1355);
and U5027 (N_5027,N_2174,N_2358);
and U5028 (N_5028,N_3734,N_321);
and U5029 (N_5029,N_3906,N_3006);
or U5030 (N_5030,N_152,N_1058);
and U5031 (N_5031,N_3231,N_159);
xor U5032 (N_5032,N_120,N_2487);
or U5033 (N_5033,N_445,N_3013);
or U5034 (N_5034,N_66,N_3164);
and U5035 (N_5035,N_400,N_1805);
and U5036 (N_5036,N_1470,N_3455);
nand U5037 (N_5037,N_3785,N_2918);
xnor U5038 (N_5038,N_2856,N_2088);
and U5039 (N_5039,N_200,N_721);
or U5040 (N_5040,N_1654,N_2064);
nor U5041 (N_5041,N_2814,N_1192);
nor U5042 (N_5042,N_2767,N_2026);
and U5043 (N_5043,N_3012,N_2957);
or U5044 (N_5044,N_734,N_97);
nor U5045 (N_5045,N_3813,N_3100);
xor U5046 (N_5046,N_2637,N_1832);
and U5047 (N_5047,N_1916,N_158);
nor U5048 (N_5048,N_589,N_2654);
nor U5049 (N_5049,N_657,N_737);
xnor U5050 (N_5050,N_429,N_3212);
nor U5051 (N_5051,N_3221,N_3881);
xor U5052 (N_5052,N_1726,N_448);
nor U5053 (N_5053,N_2328,N_1882);
xnor U5054 (N_5054,N_530,N_1790);
nor U5055 (N_5055,N_965,N_2913);
xnor U5056 (N_5056,N_1032,N_1527);
nand U5057 (N_5057,N_1611,N_45);
xnor U5058 (N_5058,N_3311,N_182);
xor U5059 (N_5059,N_3581,N_3288);
xnor U5060 (N_5060,N_3855,N_2883);
xnor U5061 (N_5061,N_709,N_2344);
nand U5062 (N_5062,N_3330,N_3507);
xor U5063 (N_5063,N_516,N_3069);
or U5064 (N_5064,N_1740,N_1743);
nor U5065 (N_5065,N_3068,N_602);
or U5066 (N_5066,N_1648,N_2852);
nor U5067 (N_5067,N_1581,N_2510);
nand U5068 (N_5068,N_1634,N_483);
or U5069 (N_5069,N_1376,N_3326);
nor U5070 (N_5070,N_1953,N_2634);
nor U5071 (N_5071,N_2453,N_410);
nor U5072 (N_5072,N_1647,N_3416);
or U5073 (N_5073,N_3498,N_252);
nand U5074 (N_5074,N_2661,N_2556);
nor U5075 (N_5075,N_777,N_1084);
nor U5076 (N_5076,N_2973,N_213);
nand U5077 (N_5077,N_2921,N_1857);
nand U5078 (N_5078,N_2261,N_437);
and U5079 (N_5079,N_263,N_2520);
and U5080 (N_5080,N_1481,N_1865);
nor U5081 (N_5081,N_398,N_1656);
nand U5082 (N_5082,N_2924,N_1640);
nand U5083 (N_5083,N_1448,N_1059);
nor U5084 (N_5084,N_1826,N_413);
nand U5085 (N_5085,N_951,N_2596);
xor U5086 (N_5086,N_3661,N_3081);
nand U5087 (N_5087,N_1846,N_2722);
nand U5088 (N_5088,N_1468,N_2356);
nand U5089 (N_5089,N_1875,N_1957);
nor U5090 (N_5090,N_1672,N_299);
nor U5091 (N_5091,N_1879,N_2286);
nand U5092 (N_5092,N_482,N_944);
and U5093 (N_5093,N_2583,N_13);
nand U5094 (N_5094,N_73,N_1528);
nor U5095 (N_5095,N_1596,N_3393);
nor U5096 (N_5096,N_2434,N_33);
and U5097 (N_5097,N_3720,N_383);
or U5098 (N_5098,N_2765,N_861);
nand U5099 (N_5099,N_1577,N_2338);
nor U5100 (N_5100,N_2561,N_2787);
and U5101 (N_5101,N_1909,N_1267);
or U5102 (N_5102,N_1742,N_3944);
or U5103 (N_5103,N_680,N_753);
nor U5104 (N_5104,N_101,N_561);
xor U5105 (N_5105,N_3808,N_2946);
nor U5106 (N_5106,N_3205,N_459);
or U5107 (N_5107,N_2007,N_517);
xor U5108 (N_5108,N_997,N_2906);
xnor U5109 (N_5109,N_2210,N_2864);
and U5110 (N_5110,N_2267,N_2479);
nand U5111 (N_5111,N_630,N_586);
or U5112 (N_5112,N_3770,N_2364);
or U5113 (N_5113,N_1220,N_1054);
or U5114 (N_5114,N_114,N_3113);
and U5115 (N_5115,N_801,N_2233);
xnor U5116 (N_5116,N_884,N_139);
or U5117 (N_5117,N_3108,N_2798);
xnor U5118 (N_5118,N_2689,N_2926);
nand U5119 (N_5119,N_3011,N_424);
nand U5120 (N_5120,N_800,N_2779);
and U5121 (N_5121,N_2191,N_879);
xor U5122 (N_5122,N_165,N_689);
xor U5123 (N_5123,N_3209,N_1929);
or U5124 (N_5124,N_2251,N_2316);
nor U5125 (N_5125,N_3036,N_3772);
nor U5126 (N_5126,N_2611,N_1372);
and U5127 (N_5127,N_2747,N_2548);
and U5128 (N_5128,N_1903,N_2919);
or U5129 (N_5129,N_3166,N_585);
nor U5130 (N_5130,N_2613,N_1584);
nand U5131 (N_5131,N_3279,N_1158);
nor U5132 (N_5132,N_3095,N_3356);
nand U5133 (N_5133,N_3952,N_1902);
nand U5134 (N_5134,N_2658,N_3004);
nor U5135 (N_5135,N_2162,N_3438);
nor U5136 (N_5136,N_3731,N_1276);
xnor U5137 (N_5137,N_3579,N_3960);
nand U5138 (N_5138,N_3361,N_3304);
nand U5139 (N_5139,N_3714,N_201);
xnor U5140 (N_5140,N_3765,N_1315);
nand U5141 (N_5141,N_2844,N_2522);
nand U5142 (N_5142,N_3222,N_851);
and U5143 (N_5143,N_2901,N_3228);
and U5144 (N_5144,N_813,N_3938);
nor U5145 (N_5145,N_855,N_3701);
and U5146 (N_5146,N_1410,N_2441);
nor U5147 (N_5147,N_975,N_2903);
nor U5148 (N_5148,N_2813,N_102);
nand U5149 (N_5149,N_1738,N_1605);
nand U5150 (N_5150,N_2841,N_2443);
nor U5151 (N_5151,N_3354,N_3741);
or U5152 (N_5152,N_2954,N_3206);
nor U5153 (N_5153,N_1370,N_3578);
xnor U5154 (N_5154,N_352,N_1354);
or U5155 (N_5155,N_1171,N_278);
and U5156 (N_5156,N_3450,N_1487);
xor U5157 (N_5157,N_618,N_829);
xnor U5158 (N_5158,N_3191,N_1715);
and U5159 (N_5159,N_707,N_2473);
and U5160 (N_5160,N_270,N_3127);
and U5161 (N_5161,N_130,N_1418);
nand U5162 (N_5162,N_1229,N_54);
and U5163 (N_5163,N_335,N_1907);
nand U5164 (N_5164,N_1891,N_1606);
xnor U5165 (N_5165,N_1427,N_513);
and U5166 (N_5166,N_2010,N_587);
and U5167 (N_5167,N_3698,N_2276);
or U5168 (N_5168,N_3177,N_2396);
or U5169 (N_5169,N_3713,N_3119);
nand U5170 (N_5170,N_3513,N_536);
nand U5171 (N_5171,N_2322,N_3400);
or U5172 (N_5172,N_3689,N_3480);
or U5173 (N_5173,N_1838,N_772);
or U5174 (N_5174,N_2833,N_1009);
xor U5175 (N_5175,N_3040,N_759);
and U5176 (N_5176,N_408,N_3088);
and U5177 (N_5177,N_3744,N_3378);
nor U5178 (N_5178,N_2377,N_1511);
or U5179 (N_5179,N_3010,N_2742);
or U5180 (N_5180,N_125,N_754);
nand U5181 (N_5181,N_993,N_1034);
xnor U5182 (N_5182,N_1393,N_1827);
xor U5183 (N_5183,N_1438,N_1209);
nand U5184 (N_5184,N_10,N_1824);
nand U5185 (N_5185,N_1288,N_2138);
xor U5186 (N_5186,N_1352,N_2222);
nand U5187 (N_5187,N_3755,N_735);
nor U5188 (N_5188,N_650,N_283);
nor U5189 (N_5189,N_34,N_226);
xor U5190 (N_5190,N_3641,N_3668);
nand U5191 (N_5191,N_3614,N_2590);
or U5192 (N_5192,N_1519,N_2693);
xnor U5193 (N_5193,N_576,N_1227);
nand U5194 (N_5194,N_3533,N_3801);
xor U5195 (N_5195,N_2925,N_3071);
nor U5196 (N_5196,N_2641,N_3155);
xnor U5197 (N_5197,N_869,N_3079);
nor U5198 (N_5198,N_3907,N_2323);
xnor U5199 (N_5199,N_3707,N_2436);
nor U5200 (N_5200,N_654,N_3646);
nand U5201 (N_5201,N_3053,N_2838);
or U5202 (N_5202,N_3458,N_745);
xnor U5203 (N_5203,N_3914,N_1208);
xnor U5204 (N_5204,N_785,N_2528);
nor U5205 (N_5205,N_379,N_2189);
xnor U5206 (N_5206,N_3299,N_3740);
xnor U5207 (N_5207,N_2295,N_3783);
xnor U5208 (N_5208,N_2985,N_493);
and U5209 (N_5209,N_1859,N_3211);
nand U5210 (N_5210,N_2604,N_2999);
xor U5211 (N_5211,N_1103,N_2978);
xnor U5212 (N_5212,N_2289,N_312);
nand U5213 (N_5213,N_78,N_1316);
nor U5214 (N_5214,N_1993,N_1168);
nand U5215 (N_5215,N_93,N_1499);
and U5216 (N_5216,N_3082,N_2140);
nor U5217 (N_5217,N_2896,N_3540);
or U5218 (N_5218,N_2303,N_3989);
and U5219 (N_5219,N_3334,N_642);
and U5220 (N_5220,N_1657,N_2601);
nor U5221 (N_5221,N_1542,N_767);
nand U5222 (N_5222,N_3314,N_2674);
nor U5223 (N_5223,N_2599,N_3431);
xor U5224 (N_5224,N_100,N_2056);
or U5225 (N_5225,N_622,N_893);
or U5226 (N_5226,N_2766,N_1958);
xnor U5227 (N_5227,N_1474,N_2023);
and U5228 (N_5228,N_2807,N_2440);
xnor U5229 (N_5229,N_3007,N_3859);
nor U5230 (N_5230,N_3054,N_2905);
nand U5231 (N_5231,N_3162,N_1885);
and U5232 (N_5232,N_3284,N_676);
or U5233 (N_5233,N_2447,N_1586);
nand U5234 (N_5234,N_378,N_3677);
nand U5235 (N_5235,N_3457,N_1525);
nor U5236 (N_5236,N_727,N_1721);
or U5237 (N_5237,N_791,N_1231);
and U5238 (N_5238,N_3233,N_3562);
or U5239 (N_5239,N_2584,N_3566);
and U5240 (N_5240,N_2466,N_2666);
nand U5241 (N_5241,N_2821,N_1847);
or U5242 (N_5242,N_3418,N_1266);
and U5243 (N_5243,N_3469,N_2047);
xor U5244 (N_5244,N_85,N_3190);
and U5245 (N_5245,N_2962,N_3563);
nand U5246 (N_5246,N_1215,N_1428);
xor U5247 (N_5247,N_2511,N_685);
xnor U5248 (N_5248,N_3747,N_2594);
nand U5249 (N_5249,N_740,N_1833);
nor U5250 (N_5250,N_2015,N_617);
xnor U5251 (N_5251,N_3294,N_3921);
or U5252 (N_5252,N_2667,N_1928);
nor U5253 (N_5253,N_407,N_1473);
and U5254 (N_5254,N_1284,N_1604);
nor U5255 (N_5255,N_2663,N_2573);
or U5256 (N_5256,N_2809,N_3104);
nand U5257 (N_5257,N_2273,N_1797);
nand U5258 (N_5258,N_3246,N_3543);
or U5259 (N_5259,N_3670,N_552);
xor U5260 (N_5260,N_546,N_1989);
nor U5261 (N_5261,N_1782,N_877);
nand U5262 (N_5262,N_1207,N_2113);
nor U5263 (N_5263,N_526,N_2386);
or U5264 (N_5264,N_555,N_227);
and U5265 (N_5265,N_3549,N_2907);
xnor U5266 (N_5266,N_1780,N_405);
xnor U5267 (N_5267,N_1256,N_1982);
xor U5268 (N_5268,N_3798,N_240);
and U5269 (N_5269,N_2580,N_3242);
or U5270 (N_5270,N_3374,N_154);
or U5271 (N_5271,N_842,N_2517);
xnor U5272 (N_5272,N_1776,N_2824);
nor U5273 (N_5273,N_1592,N_3918);
xor U5274 (N_5274,N_3484,N_2953);
nor U5275 (N_5275,N_876,N_151);
and U5276 (N_5276,N_469,N_3339);
or U5277 (N_5277,N_1037,N_3335);
xor U5278 (N_5278,N_2525,N_2829);
or U5279 (N_5279,N_2759,N_69);
nor U5280 (N_5280,N_3643,N_2908);
nand U5281 (N_5281,N_1086,N_1236);
nor U5282 (N_5282,N_1927,N_3238);
nor U5283 (N_5283,N_2987,N_2659);
nor U5284 (N_5284,N_290,N_2118);
and U5285 (N_5285,N_875,N_2484);
and U5286 (N_5286,N_3943,N_357);
nand U5287 (N_5287,N_1123,N_1087);
or U5288 (N_5288,N_1936,N_2871);
or U5289 (N_5289,N_40,N_3249);
nand U5290 (N_5290,N_713,N_63);
nand U5291 (N_5291,N_3086,N_3830);
nor U5292 (N_5292,N_3764,N_3592);
or U5293 (N_5293,N_2855,N_157);
or U5294 (N_5294,N_1259,N_902);
nand U5295 (N_5295,N_3454,N_1046);
nor U5296 (N_5296,N_1402,N_910);
nor U5297 (N_5297,N_1822,N_3650);
or U5298 (N_5298,N_2728,N_1318);
or U5299 (N_5299,N_1603,N_2357);
and U5300 (N_5300,N_1312,N_205);
and U5301 (N_5301,N_3106,N_1808);
nand U5302 (N_5302,N_1587,N_1547);
or U5303 (N_5303,N_1120,N_2365);
nand U5304 (N_5304,N_1849,N_2523);
xnor U5305 (N_5305,N_2244,N_2639);
nand U5306 (N_5306,N_2370,N_1748);
and U5307 (N_5307,N_1778,N_1585);
xor U5308 (N_5308,N_2859,N_1961);
nor U5309 (N_5309,N_1517,N_2275);
nand U5310 (N_5310,N_3383,N_3343);
nand U5311 (N_5311,N_1996,N_2458);
or U5312 (N_5312,N_3442,N_1889);
nand U5313 (N_5313,N_3891,N_128);
nand U5314 (N_5314,N_3877,N_3200);
or U5315 (N_5315,N_3788,N_442);
nand U5316 (N_5316,N_1579,N_339);
and U5317 (N_5317,N_2455,N_1351);
or U5318 (N_5318,N_1716,N_1007);
xor U5319 (N_5319,N_1329,N_682);
nand U5320 (N_5320,N_2612,N_3230);
xnor U5321 (N_5321,N_3470,N_27);
xor U5322 (N_5322,N_2777,N_1655);
or U5323 (N_5323,N_1920,N_1368);
nor U5324 (N_5324,N_817,N_638);
nand U5325 (N_5325,N_441,N_982);
nor U5326 (N_5326,N_1154,N_1232);
or U5327 (N_5327,N_2544,N_978);
and U5328 (N_5328,N_1280,N_280);
and U5329 (N_5329,N_166,N_367);
xor U5330 (N_5330,N_3962,N_2478);
xnor U5331 (N_5331,N_2734,N_2307);
nor U5332 (N_5332,N_920,N_569);
nor U5333 (N_5333,N_485,N_2027);
nand U5334 (N_5334,N_231,N_963);
and U5335 (N_5335,N_3215,N_1320);
or U5336 (N_5336,N_214,N_1401);
nor U5337 (N_5337,N_572,N_2168);
xnor U5338 (N_5338,N_2403,N_3872);
or U5339 (N_5339,N_1763,N_155);
nand U5340 (N_5340,N_1148,N_313);
nand U5341 (N_5341,N_2164,N_1652);
nor U5342 (N_5342,N_600,N_3490);
nand U5343 (N_5343,N_1301,N_350);
nand U5344 (N_5344,N_2868,N_3865);
nor U5345 (N_5345,N_1869,N_3502);
nand U5346 (N_5346,N_2536,N_363);
or U5347 (N_5347,N_1271,N_2900);
nor U5348 (N_5348,N_30,N_2086);
nor U5349 (N_5349,N_3717,N_3277);
and U5350 (N_5350,N_1588,N_2678);
and U5351 (N_5351,N_2876,N_1455);
nor U5352 (N_5352,N_3752,N_2803);
or U5353 (N_5353,N_3603,N_2756);
xnor U5354 (N_5354,N_2280,N_1150);
and U5355 (N_5355,N_1730,N_1281);
and U5356 (N_5356,N_3652,N_3761);
nor U5357 (N_5357,N_1491,N_3120);
and U5358 (N_5358,N_658,N_186);
or U5359 (N_5359,N_1371,N_1126);
nor U5360 (N_5360,N_980,N_3350);
nor U5361 (N_5361,N_1020,N_2084);
nor U5362 (N_5362,N_809,N_2795);
xnor U5363 (N_5363,N_1443,N_2818);
or U5364 (N_5364,N_425,N_371);
nand U5365 (N_5365,N_3122,N_3756);
xnor U5366 (N_5366,N_702,N_3389);
nand U5367 (N_5367,N_2063,N_2785);
or U5368 (N_5368,N_3957,N_2298);
xnor U5369 (N_5369,N_529,N_3993);
nand U5370 (N_5370,N_2350,N_1692);
nand U5371 (N_5371,N_1040,N_1189);
or U5372 (N_5372,N_1166,N_3887);
xor U5373 (N_5373,N_1321,N_1676);
nand U5374 (N_5374,N_596,N_3261);
nand U5375 (N_5375,N_1675,N_475);
nor U5376 (N_5376,N_1549,N_1934);
nand U5377 (N_5377,N_2755,N_2234);
nand U5378 (N_5378,N_3315,N_1391);
nand U5379 (N_5379,N_2431,N_3647);
xor U5380 (N_5380,N_3255,N_807);
and U5381 (N_5381,N_2676,N_1990);
nand U5382 (N_5382,N_250,N_1723);
and U5383 (N_5383,N_1362,N_3364);
xnor U5384 (N_5384,N_1228,N_3055);
xor U5385 (N_5385,N_2989,N_3058);
xnor U5386 (N_5386,N_1751,N_1623);
or U5387 (N_5387,N_956,N_277);
xor U5388 (N_5388,N_82,N_1310);
and U5389 (N_5389,N_1331,N_3178);
nand U5390 (N_5390,N_2277,N_2754);
and U5391 (N_5391,N_2764,N_2032);
xor U5392 (N_5392,N_135,N_296);
nor U5393 (N_5393,N_948,N_3027);
nor U5394 (N_5394,N_1456,N_2960);
xnor U5395 (N_5395,N_700,N_3570);
nand U5396 (N_5396,N_264,N_3260);
nand U5397 (N_5397,N_315,N_924);
nor U5398 (N_5398,N_3936,N_2662);
or U5399 (N_5399,N_3448,N_92);
nand U5400 (N_5400,N_1373,N_1407);
or U5401 (N_5401,N_964,N_3170);
nor U5402 (N_5402,N_3754,N_1445);
nor U5403 (N_5403,N_3998,N_3615);
and U5404 (N_5404,N_3935,N_1632);
or U5405 (N_5405,N_827,N_1622);
nand U5406 (N_5406,N_2379,N_3919);
nor U5407 (N_5407,N_1255,N_537);
and U5408 (N_5408,N_2816,N_2723);
nand U5409 (N_5409,N_898,N_134);
xor U5410 (N_5410,N_1218,N_2284);
xnor U5411 (N_5411,N_1118,N_2493);
nand U5412 (N_5412,N_2694,N_145);
and U5413 (N_5413,N_3977,N_103);
and U5414 (N_5414,N_773,N_664);
nand U5415 (N_5415,N_2016,N_3536);
xor U5416 (N_5416,N_3336,N_3137);
nand U5417 (N_5417,N_1733,N_2018);
nor U5418 (N_5418,N_1397,N_2136);
nand U5419 (N_5419,N_1380,N_2311);
nand U5420 (N_5420,N_403,N_3271);
xor U5421 (N_5421,N_3728,N_306);
or U5422 (N_5422,N_129,N_3711);
and U5423 (N_5423,N_3799,N_2873);
and U5424 (N_5424,N_2452,N_1247);
nand U5425 (N_5425,N_2739,N_59);
xnor U5426 (N_5426,N_3169,N_1886);
or U5427 (N_5427,N_3247,N_2423);
nand U5428 (N_5428,N_462,N_1668);
nand U5429 (N_5429,N_891,N_1178);
or U5430 (N_5430,N_178,N_251);
nand U5431 (N_5431,N_2494,N_3696);
nand U5432 (N_5432,N_219,N_2378);
xnor U5433 (N_5433,N_1234,N_3370);
nor U5434 (N_5434,N_566,N_1638);
nand U5435 (N_5435,N_358,N_2524);
or U5436 (N_5436,N_1630,N_3574);
or U5437 (N_5437,N_3544,N_1750);
nand U5438 (N_5438,N_3987,N_108);
and U5439 (N_5439,N_3160,N_3219);
or U5440 (N_5440,N_402,N_1333);
nor U5441 (N_5441,N_2230,N_2932);
nand U5442 (N_5442,N_1490,N_3465);
nand U5443 (N_5443,N_1353,N_764);
xnor U5444 (N_5444,N_1263,N_1520);
xnor U5445 (N_5445,N_3932,N_2111);
xnor U5446 (N_5446,N_1755,N_1332);
or U5447 (N_5447,N_297,N_3037);
nand U5448 (N_5448,N_1793,N_2530);
and U5449 (N_5449,N_2260,N_2929);
xnor U5450 (N_5450,N_116,N_3477);
and U5451 (N_5451,N_2448,N_3913);
xor U5452 (N_5452,N_3905,N_3767);
xor U5453 (N_5453,N_1613,N_1069);
xnor U5454 (N_5454,N_761,N_2424);
nor U5455 (N_5455,N_43,N_790);
xnor U5456 (N_5456,N_349,N_3340);
nor U5457 (N_5457,N_449,N_1756);
and U5458 (N_5458,N_3506,N_2421);
nor U5459 (N_5459,N_1823,N_1369);
nand U5460 (N_5460,N_1976,N_2310);
nor U5461 (N_5461,N_404,N_1302);
xnor U5462 (N_5462,N_1667,N_3278);
or U5463 (N_5463,N_1661,N_474);
nor U5464 (N_5464,N_1167,N_2743);
nand U5465 (N_5465,N_348,N_3748);
xor U5466 (N_5466,N_3842,N_2931);
and U5467 (N_5467,N_2951,N_1683);
nor U5468 (N_5468,N_2834,N_1862);
nand U5469 (N_5469,N_711,N_3301);
xor U5470 (N_5470,N_3535,N_3276);
xor U5471 (N_5471,N_2687,N_2184);
xnor U5472 (N_5472,N_1089,N_2920);
or U5473 (N_5473,N_2070,N_2306);
or U5474 (N_5474,N_3115,N_2241);
xor U5475 (N_5475,N_440,N_3172);
nor U5476 (N_5476,N_1508,N_3098);
nand U5477 (N_5477,N_961,N_776);
xor U5478 (N_5478,N_3142,N_1980);
nor U5479 (N_5479,N_2314,N_3432);
and U5480 (N_5480,N_2391,N_3375);
nor U5481 (N_5481,N_2851,N_189);
xor U5482 (N_5482,N_3410,N_2141);
xnor U5483 (N_5483,N_2321,N_523);
nor U5484 (N_5484,N_2054,N_3180);
or U5485 (N_5485,N_3150,N_3782);
nand U5486 (N_5486,N_2499,N_3181);
nand U5487 (N_5487,N_857,N_1017);
and U5488 (N_5488,N_1199,N_3377);
xor U5489 (N_5489,N_2354,N_2521);
nor U5490 (N_5490,N_3346,N_3902);
or U5491 (N_5491,N_3047,N_2598);
nand U5492 (N_5492,N_2109,N_533);
nor U5493 (N_5493,N_766,N_249);
nand U5494 (N_5494,N_3274,N_2961);
xor U5495 (N_5495,N_2467,N_2781);
nand U5496 (N_5496,N_974,N_2751);
xnor U5497 (N_5497,N_852,N_708);
nor U5498 (N_5498,N_1177,N_2165);
or U5499 (N_5499,N_1081,N_1221);
xor U5500 (N_5500,N_1071,N_2020);
xnor U5501 (N_5501,N_786,N_4);
and U5502 (N_5502,N_714,N_1831);
nand U5503 (N_5503,N_1513,N_292);
nor U5504 (N_5504,N_2235,N_2837);
nand U5505 (N_5505,N_3390,N_2123);
nor U5506 (N_5506,N_3635,N_3520);
or U5507 (N_5507,N_3325,N_480);
and U5508 (N_5508,N_2096,N_804);
and U5509 (N_5509,N_284,N_1850);
nor U5510 (N_5510,N_3923,N_2203);
nand U5511 (N_5511,N_1272,N_1974);
nand U5512 (N_5512,N_1113,N_2591);
nand U5513 (N_5513,N_2516,N_2847);
xnor U5514 (N_5514,N_3196,N_1014);
xnor U5515 (N_5515,N_1196,N_433);
nand U5516 (N_5516,N_1999,N_1546);
xnor U5517 (N_5517,N_991,N_1514);
nand U5518 (N_5518,N_2160,N_511);
and U5519 (N_5519,N_3493,N_384);
or U5520 (N_5520,N_2545,N_1444);
or U5521 (N_5521,N_2863,N_463);
or U5522 (N_5522,N_419,N_698);
nand U5523 (N_5523,N_904,N_1754);
nor U5524 (N_5524,N_3663,N_3397);
nor U5525 (N_5525,N_1433,N_841);
nand U5526 (N_5526,N_2215,N_479);
or U5527 (N_5527,N_162,N_3153);
or U5528 (N_5528,N_3745,N_1294);
xor U5529 (N_5529,N_362,N_2914);
xor U5530 (N_5530,N_3537,N_1251);
or U5531 (N_5531,N_1297,N_1669);
or U5532 (N_5532,N_3996,N_3253);
nor U5533 (N_5533,N_3372,N_1734);
nand U5534 (N_5534,N_67,N_1295);
and U5535 (N_5535,N_609,N_3555);
or U5536 (N_5536,N_2508,N_168);
or U5537 (N_5537,N_390,N_2353);
xnor U5538 (N_5538,N_347,N_2532);
or U5539 (N_5539,N_1119,N_1042);
or U5540 (N_5540,N_1142,N_3056);
xnor U5541 (N_5541,N_2571,N_1766);
nor U5542 (N_5542,N_211,N_3290);
nor U5543 (N_5543,N_3700,N_2812);
nand U5544 (N_5544,N_3941,N_899);
xnor U5545 (N_5545,N_3559,N_1798);
xor U5546 (N_5546,N_1277,N_3268);
nand U5547 (N_5547,N_1233,N_2626);
nand U5548 (N_5548,N_2860,N_1904);
nand U5549 (N_5549,N_3999,N_1324);
nand U5550 (N_5550,N_3558,N_3412);
or U5551 (N_5551,N_2102,N_2646);
nand U5552 (N_5552,N_414,N_2359);
nor U5553 (N_5553,N_1080,N_57);
or U5554 (N_5554,N_2836,N_318);
xor U5555 (N_5555,N_2347,N_723);
nand U5556 (N_5556,N_3320,N_3381);
xor U5557 (N_5557,N_901,N_1526);
and U5558 (N_5558,N_1650,N_2217);
nand U5559 (N_5559,N_1599,N_952);
or U5560 (N_5560,N_3264,N_2430);
or U5561 (N_5561,N_2910,N_2290);
xor U5562 (N_5562,N_571,N_396);
or U5563 (N_5563,N_2419,N_3858);
or U5564 (N_5564,N_818,N_221);
or U5565 (N_5565,N_874,N_2515);
or U5566 (N_5566,N_3854,N_2887);
nand U5567 (N_5567,N_2762,N_3532);
or U5568 (N_5568,N_261,N_2991);
and U5569 (N_5569,N_1296,N_2984);
xor U5570 (N_5570,N_2226,N_1061);
or U5571 (N_5571,N_2446,N_726);
xor U5572 (N_5572,N_3305,N_99);
xnor U5573 (N_5573,N_258,N_1627);
nor U5574 (N_5574,N_1348,N_3345);
nor U5575 (N_5575,N_1709,N_1201);
nand U5576 (N_5576,N_218,N_2130);
xnor U5577 (N_5577,N_932,N_2464);
and U5578 (N_5578,N_175,N_2939);
nand U5579 (N_5579,N_121,N_2990);
nand U5580 (N_5580,N_1696,N_830);
and U5581 (N_5581,N_1789,N_3131);
xnor U5582 (N_5582,N_450,N_2019);
nand U5583 (N_5583,N_1346,N_2268);
nand U5584 (N_5584,N_2605,N_1784);
nor U5585 (N_5585,N_3900,N_238);
nand U5586 (N_5586,N_943,N_3595);
and U5587 (N_5587,N_1994,N_2560);
and U5588 (N_5588,N_2780,N_1403);
nand U5589 (N_5589,N_931,N_1690);
or U5590 (N_5590,N_1421,N_193);
nor U5591 (N_5591,N_3526,N_3529);
or U5592 (N_5592,N_235,N_543);
nor U5593 (N_5593,N_3141,N_141);
or U5594 (N_5594,N_1641,N_1626);
and U5595 (N_5595,N_3248,N_1752);
and U5596 (N_5596,N_506,N_3497);
xnor U5597 (N_5597,N_336,N_3664);
xor U5598 (N_5598,N_514,N_3130);
or U5599 (N_5599,N_747,N_3712);
or U5600 (N_5600,N_2444,N_1115);
nor U5601 (N_5601,N_1205,N_2037);
or U5602 (N_5602,N_174,N_3853);
nor U5603 (N_5603,N_3224,N_2881);
nor U5604 (N_5604,N_2406,N_2582);
nand U5605 (N_5605,N_959,N_1809);
or U5606 (N_5606,N_1413,N_578);
nand U5607 (N_5607,N_553,N_1770);
nor U5608 (N_5608,N_2709,N_2336);
nand U5609 (N_5609,N_2616,N_1724);
and U5610 (N_5610,N_338,N_687);
xnor U5611 (N_5611,N_907,N_2239);
xor U5612 (N_5612,N_2771,N_3585);
and U5613 (N_5613,N_1472,N_453);
xor U5614 (N_5614,N_50,N_262);
or U5615 (N_5615,N_583,N_2757);
xor U5616 (N_5616,N_2262,N_401);
or U5617 (N_5617,N_3606,N_3110);
nand U5618 (N_5618,N_320,N_1489);
xor U5619 (N_5619,N_3310,N_2004);
and U5620 (N_5620,N_3704,N_2134);
or U5621 (N_5621,N_2535,N_3183);
nand U5622 (N_5622,N_2000,N_814);
xor U5623 (N_5623,N_1282,N_1360);
or U5624 (N_5624,N_1967,N_3780);
and U5625 (N_5625,N_3376,N_1569);
xnor U5626 (N_5626,N_3814,N_3920);
and U5627 (N_5627,N_3292,N_573);
nand U5628 (N_5628,N_307,N_232);
and U5629 (N_5629,N_3693,N_7);
or U5630 (N_5630,N_3093,N_3420);
or U5631 (N_5631,N_3797,N_3924);
and U5632 (N_5632,N_3685,N_3159);
nand U5633 (N_5633,N_1306,N_3686);
or U5634 (N_5634,N_539,N_3903);
or U5635 (N_5635,N_1206,N_2769);
nor U5636 (N_5636,N_2972,N_3175);
or U5637 (N_5637,N_1463,N_645);
xor U5638 (N_5638,N_1496,N_1292);
nor U5639 (N_5639,N_2258,N_730);
or U5640 (N_5640,N_2472,N_2451);
and U5641 (N_5641,N_3561,N_3955);
nor U5642 (N_5642,N_3407,N_3710);
nand U5643 (N_5643,N_806,N_538);
or U5644 (N_5644,N_2204,N_750);
nand U5645 (N_5645,N_1671,N_1486);
or U5646 (N_5646,N_3039,N_1289);
xor U5647 (N_5647,N_1132,N_3888);
nor U5648 (N_5648,N_331,N_716);
and U5649 (N_5649,N_2570,N_2305);
or U5650 (N_5650,N_3195,N_1649);
and U5651 (N_5651,N_314,N_3856);
xor U5652 (N_5652,N_1968,N_1946);
nor U5653 (N_5653,N_3426,N_156);
nor U5654 (N_5654,N_544,N_1877);
xor U5655 (N_5655,N_3975,N_3358);
xnor U5656 (N_5656,N_3964,N_1883);
nand U5657 (N_5657,N_870,N_1431);
nor U5658 (N_5658,N_3051,N_1153);
nor U5659 (N_5659,N_26,N_3642);
xor U5660 (N_5660,N_605,N_1504);
nor U5661 (N_5661,N_3557,N_2199);
nand U5662 (N_5662,N_3787,N_3029);
xnor U5663 (N_5663,N_1500,N_3092);
or U5664 (N_5664,N_198,N_2116);
and U5665 (N_5665,N_1777,N_2553);
nor U5666 (N_5666,N_2748,N_1275);
nor U5667 (N_5667,N_1914,N_3463);
or U5668 (N_5668,N_815,N_2326);
xor U5669 (N_5669,N_2376,N_955);
xnor U5670 (N_5670,N_3124,N_6);
nand U5671 (N_5671,N_353,N_3022);
xor U5672 (N_5672,N_2677,N_757);
and U5673 (N_5673,N_3064,N_1319);
or U5674 (N_5674,N_281,N_2119);
nand U5675 (N_5675,N_1349,N_1308);
nor U5676 (N_5676,N_2014,N_1030);
and U5677 (N_5677,N_428,N_1156);
and U5678 (N_5678,N_330,N_2293);
xnor U5679 (N_5679,N_2195,N_3868);
and U5680 (N_5680,N_3380,N_1423);
or U5681 (N_5681,N_2643,N_3348);
nand U5682 (N_5682,N_366,N_3425);
nor U5683 (N_5683,N_3658,N_887);
nor U5684 (N_5684,N_3478,N_1576);
or U5685 (N_5685,N_1001,N_3483);
nand U5686 (N_5686,N_1767,N_340);
nand U5687 (N_5687,N_3521,N_2097);
and U5688 (N_5688,N_1684,N_2698);
xor U5689 (N_5689,N_2107,N_2214);
nor U5690 (N_5690,N_3024,N_1378);
and U5691 (N_5691,N_1686,N_21);
and U5692 (N_5692,N_1518,N_686);
nand U5693 (N_5693,N_1918,N_203);
xor U5694 (N_5694,N_915,N_3699);
nor U5695 (N_5695,N_704,N_3223);
nand U5696 (N_5696,N_58,N_548);
xor U5697 (N_5697,N_2143,N_2805);
or U5698 (N_5698,N_1457,N_2519);
nand U5699 (N_5699,N_1532,N_725);
xor U5700 (N_5700,N_423,N_2067);
nand U5701 (N_5701,N_3321,N_411);
or U5702 (N_5702,N_1045,N_957);
nand U5703 (N_5703,N_1260,N_3282);
or U5704 (N_5704,N_2414,N_3275);
nor U5705 (N_5705,N_2005,N_1244);
nor U5706 (N_5706,N_3607,N_2031);
nand U5707 (N_5707,N_554,N_2526);
nor U5708 (N_5708,N_197,N_1025);
nor U5709 (N_5709,N_1662,N_2947);
or U5710 (N_5710,N_3857,N_1732);
or U5711 (N_5711,N_2139,N_556);
nor U5712 (N_5712,N_2301,N_2736);
nand U5713 (N_5713,N_542,N_3757);
xnor U5714 (N_5714,N_1137,N_260);
xnor U5715 (N_5715,N_345,N_2842);
or U5716 (N_5716,N_528,N_2970);
nor U5717 (N_5717,N_212,N_981);
nand U5718 (N_5718,N_1618,N_1541);
or U5719 (N_5719,N_947,N_3528);
nor U5720 (N_5720,N_744,N_1819);
and U5721 (N_5721,N_3867,N_2137);
nor U5722 (N_5722,N_1731,N_2149);
xnor U5723 (N_5723,N_1697,N_2050);
nor U5724 (N_5724,N_3045,N_1567);
nand U5725 (N_5725,N_2167,N_1110);
xor U5726 (N_5726,N_2439,N_3886);
xor U5727 (N_5727,N_2427,N_1682);
nand U5728 (N_5728,N_254,N_2380);
and U5729 (N_5729,N_2433,N_2941);
xnor U5730 (N_5730,N_369,N_3262);
xor U5731 (N_5731,N_3067,N_2529);
nand U5732 (N_5732,N_324,N_3836);
nand U5733 (N_5733,N_2554,N_1568);
or U5734 (N_5734,N_1645,N_3988);
nor U5735 (N_5735,N_1063,N_208);
xor U5736 (N_5736,N_3848,N_3899);
nor U5737 (N_5737,N_2711,N_3632);
and U5738 (N_5738,N_1285,N_580);
nand U5739 (N_5739,N_1488,N_3727);
xnor U5740 (N_5740,N_781,N_446);
xnor U5741 (N_5741,N_1303,N_3820);
and U5742 (N_5742,N_850,N_1015);
nor U5743 (N_5743,N_3687,N_1956);
and U5744 (N_5744,N_1493,N_3351);
nand U5745 (N_5745,N_2672,N_394);
xnor U5746 (N_5746,N_743,N_2154);
and U5747 (N_5747,N_661,N_1483);
nor U5748 (N_5748,N_3937,N_3605);
xnor U5749 (N_5749,N_2870,N_1449);
nand U5750 (N_5750,N_3203,N_3020);
nand U5751 (N_5751,N_732,N_106);
and U5752 (N_5752,N_3157,N_833);
nand U5753 (N_5753,N_282,N_1197);
and U5754 (N_5754,N_3218,N_1060);
and U5755 (N_5755,N_2964,N_896);
xnor U5756 (N_5756,N_2974,N_1708);
xnor U5757 (N_5757,N_2078,N_2065);
nand U5758 (N_5758,N_3541,N_2457);
nor U5759 (N_5759,N_329,N_2514);
and U5760 (N_5760,N_360,N_1959);
xnor U5761 (N_5761,N_2271,N_1469);
xor U5762 (N_5762,N_2351,N_2490);
xor U5763 (N_5763,N_3800,N_3075);
xnor U5764 (N_5764,N_1313,N_3845);
or U5765 (N_5765,N_188,N_987);
xor U5766 (N_5766,N_487,N_3792);
nand U5767 (N_5767,N_3576,N_1085);
xnor U5768 (N_5768,N_1048,N_3827);
xnor U5769 (N_5769,N_892,N_204);
or U5770 (N_5770,N_675,N_3925);
or U5771 (N_5771,N_117,N_1342);
and U5772 (N_5772,N_3163,N_1615);
and U5773 (N_5773,N_2622,N_1867);
and U5774 (N_5774,N_3835,N_979);
and U5775 (N_5775,N_2533,N_3384);
xnor U5776 (N_5776,N_3298,N_2949);
nand U5777 (N_5777,N_2142,N_2552);
and U5778 (N_5778,N_461,N_1170);
and U5779 (N_5779,N_3824,N_1091);
or U5780 (N_5780,N_2060,N_1395);
and U5781 (N_5781,N_2506,N_420);
or U5782 (N_5782,N_928,N_1454);
nor U5783 (N_5783,N_3694,N_2668);
nand U5784 (N_5784,N_2811,N_1230);
and U5785 (N_5785,N_2715,N_2428);
xnor U5786 (N_5786,N_2294,N_840);
and U5787 (N_5787,N_2312,N_298);
nand U5788 (N_5788,N_1051,N_3708);
nand U5789 (N_5789,N_3621,N_1545);
nand U5790 (N_5790,N_127,N_1580);
xor U5791 (N_5791,N_3762,N_2132);
nand U5792 (N_5792,N_3967,N_269);
nand U5793 (N_5793,N_207,N_274);
or U5794 (N_5794,N_3042,N_478);
xnor U5795 (N_5795,N_1954,N_1035);
nor U5796 (N_5796,N_844,N_1257);
xnor U5797 (N_5797,N_3672,N_180);
nand U5798 (N_5798,N_1043,N_1248);
nand U5799 (N_5799,N_864,N_3774);
xnor U5800 (N_5800,N_2603,N_1096);
and U5801 (N_5801,N_2802,N_426);
xnor U5802 (N_5802,N_1304,N_2238);
xnor U5803 (N_5803,N_1268,N_2272);
nand U5804 (N_5804,N_1184,N_2095);
nor U5805 (N_5805,N_3933,N_1152);
nand U5806 (N_5806,N_996,N_376);
or U5807 (N_5807,N_146,N_755);
or U5808 (N_5808,N_2090,N_2936);
nand U5809 (N_5809,N_2656,N_3363);
nand U5810 (N_5810,N_2607,N_2720);
and U5811 (N_5811,N_2564,N_1131);
or U5812 (N_5812,N_3422,N_1141);
nand U5813 (N_5813,N_2718,N_2684);
or U5814 (N_5814,N_2513,N_2606);
nor U5815 (N_5815,N_3733,N_72);
nor U5816 (N_5816,N_3703,N_597);
xor U5817 (N_5817,N_3572,N_3850);
or U5818 (N_5818,N_648,N_1972);
and U5819 (N_5819,N_1521,N_2823);
or U5820 (N_5820,N_2062,N_1066);
and U5821 (N_5821,N_796,N_2758);
and U5822 (N_5822,N_1768,N_492);
and U5823 (N_5823,N_2125,N_1162);
and U5824 (N_5824,N_2003,N_1365);
or U5825 (N_5825,N_1018,N_1022);
nor U5826 (N_5826,N_3306,N_265);
or U5827 (N_5827,N_2854,N_2039);
nand U5828 (N_5828,N_3847,N_1860);
nand U5829 (N_5829,N_1262,N_1617);
xnor U5830 (N_5830,N_501,N_2577);
and U5831 (N_5831,N_1593,N_2361);
nand U5832 (N_5832,N_244,N_17);
or U5833 (N_5833,N_2126,N_2669);
nand U5834 (N_5834,N_3154,N_2700);
nand U5835 (N_5835,N_3610,N_3225);
nor U5836 (N_5836,N_559,N_2944);
xor U5837 (N_5837,N_507,N_1983);
or U5838 (N_5838,N_2017,N_3873);
nor U5839 (N_5839,N_1963,N_705);
or U5840 (N_5840,N_803,N_1055);
nand U5841 (N_5841,N_3078,N_132);
nor U5842 (N_5842,N_2846,N_3116);
nand U5843 (N_5843,N_2673,N_1450);
nor U5844 (N_5844,N_2937,N_434);
or U5845 (N_5845,N_2632,N_816);
nand U5846 (N_5846,N_1340,N_356);
and U5847 (N_5847,N_2008,N_1817);
and U5848 (N_5848,N_847,N_39);
nand U5849 (N_5849,N_2786,N_2327);
and U5850 (N_5850,N_2495,N_305);
nor U5851 (N_5851,N_1477,N_1143);
nand U5852 (N_5852,N_1138,N_2744);
nor U5853 (N_5853,N_3512,N_1439);
and U5854 (N_5854,N_1317,N_2400);
xor U5855 (N_5855,N_3736,N_74);
and U5856 (N_5856,N_625,N_1987);
nor U5857 (N_5857,N_3102,N_655);
and U5858 (N_5858,N_3355,N_3091);
xnor U5859 (N_5859,N_2745,N_1217);
nor U5860 (N_5860,N_3961,N_288);
or U5861 (N_5861,N_3889,N_1729);
xor U5862 (N_5862,N_2889,N_1801);
or U5863 (N_5863,N_2952,N_903);
nand U5864 (N_5864,N_3522,N_37);
and U5865 (N_5865,N_611,N_2445);
and U5866 (N_5866,N_2977,N_370);
xnor U5867 (N_5867,N_2269,N_1608);
nor U5868 (N_5868,N_835,N_1193);
and U5869 (N_5869,N_3684,N_393);
nor U5870 (N_5870,N_2442,N_3586);
or U5871 (N_5871,N_3874,N_1430);
or U5872 (N_5872,N_342,N_1364);
nand U5873 (N_5873,N_1893,N_3878);
xnor U5874 (N_5874,N_3368,N_3);
nor U5875 (N_5875,N_2401,N_2252);
or U5876 (N_5876,N_2461,N_2614);
nor U5877 (N_5877,N_3111,N_3775);
nand U5878 (N_5878,N_3518,N_2796);
nor U5879 (N_5879,N_1254,N_3897);
xor U5880 (N_5880,N_2651,N_418);
xor U5881 (N_5881,N_3072,N_2927);
and U5882 (N_5882,N_929,N_3399);
nand U5883 (N_5883,N_1052,N_3099);
nand U5884 (N_5884,N_3446,N_584);
or U5885 (N_5885,N_1461,N_3237);
nor U5886 (N_5886,N_3638,N_2539);
or U5887 (N_5887,N_185,N_3329);
or U5888 (N_5888,N_124,N_3860);
nand U5889 (N_5889,N_939,N_1772);
or U5890 (N_5890,N_3619,N_594);
nor U5891 (N_5891,N_1629,N_1858);
nand U5892 (N_5892,N_1554,N_2685);
and U5893 (N_5893,N_3415,N_3501);
and U5894 (N_5894,N_1536,N_2059);
nor U5895 (N_5895,N_2877,N_3654);
xnor U5896 (N_5896,N_1591,N_1325);
nor U5897 (N_5897,N_2381,N_525);
nor U5898 (N_5898,N_3387,N_1501);
nand U5899 (N_5899,N_1783,N_620);
and U5900 (N_5900,N_1347,N_35);
xnor U5901 (N_5901,N_2483,N_3419);
nand U5902 (N_5902,N_2982,N_1908);
nor U5903 (N_5903,N_3602,N_1736);
or U5904 (N_5904,N_385,N_1314);
and U5905 (N_5905,N_3066,N_2981);
nand U5906 (N_5906,N_1105,N_2099);
and U5907 (N_5907,N_2950,N_12);
nor U5908 (N_5908,N_3174,N_3828);
nand U5909 (N_5909,N_3052,N_2363);
and U5910 (N_5910,N_2385,N_1688);
nor U5911 (N_5911,N_2815,N_1658);
or U5912 (N_5912,N_3144,N_880);
nor U5913 (N_5913,N_762,N_2475);
and U5914 (N_5914,N_1973,N_795);
xnor U5915 (N_5915,N_1844,N_1124);
or U5916 (N_5916,N_1912,N_3133);
nand U5917 (N_5917,N_3898,N_1175);
or U5918 (N_5918,N_678,N_3208);
nor U5919 (N_5919,N_652,N_2830);
nand U5920 (N_5920,N_608,N_2899);
and U5921 (N_5921,N_183,N_2368);
and U5922 (N_5922,N_3270,N_2878);
and U5923 (N_5923,N_1130,N_343);
or U5924 (N_5924,N_1385,N_3816);
or U5925 (N_5925,N_224,N_181);
nand U5926 (N_5926,N_3674,N_1938);
nand U5927 (N_5927,N_1932,N_524);
or U5928 (N_5928,N_1803,N_53);
nand U5929 (N_5929,N_649,N_1211);
or U5930 (N_5930,N_839,N_1102);
xor U5931 (N_5931,N_2274,N_3189);
nor U5932 (N_5932,N_793,N_838);
or U5933 (N_5933,N_177,N_2013);
nor U5934 (N_5934,N_3523,N_1548);
and U5935 (N_5935,N_1759,N_3267);
xnor U5936 (N_5936,N_568,N_3353);
and U5937 (N_5937,N_3061,N_949);
nor U5938 (N_5938,N_3447,N_1396);
nor U5939 (N_5939,N_3496,N_1505);
or U5940 (N_5940,N_3143,N_451);
or U5941 (N_5941,N_2253,N_3050);
nand U5942 (N_5942,N_94,N_2308);
xor U5943 (N_5943,N_24,N_3623);
nand U5944 (N_5944,N_3185,N_1434);
nand U5945 (N_5945,N_3089,N_3862);
or U5946 (N_5946,N_3475,N_780);
nand U5947 (N_5947,N_3328,N_3645);
nand U5948 (N_5948,N_1112,N_779);
nor U5949 (N_5949,N_3904,N_2568);
nand U5950 (N_5950,N_2538,N_417);
xnor U5951 (N_5951,N_3759,N_2061);
xor U5952 (N_5952,N_2171,N_346);
xor U5953 (N_5953,N_484,N_3018);
or U5954 (N_5954,N_2463,N_2609);
and U5955 (N_5955,N_1338,N_1065);
nor U5956 (N_5956,N_591,N_3839);
or U5957 (N_5957,N_1515,N_1853);
and U5958 (N_5958,N_3869,N_1829);
nor U5959 (N_5959,N_1854,N_774);
or U5960 (N_5960,N_653,N_3590);
nor U5961 (N_5961,N_334,N_3487);
nor U5962 (N_5962,N_2197,N_2586);
nand U5963 (N_5963,N_3156,N_3360);
nand U5964 (N_5964,N_1722,N_3986);
xnor U5965 (N_5965,N_18,N_2861);
or U5966 (N_5966,N_3227,N_1947);
or U5967 (N_5967,N_2242,N_1334);
or U5968 (N_5968,N_756,N_29);
and U5969 (N_5969,N_84,N_3359);
nor U5970 (N_5970,N_2420,N_2776);
xor U5971 (N_5971,N_1799,N_1079);
or U5972 (N_5972,N_3773,N_3593);
nor U5973 (N_5973,N_2340,N_1460);
or U5974 (N_5974,N_2968,N_1462);
nor U5975 (N_5975,N_3019,N_2148);
nor U5976 (N_5976,N_3637,N_2822);
and U5977 (N_5977,N_3489,N_668);
xnor U5978 (N_5978,N_2263,N_228);
xnor U5979 (N_5979,N_1252,N_409);
or U5980 (N_5980,N_1399,N_1157);
or U5981 (N_5981,N_3849,N_1666);
xnor U5982 (N_5982,N_2150,N_908);
and U5983 (N_5983,N_3922,N_962);
or U5984 (N_5984,N_3959,N_2425);
nand U5985 (N_5985,N_220,N_456);
and U5986 (N_5986,N_172,N_355);
and U5987 (N_5987,N_3285,N_2888);
and U5988 (N_5988,N_3653,N_3973);
xor U5989 (N_5989,N_498,N_486);
nand U5990 (N_5990,N_1179,N_1210);
or U5991 (N_5991,N_1602,N_2886);
xnor U5992 (N_5992,N_1226,N_1136);
or U5993 (N_5993,N_2806,N_897);
and U5994 (N_5994,N_3440,N_926);
and U5995 (N_5995,N_2527,N_2145);
nand U5996 (N_5996,N_1747,N_1174);
nand U5997 (N_5997,N_748,N_2680);
and U5998 (N_5998,N_1892,N_1186);
or U5999 (N_5999,N_2404,N_3245);
nand U6000 (N_6000,N_1683,N_685);
nand U6001 (N_6001,N_3989,N_68);
xor U6002 (N_6002,N_2269,N_184);
xor U6003 (N_6003,N_1573,N_2201);
xor U6004 (N_6004,N_1356,N_1248);
and U6005 (N_6005,N_2847,N_1494);
nand U6006 (N_6006,N_2969,N_1350);
nand U6007 (N_6007,N_53,N_474);
nor U6008 (N_6008,N_3023,N_787);
xor U6009 (N_6009,N_208,N_800);
nand U6010 (N_6010,N_1063,N_2785);
or U6011 (N_6011,N_1287,N_2611);
and U6012 (N_6012,N_1334,N_475);
xor U6013 (N_6013,N_1352,N_2342);
or U6014 (N_6014,N_2161,N_209);
and U6015 (N_6015,N_1231,N_1744);
nor U6016 (N_6016,N_2345,N_754);
and U6017 (N_6017,N_3727,N_1079);
and U6018 (N_6018,N_2294,N_3293);
and U6019 (N_6019,N_1429,N_1721);
nor U6020 (N_6020,N_22,N_3129);
and U6021 (N_6021,N_2314,N_3644);
nand U6022 (N_6022,N_2981,N_1987);
or U6023 (N_6023,N_2870,N_1058);
nand U6024 (N_6024,N_731,N_2814);
nand U6025 (N_6025,N_1015,N_299);
nand U6026 (N_6026,N_3435,N_204);
xnor U6027 (N_6027,N_1123,N_680);
or U6028 (N_6028,N_2978,N_1525);
xor U6029 (N_6029,N_508,N_2035);
nor U6030 (N_6030,N_1261,N_708);
nand U6031 (N_6031,N_2180,N_898);
xor U6032 (N_6032,N_1221,N_310);
nand U6033 (N_6033,N_1154,N_7);
nor U6034 (N_6034,N_1703,N_743);
nor U6035 (N_6035,N_11,N_962);
or U6036 (N_6036,N_1418,N_3025);
nand U6037 (N_6037,N_2047,N_396);
xnor U6038 (N_6038,N_2200,N_681);
or U6039 (N_6039,N_3236,N_674);
nand U6040 (N_6040,N_3875,N_3014);
nor U6041 (N_6041,N_3043,N_1762);
nand U6042 (N_6042,N_79,N_1167);
xor U6043 (N_6043,N_3047,N_2834);
or U6044 (N_6044,N_340,N_2819);
nor U6045 (N_6045,N_1499,N_1885);
nand U6046 (N_6046,N_354,N_708);
nor U6047 (N_6047,N_26,N_67);
xor U6048 (N_6048,N_2559,N_1662);
xnor U6049 (N_6049,N_716,N_1275);
nor U6050 (N_6050,N_2352,N_1668);
xnor U6051 (N_6051,N_1858,N_2724);
nor U6052 (N_6052,N_562,N_851);
nand U6053 (N_6053,N_3615,N_2652);
or U6054 (N_6054,N_3334,N_1435);
nand U6055 (N_6055,N_1440,N_3623);
nor U6056 (N_6056,N_3699,N_735);
nand U6057 (N_6057,N_2269,N_220);
and U6058 (N_6058,N_1998,N_1281);
xnor U6059 (N_6059,N_153,N_796);
and U6060 (N_6060,N_2,N_2052);
and U6061 (N_6061,N_861,N_2025);
nand U6062 (N_6062,N_3957,N_518);
xor U6063 (N_6063,N_829,N_2714);
nand U6064 (N_6064,N_2159,N_2529);
nor U6065 (N_6065,N_714,N_1620);
or U6066 (N_6066,N_2320,N_290);
xnor U6067 (N_6067,N_1208,N_3847);
nor U6068 (N_6068,N_2992,N_2681);
nor U6069 (N_6069,N_131,N_3194);
xnor U6070 (N_6070,N_3158,N_2988);
or U6071 (N_6071,N_2084,N_2424);
and U6072 (N_6072,N_2548,N_1828);
nand U6073 (N_6073,N_3783,N_1076);
xor U6074 (N_6074,N_2454,N_3249);
nor U6075 (N_6075,N_1331,N_1875);
and U6076 (N_6076,N_127,N_1181);
and U6077 (N_6077,N_2518,N_670);
xor U6078 (N_6078,N_3988,N_3526);
xnor U6079 (N_6079,N_1778,N_3798);
nand U6080 (N_6080,N_1439,N_1900);
or U6081 (N_6081,N_3425,N_1626);
nor U6082 (N_6082,N_629,N_2005);
nand U6083 (N_6083,N_975,N_1308);
and U6084 (N_6084,N_1052,N_3334);
nand U6085 (N_6085,N_2320,N_162);
nand U6086 (N_6086,N_2308,N_1102);
or U6087 (N_6087,N_1160,N_3414);
nor U6088 (N_6088,N_914,N_3854);
xor U6089 (N_6089,N_3136,N_2756);
and U6090 (N_6090,N_3215,N_1701);
or U6091 (N_6091,N_3743,N_2276);
and U6092 (N_6092,N_674,N_3554);
xnor U6093 (N_6093,N_975,N_2939);
xnor U6094 (N_6094,N_708,N_1506);
xnor U6095 (N_6095,N_3857,N_2178);
xnor U6096 (N_6096,N_2429,N_3680);
or U6097 (N_6097,N_3383,N_338);
nand U6098 (N_6098,N_2067,N_3801);
and U6099 (N_6099,N_1275,N_1769);
and U6100 (N_6100,N_2792,N_1770);
nor U6101 (N_6101,N_2515,N_2987);
or U6102 (N_6102,N_2397,N_2441);
or U6103 (N_6103,N_2143,N_2526);
nand U6104 (N_6104,N_3200,N_3395);
and U6105 (N_6105,N_2389,N_3780);
nand U6106 (N_6106,N_2651,N_3045);
nand U6107 (N_6107,N_3521,N_1145);
nor U6108 (N_6108,N_2603,N_1735);
and U6109 (N_6109,N_3229,N_2106);
or U6110 (N_6110,N_1699,N_3503);
or U6111 (N_6111,N_2320,N_923);
nand U6112 (N_6112,N_2874,N_907);
and U6113 (N_6113,N_1297,N_465);
nor U6114 (N_6114,N_1027,N_829);
nand U6115 (N_6115,N_847,N_1959);
nor U6116 (N_6116,N_3199,N_2953);
nor U6117 (N_6117,N_785,N_3421);
and U6118 (N_6118,N_709,N_51);
nor U6119 (N_6119,N_949,N_3108);
nand U6120 (N_6120,N_828,N_3903);
nor U6121 (N_6121,N_611,N_2646);
xor U6122 (N_6122,N_91,N_1626);
nand U6123 (N_6123,N_3342,N_827);
xor U6124 (N_6124,N_93,N_3779);
xnor U6125 (N_6125,N_1396,N_1161);
or U6126 (N_6126,N_3948,N_109);
or U6127 (N_6127,N_730,N_727);
xnor U6128 (N_6128,N_1453,N_874);
and U6129 (N_6129,N_1687,N_267);
nand U6130 (N_6130,N_3405,N_564);
and U6131 (N_6131,N_2975,N_1487);
or U6132 (N_6132,N_420,N_474);
nand U6133 (N_6133,N_3964,N_1475);
nor U6134 (N_6134,N_1536,N_1306);
nand U6135 (N_6135,N_1241,N_1308);
nand U6136 (N_6136,N_3667,N_2692);
and U6137 (N_6137,N_735,N_2337);
nand U6138 (N_6138,N_954,N_2836);
and U6139 (N_6139,N_1475,N_434);
or U6140 (N_6140,N_435,N_2529);
nand U6141 (N_6141,N_3341,N_1245);
xor U6142 (N_6142,N_2367,N_3063);
nor U6143 (N_6143,N_2605,N_3060);
xnor U6144 (N_6144,N_3529,N_2330);
or U6145 (N_6145,N_515,N_3565);
and U6146 (N_6146,N_706,N_2375);
nor U6147 (N_6147,N_1050,N_1905);
and U6148 (N_6148,N_1609,N_1762);
xor U6149 (N_6149,N_2429,N_2070);
nand U6150 (N_6150,N_980,N_2972);
and U6151 (N_6151,N_16,N_1910);
or U6152 (N_6152,N_466,N_2684);
nand U6153 (N_6153,N_1808,N_978);
nand U6154 (N_6154,N_3087,N_3813);
nor U6155 (N_6155,N_3233,N_1464);
or U6156 (N_6156,N_592,N_346);
nor U6157 (N_6157,N_533,N_3648);
nor U6158 (N_6158,N_3707,N_3322);
nor U6159 (N_6159,N_2749,N_2902);
or U6160 (N_6160,N_2599,N_685);
nor U6161 (N_6161,N_2671,N_1025);
nand U6162 (N_6162,N_1383,N_3299);
and U6163 (N_6163,N_1838,N_2716);
xor U6164 (N_6164,N_483,N_2551);
nand U6165 (N_6165,N_1842,N_1888);
and U6166 (N_6166,N_1323,N_2736);
nor U6167 (N_6167,N_296,N_908);
nand U6168 (N_6168,N_1207,N_2463);
nand U6169 (N_6169,N_849,N_3322);
xor U6170 (N_6170,N_1085,N_1087);
or U6171 (N_6171,N_1481,N_398);
and U6172 (N_6172,N_2019,N_2480);
xor U6173 (N_6173,N_1499,N_146);
and U6174 (N_6174,N_2108,N_3030);
or U6175 (N_6175,N_1457,N_3633);
nor U6176 (N_6176,N_1803,N_1184);
or U6177 (N_6177,N_602,N_2457);
nand U6178 (N_6178,N_1710,N_362);
nor U6179 (N_6179,N_2619,N_1412);
or U6180 (N_6180,N_578,N_1479);
nand U6181 (N_6181,N_3726,N_368);
xor U6182 (N_6182,N_11,N_3737);
or U6183 (N_6183,N_3622,N_2611);
xnor U6184 (N_6184,N_748,N_127);
and U6185 (N_6185,N_738,N_3838);
and U6186 (N_6186,N_1535,N_1236);
or U6187 (N_6187,N_2816,N_3811);
nor U6188 (N_6188,N_263,N_1344);
and U6189 (N_6189,N_632,N_1452);
and U6190 (N_6190,N_3423,N_3794);
or U6191 (N_6191,N_352,N_2605);
or U6192 (N_6192,N_1099,N_3081);
and U6193 (N_6193,N_1857,N_574);
nand U6194 (N_6194,N_3557,N_381);
nand U6195 (N_6195,N_2013,N_1408);
and U6196 (N_6196,N_3067,N_3318);
or U6197 (N_6197,N_1290,N_3955);
nor U6198 (N_6198,N_1605,N_3109);
nor U6199 (N_6199,N_1725,N_1174);
nand U6200 (N_6200,N_2316,N_3857);
and U6201 (N_6201,N_113,N_206);
or U6202 (N_6202,N_1662,N_3252);
or U6203 (N_6203,N_3674,N_1057);
nand U6204 (N_6204,N_301,N_2518);
and U6205 (N_6205,N_2547,N_53);
nor U6206 (N_6206,N_1808,N_3497);
and U6207 (N_6207,N_465,N_1657);
and U6208 (N_6208,N_539,N_1784);
nor U6209 (N_6209,N_189,N_1908);
or U6210 (N_6210,N_2181,N_3221);
nor U6211 (N_6211,N_2007,N_2792);
xnor U6212 (N_6212,N_2748,N_3909);
or U6213 (N_6213,N_2788,N_2559);
or U6214 (N_6214,N_3077,N_2999);
nand U6215 (N_6215,N_2863,N_1853);
and U6216 (N_6216,N_1034,N_2251);
xor U6217 (N_6217,N_2593,N_3051);
xor U6218 (N_6218,N_2608,N_3113);
xor U6219 (N_6219,N_263,N_473);
and U6220 (N_6220,N_1792,N_3030);
nor U6221 (N_6221,N_1168,N_2026);
and U6222 (N_6222,N_2946,N_1175);
nand U6223 (N_6223,N_1145,N_694);
nor U6224 (N_6224,N_249,N_3214);
nor U6225 (N_6225,N_2401,N_2154);
nor U6226 (N_6226,N_2062,N_221);
nand U6227 (N_6227,N_2840,N_3108);
xnor U6228 (N_6228,N_2202,N_2684);
xor U6229 (N_6229,N_1035,N_2378);
nand U6230 (N_6230,N_2785,N_738);
and U6231 (N_6231,N_1464,N_598);
xnor U6232 (N_6232,N_3536,N_3284);
nand U6233 (N_6233,N_130,N_2230);
xnor U6234 (N_6234,N_1703,N_2699);
xor U6235 (N_6235,N_1844,N_2551);
nor U6236 (N_6236,N_3170,N_2288);
nand U6237 (N_6237,N_3334,N_539);
and U6238 (N_6238,N_3719,N_593);
and U6239 (N_6239,N_3008,N_2783);
and U6240 (N_6240,N_1246,N_662);
and U6241 (N_6241,N_276,N_704);
nor U6242 (N_6242,N_975,N_2442);
or U6243 (N_6243,N_979,N_1385);
and U6244 (N_6244,N_1788,N_2972);
and U6245 (N_6245,N_1642,N_382);
xnor U6246 (N_6246,N_1273,N_891);
or U6247 (N_6247,N_3587,N_3670);
nand U6248 (N_6248,N_2546,N_2267);
nor U6249 (N_6249,N_386,N_1711);
xnor U6250 (N_6250,N_3586,N_235);
or U6251 (N_6251,N_3146,N_237);
and U6252 (N_6252,N_2040,N_3075);
nand U6253 (N_6253,N_3349,N_1546);
and U6254 (N_6254,N_509,N_948);
and U6255 (N_6255,N_1582,N_1951);
xor U6256 (N_6256,N_2222,N_3145);
xor U6257 (N_6257,N_2195,N_1499);
xor U6258 (N_6258,N_2695,N_2577);
xnor U6259 (N_6259,N_745,N_2611);
and U6260 (N_6260,N_2730,N_2380);
and U6261 (N_6261,N_2952,N_2567);
nand U6262 (N_6262,N_2771,N_3874);
nand U6263 (N_6263,N_3411,N_2000);
xnor U6264 (N_6264,N_2703,N_3028);
and U6265 (N_6265,N_1312,N_209);
nor U6266 (N_6266,N_2378,N_765);
nor U6267 (N_6267,N_90,N_1255);
or U6268 (N_6268,N_2009,N_710);
or U6269 (N_6269,N_149,N_1152);
xnor U6270 (N_6270,N_2441,N_3714);
nand U6271 (N_6271,N_2430,N_371);
nor U6272 (N_6272,N_569,N_3634);
or U6273 (N_6273,N_3921,N_2777);
or U6274 (N_6274,N_957,N_600);
nand U6275 (N_6275,N_2134,N_574);
xnor U6276 (N_6276,N_1279,N_3283);
xnor U6277 (N_6277,N_2075,N_1898);
xnor U6278 (N_6278,N_887,N_2998);
nand U6279 (N_6279,N_1297,N_3535);
nand U6280 (N_6280,N_1533,N_342);
and U6281 (N_6281,N_187,N_1003);
nor U6282 (N_6282,N_2810,N_3206);
or U6283 (N_6283,N_3903,N_1559);
nor U6284 (N_6284,N_2904,N_3407);
nand U6285 (N_6285,N_1450,N_3398);
and U6286 (N_6286,N_3957,N_2136);
or U6287 (N_6287,N_1135,N_2146);
nor U6288 (N_6288,N_2472,N_2480);
xor U6289 (N_6289,N_2395,N_3496);
nand U6290 (N_6290,N_2363,N_625);
xnor U6291 (N_6291,N_3641,N_3102);
nor U6292 (N_6292,N_3129,N_589);
nor U6293 (N_6293,N_3285,N_3394);
nand U6294 (N_6294,N_1512,N_1198);
and U6295 (N_6295,N_3475,N_2921);
nand U6296 (N_6296,N_2224,N_1560);
or U6297 (N_6297,N_2142,N_1412);
or U6298 (N_6298,N_2829,N_1840);
nor U6299 (N_6299,N_2434,N_477);
nor U6300 (N_6300,N_3211,N_863);
nand U6301 (N_6301,N_1505,N_2857);
or U6302 (N_6302,N_192,N_486);
nor U6303 (N_6303,N_1639,N_1490);
nand U6304 (N_6304,N_1934,N_2324);
and U6305 (N_6305,N_710,N_828);
nand U6306 (N_6306,N_3563,N_983);
xnor U6307 (N_6307,N_1667,N_3360);
xnor U6308 (N_6308,N_1375,N_3990);
nand U6309 (N_6309,N_3914,N_1741);
or U6310 (N_6310,N_3539,N_2133);
nand U6311 (N_6311,N_1455,N_3088);
nand U6312 (N_6312,N_906,N_3970);
nand U6313 (N_6313,N_1784,N_1619);
nand U6314 (N_6314,N_1751,N_3863);
or U6315 (N_6315,N_1333,N_2177);
nand U6316 (N_6316,N_3571,N_2718);
nor U6317 (N_6317,N_2886,N_1113);
or U6318 (N_6318,N_3118,N_291);
xnor U6319 (N_6319,N_3381,N_2266);
xor U6320 (N_6320,N_841,N_1623);
xnor U6321 (N_6321,N_834,N_1491);
nor U6322 (N_6322,N_2527,N_196);
nand U6323 (N_6323,N_1297,N_812);
nand U6324 (N_6324,N_2355,N_2184);
or U6325 (N_6325,N_2682,N_3567);
nor U6326 (N_6326,N_341,N_3223);
or U6327 (N_6327,N_2992,N_1394);
xor U6328 (N_6328,N_24,N_140);
and U6329 (N_6329,N_1716,N_1988);
and U6330 (N_6330,N_751,N_1777);
and U6331 (N_6331,N_18,N_2339);
xnor U6332 (N_6332,N_892,N_455);
xor U6333 (N_6333,N_458,N_2403);
and U6334 (N_6334,N_842,N_1332);
and U6335 (N_6335,N_307,N_164);
nand U6336 (N_6336,N_103,N_819);
nand U6337 (N_6337,N_2924,N_3946);
and U6338 (N_6338,N_2405,N_2353);
and U6339 (N_6339,N_2711,N_3093);
nor U6340 (N_6340,N_2407,N_1864);
nand U6341 (N_6341,N_2363,N_109);
nand U6342 (N_6342,N_558,N_900);
and U6343 (N_6343,N_1289,N_752);
nor U6344 (N_6344,N_2472,N_613);
nand U6345 (N_6345,N_1027,N_2933);
nor U6346 (N_6346,N_1172,N_61);
nor U6347 (N_6347,N_3260,N_1954);
and U6348 (N_6348,N_1846,N_3024);
xor U6349 (N_6349,N_2559,N_1240);
and U6350 (N_6350,N_1535,N_1262);
and U6351 (N_6351,N_774,N_1277);
xnor U6352 (N_6352,N_3636,N_2748);
and U6353 (N_6353,N_3802,N_654);
and U6354 (N_6354,N_692,N_1964);
and U6355 (N_6355,N_923,N_3522);
nand U6356 (N_6356,N_1726,N_583);
nor U6357 (N_6357,N_652,N_3169);
nand U6358 (N_6358,N_715,N_2757);
nor U6359 (N_6359,N_42,N_1801);
nand U6360 (N_6360,N_530,N_3608);
xor U6361 (N_6361,N_1367,N_2168);
and U6362 (N_6362,N_2441,N_3006);
or U6363 (N_6363,N_2770,N_2914);
nand U6364 (N_6364,N_3743,N_3759);
nand U6365 (N_6365,N_3313,N_2808);
or U6366 (N_6366,N_3061,N_2916);
nand U6367 (N_6367,N_1036,N_1258);
xnor U6368 (N_6368,N_3895,N_676);
nand U6369 (N_6369,N_1569,N_2849);
xnor U6370 (N_6370,N_2474,N_2483);
nor U6371 (N_6371,N_3384,N_578);
and U6372 (N_6372,N_815,N_876);
and U6373 (N_6373,N_2216,N_1559);
nand U6374 (N_6374,N_824,N_2079);
and U6375 (N_6375,N_274,N_1664);
and U6376 (N_6376,N_3598,N_3891);
nand U6377 (N_6377,N_227,N_2060);
or U6378 (N_6378,N_2650,N_331);
and U6379 (N_6379,N_724,N_2434);
nor U6380 (N_6380,N_276,N_3922);
or U6381 (N_6381,N_2321,N_2564);
or U6382 (N_6382,N_1285,N_3259);
nand U6383 (N_6383,N_2640,N_2209);
xnor U6384 (N_6384,N_35,N_2051);
nand U6385 (N_6385,N_3601,N_2344);
nand U6386 (N_6386,N_1704,N_1255);
nand U6387 (N_6387,N_1216,N_2843);
nor U6388 (N_6388,N_3759,N_3392);
and U6389 (N_6389,N_719,N_1346);
nor U6390 (N_6390,N_2769,N_1310);
nand U6391 (N_6391,N_2689,N_3364);
and U6392 (N_6392,N_3401,N_3937);
nand U6393 (N_6393,N_378,N_751);
nand U6394 (N_6394,N_2215,N_2682);
and U6395 (N_6395,N_2779,N_388);
nand U6396 (N_6396,N_3970,N_1439);
xnor U6397 (N_6397,N_1940,N_2130);
nor U6398 (N_6398,N_924,N_2547);
nor U6399 (N_6399,N_3510,N_534);
or U6400 (N_6400,N_1645,N_2855);
nor U6401 (N_6401,N_460,N_2286);
or U6402 (N_6402,N_3307,N_208);
xnor U6403 (N_6403,N_177,N_3924);
xnor U6404 (N_6404,N_2530,N_316);
and U6405 (N_6405,N_971,N_383);
xnor U6406 (N_6406,N_2621,N_2397);
nor U6407 (N_6407,N_1476,N_1780);
xnor U6408 (N_6408,N_530,N_2634);
or U6409 (N_6409,N_3398,N_3352);
xor U6410 (N_6410,N_1702,N_1277);
xor U6411 (N_6411,N_3701,N_3613);
nand U6412 (N_6412,N_1499,N_2447);
or U6413 (N_6413,N_2202,N_369);
nand U6414 (N_6414,N_516,N_1795);
xnor U6415 (N_6415,N_1613,N_837);
or U6416 (N_6416,N_3876,N_3162);
or U6417 (N_6417,N_1002,N_3736);
xnor U6418 (N_6418,N_136,N_2223);
nand U6419 (N_6419,N_2393,N_3185);
nand U6420 (N_6420,N_2405,N_3923);
nand U6421 (N_6421,N_539,N_3928);
nor U6422 (N_6422,N_1568,N_2511);
and U6423 (N_6423,N_1606,N_160);
nand U6424 (N_6424,N_2895,N_900);
nand U6425 (N_6425,N_638,N_603);
nor U6426 (N_6426,N_1494,N_2195);
xor U6427 (N_6427,N_2221,N_1012);
nand U6428 (N_6428,N_3658,N_2992);
or U6429 (N_6429,N_2977,N_2244);
or U6430 (N_6430,N_873,N_184);
nand U6431 (N_6431,N_1684,N_905);
nor U6432 (N_6432,N_1401,N_1896);
or U6433 (N_6433,N_3728,N_3468);
xor U6434 (N_6434,N_2646,N_0);
xnor U6435 (N_6435,N_3703,N_1419);
nand U6436 (N_6436,N_1863,N_1602);
nand U6437 (N_6437,N_831,N_2743);
nor U6438 (N_6438,N_2987,N_1123);
xnor U6439 (N_6439,N_732,N_1482);
and U6440 (N_6440,N_411,N_3833);
xor U6441 (N_6441,N_785,N_327);
and U6442 (N_6442,N_3776,N_3351);
xnor U6443 (N_6443,N_2306,N_1995);
and U6444 (N_6444,N_1987,N_547);
and U6445 (N_6445,N_1140,N_2714);
nand U6446 (N_6446,N_2481,N_2778);
nor U6447 (N_6447,N_544,N_1855);
xor U6448 (N_6448,N_581,N_61);
nand U6449 (N_6449,N_299,N_1860);
nand U6450 (N_6450,N_2380,N_1194);
and U6451 (N_6451,N_2142,N_145);
xor U6452 (N_6452,N_3146,N_3917);
nand U6453 (N_6453,N_3619,N_972);
nor U6454 (N_6454,N_2684,N_2708);
or U6455 (N_6455,N_2942,N_3597);
nor U6456 (N_6456,N_858,N_3451);
nand U6457 (N_6457,N_768,N_3824);
and U6458 (N_6458,N_3505,N_118);
xor U6459 (N_6459,N_3174,N_875);
or U6460 (N_6460,N_3620,N_2573);
or U6461 (N_6461,N_2817,N_1609);
and U6462 (N_6462,N_2789,N_16);
nor U6463 (N_6463,N_2065,N_1580);
or U6464 (N_6464,N_3267,N_1063);
xnor U6465 (N_6465,N_1682,N_2009);
xor U6466 (N_6466,N_2662,N_3950);
xnor U6467 (N_6467,N_2941,N_3096);
xnor U6468 (N_6468,N_3994,N_2835);
or U6469 (N_6469,N_3082,N_2155);
xor U6470 (N_6470,N_3526,N_447);
and U6471 (N_6471,N_3835,N_3983);
or U6472 (N_6472,N_3996,N_1209);
nor U6473 (N_6473,N_3311,N_200);
nand U6474 (N_6474,N_257,N_572);
nand U6475 (N_6475,N_1615,N_2192);
and U6476 (N_6476,N_241,N_2598);
nor U6477 (N_6477,N_1915,N_2752);
or U6478 (N_6478,N_216,N_2099);
nor U6479 (N_6479,N_3876,N_90);
xnor U6480 (N_6480,N_1095,N_1589);
or U6481 (N_6481,N_842,N_2659);
xor U6482 (N_6482,N_2699,N_1819);
xor U6483 (N_6483,N_3492,N_577);
and U6484 (N_6484,N_3790,N_3279);
nand U6485 (N_6485,N_211,N_3871);
or U6486 (N_6486,N_961,N_2710);
nor U6487 (N_6487,N_256,N_549);
xnor U6488 (N_6488,N_1654,N_1905);
and U6489 (N_6489,N_2124,N_1247);
and U6490 (N_6490,N_1244,N_3847);
or U6491 (N_6491,N_3142,N_2103);
nor U6492 (N_6492,N_2846,N_3352);
nor U6493 (N_6493,N_809,N_2875);
nand U6494 (N_6494,N_2518,N_1842);
and U6495 (N_6495,N_3202,N_2679);
or U6496 (N_6496,N_3075,N_2365);
nor U6497 (N_6497,N_321,N_569);
nand U6498 (N_6498,N_3709,N_1510);
nor U6499 (N_6499,N_3999,N_3383);
xnor U6500 (N_6500,N_3185,N_2876);
nor U6501 (N_6501,N_1094,N_1048);
nand U6502 (N_6502,N_1305,N_926);
and U6503 (N_6503,N_3148,N_348);
and U6504 (N_6504,N_216,N_3996);
or U6505 (N_6505,N_2177,N_621);
or U6506 (N_6506,N_2954,N_2706);
xor U6507 (N_6507,N_553,N_1801);
xor U6508 (N_6508,N_2409,N_1119);
nand U6509 (N_6509,N_2128,N_2047);
or U6510 (N_6510,N_3928,N_650);
nand U6511 (N_6511,N_3073,N_908);
or U6512 (N_6512,N_1171,N_359);
or U6513 (N_6513,N_606,N_3644);
nand U6514 (N_6514,N_907,N_3747);
nand U6515 (N_6515,N_2239,N_2101);
and U6516 (N_6516,N_2362,N_1110);
xnor U6517 (N_6517,N_2106,N_1034);
and U6518 (N_6518,N_1913,N_1124);
nand U6519 (N_6519,N_1521,N_392);
nor U6520 (N_6520,N_999,N_3043);
or U6521 (N_6521,N_790,N_196);
nand U6522 (N_6522,N_357,N_2140);
and U6523 (N_6523,N_3128,N_1127);
nand U6524 (N_6524,N_488,N_2513);
nand U6525 (N_6525,N_3461,N_455);
or U6526 (N_6526,N_1788,N_3539);
or U6527 (N_6527,N_1509,N_3791);
xnor U6528 (N_6528,N_111,N_3085);
or U6529 (N_6529,N_116,N_2378);
nor U6530 (N_6530,N_369,N_862);
nand U6531 (N_6531,N_1087,N_2462);
nand U6532 (N_6532,N_2859,N_2526);
nand U6533 (N_6533,N_852,N_2787);
nand U6534 (N_6534,N_2011,N_2937);
or U6535 (N_6535,N_2286,N_2446);
and U6536 (N_6536,N_1368,N_687);
xnor U6537 (N_6537,N_844,N_2406);
xor U6538 (N_6538,N_1753,N_3261);
xnor U6539 (N_6539,N_912,N_2715);
xnor U6540 (N_6540,N_1770,N_3072);
nand U6541 (N_6541,N_461,N_2486);
nor U6542 (N_6542,N_710,N_2061);
or U6543 (N_6543,N_2406,N_1863);
xnor U6544 (N_6544,N_745,N_254);
or U6545 (N_6545,N_844,N_2194);
nand U6546 (N_6546,N_3489,N_2048);
nand U6547 (N_6547,N_3163,N_193);
or U6548 (N_6548,N_595,N_1596);
nor U6549 (N_6549,N_3441,N_1123);
nor U6550 (N_6550,N_2979,N_251);
nand U6551 (N_6551,N_3900,N_2594);
or U6552 (N_6552,N_2845,N_2201);
nor U6553 (N_6553,N_592,N_505);
xnor U6554 (N_6554,N_1587,N_3800);
and U6555 (N_6555,N_2018,N_2683);
xor U6556 (N_6556,N_2107,N_1375);
and U6557 (N_6557,N_270,N_2584);
xor U6558 (N_6558,N_3881,N_2580);
or U6559 (N_6559,N_788,N_516);
nand U6560 (N_6560,N_347,N_1547);
xnor U6561 (N_6561,N_1463,N_1751);
or U6562 (N_6562,N_3232,N_639);
nand U6563 (N_6563,N_607,N_2814);
nor U6564 (N_6564,N_1124,N_1174);
nand U6565 (N_6565,N_1772,N_1778);
xor U6566 (N_6566,N_220,N_59);
xor U6567 (N_6567,N_3012,N_3200);
nand U6568 (N_6568,N_3904,N_936);
or U6569 (N_6569,N_1132,N_1491);
xnor U6570 (N_6570,N_2117,N_1810);
nor U6571 (N_6571,N_590,N_2995);
nor U6572 (N_6572,N_1138,N_1993);
and U6573 (N_6573,N_2696,N_2406);
or U6574 (N_6574,N_1791,N_1994);
nor U6575 (N_6575,N_328,N_1681);
xnor U6576 (N_6576,N_3997,N_3705);
or U6577 (N_6577,N_1496,N_3761);
and U6578 (N_6578,N_3566,N_2077);
nor U6579 (N_6579,N_3706,N_2093);
and U6580 (N_6580,N_1054,N_3393);
and U6581 (N_6581,N_1142,N_2652);
nand U6582 (N_6582,N_2030,N_446);
and U6583 (N_6583,N_2121,N_1362);
nor U6584 (N_6584,N_1789,N_3704);
nor U6585 (N_6585,N_3142,N_2292);
and U6586 (N_6586,N_2958,N_1316);
or U6587 (N_6587,N_2684,N_171);
and U6588 (N_6588,N_3595,N_967);
nand U6589 (N_6589,N_2222,N_1442);
or U6590 (N_6590,N_2874,N_662);
nand U6591 (N_6591,N_3437,N_1287);
nand U6592 (N_6592,N_1127,N_1065);
or U6593 (N_6593,N_3107,N_1960);
nand U6594 (N_6594,N_3592,N_1480);
nand U6595 (N_6595,N_2044,N_1703);
xor U6596 (N_6596,N_1664,N_1935);
or U6597 (N_6597,N_2629,N_2032);
xor U6598 (N_6598,N_3461,N_400);
nand U6599 (N_6599,N_2747,N_1525);
or U6600 (N_6600,N_2518,N_940);
or U6601 (N_6601,N_2578,N_716);
xor U6602 (N_6602,N_3516,N_2001);
nand U6603 (N_6603,N_3473,N_705);
nor U6604 (N_6604,N_923,N_2549);
or U6605 (N_6605,N_103,N_3962);
nor U6606 (N_6606,N_3154,N_1860);
and U6607 (N_6607,N_2518,N_3145);
and U6608 (N_6608,N_311,N_529);
or U6609 (N_6609,N_1135,N_1624);
or U6610 (N_6610,N_2134,N_3602);
nor U6611 (N_6611,N_2681,N_2299);
xor U6612 (N_6612,N_1448,N_497);
and U6613 (N_6613,N_2995,N_3307);
nor U6614 (N_6614,N_2972,N_808);
xnor U6615 (N_6615,N_2603,N_1366);
and U6616 (N_6616,N_2825,N_3174);
nand U6617 (N_6617,N_2598,N_1215);
nand U6618 (N_6618,N_2021,N_3964);
nor U6619 (N_6619,N_877,N_1553);
nor U6620 (N_6620,N_137,N_2775);
and U6621 (N_6621,N_3759,N_1514);
nand U6622 (N_6622,N_672,N_1624);
and U6623 (N_6623,N_716,N_3493);
or U6624 (N_6624,N_3813,N_2219);
xnor U6625 (N_6625,N_2886,N_3356);
or U6626 (N_6626,N_1444,N_300);
nor U6627 (N_6627,N_2768,N_554);
nand U6628 (N_6628,N_974,N_3149);
or U6629 (N_6629,N_1491,N_2096);
nand U6630 (N_6630,N_3678,N_2210);
or U6631 (N_6631,N_2267,N_467);
and U6632 (N_6632,N_638,N_1392);
or U6633 (N_6633,N_2271,N_1980);
or U6634 (N_6634,N_3705,N_1146);
nor U6635 (N_6635,N_1246,N_3332);
or U6636 (N_6636,N_3035,N_3577);
or U6637 (N_6637,N_969,N_869);
xnor U6638 (N_6638,N_2685,N_3426);
nor U6639 (N_6639,N_1976,N_1380);
nand U6640 (N_6640,N_3038,N_986);
nand U6641 (N_6641,N_15,N_2783);
nand U6642 (N_6642,N_292,N_3100);
nand U6643 (N_6643,N_599,N_1989);
nand U6644 (N_6644,N_1734,N_2592);
and U6645 (N_6645,N_2147,N_2267);
nand U6646 (N_6646,N_3182,N_1615);
nand U6647 (N_6647,N_1032,N_898);
nor U6648 (N_6648,N_2902,N_2930);
nand U6649 (N_6649,N_2343,N_718);
or U6650 (N_6650,N_1843,N_3544);
xnor U6651 (N_6651,N_3807,N_2159);
nand U6652 (N_6652,N_1523,N_1143);
nand U6653 (N_6653,N_3263,N_2392);
nor U6654 (N_6654,N_2388,N_1810);
or U6655 (N_6655,N_2386,N_3179);
nand U6656 (N_6656,N_1179,N_3259);
nor U6657 (N_6657,N_53,N_2293);
xnor U6658 (N_6658,N_1908,N_1367);
and U6659 (N_6659,N_1637,N_2477);
and U6660 (N_6660,N_3024,N_3078);
nand U6661 (N_6661,N_717,N_2685);
nand U6662 (N_6662,N_2363,N_839);
nor U6663 (N_6663,N_684,N_960);
or U6664 (N_6664,N_3670,N_2271);
nand U6665 (N_6665,N_2532,N_59);
or U6666 (N_6666,N_3694,N_2995);
and U6667 (N_6667,N_1057,N_791);
nand U6668 (N_6668,N_2913,N_807);
xor U6669 (N_6669,N_2082,N_2435);
or U6670 (N_6670,N_2185,N_3081);
nor U6671 (N_6671,N_1599,N_2683);
or U6672 (N_6672,N_2351,N_1392);
xor U6673 (N_6673,N_1138,N_533);
and U6674 (N_6674,N_3458,N_1346);
xor U6675 (N_6675,N_1721,N_2908);
and U6676 (N_6676,N_2409,N_1064);
nand U6677 (N_6677,N_1719,N_2829);
xor U6678 (N_6678,N_1043,N_3691);
nor U6679 (N_6679,N_773,N_2041);
xnor U6680 (N_6680,N_1983,N_218);
or U6681 (N_6681,N_379,N_3225);
and U6682 (N_6682,N_3124,N_2933);
nand U6683 (N_6683,N_3184,N_2524);
or U6684 (N_6684,N_67,N_549);
nor U6685 (N_6685,N_173,N_1098);
nor U6686 (N_6686,N_2772,N_3702);
and U6687 (N_6687,N_3080,N_2973);
or U6688 (N_6688,N_2495,N_1298);
nand U6689 (N_6689,N_2996,N_3261);
nor U6690 (N_6690,N_2412,N_409);
and U6691 (N_6691,N_1118,N_1067);
and U6692 (N_6692,N_3314,N_2072);
or U6693 (N_6693,N_423,N_1776);
xor U6694 (N_6694,N_2184,N_442);
nor U6695 (N_6695,N_3537,N_2681);
nand U6696 (N_6696,N_510,N_3816);
and U6697 (N_6697,N_3757,N_1182);
nor U6698 (N_6698,N_3243,N_2939);
xor U6699 (N_6699,N_71,N_1821);
nor U6700 (N_6700,N_3421,N_1459);
nor U6701 (N_6701,N_2440,N_3817);
nand U6702 (N_6702,N_2982,N_143);
or U6703 (N_6703,N_1330,N_2536);
nand U6704 (N_6704,N_2584,N_182);
nand U6705 (N_6705,N_3629,N_3398);
nor U6706 (N_6706,N_488,N_3442);
and U6707 (N_6707,N_1750,N_2812);
or U6708 (N_6708,N_1670,N_2541);
xor U6709 (N_6709,N_112,N_281);
nand U6710 (N_6710,N_2494,N_1098);
nor U6711 (N_6711,N_1437,N_3667);
or U6712 (N_6712,N_2580,N_1196);
xnor U6713 (N_6713,N_1963,N_1921);
nor U6714 (N_6714,N_3097,N_3355);
xor U6715 (N_6715,N_1751,N_3497);
xor U6716 (N_6716,N_1321,N_3728);
nor U6717 (N_6717,N_122,N_521);
and U6718 (N_6718,N_2993,N_1453);
nor U6719 (N_6719,N_3254,N_3768);
xnor U6720 (N_6720,N_2278,N_1206);
and U6721 (N_6721,N_1342,N_409);
or U6722 (N_6722,N_1998,N_2280);
and U6723 (N_6723,N_2934,N_1733);
and U6724 (N_6724,N_127,N_407);
and U6725 (N_6725,N_3489,N_1448);
or U6726 (N_6726,N_452,N_2012);
nand U6727 (N_6727,N_3912,N_494);
xnor U6728 (N_6728,N_52,N_3914);
and U6729 (N_6729,N_1198,N_429);
nor U6730 (N_6730,N_1337,N_3955);
or U6731 (N_6731,N_1999,N_1723);
xor U6732 (N_6732,N_1363,N_1231);
and U6733 (N_6733,N_55,N_1484);
xor U6734 (N_6734,N_788,N_88);
nand U6735 (N_6735,N_3878,N_776);
nor U6736 (N_6736,N_824,N_2978);
or U6737 (N_6737,N_3526,N_44);
nand U6738 (N_6738,N_1147,N_1771);
or U6739 (N_6739,N_2619,N_36);
and U6740 (N_6740,N_2126,N_1293);
or U6741 (N_6741,N_792,N_693);
nor U6742 (N_6742,N_2163,N_2192);
and U6743 (N_6743,N_459,N_3102);
nand U6744 (N_6744,N_2609,N_156);
or U6745 (N_6745,N_1616,N_3752);
nor U6746 (N_6746,N_296,N_2459);
nor U6747 (N_6747,N_2621,N_2004);
xnor U6748 (N_6748,N_1359,N_1498);
or U6749 (N_6749,N_89,N_2865);
nand U6750 (N_6750,N_2749,N_1224);
nand U6751 (N_6751,N_2651,N_1885);
or U6752 (N_6752,N_1462,N_586);
or U6753 (N_6753,N_2640,N_2816);
and U6754 (N_6754,N_1777,N_1714);
or U6755 (N_6755,N_313,N_25);
nand U6756 (N_6756,N_3224,N_2952);
and U6757 (N_6757,N_268,N_2949);
nor U6758 (N_6758,N_44,N_2927);
xor U6759 (N_6759,N_3290,N_3043);
or U6760 (N_6760,N_609,N_2125);
and U6761 (N_6761,N_835,N_1143);
nand U6762 (N_6762,N_124,N_2744);
xor U6763 (N_6763,N_1076,N_648);
or U6764 (N_6764,N_1867,N_3004);
nor U6765 (N_6765,N_3487,N_1263);
or U6766 (N_6766,N_1310,N_1304);
nand U6767 (N_6767,N_948,N_3000);
xor U6768 (N_6768,N_2113,N_3047);
xor U6769 (N_6769,N_2736,N_3627);
nand U6770 (N_6770,N_2803,N_2925);
or U6771 (N_6771,N_447,N_519);
nand U6772 (N_6772,N_3936,N_2317);
or U6773 (N_6773,N_1000,N_521);
nor U6774 (N_6774,N_2435,N_3723);
or U6775 (N_6775,N_139,N_738);
or U6776 (N_6776,N_2149,N_602);
and U6777 (N_6777,N_3336,N_3088);
and U6778 (N_6778,N_3579,N_2512);
nand U6779 (N_6779,N_1777,N_2455);
or U6780 (N_6780,N_3324,N_981);
nor U6781 (N_6781,N_1415,N_1178);
nor U6782 (N_6782,N_762,N_952);
nand U6783 (N_6783,N_633,N_736);
nand U6784 (N_6784,N_2242,N_3596);
nand U6785 (N_6785,N_523,N_1519);
or U6786 (N_6786,N_2011,N_1001);
nor U6787 (N_6787,N_111,N_212);
or U6788 (N_6788,N_3047,N_1540);
nand U6789 (N_6789,N_1874,N_2028);
xnor U6790 (N_6790,N_1392,N_2977);
or U6791 (N_6791,N_815,N_2189);
and U6792 (N_6792,N_924,N_3089);
xor U6793 (N_6793,N_3098,N_1079);
or U6794 (N_6794,N_3203,N_2103);
nand U6795 (N_6795,N_1994,N_2411);
or U6796 (N_6796,N_2376,N_2556);
nand U6797 (N_6797,N_1987,N_2283);
nor U6798 (N_6798,N_3106,N_3122);
nand U6799 (N_6799,N_112,N_3153);
or U6800 (N_6800,N_2870,N_363);
nor U6801 (N_6801,N_3224,N_3716);
nand U6802 (N_6802,N_827,N_2853);
nand U6803 (N_6803,N_3575,N_2566);
nand U6804 (N_6804,N_1512,N_1913);
nor U6805 (N_6805,N_1701,N_3898);
nand U6806 (N_6806,N_1426,N_2778);
nor U6807 (N_6807,N_1027,N_876);
or U6808 (N_6808,N_2400,N_1543);
or U6809 (N_6809,N_1520,N_3025);
or U6810 (N_6810,N_3960,N_2907);
nand U6811 (N_6811,N_3635,N_671);
xnor U6812 (N_6812,N_1969,N_3004);
xnor U6813 (N_6813,N_1885,N_1839);
or U6814 (N_6814,N_1178,N_2945);
nand U6815 (N_6815,N_2392,N_2081);
nand U6816 (N_6816,N_3072,N_3340);
xnor U6817 (N_6817,N_1056,N_1398);
nand U6818 (N_6818,N_2052,N_2349);
xor U6819 (N_6819,N_719,N_2402);
or U6820 (N_6820,N_1484,N_1074);
or U6821 (N_6821,N_734,N_3263);
nor U6822 (N_6822,N_1001,N_322);
nor U6823 (N_6823,N_416,N_3780);
or U6824 (N_6824,N_3735,N_701);
and U6825 (N_6825,N_2333,N_932);
nor U6826 (N_6826,N_2825,N_620);
or U6827 (N_6827,N_1171,N_487);
and U6828 (N_6828,N_2828,N_3662);
and U6829 (N_6829,N_478,N_2254);
xor U6830 (N_6830,N_660,N_2960);
nor U6831 (N_6831,N_1990,N_3990);
nand U6832 (N_6832,N_851,N_2486);
and U6833 (N_6833,N_3090,N_889);
and U6834 (N_6834,N_3452,N_2252);
and U6835 (N_6835,N_933,N_457);
nor U6836 (N_6836,N_839,N_2626);
xnor U6837 (N_6837,N_1519,N_2295);
or U6838 (N_6838,N_1843,N_490);
xor U6839 (N_6839,N_275,N_1532);
and U6840 (N_6840,N_869,N_3211);
nand U6841 (N_6841,N_1588,N_1218);
xor U6842 (N_6842,N_2438,N_2936);
nor U6843 (N_6843,N_2243,N_2866);
and U6844 (N_6844,N_3531,N_2806);
and U6845 (N_6845,N_2206,N_1207);
nand U6846 (N_6846,N_3142,N_204);
nor U6847 (N_6847,N_478,N_1981);
xnor U6848 (N_6848,N_2009,N_2125);
and U6849 (N_6849,N_1683,N_1823);
and U6850 (N_6850,N_2438,N_721);
and U6851 (N_6851,N_2130,N_2418);
xor U6852 (N_6852,N_3396,N_773);
nor U6853 (N_6853,N_3530,N_3439);
nor U6854 (N_6854,N_1759,N_324);
xnor U6855 (N_6855,N_3823,N_3906);
or U6856 (N_6856,N_790,N_3986);
nand U6857 (N_6857,N_3762,N_804);
xor U6858 (N_6858,N_2768,N_74);
nor U6859 (N_6859,N_1793,N_2491);
xnor U6860 (N_6860,N_3279,N_2155);
xnor U6861 (N_6861,N_38,N_1589);
or U6862 (N_6862,N_1386,N_2429);
nand U6863 (N_6863,N_167,N_1484);
xnor U6864 (N_6864,N_126,N_253);
and U6865 (N_6865,N_3012,N_1003);
or U6866 (N_6866,N_3957,N_1320);
or U6867 (N_6867,N_1912,N_2384);
xor U6868 (N_6868,N_2889,N_1856);
xor U6869 (N_6869,N_507,N_2964);
or U6870 (N_6870,N_861,N_3754);
nand U6871 (N_6871,N_3985,N_374);
or U6872 (N_6872,N_1863,N_616);
xor U6873 (N_6873,N_1415,N_1956);
xor U6874 (N_6874,N_2888,N_613);
xor U6875 (N_6875,N_3074,N_3892);
xnor U6876 (N_6876,N_3510,N_3658);
or U6877 (N_6877,N_2311,N_3949);
xor U6878 (N_6878,N_3024,N_2074);
xnor U6879 (N_6879,N_1683,N_601);
nand U6880 (N_6880,N_1177,N_1369);
nor U6881 (N_6881,N_2967,N_646);
nor U6882 (N_6882,N_2743,N_504);
and U6883 (N_6883,N_293,N_434);
and U6884 (N_6884,N_3116,N_2346);
nand U6885 (N_6885,N_560,N_1602);
nand U6886 (N_6886,N_2188,N_2558);
and U6887 (N_6887,N_3394,N_1615);
and U6888 (N_6888,N_1309,N_1457);
xnor U6889 (N_6889,N_2534,N_1172);
and U6890 (N_6890,N_470,N_3918);
xor U6891 (N_6891,N_3438,N_3060);
nor U6892 (N_6892,N_2119,N_2449);
or U6893 (N_6893,N_3156,N_17);
and U6894 (N_6894,N_3549,N_318);
or U6895 (N_6895,N_3184,N_3105);
nor U6896 (N_6896,N_2086,N_3111);
xnor U6897 (N_6897,N_1656,N_3115);
nand U6898 (N_6898,N_2447,N_251);
nand U6899 (N_6899,N_3107,N_1269);
nand U6900 (N_6900,N_1640,N_3984);
nor U6901 (N_6901,N_1826,N_307);
xnor U6902 (N_6902,N_15,N_2938);
nand U6903 (N_6903,N_1930,N_532);
and U6904 (N_6904,N_801,N_2477);
nand U6905 (N_6905,N_3687,N_743);
nor U6906 (N_6906,N_2290,N_3094);
xnor U6907 (N_6907,N_3194,N_857);
or U6908 (N_6908,N_1987,N_1100);
nor U6909 (N_6909,N_22,N_504);
nand U6910 (N_6910,N_3695,N_2489);
nor U6911 (N_6911,N_49,N_1159);
xnor U6912 (N_6912,N_2318,N_505);
xnor U6913 (N_6913,N_2970,N_3781);
xor U6914 (N_6914,N_2999,N_627);
or U6915 (N_6915,N_3883,N_2777);
or U6916 (N_6916,N_577,N_896);
or U6917 (N_6917,N_3025,N_319);
and U6918 (N_6918,N_1726,N_1695);
nand U6919 (N_6919,N_2676,N_2548);
or U6920 (N_6920,N_2943,N_3555);
nor U6921 (N_6921,N_3121,N_1312);
nand U6922 (N_6922,N_1750,N_3666);
or U6923 (N_6923,N_2419,N_2258);
nand U6924 (N_6924,N_1394,N_832);
and U6925 (N_6925,N_2913,N_854);
nand U6926 (N_6926,N_540,N_513);
and U6927 (N_6927,N_2621,N_2406);
nor U6928 (N_6928,N_2568,N_1525);
nor U6929 (N_6929,N_1131,N_1304);
and U6930 (N_6930,N_2408,N_1233);
nor U6931 (N_6931,N_3301,N_3992);
or U6932 (N_6932,N_3256,N_3854);
nor U6933 (N_6933,N_3171,N_2821);
nor U6934 (N_6934,N_269,N_1497);
and U6935 (N_6935,N_2944,N_2435);
or U6936 (N_6936,N_1197,N_582);
or U6937 (N_6937,N_426,N_121);
nand U6938 (N_6938,N_1445,N_1861);
or U6939 (N_6939,N_1966,N_3380);
and U6940 (N_6940,N_1568,N_3212);
xnor U6941 (N_6941,N_3055,N_3280);
nor U6942 (N_6942,N_1284,N_133);
nor U6943 (N_6943,N_923,N_1092);
or U6944 (N_6944,N_2165,N_3776);
or U6945 (N_6945,N_1907,N_270);
nand U6946 (N_6946,N_2732,N_2444);
and U6947 (N_6947,N_3644,N_2749);
nand U6948 (N_6948,N_351,N_3130);
and U6949 (N_6949,N_3849,N_3045);
and U6950 (N_6950,N_3208,N_1486);
xnor U6951 (N_6951,N_2882,N_3091);
and U6952 (N_6952,N_2888,N_3593);
nor U6953 (N_6953,N_116,N_3902);
and U6954 (N_6954,N_1738,N_2873);
nand U6955 (N_6955,N_3499,N_1548);
nand U6956 (N_6956,N_3769,N_3617);
xnor U6957 (N_6957,N_750,N_3177);
nor U6958 (N_6958,N_338,N_47);
xor U6959 (N_6959,N_2878,N_3950);
and U6960 (N_6960,N_3672,N_2840);
xnor U6961 (N_6961,N_3815,N_523);
xnor U6962 (N_6962,N_1640,N_1084);
and U6963 (N_6963,N_44,N_273);
or U6964 (N_6964,N_2869,N_2726);
xnor U6965 (N_6965,N_2391,N_1212);
and U6966 (N_6966,N_3455,N_3572);
nand U6967 (N_6967,N_2238,N_1052);
nor U6968 (N_6968,N_2071,N_1834);
nor U6969 (N_6969,N_2065,N_3427);
or U6970 (N_6970,N_3367,N_224);
and U6971 (N_6971,N_1283,N_1025);
or U6972 (N_6972,N_3575,N_3659);
nor U6973 (N_6973,N_772,N_435);
and U6974 (N_6974,N_11,N_2595);
and U6975 (N_6975,N_3437,N_15);
nor U6976 (N_6976,N_3081,N_1718);
or U6977 (N_6977,N_3335,N_2859);
xor U6978 (N_6978,N_177,N_2309);
or U6979 (N_6979,N_1350,N_3386);
xnor U6980 (N_6980,N_410,N_3333);
xnor U6981 (N_6981,N_1990,N_2441);
xor U6982 (N_6982,N_1083,N_340);
or U6983 (N_6983,N_2314,N_1732);
or U6984 (N_6984,N_2873,N_3304);
nor U6985 (N_6985,N_3121,N_1663);
xnor U6986 (N_6986,N_124,N_1516);
and U6987 (N_6987,N_2569,N_2405);
nand U6988 (N_6988,N_1727,N_25);
and U6989 (N_6989,N_2234,N_361);
nor U6990 (N_6990,N_2850,N_3934);
nand U6991 (N_6991,N_94,N_79);
and U6992 (N_6992,N_3187,N_1638);
and U6993 (N_6993,N_832,N_3111);
and U6994 (N_6994,N_3257,N_2074);
or U6995 (N_6995,N_838,N_1987);
or U6996 (N_6996,N_2468,N_739);
nand U6997 (N_6997,N_1040,N_3177);
xnor U6998 (N_6998,N_517,N_3623);
nor U6999 (N_6999,N_2353,N_3571);
and U7000 (N_7000,N_3791,N_1834);
nor U7001 (N_7001,N_2101,N_1709);
or U7002 (N_7002,N_412,N_3345);
xnor U7003 (N_7003,N_649,N_565);
nor U7004 (N_7004,N_3142,N_755);
nor U7005 (N_7005,N_225,N_295);
nor U7006 (N_7006,N_2041,N_1949);
or U7007 (N_7007,N_418,N_162);
nand U7008 (N_7008,N_721,N_3301);
or U7009 (N_7009,N_2470,N_2913);
and U7010 (N_7010,N_1456,N_1240);
xnor U7011 (N_7011,N_1786,N_3703);
and U7012 (N_7012,N_2631,N_3581);
xnor U7013 (N_7013,N_1501,N_1614);
nand U7014 (N_7014,N_1609,N_3348);
xor U7015 (N_7015,N_1456,N_839);
or U7016 (N_7016,N_1019,N_3954);
and U7017 (N_7017,N_1957,N_3970);
nor U7018 (N_7018,N_3856,N_3367);
nor U7019 (N_7019,N_91,N_1299);
or U7020 (N_7020,N_1925,N_1462);
or U7021 (N_7021,N_1320,N_3598);
nor U7022 (N_7022,N_3758,N_3198);
nor U7023 (N_7023,N_162,N_2637);
and U7024 (N_7024,N_517,N_893);
or U7025 (N_7025,N_2405,N_3722);
and U7026 (N_7026,N_654,N_1703);
nand U7027 (N_7027,N_2500,N_1388);
or U7028 (N_7028,N_3724,N_2437);
and U7029 (N_7029,N_1278,N_2750);
xor U7030 (N_7030,N_325,N_3593);
or U7031 (N_7031,N_2909,N_1070);
nor U7032 (N_7032,N_225,N_1377);
or U7033 (N_7033,N_717,N_2117);
or U7034 (N_7034,N_2755,N_1534);
nor U7035 (N_7035,N_3736,N_3615);
xnor U7036 (N_7036,N_2721,N_3454);
xnor U7037 (N_7037,N_3897,N_3334);
and U7038 (N_7038,N_450,N_2131);
and U7039 (N_7039,N_2420,N_3193);
and U7040 (N_7040,N_461,N_3080);
nand U7041 (N_7041,N_994,N_182);
nor U7042 (N_7042,N_2407,N_3330);
nor U7043 (N_7043,N_1975,N_2116);
xor U7044 (N_7044,N_3368,N_2530);
or U7045 (N_7045,N_1016,N_2058);
and U7046 (N_7046,N_645,N_2846);
nor U7047 (N_7047,N_537,N_1933);
and U7048 (N_7048,N_1199,N_3788);
and U7049 (N_7049,N_59,N_1031);
or U7050 (N_7050,N_1953,N_3492);
nor U7051 (N_7051,N_607,N_2446);
xnor U7052 (N_7052,N_3991,N_367);
or U7053 (N_7053,N_525,N_79);
or U7054 (N_7054,N_1520,N_3220);
nand U7055 (N_7055,N_1870,N_2344);
nor U7056 (N_7056,N_3976,N_3199);
nor U7057 (N_7057,N_2065,N_1268);
and U7058 (N_7058,N_2586,N_3463);
xor U7059 (N_7059,N_1533,N_279);
nor U7060 (N_7060,N_1114,N_3569);
or U7061 (N_7061,N_2696,N_3503);
xor U7062 (N_7062,N_308,N_24);
and U7063 (N_7063,N_378,N_893);
xor U7064 (N_7064,N_1730,N_1223);
and U7065 (N_7065,N_2100,N_956);
or U7066 (N_7066,N_1417,N_622);
nand U7067 (N_7067,N_1265,N_725);
xor U7068 (N_7068,N_3741,N_3496);
nand U7069 (N_7069,N_3524,N_2107);
nand U7070 (N_7070,N_3566,N_2040);
nor U7071 (N_7071,N_2452,N_784);
nor U7072 (N_7072,N_1909,N_788);
and U7073 (N_7073,N_276,N_2502);
nor U7074 (N_7074,N_2329,N_3599);
and U7075 (N_7075,N_3636,N_951);
nor U7076 (N_7076,N_2027,N_3708);
nand U7077 (N_7077,N_388,N_3249);
and U7078 (N_7078,N_1943,N_3501);
or U7079 (N_7079,N_2689,N_3663);
nor U7080 (N_7080,N_2223,N_3390);
and U7081 (N_7081,N_620,N_1888);
nand U7082 (N_7082,N_1036,N_154);
xor U7083 (N_7083,N_1094,N_2205);
nor U7084 (N_7084,N_1479,N_3410);
nor U7085 (N_7085,N_2946,N_267);
nand U7086 (N_7086,N_564,N_1955);
xnor U7087 (N_7087,N_3440,N_3228);
nand U7088 (N_7088,N_1986,N_2800);
nand U7089 (N_7089,N_3747,N_1026);
and U7090 (N_7090,N_3036,N_3002);
nor U7091 (N_7091,N_3474,N_1323);
and U7092 (N_7092,N_1850,N_2774);
xnor U7093 (N_7093,N_574,N_2699);
nand U7094 (N_7094,N_266,N_3532);
or U7095 (N_7095,N_3851,N_2025);
nand U7096 (N_7096,N_3012,N_2301);
nor U7097 (N_7097,N_1954,N_3458);
xnor U7098 (N_7098,N_749,N_1224);
or U7099 (N_7099,N_2885,N_977);
or U7100 (N_7100,N_2911,N_2804);
and U7101 (N_7101,N_167,N_3984);
nand U7102 (N_7102,N_1218,N_3314);
xor U7103 (N_7103,N_1916,N_3939);
and U7104 (N_7104,N_1298,N_3663);
nor U7105 (N_7105,N_929,N_3276);
xnor U7106 (N_7106,N_797,N_1668);
nand U7107 (N_7107,N_1508,N_2401);
and U7108 (N_7108,N_1308,N_255);
xor U7109 (N_7109,N_522,N_3796);
nand U7110 (N_7110,N_403,N_1735);
nor U7111 (N_7111,N_2836,N_1201);
nand U7112 (N_7112,N_453,N_1814);
nor U7113 (N_7113,N_2742,N_3304);
and U7114 (N_7114,N_2131,N_702);
nand U7115 (N_7115,N_2657,N_3643);
or U7116 (N_7116,N_3570,N_3042);
and U7117 (N_7117,N_2574,N_1415);
nor U7118 (N_7118,N_2975,N_1941);
xnor U7119 (N_7119,N_2832,N_1356);
and U7120 (N_7120,N_770,N_1499);
nand U7121 (N_7121,N_358,N_3337);
nand U7122 (N_7122,N_1905,N_2075);
and U7123 (N_7123,N_325,N_613);
and U7124 (N_7124,N_539,N_837);
nor U7125 (N_7125,N_993,N_138);
nand U7126 (N_7126,N_2833,N_351);
nor U7127 (N_7127,N_3786,N_2520);
nand U7128 (N_7128,N_3651,N_2679);
and U7129 (N_7129,N_188,N_2055);
nand U7130 (N_7130,N_1970,N_215);
nand U7131 (N_7131,N_3076,N_3315);
nand U7132 (N_7132,N_828,N_39);
xnor U7133 (N_7133,N_3077,N_388);
nand U7134 (N_7134,N_36,N_3449);
nor U7135 (N_7135,N_2992,N_2184);
nor U7136 (N_7136,N_36,N_854);
xor U7137 (N_7137,N_173,N_832);
or U7138 (N_7138,N_3745,N_2564);
xnor U7139 (N_7139,N_1236,N_3034);
or U7140 (N_7140,N_923,N_3389);
xor U7141 (N_7141,N_635,N_238);
nor U7142 (N_7142,N_2941,N_384);
and U7143 (N_7143,N_3701,N_1315);
and U7144 (N_7144,N_770,N_26);
and U7145 (N_7145,N_1120,N_1235);
nor U7146 (N_7146,N_737,N_2993);
xor U7147 (N_7147,N_576,N_3080);
nand U7148 (N_7148,N_1378,N_3844);
and U7149 (N_7149,N_1820,N_1944);
and U7150 (N_7150,N_1321,N_881);
xor U7151 (N_7151,N_2950,N_3489);
and U7152 (N_7152,N_765,N_3887);
or U7153 (N_7153,N_422,N_2944);
and U7154 (N_7154,N_1675,N_226);
xnor U7155 (N_7155,N_666,N_1413);
xor U7156 (N_7156,N_422,N_2875);
nand U7157 (N_7157,N_1607,N_1485);
xnor U7158 (N_7158,N_1105,N_1165);
and U7159 (N_7159,N_791,N_2424);
nor U7160 (N_7160,N_1815,N_1863);
nor U7161 (N_7161,N_1612,N_1093);
and U7162 (N_7162,N_3062,N_2125);
nand U7163 (N_7163,N_2370,N_404);
or U7164 (N_7164,N_1418,N_2260);
nor U7165 (N_7165,N_1184,N_1593);
and U7166 (N_7166,N_3440,N_3794);
nand U7167 (N_7167,N_551,N_3484);
nand U7168 (N_7168,N_52,N_2860);
xor U7169 (N_7169,N_400,N_1631);
xnor U7170 (N_7170,N_1448,N_2065);
xor U7171 (N_7171,N_305,N_3075);
and U7172 (N_7172,N_3247,N_3154);
and U7173 (N_7173,N_1365,N_1910);
or U7174 (N_7174,N_3510,N_3911);
xor U7175 (N_7175,N_1598,N_3906);
xnor U7176 (N_7176,N_846,N_1748);
nor U7177 (N_7177,N_1061,N_2234);
nor U7178 (N_7178,N_3005,N_2166);
or U7179 (N_7179,N_910,N_1030);
and U7180 (N_7180,N_865,N_1267);
or U7181 (N_7181,N_2209,N_2616);
nor U7182 (N_7182,N_1928,N_2712);
xnor U7183 (N_7183,N_2888,N_1901);
nor U7184 (N_7184,N_2239,N_1535);
xor U7185 (N_7185,N_1421,N_3793);
or U7186 (N_7186,N_1268,N_2053);
or U7187 (N_7187,N_3969,N_68);
xor U7188 (N_7188,N_3531,N_1514);
nand U7189 (N_7189,N_2591,N_1087);
or U7190 (N_7190,N_129,N_931);
xnor U7191 (N_7191,N_2301,N_2895);
or U7192 (N_7192,N_787,N_924);
and U7193 (N_7193,N_2552,N_577);
or U7194 (N_7194,N_98,N_1521);
nor U7195 (N_7195,N_3113,N_2546);
nor U7196 (N_7196,N_3737,N_750);
nor U7197 (N_7197,N_107,N_2555);
or U7198 (N_7198,N_1717,N_970);
nor U7199 (N_7199,N_3900,N_3115);
nor U7200 (N_7200,N_1860,N_3635);
nand U7201 (N_7201,N_2238,N_2281);
or U7202 (N_7202,N_192,N_659);
nor U7203 (N_7203,N_2909,N_3946);
and U7204 (N_7204,N_3230,N_3600);
and U7205 (N_7205,N_3515,N_2894);
xnor U7206 (N_7206,N_3617,N_306);
xnor U7207 (N_7207,N_1031,N_1751);
nor U7208 (N_7208,N_1591,N_1982);
and U7209 (N_7209,N_414,N_1390);
nand U7210 (N_7210,N_3183,N_974);
nor U7211 (N_7211,N_465,N_268);
and U7212 (N_7212,N_1019,N_2210);
nor U7213 (N_7213,N_2115,N_3463);
and U7214 (N_7214,N_1393,N_2089);
and U7215 (N_7215,N_1592,N_2350);
nor U7216 (N_7216,N_724,N_2232);
or U7217 (N_7217,N_2950,N_2529);
or U7218 (N_7218,N_3255,N_759);
or U7219 (N_7219,N_949,N_3080);
or U7220 (N_7220,N_123,N_3647);
or U7221 (N_7221,N_1563,N_2609);
xor U7222 (N_7222,N_1972,N_3444);
nand U7223 (N_7223,N_8,N_2092);
xnor U7224 (N_7224,N_347,N_1487);
nand U7225 (N_7225,N_3724,N_2696);
and U7226 (N_7226,N_33,N_98);
or U7227 (N_7227,N_1780,N_3881);
or U7228 (N_7228,N_291,N_3628);
nor U7229 (N_7229,N_635,N_652);
xor U7230 (N_7230,N_3247,N_1095);
xnor U7231 (N_7231,N_2552,N_2455);
xnor U7232 (N_7232,N_3477,N_3985);
and U7233 (N_7233,N_1402,N_1358);
and U7234 (N_7234,N_0,N_1473);
xnor U7235 (N_7235,N_2661,N_3843);
xor U7236 (N_7236,N_309,N_2613);
nand U7237 (N_7237,N_459,N_879);
and U7238 (N_7238,N_2288,N_557);
nand U7239 (N_7239,N_1450,N_3678);
nor U7240 (N_7240,N_2948,N_3119);
nor U7241 (N_7241,N_3510,N_1505);
and U7242 (N_7242,N_1316,N_2411);
xnor U7243 (N_7243,N_3918,N_3163);
nor U7244 (N_7244,N_2491,N_3768);
xor U7245 (N_7245,N_439,N_1759);
or U7246 (N_7246,N_1728,N_2795);
or U7247 (N_7247,N_2485,N_1437);
nor U7248 (N_7248,N_83,N_959);
xnor U7249 (N_7249,N_3754,N_3564);
nand U7250 (N_7250,N_2570,N_3895);
and U7251 (N_7251,N_833,N_2659);
xnor U7252 (N_7252,N_2811,N_24);
and U7253 (N_7253,N_3382,N_2688);
nor U7254 (N_7254,N_2083,N_506);
xnor U7255 (N_7255,N_127,N_2939);
and U7256 (N_7256,N_2184,N_3100);
nor U7257 (N_7257,N_2051,N_518);
and U7258 (N_7258,N_1798,N_3475);
nand U7259 (N_7259,N_940,N_3352);
nor U7260 (N_7260,N_1224,N_2803);
xor U7261 (N_7261,N_3702,N_885);
nor U7262 (N_7262,N_3576,N_2127);
nand U7263 (N_7263,N_3201,N_2383);
and U7264 (N_7264,N_1124,N_3102);
or U7265 (N_7265,N_3026,N_2344);
or U7266 (N_7266,N_3976,N_192);
nand U7267 (N_7267,N_3846,N_2500);
and U7268 (N_7268,N_3261,N_1420);
or U7269 (N_7269,N_3441,N_2159);
or U7270 (N_7270,N_3797,N_3046);
nand U7271 (N_7271,N_3887,N_2287);
xnor U7272 (N_7272,N_754,N_1653);
nand U7273 (N_7273,N_3548,N_3152);
or U7274 (N_7274,N_1156,N_562);
and U7275 (N_7275,N_2236,N_2996);
xnor U7276 (N_7276,N_2932,N_2488);
xnor U7277 (N_7277,N_3142,N_583);
and U7278 (N_7278,N_3198,N_3296);
nand U7279 (N_7279,N_3693,N_1462);
nand U7280 (N_7280,N_1053,N_2544);
and U7281 (N_7281,N_3031,N_2600);
nand U7282 (N_7282,N_1978,N_303);
and U7283 (N_7283,N_2895,N_2796);
or U7284 (N_7284,N_1898,N_2093);
nand U7285 (N_7285,N_3020,N_1851);
or U7286 (N_7286,N_227,N_1535);
xnor U7287 (N_7287,N_2995,N_1210);
and U7288 (N_7288,N_2703,N_2333);
nor U7289 (N_7289,N_2370,N_252);
nor U7290 (N_7290,N_1765,N_100);
xnor U7291 (N_7291,N_1922,N_739);
nor U7292 (N_7292,N_2375,N_1129);
and U7293 (N_7293,N_3467,N_2549);
or U7294 (N_7294,N_2012,N_3338);
and U7295 (N_7295,N_3132,N_2618);
xnor U7296 (N_7296,N_631,N_1401);
nor U7297 (N_7297,N_727,N_526);
or U7298 (N_7298,N_2156,N_2563);
nand U7299 (N_7299,N_342,N_3342);
nor U7300 (N_7300,N_627,N_3165);
or U7301 (N_7301,N_2303,N_3946);
nor U7302 (N_7302,N_3128,N_2698);
nor U7303 (N_7303,N_1275,N_2176);
and U7304 (N_7304,N_2954,N_2898);
nand U7305 (N_7305,N_286,N_2091);
xor U7306 (N_7306,N_1266,N_3253);
xnor U7307 (N_7307,N_2952,N_1679);
nand U7308 (N_7308,N_3575,N_1883);
nand U7309 (N_7309,N_1059,N_1359);
xnor U7310 (N_7310,N_256,N_2705);
nand U7311 (N_7311,N_300,N_1054);
nand U7312 (N_7312,N_3597,N_2751);
nand U7313 (N_7313,N_3644,N_615);
nand U7314 (N_7314,N_2897,N_2625);
nor U7315 (N_7315,N_2606,N_1150);
nand U7316 (N_7316,N_516,N_1789);
xnor U7317 (N_7317,N_614,N_789);
or U7318 (N_7318,N_1626,N_1274);
or U7319 (N_7319,N_520,N_2841);
and U7320 (N_7320,N_113,N_47);
xor U7321 (N_7321,N_701,N_3532);
nand U7322 (N_7322,N_490,N_3640);
xnor U7323 (N_7323,N_1624,N_1698);
nand U7324 (N_7324,N_3027,N_3037);
or U7325 (N_7325,N_3110,N_3676);
xnor U7326 (N_7326,N_923,N_2479);
nand U7327 (N_7327,N_3216,N_1518);
or U7328 (N_7328,N_1088,N_392);
nor U7329 (N_7329,N_678,N_2600);
nor U7330 (N_7330,N_1207,N_2335);
nand U7331 (N_7331,N_2816,N_3427);
xnor U7332 (N_7332,N_986,N_273);
and U7333 (N_7333,N_283,N_1948);
nor U7334 (N_7334,N_2542,N_1371);
xor U7335 (N_7335,N_1784,N_2154);
nand U7336 (N_7336,N_194,N_3304);
xnor U7337 (N_7337,N_665,N_663);
and U7338 (N_7338,N_3065,N_2819);
nand U7339 (N_7339,N_2967,N_1574);
and U7340 (N_7340,N_2449,N_1710);
and U7341 (N_7341,N_3354,N_786);
nor U7342 (N_7342,N_3473,N_942);
or U7343 (N_7343,N_500,N_780);
nor U7344 (N_7344,N_916,N_1439);
nor U7345 (N_7345,N_523,N_1653);
nand U7346 (N_7346,N_2853,N_2454);
or U7347 (N_7347,N_2315,N_1021);
or U7348 (N_7348,N_1075,N_3236);
or U7349 (N_7349,N_376,N_3966);
nor U7350 (N_7350,N_3787,N_486);
nand U7351 (N_7351,N_2769,N_2504);
or U7352 (N_7352,N_19,N_551);
nand U7353 (N_7353,N_2335,N_2688);
or U7354 (N_7354,N_3413,N_3108);
or U7355 (N_7355,N_1762,N_3426);
or U7356 (N_7356,N_1952,N_2545);
nor U7357 (N_7357,N_2389,N_505);
nand U7358 (N_7358,N_1172,N_2564);
nor U7359 (N_7359,N_1403,N_173);
nand U7360 (N_7360,N_3600,N_1774);
or U7361 (N_7361,N_2020,N_687);
nand U7362 (N_7362,N_2804,N_2592);
nand U7363 (N_7363,N_390,N_1005);
or U7364 (N_7364,N_1142,N_2850);
nor U7365 (N_7365,N_3878,N_3591);
nor U7366 (N_7366,N_1610,N_1877);
nor U7367 (N_7367,N_3014,N_1908);
or U7368 (N_7368,N_778,N_3872);
nor U7369 (N_7369,N_2508,N_1192);
and U7370 (N_7370,N_1584,N_1110);
nand U7371 (N_7371,N_3133,N_2739);
and U7372 (N_7372,N_3534,N_3110);
and U7373 (N_7373,N_3702,N_565);
and U7374 (N_7374,N_3165,N_3104);
or U7375 (N_7375,N_3648,N_2021);
xnor U7376 (N_7376,N_2889,N_1302);
and U7377 (N_7377,N_3557,N_1762);
or U7378 (N_7378,N_2988,N_3059);
nor U7379 (N_7379,N_3078,N_1870);
nand U7380 (N_7380,N_205,N_2346);
and U7381 (N_7381,N_1047,N_1350);
nand U7382 (N_7382,N_2091,N_1291);
xnor U7383 (N_7383,N_3353,N_1886);
nor U7384 (N_7384,N_1621,N_2471);
and U7385 (N_7385,N_3048,N_633);
xnor U7386 (N_7386,N_3949,N_70);
or U7387 (N_7387,N_1029,N_3191);
nor U7388 (N_7388,N_1932,N_1939);
nor U7389 (N_7389,N_2611,N_2485);
nand U7390 (N_7390,N_2878,N_1488);
xor U7391 (N_7391,N_2905,N_2287);
nand U7392 (N_7392,N_1445,N_2915);
xor U7393 (N_7393,N_2359,N_1248);
and U7394 (N_7394,N_2253,N_3858);
xor U7395 (N_7395,N_2920,N_3645);
and U7396 (N_7396,N_814,N_3536);
nor U7397 (N_7397,N_246,N_3487);
nor U7398 (N_7398,N_365,N_3455);
nand U7399 (N_7399,N_2025,N_967);
and U7400 (N_7400,N_1414,N_740);
and U7401 (N_7401,N_1466,N_3156);
or U7402 (N_7402,N_1116,N_654);
nand U7403 (N_7403,N_1535,N_1739);
nand U7404 (N_7404,N_3270,N_1200);
nand U7405 (N_7405,N_3234,N_48);
xor U7406 (N_7406,N_2966,N_243);
nand U7407 (N_7407,N_252,N_359);
or U7408 (N_7408,N_2313,N_3677);
xor U7409 (N_7409,N_106,N_450);
nor U7410 (N_7410,N_3248,N_1510);
nor U7411 (N_7411,N_2136,N_2636);
nor U7412 (N_7412,N_3258,N_504);
xor U7413 (N_7413,N_2561,N_1091);
nand U7414 (N_7414,N_1076,N_1734);
and U7415 (N_7415,N_2135,N_3722);
and U7416 (N_7416,N_2237,N_3784);
or U7417 (N_7417,N_311,N_2570);
and U7418 (N_7418,N_3361,N_1828);
xnor U7419 (N_7419,N_1333,N_2479);
nand U7420 (N_7420,N_801,N_3651);
nor U7421 (N_7421,N_634,N_3075);
nor U7422 (N_7422,N_788,N_3582);
and U7423 (N_7423,N_1448,N_343);
and U7424 (N_7424,N_2981,N_3450);
or U7425 (N_7425,N_3909,N_1036);
and U7426 (N_7426,N_1789,N_2400);
and U7427 (N_7427,N_1808,N_3359);
nand U7428 (N_7428,N_2641,N_1571);
xnor U7429 (N_7429,N_1137,N_2422);
xor U7430 (N_7430,N_1653,N_2535);
nor U7431 (N_7431,N_3367,N_924);
and U7432 (N_7432,N_3655,N_3233);
nor U7433 (N_7433,N_2702,N_3950);
or U7434 (N_7434,N_2238,N_3193);
and U7435 (N_7435,N_2755,N_3792);
nand U7436 (N_7436,N_1390,N_1524);
nor U7437 (N_7437,N_1209,N_1604);
and U7438 (N_7438,N_1076,N_3311);
or U7439 (N_7439,N_2454,N_2419);
nor U7440 (N_7440,N_3663,N_780);
nor U7441 (N_7441,N_234,N_685);
nand U7442 (N_7442,N_153,N_2463);
nand U7443 (N_7443,N_1074,N_2242);
and U7444 (N_7444,N_3689,N_1429);
xor U7445 (N_7445,N_314,N_3178);
xor U7446 (N_7446,N_2708,N_1355);
nand U7447 (N_7447,N_3428,N_2633);
or U7448 (N_7448,N_3102,N_707);
nand U7449 (N_7449,N_3025,N_3169);
and U7450 (N_7450,N_2425,N_453);
nand U7451 (N_7451,N_2603,N_2123);
nand U7452 (N_7452,N_294,N_3946);
xor U7453 (N_7453,N_991,N_2076);
nand U7454 (N_7454,N_3462,N_544);
xnor U7455 (N_7455,N_1741,N_1312);
nor U7456 (N_7456,N_3674,N_393);
or U7457 (N_7457,N_3009,N_913);
nand U7458 (N_7458,N_3650,N_416);
nor U7459 (N_7459,N_3556,N_2950);
or U7460 (N_7460,N_1377,N_508);
and U7461 (N_7461,N_2820,N_3571);
nor U7462 (N_7462,N_2253,N_731);
nand U7463 (N_7463,N_3887,N_1575);
xor U7464 (N_7464,N_2308,N_248);
and U7465 (N_7465,N_3951,N_811);
nor U7466 (N_7466,N_1554,N_3452);
or U7467 (N_7467,N_2752,N_1472);
or U7468 (N_7468,N_3067,N_2331);
nor U7469 (N_7469,N_1020,N_3730);
or U7470 (N_7470,N_935,N_3756);
nand U7471 (N_7471,N_896,N_569);
xor U7472 (N_7472,N_2365,N_1492);
nor U7473 (N_7473,N_1016,N_3574);
and U7474 (N_7474,N_450,N_3651);
nor U7475 (N_7475,N_3663,N_2695);
nand U7476 (N_7476,N_3433,N_3224);
nand U7477 (N_7477,N_2155,N_259);
xnor U7478 (N_7478,N_2507,N_3862);
nor U7479 (N_7479,N_3016,N_2964);
nor U7480 (N_7480,N_3626,N_63);
nor U7481 (N_7481,N_1442,N_982);
or U7482 (N_7482,N_577,N_1185);
nand U7483 (N_7483,N_3370,N_2425);
nor U7484 (N_7484,N_1971,N_2255);
xnor U7485 (N_7485,N_3523,N_219);
nand U7486 (N_7486,N_1682,N_1881);
xnor U7487 (N_7487,N_2730,N_3742);
nor U7488 (N_7488,N_2242,N_1342);
nor U7489 (N_7489,N_372,N_233);
xor U7490 (N_7490,N_451,N_697);
nor U7491 (N_7491,N_2520,N_2260);
nand U7492 (N_7492,N_455,N_826);
and U7493 (N_7493,N_650,N_3151);
nand U7494 (N_7494,N_3632,N_719);
xnor U7495 (N_7495,N_2430,N_2606);
or U7496 (N_7496,N_2428,N_1602);
and U7497 (N_7497,N_2349,N_1317);
and U7498 (N_7498,N_3765,N_1157);
and U7499 (N_7499,N_2152,N_2877);
nand U7500 (N_7500,N_1314,N_32);
nor U7501 (N_7501,N_2939,N_2925);
nand U7502 (N_7502,N_663,N_1286);
and U7503 (N_7503,N_3804,N_2286);
or U7504 (N_7504,N_3200,N_1744);
and U7505 (N_7505,N_45,N_3061);
xor U7506 (N_7506,N_2817,N_2965);
and U7507 (N_7507,N_1956,N_2241);
xor U7508 (N_7508,N_2005,N_2375);
nand U7509 (N_7509,N_3219,N_424);
nor U7510 (N_7510,N_3810,N_3225);
nand U7511 (N_7511,N_1153,N_2400);
nor U7512 (N_7512,N_1529,N_913);
xor U7513 (N_7513,N_594,N_1079);
nor U7514 (N_7514,N_1917,N_1782);
nor U7515 (N_7515,N_2062,N_1824);
or U7516 (N_7516,N_3608,N_1388);
nor U7517 (N_7517,N_2515,N_529);
and U7518 (N_7518,N_2344,N_2556);
nor U7519 (N_7519,N_1584,N_2162);
or U7520 (N_7520,N_2174,N_1931);
nor U7521 (N_7521,N_3806,N_217);
and U7522 (N_7522,N_2860,N_3345);
xnor U7523 (N_7523,N_1181,N_969);
nor U7524 (N_7524,N_3758,N_2749);
or U7525 (N_7525,N_3554,N_1188);
or U7526 (N_7526,N_1886,N_2366);
nand U7527 (N_7527,N_2291,N_624);
nor U7528 (N_7528,N_2781,N_2365);
nor U7529 (N_7529,N_3727,N_487);
nor U7530 (N_7530,N_1314,N_3195);
nor U7531 (N_7531,N_2945,N_765);
nor U7532 (N_7532,N_3104,N_658);
or U7533 (N_7533,N_227,N_1797);
nand U7534 (N_7534,N_1286,N_2405);
or U7535 (N_7535,N_3991,N_140);
nand U7536 (N_7536,N_5,N_3396);
nand U7537 (N_7537,N_1756,N_1039);
or U7538 (N_7538,N_2951,N_3013);
nand U7539 (N_7539,N_1936,N_3685);
nand U7540 (N_7540,N_1488,N_641);
xor U7541 (N_7541,N_3802,N_1168);
nor U7542 (N_7542,N_3637,N_667);
xor U7543 (N_7543,N_2995,N_2615);
nor U7544 (N_7544,N_3464,N_3845);
xnor U7545 (N_7545,N_496,N_3227);
xor U7546 (N_7546,N_1105,N_1139);
xor U7547 (N_7547,N_1906,N_1397);
and U7548 (N_7548,N_990,N_431);
or U7549 (N_7549,N_2448,N_1309);
xor U7550 (N_7550,N_1294,N_1986);
or U7551 (N_7551,N_3360,N_727);
or U7552 (N_7552,N_3752,N_2034);
or U7553 (N_7553,N_864,N_578);
xnor U7554 (N_7554,N_204,N_715);
and U7555 (N_7555,N_2422,N_358);
or U7556 (N_7556,N_3056,N_293);
or U7557 (N_7557,N_1158,N_2754);
or U7558 (N_7558,N_1464,N_1065);
nor U7559 (N_7559,N_1791,N_1628);
or U7560 (N_7560,N_2520,N_3034);
and U7561 (N_7561,N_458,N_1663);
or U7562 (N_7562,N_395,N_209);
nor U7563 (N_7563,N_1474,N_268);
nor U7564 (N_7564,N_1404,N_1117);
xnor U7565 (N_7565,N_2436,N_142);
nor U7566 (N_7566,N_26,N_909);
nand U7567 (N_7567,N_71,N_2816);
nor U7568 (N_7568,N_1133,N_3763);
and U7569 (N_7569,N_1977,N_1206);
xnor U7570 (N_7570,N_2871,N_2972);
and U7571 (N_7571,N_2413,N_1534);
nor U7572 (N_7572,N_2452,N_314);
xnor U7573 (N_7573,N_1736,N_2381);
or U7574 (N_7574,N_49,N_154);
nor U7575 (N_7575,N_2900,N_2770);
nor U7576 (N_7576,N_1455,N_3244);
nand U7577 (N_7577,N_609,N_1809);
nor U7578 (N_7578,N_3083,N_2262);
and U7579 (N_7579,N_1792,N_1117);
or U7580 (N_7580,N_1602,N_1687);
nand U7581 (N_7581,N_3048,N_3103);
nor U7582 (N_7582,N_1248,N_3196);
xnor U7583 (N_7583,N_962,N_2488);
nor U7584 (N_7584,N_1578,N_2113);
xor U7585 (N_7585,N_2267,N_2091);
nand U7586 (N_7586,N_1888,N_3254);
xor U7587 (N_7587,N_3081,N_1956);
or U7588 (N_7588,N_2858,N_111);
nor U7589 (N_7589,N_472,N_744);
or U7590 (N_7590,N_884,N_2005);
or U7591 (N_7591,N_1424,N_3042);
or U7592 (N_7592,N_260,N_948);
xnor U7593 (N_7593,N_1339,N_959);
xor U7594 (N_7594,N_3744,N_2151);
and U7595 (N_7595,N_2877,N_2869);
or U7596 (N_7596,N_1572,N_2379);
xor U7597 (N_7597,N_2501,N_159);
or U7598 (N_7598,N_2027,N_2921);
and U7599 (N_7599,N_3306,N_621);
and U7600 (N_7600,N_3093,N_441);
xor U7601 (N_7601,N_3810,N_948);
nand U7602 (N_7602,N_2630,N_3845);
nor U7603 (N_7603,N_2086,N_3238);
nor U7604 (N_7604,N_3465,N_202);
nor U7605 (N_7605,N_3601,N_3284);
nand U7606 (N_7606,N_3775,N_1103);
xor U7607 (N_7607,N_2302,N_395);
or U7608 (N_7608,N_190,N_323);
and U7609 (N_7609,N_1433,N_1302);
nor U7610 (N_7610,N_353,N_115);
nand U7611 (N_7611,N_2743,N_2477);
xnor U7612 (N_7612,N_3689,N_1362);
or U7613 (N_7613,N_2350,N_1363);
xnor U7614 (N_7614,N_3531,N_2206);
or U7615 (N_7615,N_3859,N_3773);
and U7616 (N_7616,N_2993,N_3650);
nor U7617 (N_7617,N_1649,N_3233);
nor U7618 (N_7618,N_3231,N_203);
nor U7619 (N_7619,N_1112,N_3386);
nor U7620 (N_7620,N_2522,N_1365);
or U7621 (N_7621,N_279,N_1990);
or U7622 (N_7622,N_1592,N_1604);
nor U7623 (N_7623,N_2501,N_693);
xor U7624 (N_7624,N_1456,N_3926);
or U7625 (N_7625,N_2846,N_3531);
nand U7626 (N_7626,N_2796,N_1130);
nand U7627 (N_7627,N_920,N_213);
nor U7628 (N_7628,N_781,N_3027);
nand U7629 (N_7629,N_3755,N_3221);
nor U7630 (N_7630,N_1822,N_1317);
or U7631 (N_7631,N_2568,N_2514);
or U7632 (N_7632,N_2719,N_3562);
or U7633 (N_7633,N_2597,N_89);
nand U7634 (N_7634,N_577,N_220);
or U7635 (N_7635,N_32,N_313);
or U7636 (N_7636,N_302,N_909);
nor U7637 (N_7637,N_1119,N_1164);
xor U7638 (N_7638,N_3403,N_2921);
nand U7639 (N_7639,N_3033,N_2058);
or U7640 (N_7640,N_3842,N_3485);
nand U7641 (N_7641,N_1950,N_1615);
xor U7642 (N_7642,N_3340,N_2145);
and U7643 (N_7643,N_2632,N_1406);
nand U7644 (N_7644,N_983,N_347);
and U7645 (N_7645,N_2149,N_785);
and U7646 (N_7646,N_198,N_684);
and U7647 (N_7647,N_1467,N_2591);
nor U7648 (N_7648,N_2966,N_2940);
or U7649 (N_7649,N_1378,N_1212);
nor U7650 (N_7650,N_236,N_1697);
and U7651 (N_7651,N_2705,N_487);
or U7652 (N_7652,N_793,N_1822);
nand U7653 (N_7653,N_804,N_1554);
nand U7654 (N_7654,N_3244,N_3493);
or U7655 (N_7655,N_3483,N_3316);
or U7656 (N_7656,N_591,N_3000);
nand U7657 (N_7657,N_3970,N_627);
and U7658 (N_7658,N_2277,N_3142);
nor U7659 (N_7659,N_2420,N_159);
nor U7660 (N_7660,N_428,N_1847);
nand U7661 (N_7661,N_1304,N_1342);
xnor U7662 (N_7662,N_3957,N_357);
nor U7663 (N_7663,N_3280,N_3550);
or U7664 (N_7664,N_1667,N_3653);
nand U7665 (N_7665,N_2482,N_547);
nor U7666 (N_7666,N_3877,N_2812);
and U7667 (N_7667,N_2973,N_2503);
nor U7668 (N_7668,N_1349,N_644);
nand U7669 (N_7669,N_2722,N_270);
nor U7670 (N_7670,N_2662,N_1768);
xnor U7671 (N_7671,N_2504,N_3102);
and U7672 (N_7672,N_818,N_3551);
or U7673 (N_7673,N_864,N_1748);
xnor U7674 (N_7674,N_2515,N_1007);
and U7675 (N_7675,N_2318,N_1268);
nand U7676 (N_7676,N_2222,N_1048);
and U7677 (N_7677,N_2627,N_1799);
and U7678 (N_7678,N_1420,N_1558);
xnor U7679 (N_7679,N_344,N_1825);
nor U7680 (N_7680,N_3953,N_407);
nand U7681 (N_7681,N_314,N_765);
xor U7682 (N_7682,N_2970,N_1131);
nand U7683 (N_7683,N_1383,N_3768);
and U7684 (N_7684,N_1537,N_199);
or U7685 (N_7685,N_659,N_1464);
and U7686 (N_7686,N_2985,N_3795);
xnor U7687 (N_7687,N_1082,N_1534);
nand U7688 (N_7688,N_615,N_3971);
nand U7689 (N_7689,N_315,N_791);
and U7690 (N_7690,N_995,N_1593);
and U7691 (N_7691,N_3056,N_1357);
and U7692 (N_7692,N_289,N_2813);
or U7693 (N_7693,N_8,N_3035);
and U7694 (N_7694,N_375,N_2545);
and U7695 (N_7695,N_1361,N_683);
xor U7696 (N_7696,N_2880,N_390);
and U7697 (N_7697,N_3861,N_842);
nand U7698 (N_7698,N_2005,N_3997);
nand U7699 (N_7699,N_3175,N_2015);
nor U7700 (N_7700,N_324,N_508);
xnor U7701 (N_7701,N_1403,N_1002);
nand U7702 (N_7702,N_2673,N_1345);
and U7703 (N_7703,N_526,N_71);
and U7704 (N_7704,N_876,N_1312);
or U7705 (N_7705,N_321,N_3475);
or U7706 (N_7706,N_574,N_1051);
and U7707 (N_7707,N_1318,N_611);
xnor U7708 (N_7708,N_325,N_3033);
or U7709 (N_7709,N_3082,N_3667);
nor U7710 (N_7710,N_2129,N_3542);
nand U7711 (N_7711,N_620,N_153);
nand U7712 (N_7712,N_2575,N_697);
and U7713 (N_7713,N_3132,N_2935);
or U7714 (N_7714,N_1555,N_2481);
and U7715 (N_7715,N_2048,N_902);
nor U7716 (N_7716,N_3923,N_3818);
or U7717 (N_7717,N_203,N_3869);
or U7718 (N_7718,N_3989,N_2696);
and U7719 (N_7719,N_350,N_574);
and U7720 (N_7720,N_1005,N_111);
nor U7721 (N_7721,N_1248,N_2916);
nor U7722 (N_7722,N_2294,N_1173);
and U7723 (N_7723,N_1090,N_1049);
nand U7724 (N_7724,N_194,N_2776);
or U7725 (N_7725,N_3099,N_2685);
nand U7726 (N_7726,N_930,N_3890);
or U7727 (N_7727,N_2991,N_828);
xor U7728 (N_7728,N_2245,N_3397);
xor U7729 (N_7729,N_2353,N_993);
nor U7730 (N_7730,N_882,N_2182);
or U7731 (N_7731,N_3769,N_2193);
or U7732 (N_7732,N_2811,N_2930);
xnor U7733 (N_7733,N_2269,N_2550);
xnor U7734 (N_7734,N_3414,N_3429);
nand U7735 (N_7735,N_1036,N_46);
nor U7736 (N_7736,N_657,N_2936);
nor U7737 (N_7737,N_2477,N_2822);
nand U7738 (N_7738,N_1974,N_2963);
or U7739 (N_7739,N_3085,N_2189);
nand U7740 (N_7740,N_2874,N_1782);
nand U7741 (N_7741,N_469,N_3036);
nand U7742 (N_7742,N_448,N_3446);
xnor U7743 (N_7743,N_3948,N_510);
or U7744 (N_7744,N_3068,N_3992);
nand U7745 (N_7745,N_437,N_906);
nor U7746 (N_7746,N_1975,N_11);
and U7747 (N_7747,N_3320,N_1769);
nor U7748 (N_7748,N_2263,N_2926);
and U7749 (N_7749,N_1480,N_916);
nand U7750 (N_7750,N_1419,N_2986);
and U7751 (N_7751,N_3614,N_290);
and U7752 (N_7752,N_215,N_3137);
or U7753 (N_7753,N_2714,N_3305);
xor U7754 (N_7754,N_3646,N_1000);
and U7755 (N_7755,N_2172,N_2904);
and U7756 (N_7756,N_2224,N_3999);
nand U7757 (N_7757,N_3273,N_310);
xor U7758 (N_7758,N_367,N_2615);
nor U7759 (N_7759,N_697,N_1169);
nor U7760 (N_7760,N_2409,N_1929);
or U7761 (N_7761,N_3835,N_1048);
and U7762 (N_7762,N_3791,N_875);
or U7763 (N_7763,N_1113,N_63);
nand U7764 (N_7764,N_3867,N_2659);
nand U7765 (N_7765,N_1650,N_2332);
or U7766 (N_7766,N_1972,N_3596);
xor U7767 (N_7767,N_2549,N_250);
xnor U7768 (N_7768,N_567,N_2791);
or U7769 (N_7769,N_1131,N_384);
nand U7770 (N_7770,N_413,N_2391);
xor U7771 (N_7771,N_2689,N_2);
nand U7772 (N_7772,N_1338,N_3140);
or U7773 (N_7773,N_2969,N_845);
and U7774 (N_7774,N_3232,N_1296);
or U7775 (N_7775,N_2018,N_1207);
or U7776 (N_7776,N_398,N_1765);
xnor U7777 (N_7777,N_188,N_2018);
xnor U7778 (N_7778,N_3491,N_902);
and U7779 (N_7779,N_2673,N_1333);
nor U7780 (N_7780,N_266,N_1669);
and U7781 (N_7781,N_3850,N_2678);
xnor U7782 (N_7782,N_2,N_3956);
nand U7783 (N_7783,N_3608,N_1358);
nor U7784 (N_7784,N_1879,N_18);
xor U7785 (N_7785,N_2723,N_486);
or U7786 (N_7786,N_3550,N_1568);
nand U7787 (N_7787,N_2604,N_2725);
and U7788 (N_7788,N_2142,N_902);
and U7789 (N_7789,N_3736,N_3695);
nor U7790 (N_7790,N_2359,N_2882);
nor U7791 (N_7791,N_138,N_552);
nor U7792 (N_7792,N_1938,N_3011);
nand U7793 (N_7793,N_3437,N_1305);
nor U7794 (N_7794,N_3675,N_3915);
or U7795 (N_7795,N_3956,N_1237);
and U7796 (N_7796,N_100,N_19);
nand U7797 (N_7797,N_3967,N_3211);
nor U7798 (N_7798,N_1797,N_91);
xor U7799 (N_7799,N_112,N_2924);
nand U7800 (N_7800,N_2204,N_2350);
xor U7801 (N_7801,N_2674,N_2822);
nand U7802 (N_7802,N_2790,N_3748);
and U7803 (N_7803,N_1729,N_688);
xor U7804 (N_7804,N_440,N_74);
nand U7805 (N_7805,N_2118,N_2784);
nand U7806 (N_7806,N_1926,N_274);
or U7807 (N_7807,N_2741,N_1308);
nor U7808 (N_7808,N_682,N_3498);
nand U7809 (N_7809,N_204,N_1934);
nand U7810 (N_7810,N_3878,N_1783);
or U7811 (N_7811,N_2148,N_3139);
or U7812 (N_7812,N_1072,N_3107);
nor U7813 (N_7813,N_316,N_3389);
xor U7814 (N_7814,N_535,N_3468);
nor U7815 (N_7815,N_184,N_56);
nor U7816 (N_7816,N_3405,N_916);
xor U7817 (N_7817,N_198,N_1158);
nand U7818 (N_7818,N_1960,N_128);
and U7819 (N_7819,N_2274,N_1896);
nand U7820 (N_7820,N_3574,N_3107);
nor U7821 (N_7821,N_634,N_3406);
nand U7822 (N_7822,N_2949,N_3535);
nand U7823 (N_7823,N_3392,N_3579);
nor U7824 (N_7824,N_1531,N_2784);
nand U7825 (N_7825,N_3060,N_234);
nor U7826 (N_7826,N_223,N_794);
nand U7827 (N_7827,N_1432,N_649);
nor U7828 (N_7828,N_2849,N_449);
or U7829 (N_7829,N_2608,N_3989);
nor U7830 (N_7830,N_2442,N_2995);
or U7831 (N_7831,N_3289,N_324);
and U7832 (N_7832,N_3645,N_184);
and U7833 (N_7833,N_1814,N_3706);
nand U7834 (N_7834,N_1533,N_3276);
or U7835 (N_7835,N_2345,N_3088);
nor U7836 (N_7836,N_1166,N_2437);
and U7837 (N_7837,N_974,N_1144);
xor U7838 (N_7838,N_3067,N_1561);
nor U7839 (N_7839,N_1539,N_3053);
nand U7840 (N_7840,N_3642,N_156);
xor U7841 (N_7841,N_2435,N_3932);
or U7842 (N_7842,N_2016,N_1125);
or U7843 (N_7843,N_3835,N_1026);
nand U7844 (N_7844,N_1752,N_1580);
xor U7845 (N_7845,N_3732,N_3173);
xor U7846 (N_7846,N_166,N_3862);
nand U7847 (N_7847,N_2507,N_234);
nor U7848 (N_7848,N_2521,N_3698);
xnor U7849 (N_7849,N_780,N_3472);
xor U7850 (N_7850,N_3557,N_1967);
and U7851 (N_7851,N_3823,N_1260);
and U7852 (N_7852,N_1358,N_1019);
nor U7853 (N_7853,N_2247,N_3671);
nor U7854 (N_7854,N_2483,N_1973);
nand U7855 (N_7855,N_3293,N_2193);
or U7856 (N_7856,N_26,N_2832);
xor U7857 (N_7857,N_3761,N_3376);
and U7858 (N_7858,N_2158,N_2315);
nor U7859 (N_7859,N_643,N_850);
nor U7860 (N_7860,N_2924,N_1431);
and U7861 (N_7861,N_731,N_1133);
nor U7862 (N_7862,N_285,N_2028);
nand U7863 (N_7863,N_2644,N_3692);
xnor U7864 (N_7864,N_3726,N_1216);
or U7865 (N_7865,N_2908,N_3751);
and U7866 (N_7866,N_2322,N_2548);
nand U7867 (N_7867,N_337,N_1217);
xor U7868 (N_7868,N_574,N_3575);
and U7869 (N_7869,N_3272,N_142);
nand U7870 (N_7870,N_1696,N_3096);
xor U7871 (N_7871,N_2259,N_2522);
xor U7872 (N_7872,N_2252,N_977);
nor U7873 (N_7873,N_1571,N_334);
and U7874 (N_7874,N_2268,N_1148);
nor U7875 (N_7875,N_3394,N_1576);
or U7876 (N_7876,N_2156,N_3287);
or U7877 (N_7877,N_1911,N_2892);
nand U7878 (N_7878,N_3339,N_1905);
nor U7879 (N_7879,N_532,N_1312);
xor U7880 (N_7880,N_735,N_3114);
xnor U7881 (N_7881,N_1063,N_3065);
nor U7882 (N_7882,N_3753,N_2051);
nor U7883 (N_7883,N_2683,N_1598);
xor U7884 (N_7884,N_244,N_543);
xnor U7885 (N_7885,N_3985,N_3231);
nand U7886 (N_7886,N_2140,N_2220);
nor U7887 (N_7887,N_1224,N_594);
nand U7888 (N_7888,N_1199,N_1890);
xor U7889 (N_7889,N_3816,N_3726);
xor U7890 (N_7890,N_3799,N_3190);
nand U7891 (N_7891,N_2734,N_3490);
and U7892 (N_7892,N_294,N_1606);
nand U7893 (N_7893,N_1843,N_1996);
or U7894 (N_7894,N_481,N_156);
and U7895 (N_7895,N_103,N_2540);
xor U7896 (N_7896,N_3454,N_3868);
or U7897 (N_7897,N_1374,N_1149);
nor U7898 (N_7898,N_1061,N_1218);
nand U7899 (N_7899,N_1659,N_3569);
and U7900 (N_7900,N_47,N_3840);
nand U7901 (N_7901,N_3015,N_2761);
nor U7902 (N_7902,N_2494,N_2092);
nand U7903 (N_7903,N_2953,N_1607);
or U7904 (N_7904,N_3697,N_432);
or U7905 (N_7905,N_1579,N_1712);
nand U7906 (N_7906,N_3380,N_3978);
and U7907 (N_7907,N_872,N_3431);
xnor U7908 (N_7908,N_2509,N_1410);
and U7909 (N_7909,N_3525,N_1528);
nor U7910 (N_7910,N_3234,N_3709);
nand U7911 (N_7911,N_216,N_3098);
nor U7912 (N_7912,N_1207,N_1028);
and U7913 (N_7913,N_1644,N_1625);
xnor U7914 (N_7914,N_1945,N_36);
nand U7915 (N_7915,N_60,N_240);
nand U7916 (N_7916,N_1666,N_1810);
nor U7917 (N_7917,N_2840,N_1498);
and U7918 (N_7918,N_1325,N_3955);
xnor U7919 (N_7919,N_1290,N_2400);
xnor U7920 (N_7920,N_1369,N_885);
nand U7921 (N_7921,N_688,N_2941);
and U7922 (N_7922,N_372,N_3290);
and U7923 (N_7923,N_759,N_2524);
and U7924 (N_7924,N_523,N_2874);
xnor U7925 (N_7925,N_1196,N_3433);
and U7926 (N_7926,N_3785,N_1475);
nor U7927 (N_7927,N_2761,N_3296);
and U7928 (N_7928,N_2118,N_1170);
nor U7929 (N_7929,N_1598,N_2076);
and U7930 (N_7930,N_1515,N_3018);
nand U7931 (N_7931,N_653,N_3250);
and U7932 (N_7932,N_1407,N_1966);
and U7933 (N_7933,N_3015,N_103);
or U7934 (N_7934,N_2216,N_3046);
nor U7935 (N_7935,N_1369,N_3959);
or U7936 (N_7936,N_3473,N_996);
nor U7937 (N_7937,N_2511,N_3144);
and U7938 (N_7938,N_2006,N_110);
nor U7939 (N_7939,N_3545,N_1799);
and U7940 (N_7940,N_323,N_3757);
xor U7941 (N_7941,N_2530,N_3912);
nand U7942 (N_7942,N_1828,N_3250);
xnor U7943 (N_7943,N_843,N_305);
or U7944 (N_7944,N_430,N_2255);
and U7945 (N_7945,N_2398,N_10);
xor U7946 (N_7946,N_3929,N_3132);
nand U7947 (N_7947,N_640,N_3981);
xnor U7948 (N_7948,N_160,N_2271);
or U7949 (N_7949,N_3968,N_2662);
nor U7950 (N_7950,N_2045,N_2022);
nor U7951 (N_7951,N_708,N_3157);
and U7952 (N_7952,N_1711,N_2373);
nand U7953 (N_7953,N_759,N_3578);
or U7954 (N_7954,N_242,N_440);
or U7955 (N_7955,N_3648,N_1645);
nand U7956 (N_7956,N_1484,N_1383);
xnor U7957 (N_7957,N_2761,N_3860);
or U7958 (N_7958,N_219,N_2589);
nor U7959 (N_7959,N_2685,N_3736);
nand U7960 (N_7960,N_663,N_3398);
or U7961 (N_7961,N_77,N_3516);
nor U7962 (N_7962,N_955,N_2222);
and U7963 (N_7963,N_514,N_2572);
and U7964 (N_7964,N_262,N_2665);
xor U7965 (N_7965,N_2744,N_1338);
nor U7966 (N_7966,N_1440,N_1891);
and U7967 (N_7967,N_1562,N_1823);
xnor U7968 (N_7968,N_342,N_2225);
nor U7969 (N_7969,N_2515,N_2841);
nand U7970 (N_7970,N_2497,N_909);
xor U7971 (N_7971,N_1141,N_1929);
or U7972 (N_7972,N_316,N_3815);
or U7973 (N_7973,N_1361,N_3840);
nand U7974 (N_7974,N_3388,N_1077);
xor U7975 (N_7975,N_1510,N_496);
and U7976 (N_7976,N_3633,N_2826);
nor U7977 (N_7977,N_679,N_3509);
xnor U7978 (N_7978,N_66,N_1717);
nand U7979 (N_7979,N_1927,N_3516);
nand U7980 (N_7980,N_2247,N_3707);
or U7981 (N_7981,N_698,N_2257);
and U7982 (N_7982,N_2197,N_411);
nor U7983 (N_7983,N_1915,N_2705);
nor U7984 (N_7984,N_2412,N_2045);
xor U7985 (N_7985,N_2877,N_3030);
xor U7986 (N_7986,N_2085,N_2447);
nand U7987 (N_7987,N_3965,N_3845);
and U7988 (N_7988,N_2133,N_752);
nor U7989 (N_7989,N_1949,N_802);
nand U7990 (N_7990,N_345,N_3692);
or U7991 (N_7991,N_3274,N_1338);
nor U7992 (N_7992,N_1627,N_34);
or U7993 (N_7993,N_283,N_3892);
nor U7994 (N_7994,N_3309,N_3886);
nor U7995 (N_7995,N_3692,N_690);
nand U7996 (N_7996,N_3676,N_597);
nor U7997 (N_7997,N_1379,N_442);
xor U7998 (N_7998,N_1092,N_3408);
nand U7999 (N_7999,N_2416,N_870);
or U8000 (N_8000,N_4292,N_6307);
nor U8001 (N_8001,N_5935,N_4031);
xnor U8002 (N_8002,N_5992,N_4718);
nand U8003 (N_8003,N_5124,N_5296);
xor U8004 (N_8004,N_6120,N_6637);
and U8005 (N_8005,N_5790,N_4566);
nor U8006 (N_8006,N_6240,N_5174);
nor U8007 (N_8007,N_6355,N_6782);
nor U8008 (N_8008,N_5239,N_4035);
or U8009 (N_8009,N_6288,N_4772);
and U8010 (N_8010,N_6687,N_4583);
and U8011 (N_8011,N_4809,N_5156);
or U8012 (N_8012,N_4419,N_5898);
nor U8013 (N_8013,N_7544,N_6213);
xnor U8014 (N_8014,N_6962,N_5742);
and U8015 (N_8015,N_4374,N_7246);
xnor U8016 (N_8016,N_4064,N_5751);
nand U8017 (N_8017,N_7134,N_6573);
xnor U8018 (N_8018,N_5622,N_5291);
or U8019 (N_8019,N_4254,N_6456);
nor U8020 (N_8020,N_7694,N_6952);
nor U8021 (N_8021,N_6950,N_7122);
nand U8022 (N_8022,N_6802,N_5219);
nor U8023 (N_8023,N_5545,N_7535);
or U8024 (N_8024,N_7120,N_4877);
nor U8025 (N_8025,N_7732,N_5747);
and U8026 (N_8026,N_7001,N_4644);
or U8027 (N_8027,N_6423,N_6741);
nor U8028 (N_8028,N_5508,N_4965);
and U8029 (N_8029,N_4312,N_7680);
nand U8030 (N_8030,N_5894,N_5026);
nor U8031 (N_8031,N_5380,N_5674);
nand U8032 (N_8032,N_4438,N_4316);
and U8033 (N_8033,N_5815,N_5340);
xor U8034 (N_8034,N_5637,N_6984);
xor U8035 (N_8035,N_5956,N_4342);
and U8036 (N_8036,N_6908,N_7755);
or U8037 (N_8037,N_4236,N_4645);
xor U8038 (N_8038,N_5796,N_7237);
xor U8039 (N_8039,N_7356,N_6762);
or U8040 (N_8040,N_5247,N_4066);
and U8041 (N_8041,N_7287,N_4350);
nand U8042 (N_8042,N_5682,N_4859);
and U8043 (N_8043,N_5140,N_4627);
or U8044 (N_8044,N_4764,N_5726);
xor U8045 (N_8045,N_4789,N_6679);
and U8046 (N_8046,N_6860,N_7060);
or U8047 (N_8047,N_5617,N_6137);
xnor U8048 (N_8048,N_7688,N_6595);
or U8049 (N_8049,N_6246,N_6533);
nor U8050 (N_8050,N_6453,N_4516);
xnor U8051 (N_8051,N_6569,N_4737);
nor U8052 (N_8052,N_4686,N_7437);
nor U8053 (N_8053,N_5990,N_6269);
xor U8054 (N_8054,N_7880,N_5628);
nor U8055 (N_8055,N_5137,N_5338);
and U8056 (N_8056,N_4261,N_4164);
or U8057 (N_8057,N_7998,N_7005);
and U8058 (N_8058,N_7536,N_7126);
xnor U8059 (N_8059,N_5647,N_5311);
and U8060 (N_8060,N_7509,N_6194);
xor U8061 (N_8061,N_7840,N_6346);
xor U8062 (N_8062,N_4638,N_7405);
nand U8063 (N_8063,N_5408,N_7374);
or U8064 (N_8064,N_7752,N_7958);
nand U8065 (N_8065,N_5700,N_4293);
and U8066 (N_8066,N_6179,N_7964);
xor U8067 (N_8067,N_6799,N_6503);
nor U8068 (N_8068,N_6476,N_6159);
or U8069 (N_8069,N_4882,N_5080);
nand U8070 (N_8070,N_4763,N_6664);
nor U8071 (N_8071,N_7009,N_5854);
and U8072 (N_8072,N_4068,N_4571);
and U8073 (N_8073,N_6220,N_7894);
or U8074 (N_8074,N_4620,N_4541);
or U8075 (N_8075,N_5094,N_5832);
xnor U8076 (N_8076,N_7628,N_6810);
nor U8077 (N_8077,N_6534,N_7039);
or U8078 (N_8078,N_5272,N_6107);
and U8079 (N_8079,N_5928,N_4383);
xnor U8080 (N_8080,N_4576,N_7708);
nand U8081 (N_8081,N_4547,N_7625);
nand U8082 (N_8082,N_4659,N_4818);
nor U8083 (N_8083,N_6452,N_6410);
nor U8084 (N_8084,N_7472,N_7273);
or U8085 (N_8085,N_6555,N_6309);
and U8086 (N_8086,N_5615,N_7041);
or U8087 (N_8087,N_4412,N_6277);
nand U8088 (N_8088,N_5176,N_6876);
xor U8089 (N_8089,N_5781,N_7026);
nor U8090 (N_8090,N_4318,N_6302);
and U8091 (N_8091,N_6446,N_6460);
nand U8092 (N_8092,N_5441,N_5512);
nand U8093 (N_8093,N_7718,N_4949);
xnor U8094 (N_8094,N_5459,N_4218);
nor U8095 (N_8095,N_6133,N_4043);
and U8096 (N_8096,N_5131,N_6942);
xor U8097 (N_8097,N_5970,N_7845);
xor U8098 (N_8098,N_7877,N_6671);
and U8099 (N_8099,N_6459,N_7723);
nand U8100 (N_8100,N_5030,N_7502);
or U8101 (N_8101,N_4089,N_7646);
nor U8102 (N_8102,N_5933,N_7231);
xnor U8103 (N_8103,N_7100,N_4482);
nand U8104 (N_8104,N_5654,N_7985);
and U8105 (N_8105,N_5175,N_6372);
xnor U8106 (N_8106,N_5091,N_6585);
and U8107 (N_8107,N_7063,N_7201);
and U8108 (N_8108,N_4067,N_5258);
and U8109 (N_8109,N_7864,N_6182);
nor U8110 (N_8110,N_6626,N_4432);
and U8111 (N_8111,N_7158,N_4868);
nor U8112 (N_8112,N_5191,N_4952);
nor U8113 (N_8113,N_4749,N_7088);
nand U8114 (N_8114,N_5612,N_6449);
and U8115 (N_8115,N_5704,N_5973);
xor U8116 (N_8116,N_7253,N_5067);
nand U8117 (N_8117,N_7711,N_7234);
nor U8118 (N_8118,N_4022,N_7510);
and U8119 (N_8119,N_5349,N_7922);
or U8120 (N_8120,N_5911,N_5447);
xor U8121 (N_8121,N_4819,N_7681);
or U8122 (N_8122,N_6354,N_7753);
nand U8123 (N_8123,N_6963,N_6634);
xor U8124 (N_8124,N_5630,N_7553);
xor U8125 (N_8125,N_5233,N_6896);
or U8126 (N_8126,N_5955,N_7232);
xnor U8127 (N_8127,N_6365,N_6368);
or U8128 (N_8128,N_7715,N_5966);
xnor U8129 (N_8129,N_5472,N_6006);
nand U8130 (N_8130,N_5574,N_4615);
nor U8131 (N_8131,N_7298,N_6471);
nand U8132 (N_8132,N_4013,N_5871);
nor U8133 (N_8133,N_6135,N_4979);
nand U8134 (N_8134,N_4943,N_4270);
or U8135 (N_8135,N_6150,N_7630);
and U8136 (N_8136,N_4814,N_4880);
and U8137 (N_8137,N_5019,N_7395);
nor U8138 (N_8138,N_4656,N_4369);
nand U8139 (N_8139,N_6188,N_5365);
and U8140 (N_8140,N_5716,N_6168);
or U8141 (N_8141,N_6532,N_4277);
or U8142 (N_8142,N_6201,N_5982);
and U8143 (N_8143,N_5814,N_6932);
or U8144 (N_8144,N_7710,N_7187);
nand U8145 (N_8145,N_5061,N_5998);
and U8146 (N_8146,N_4307,N_6980);
nor U8147 (N_8147,N_4006,N_7609);
xnor U8148 (N_8148,N_5445,N_7062);
nor U8149 (N_8149,N_6987,N_6224);
or U8150 (N_8150,N_6378,N_4183);
nor U8151 (N_8151,N_6046,N_7386);
xnor U8152 (N_8152,N_7988,N_7926);
and U8153 (N_8153,N_5975,N_4077);
and U8154 (N_8154,N_5830,N_5535);
nor U8155 (N_8155,N_7455,N_4777);
nand U8156 (N_8156,N_6601,N_5464);
and U8157 (N_8157,N_6968,N_6698);
nor U8158 (N_8158,N_4507,N_4508);
nand U8159 (N_8159,N_6755,N_6828);
nand U8160 (N_8160,N_6348,N_4456);
and U8161 (N_8161,N_7866,N_4107);
xor U8162 (N_8162,N_6711,N_5693);
and U8163 (N_8163,N_5688,N_6743);
nand U8164 (N_8164,N_7571,N_4224);
and U8165 (N_8165,N_6290,N_7594);
and U8166 (N_8166,N_6273,N_6363);
and U8167 (N_8167,N_7826,N_4172);
or U8168 (N_8168,N_6853,N_5819);
xnor U8169 (N_8169,N_7731,N_6903);
and U8170 (N_8170,N_5188,N_6123);
nor U8171 (N_8171,N_4595,N_4247);
xnor U8172 (N_8172,N_7235,N_7180);
and U8173 (N_8173,N_7383,N_5270);
nand U8174 (N_8174,N_5125,N_5566);
or U8175 (N_8175,N_6697,N_5957);
xnor U8176 (N_8176,N_5549,N_6519);
xnor U8177 (N_8177,N_7882,N_7637);
nor U8178 (N_8178,N_5639,N_6832);
or U8179 (N_8179,N_4591,N_7130);
or U8180 (N_8180,N_5235,N_4495);
nand U8181 (N_8181,N_4460,N_5346);
and U8182 (N_8182,N_5817,N_5473);
and U8183 (N_8183,N_6037,N_6837);
nand U8184 (N_8184,N_4671,N_6023);
and U8185 (N_8185,N_4162,N_4742);
or U8186 (N_8186,N_5106,N_4084);
nor U8187 (N_8187,N_7586,N_7085);
or U8188 (N_8188,N_5037,N_4073);
or U8189 (N_8189,N_6584,N_7045);
xnor U8190 (N_8190,N_5821,N_7524);
nand U8191 (N_8191,N_6324,N_5979);
nor U8192 (N_8192,N_5243,N_4379);
xnor U8193 (N_8193,N_5748,N_7538);
and U8194 (N_8194,N_6052,N_4646);
and U8195 (N_8195,N_5727,N_7016);
nor U8196 (N_8196,N_6353,N_6063);
nor U8197 (N_8197,N_6969,N_7123);
xor U8198 (N_8198,N_6482,N_6675);
and U8199 (N_8199,N_4904,N_4058);
and U8200 (N_8200,N_7159,N_6596);
nand U8201 (N_8201,N_5586,N_7031);
and U8202 (N_8202,N_4268,N_5274);
nor U8203 (N_8203,N_4578,N_7636);
xor U8204 (N_8204,N_6631,N_6097);
nor U8205 (N_8205,N_7413,N_5944);
and U8206 (N_8206,N_6732,N_5534);
and U8207 (N_8207,N_4529,N_7893);
xnor U8208 (N_8208,N_4311,N_6017);
and U8209 (N_8209,N_6892,N_6529);
and U8210 (N_8210,N_6153,N_5558);
nand U8211 (N_8211,N_5516,N_6866);
or U8212 (N_8212,N_6380,N_5948);
nor U8213 (N_8213,N_7531,N_5964);
or U8214 (N_8214,N_4855,N_6629);
or U8215 (N_8215,N_7687,N_4228);
and U8216 (N_8216,N_4304,N_6727);
and U8217 (N_8217,N_7164,N_4746);
nand U8218 (N_8218,N_7859,N_7236);
or U8219 (N_8219,N_6299,N_5224);
nand U8220 (N_8220,N_5564,N_7701);
xnor U8221 (N_8221,N_4621,N_7938);
nor U8222 (N_8222,N_6644,N_5881);
xnor U8223 (N_8223,N_5448,N_7353);
nand U8224 (N_8224,N_5303,N_7427);
or U8225 (N_8225,N_4017,N_5392);
nand U8226 (N_8226,N_5606,N_6633);
xnor U8227 (N_8227,N_5527,N_5487);
or U8228 (N_8228,N_5684,N_5707);
nand U8229 (N_8229,N_7730,N_7286);
nand U8230 (N_8230,N_7378,N_7275);
nor U8231 (N_8231,N_6742,N_4244);
and U8232 (N_8232,N_5642,N_4094);
nand U8233 (N_8233,N_4208,N_4267);
xor U8234 (N_8234,N_5417,N_4888);
or U8235 (N_8235,N_7768,N_7573);
nor U8236 (N_8236,N_5605,N_6357);
xnor U8237 (N_8237,N_4543,N_5208);
nand U8238 (N_8238,N_6989,N_6557);
nor U8239 (N_8239,N_6259,N_6500);
or U8240 (N_8240,N_6214,N_4009);
nand U8241 (N_8241,N_4520,N_5348);
and U8242 (N_8242,N_7418,N_6759);
or U8243 (N_8243,N_5143,N_6630);
nand U8244 (N_8244,N_6436,N_7094);
and U8245 (N_8245,N_4352,N_7460);
nand U8246 (N_8246,N_7528,N_7025);
nor U8247 (N_8247,N_5240,N_7254);
or U8248 (N_8248,N_5976,N_5225);
nor U8249 (N_8249,N_5032,N_7458);
and U8250 (N_8250,N_5771,N_6775);
or U8251 (N_8251,N_5801,N_7243);
nor U8252 (N_8252,N_7098,N_5342);
nor U8253 (N_8253,N_6744,N_5685);
nand U8254 (N_8254,N_7950,N_4417);
nor U8255 (N_8255,N_6767,N_7690);
or U8256 (N_8256,N_5749,N_5362);
or U8257 (N_8257,N_6486,N_6696);
xor U8258 (N_8258,N_6493,N_7328);
xnor U8259 (N_8259,N_5020,N_6833);
xnor U8260 (N_8260,N_5552,N_7327);
nand U8261 (N_8261,N_5744,N_7284);
or U8262 (N_8262,N_7817,N_5532);
nand U8263 (N_8263,N_5287,N_6254);
or U8264 (N_8264,N_6923,N_5288);
xor U8265 (N_8265,N_7682,N_5591);
or U8266 (N_8266,N_6680,N_5205);
and U8267 (N_8267,N_4681,N_5256);
xnor U8268 (N_8268,N_5409,N_7075);
nand U8269 (N_8269,N_6538,N_6885);
and U8270 (N_8270,N_5370,N_4725);
nor U8271 (N_8271,N_6461,N_6966);
nand U8272 (N_8272,N_7279,N_4229);
or U8273 (N_8273,N_5501,N_6096);
nand U8274 (N_8274,N_7673,N_7972);
xnor U8275 (N_8275,N_6216,N_7696);
nor U8276 (N_8276,N_6547,N_4942);
or U8277 (N_8277,N_5379,N_4357);
nand U8278 (N_8278,N_6349,N_7317);
and U8279 (N_8279,N_4424,N_6341);
and U8280 (N_8280,N_6702,N_4954);
xnor U8281 (N_8281,N_6704,N_7303);
nand U8282 (N_8282,N_4488,N_6899);
or U8283 (N_8283,N_4063,N_4360);
nor U8284 (N_8284,N_6412,N_5165);
nand U8285 (N_8285,N_4905,N_6965);
nand U8286 (N_8286,N_5589,N_7067);
and U8287 (N_8287,N_5133,N_5561);
or U8288 (N_8288,N_6575,N_7911);
xnor U8289 (N_8289,N_7048,N_6893);
nor U8290 (N_8290,N_6389,N_6474);
nand U8291 (N_8291,N_4692,N_4697);
nand U8292 (N_8292,N_7017,N_5838);
nor U8293 (N_8293,N_6242,N_4110);
nor U8294 (N_8294,N_7583,N_5363);
nand U8295 (N_8295,N_4467,N_4444);
nor U8296 (N_8296,N_7358,N_4023);
nor U8297 (N_8297,N_6174,N_7487);
or U8298 (N_8298,N_6850,N_5883);
or U8299 (N_8299,N_5255,N_7526);
nor U8300 (N_8300,N_5805,N_6255);
and U8301 (N_8301,N_6838,N_4033);
xor U8302 (N_8302,N_5112,N_5946);
or U8303 (N_8303,N_7957,N_5740);
xor U8304 (N_8304,N_6870,N_7002);
and U8305 (N_8305,N_5705,N_7467);
nand U8306 (N_8306,N_5579,N_5537);
xor U8307 (N_8307,N_6959,N_6909);
or U8308 (N_8308,N_5439,N_6409);
and U8309 (N_8309,N_5197,N_6934);
xnor U8310 (N_8310,N_6847,N_5273);
and U8311 (N_8311,N_5793,N_5152);
nor U8312 (N_8312,N_7080,N_7439);
nor U8313 (N_8313,N_4521,N_5282);
xor U8314 (N_8314,N_7267,N_4329);
nor U8315 (N_8315,N_5683,N_7995);
and U8316 (N_8316,N_7647,N_7951);
and U8317 (N_8317,N_4643,N_4300);
and U8318 (N_8318,N_7978,N_4601);
nand U8319 (N_8319,N_5446,N_4472);
or U8320 (N_8320,N_5644,N_7324);
xnor U8321 (N_8321,N_4333,N_6005);
or U8322 (N_8322,N_4054,N_7268);
nand U8323 (N_8323,N_6681,N_7678);
and U8324 (N_8324,N_7970,N_6639);
nand U8325 (N_8325,N_6377,N_7357);
nor U8326 (N_8326,N_5078,N_4959);
and U8327 (N_8327,N_5024,N_5171);
nor U8328 (N_8328,N_5449,N_5643);
nor U8329 (N_8329,N_7841,N_7495);
nor U8330 (N_8330,N_6091,N_4061);
or U8331 (N_8331,N_4629,N_4186);
nand U8332 (N_8332,N_5594,N_6848);
and U8333 (N_8333,N_4505,N_6072);
nand U8334 (N_8334,N_5367,N_5358);
nor U8335 (N_8335,N_5712,N_5522);
nand U8336 (N_8336,N_6628,N_5570);
or U8337 (N_8337,N_6490,N_6401);
xor U8338 (N_8338,N_7127,N_5246);
xor U8339 (N_8339,N_7283,N_6148);
or U8340 (N_8340,N_7902,N_6935);
or U8341 (N_8341,N_5920,N_7396);
and U8342 (N_8342,N_7314,N_5936);
xnor U8343 (N_8343,N_5610,N_6071);
nor U8344 (N_8344,N_4986,N_7494);
nor U8345 (N_8345,N_4388,N_6347);
nor U8346 (N_8346,N_7415,N_7953);
nor U8347 (N_8347,N_6815,N_7908);
or U8348 (N_8348,N_4250,N_7705);
or U8349 (N_8349,N_5395,N_6880);
nand U8350 (N_8350,N_7466,N_5590);
nand U8351 (N_8351,N_5264,N_5772);
nor U8352 (N_8352,N_6811,N_6852);
and U8353 (N_8353,N_5271,N_5638);
and U8354 (N_8354,N_6798,N_6668);
or U8355 (N_8355,N_6572,N_6663);
or U8356 (N_8356,N_4288,N_5251);
nor U8357 (N_8357,N_5325,N_7720);
nor U8358 (N_8358,N_6283,N_6638);
and U8359 (N_8359,N_5050,N_7239);
xnor U8360 (N_8360,N_4226,N_4950);
nor U8361 (N_8361,N_6289,N_7740);
or U8362 (N_8362,N_7054,N_4422);
or U8363 (N_8363,N_4210,N_4512);
and U8364 (N_8364,N_5664,N_5257);
nor U8365 (N_8365,N_7672,N_6895);
xor U8366 (N_8366,N_6293,N_4849);
nand U8367 (N_8367,N_7300,N_7937);
nor U8368 (N_8368,N_4173,N_4553);
nand U8369 (N_8369,N_4452,N_4633);
or U8370 (N_8370,N_5179,N_5070);
and U8371 (N_8371,N_7564,N_7862);
nor U8372 (N_8372,N_7961,N_5714);
and U8373 (N_8373,N_4135,N_5728);
nor U8374 (N_8374,N_4474,N_5321);
or U8375 (N_8375,N_6425,N_4118);
and U8376 (N_8376,N_5785,N_4996);
nand U8377 (N_8377,N_6130,N_7621);
or U8378 (N_8378,N_6451,N_7412);
xnor U8379 (N_8379,N_6768,N_4929);
xnor U8380 (N_8380,N_7741,N_6985);
xnor U8381 (N_8381,N_5455,N_7361);
nor U8382 (N_8382,N_5857,N_6043);
xor U8383 (N_8383,N_4639,N_5283);
nand U8384 (N_8384,N_4797,N_7613);
and U8385 (N_8385,N_4124,N_6983);
nand U8386 (N_8386,N_5962,N_5598);
nand U8387 (N_8387,N_5525,N_4890);
and U8388 (N_8388,N_7533,N_5602);
xnor U8389 (N_8389,N_6297,N_4624);
nor U8390 (N_8390,N_6406,N_6276);
nor U8391 (N_8391,N_6994,N_6577);
xor U8392 (N_8392,N_6171,N_7852);
nand U8393 (N_8393,N_7527,N_4750);
or U8394 (N_8394,N_5076,N_4088);
nor U8395 (N_8395,N_6057,N_6703);
nand U8396 (N_8396,N_5666,N_6085);
or U8397 (N_8397,N_6558,N_7912);
nor U8398 (N_8398,N_6625,N_4389);
nand U8399 (N_8399,N_7059,N_7581);
xor U8400 (N_8400,N_6087,N_5294);
nand U8401 (N_8401,N_6065,N_4264);
nor U8402 (N_8402,N_7216,N_7517);
nor U8403 (N_8403,N_5876,N_5818);
or U8404 (N_8404,N_5307,N_5952);
nand U8405 (N_8405,N_5505,N_5835);
or U8406 (N_8406,N_6086,N_4168);
nor U8407 (N_8407,N_6236,N_6121);
and U8408 (N_8408,N_5186,N_7350);
xor U8409 (N_8409,N_6369,N_6192);
nand U8410 (N_8410,N_7480,N_6560);
nor U8411 (N_8411,N_5884,N_5645);
nand U8412 (N_8412,N_4720,N_7560);
nor U8413 (N_8413,N_4978,N_4145);
nand U8414 (N_8414,N_7401,N_7762);
nand U8415 (N_8415,N_7373,N_6082);
xnor U8416 (N_8416,N_5231,N_7649);
nor U8417 (N_8417,N_5611,N_5426);
nand U8418 (N_8418,N_5902,N_6986);
nor U8419 (N_8419,N_7505,N_7256);
xnor U8420 (N_8420,N_6498,N_4745);
xnor U8421 (N_8421,N_4668,N_7722);
nor U8422 (N_8422,N_4913,N_7241);
nand U8423 (N_8423,N_6954,N_7733);
and U8424 (N_8424,N_4885,N_7053);
nor U8425 (N_8425,N_6588,N_4399);
or U8426 (N_8426,N_5985,N_4366);
nand U8427 (N_8427,N_4446,N_4705);
and U8428 (N_8428,N_7179,N_5187);
or U8429 (N_8429,N_6937,N_5937);
nor U8430 (N_8430,N_4425,N_4353);
and U8431 (N_8431,N_6705,N_6215);
and U8432 (N_8432,N_7290,N_5132);
xor U8433 (N_8433,N_6800,N_7295);
and U8434 (N_8434,N_4121,N_5721);
nor U8435 (N_8435,N_5298,N_4744);
xor U8436 (N_8436,N_6287,N_5382);
nand U8437 (N_8437,N_4572,N_7962);
or U8438 (N_8438,N_5870,N_7233);
nor U8439 (N_8439,N_7148,N_6008);
nand U8440 (N_8440,N_5092,N_6310);
and U8441 (N_8441,N_7887,N_7345);
xor U8442 (N_8442,N_6241,N_6157);
or U8443 (N_8443,N_4728,N_7251);
or U8444 (N_8444,N_7457,N_5119);
and U8445 (N_8445,N_7803,N_5368);
or U8446 (N_8446,N_5897,N_4984);
and U8447 (N_8447,N_7843,N_6292);
xnor U8448 (N_8448,N_4176,N_4569);
nor U8449 (N_8449,N_4866,N_7567);
xnor U8450 (N_8450,N_5006,N_5347);
nand U8451 (N_8451,N_5461,N_7546);
nor U8452 (N_8452,N_6660,N_4328);
and U8453 (N_8453,N_7804,N_6695);
nand U8454 (N_8454,N_6432,N_4730);
and U8455 (N_8455,N_7656,N_5322);
xor U8456 (N_8456,N_5227,N_4149);
or U8457 (N_8457,N_7810,N_6865);
nand U8458 (N_8458,N_7116,N_5045);
and U8459 (N_8459,N_6092,N_4606);
nand U8460 (N_8460,N_7568,N_7523);
nor U8461 (N_8461,N_4455,N_5249);
nor U8462 (N_8462,N_4617,N_6499);
xnor U8463 (N_8463,N_5969,N_4171);
xor U8464 (N_8464,N_6518,N_7677);
or U8465 (N_8465,N_5064,N_5977);
nor U8466 (N_8466,N_6877,N_4046);
and U8467 (N_8467,N_6763,N_4331);
nor U8468 (N_8468,N_5162,N_6677);
and U8469 (N_8469,N_6325,N_7305);
and U8470 (N_8470,N_5791,N_4439);
xor U8471 (N_8471,N_5318,N_4498);
and U8472 (N_8472,N_4871,N_7477);
or U8473 (N_8473,N_5351,N_5300);
nand U8474 (N_8474,N_7102,N_6941);
and U8475 (N_8475,N_5277,N_6394);
and U8476 (N_8476,N_5405,N_5483);
and U8477 (N_8477,N_4497,N_5048);
or U8478 (N_8478,N_6846,N_5324);
xnor U8479 (N_8479,N_4309,N_5978);
and U8480 (N_8480,N_7529,N_4458);
or U8481 (N_8481,N_6155,N_7081);
and U8482 (N_8482,N_5345,N_6882);
nor U8483 (N_8483,N_7616,N_6897);
or U8484 (N_8484,N_4448,N_6278);
nand U8485 (N_8485,N_4287,N_4775);
or U8486 (N_8486,N_4131,N_4504);
nor U8487 (N_8487,N_4781,N_6080);
xor U8488 (N_8488,N_4807,N_7097);
nand U8489 (N_8489,N_6505,N_6614);
or U8490 (N_8490,N_4754,N_7624);
xor U8491 (N_8491,N_7749,N_7389);
nor U8492 (N_8492,N_4280,N_4144);
and U8493 (N_8493,N_6258,N_7868);
or U8494 (N_8494,N_7445,N_5960);
xnor U8495 (N_8495,N_7023,N_6976);
xor U8496 (N_8496,N_6274,N_6167);
nand U8497 (N_8497,N_7934,N_5326);
and U8498 (N_8498,N_7598,N_4204);
and U8499 (N_8499,N_6624,N_7113);
nand U8500 (N_8500,N_5673,N_6340);
or U8501 (N_8501,N_5432,N_6454);
nor U8502 (N_8502,N_5916,N_7092);
nand U8503 (N_8503,N_6039,N_6612);
xnor U8504 (N_8504,N_7796,N_4815);
or U8505 (N_8505,N_6203,N_6011);
or U8506 (N_8506,N_7042,N_7576);
and U8507 (N_8507,N_4294,N_5344);
nand U8508 (N_8508,N_5289,N_5115);
nor U8509 (N_8509,N_5603,N_7744);
or U8510 (N_8510,N_7674,N_5044);
nand U8511 (N_8511,N_7490,N_4182);
or U8512 (N_8512,N_6266,N_6227);
nand U8513 (N_8513,N_5263,N_6308);
and U8514 (N_8514,N_4394,N_5556);
nor U8515 (N_8515,N_6661,N_7227);
nand U8516 (N_8516,N_4808,N_7813);
nor U8517 (N_8517,N_7883,N_4873);
nand U8518 (N_8518,N_4729,N_4833);
or U8519 (N_8519,N_6279,N_6706);
xor U8520 (N_8520,N_6824,N_5889);
xor U8521 (N_8521,N_5230,N_5077);
nor U8522 (N_8522,N_6604,N_6864);
and U8523 (N_8523,N_6718,N_5378);
and U8524 (N_8524,N_7955,N_5265);
or U8525 (N_8525,N_7842,N_5416);
and U8526 (N_8526,N_5433,N_4551);
and U8527 (N_8527,N_7865,N_7408);
nand U8528 (N_8528,N_6233,N_4874);
nor U8529 (N_8529,N_4381,N_6462);
nand U8530 (N_8530,N_6015,N_6669);
and U8531 (N_8531,N_4271,N_5047);
or U8532 (N_8532,N_5085,N_6749);
xnor U8533 (N_8533,N_4972,N_4096);
nor U8534 (N_8534,N_5576,N_4079);
and U8535 (N_8535,N_5073,N_5074);
nand U8536 (N_8536,N_7947,N_4533);
xnor U8537 (N_8537,N_4678,N_6665);
nor U8538 (N_8538,N_6536,N_7837);
nand U8539 (N_8539,N_5309,N_5752);
nor U8540 (N_8540,N_4510,N_5734);
nor U8541 (N_8541,N_6685,N_6186);
xor U8542 (N_8542,N_4989,N_5057);
or U8543 (N_8543,N_7872,N_6527);
nand U8544 (N_8544,N_7593,N_4349);
nand U8545 (N_8545,N_4604,N_5923);
and U8546 (N_8546,N_7819,N_7109);
nand U8547 (N_8547,N_7663,N_5178);
and U8548 (N_8548,N_4092,N_7056);
xor U8549 (N_8549,N_7914,N_5994);
and U8550 (N_8550,N_4526,N_4714);
and U8551 (N_8551,N_6012,N_6715);
or U8552 (N_8552,N_7362,N_4491);
and U8553 (N_8553,N_4704,N_4246);
xor U8554 (N_8554,N_5477,N_7795);
nor U8555 (N_8555,N_6791,N_4517);
and U8556 (N_8556,N_4194,N_6021);
nand U8557 (N_8557,N_5823,N_7065);
or U8558 (N_8558,N_5577,N_4918);
or U8559 (N_8559,N_6344,N_4605);
nor U8560 (N_8560,N_4637,N_4941);
nand U8561 (N_8561,N_5198,N_6922);
nor U8562 (N_8562,N_4593,N_7029);
xnor U8563 (N_8563,N_6772,N_4922);
or U8564 (N_8564,N_5765,N_4203);
and U8565 (N_8565,N_7518,N_6801);
xnor U8566 (N_8566,N_4515,N_7631);
xnor U8567 (N_8567,N_5706,N_6956);
and U8568 (N_8568,N_7247,N_6939);
xnor U8569 (N_8569,N_5023,N_7105);
or U8570 (N_8570,N_6465,N_7507);
xnor U8571 (N_8571,N_7166,N_5136);
nor U8572 (N_8572,N_7549,N_5601);
nor U8573 (N_8573,N_6049,N_4122);
nor U8574 (N_8574,N_6602,N_4796);
nand U8575 (N_8575,N_6090,N_4211);
and U8576 (N_8576,N_6177,N_5138);
and U8577 (N_8577,N_6701,N_7438);
xor U8578 (N_8578,N_6520,N_7774);
or U8579 (N_8579,N_5524,N_5496);
and U8580 (N_8580,N_7860,N_5901);
nand U8581 (N_8581,N_6765,N_6373);
or U8582 (N_8582,N_4485,N_4302);
xor U8583 (N_8583,N_5528,N_6291);
and U8584 (N_8584,N_7695,N_5457);
and U8585 (N_8585,N_6112,N_7190);
nor U8586 (N_8586,N_6925,N_6285);
and U8587 (N_8587,N_4588,N_4716);
or U8588 (N_8588,N_4848,N_4751);
and U8589 (N_8589,N_7793,N_6058);
nand U8590 (N_8590,N_5531,N_5631);
nand U8591 (N_8591,N_5538,N_6352);
nand U8592 (N_8592,N_4560,N_6656);
nand U8593 (N_8593,N_7443,N_7311);
or U8594 (N_8594,N_4050,N_4915);
nor U8595 (N_8595,N_7262,N_6332);
and U8596 (N_8596,N_6542,N_6504);
nor U8597 (N_8597,N_4713,N_7585);
xnor U8598 (N_8598,N_6424,N_6163);
xor U8599 (N_8599,N_6078,N_6371);
nor U8600 (N_8600,N_5497,N_7221);
xnor U8601 (N_8601,N_4683,N_7765);
nor U8602 (N_8602,N_5142,N_4380);
or U8603 (N_8603,N_6145,N_7064);
or U8604 (N_8604,N_7556,N_7642);
and U8605 (N_8605,N_4128,N_5813);
nor U8606 (N_8606,N_6313,N_4008);
or U8607 (N_8607,N_5411,N_4103);
nor U8608 (N_8608,N_4049,N_7493);
nor U8609 (N_8609,N_5810,N_5914);
and U8610 (N_8610,N_5245,N_6075);
nand U8611 (N_8611,N_5795,N_5567);
nor U8612 (N_8612,N_4788,N_4799);
nor U8613 (N_8613,N_7337,N_7871);
or U8614 (N_8614,N_5129,N_5252);
xor U8615 (N_8615,N_7555,N_4177);
and U8616 (N_8616,N_7541,N_4223);
nor U8617 (N_8617,N_5502,N_4528);
and U8618 (N_8618,N_6433,N_4825);
nand U8619 (N_8619,N_4939,N_4976);
nor U8620 (N_8620,N_5784,N_5940);
or U8621 (N_8621,N_7326,N_4231);
or U8622 (N_8622,N_5002,N_4732);
and U8623 (N_8623,N_4199,N_4863);
xor U8624 (N_8624,N_6404,N_6996);
and U8625 (N_8625,N_7787,N_4493);
nand U8626 (N_8626,N_7689,N_4894);
or U8627 (N_8627,N_6651,N_6546);
nand U8628 (N_8628,N_5520,N_5158);
and U8629 (N_8629,N_4308,N_4405);
nand U8630 (N_8630,N_7836,N_7354);
or U8631 (N_8631,N_4057,N_7479);
and U8632 (N_8632,N_6928,N_4655);
nand U8633 (N_8633,N_4195,N_6180);
nor U8634 (N_8634,N_4420,N_6507);
xor U8635 (N_8635,N_4150,N_5012);
nor U8636 (N_8636,N_7686,N_4711);
nand U8637 (N_8637,N_7206,N_6600);
or U8638 (N_8638,N_6463,N_7878);
nor U8639 (N_8639,N_7579,N_4385);
xnor U8640 (N_8640,N_5836,N_5438);
xnor U8641 (N_8641,N_7724,N_6339);
or U8642 (N_8642,N_6257,N_4459);
nand U8643 (N_8643,N_4870,N_6879);
nand U8644 (N_8644,N_4296,N_6126);
or U8645 (N_8645,N_4648,N_6305);
or U8646 (N_8646,N_4895,N_7035);
nor U8647 (N_8647,N_6181,N_5018);
nand U8648 (N_8648,N_7101,N_5825);
nor U8649 (N_8649,N_4886,N_6235);
and U8650 (N_8650,N_4523,N_4060);
nand U8651 (N_8651,N_6228,N_5121);
nand U8652 (N_8652,N_5183,N_6358);
and U8653 (N_8653,N_7948,N_4235);
nand U8654 (N_8654,N_7154,N_6961);
nor U8655 (N_8655,N_4140,N_5972);
and U8656 (N_8656,N_4717,N_4891);
and U8657 (N_8657,N_7521,N_5093);
or U8658 (N_8658,N_4411,N_5425);
and U8659 (N_8659,N_6829,N_5550);
nor U8660 (N_8660,N_6793,N_7258);
xor U8661 (N_8661,N_7921,N_5655);
or U8662 (N_8662,N_6329,N_4025);
and U8663 (N_8663,N_4919,N_5947);
xnor U8664 (N_8664,N_6051,N_7770);
xor U8665 (N_8665,N_4243,N_6418);
nand U8666 (N_8666,N_7773,N_7945);
nor U8667 (N_8667,N_5646,N_5027);
nor U8668 (N_8668,N_4015,N_4492);
and U8669 (N_8669,N_4707,N_5743);
xnor U8670 (N_8670,N_5199,N_4259);
nor U8671 (N_8671,N_6918,N_5120);
and U8672 (N_8672,N_4765,N_6884);
nor U8673 (N_8673,N_4161,N_5401);
or U8674 (N_8674,N_5746,N_4373);
nor U8675 (N_8675,N_6264,N_5109);
and U8676 (N_8676,N_4346,N_5335);
xnor U8677 (N_8677,N_5377,N_6861);
nand U8678 (N_8678,N_5562,N_5100);
nor U8679 (N_8679,N_4597,N_4305);
nor U8680 (N_8680,N_6977,N_6991);
and U8681 (N_8681,N_6618,N_7889);
nor U8682 (N_8682,N_7569,N_6683);
nor U8683 (N_8683,N_6069,N_4070);
or U8684 (N_8684,N_5519,N_5922);
nor U8685 (N_8685,N_7366,N_6261);
nor U8686 (N_8686,N_5398,N_7384);
and U8687 (N_8687,N_4650,N_6946);
xor U8688 (N_8688,N_4845,N_6881);
nor U8689 (N_8689,N_7539,N_7618);
and U8690 (N_8690,N_5260,N_4626);
or U8691 (N_8691,N_5938,N_5518);
nand U8692 (N_8692,N_5015,N_7750);
nor U8693 (N_8693,N_5369,N_7994);
nand U8694 (N_8694,N_7093,N_7965);
or U8695 (N_8695,N_4946,N_4565);
and U8696 (N_8696,N_6251,N_5993);
nor U8697 (N_8697,N_7946,N_5202);
nand U8698 (N_8698,N_5204,N_6303);
nor U8699 (N_8699,N_7820,N_6834);
or U8700 (N_8700,N_4971,N_4719);
nand U8701 (N_8701,N_6102,N_5402);
nand U8702 (N_8702,N_7604,N_6200);
nor U8703 (N_8703,N_4921,N_7622);
or U8704 (N_8704,N_5942,N_5430);
nor U8705 (N_8705,N_7540,N_7066);
or U8706 (N_8706,N_6398,N_6568);
and U8707 (N_8707,N_7084,N_4091);
nand U8708 (N_8708,N_7335,N_6083);
or U8709 (N_8709,N_4867,N_5254);
or U8710 (N_8710,N_4037,N_5539);
nand U8711 (N_8711,N_4371,N_7107);
and U8712 (N_8712,N_4827,N_7073);
nor U8713 (N_8713,N_7484,N_7808);
or U8714 (N_8714,N_5867,N_7008);
nand U8715 (N_8715,N_5997,N_6891);
nand U8716 (N_8716,N_5241,N_5757);
or U8717 (N_8717,N_5544,N_6806);
and U8718 (N_8718,N_7446,N_4851);
nand U8719 (N_8719,N_7794,N_7769);
or U8720 (N_8720,N_4397,N_4847);
xnor U8721 (N_8721,N_7522,N_5068);
or U8722 (N_8722,N_4787,N_4875);
nand U8723 (N_8723,N_4828,N_4557);
nand U8724 (N_8724,N_5075,N_5945);
and U8725 (N_8725,N_5305,N_6487);
or U8726 (N_8726,N_4454,N_6088);
xnor U8727 (N_8727,N_4619,N_6245);
nor U8728 (N_8728,N_5702,N_7790);
xnor U8729 (N_8729,N_5134,N_5194);
and U8730 (N_8730,N_5614,N_7940);
nor U8731 (N_8731,N_4215,N_6405);
nor U8732 (N_8732,N_6587,N_6658);
xnor U8733 (N_8733,N_4074,N_5293);
or U8734 (N_8734,N_6502,N_7513);
nor U8735 (N_8735,N_7504,N_7830);
nor U8736 (N_8736,N_5849,N_5475);
and U8737 (N_8737,N_4675,N_4932);
xnor U8738 (N_8738,N_4857,N_5145);
nand U8739 (N_8739,N_6726,N_7468);
or U8740 (N_8740,N_4447,N_4165);
nand U8741 (N_8741,N_7320,N_6382);
nor U8742 (N_8742,N_5450,N_6617);
nand U8743 (N_8743,N_6565,N_6990);
or U8744 (N_8744,N_6689,N_4213);
nor U8745 (N_8745,N_4839,N_6333);
nand U8746 (N_8746,N_6469,N_6635);
and U8747 (N_8747,N_4403,N_6109);
xor U8748 (N_8748,N_6608,N_6491);
nor U8749 (N_8749,N_7402,N_7342);
nand U8750 (N_8750,N_7230,N_5200);
and U8751 (N_8751,N_7004,N_5114);
nor U8752 (N_8752,N_5761,N_7344);
nor U8753 (N_8753,N_4297,N_5653);
or U8754 (N_8754,N_5839,N_7824);
and U8755 (N_8755,N_6515,N_4802);
or U8756 (N_8756,N_5281,N_7333);
and U8757 (N_8757,N_4960,N_6590);
nor U8758 (N_8758,N_5511,N_7217);
and U8759 (N_8759,N_6890,N_5168);
nor U8760 (N_8760,N_5580,N_5953);
nor U8761 (N_8761,N_6431,N_5833);
or U8762 (N_8762,N_5600,N_7173);
and U8763 (N_8763,N_6878,N_4842);
and U8764 (N_8764,N_6953,N_6528);
nor U8765 (N_8765,N_7605,N_4727);
xor U8766 (N_8766,N_5533,N_5907);
xor U8767 (N_8767,N_6384,N_4916);
xnor U8768 (N_8768,N_5858,N_7491);
nand U8769 (N_8769,N_5678,N_5229);
or U8770 (N_8770,N_7662,N_5811);
nand U8771 (N_8771,N_7547,N_4536);
and U8772 (N_8772,N_4722,N_6280);
nand U8773 (N_8773,N_5530,N_4018);
xor U8774 (N_8774,N_6710,N_4273);
xnor U8775 (N_8775,N_6773,N_4206);
nor U8776 (N_8776,N_6649,N_4738);
nand U8777 (N_8777,N_5206,N_7739);
nand U8778 (N_8778,N_7551,N_5454);
and U8779 (N_8779,N_4029,N_7103);
nor U8780 (N_8780,N_4562,N_4468);
nor U8781 (N_8781,N_4514,N_4153);
nor U8782 (N_8782,N_5676,N_7370);
nor U8783 (N_8783,N_7077,N_6314);
xor U8784 (N_8784,N_7881,N_6345);
or U8785 (N_8785,N_5128,N_5872);
and U8786 (N_8786,N_7352,N_7748);
or U8787 (N_8787,N_6988,N_4175);
or U8788 (N_8788,N_7111,N_5681);
xnor U8789 (N_8789,N_6501,N_7834);
and U8790 (N_8790,N_7315,N_7959);
xor U8791 (N_8791,N_5005,N_6550);
nor U8792 (N_8792,N_7875,N_7322);
nor U8793 (N_8793,N_4441,N_5372);
and U8794 (N_8794,N_7124,N_5051);
nor U8795 (N_8795,N_7184,N_6204);
xnor U8796 (N_8796,N_7447,N_4524);
nor U8797 (N_8797,N_4453,N_4298);
nor U8798 (N_8798,N_7989,N_6777);
or U8799 (N_8799,N_4163,N_5480);
nand U8800 (N_8800,N_5895,N_7379);
nand U8801 (N_8801,N_6400,N_6676);
and U8802 (N_8802,N_7069,N_7404);
and U8803 (N_8803,N_4086,N_6611);
and U8804 (N_8804,N_5299,N_6402);
or U8805 (N_8805,N_4771,N_6855);
or U8806 (N_8806,N_4184,N_7334);
and U8807 (N_8807,N_4766,N_5557);
nor U8808 (N_8808,N_6330,N_7660);
xnor U8809 (N_8809,N_6362,N_7980);
nor U8810 (N_8810,N_4936,N_7767);
nor U8811 (N_8811,N_7086,N_7338);
nand U8812 (N_8812,N_4824,N_4167);
nand U8813 (N_8813,N_6064,N_5669);
and U8814 (N_8814,N_7406,N_5403);
and U8815 (N_8815,N_5724,N_5672);
or U8816 (N_8816,N_7425,N_6686);
and U8817 (N_8817,N_5593,N_7590);
nand U8818 (N_8818,N_4682,N_7855);
nor U8819 (N_8819,N_6124,N_7987);
nand U8820 (N_8820,N_6805,N_4657);
and U8821 (N_8821,N_4071,N_4923);
nor U8822 (N_8822,N_5711,N_7426);
or U8823 (N_8823,N_7456,N_7274);
nor U8824 (N_8824,N_6084,N_4721);
xor U8825 (N_8825,N_6435,N_5317);
or U8826 (N_8826,N_6320,N_4525);
nor U8827 (N_8827,N_4284,N_4858);
xor U8828 (N_8828,N_7827,N_7736);
xnor U8829 (N_8829,N_5657,N_6218);
nor U8830 (N_8830,N_4227,N_4677);
or U8831 (N_8831,N_5110,N_5658);
nor U8832 (N_8832,N_5853,N_4166);
or U8833 (N_8833,N_5651,N_6045);
xnor U8834 (N_8834,N_6545,N_4974);
and U8835 (N_8835,N_4558,N_7204);
or U8836 (N_8836,N_6311,N_7465);
nor U8837 (N_8837,N_7779,N_4174);
nand U8838 (N_8838,N_4040,N_5276);
nand U8839 (N_8839,N_4613,N_4967);
nand U8840 (N_8840,N_7000,N_5269);
nor U8841 (N_8841,N_6367,N_5691);
or U8842 (N_8842,N_7222,N_4185);
nor U8843 (N_8843,N_6960,N_5799);
or U8844 (N_8844,N_4793,N_5626);
nor U8845 (N_8845,N_5627,N_7726);
and U8846 (N_8846,N_7728,N_4120);
nor U8847 (N_8847,N_5662,N_5932);
and U8848 (N_8848,N_4368,N_4179);
and U8849 (N_8849,N_6429,N_6196);
nor U8850 (N_8850,N_4783,N_6068);
nand U8851 (N_8851,N_4429,N_5689);
and U8852 (N_8852,N_6335,N_7276);
nand U8853 (N_8853,N_7534,N_5242);
or U8854 (N_8854,N_5542,N_7229);
or U8855 (N_8855,N_5910,N_7482);
nor U8856 (N_8856,N_6105,N_6819);
or U8857 (N_8857,N_5578,N_6304);
or U8858 (N_8858,N_4542,N_4085);
nor U8859 (N_8859,N_5690,N_5150);
xor U8860 (N_8860,N_7058,N_6862);
nor U8861 (N_8861,N_7918,N_4679);
xor U8862 (N_8862,N_5708,N_4496);
nor U8863 (N_8863,N_7133,N_4052);
nand U8864 (N_8864,N_6657,N_5925);
or U8865 (N_8865,N_5146,N_4676);
or U8866 (N_8866,N_5096,N_5974);
and U8867 (N_8867,N_6851,N_6915);
nand U8868 (N_8868,N_7293,N_4111);
and U8869 (N_8869,N_7968,N_5687);
nand U8870 (N_8870,N_6443,N_7440);
and U8871 (N_8871,N_4532,N_7095);
xnor U8872 (N_8872,N_6745,N_6166);
or U8873 (N_8873,N_7331,N_7071);
xor U8874 (N_8874,N_5764,N_5851);
nand U8875 (N_8875,N_6106,N_6391);
xor U8876 (N_8876,N_7910,N_7244);
and U8877 (N_8877,N_6643,N_5756);
xnor U8878 (N_8878,N_6445,N_4689);
or U8879 (N_8879,N_5153,N_5389);
nor U8880 (N_8880,N_6116,N_4486);
or U8881 (N_8881,N_6863,N_6551);
xnor U8882 (N_8882,N_5783,N_5193);
nor U8883 (N_8883,N_4554,N_6926);
nand U8884 (N_8884,N_5722,N_4610);
nor U8885 (N_8885,N_4843,N_7325);
nand U8886 (N_8886,N_5618,N_6478);
nand U8887 (N_8887,N_5903,N_7758);
nand U8888 (N_8888,N_7610,N_5217);
nor U8889 (N_8889,N_7849,N_4854);
nor U8890 (N_8890,N_6327,N_6338);
and U8891 (N_8891,N_7218,N_6992);
nor U8892 (N_8892,N_4641,N_5017);
and U8893 (N_8893,N_5840,N_4030);
xnor U8894 (N_8894,N_5451,N_6464);
or U8895 (N_8895,N_6906,N_5906);
xnor U8896 (N_8896,N_6607,N_4961);
nor U8897 (N_8897,N_7811,N_7971);
nor U8898 (N_8898,N_7885,N_5798);
or U8899 (N_8899,N_6621,N_7983);
and U8900 (N_8900,N_4816,N_4012);
xnor U8901 (N_8901,N_4735,N_6830);
nand U8902 (N_8902,N_6262,N_5033);
nor U8903 (N_8903,N_7444,N_4977);
xnor U8904 (N_8904,N_5108,N_4233);
nor U8905 (N_8905,N_6393,N_7906);
nor U8906 (N_8906,N_4609,N_5421);
and U8907 (N_8907,N_5058,N_4622);
and U8908 (N_8908,N_5668,N_6781);
xor U8909 (N_8909,N_7896,N_6511);
or U8910 (N_8910,N_7992,N_5216);
and U8911 (N_8911,N_5896,N_4005);
xor U8912 (N_8912,N_7037,N_7716);
nand U8913 (N_8913,N_6387,N_5904);
xnor U8914 (N_8914,N_5769,N_5236);
xor U8915 (N_8915,N_4734,N_7266);
and U8916 (N_8916,N_5554,N_4549);
nand U8917 (N_8917,N_7061,N_5850);
xnor U8918 (N_8918,N_6169,N_4500);
nand U8919 (N_8919,N_4098,N_5999);
nand U8920 (N_8920,N_4141,N_6856);
nor U8921 (N_8921,N_5049,N_6647);
xor U8922 (N_8922,N_7189,N_4694);
xor U8923 (N_8923,N_5034,N_4398);
xor U8924 (N_8924,N_7052,N_6875);
and U8925 (N_8925,N_5105,N_7671);
and U8926 (N_8926,N_4036,N_4169);
or U8927 (N_8927,N_4102,N_7441);
and U8928 (N_8928,N_5989,N_4143);
nand U8929 (N_8929,N_7932,N_7177);
or U8930 (N_8930,N_7707,N_5334);
nor U8931 (N_8931,N_5021,N_4958);
nand U8932 (N_8932,N_4278,N_4951);
and U8933 (N_8933,N_4069,N_6995);
nand U8934 (N_8934,N_7083,N_6544);
xnor U8935 (N_8935,N_6945,N_7617);
xor U8936 (N_8936,N_4647,N_5482);
or U8937 (N_8937,N_4489,N_7161);
xor U8938 (N_8938,N_6836,N_4387);
nor U8939 (N_8939,N_5859,N_4599);
xnor U8940 (N_8940,N_4076,N_5196);
nand U8941 (N_8941,N_5062,N_5788);
or U8942 (N_8942,N_6027,N_7172);
nor U8943 (N_8943,N_5780,N_4156);
or U8944 (N_8944,N_7118,N_5847);
nor U8945 (N_8945,N_7022,N_4003);
nor U8946 (N_8946,N_6127,N_7515);
xnor U8947 (N_8947,N_6033,N_6812);
and U8948 (N_8948,N_6739,N_4869);
and U8949 (N_8949,N_4378,N_5927);
xnor U8950 (N_8950,N_7481,N_6267);
and U8951 (N_8951,N_5052,N_4126);
xnor U8952 (N_8952,N_5919,N_6816);
nand U8953 (N_8953,N_4887,N_4401);
nor U8954 (N_8954,N_6894,N_7007);
or U8955 (N_8955,N_6397,N_4577);
nor U8956 (N_8956,N_4658,N_5592);
nor U8957 (N_8957,N_7916,N_4582);
or U8958 (N_8958,N_6868,N_5513);
xnor U8959 (N_8959,N_4672,N_5428);
xnor U8960 (N_8960,N_6752,N_5632);
xor U8961 (N_8961,N_6738,N_5875);
or U8962 (N_8962,N_5319,N_6785);
and U8963 (N_8963,N_7563,N_6480);
xor U8964 (N_8964,N_7355,N_7778);
nand U8965 (N_8965,N_6673,N_4427);
or U8966 (N_8966,N_5584,N_6047);
nor U8967 (N_8967,N_4684,N_6270);
xnor U8968 (N_8968,N_5327,N_4853);
nor U8969 (N_8969,N_7486,N_6540);
and U8970 (N_8970,N_6804,N_4931);
nor U8971 (N_8971,N_6822,N_6691);
xnor U8972 (N_8972,N_6020,N_4423);
nor U8973 (N_8973,N_6567,N_5084);
nor U8974 (N_8974,N_6902,N_4674);
nor U8975 (N_8975,N_4241,N_5185);
nand U8976 (N_8976,N_6234,N_7776);
xnor U8977 (N_8977,N_4544,N_7658);
nand U8978 (N_8978,N_6780,N_5621);
and U8979 (N_8979,N_4723,N_6184);
or U8980 (N_8980,N_5151,N_5648);
nor U8981 (N_8981,N_5101,N_6958);
nor U8982 (N_8982,N_4782,N_7558);
nor U8983 (N_8983,N_6859,N_7892);
and U8984 (N_8984,N_4513,N_4511);
or U8985 (N_8985,N_6943,N_6427);
xor U8986 (N_8986,N_6562,N_4790);
xor U8987 (N_8987,N_7895,N_5968);
and U8988 (N_8988,N_5025,N_6485);
xor U8989 (N_8989,N_6056,N_6013);
xor U8990 (N_8990,N_7917,N_4326);
and U8991 (N_8991,N_4232,N_7392);
nor U8992 (N_8992,N_6294,N_6114);
nor U8993 (N_8993,N_6904,N_4257);
nor U8994 (N_8994,N_7943,N_4408);
nor U8995 (N_8995,N_6477,N_6857);
or U8996 (N_8996,N_7582,N_7870);
xor U8997 (N_8997,N_7775,N_4376);
nand U8998 (N_8998,N_6933,N_7341);
and U8999 (N_8999,N_6472,N_5759);
and U9000 (N_9000,N_4127,N_4266);
nand U9001 (N_9001,N_7713,N_5427);
xor U9002 (N_9002,N_5492,N_6623);
xor U9003 (N_9003,N_5144,N_7511);
nand U9004 (N_9004,N_6031,N_6399);
nand U9005 (N_9005,N_4881,N_7999);
nor U9006 (N_9006,N_7615,N_6484);
or U9007 (N_9007,N_6641,N_5385);
or U9008 (N_9008,N_6042,N_5961);
or U9009 (N_9009,N_4189,N_7208);
and U9010 (N_9010,N_5489,N_7815);
nand U9011 (N_9011,N_5419,N_5873);
and U9012 (N_9012,N_7854,N_6434);
nand U9013 (N_9013,N_5170,N_5634);
xor U9014 (N_9014,N_4106,N_7927);
and U9015 (N_9015,N_7606,N_7734);
xor U9016 (N_9016,N_7421,N_6901);
xnor U9017 (N_9017,N_4134,N_7492);
nor U9018 (N_9018,N_6642,N_5376);
and U9019 (N_9019,N_4935,N_4451);
and U9020 (N_9020,N_7800,N_7869);
and U9021 (N_9021,N_4980,N_7194);
or U9022 (N_9022,N_6066,N_6981);
and U9023 (N_9023,N_7942,N_4104);
nor U9024 (N_9024,N_6849,N_5102);
nor U9025 (N_9025,N_7589,N_7956);
nor U9026 (N_9026,N_5710,N_5160);
xnor U9027 (N_9027,N_7340,N_4550);
nand U9028 (N_9028,N_5921,N_7520);
nor U9029 (N_9029,N_7489,N_4026);
nor U9030 (N_9030,N_7450,N_5413);
xor U9031 (N_9031,N_7925,N_6444);
nand U9032 (N_9032,N_5434,N_7264);
and U9033 (N_9033,N_5011,N_6931);
and U9034 (N_9034,N_4180,N_6883);
or U9035 (N_9035,N_6910,N_5436);
nand U9036 (N_9036,N_5913,N_7175);
or U9037 (N_9037,N_7297,N_4592);
and U9038 (N_9038,N_6396,N_6470);
or U9039 (N_9039,N_5909,N_7764);
and U9040 (N_9040,N_5407,N_4556);
or U9041 (N_9041,N_4115,N_6826);
nand U9042 (N_9042,N_7296,N_6779);
or U9043 (N_9043,N_6599,N_7198);
xor U9044 (N_9044,N_4306,N_4724);
and U9045 (N_9045,N_5717,N_5861);
xor U9046 (N_9046,N_6887,N_6999);
or U9047 (N_9047,N_5043,N_4119);
nor U9048 (N_9048,N_4795,N_7011);
xor U9049 (N_9049,N_7756,N_6317);
or U9050 (N_9050,N_6244,N_7226);
and U9051 (N_9051,N_6841,N_7858);
nand U9052 (N_9052,N_4669,N_4726);
or U9053 (N_9053,N_6243,N_5004);
nand U9054 (N_9054,N_6392,N_5504);
nand U9055 (N_9055,N_7623,N_5640);
and U9056 (N_9056,N_6766,N_5892);
xor U9057 (N_9057,N_7634,N_5663);
and U9058 (N_9058,N_5595,N_7146);
xor U9059 (N_9059,N_6173,N_7501);
nand U9060 (N_9060,N_4020,N_4983);
nand U9061 (N_9061,N_5844,N_7381);
or U9062 (N_9062,N_6430,N_5177);
nor U9063 (N_9063,N_7792,N_7036);
or U9064 (N_9064,N_7783,N_4187);
xor U9065 (N_9065,N_4567,N_7818);
xor U9066 (N_9066,N_7805,N_4813);
xnor U9067 (N_9067,N_6719,N_6111);
and U9068 (N_9068,N_6730,N_4114);
nand U9069 (N_9069,N_4426,N_4415);
nand U9070 (N_9070,N_5568,N_6605);
xor U9071 (N_9071,N_6873,N_4708);
and U9072 (N_9072,N_6554,N_4534);
xnor U9073 (N_9073,N_7600,N_4407);
xor U9074 (N_9074,N_6250,N_4555);
nand U9075 (N_9075,N_4640,N_5984);
and U9076 (N_9076,N_4897,N_4700);
nand U9077 (N_9077,N_5623,N_6040);
xor U9078 (N_9078,N_7434,N_7137);
nand U9079 (N_9079,N_6016,N_6128);
nand U9080 (N_9080,N_7463,N_6374);
and U9081 (N_9081,N_4370,N_4670);
nor U9082 (N_9082,N_7104,N_4548);
nor U9083 (N_9083,N_6734,N_4234);
xnor U9084 (N_9084,N_5900,N_4861);
or U9085 (N_9085,N_7823,N_6889);
nor U9086 (N_9086,N_7292,N_5954);
and U9087 (N_9087,N_7641,N_7781);
xor U9088 (N_9088,N_6674,N_5460);
nand U9089 (N_9089,N_7519,N_5022);
nand U9090 (N_9090,N_7224,N_4944);
xnor U9091 (N_9091,N_4778,N_4581);
xor U9092 (N_9092,N_4290,N_7653);
nand U9093 (N_9093,N_7907,N_5054);
nand U9094 (N_9094,N_4806,N_4469);
xor U9095 (N_9095,N_6729,N_4844);
nor U9096 (N_9096,N_5787,N_4506);
or U9097 (N_9097,N_5514,N_4494);
nor U9098 (N_9098,N_4466,N_4258);
nor U9099 (N_9099,N_5804,N_6662);
or U9100 (N_9100,N_5394,N_4445);
and U9101 (N_9101,N_6140,N_4072);
xor U9102 (N_9102,N_7010,N_7429);
and U9103 (N_9103,N_7431,N_6165);
or U9104 (N_9104,N_5337,N_5086);
nor U9105 (N_9105,N_5755,N_7207);
nand U9106 (N_9106,N_7602,N_7400);
or U9107 (N_9107,N_7941,N_5800);
or U9108 (N_9108,N_4699,N_5686);
nand U9109 (N_9109,N_5228,N_7761);
nor U9110 (N_9110,N_7839,N_4900);
xor U9111 (N_9111,N_6239,N_5341);
or U9112 (N_9112,N_7261,N_5951);
and U9113 (N_9113,N_7414,N_6938);
xnor U9114 (N_9114,N_7196,N_7289);
nand U9115 (N_9115,N_7079,N_5987);
or U9116 (N_9116,N_6142,N_7454);
nor U9117 (N_9117,N_5526,N_6077);
xnor U9118 (N_9118,N_4933,N_6110);
and U9119 (N_9119,N_7717,N_6764);
and U9120 (N_9120,N_4087,N_6035);
xor U9121 (N_9121,N_6009,N_6370);
nand U9122 (N_9122,N_4574,N_5569);
xnor U9123 (N_9123,N_4987,N_6439);
or U9124 (N_9124,N_6366,N_5207);
nand U9125 (N_9125,N_4242,N_5943);
xor U9126 (N_9126,N_6509,N_4635);
nor U9127 (N_9127,N_7709,N_7200);
nand U9128 (N_9128,N_7459,N_4483);
or U9129 (N_9129,N_5767,N_4001);
xnor U9130 (N_9130,N_4600,N_7388);
nor U9131 (N_9131,N_6508,N_4995);
nand U9132 (N_9132,N_5778,N_5088);
and U9133 (N_9133,N_4260,N_5393);
nor U9134 (N_9134,N_4910,N_5822);
nor U9135 (N_9135,N_6973,N_7498);
and U9136 (N_9136,N_6740,N_7901);
nand U9137 (N_9137,N_6407,N_7225);
and U9138 (N_9138,N_4546,N_4688);
or U9139 (N_9139,N_4093,N_6754);
and U9140 (N_9140,N_5536,N_7360);
xor U9141 (N_9141,N_5082,N_7851);
nand U9142 (N_9142,N_4712,N_5829);
or U9143 (N_9143,N_7595,N_6059);
xnor U9144 (N_9144,N_6495,N_7976);
or U9145 (N_9145,N_6944,N_7990);
nand U9146 (N_9146,N_5330,N_6620);
or U9147 (N_9147,N_5028,N_5320);
nand U9148 (N_9148,N_5499,N_7557);
xnor U9149 (N_9149,N_7692,N_4034);
nor U9150 (N_9150,N_7867,N_7777);
xor U9151 (N_9151,N_7182,N_7391);
and U9152 (N_9152,N_7128,N_5212);
nand U9153 (N_9153,N_6319,N_5899);
or U9154 (N_9154,N_7898,N_5476);
and U9155 (N_9155,N_5268,N_7666);
or U9156 (N_9156,N_6709,N_4457);
and U9157 (N_9157,N_7737,N_6428);
xor U9158 (N_9158,N_5741,N_6758);
or U9159 (N_9159,N_7847,N_6622);
nor U9160 (N_9160,N_5310,N_4872);
nor U9161 (N_9161,N_4736,N_6886);
nand U9162 (N_9162,N_6613,N_6206);
or U9163 (N_9163,N_4251,N_7397);
xor U9164 (N_9164,N_6929,N_7351);
nand U9165 (N_9165,N_7838,N_5308);
or U9166 (N_9166,N_6576,N_4817);
nor U9167 (N_9167,N_7712,N_4878);
or U9168 (N_9168,N_4027,N_6975);
or U9169 (N_9169,N_6525,N_6840);
nand U9170 (N_9170,N_6921,N_4367);
and U9171 (N_9171,N_5494,N_5180);
nor U9172 (N_9172,N_4826,N_6594);
nand U9173 (N_9173,N_6312,N_7974);
xnor U9174 (N_9174,N_5507,N_6940);
or U9175 (N_9175,N_7363,N_4835);
nand U9176 (N_9176,N_6375,N_4428);
or U9177 (N_9177,N_5760,N_6670);
xnor U9178 (N_9178,N_6104,N_7178);
nor U9179 (N_9179,N_4792,N_4042);
nand U9180 (N_9180,N_6275,N_4696);
or U9181 (N_9181,N_7735,N_6252);
nand U9182 (N_9182,N_7575,N_5371);
nor U9183 (N_9183,N_6103,N_6757);
and U9184 (N_9184,N_7114,N_5608);
nor U9185 (N_9185,N_7428,N_6632);
and U9186 (N_9186,N_5963,N_7451);
xor U9187 (N_9187,N_6510,N_5891);
and U9188 (N_9188,N_5729,N_5863);
and U9189 (N_9189,N_6690,N_5782);
and U9190 (N_9190,N_7369,N_4230);
and U9191 (N_9191,N_6113,N_5098);
or U9192 (N_9192,N_7330,N_5843);
or U9193 (N_9193,N_7788,N_4575);
nand U9194 (N_9194,N_6422,N_5415);
and U9195 (N_9195,N_5203,N_7760);
nand U9196 (N_9196,N_4433,N_5423);
nand U9197 (N_9197,N_6411,N_7203);
and U9198 (N_9198,N_6570,N_4252);
xor U9199 (N_9199,N_4812,N_5862);
nand U9200 (N_9200,N_6067,N_6496);
or U9201 (N_9201,N_5332,N_7399);
xnor U9202 (N_9202,N_7500,N_7163);
nand U9203 (N_9203,N_7935,N_6448);
xor U9204 (N_9204,N_5173,N_5328);
and U9205 (N_9205,N_4384,N_7057);
xor U9206 (N_9206,N_7607,N_6079);
nand U9207 (N_9207,N_7508,N_6050);
and U9208 (N_9208,N_7027,N_5918);
xnor U9209 (N_9209,N_5031,N_7929);
and U9210 (N_9210,N_7117,N_5148);
xor U9211 (N_9211,N_7306,N_4988);
or U9212 (N_9212,N_7612,N_7844);
nand U9213 (N_9213,N_7742,N_5478);
xnor U9214 (N_9214,N_5059,N_6232);
nand U9215 (N_9215,N_7195,N_6972);
nor U9216 (N_9216,N_6026,N_5237);
xnor U9217 (N_9217,N_4044,N_4911);
nor U9218 (N_9218,N_4317,N_7969);
xor U9219 (N_9219,N_5390,N_4994);
xor U9220 (N_9220,N_6229,N_4279);
nor U9221 (N_9221,N_4053,N_5649);
nor U9222 (N_9222,N_5934,N_7809);
and U9223 (N_9223,N_5155,N_5479);
nand U9224 (N_9224,N_6900,N_5099);
and U9225 (N_9225,N_4123,N_4889);
and U9226 (N_9226,N_7162,N_5571);
xnor U9227 (N_9227,N_6268,N_6583);
or U9228 (N_9228,N_6416,N_4479);
or U9229 (N_9229,N_6326,N_4698);
nand U9230 (N_9230,N_7789,N_7580);
nor U9231 (N_9231,N_6736,N_7223);
xor U9232 (N_9232,N_5619,N_7806);
xnor U9233 (N_9233,N_7304,N_4519);
nor U9234 (N_9234,N_7638,N_5758);
and U9235 (N_9235,N_4133,N_5924);
xnor U9236 (N_9236,N_4391,N_4801);
nor U9237 (N_9237,N_7863,N_5001);
and U9238 (N_9238,N_6323,N_7153);
nor U9239 (N_9239,N_7423,N_4400);
nand U9240 (N_9240,N_7897,N_4217);
and U9241 (N_9241,N_5267,N_5361);
xnor U9242 (N_9242,N_4435,N_4263);
xnor U9243 (N_9243,N_5996,N_6351);
nor U9244 (N_9244,N_6217,N_6817);
xor U9245 (N_9245,N_4798,N_7485);
and U9246 (N_9246,N_5827,N_6678);
nor U9247 (N_9247,N_7802,N_7197);
and U9248 (N_9248,N_7257,N_5886);
or U9249 (N_9249,N_5181,N_7587);
nor U9250 (N_9250,N_4443,N_4907);
and U9251 (N_9251,N_7288,N_4841);
and U9252 (N_9252,N_4810,N_4618);
xor U9253 (N_9253,N_6526,N_6256);
xnor U9254 (N_9254,N_4222,N_4968);
xor U9255 (N_9255,N_4430,N_6982);
or U9256 (N_9256,N_5792,N_7160);
xnor U9257 (N_9257,N_7099,N_7561);
nor U9258 (N_9258,N_7272,N_6343);
nor U9259 (N_9259,N_4780,N_7714);
nor U9260 (N_9260,N_4940,N_6803);
xnor U9261 (N_9261,N_5159,N_5775);
or U9262 (N_9262,N_6221,N_5422);
xor U9263 (N_9263,N_4879,N_4666);
nand U9264 (N_9264,N_7006,N_4314);
xor U9265 (N_9265,N_6154,N_7559);
nand U9266 (N_9266,N_5739,N_4319);
and U9267 (N_9267,N_6713,N_4616);
or U9268 (N_9268,N_6820,N_4632);
or U9269 (N_9269,N_5013,N_6714);
or U9270 (N_9270,N_4838,N_4181);
xor U9271 (N_9271,N_7588,N_4701);
and U9272 (N_9272,N_4898,N_5809);
xor U9273 (N_9273,N_5633,N_4773);
or U9274 (N_9274,N_7537,N_5620);
and U9275 (N_9275,N_4157,N_7890);
or U9276 (N_9276,N_6581,N_7903);
and U9277 (N_9277,N_6930,N_4860);
nand U9278 (N_9278,N_7076,N_7997);
and U9279 (N_9279,N_7043,N_7798);
and U9280 (N_9280,N_4779,N_5803);
and U9281 (N_9281,N_6225,N_4762);
xor U9282 (N_9282,N_7055,N_5723);
nand U9283 (N_9283,N_6839,N_7329);
nor U9284 (N_9284,N_5939,N_4048);
nor U9285 (N_9285,N_5878,N_4985);
nor U9286 (N_9286,N_4136,N_6361);
nand U9287 (N_9287,N_7759,N_5736);
xnor U9288 (N_9288,N_5692,N_6541);
nor U9289 (N_9289,N_5725,N_4325);
nor U9290 (N_9290,N_7436,N_7936);
and U9291 (N_9291,N_5730,N_4356);
nand U9292 (N_9292,N_6920,N_5095);
nor U9293 (N_9293,N_6197,N_6655);
xor U9294 (N_9294,N_5414,N_7833);
xnor U9295 (N_9295,N_7171,N_6619);
nand U9296 (N_9296,N_4834,N_4667);
or U9297 (N_9297,N_6328,N_6778);
xnor U9298 (N_9298,N_4580,N_4587);
or U9299 (N_9299,N_5864,N_4062);
xor U9300 (N_9300,N_6530,N_4406);
or U9301 (N_9301,N_6814,N_4509);
and U9302 (N_9302,N_5773,N_6019);
nand U9303 (N_9303,N_7255,N_6024);
nand U9304 (N_9304,N_7920,N_6917);
nand U9305 (N_9305,N_6786,N_5316);
xor U9306 (N_9306,N_6350,N_6004);
nor U9307 (N_9307,N_5169,N_6028);
nor U9308 (N_9308,N_5359,N_7152);
nand U9309 (N_9309,N_4323,N_6034);
xor U9310 (N_9310,N_6936,N_6783);
xor U9311 (N_9311,N_7923,N_4437);
nand U9312 (N_9312,N_4865,N_6060);
and U9313 (N_9313,N_7931,N_4709);
xor U9314 (N_9314,N_7635,N_7574);
and U9315 (N_9315,N_5624,N_7655);
or U9316 (N_9316,N_5848,N_6131);
or U9317 (N_9317,N_6386,N_6089);
nor U9318 (N_9318,N_4660,N_5820);
xor U9319 (N_9319,N_5354,N_5802);
and U9320 (N_9320,N_6724,N_5081);
and U9321 (N_9321,N_5671,N_7554);
nand U9322 (N_9322,N_7780,N_6589);
xnor U9323 (N_9323,N_7578,N_7659);
or U9324 (N_9324,N_7471,N_7215);
or U9325 (N_9325,N_6760,N_5887);
xor U9326 (N_9326,N_6627,N_4928);
nor U9327 (N_9327,N_6746,N_4631);
nor U9328 (N_9328,N_6650,N_7013);
and U9329 (N_9329,N_6138,N_7074);
or U9330 (N_9330,N_5381,N_5462);
and U9331 (N_9331,N_6467,N_5762);
nor U9332 (N_9332,N_4375,N_5652);
and U9333 (N_9333,N_4934,N_6874);
or U9334 (N_9334,N_6694,N_4570);
nor U9335 (N_9335,N_6473,N_5981);
nor U9336 (N_9336,N_5738,N_4703);
and U9337 (N_9337,N_6653,N_5468);
and U9338 (N_9338,N_4004,N_4269);
or U9339 (N_9339,N_6796,N_7393);
nor U9340 (N_9340,N_5547,N_7068);
nand U9341 (N_9341,N_6141,N_5625);
nor U9342 (N_9342,N_5195,N_5238);
xnor U9343 (N_9343,N_4748,N_7825);
and U9344 (N_9344,N_6161,N_4836);
nor U9345 (N_9345,N_4475,N_4975);
xor U9346 (N_9346,N_4776,N_4964);
or U9347 (N_9347,N_7228,N_7090);
nor U9348 (N_9348,N_7657,N_5087);
xor U9349 (N_9349,N_4832,N_4395);
xnor U9350 (N_9350,N_4757,N_4416);
or U9351 (N_9351,N_5597,N_4345);
nand U9352 (N_9352,N_6717,N_7151);
nand U9353 (N_9353,N_4014,N_4981);
xor U9354 (N_9354,N_7038,N_6438);
nand U9355 (N_9355,N_7199,N_7801);
and U9356 (N_9356,N_4612,N_4786);
and U9357 (N_9357,N_5467,N_5387);
and U9358 (N_9358,N_6007,N_7110);
and U9359 (N_9359,N_6030,N_6582);
xor U9360 (N_9360,N_4421,N_5149);
and U9361 (N_9361,N_7051,N_5541);
or U9362 (N_9362,N_4363,N_6247);
and U9363 (N_9363,N_4332,N_5599);
and U9364 (N_9364,N_4480,N_4248);
and U9365 (N_9365,N_5141,N_6286);
nor U9366 (N_9366,N_6606,N_6178);
xnor U9367 (N_9367,N_7981,N_6835);
xnor U9368 (N_9368,N_6970,N_5474);
or U9369 (N_9369,N_4409,N_6282);
nand U9370 (N_9370,N_4274,N_5313);
xor U9371 (N_9371,N_4602,N_7721);
xor U9372 (N_9372,N_7543,N_6770);
nand U9373 (N_9373,N_6610,N_7186);
nor U9374 (N_9374,N_4155,N_6249);
nor U9375 (N_9375,N_5429,N_4731);
nand U9376 (N_9376,N_5616,N_5103);
and U9377 (N_9377,N_7242,N_6115);
and U9378 (N_9378,N_6913,N_5466);
nor U9379 (N_9379,N_4892,N_6776);
nor U9380 (N_9380,N_5286,N_6654);
or U9381 (N_9381,N_7702,N_5503);
or U9382 (N_9382,N_7900,N_5824);
xnor U9383 (N_9383,N_6238,N_4906);
and U9384 (N_9384,N_7348,N_4303);
nor U9385 (N_9385,N_5014,N_6226);
nor U9386 (N_9386,N_5323,N_4051);
nand U9387 (N_9387,N_6548,N_4214);
or U9388 (N_9388,N_4563,N_4343);
xnor U9389 (N_9389,N_5116,N_7430);
xor U9390 (N_9390,N_4473,N_4759);
or U9391 (N_9391,N_7211,N_6888);
and U9392 (N_9392,N_5991,N_7321);
or U9393 (N_9393,N_5126,N_4741);
nand U9394 (N_9394,N_6788,N_5166);
and U9395 (N_9395,N_7514,N_7302);
or U9396 (N_9396,N_4791,N_5613);
xnor U9397 (N_9397,N_6306,N_7474);
or U9398 (N_9398,N_6230,N_7614);
or U9399 (N_9399,N_7462,N_6301);
nor U9400 (N_9400,N_6098,N_7260);
xnor U9401 (N_9401,N_7706,N_4081);
nand U9402 (N_9402,N_6457,N_7782);
nor U9403 (N_9403,N_6211,N_5879);
nor U9404 (N_9404,N_4768,N_4197);
nand U9405 (N_9405,N_4710,N_5285);
nand U9406 (N_9406,N_7619,N_7249);
xor U9407 (N_9407,N_4490,N_5139);
nand U9408 (N_9408,N_7784,N_7496);
xnor U9409 (N_9409,N_7240,N_4920);
xnor U9410 (N_9410,N_7168,N_4568);
nand U9411 (N_9411,N_4561,N_6700);
or U9412 (N_9412,N_7140,N_7365);
nand U9413 (N_9413,N_6912,N_6845);
or U9414 (N_9414,N_5384,N_7313);
nand U9415 (N_9415,N_4000,N_6728);
and U9416 (N_9416,N_4501,N_7343);
nand U9417 (N_9417,N_4926,N_4355);
nand U9418 (N_9418,N_4991,N_5388);
nand U9419 (N_9419,N_5223,N_5278);
or U9420 (N_9420,N_6549,N_5941);
or U9421 (N_9421,N_4372,N_4099);
nand U9422 (N_9422,N_5275,N_7419);
xnor U9423 (N_9423,N_6488,N_7683);
xor U9424 (N_9424,N_6117,N_6827);
nand U9425 (N_9425,N_6720,N_5555);
and U9426 (N_9426,N_6916,N_6597);
or U9427 (N_9427,N_4970,N_7210);
nor U9428 (N_9428,N_4998,N_6579);
or U9429 (N_9429,N_7831,N_7993);
or U9430 (N_9430,N_7049,N_4831);
nor U9431 (N_9431,N_6170,N_6666);
xnor U9432 (N_9432,N_4856,N_7608);
or U9433 (N_9433,N_4116,N_4359);
xor U9434 (N_9434,N_6531,N_5383);
and U9435 (N_9435,N_7668,N_4623);
nand U9436 (N_9436,N_4344,N_7385);
nor U9437 (N_9437,N_4884,N_5715);
xnor U9438 (N_9438,N_7220,N_5465);
xnor U9439 (N_9439,N_6539,N_6044);
nand U9440 (N_9440,N_6807,N_5259);
xor U9441 (N_9441,N_7814,N_4154);
xnor U9442 (N_9442,N_5481,N_7949);
and U9443 (N_9443,N_7349,N_4138);
and U9444 (N_9444,N_5695,N_5154);
or U9445 (N_9445,N_6193,N_6219);
nor U9446 (N_9446,N_7192,N_6652);
and U9447 (N_9447,N_7661,N_5189);
and U9448 (N_9448,N_4715,N_7643);
nand U9449 (N_9449,N_4285,N_6537);
xnor U9450 (N_9450,N_6998,N_7307);
nor U9451 (N_9451,N_7488,N_4800);
xnor U9452 (N_9452,N_6561,N_6672);
nand U9453 (N_9453,N_7596,N_6119);
nor U9454 (N_9454,N_4589,N_5506);
xnor U9455 (N_9455,N_5343,N_4761);
or U9456 (N_9456,N_4693,N_5060);
and U9457 (N_9457,N_7924,N_7960);
nand U9458 (N_9458,N_6481,N_5581);
xor U9459 (N_9459,N_4465,N_7873);
and U9460 (N_9460,N_6761,N_5573);
nand U9461 (N_9461,N_5808,N_7145);
xor U9462 (N_9462,N_6566,N_6403);
nand U9463 (N_9463,N_5486,N_7640);
or U9464 (N_9464,N_5039,N_4436);
nor U9465 (N_9465,N_7155,N_6003);
or U9466 (N_9466,N_6914,N_4603);
xor U9467 (N_9467,N_4105,N_6383);
or U9468 (N_9468,N_4286,N_5720);
nand U9469 (N_9469,N_4925,N_5104);
and U9470 (N_9470,N_6076,N_6475);
nor U9471 (N_9471,N_6512,N_7033);
xnor U9472 (N_9472,N_4212,N_7409);
nor U9473 (N_9473,N_7149,N_5665);
nor U9474 (N_9474,N_4785,N_6466);
nand U9475 (N_9475,N_6152,N_5035);
nand U9476 (N_9476,N_4440,N_5517);
or U9477 (N_9477,N_7545,N_5560);
nor U9478 (N_9478,N_7570,N_5041);
and U9479 (N_9479,N_7727,N_6061);
xor U9480 (N_9480,N_7265,N_7346);
xnor U9481 (N_9481,N_4893,N_5209);
or U9482 (N_9482,N_4733,N_7285);
nand U9483 (N_9483,N_6342,N_5493);
xor U9484 (N_9484,N_4767,N_5331);
nand U9485 (N_9485,N_4774,N_7050);
nor U9486 (N_9486,N_5452,N_4080);
and U9487 (N_9487,N_4392,N_4276);
nor U9488 (N_9488,N_4901,N_6364);
or U9489 (N_9489,N_7704,N_6479);
and U9490 (N_9490,N_4559,N_5551);
and U9491 (N_9491,N_7700,N_5766);
nor U9492 (N_9492,N_6160,N_5660);
xnor U9493 (N_9493,N_7390,N_5670);
and U9494 (N_9494,N_4402,N_7047);
xor U9495 (N_9495,N_6272,N_5130);
nand U9496 (N_9496,N_7665,N_5453);
or U9497 (N_9497,N_7291,N_5515);
and U9498 (N_9498,N_6222,N_7433);
nor U9499 (N_9499,N_5214,N_5846);
or U9500 (N_9500,N_7503,N_5463);
nor U9501 (N_9501,N_7142,N_4413);
xor U9502 (N_9502,N_6756,N_5659);
nor U9503 (N_9503,N_5400,N_4059);
or U9504 (N_9504,N_6001,N_4864);
xnor U9505 (N_9505,N_5210,N_7131);
and U9506 (N_9506,N_7725,N_6271);
nor U9507 (N_9507,N_5831,N_7461);
nand U9508 (N_9508,N_6440,N_4664);
and U9509 (N_9509,N_4484,N_6054);
xnor U9510 (N_9510,N_6381,N_6455);
nor U9511 (N_9511,N_6693,N_5333);
or U9512 (N_9512,N_7766,N_6183);
or U9513 (N_9513,N_5915,N_6927);
nand U9514 (N_9514,N_6552,N_6553);
nor U9515 (N_9515,N_7591,N_5117);
nand U9516 (N_9516,N_6494,N_4948);
nor U9517 (N_9517,N_7698,N_7193);
xor U9518 (N_9518,N_4740,N_7850);
xnor U9519 (N_9519,N_5157,N_4334);
or U9520 (N_9520,N_6722,N_5147);
nand U9521 (N_9521,N_4147,N_6514);
nand U9522 (N_9522,N_6955,N_6447);
nor U9523 (N_9523,N_7763,N_5498);
xor U9524 (N_9524,N_7670,N_7611);
nor U9525 (N_9525,N_4291,N_4661);
or U9526 (N_9526,N_6712,N_5261);
nor U9527 (N_9527,N_5211,N_6843);
or U9528 (N_9528,N_7532,N_4966);
or U9529 (N_9529,N_4137,N_6014);
and U9530 (N_9530,N_7147,N_6415);
nor U9531 (N_9531,N_4846,N_6144);
and U9532 (N_9532,N_7212,N_7132);
nor U9533 (N_9533,N_6207,N_5868);
nand U9534 (N_9534,N_5582,N_6101);
xnor U9535 (N_9535,N_4899,N_4503);
and U9536 (N_9536,N_5396,N_6205);
xor U9537 (N_9537,N_4282,N_6426);
and U9538 (N_9538,N_6497,N_6295);
or U9539 (N_9539,N_5807,N_4530);
xnor U9540 (N_9540,N_6185,N_5444);
or U9541 (N_9541,N_4348,N_5374);
nor U9542 (N_9542,N_5572,N_4010);
xnor U9543 (N_9543,N_4101,N_5930);
nand U9544 (N_9544,N_7516,N_7034);
nor U9545 (N_9545,N_7301,N_5816);
xnor U9546 (N_9546,N_4837,N_6237);
xor U9547 (N_9547,N_5357,N_7299);
and U9548 (N_9548,N_7250,N_6707);
nor U9549 (N_9549,N_5929,N_5959);
and U9550 (N_9550,N_6580,N_5488);
xor U9551 (N_9551,N_4784,N_4539);
or U9552 (N_9552,N_5456,N_6421);
xnor U9553 (N_9553,N_4862,N_6095);
or U9554 (N_9554,N_4097,N_4190);
nor U9555 (N_9555,N_5226,N_6636);
nand U9556 (N_9556,N_5699,N_4196);
and U9557 (N_9557,N_7368,N_6036);
nor U9558 (N_9558,N_5905,N_5184);
nor U9559 (N_9559,N_6872,N_6905);
xnor U9560 (N_9560,N_6420,N_5701);
nand U9561 (N_9561,N_4982,N_5302);
nand U9562 (N_9562,N_7202,N_5546);
nor U9563 (N_9563,N_6771,N_7620);
or U9564 (N_9564,N_7312,N_7856);
xor U9565 (N_9565,N_7269,N_4963);
xnor U9566 (N_9566,N_4377,N_4973);
xor U9567 (N_9567,N_6139,N_7676);
xnor U9568 (N_9568,N_5826,N_4794);
or U9569 (N_9569,N_5650,N_5890);
and U9570 (N_9570,N_6563,N_4361);
or U9571 (N_9571,N_5860,N_6162);
nor U9572 (N_9572,N_4320,N_4351);
nor U9573 (N_9573,N_7259,N_7394);
xnor U9574 (N_9574,N_4912,N_5250);
or U9575 (N_9575,N_5718,N_7654);
or U9576 (N_9576,N_6062,N_5029);
nand U9577 (N_9577,N_4205,N_4538);
and U9578 (N_9578,N_5164,N_4470);
or U9579 (N_9579,N_6334,N_4850);
and U9580 (N_9580,N_4245,N_4527);
nor U9581 (N_9581,N_5055,N_4695);
or U9582 (N_9582,N_5789,N_6747);
or U9583 (N_9583,N_7143,N_4903);
or U9584 (N_9584,N_5908,N_7323);
xnor U9585 (N_9585,N_4219,N_5754);
or U9586 (N_9586,N_6737,N_4930);
nor U9587 (N_9587,N_6151,N_7318);
xnor U9588 (N_9588,N_7020,N_6948);
nor U9589 (N_9589,N_5375,N_7319);
or U9590 (N_9590,N_7915,N_7377);
xnor U9591 (N_9591,N_5218,N_4041);
and U9592 (N_9592,N_6492,N_4908);
xor U9593 (N_9593,N_6869,N_6437);
nor U9594 (N_9594,N_7435,N_4653);
or U9595 (N_9595,N_7308,N_4112);
or U9596 (N_9596,N_7584,N_7876);
xnor U9597 (N_9597,N_7562,N_7785);
xnor U9598 (N_9598,N_7738,N_7797);
or U9599 (N_9599,N_6136,N_4535);
nand U9600 (N_9600,N_6175,N_5575);
nor U9601 (N_9601,N_7905,N_6842);
or U9602 (N_9602,N_6949,N_5696);
nand U9603 (N_9603,N_5877,N_5986);
xor U9604 (N_9604,N_6032,N_4047);
and U9605 (N_9605,N_5786,N_4883);
nand U9606 (N_9606,N_6523,N_4590);
nor U9607 (N_9607,N_7542,N_5882);
xor U9608 (N_9608,N_4108,N_7743);
or U9609 (N_9609,N_4598,N_5768);
nand U9610 (N_9610,N_4829,N_6818);
nand U9611 (N_9611,N_6521,N_5776);
and U9612 (N_9612,N_4625,N_5797);
nand U9613 (N_9613,N_4947,N_4337);
nor U9614 (N_9614,N_5420,N_4159);
nand U9615 (N_9615,N_7754,N_5885);
nand U9616 (N_9616,N_6645,N_6189);
and U9617 (N_9617,N_5604,N_4255);
and U9618 (N_9618,N_4396,N_5750);
xor U9619 (N_9619,N_5912,N_6199);
xor U9620 (N_9620,N_6522,N_7550);
or U9621 (N_9621,N_7651,N_7691);
and U9622 (N_9622,N_6248,N_5931);
or U9623 (N_9623,N_4192,N_7669);
nor U9624 (N_9624,N_4338,N_6592);
or U9625 (N_9625,N_6769,N_6322);
nand U9626 (N_9626,N_7424,N_7270);
and U9627 (N_9627,N_6821,N_5661);
or U9628 (N_9628,N_7339,N_7675);
or U9629 (N_9629,N_7552,N_7139);
nand U9630 (N_9630,N_4690,N_7252);
xor U9631 (N_9631,N_6146,N_4038);
or U9632 (N_9632,N_4476,N_7219);
nor U9633 (N_9633,N_6331,N_6733);
nor U9634 (N_9634,N_4585,N_6753);
and U9635 (N_9635,N_4442,N_6898);
xor U9636 (N_9636,N_4649,N_6041);
or U9637 (N_9637,N_7096,N_7089);
or U9638 (N_9638,N_5763,N_7205);
nand U9639 (N_9639,N_7967,N_5636);
or U9640 (N_9640,N_7478,N_4347);
and U9641 (N_9641,N_7082,N_4471);
and U9642 (N_9642,N_5874,N_6336);
nand U9643 (N_9643,N_6187,N_6784);
or U9644 (N_9644,N_7156,N_4758);
nor U9645 (N_9645,N_6517,N_5828);
nor U9646 (N_9646,N_7012,N_5352);
nand U9647 (N_9647,N_7248,N_6792);
and U9648 (N_9648,N_7986,N_5040);
nor U9649 (N_9649,N_4586,N_5719);
or U9650 (N_9650,N_5221,N_4803);
or U9651 (N_9651,N_4990,N_7473);
and U9652 (N_9652,N_6129,N_4805);
or U9653 (N_9653,N_6223,N_7416);
or U9654 (N_9654,N_4955,N_5418);
nor U9655 (N_9655,N_5852,N_6979);
and U9656 (N_9656,N_4021,N_4464);
nor U9657 (N_9657,N_6038,N_4130);
xor U9658 (N_9658,N_7072,N_5339);
nand U9659 (N_9659,N_7483,N_7191);
or U9660 (N_9660,N_7512,N_6388);
nand U9661 (N_9661,N_6751,N_6210);
nand U9662 (N_9662,N_5856,N_7791);
and U9663 (N_9663,N_4760,N_4596);
xnor U9664 (N_9664,N_4354,N_4663);
nand U9665 (N_9665,N_5733,N_5373);
nand U9666 (N_9666,N_5980,N_4431);
and U9667 (N_9667,N_6212,N_4404);
nor U9668 (N_9668,N_4969,N_4477);
and U9669 (N_9669,N_4651,N_6073);
xnor U9670 (N_9670,N_6735,N_4450);
nand U9671 (N_9671,N_5995,N_7411);
and U9672 (N_9672,N_5297,N_7382);
nand U9673 (N_9673,N_7387,N_6825);
or U9674 (N_9674,N_6516,N_4200);
nor U9675 (N_9675,N_5424,N_5295);
nand U9676 (N_9676,N_7822,N_7928);
xnor U9677 (N_9677,N_6997,N_7347);
and U9678 (N_9678,N_5698,N_6010);
or U9679 (N_9679,N_6143,N_5967);
or U9680 (N_9680,N_7832,N_7280);
nand U9681 (N_9681,N_6093,N_7979);
xor U9682 (N_9682,N_5893,N_5063);
nor U9683 (N_9683,N_4148,N_5069);
nor U9684 (N_9684,N_7125,N_7650);
or U9685 (N_9685,N_5038,N_4362);
xor U9686 (N_9686,N_4752,N_7278);
xor U9687 (N_9687,N_7018,N_4075);
xnor U9688 (N_9688,N_5314,N_7699);
or U9689 (N_9689,N_6795,N_4158);
xnor U9690 (N_9690,N_4770,N_5845);
or U9691 (N_9691,N_6947,N_5753);
and U9692 (N_9692,N_4487,N_5053);
xor U9693 (N_9693,N_6615,N_6265);
xor U9694 (N_9694,N_4256,N_4823);
or U9695 (N_9695,N_4434,N_6640);
xnor U9696 (N_9696,N_5304,N_6147);
nor U9697 (N_9697,N_5290,N_7807);
nor U9698 (N_9698,N_6591,N_5629);
or U9699 (N_9699,N_5010,N_5855);
or U9700 (N_9700,N_5596,N_7648);
nor U9701 (N_9701,N_5540,N_6911);
xor U9702 (N_9702,N_4997,N_5065);
xor U9703 (N_9703,N_5123,N_7626);
xnor U9704 (N_9704,N_7157,N_7652);
and U9705 (N_9705,N_4335,N_5794);
nor U9706 (N_9706,N_5279,N_7719);
xnor U9707 (N_9707,N_5510,N_6723);
nand U9708 (N_9708,N_5122,N_6118);
nor U9709 (N_9709,N_5774,N_5491);
nor U9710 (N_9710,N_6831,N_5135);
xnor U9711 (N_9711,N_7410,N_5391);
nand U9712 (N_9712,N_7238,N_5866);
xor U9713 (N_9713,N_5253,N_4945);
or U9714 (N_9714,N_4129,N_4113);
nor U9715 (N_9715,N_7644,N_5709);
and U9716 (N_9716,N_6002,N_7592);
and U9717 (N_9717,N_4642,N_4478);
nor U9718 (N_9718,N_5548,N_6684);
nor U9719 (N_9719,N_4820,N_5565);
and U9720 (N_9720,N_7639,N_7135);
and U9721 (N_9721,N_6284,N_4607);
or U9722 (N_9722,N_7772,N_6316);
xnor U9723 (N_9723,N_6190,N_5118);
nor U9724 (N_9724,N_4339,N_6281);
xnor U9725 (N_9725,N_5585,N_5950);
or U9726 (N_9726,N_5559,N_5495);
nand U9727 (N_9727,N_5284,N_4178);
nor U9728 (N_9728,N_4390,N_4579);
or U9729 (N_9729,N_4315,N_7376);
and U9730 (N_9730,N_4330,N_7751);
nand U9731 (N_9731,N_5965,N_4032);
and U9732 (N_9732,N_5656,N_7024);
or U9733 (N_9733,N_5458,N_7729);
nor U9734 (N_9734,N_7601,N_4272);
xnor U9735 (N_9735,N_4957,N_5312);
nor U9736 (N_9736,N_5440,N_4299);
nor U9737 (N_9737,N_4275,N_4249);
xor U9738 (N_9738,N_4082,N_7954);
nor U9739 (N_9739,N_4811,N_4237);
or U9740 (N_9740,N_5588,N_4019);
xor U9741 (N_9741,N_4056,N_4999);
and U9742 (N_9742,N_5880,N_7183);
or U9743 (N_9743,N_7078,N_6774);
xnor U9744 (N_9744,N_4924,N_6337);
xor U9745 (N_9745,N_6094,N_7138);
nand U9746 (N_9746,N_4769,N_4706);
nand U9747 (N_9747,N_4100,N_5042);
nand U9748 (N_9748,N_7420,N_7040);
xor U9749 (N_9749,N_4152,N_4756);
nor U9750 (N_9750,N_7599,N_5737);
nand U9751 (N_9751,N_4462,N_5007);
and U9752 (N_9752,N_4584,N_7030);
or U9753 (N_9753,N_6134,N_5777);
nand U9754 (N_9754,N_4687,N_6809);
or U9755 (N_9755,N_7170,N_4240);
or U9756 (N_9756,N_7884,N_7829);
or U9757 (N_9757,N_5806,N_7899);
and U9758 (N_9758,N_4611,N_4146);
nand U9759 (N_9759,N_5315,N_6907);
or U9760 (N_9760,N_7336,N_7982);
nand U9761 (N_9761,N_7846,N_5842);
and U9762 (N_9762,N_7879,N_7952);
or U9763 (N_9763,N_4753,N_7475);
nor U9764 (N_9764,N_5745,N_7693);
nand U9765 (N_9765,N_7848,N_7380);
xnor U9766 (N_9766,N_5471,N_6122);
nor U9767 (N_9767,N_7309,N_4045);
xnor U9768 (N_9768,N_5220,N_4614);
nand U9769 (N_9769,N_5016,N_5036);
and U9770 (N_9770,N_5949,N_7209);
and U9771 (N_9771,N_4301,N_6390);
xnor U9772 (N_9772,N_6321,N_6797);
xnor U9773 (N_9773,N_7372,N_7422);
nor U9774 (N_9774,N_6260,N_5353);
nor U9775 (N_9775,N_6417,N_6578);
nand U9776 (N_9776,N_4937,N_7566);
xnor U9777 (N_9777,N_5667,N_5609);
or U9778 (N_9778,N_6413,N_6315);
or U9779 (N_9779,N_7991,N_7861);
and U9780 (N_9780,N_6844,N_4125);
nor U9781 (N_9781,N_5215,N_7919);
nand U9782 (N_9782,N_4225,N_5355);
and U9783 (N_9783,N_4393,N_5490);
xnor U9784 (N_9784,N_5412,N_6022);
xnor U9785 (N_9785,N_7816,N_5841);
and U9786 (N_9786,N_7028,N_4636);
xor U9787 (N_9787,N_7627,N_4685);
or U9788 (N_9788,N_7294,N_7185);
or U9789 (N_9789,N_6408,N_5192);
nand U9790 (N_9790,N_6748,N_7973);
nor U9791 (N_9791,N_7499,N_7745);
and U9792 (N_9792,N_7141,N_6360);
nor U9793 (N_9793,N_4992,N_4821);
nand U9794 (N_9794,N_5435,N_7939);
or U9795 (N_9795,N_4573,N_4095);
xnor U9796 (N_9796,N_7853,N_5587);
and U9797 (N_9797,N_5248,N_7150);
nand U9798 (N_9798,N_5056,N_6191);
nand U9799 (N_9799,N_4002,N_6951);
nor U9800 (N_9800,N_7119,N_4652);
nor U9801 (N_9801,N_4630,N_6586);
xor U9802 (N_9802,N_4449,N_6108);
nand U9803 (N_9803,N_6967,N_5356);
and U9804 (N_9804,N_6571,N_7506);
nand U9805 (N_9805,N_5222,N_5066);
nand U9806 (N_9806,N_7597,N_7664);
nand U9807 (N_9807,N_5163,N_5523);
nor U9808 (N_9808,N_6158,N_7367);
xor U9809 (N_9809,N_6919,N_7685);
and U9810 (N_9810,N_4324,N_4481);
nor U9811 (N_9811,N_5266,N_7332);
nor U9812 (N_9812,N_7909,N_7684);
nor U9813 (N_9813,N_7975,N_5364);
nand U9814 (N_9814,N_5635,N_7930);
nor U9815 (N_9815,N_7046,N_4876);
xor U9816 (N_9816,N_7121,N_7245);
and U9817 (N_9817,N_6924,N_5983);
nand U9818 (N_9818,N_4028,N_7015);
nor U9819 (N_9819,N_5280,N_6379);
and U9820 (N_9820,N_7442,N_5703);
nand U9821 (N_9821,N_7828,N_7996);
xor U9822 (N_9822,N_7572,N_6708);
nor U9823 (N_9823,N_5679,N_7633);
nor U9824 (N_9824,N_7115,N_7403);
nand U9825 (N_9825,N_6731,N_5201);
nor U9826 (N_9826,N_4804,N_6506);
xnor U9827 (N_9827,N_7821,N_5113);
xor U9828 (N_9828,N_7453,N_5306);
and U9829 (N_9829,N_6659,N_5336);
nor U9830 (N_9830,N_5563,N_7812);
or U9831 (N_9831,N_6395,N_5111);
or U9832 (N_9832,N_4117,N_7091);
or U9833 (N_9833,N_4216,N_7679);
xor U9834 (N_9834,N_7786,N_6164);
xnor U9835 (N_9835,N_6149,N_5046);
and U9836 (N_9836,N_4909,N_6296);
nor U9837 (N_9837,N_5410,N_7129);
or U9838 (N_9838,N_4209,N_5713);
xnor U9839 (N_9839,N_5484,N_7464);
nand U9840 (N_9840,N_7746,N_7144);
xnor U9841 (N_9841,N_6198,N_4564);
nor U9842 (N_9842,N_4188,N_4039);
or U9843 (N_9843,N_6794,N_4024);
and U9844 (N_9844,N_7432,N_6300);
and U9845 (N_9845,N_4083,N_6025);
and U9846 (N_9846,N_7857,N_5071);
and U9847 (N_9847,N_4011,N_4386);
nand U9848 (N_9848,N_7271,N_6667);
nand U9849 (N_9849,N_7697,N_7548);
or U9850 (N_9850,N_4220,N_6385);
and U9851 (N_9851,N_7169,N_6858);
or U9852 (N_9852,N_4522,N_5837);
or U9853 (N_9853,N_7108,N_6263);
nor U9854 (N_9854,N_5107,N_6253);
xor U9855 (N_9855,N_7632,N_5008);
or U9856 (N_9856,N_7282,N_5869);
nor U9857 (N_9857,N_7214,N_5182);
nand U9858 (N_9858,N_7003,N_4340);
nor U9859 (N_9859,N_5443,N_6556);
nor U9860 (N_9860,N_7176,N_5779);
nand U9861 (N_9861,N_6489,N_7747);
nand U9862 (N_9862,N_4289,N_4840);
xor U9863 (N_9863,N_6598,N_6750);
xnor U9864 (N_9864,N_6099,N_6957);
or U9865 (N_9865,N_4755,N_4055);
nor U9866 (N_9866,N_4662,N_5607);
or U9867 (N_9867,N_5521,N_5971);
and U9868 (N_9868,N_6721,N_6574);
nand U9869 (N_9869,N_6132,N_5329);
and U9870 (N_9870,N_5404,N_4962);
or U9871 (N_9871,N_5161,N_7364);
xor U9872 (N_9872,N_5442,N_4207);
nand U9873 (N_9873,N_6053,N_5090);
and U9874 (N_9874,N_4221,N_4608);
nand U9875 (N_9875,N_6543,N_4463);
and U9876 (N_9876,N_4327,N_7577);
nand U9877 (N_9877,N_6483,N_5244);
or U9878 (N_9878,N_4634,N_5677);
and U9879 (N_9879,N_4313,N_4531);
nand U9880 (N_9880,N_4956,N_4322);
and U9881 (N_9881,N_7407,N_4739);
and U9882 (N_9882,N_6646,N_4358);
xnor U9883 (N_9883,N_7667,N_6048);
and U9884 (N_9884,N_6789,N_7977);
or U9885 (N_9885,N_7359,N_7021);
xnor U9886 (N_9886,N_5917,N_7629);
and U9887 (N_9887,N_7019,N_4830);
nand U9888 (N_9888,N_7452,N_7281);
and U9889 (N_9889,N_7106,N_7835);
and U9890 (N_9890,N_4461,N_5553);
xnor U9891 (N_9891,N_6559,N_4007);
nor U9892 (N_9892,N_7213,N_5437);
nor U9893 (N_9893,N_4191,N_5292);
or U9894 (N_9894,N_4321,N_6725);
and U9895 (N_9895,N_5770,N_5731);
and U9896 (N_9896,N_4336,N_6535);
or U9897 (N_9897,N_6993,N_6318);
nor U9898 (N_9898,N_4016,N_4654);
nand U9899 (N_9899,N_6055,N_5079);
nor U9900 (N_9900,N_5958,N_5406);
xor U9901 (N_9901,N_5397,N_4365);
or U9902 (N_9902,N_6029,N_6871);
xor U9903 (N_9903,N_7277,N_5213);
or U9904 (N_9904,N_7112,N_6208);
or U9905 (N_9905,N_4822,N_4265);
nand U9906 (N_9906,N_6854,N_7757);
and U9907 (N_9907,N_6070,N_5262);
nor U9908 (N_9908,N_4410,N_7966);
nor U9909 (N_9909,N_7165,N_7603);
and U9910 (N_9910,N_7799,N_6978);
or U9911 (N_9911,N_5072,N_6692);
and U9912 (N_9912,N_5399,N_4414);
nor U9913 (N_9913,N_7703,N_7891);
nor U9914 (N_9914,N_4090,N_6298);
xor U9915 (N_9915,N_6524,N_6081);
nand U9916 (N_9916,N_6790,N_7944);
and U9917 (N_9917,N_6823,N_7771);
xnor U9918 (N_9918,N_4502,N_6000);
xnor U9919 (N_9919,N_4594,N_6172);
nand U9920 (N_9920,N_6468,N_6156);
and U9921 (N_9921,N_7181,N_6356);
and U9922 (N_9922,N_5469,N_4702);
or U9923 (N_9923,N_5190,N_4151);
xnor U9924 (N_9924,N_4382,N_7032);
nand U9925 (N_9925,N_5172,N_4852);
nor U9926 (N_9926,N_7398,N_4545);
xor U9927 (N_9927,N_7476,N_7470);
and U9928 (N_9928,N_5926,N_4364);
or U9929 (N_9929,N_6867,N_7469);
or U9930 (N_9930,N_7310,N_7913);
nand U9931 (N_9931,N_4142,N_5543);
xnor U9932 (N_9932,N_7645,N_7371);
and U9933 (N_9933,N_7933,N_5000);
nor U9934 (N_9934,N_6458,N_5865);
nand U9935 (N_9935,N_4665,N_4896);
nand U9936 (N_9936,N_5509,N_4552);
nor U9937 (N_9937,N_6125,N_7263);
nor U9938 (N_9938,N_4239,N_6682);
nand U9939 (N_9939,N_4499,N_4902);
xnor U9940 (N_9940,N_6787,N_4747);
or U9941 (N_9941,N_7497,N_4680);
xor U9942 (N_9942,N_7565,N_4078);
nor U9943 (N_9943,N_4518,N_5350);
or U9944 (N_9944,N_5485,N_4198);
or U9945 (N_9945,N_7188,N_6231);
nor U9946 (N_9946,N_5431,N_7136);
and U9947 (N_9947,N_5009,N_7530);
and U9948 (N_9948,N_4993,N_6441);
nand U9949 (N_9949,N_7417,N_7886);
and U9950 (N_9950,N_7375,N_6813);
xor U9951 (N_9951,N_5732,N_5988);
nand U9952 (N_9952,N_4938,N_5003);
nor U9953 (N_9953,N_5675,N_7167);
or U9954 (N_9954,N_4295,N_4927);
nor U9955 (N_9955,N_4109,N_4743);
or U9956 (N_9956,N_4540,N_4418);
nand U9957 (N_9957,N_7174,N_6100);
nand U9958 (N_9958,N_4132,N_7070);
xnor U9959 (N_9959,N_4065,N_6414);
nand U9960 (N_9960,N_6195,N_5697);
or U9961 (N_9961,N_6593,N_5127);
or U9962 (N_9962,N_5234,N_5167);
or U9963 (N_9963,N_7963,N_4310);
xnor U9964 (N_9964,N_4537,N_6202);
or U9965 (N_9965,N_4917,N_4238);
or U9966 (N_9966,N_6359,N_5834);
nand U9967 (N_9967,N_6419,N_7888);
nand U9968 (N_9968,N_4253,N_5812);
and U9969 (N_9969,N_6209,N_5888);
xnor U9970 (N_9970,N_4139,N_5232);
and U9971 (N_9971,N_6018,N_5386);
and U9972 (N_9972,N_7044,N_5583);
or U9973 (N_9973,N_4193,N_7874);
nor U9974 (N_9974,N_6974,N_6808);
and U9975 (N_9975,N_4341,N_6688);
nor U9976 (N_9976,N_5735,N_7448);
xor U9977 (N_9977,N_6603,N_6513);
or U9978 (N_9978,N_6376,N_5097);
or U9979 (N_9979,N_7449,N_7014);
xor U9980 (N_9980,N_4170,N_7984);
xnor U9981 (N_9981,N_5641,N_6074);
or U9982 (N_9982,N_7087,N_5360);
and U9983 (N_9983,N_6176,N_6699);
nor U9984 (N_9984,N_5366,N_4202);
or U9985 (N_9985,N_7904,N_5529);
xnor U9986 (N_9986,N_5500,N_6609);
or U9987 (N_9987,N_4262,N_5301);
xnor U9988 (N_9988,N_4628,N_5083);
xnor U9989 (N_9989,N_6971,N_4953);
nand U9990 (N_9990,N_5470,N_4201);
xor U9991 (N_9991,N_4691,N_7316);
xor U9992 (N_9992,N_4283,N_5089);
and U9993 (N_9993,N_6564,N_4281);
nand U9994 (N_9994,N_4673,N_4914);
nand U9995 (N_9995,N_6648,N_5680);
nand U9996 (N_9996,N_6616,N_7525);
xor U9997 (N_9997,N_6450,N_6964);
nand U9998 (N_9998,N_4160,N_5694);
and U9999 (N_9999,N_6442,N_6716);
nor U10000 (N_10000,N_5952,N_6467);
nand U10001 (N_10001,N_6931,N_4520);
nor U10002 (N_10002,N_5639,N_6965);
xor U10003 (N_10003,N_7462,N_4551);
and U10004 (N_10004,N_6088,N_6675);
nor U10005 (N_10005,N_4146,N_4978);
nor U10006 (N_10006,N_5778,N_6655);
and U10007 (N_10007,N_7796,N_7582);
xor U10008 (N_10008,N_4647,N_5472);
nor U10009 (N_10009,N_7252,N_7296);
nand U10010 (N_10010,N_6199,N_4637);
xnor U10011 (N_10011,N_6143,N_7296);
nand U10012 (N_10012,N_4504,N_4042);
nor U10013 (N_10013,N_6240,N_4409);
nor U10014 (N_10014,N_7387,N_5359);
xor U10015 (N_10015,N_7771,N_6258);
xnor U10016 (N_10016,N_6821,N_5742);
xnor U10017 (N_10017,N_4685,N_4623);
and U10018 (N_10018,N_7906,N_6783);
nand U10019 (N_10019,N_6744,N_6907);
xor U10020 (N_10020,N_6903,N_7231);
nor U10021 (N_10021,N_5046,N_7138);
or U10022 (N_10022,N_4502,N_6740);
nor U10023 (N_10023,N_7910,N_6632);
or U10024 (N_10024,N_4442,N_6192);
xor U10025 (N_10025,N_6885,N_7038);
or U10026 (N_10026,N_6995,N_5765);
and U10027 (N_10027,N_7499,N_5645);
and U10028 (N_10028,N_6688,N_4134);
or U10029 (N_10029,N_7309,N_6803);
nor U10030 (N_10030,N_7964,N_5572);
nand U10031 (N_10031,N_4858,N_7329);
or U10032 (N_10032,N_7570,N_4132);
or U10033 (N_10033,N_4782,N_7202);
nor U10034 (N_10034,N_4256,N_4434);
or U10035 (N_10035,N_4690,N_4938);
and U10036 (N_10036,N_4671,N_5515);
nand U10037 (N_10037,N_4559,N_4377);
nand U10038 (N_10038,N_6333,N_7708);
nand U10039 (N_10039,N_4823,N_6420);
nand U10040 (N_10040,N_6568,N_6612);
xor U10041 (N_10041,N_7171,N_5998);
or U10042 (N_10042,N_6981,N_5052);
nand U10043 (N_10043,N_5067,N_5394);
and U10044 (N_10044,N_5168,N_7635);
or U10045 (N_10045,N_6047,N_6699);
or U10046 (N_10046,N_5566,N_5539);
and U10047 (N_10047,N_7049,N_4665);
xnor U10048 (N_10048,N_4877,N_7828);
and U10049 (N_10049,N_6394,N_4625);
nand U10050 (N_10050,N_4156,N_7913);
nand U10051 (N_10051,N_5899,N_7020);
or U10052 (N_10052,N_4987,N_7397);
xor U10053 (N_10053,N_4325,N_5618);
nand U10054 (N_10054,N_4562,N_4319);
nor U10055 (N_10055,N_4652,N_6729);
nor U10056 (N_10056,N_5198,N_4683);
xor U10057 (N_10057,N_7460,N_4158);
and U10058 (N_10058,N_6256,N_7061);
or U10059 (N_10059,N_4535,N_6673);
xnor U10060 (N_10060,N_4248,N_6302);
xnor U10061 (N_10061,N_5408,N_6580);
nor U10062 (N_10062,N_6667,N_5944);
nand U10063 (N_10063,N_4397,N_4941);
and U10064 (N_10064,N_4423,N_5327);
nor U10065 (N_10065,N_5738,N_5075);
nand U10066 (N_10066,N_7779,N_7257);
and U10067 (N_10067,N_4944,N_7870);
or U10068 (N_10068,N_6302,N_5021);
or U10069 (N_10069,N_5667,N_7843);
and U10070 (N_10070,N_5680,N_5926);
or U10071 (N_10071,N_7058,N_7218);
nor U10072 (N_10072,N_6678,N_6411);
nor U10073 (N_10073,N_5782,N_5781);
nor U10074 (N_10074,N_4846,N_6106);
xnor U10075 (N_10075,N_6917,N_6753);
nor U10076 (N_10076,N_5934,N_6629);
nor U10077 (N_10077,N_5461,N_7550);
nand U10078 (N_10078,N_5488,N_5400);
and U10079 (N_10079,N_5158,N_4512);
nor U10080 (N_10080,N_5049,N_7272);
xnor U10081 (N_10081,N_6771,N_7911);
or U10082 (N_10082,N_5847,N_4325);
nand U10083 (N_10083,N_4732,N_6844);
or U10084 (N_10084,N_4764,N_6602);
and U10085 (N_10085,N_7015,N_5035);
xnor U10086 (N_10086,N_5017,N_4496);
or U10087 (N_10087,N_7981,N_7532);
and U10088 (N_10088,N_5319,N_5231);
and U10089 (N_10089,N_4219,N_4857);
or U10090 (N_10090,N_4401,N_7483);
or U10091 (N_10091,N_5217,N_5279);
and U10092 (N_10092,N_6778,N_7706);
nand U10093 (N_10093,N_6878,N_6577);
xor U10094 (N_10094,N_7400,N_6096);
nor U10095 (N_10095,N_7649,N_4045);
nor U10096 (N_10096,N_7203,N_6447);
and U10097 (N_10097,N_7651,N_5726);
nand U10098 (N_10098,N_5333,N_7327);
xor U10099 (N_10099,N_4740,N_7999);
nor U10100 (N_10100,N_5071,N_6342);
nor U10101 (N_10101,N_7391,N_7599);
or U10102 (N_10102,N_4130,N_6020);
xnor U10103 (N_10103,N_4253,N_6017);
nand U10104 (N_10104,N_5054,N_5484);
nand U10105 (N_10105,N_4834,N_4227);
or U10106 (N_10106,N_6274,N_5510);
xor U10107 (N_10107,N_6322,N_7733);
xor U10108 (N_10108,N_5950,N_7780);
and U10109 (N_10109,N_4996,N_5145);
nand U10110 (N_10110,N_7332,N_7055);
xor U10111 (N_10111,N_6490,N_6547);
and U10112 (N_10112,N_7346,N_4750);
nor U10113 (N_10113,N_7461,N_4197);
and U10114 (N_10114,N_4877,N_7118);
nand U10115 (N_10115,N_5841,N_6978);
xnor U10116 (N_10116,N_4212,N_5827);
nand U10117 (N_10117,N_4481,N_5712);
xnor U10118 (N_10118,N_6811,N_4835);
nor U10119 (N_10119,N_4254,N_6601);
xnor U10120 (N_10120,N_7735,N_7292);
nand U10121 (N_10121,N_4443,N_4310);
nor U10122 (N_10122,N_5041,N_7463);
nor U10123 (N_10123,N_7436,N_7837);
xnor U10124 (N_10124,N_4699,N_4342);
and U10125 (N_10125,N_4514,N_7400);
or U10126 (N_10126,N_7696,N_4862);
or U10127 (N_10127,N_4569,N_7200);
nor U10128 (N_10128,N_7370,N_7700);
or U10129 (N_10129,N_6454,N_7891);
and U10130 (N_10130,N_4913,N_5589);
or U10131 (N_10131,N_6804,N_5327);
nand U10132 (N_10132,N_6878,N_7789);
nor U10133 (N_10133,N_6542,N_6221);
or U10134 (N_10134,N_5449,N_5190);
nor U10135 (N_10135,N_7865,N_5114);
xor U10136 (N_10136,N_6998,N_4644);
nor U10137 (N_10137,N_7175,N_4189);
and U10138 (N_10138,N_4754,N_4781);
nand U10139 (N_10139,N_7476,N_4437);
xnor U10140 (N_10140,N_5504,N_7076);
xor U10141 (N_10141,N_6267,N_6835);
nand U10142 (N_10142,N_6167,N_5151);
nand U10143 (N_10143,N_6460,N_6335);
nand U10144 (N_10144,N_4409,N_7105);
xnor U10145 (N_10145,N_7549,N_5576);
nor U10146 (N_10146,N_6865,N_5570);
or U10147 (N_10147,N_6887,N_5645);
nand U10148 (N_10148,N_7569,N_6867);
xor U10149 (N_10149,N_5121,N_6779);
nor U10150 (N_10150,N_7370,N_7042);
or U10151 (N_10151,N_5162,N_7359);
nor U10152 (N_10152,N_5651,N_4137);
nand U10153 (N_10153,N_7297,N_4972);
and U10154 (N_10154,N_6777,N_6263);
nand U10155 (N_10155,N_4225,N_6183);
or U10156 (N_10156,N_4578,N_6410);
nand U10157 (N_10157,N_6538,N_5931);
xnor U10158 (N_10158,N_5666,N_4642);
or U10159 (N_10159,N_4471,N_5342);
nor U10160 (N_10160,N_6265,N_5209);
nand U10161 (N_10161,N_4087,N_7834);
and U10162 (N_10162,N_6955,N_4525);
and U10163 (N_10163,N_6435,N_4659);
nand U10164 (N_10164,N_6557,N_6621);
or U10165 (N_10165,N_5752,N_6064);
xor U10166 (N_10166,N_6755,N_5079);
or U10167 (N_10167,N_6228,N_6898);
nor U10168 (N_10168,N_6542,N_4458);
xor U10169 (N_10169,N_4046,N_5279);
and U10170 (N_10170,N_6578,N_6231);
xnor U10171 (N_10171,N_4731,N_4985);
xnor U10172 (N_10172,N_4361,N_7291);
xnor U10173 (N_10173,N_5297,N_6951);
or U10174 (N_10174,N_6801,N_4337);
nand U10175 (N_10175,N_6215,N_7439);
or U10176 (N_10176,N_4911,N_5320);
nand U10177 (N_10177,N_4422,N_7854);
or U10178 (N_10178,N_6640,N_6368);
nand U10179 (N_10179,N_6983,N_5361);
and U10180 (N_10180,N_7529,N_7784);
or U10181 (N_10181,N_6345,N_4717);
and U10182 (N_10182,N_4987,N_6572);
xnor U10183 (N_10183,N_6918,N_4640);
nand U10184 (N_10184,N_4462,N_7669);
and U10185 (N_10185,N_4744,N_5148);
or U10186 (N_10186,N_6267,N_4220);
and U10187 (N_10187,N_4942,N_7046);
and U10188 (N_10188,N_4878,N_7822);
or U10189 (N_10189,N_7643,N_6679);
nand U10190 (N_10190,N_5267,N_4987);
nor U10191 (N_10191,N_5255,N_6518);
nand U10192 (N_10192,N_5425,N_7934);
or U10193 (N_10193,N_6414,N_4226);
nor U10194 (N_10194,N_7473,N_4336);
nand U10195 (N_10195,N_7585,N_5899);
nand U10196 (N_10196,N_7267,N_6236);
xor U10197 (N_10197,N_5576,N_7861);
nor U10198 (N_10198,N_7506,N_7846);
and U10199 (N_10199,N_7701,N_5947);
xnor U10200 (N_10200,N_4532,N_6763);
nand U10201 (N_10201,N_7204,N_4096);
and U10202 (N_10202,N_7819,N_6021);
and U10203 (N_10203,N_6796,N_4352);
nor U10204 (N_10204,N_4956,N_7122);
nor U10205 (N_10205,N_5424,N_7679);
and U10206 (N_10206,N_4119,N_6547);
xnor U10207 (N_10207,N_7210,N_5755);
xor U10208 (N_10208,N_7829,N_4687);
or U10209 (N_10209,N_5754,N_7992);
xor U10210 (N_10210,N_7015,N_4178);
xnor U10211 (N_10211,N_4067,N_7127);
nor U10212 (N_10212,N_7870,N_5566);
nand U10213 (N_10213,N_7074,N_6998);
nand U10214 (N_10214,N_6786,N_5552);
nand U10215 (N_10215,N_7865,N_4675);
or U10216 (N_10216,N_7470,N_6507);
nor U10217 (N_10217,N_7998,N_7654);
nor U10218 (N_10218,N_4982,N_4352);
or U10219 (N_10219,N_7863,N_4724);
and U10220 (N_10220,N_4872,N_7584);
nor U10221 (N_10221,N_6375,N_6873);
xor U10222 (N_10222,N_6015,N_5685);
nand U10223 (N_10223,N_4463,N_5307);
nand U10224 (N_10224,N_5853,N_6456);
nor U10225 (N_10225,N_4701,N_4718);
nor U10226 (N_10226,N_6268,N_4576);
nor U10227 (N_10227,N_5740,N_5837);
and U10228 (N_10228,N_7207,N_6025);
xnor U10229 (N_10229,N_6669,N_4033);
nand U10230 (N_10230,N_6811,N_6741);
and U10231 (N_10231,N_7697,N_6735);
and U10232 (N_10232,N_5966,N_5887);
and U10233 (N_10233,N_4091,N_4021);
nand U10234 (N_10234,N_6462,N_6952);
or U10235 (N_10235,N_6950,N_7908);
and U10236 (N_10236,N_6958,N_7631);
nor U10237 (N_10237,N_4951,N_5627);
nand U10238 (N_10238,N_7729,N_7932);
or U10239 (N_10239,N_5672,N_4317);
and U10240 (N_10240,N_6693,N_5735);
nand U10241 (N_10241,N_7198,N_7608);
nor U10242 (N_10242,N_5151,N_7744);
and U10243 (N_10243,N_6847,N_6228);
nor U10244 (N_10244,N_6348,N_5948);
and U10245 (N_10245,N_4997,N_6082);
nand U10246 (N_10246,N_5079,N_7384);
and U10247 (N_10247,N_4262,N_4507);
nand U10248 (N_10248,N_7605,N_5523);
nor U10249 (N_10249,N_5970,N_4034);
xor U10250 (N_10250,N_5346,N_5855);
or U10251 (N_10251,N_6914,N_6124);
and U10252 (N_10252,N_6116,N_4897);
xnor U10253 (N_10253,N_4589,N_4512);
and U10254 (N_10254,N_6229,N_4394);
nand U10255 (N_10255,N_5746,N_4619);
nor U10256 (N_10256,N_7018,N_7496);
xor U10257 (N_10257,N_7887,N_4012);
nand U10258 (N_10258,N_6297,N_5147);
or U10259 (N_10259,N_5277,N_6341);
xnor U10260 (N_10260,N_5430,N_7770);
nor U10261 (N_10261,N_6773,N_5219);
nor U10262 (N_10262,N_4463,N_4809);
nor U10263 (N_10263,N_5554,N_4902);
nor U10264 (N_10264,N_4843,N_5176);
nor U10265 (N_10265,N_6172,N_7118);
or U10266 (N_10266,N_4984,N_6758);
xnor U10267 (N_10267,N_4256,N_6328);
and U10268 (N_10268,N_4239,N_6128);
nand U10269 (N_10269,N_4257,N_6128);
nor U10270 (N_10270,N_6545,N_6757);
or U10271 (N_10271,N_4017,N_7706);
xnor U10272 (N_10272,N_6008,N_5969);
nor U10273 (N_10273,N_4573,N_4412);
xor U10274 (N_10274,N_6673,N_4853);
nor U10275 (N_10275,N_4346,N_4002);
nand U10276 (N_10276,N_5659,N_5558);
nor U10277 (N_10277,N_7778,N_6167);
nand U10278 (N_10278,N_4786,N_6018);
or U10279 (N_10279,N_6430,N_7663);
and U10280 (N_10280,N_5368,N_5631);
nor U10281 (N_10281,N_5187,N_6753);
nand U10282 (N_10282,N_7053,N_5755);
nor U10283 (N_10283,N_5250,N_6431);
nor U10284 (N_10284,N_6824,N_7335);
nand U10285 (N_10285,N_4277,N_4313);
nand U10286 (N_10286,N_5351,N_4122);
and U10287 (N_10287,N_7996,N_6050);
nor U10288 (N_10288,N_6315,N_5716);
nand U10289 (N_10289,N_7381,N_6253);
nand U10290 (N_10290,N_4394,N_4452);
nand U10291 (N_10291,N_5310,N_4081);
nor U10292 (N_10292,N_4921,N_7344);
xnor U10293 (N_10293,N_4416,N_5281);
and U10294 (N_10294,N_4646,N_4628);
xnor U10295 (N_10295,N_4270,N_4762);
and U10296 (N_10296,N_5346,N_4169);
or U10297 (N_10297,N_7488,N_6823);
nand U10298 (N_10298,N_4629,N_5871);
or U10299 (N_10299,N_5422,N_6588);
nand U10300 (N_10300,N_5103,N_5659);
xor U10301 (N_10301,N_6953,N_6932);
nand U10302 (N_10302,N_4919,N_5228);
nor U10303 (N_10303,N_4640,N_6737);
or U10304 (N_10304,N_6946,N_6219);
and U10305 (N_10305,N_4666,N_4458);
nor U10306 (N_10306,N_4561,N_7483);
and U10307 (N_10307,N_6383,N_6694);
nor U10308 (N_10308,N_4537,N_7788);
nand U10309 (N_10309,N_5339,N_7043);
xor U10310 (N_10310,N_7434,N_4200);
xor U10311 (N_10311,N_5465,N_6089);
nand U10312 (N_10312,N_4015,N_7092);
nand U10313 (N_10313,N_4967,N_7545);
nand U10314 (N_10314,N_6724,N_6913);
nand U10315 (N_10315,N_4213,N_5599);
nor U10316 (N_10316,N_7855,N_7200);
and U10317 (N_10317,N_7339,N_6301);
nor U10318 (N_10318,N_6491,N_7196);
xor U10319 (N_10319,N_5386,N_5777);
nor U10320 (N_10320,N_5110,N_5091);
nor U10321 (N_10321,N_7141,N_4848);
nor U10322 (N_10322,N_6694,N_5177);
and U10323 (N_10323,N_7082,N_6669);
or U10324 (N_10324,N_4783,N_6108);
xnor U10325 (N_10325,N_6207,N_7831);
or U10326 (N_10326,N_7366,N_6096);
or U10327 (N_10327,N_6734,N_4619);
nand U10328 (N_10328,N_7892,N_7877);
or U10329 (N_10329,N_7022,N_7227);
nor U10330 (N_10330,N_6958,N_7675);
nor U10331 (N_10331,N_6293,N_7067);
and U10332 (N_10332,N_7504,N_7730);
nor U10333 (N_10333,N_5654,N_6438);
xor U10334 (N_10334,N_7771,N_6358);
nand U10335 (N_10335,N_5918,N_6428);
nor U10336 (N_10336,N_4870,N_6867);
and U10337 (N_10337,N_6853,N_6426);
xnor U10338 (N_10338,N_6308,N_5806);
xnor U10339 (N_10339,N_7027,N_5020);
nand U10340 (N_10340,N_5250,N_6619);
or U10341 (N_10341,N_4917,N_6988);
or U10342 (N_10342,N_7878,N_6979);
xor U10343 (N_10343,N_4035,N_4767);
xor U10344 (N_10344,N_5907,N_5634);
nand U10345 (N_10345,N_7175,N_6021);
and U10346 (N_10346,N_6888,N_4880);
nor U10347 (N_10347,N_5077,N_7696);
nor U10348 (N_10348,N_6282,N_6133);
xnor U10349 (N_10349,N_7805,N_4832);
xor U10350 (N_10350,N_5815,N_6533);
nand U10351 (N_10351,N_6181,N_6280);
xnor U10352 (N_10352,N_7428,N_5332);
nand U10353 (N_10353,N_5865,N_5825);
xor U10354 (N_10354,N_5628,N_6326);
and U10355 (N_10355,N_7612,N_4700);
xnor U10356 (N_10356,N_5401,N_5602);
nand U10357 (N_10357,N_6719,N_6707);
xor U10358 (N_10358,N_5575,N_6923);
or U10359 (N_10359,N_4030,N_7446);
nor U10360 (N_10360,N_6860,N_4096);
nand U10361 (N_10361,N_6586,N_7119);
nand U10362 (N_10362,N_7499,N_7510);
xor U10363 (N_10363,N_6479,N_7326);
and U10364 (N_10364,N_7539,N_4066);
or U10365 (N_10365,N_4994,N_6014);
xnor U10366 (N_10366,N_6133,N_7076);
nor U10367 (N_10367,N_6462,N_5318);
nor U10368 (N_10368,N_7104,N_6174);
nor U10369 (N_10369,N_7923,N_6720);
xnor U10370 (N_10370,N_6102,N_7340);
nand U10371 (N_10371,N_5565,N_6813);
or U10372 (N_10372,N_5712,N_6547);
or U10373 (N_10373,N_7027,N_4102);
or U10374 (N_10374,N_5164,N_7401);
nand U10375 (N_10375,N_7432,N_7901);
xor U10376 (N_10376,N_4481,N_5884);
or U10377 (N_10377,N_6850,N_5941);
nand U10378 (N_10378,N_6018,N_6392);
nand U10379 (N_10379,N_6252,N_5338);
nand U10380 (N_10380,N_6818,N_6924);
and U10381 (N_10381,N_4843,N_5354);
nor U10382 (N_10382,N_6106,N_6009);
and U10383 (N_10383,N_6495,N_4315);
xnor U10384 (N_10384,N_4223,N_4275);
or U10385 (N_10385,N_4536,N_4753);
and U10386 (N_10386,N_4699,N_6476);
nor U10387 (N_10387,N_5799,N_4152);
and U10388 (N_10388,N_7439,N_7920);
and U10389 (N_10389,N_4244,N_4988);
and U10390 (N_10390,N_5459,N_4757);
nand U10391 (N_10391,N_4733,N_6185);
or U10392 (N_10392,N_4891,N_5308);
nor U10393 (N_10393,N_7019,N_4991);
xor U10394 (N_10394,N_7199,N_4451);
or U10395 (N_10395,N_6680,N_6866);
xor U10396 (N_10396,N_6198,N_6647);
and U10397 (N_10397,N_5056,N_7094);
nand U10398 (N_10398,N_4786,N_4981);
and U10399 (N_10399,N_5628,N_5229);
xnor U10400 (N_10400,N_5393,N_7843);
or U10401 (N_10401,N_4900,N_5433);
or U10402 (N_10402,N_6143,N_6162);
or U10403 (N_10403,N_5401,N_5037);
nand U10404 (N_10404,N_6156,N_6182);
or U10405 (N_10405,N_7332,N_6869);
nor U10406 (N_10406,N_7786,N_7950);
nor U10407 (N_10407,N_4376,N_7206);
nor U10408 (N_10408,N_6950,N_7154);
xor U10409 (N_10409,N_4718,N_7542);
nor U10410 (N_10410,N_7252,N_4414);
and U10411 (N_10411,N_4909,N_7283);
xor U10412 (N_10412,N_5617,N_7106);
xor U10413 (N_10413,N_5676,N_5439);
and U10414 (N_10414,N_7636,N_5717);
and U10415 (N_10415,N_5868,N_5247);
and U10416 (N_10416,N_6041,N_6033);
nand U10417 (N_10417,N_6156,N_4093);
nor U10418 (N_10418,N_6034,N_5122);
xor U10419 (N_10419,N_7835,N_7261);
nand U10420 (N_10420,N_5161,N_4361);
or U10421 (N_10421,N_4224,N_6285);
and U10422 (N_10422,N_4406,N_6780);
and U10423 (N_10423,N_5387,N_7884);
xnor U10424 (N_10424,N_7577,N_6231);
nor U10425 (N_10425,N_6048,N_4944);
xor U10426 (N_10426,N_6210,N_5618);
nand U10427 (N_10427,N_6355,N_5701);
nand U10428 (N_10428,N_7910,N_5637);
or U10429 (N_10429,N_5388,N_5179);
xnor U10430 (N_10430,N_6781,N_7280);
nand U10431 (N_10431,N_6787,N_7412);
or U10432 (N_10432,N_5125,N_4197);
nand U10433 (N_10433,N_6509,N_4760);
xnor U10434 (N_10434,N_6443,N_7449);
nand U10435 (N_10435,N_4797,N_6831);
nand U10436 (N_10436,N_4126,N_5078);
nand U10437 (N_10437,N_5575,N_5916);
xor U10438 (N_10438,N_7669,N_5055);
xor U10439 (N_10439,N_4196,N_7161);
or U10440 (N_10440,N_4568,N_5398);
or U10441 (N_10441,N_7705,N_5081);
xnor U10442 (N_10442,N_7632,N_6858);
and U10443 (N_10443,N_7430,N_5825);
or U10444 (N_10444,N_7949,N_5697);
xnor U10445 (N_10445,N_6438,N_5743);
or U10446 (N_10446,N_5431,N_4354);
nand U10447 (N_10447,N_6415,N_6706);
nand U10448 (N_10448,N_4374,N_5075);
nand U10449 (N_10449,N_7351,N_5163);
and U10450 (N_10450,N_5420,N_5506);
nand U10451 (N_10451,N_7597,N_5700);
nand U10452 (N_10452,N_5429,N_5962);
and U10453 (N_10453,N_7883,N_4576);
nor U10454 (N_10454,N_6989,N_5410);
xnor U10455 (N_10455,N_5945,N_6273);
nand U10456 (N_10456,N_7738,N_5018);
nor U10457 (N_10457,N_7819,N_4975);
nand U10458 (N_10458,N_4114,N_7372);
and U10459 (N_10459,N_7739,N_5194);
nor U10460 (N_10460,N_7176,N_7419);
xor U10461 (N_10461,N_7783,N_6131);
xnor U10462 (N_10462,N_7335,N_5964);
xor U10463 (N_10463,N_7213,N_7974);
or U10464 (N_10464,N_7837,N_5398);
nor U10465 (N_10465,N_4657,N_6324);
nor U10466 (N_10466,N_5467,N_5185);
nor U10467 (N_10467,N_7213,N_4319);
xnor U10468 (N_10468,N_7373,N_7985);
and U10469 (N_10469,N_5933,N_4683);
xor U10470 (N_10470,N_6364,N_4393);
xor U10471 (N_10471,N_5420,N_4174);
and U10472 (N_10472,N_4047,N_4914);
xor U10473 (N_10473,N_4677,N_4335);
or U10474 (N_10474,N_7390,N_5303);
xnor U10475 (N_10475,N_5606,N_6234);
xor U10476 (N_10476,N_5716,N_4046);
and U10477 (N_10477,N_4671,N_4274);
xnor U10478 (N_10478,N_7766,N_5537);
xor U10479 (N_10479,N_7152,N_4318);
nor U10480 (N_10480,N_7855,N_6731);
or U10481 (N_10481,N_7510,N_6053);
nor U10482 (N_10482,N_7532,N_6544);
xnor U10483 (N_10483,N_5733,N_5363);
nor U10484 (N_10484,N_6364,N_5757);
and U10485 (N_10485,N_5430,N_5969);
or U10486 (N_10486,N_7165,N_5714);
nand U10487 (N_10487,N_7512,N_6297);
nand U10488 (N_10488,N_4570,N_7972);
or U10489 (N_10489,N_4526,N_4780);
nor U10490 (N_10490,N_5788,N_4264);
nand U10491 (N_10491,N_5123,N_7867);
nand U10492 (N_10492,N_5056,N_4070);
or U10493 (N_10493,N_4056,N_5272);
nor U10494 (N_10494,N_7287,N_6009);
xor U10495 (N_10495,N_7198,N_4344);
or U10496 (N_10496,N_6886,N_5967);
nor U10497 (N_10497,N_5864,N_5721);
nand U10498 (N_10498,N_5658,N_6466);
nand U10499 (N_10499,N_5842,N_6333);
nor U10500 (N_10500,N_5814,N_5377);
or U10501 (N_10501,N_5287,N_5331);
nand U10502 (N_10502,N_4859,N_4325);
xor U10503 (N_10503,N_7256,N_4755);
xor U10504 (N_10504,N_7714,N_6046);
or U10505 (N_10505,N_6751,N_4472);
xnor U10506 (N_10506,N_6853,N_6135);
xor U10507 (N_10507,N_4781,N_4187);
nor U10508 (N_10508,N_4731,N_7723);
nor U10509 (N_10509,N_4102,N_4545);
xor U10510 (N_10510,N_7912,N_6427);
xor U10511 (N_10511,N_4772,N_5015);
nor U10512 (N_10512,N_6976,N_7936);
xnor U10513 (N_10513,N_7427,N_7334);
and U10514 (N_10514,N_7370,N_5197);
and U10515 (N_10515,N_6867,N_5309);
or U10516 (N_10516,N_5753,N_6798);
nand U10517 (N_10517,N_6965,N_7410);
nor U10518 (N_10518,N_4355,N_5737);
nand U10519 (N_10519,N_6356,N_4959);
or U10520 (N_10520,N_5957,N_4440);
xor U10521 (N_10521,N_4866,N_7033);
xnor U10522 (N_10522,N_7478,N_5560);
nand U10523 (N_10523,N_6774,N_7885);
nand U10524 (N_10524,N_6523,N_5931);
and U10525 (N_10525,N_5699,N_7575);
nand U10526 (N_10526,N_6113,N_6982);
and U10527 (N_10527,N_6334,N_4531);
and U10528 (N_10528,N_5456,N_7529);
xnor U10529 (N_10529,N_5975,N_6948);
nand U10530 (N_10530,N_4028,N_7884);
nor U10531 (N_10531,N_5845,N_7252);
and U10532 (N_10532,N_6134,N_6790);
and U10533 (N_10533,N_4971,N_5480);
xnor U10534 (N_10534,N_7799,N_5355);
nand U10535 (N_10535,N_6196,N_5252);
and U10536 (N_10536,N_5744,N_6356);
nand U10537 (N_10537,N_5345,N_7343);
and U10538 (N_10538,N_4522,N_5593);
xnor U10539 (N_10539,N_4716,N_5489);
nor U10540 (N_10540,N_6846,N_5521);
nand U10541 (N_10541,N_7027,N_5580);
and U10542 (N_10542,N_5356,N_4530);
nand U10543 (N_10543,N_7763,N_6742);
xor U10544 (N_10544,N_6830,N_5013);
nor U10545 (N_10545,N_6511,N_4143);
nand U10546 (N_10546,N_4939,N_6349);
nand U10547 (N_10547,N_6017,N_4091);
or U10548 (N_10548,N_6239,N_5324);
or U10549 (N_10549,N_7376,N_4930);
or U10550 (N_10550,N_5994,N_5601);
or U10551 (N_10551,N_7242,N_6083);
xor U10552 (N_10552,N_6723,N_4529);
xor U10553 (N_10553,N_7187,N_6597);
xor U10554 (N_10554,N_4772,N_4427);
nor U10555 (N_10555,N_7375,N_6964);
nor U10556 (N_10556,N_5197,N_5202);
and U10557 (N_10557,N_7589,N_5387);
nor U10558 (N_10558,N_6904,N_6103);
nor U10559 (N_10559,N_4426,N_5172);
and U10560 (N_10560,N_6231,N_4377);
and U10561 (N_10561,N_5147,N_6117);
xnor U10562 (N_10562,N_6443,N_6902);
or U10563 (N_10563,N_4951,N_6231);
nor U10564 (N_10564,N_7524,N_5801);
or U10565 (N_10565,N_4756,N_7843);
or U10566 (N_10566,N_7045,N_7154);
and U10567 (N_10567,N_4364,N_7952);
nand U10568 (N_10568,N_7006,N_4253);
or U10569 (N_10569,N_7767,N_5903);
nand U10570 (N_10570,N_7390,N_4841);
xnor U10571 (N_10571,N_7263,N_4044);
xnor U10572 (N_10572,N_5230,N_7934);
and U10573 (N_10573,N_7844,N_4154);
or U10574 (N_10574,N_7637,N_5526);
nor U10575 (N_10575,N_7315,N_5167);
and U10576 (N_10576,N_6677,N_4332);
or U10577 (N_10577,N_5850,N_7269);
xnor U10578 (N_10578,N_4371,N_5002);
and U10579 (N_10579,N_7285,N_7972);
xnor U10580 (N_10580,N_6878,N_4164);
or U10581 (N_10581,N_5759,N_4843);
xnor U10582 (N_10582,N_4749,N_4984);
or U10583 (N_10583,N_7482,N_5001);
nor U10584 (N_10584,N_4358,N_5860);
xnor U10585 (N_10585,N_6705,N_4486);
nand U10586 (N_10586,N_4863,N_6418);
or U10587 (N_10587,N_7133,N_6843);
nor U10588 (N_10588,N_5595,N_5489);
nand U10589 (N_10589,N_5616,N_4912);
and U10590 (N_10590,N_7566,N_6045);
xnor U10591 (N_10591,N_5880,N_7285);
xor U10592 (N_10592,N_7923,N_7851);
nand U10593 (N_10593,N_4975,N_4340);
nor U10594 (N_10594,N_7056,N_6675);
xor U10595 (N_10595,N_5368,N_7957);
nand U10596 (N_10596,N_4201,N_4615);
and U10597 (N_10597,N_4474,N_4609);
nor U10598 (N_10598,N_5423,N_5896);
xor U10599 (N_10599,N_6410,N_6580);
xnor U10600 (N_10600,N_4940,N_4618);
nor U10601 (N_10601,N_5752,N_7470);
nand U10602 (N_10602,N_4634,N_6768);
xor U10603 (N_10603,N_4830,N_6319);
xor U10604 (N_10604,N_6712,N_4696);
xor U10605 (N_10605,N_6533,N_6931);
nand U10606 (N_10606,N_4050,N_7690);
and U10607 (N_10607,N_7634,N_7263);
nand U10608 (N_10608,N_7432,N_5592);
nand U10609 (N_10609,N_5264,N_6400);
nand U10610 (N_10610,N_7185,N_6257);
or U10611 (N_10611,N_6913,N_4648);
xnor U10612 (N_10612,N_7325,N_4933);
or U10613 (N_10613,N_7367,N_7276);
or U10614 (N_10614,N_4555,N_7211);
nand U10615 (N_10615,N_7750,N_5979);
xnor U10616 (N_10616,N_4028,N_5415);
xnor U10617 (N_10617,N_4540,N_4742);
nor U10618 (N_10618,N_6484,N_4362);
and U10619 (N_10619,N_4001,N_5984);
and U10620 (N_10620,N_5747,N_5116);
nand U10621 (N_10621,N_5566,N_6634);
xnor U10622 (N_10622,N_5394,N_7111);
nand U10623 (N_10623,N_5078,N_4370);
and U10624 (N_10624,N_6839,N_5066);
nor U10625 (N_10625,N_7992,N_5649);
and U10626 (N_10626,N_6505,N_5551);
or U10627 (N_10627,N_6055,N_5950);
or U10628 (N_10628,N_4018,N_4934);
nor U10629 (N_10629,N_4338,N_7466);
xnor U10630 (N_10630,N_4492,N_7156);
and U10631 (N_10631,N_6778,N_4152);
xor U10632 (N_10632,N_6940,N_7473);
nor U10633 (N_10633,N_5198,N_7165);
nand U10634 (N_10634,N_5176,N_7647);
nor U10635 (N_10635,N_6748,N_6620);
and U10636 (N_10636,N_5280,N_4982);
xor U10637 (N_10637,N_7386,N_5100);
and U10638 (N_10638,N_5563,N_7622);
or U10639 (N_10639,N_5874,N_7751);
nor U10640 (N_10640,N_6612,N_4861);
and U10641 (N_10641,N_7242,N_4901);
and U10642 (N_10642,N_5197,N_4872);
nand U10643 (N_10643,N_6777,N_7118);
and U10644 (N_10644,N_4554,N_6159);
nand U10645 (N_10645,N_4227,N_5992);
nand U10646 (N_10646,N_4927,N_7973);
nand U10647 (N_10647,N_5565,N_5408);
and U10648 (N_10648,N_6731,N_6234);
xnor U10649 (N_10649,N_6245,N_7895);
or U10650 (N_10650,N_5243,N_4498);
nand U10651 (N_10651,N_5044,N_7667);
nor U10652 (N_10652,N_7885,N_5815);
and U10653 (N_10653,N_4666,N_7078);
nor U10654 (N_10654,N_6872,N_6141);
nor U10655 (N_10655,N_4981,N_4742);
or U10656 (N_10656,N_7074,N_4796);
xor U10657 (N_10657,N_7608,N_6875);
and U10658 (N_10658,N_5994,N_7024);
nand U10659 (N_10659,N_4181,N_5791);
nor U10660 (N_10660,N_5602,N_7960);
and U10661 (N_10661,N_5196,N_6713);
and U10662 (N_10662,N_6147,N_7160);
and U10663 (N_10663,N_4574,N_5670);
or U10664 (N_10664,N_7536,N_4425);
and U10665 (N_10665,N_5925,N_5547);
nor U10666 (N_10666,N_5755,N_6604);
xor U10667 (N_10667,N_4545,N_7252);
nor U10668 (N_10668,N_4717,N_7809);
or U10669 (N_10669,N_5705,N_5355);
or U10670 (N_10670,N_5573,N_5575);
xnor U10671 (N_10671,N_5664,N_4511);
xnor U10672 (N_10672,N_5055,N_6659);
nor U10673 (N_10673,N_7505,N_4914);
nand U10674 (N_10674,N_6336,N_7995);
xor U10675 (N_10675,N_7931,N_5908);
xnor U10676 (N_10676,N_7591,N_7105);
and U10677 (N_10677,N_6400,N_6183);
nand U10678 (N_10678,N_4504,N_5186);
nor U10679 (N_10679,N_7275,N_7534);
nor U10680 (N_10680,N_4802,N_6669);
nand U10681 (N_10681,N_6947,N_7206);
nor U10682 (N_10682,N_5614,N_7090);
nor U10683 (N_10683,N_4869,N_7888);
or U10684 (N_10684,N_4848,N_7451);
and U10685 (N_10685,N_5877,N_5687);
and U10686 (N_10686,N_5208,N_6117);
or U10687 (N_10687,N_7155,N_6251);
xor U10688 (N_10688,N_4968,N_4977);
nor U10689 (N_10689,N_6534,N_4542);
and U10690 (N_10690,N_5365,N_5507);
and U10691 (N_10691,N_4497,N_5913);
nor U10692 (N_10692,N_5957,N_4686);
or U10693 (N_10693,N_5775,N_7348);
nand U10694 (N_10694,N_6507,N_5666);
or U10695 (N_10695,N_6339,N_6425);
nand U10696 (N_10696,N_7241,N_4060);
and U10697 (N_10697,N_4852,N_6221);
nand U10698 (N_10698,N_7206,N_4225);
and U10699 (N_10699,N_4984,N_4569);
and U10700 (N_10700,N_6266,N_6592);
and U10701 (N_10701,N_7299,N_4796);
nand U10702 (N_10702,N_4509,N_7384);
xor U10703 (N_10703,N_6011,N_6875);
xor U10704 (N_10704,N_4337,N_4039);
and U10705 (N_10705,N_4043,N_6077);
nand U10706 (N_10706,N_7810,N_5551);
and U10707 (N_10707,N_5649,N_7757);
xor U10708 (N_10708,N_5782,N_5120);
and U10709 (N_10709,N_4204,N_7842);
nor U10710 (N_10710,N_7137,N_4210);
xnor U10711 (N_10711,N_4233,N_6968);
or U10712 (N_10712,N_6577,N_7144);
xor U10713 (N_10713,N_6950,N_5020);
nor U10714 (N_10714,N_6891,N_7407);
xor U10715 (N_10715,N_5069,N_4219);
xor U10716 (N_10716,N_7396,N_7423);
xnor U10717 (N_10717,N_6576,N_6744);
nor U10718 (N_10718,N_4634,N_4169);
xnor U10719 (N_10719,N_4319,N_4477);
nor U10720 (N_10720,N_7707,N_5106);
nor U10721 (N_10721,N_6884,N_5612);
nand U10722 (N_10722,N_7543,N_6048);
xnor U10723 (N_10723,N_4837,N_4709);
nor U10724 (N_10724,N_6240,N_6093);
nor U10725 (N_10725,N_5385,N_4301);
nand U10726 (N_10726,N_5542,N_6240);
xnor U10727 (N_10727,N_5190,N_6825);
or U10728 (N_10728,N_4022,N_4700);
nor U10729 (N_10729,N_5407,N_7961);
or U10730 (N_10730,N_7573,N_5826);
nand U10731 (N_10731,N_5703,N_5522);
and U10732 (N_10732,N_6668,N_4553);
nor U10733 (N_10733,N_4897,N_7268);
nor U10734 (N_10734,N_6041,N_6393);
xor U10735 (N_10735,N_4819,N_4890);
and U10736 (N_10736,N_4359,N_6779);
or U10737 (N_10737,N_4731,N_6996);
xor U10738 (N_10738,N_6269,N_5416);
or U10739 (N_10739,N_4161,N_7991);
xor U10740 (N_10740,N_5410,N_5765);
or U10741 (N_10741,N_4283,N_5484);
nand U10742 (N_10742,N_4971,N_5693);
xor U10743 (N_10743,N_7616,N_4172);
nand U10744 (N_10744,N_7837,N_7488);
nand U10745 (N_10745,N_4686,N_6615);
xnor U10746 (N_10746,N_7850,N_5620);
and U10747 (N_10747,N_7457,N_6116);
nand U10748 (N_10748,N_7118,N_4267);
nor U10749 (N_10749,N_5789,N_4029);
nor U10750 (N_10750,N_4116,N_4897);
xor U10751 (N_10751,N_4094,N_7552);
nand U10752 (N_10752,N_5233,N_4020);
and U10753 (N_10753,N_5178,N_4015);
nor U10754 (N_10754,N_6221,N_7565);
and U10755 (N_10755,N_6860,N_6132);
nand U10756 (N_10756,N_6043,N_4711);
or U10757 (N_10757,N_6386,N_6871);
nor U10758 (N_10758,N_6502,N_6103);
xnor U10759 (N_10759,N_5031,N_6587);
nand U10760 (N_10760,N_6269,N_7364);
and U10761 (N_10761,N_4252,N_5815);
or U10762 (N_10762,N_7554,N_7470);
xnor U10763 (N_10763,N_5557,N_4819);
or U10764 (N_10764,N_4105,N_7907);
nand U10765 (N_10765,N_6335,N_6456);
or U10766 (N_10766,N_7425,N_5150);
xor U10767 (N_10767,N_4508,N_6413);
nor U10768 (N_10768,N_5141,N_6510);
and U10769 (N_10769,N_7318,N_5999);
nand U10770 (N_10770,N_5315,N_4677);
or U10771 (N_10771,N_5540,N_4757);
xnor U10772 (N_10772,N_6381,N_6931);
nor U10773 (N_10773,N_7971,N_4382);
or U10774 (N_10774,N_7425,N_6301);
xor U10775 (N_10775,N_7264,N_5081);
and U10776 (N_10776,N_4326,N_4578);
nor U10777 (N_10777,N_4089,N_6688);
nor U10778 (N_10778,N_6478,N_6573);
and U10779 (N_10779,N_4825,N_6549);
nand U10780 (N_10780,N_4606,N_5314);
nor U10781 (N_10781,N_7984,N_4990);
or U10782 (N_10782,N_5822,N_7410);
and U10783 (N_10783,N_5450,N_6405);
nor U10784 (N_10784,N_5132,N_7342);
nand U10785 (N_10785,N_4216,N_7609);
xor U10786 (N_10786,N_7344,N_5573);
and U10787 (N_10787,N_6804,N_6934);
nor U10788 (N_10788,N_4551,N_7762);
or U10789 (N_10789,N_6337,N_7817);
or U10790 (N_10790,N_7555,N_5560);
xnor U10791 (N_10791,N_7461,N_7221);
nand U10792 (N_10792,N_4466,N_5407);
or U10793 (N_10793,N_5533,N_5312);
and U10794 (N_10794,N_7260,N_7478);
nand U10795 (N_10795,N_5686,N_4707);
nor U10796 (N_10796,N_7552,N_7367);
nand U10797 (N_10797,N_7605,N_5521);
or U10798 (N_10798,N_5356,N_6468);
nand U10799 (N_10799,N_7656,N_5191);
and U10800 (N_10800,N_6593,N_6837);
xnor U10801 (N_10801,N_4508,N_6826);
xnor U10802 (N_10802,N_6253,N_6705);
nand U10803 (N_10803,N_6472,N_7535);
nand U10804 (N_10804,N_4748,N_6043);
xnor U10805 (N_10805,N_7798,N_6534);
nand U10806 (N_10806,N_6260,N_7145);
xor U10807 (N_10807,N_7667,N_5119);
and U10808 (N_10808,N_5305,N_7738);
nor U10809 (N_10809,N_7437,N_5650);
nand U10810 (N_10810,N_7595,N_4929);
or U10811 (N_10811,N_6026,N_7457);
nor U10812 (N_10812,N_7546,N_4361);
nand U10813 (N_10813,N_4638,N_5587);
xor U10814 (N_10814,N_5517,N_4940);
nand U10815 (N_10815,N_5795,N_5693);
nor U10816 (N_10816,N_4972,N_4147);
and U10817 (N_10817,N_7587,N_5427);
and U10818 (N_10818,N_7155,N_7643);
or U10819 (N_10819,N_6656,N_5000);
nor U10820 (N_10820,N_5666,N_5174);
nor U10821 (N_10821,N_6517,N_7314);
or U10822 (N_10822,N_4073,N_7432);
xor U10823 (N_10823,N_5854,N_4553);
or U10824 (N_10824,N_5980,N_4586);
nor U10825 (N_10825,N_6772,N_6294);
xor U10826 (N_10826,N_7901,N_4593);
nand U10827 (N_10827,N_5798,N_4003);
nand U10828 (N_10828,N_5215,N_5363);
nor U10829 (N_10829,N_7917,N_6493);
nor U10830 (N_10830,N_4874,N_5754);
and U10831 (N_10831,N_5153,N_4720);
nor U10832 (N_10832,N_4842,N_4357);
xor U10833 (N_10833,N_4454,N_4238);
or U10834 (N_10834,N_7562,N_7882);
nor U10835 (N_10835,N_7806,N_7424);
nor U10836 (N_10836,N_7731,N_5696);
xor U10837 (N_10837,N_7841,N_6769);
xnor U10838 (N_10838,N_4423,N_7755);
nand U10839 (N_10839,N_7525,N_5524);
xor U10840 (N_10840,N_6458,N_4414);
and U10841 (N_10841,N_5237,N_5644);
xnor U10842 (N_10842,N_4193,N_7901);
nand U10843 (N_10843,N_4258,N_4293);
or U10844 (N_10844,N_6459,N_5944);
and U10845 (N_10845,N_6186,N_5070);
nor U10846 (N_10846,N_5699,N_7083);
nand U10847 (N_10847,N_5257,N_4703);
or U10848 (N_10848,N_4686,N_4922);
nor U10849 (N_10849,N_7322,N_7056);
nor U10850 (N_10850,N_4416,N_7960);
nand U10851 (N_10851,N_4457,N_4224);
nand U10852 (N_10852,N_5289,N_6157);
nand U10853 (N_10853,N_7070,N_7827);
nor U10854 (N_10854,N_4857,N_5131);
nor U10855 (N_10855,N_5251,N_4534);
xor U10856 (N_10856,N_7729,N_7766);
or U10857 (N_10857,N_4394,N_4405);
nand U10858 (N_10858,N_4201,N_4925);
nor U10859 (N_10859,N_4523,N_4294);
or U10860 (N_10860,N_5112,N_5784);
xnor U10861 (N_10861,N_7106,N_5783);
or U10862 (N_10862,N_7471,N_7289);
or U10863 (N_10863,N_7979,N_4615);
and U10864 (N_10864,N_6072,N_5023);
nand U10865 (N_10865,N_7365,N_5128);
nand U10866 (N_10866,N_5928,N_6094);
nand U10867 (N_10867,N_5910,N_4133);
or U10868 (N_10868,N_5275,N_6028);
nand U10869 (N_10869,N_4704,N_7164);
xnor U10870 (N_10870,N_4257,N_7408);
nand U10871 (N_10871,N_4524,N_5753);
nand U10872 (N_10872,N_7551,N_7628);
nor U10873 (N_10873,N_6589,N_7046);
and U10874 (N_10874,N_6245,N_5058);
xor U10875 (N_10875,N_6639,N_6170);
nand U10876 (N_10876,N_6795,N_6037);
nand U10877 (N_10877,N_5239,N_4107);
nor U10878 (N_10878,N_4750,N_5110);
nor U10879 (N_10879,N_5721,N_4010);
nor U10880 (N_10880,N_7626,N_5849);
nor U10881 (N_10881,N_4916,N_7759);
xnor U10882 (N_10882,N_5177,N_6100);
xor U10883 (N_10883,N_5367,N_7005);
or U10884 (N_10884,N_5990,N_6545);
xor U10885 (N_10885,N_4069,N_6062);
nor U10886 (N_10886,N_6458,N_7836);
and U10887 (N_10887,N_4389,N_6797);
xnor U10888 (N_10888,N_6444,N_6953);
and U10889 (N_10889,N_4843,N_5024);
and U10890 (N_10890,N_6531,N_7160);
nand U10891 (N_10891,N_5108,N_7841);
and U10892 (N_10892,N_4834,N_6608);
and U10893 (N_10893,N_4082,N_6119);
nor U10894 (N_10894,N_5256,N_7914);
xnor U10895 (N_10895,N_7548,N_6429);
or U10896 (N_10896,N_4233,N_4929);
nor U10897 (N_10897,N_5296,N_4763);
xor U10898 (N_10898,N_7155,N_5306);
or U10899 (N_10899,N_7650,N_4131);
and U10900 (N_10900,N_6136,N_4789);
nand U10901 (N_10901,N_6886,N_5485);
nor U10902 (N_10902,N_5157,N_6260);
nand U10903 (N_10903,N_7212,N_7994);
and U10904 (N_10904,N_5345,N_7188);
xor U10905 (N_10905,N_6569,N_6307);
nor U10906 (N_10906,N_7829,N_7793);
xnor U10907 (N_10907,N_5284,N_4109);
or U10908 (N_10908,N_4410,N_5075);
or U10909 (N_10909,N_5029,N_5652);
and U10910 (N_10910,N_5244,N_4266);
or U10911 (N_10911,N_6213,N_4576);
nand U10912 (N_10912,N_5018,N_4655);
nand U10913 (N_10913,N_4203,N_5850);
nand U10914 (N_10914,N_7373,N_7290);
xor U10915 (N_10915,N_4685,N_7313);
xor U10916 (N_10916,N_7019,N_4860);
or U10917 (N_10917,N_5205,N_5670);
or U10918 (N_10918,N_5873,N_4078);
nor U10919 (N_10919,N_5195,N_4350);
xnor U10920 (N_10920,N_5976,N_6427);
nand U10921 (N_10921,N_5543,N_4667);
nand U10922 (N_10922,N_4913,N_7858);
nor U10923 (N_10923,N_4566,N_6032);
xnor U10924 (N_10924,N_7643,N_7040);
xnor U10925 (N_10925,N_7477,N_6168);
nor U10926 (N_10926,N_7062,N_5914);
nand U10927 (N_10927,N_6419,N_4435);
xnor U10928 (N_10928,N_7700,N_4375);
xnor U10929 (N_10929,N_7286,N_5774);
nand U10930 (N_10930,N_5554,N_4959);
and U10931 (N_10931,N_7113,N_5213);
and U10932 (N_10932,N_5827,N_4417);
or U10933 (N_10933,N_4170,N_7695);
or U10934 (N_10934,N_4230,N_6061);
or U10935 (N_10935,N_4739,N_7104);
nand U10936 (N_10936,N_5364,N_6349);
xnor U10937 (N_10937,N_6858,N_5027);
or U10938 (N_10938,N_5885,N_5363);
xor U10939 (N_10939,N_4439,N_6215);
and U10940 (N_10940,N_7960,N_6602);
nor U10941 (N_10941,N_4219,N_7248);
nand U10942 (N_10942,N_4627,N_5502);
or U10943 (N_10943,N_4581,N_4369);
or U10944 (N_10944,N_5876,N_4144);
or U10945 (N_10945,N_5665,N_5242);
nor U10946 (N_10946,N_4497,N_5271);
nor U10947 (N_10947,N_4086,N_6762);
nor U10948 (N_10948,N_7160,N_6640);
nor U10949 (N_10949,N_6345,N_6046);
nand U10950 (N_10950,N_4761,N_7652);
nor U10951 (N_10951,N_4346,N_4653);
xnor U10952 (N_10952,N_6064,N_7077);
nor U10953 (N_10953,N_7777,N_6513);
xor U10954 (N_10954,N_6100,N_4569);
nand U10955 (N_10955,N_7253,N_5630);
xor U10956 (N_10956,N_4093,N_5607);
and U10957 (N_10957,N_7548,N_7859);
nand U10958 (N_10958,N_7618,N_5462);
nor U10959 (N_10959,N_4415,N_4113);
xor U10960 (N_10960,N_5906,N_6192);
and U10961 (N_10961,N_5927,N_5410);
or U10962 (N_10962,N_5441,N_4088);
and U10963 (N_10963,N_5683,N_6892);
or U10964 (N_10964,N_7121,N_6948);
xor U10965 (N_10965,N_5462,N_5291);
or U10966 (N_10966,N_5987,N_5880);
xnor U10967 (N_10967,N_6155,N_7454);
or U10968 (N_10968,N_5223,N_7900);
nor U10969 (N_10969,N_6272,N_7559);
xnor U10970 (N_10970,N_6752,N_5776);
xnor U10971 (N_10971,N_7271,N_4094);
or U10972 (N_10972,N_4774,N_7563);
nand U10973 (N_10973,N_4321,N_7852);
xnor U10974 (N_10974,N_6587,N_6487);
and U10975 (N_10975,N_7044,N_5730);
and U10976 (N_10976,N_7626,N_7666);
xor U10977 (N_10977,N_7892,N_5353);
nand U10978 (N_10978,N_5751,N_6050);
nand U10979 (N_10979,N_6192,N_5156);
or U10980 (N_10980,N_5702,N_4584);
or U10981 (N_10981,N_7449,N_7444);
nand U10982 (N_10982,N_4472,N_5902);
nor U10983 (N_10983,N_4066,N_6755);
or U10984 (N_10984,N_7948,N_7279);
and U10985 (N_10985,N_4110,N_5121);
xnor U10986 (N_10986,N_7468,N_4700);
nand U10987 (N_10987,N_7860,N_5595);
and U10988 (N_10988,N_7042,N_4037);
and U10989 (N_10989,N_4071,N_5870);
nand U10990 (N_10990,N_7896,N_5913);
and U10991 (N_10991,N_7713,N_7845);
or U10992 (N_10992,N_4268,N_5167);
or U10993 (N_10993,N_4633,N_7136);
nand U10994 (N_10994,N_6965,N_6802);
and U10995 (N_10995,N_7648,N_6309);
and U10996 (N_10996,N_5765,N_6040);
nor U10997 (N_10997,N_4283,N_6448);
or U10998 (N_10998,N_7780,N_5505);
xor U10999 (N_10999,N_4882,N_6313);
nand U11000 (N_11000,N_5978,N_6627);
nand U11001 (N_11001,N_5453,N_6551);
xnor U11002 (N_11002,N_5355,N_4755);
xor U11003 (N_11003,N_5986,N_5639);
nor U11004 (N_11004,N_6568,N_5107);
and U11005 (N_11005,N_6319,N_7676);
xnor U11006 (N_11006,N_4291,N_5272);
or U11007 (N_11007,N_4035,N_4809);
or U11008 (N_11008,N_7896,N_6223);
nand U11009 (N_11009,N_4729,N_6349);
nor U11010 (N_11010,N_6395,N_4400);
xor U11011 (N_11011,N_6021,N_5669);
nand U11012 (N_11012,N_5912,N_4544);
nand U11013 (N_11013,N_5846,N_7358);
nand U11014 (N_11014,N_6749,N_5913);
xnor U11015 (N_11015,N_6060,N_6037);
nor U11016 (N_11016,N_5886,N_4424);
or U11017 (N_11017,N_7235,N_6546);
and U11018 (N_11018,N_6067,N_7941);
nor U11019 (N_11019,N_4439,N_4522);
xor U11020 (N_11020,N_4000,N_5973);
nor U11021 (N_11021,N_6155,N_7011);
xor U11022 (N_11022,N_6389,N_6731);
nand U11023 (N_11023,N_5328,N_5025);
and U11024 (N_11024,N_4503,N_5578);
xnor U11025 (N_11025,N_5466,N_6604);
xor U11026 (N_11026,N_5824,N_4730);
nor U11027 (N_11027,N_6417,N_7382);
xnor U11028 (N_11028,N_5327,N_5506);
nor U11029 (N_11029,N_6133,N_7526);
or U11030 (N_11030,N_5648,N_6746);
or U11031 (N_11031,N_4022,N_6852);
nor U11032 (N_11032,N_5673,N_6277);
xor U11033 (N_11033,N_4426,N_7781);
nand U11034 (N_11034,N_5123,N_4594);
xor U11035 (N_11035,N_5524,N_5061);
or U11036 (N_11036,N_7953,N_4150);
or U11037 (N_11037,N_7537,N_7678);
and U11038 (N_11038,N_4364,N_6982);
nor U11039 (N_11039,N_4694,N_7676);
nor U11040 (N_11040,N_7376,N_6741);
or U11041 (N_11041,N_5493,N_7133);
or U11042 (N_11042,N_5102,N_6745);
xor U11043 (N_11043,N_7281,N_5118);
nand U11044 (N_11044,N_5641,N_6085);
nand U11045 (N_11045,N_6246,N_5557);
and U11046 (N_11046,N_6958,N_6720);
and U11047 (N_11047,N_5353,N_7569);
nand U11048 (N_11048,N_4865,N_5233);
xor U11049 (N_11049,N_5608,N_5589);
nand U11050 (N_11050,N_7240,N_6026);
nor U11051 (N_11051,N_5697,N_7282);
or U11052 (N_11052,N_6070,N_5429);
nand U11053 (N_11053,N_6770,N_6471);
and U11054 (N_11054,N_7720,N_7002);
or U11055 (N_11055,N_6920,N_7062);
nand U11056 (N_11056,N_6971,N_4305);
and U11057 (N_11057,N_7916,N_5238);
nand U11058 (N_11058,N_4996,N_4758);
nor U11059 (N_11059,N_6574,N_5895);
xnor U11060 (N_11060,N_5192,N_6674);
or U11061 (N_11061,N_7793,N_7077);
and U11062 (N_11062,N_4165,N_5483);
nor U11063 (N_11063,N_5739,N_7666);
nor U11064 (N_11064,N_5807,N_6139);
nor U11065 (N_11065,N_5493,N_4919);
nor U11066 (N_11066,N_5035,N_7175);
and U11067 (N_11067,N_7220,N_4024);
nor U11068 (N_11068,N_6051,N_7444);
and U11069 (N_11069,N_7162,N_6773);
nand U11070 (N_11070,N_4420,N_4205);
nor U11071 (N_11071,N_6034,N_4859);
or U11072 (N_11072,N_5244,N_4913);
nor U11073 (N_11073,N_6690,N_4500);
nor U11074 (N_11074,N_4524,N_7415);
or U11075 (N_11075,N_4809,N_6165);
nand U11076 (N_11076,N_4885,N_5265);
or U11077 (N_11077,N_6516,N_7332);
xor U11078 (N_11078,N_4923,N_7257);
nor U11079 (N_11079,N_5610,N_7688);
nor U11080 (N_11080,N_7321,N_6156);
nand U11081 (N_11081,N_5736,N_4950);
nor U11082 (N_11082,N_5624,N_5933);
nand U11083 (N_11083,N_6374,N_7239);
nand U11084 (N_11084,N_7738,N_5952);
nor U11085 (N_11085,N_6202,N_4347);
nor U11086 (N_11086,N_6889,N_4196);
nand U11087 (N_11087,N_7273,N_6215);
or U11088 (N_11088,N_5348,N_4422);
xnor U11089 (N_11089,N_4853,N_5371);
or U11090 (N_11090,N_5499,N_6399);
xnor U11091 (N_11091,N_4481,N_5770);
xnor U11092 (N_11092,N_5945,N_6610);
nand U11093 (N_11093,N_5226,N_5612);
xor U11094 (N_11094,N_4245,N_6753);
nand U11095 (N_11095,N_5190,N_4152);
xor U11096 (N_11096,N_5562,N_4497);
nor U11097 (N_11097,N_5842,N_4685);
and U11098 (N_11098,N_4544,N_6549);
nand U11099 (N_11099,N_7094,N_7230);
nand U11100 (N_11100,N_6418,N_5775);
nor U11101 (N_11101,N_5260,N_4841);
xnor U11102 (N_11102,N_5582,N_6774);
or U11103 (N_11103,N_7033,N_4416);
xnor U11104 (N_11104,N_5220,N_4765);
or U11105 (N_11105,N_4420,N_4714);
nand U11106 (N_11106,N_5500,N_7709);
nor U11107 (N_11107,N_5350,N_6410);
and U11108 (N_11108,N_6088,N_5799);
or U11109 (N_11109,N_4641,N_5907);
and U11110 (N_11110,N_4866,N_6294);
and U11111 (N_11111,N_6268,N_5699);
nor U11112 (N_11112,N_6584,N_5579);
or U11113 (N_11113,N_5126,N_6355);
or U11114 (N_11114,N_7088,N_4122);
and U11115 (N_11115,N_6457,N_6339);
xor U11116 (N_11116,N_5461,N_6535);
xnor U11117 (N_11117,N_4002,N_7068);
xnor U11118 (N_11118,N_4375,N_6830);
and U11119 (N_11119,N_4578,N_4390);
and U11120 (N_11120,N_6597,N_4419);
nand U11121 (N_11121,N_5317,N_4449);
nor U11122 (N_11122,N_6653,N_5451);
or U11123 (N_11123,N_5815,N_6944);
nand U11124 (N_11124,N_7173,N_4244);
or U11125 (N_11125,N_6477,N_5298);
xnor U11126 (N_11126,N_6247,N_7078);
xor U11127 (N_11127,N_4121,N_5719);
nor U11128 (N_11128,N_4485,N_7610);
xnor U11129 (N_11129,N_5458,N_4236);
or U11130 (N_11130,N_7475,N_7437);
or U11131 (N_11131,N_6985,N_5513);
and U11132 (N_11132,N_5037,N_5033);
nand U11133 (N_11133,N_6234,N_6462);
nor U11134 (N_11134,N_5866,N_4972);
and U11135 (N_11135,N_6080,N_6160);
xnor U11136 (N_11136,N_4316,N_4325);
xor U11137 (N_11137,N_5241,N_6747);
xnor U11138 (N_11138,N_4170,N_6500);
and U11139 (N_11139,N_5002,N_4339);
and U11140 (N_11140,N_4131,N_5389);
nor U11141 (N_11141,N_5400,N_7247);
and U11142 (N_11142,N_5498,N_4745);
and U11143 (N_11143,N_6514,N_7878);
nand U11144 (N_11144,N_6104,N_7973);
nand U11145 (N_11145,N_7634,N_4097);
nand U11146 (N_11146,N_7473,N_5835);
nand U11147 (N_11147,N_4551,N_4620);
xor U11148 (N_11148,N_6306,N_4226);
or U11149 (N_11149,N_5742,N_4221);
or U11150 (N_11150,N_4829,N_5518);
nor U11151 (N_11151,N_6000,N_7640);
xnor U11152 (N_11152,N_5937,N_7706);
nand U11153 (N_11153,N_7944,N_5312);
nor U11154 (N_11154,N_4323,N_7666);
nor U11155 (N_11155,N_4740,N_7402);
nand U11156 (N_11156,N_4451,N_4967);
or U11157 (N_11157,N_7311,N_6443);
nor U11158 (N_11158,N_7873,N_6131);
nor U11159 (N_11159,N_6183,N_6863);
or U11160 (N_11160,N_4587,N_5827);
nand U11161 (N_11161,N_4946,N_6284);
xor U11162 (N_11162,N_6970,N_6888);
nand U11163 (N_11163,N_4668,N_5279);
xor U11164 (N_11164,N_4558,N_6112);
xor U11165 (N_11165,N_4882,N_5929);
and U11166 (N_11166,N_4714,N_6245);
nand U11167 (N_11167,N_4517,N_4110);
nand U11168 (N_11168,N_6399,N_5312);
xnor U11169 (N_11169,N_5042,N_5259);
nand U11170 (N_11170,N_4125,N_7016);
and U11171 (N_11171,N_6664,N_6049);
nand U11172 (N_11172,N_4606,N_7297);
or U11173 (N_11173,N_5945,N_7662);
nand U11174 (N_11174,N_5636,N_4492);
nor U11175 (N_11175,N_7584,N_7499);
nand U11176 (N_11176,N_4411,N_7069);
nand U11177 (N_11177,N_4587,N_7646);
and U11178 (N_11178,N_6278,N_6651);
xnor U11179 (N_11179,N_5078,N_4582);
nand U11180 (N_11180,N_5453,N_7689);
nor U11181 (N_11181,N_6330,N_4334);
nand U11182 (N_11182,N_7185,N_6765);
and U11183 (N_11183,N_5483,N_4799);
xor U11184 (N_11184,N_7983,N_7413);
or U11185 (N_11185,N_5029,N_6470);
or U11186 (N_11186,N_5859,N_7254);
nand U11187 (N_11187,N_4054,N_6224);
xor U11188 (N_11188,N_7577,N_4082);
nor U11189 (N_11189,N_7640,N_6196);
nor U11190 (N_11190,N_6458,N_7337);
and U11191 (N_11191,N_7275,N_5567);
nor U11192 (N_11192,N_5531,N_4138);
or U11193 (N_11193,N_6387,N_5720);
or U11194 (N_11194,N_7968,N_4761);
and U11195 (N_11195,N_6325,N_5841);
nand U11196 (N_11196,N_5054,N_5144);
or U11197 (N_11197,N_4126,N_4223);
xnor U11198 (N_11198,N_7935,N_7111);
or U11199 (N_11199,N_7686,N_6504);
nand U11200 (N_11200,N_7063,N_4943);
xor U11201 (N_11201,N_7875,N_4193);
nor U11202 (N_11202,N_6316,N_5155);
nor U11203 (N_11203,N_4007,N_4401);
nor U11204 (N_11204,N_7351,N_4451);
nor U11205 (N_11205,N_6586,N_6874);
xnor U11206 (N_11206,N_4640,N_7719);
xor U11207 (N_11207,N_5573,N_7985);
nor U11208 (N_11208,N_7494,N_5022);
and U11209 (N_11209,N_5170,N_7115);
or U11210 (N_11210,N_5250,N_6381);
xnor U11211 (N_11211,N_6521,N_4030);
nand U11212 (N_11212,N_6048,N_4997);
and U11213 (N_11213,N_5764,N_5405);
and U11214 (N_11214,N_4860,N_6632);
xnor U11215 (N_11215,N_7920,N_4218);
xor U11216 (N_11216,N_6170,N_6531);
and U11217 (N_11217,N_4345,N_5847);
nand U11218 (N_11218,N_5107,N_4361);
and U11219 (N_11219,N_6409,N_6927);
or U11220 (N_11220,N_6967,N_6743);
or U11221 (N_11221,N_6323,N_5136);
or U11222 (N_11222,N_7452,N_5756);
nand U11223 (N_11223,N_5691,N_5398);
nor U11224 (N_11224,N_5401,N_5420);
nor U11225 (N_11225,N_7966,N_4559);
and U11226 (N_11226,N_7569,N_7062);
xor U11227 (N_11227,N_6748,N_6437);
nor U11228 (N_11228,N_7812,N_7365);
and U11229 (N_11229,N_4925,N_7754);
xnor U11230 (N_11230,N_7681,N_6392);
nand U11231 (N_11231,N_5611,N_6996);
nand U11232 (N_11232,N_4031,N_6212);
nor U11233 (N_11233,N_7972,N_5274);
nand U11234 (N_11234,N_7668,N_4235);
nand U11235 (N_11235,N_4898,N_7369);
nor U11236 (N_11236,N_7789,N_7735);
xor U11237 (N_11237,N_4819,N_7771);
xor U11238 (N_11238,N_4582,N_6449);
nor U11239 (N_11239,N_4941,N_4536);
or U11240 (N_11240,N_7385,N_5632);
nand U11241 (N_11241,N_5632,N_5910);
or U11242 (N_11242,N_4350,N_7045);
or U11243 (N_11243,N_7448,N_6956);
nor U11244 (N_11244,N_5741,N_5790);
xor U11245 (N_11245,N_7178,N_5942);
or U11246 (N_11246,N_4025,N_7048);
nand U11247 (N_11247,N_7717,N_7532);
or U11248 (N_11248,N_5550,N_7380);
nand U11249 (N_11249,N_5727,N_4082);
xor U11250 (N_11250,N_7530,N_7004);
or U11251 (N_11251,N_7499,N_4392);
nor U11252 (N_11252,N_5183,N_7592);
and U11253 (N_11253,N_7132,N_5209);
or U11254 (N_11254,N_6226,N_5611);
or U11255 (N_11255,N_7893,N_4809);
xor U11256 (N_11256,N_7399,N_4790);
nand U11257 (N_11257,N_6513,N_6771);
nor U11258 (N_11258,N_5822,N_6235);
xnor U11259 (N_11259,N_7311,N_4221);
or U11260 (N_11260,N_6433,N_4349);
or U11261 (N_11261,N_5475,N_5280);
or U11262 (N_11262,N_4188,N_5064);
nor U11263 (N_11263,N_7978,N_5484);
nand U11264 (N_11264,N_7489,N_7581);
or U11265 (N_11265,N_7592,N_4432);
xor U11266 (N_11266,N_6251,N_4803);
nand U11267 (N_11267,N_6246,N_7798);
or U11268 (N_11268,N_5516,N_5838);
and U11269 (N_11269,N_7416,N_7392);
or U11270 (N_11270,N_7348,N_6733);
or U11271 (N_11271,N_5240,N_7882);
xor U11272 (N_11272,N_6441,N_5321);
or U11273 (N_11273,N_5850,N_5840);
or U11274 (N_11274,N_5684,N_7871);
xnor U11275 (N_11275,N_6860,N_4781);
xnor U11276 (N_11276,N_4211,N_6317);
nor U11277 (N_11277,N_5692,N_5502);
xor U11278 (N_11278,N_4962,N_6476);
nor U11279 (N_11279,N_4054,N_4438);
nand U11280 (N_11280,N_4655,N_4031);
and U11281 (N_11281,N_6493,N_6876);
xnor U11282 (N_11282,N_5584,N_4028);
nand U11283 (N_11283,N_4720,N_6472);
or U11284 (N_11284,N_5507,N_5354);
nand U11285 (N_11285,N_6775,N_5775);
xor U11286 (N_11286,N_6002,N_6974);
xnor U11287 (N_11287,N_7803,N_5289);
xnor U11288 (N_11288,N_7130,N_7006);
xor U11289 (N_11289,N_6733,N_7142);
and U11290 (N_11290,N_5159,N_7203);
xor U11291 (N_11291,N_5630,N_4968);
nor U11292 (N_11292,N_6176,N_4750);
nor U11293 (N_11293,N_6173,N_6444);
xor U11294 (N_11294,N_7523,N_5818);
nor U11295 (N_11295,N_6906,N_5714);
xor U11296 (N_11296,N_5878,N_5580);
or U11297 (N_11297,N_5470,N_5142);
nand U11298 (N_11298,N_6267,N_7303);
nor U11299 (N_11299,N_7014,N_4563);
or U11300 (N_11300,N_7844,N_4014);
nand U11301 (N_11301,N_4591,N_7623);
xnor U11302 (N_11302,N_4374,N_5994);
nor U11303 (N_11303,N_6772,N_4561);
and U11304 (N_11304,N_4269,N_5877);
or U11305 (N_11305,N_4540,N_4360);
nand U11306 (N_11306,N_6978,N_7056);
nor U11307 (N_11307,N_7918,N_5738);
xor U11308 (N_11308,N_7396,N_7107);
xor U11309 (N_11309,N_5206,N_4544);
nor U11310 (N_11310,N_7238,N_7980);
and U11311 (N_11311,N_7192,N_4214);
nand U11312 (N_11312,N_6730,N_4100);
xor U11313 (N_11313,N_7577,N_7099);
nor U11314 (N_11314,N_7381,N_5350);
xor U11315 (N_11315,N_7777,N_7413);
nor U11316 (N_11316,N_7893,N_6700);
nor U11317 (N_11317,N_7552,N_5323);
xor U11318 (N_11318,N_7251,N_4196);
and U11319 (N_11319,N_7443,N_5385);
nand U11320 (N_11320,N_7617,N_4617);
or U11321 (N_11321,N_5578,N_6359);
xor U11322 (N_11322,N_5125,N_7963);
xnor U11323 (N_11323,N_5995,N_4407);
xnor U11324 (N_11324,N_6480,N_4287);
nand U11325 (N_11325,N_5613,N_4478);
xor U11326 (N_11326,N_7947,N_5278);
nor U11327 (N_11327,N_7825,N_4003);
xor U11328 (N_11328,N_6594,N_4248);
nand U11329 (N_11329,N_6718,N_7951);
nand U11330 (N_11330,N_5141,N_6668);
xor U11331 (N_11331,N_4793,N_6292);
nor U11332 (N_11332,N_4226,N_6400);
nand U11333 (N_11333,N_5043,N_6164);
nor U11334 (N_11334,N_4593,N_5735);
nand U11335 (N_11335,N_6460,N_6625);
xnor U11336 (N_11336,N_5657,N_5759);
or U11337 (N_11337,N_5136,N_6918);
nor U11338 (N_11338,N_5113,N_5171);
xor U11339 (N_11339,N_7287,N_5996);
nor U11340 (N_11340,N_5522,N_5885);
nand U11341 (N_11341,N_5207,N_6992);
xor U11342 (N_11342,N_6499,N_6650);
or U11343 (N_11343,N_7244,N_5711);
and U11344 (N_11344,N_5609,N_6667);
and U11345 (N_11345,N_4182,N_5543);
xnor U11346 (N_11346,N_5848,N_5393);
nand U11347 (N_11347,N_6665,N_7326);
xor U11348 (N_11348,N_5428,N_7010);
xor U11349 (N_11349,N_6664,N_6646);
xnor U11350 (N_11350,N_7926,N_6865);
nand U11351 (N_11351,N_6273,N_5358);
xor U11352 (N_11352,N_4328,N_4940);
and U11353 (N_11353,N_6267,N_4559);
nor U11354 (N_11354,N_7203,N_4850);
and U11355 (N_11355,N_4786,N_7205);
and U11356 (N_11356,N_5008,N_7999);
nand U11357 (N_11357,N_5366,N_7881);
xnor U11358 (N_11358,N_7088,N_5312);
nor U11359 (N_11359,N_4552,N_4570);
nor U11360 (N_11360,N_4108,N_7800);
or U11361 (N_11361,N_4302,N_4863);
nand U11362 (N_11362,N_6885,N_6061);
and U11363 (N_11363,N_7737,N_4701);
or U11364 (N_11364,N_7778,N_6153);
xnor U11365 (N_11365,N_6575,N_5669);
and U11366 (N_11366,N_5576,N_7466);
nand U11367 (N_11367,N_6979,N_7279);
xor U11368 (N_11368,N_6835,N_7103);
nor U11369 (N_11369,N_7641,N_4088);
nor U11370 (N_11370,N_5165,N_7442);
xor U11371 (N_11371,N_5478,N_7895);
nand U11372 (N_11372,N_6200,N_5141);
or U11373 (N_11373,N_6912,N_5229);
or U11374 (N_11374,N_4702,N_7847);
nand U11375 (N_11375,N_6811,N_7502);
nand U11376 (N_11376,N_6299,N_6348);
nor U11377 (N_11377,N_7068,N_4086);
or U11378 (N_11378,N_5484,N_4365);
nand U11379 (N_11379,N_7627,N_7528);
nand U11380 (N_11380,N_4824,N_5516);
nand U11381 (N_11381,N_7225,N_5264);
xor U11382 (N_11382,N_4832,N_5969);
nand U11383 (N_11383,N_7057,N_7306);
xor U11384 (N_11384,N_4983,N_7233);
nand U11385 (N_11385,N_7129,N_5711);
or U11386 (N_11386,N_5691,N_5134);
and U11387 (N_11387,N_6114,N_6591);
and U11388 (N_11388,N_7939,N_4383);
and U11389 (N_11389,N_6743,N_7286);
or U11390 (N_11390,N_7660,N_6623);
xnor U11391 (N_11391,N_6645,N_4033);
and U11392 (N_11392,N_5681,N_6347);
nor U11393 (N_11393,N_6435,N_5599);
or U11394 (N_11394,N_5676,N_7278);
and U11395 (N_11395,N_4045,N_6945);
or U11396 (N_11396,N_7688,N_6853);
xnor U11397 (N_11397,N_6810,N_5817);
xor U11398 (N_11398,N_7719,N_4128);
nor U11399 (N_11399,N_7460,N_7177);
and U11400 (N_11400,N_4603,N_7870);
or U11401 (N_11401,N_4011,N_5805);
nand U11402 (N_11402,N_4357,N_4879);
and U11403 (N_11403,N_7195,N_6596);
or U11404 (N_11404,N_6326,N_4253);
or U11405 (N_11405,N_5767,N_6460);
nor U11406 (N_11406,N_6081,N_6528);
or U11407 (N_11407,N_5658,N_4445);
nor U11408 (N_11408,N_6922,N_6849);
nand U11409 (N_11409,N_7214,N_6537);
xor U11410 (N_11410,N_6214,N_6180);
and U11411 (N_11411,N_6410,N_4652);
nor U11412 (N_11412,N_7127,N_7744);
nand U11413 (N_11413,N_5819,N_7165);
nor U11414 (N_11414,N_7549,N_7172);
nor U11415 (N_11415,N_7382,N_7282);
xor U11416 (N_11416,N_7715,N_5173);
nor U11417 (N_11417,N_7729,N_7476);
and U11418 (N_11418,N_5066,N_4798);
nor U11419 (N_11419,N_4284,N_6080);
xor U11420 (N_11420,N_5640,N_6543);
or U11421 (N_11421,N_4247,N_5067);
nand U11422 (N_11422,N_7230,N_6297);
or U11423 (N_11423,N_5405,N_5557);
nand U11424 (N_11424,N_7867,N_7352);
or U11425 (N_11425,N_7092,N_7321);
nand U11426 (N_11426,N_5908,N_7963);
or U11427 (N_11427,N_4377,N_5358);
or U11428 (N_11428,N_5409,N_5629);
nor U11429 (N_11429,N_6752,N_6440);
nor U11430 (N_11430,N_4156,N_6262);
nor U11431 (N_11431,N_4053,N_7537);
or U11432 (N_11432,N_6889,N_5426);
nor U11433 (N_11433,N_5952,N_5397);
and U11434 (N_11434,N_4738,N_5459);
nand U11435 (N_11435,N_6143,N_7080);
xnor U11436 (N_11436,N_4565,N_6721);
and U11437 (N_11437,N_6932,N_7143);
nor U11438 (N_11438,N_6246,N_5758);
or U11439 (N_11439,N_4190,N_7185);
nand U11440 (N_11440,N_7885,N_7566);
nor U11441 (N_11441,N_4887,N_4197);
xnor U11442 (N_11442,N_4781,N_4004);
nor U11443 (N_11443,N_4573,N_7789);
nand U11444 (N_11444,N_4345,N_6800);
nand U11445 (N_11445,N_7191,N_5681);
nor U11446 (N_11446,N_5207,N_4087);
nand U11447 (N_11447,N_7037,N_7644);
xor U11448 (N_11448,N_5145,N_6222);
and U11449 (N_11449,N_6000,N_7580);
or U11450 (N_11450,N_5418,N_4014);
and U11451 (N_11451,N_5452,N_6614);
or U11452 (N_11452,N_5437,N_5805);
nand U11453 (N_11453,N_6407,N_4826);
or U11454 (N_11454,N_4834,N_5002);
nand U11455 (N_11455,N_7473,N_5123);
nand U11456 (N_11456,N_7777,N_5898);
nor U11457 (N_11457,N_5693,N_7259);
nor U11458 (N_11458,N_6003,N_7145);
xor U11459 (N_11459,N_4576,N_4802);
or U11460 (N_11460,N_5692,N_5879);
xnor U11461 (N_11461,N_7743,N_7361);
nand U11462 (N_11462,N_5168,N_7485);
or U11463 (N_11463,N_7512,N_5966);
and U11464 (N_11464,N_6260,N_5011);
xnor U11465 (N_11465,N_4829,N_5429);
nor U11466 (N_11466,N_4637,N_4587);
nand U11467 (N_11467,N_5814,N_4146);
xnor U11468 (N_11468,N_4153,N_7650);
xor U11469 (N_11469,N_7739,N_4473);
or U11470 (N_11470,N_6866,N_7913);
or U11471 (N_11471,N_7058,N_6907);
nand U11472 (N_11472,N_4522,N_7667);
xnor U11473 (N_11473,N_4208,N_6173);
xor U11474 (N_11474,N_6900,N_4012);
xnor U11475 (N_11475,N_4673,N_6805);
nand U11476 (N_11476,N_6553,N_5523);
nand U11477 (N_11477,N_7296,N_7391);
and U11478 (N_11478,N_5342,N_4281);
nand U11479 (N_11479,N_5527,N_6826);
and U11480 (N_11480,N_6664,N_6255);
xor U11481 (N_11481,N_6727,N_4273);
xnor U11482 (N_11482,N_4944,N_5139);
or U11483 (N_11483,N_6717,N_7964);
and U11484 (N_11484,N_7673,N_7126);
nand U11485 (N_11485,N_5466,N_6361);
and U11486 (N_11486,N_7466,N_7349);
and U11487 (N_11487,N_4099,N_6989);
and U11488 (N_11488,N_7757,N_6815);
nand U11489 (N_11489,N_6699,N_6190);
xnor U11490 (N_11490,N_7236,N_6709);
and U11491 (N_11491,N_4900,N_7437);
or U11492 (N_11492,N_4147,N_4206);
nand U11493 (N_11493,N_6832,N_4082);
and U11494 (N_11494,N_6714,N_4342);
xnor U11495 (N_11495,N_4629,N_4542);
or U11496 (N_11496,N_6982,N_4284);
xnor U11497 (N_11497,N_7882,N_7362);
or U11498 (N_11498,N_4867,N_6938);
nand U11499 (N_11499,N_4392,N_5701);
nor U11500 (N_11500,N_4152,N_7391);
nor U11501 (N_11501,N_7823,N_4225);
or U11502 (N_11502,N_6515,N_5582);
xor U11503 (N_11503,N_4964,N_5127);
and U11504 (N_11504,N_6668,N_4904);
and U11505 (N_11505,N_4311,N_4021);
nand U11506 (N_11506,N_7445,N_6251);
or U11507 (N_11507,N_4568,N_4576);
xnor U11508 (N_11508,N_5461,N_6337);
xnor U11509 (N_11509,N_6614,N_4800);
nor U11510 (N_11510,N_7477,N_7924);
or U11511 (N_11511,N_5925,N_5120);
and U11512 (N_11512,N_4015,N_6988);
xor U11513 (N_11513,N_4362,N_4489);
and U11514 (N_11514,N_5441,N_4026);
or U11515 (N_11515,N_7148,N_4838);
xor U11516 (N_11516,N_6869,N_6281);
or U11517 (N_11517,N_7193,N_4666);
nor U11518 (N_11518,N_6903,N_7177);
and U11519 (N_11519,N_6663,N_7050);
xnor U11520 (N_11520,N_5044,N_4541);
and U11521 (N_11521,N_6564,N_5848);
nor U11522 (N_11522,N_5769,N_7857);
nor U11523 (N_11523,N_7358,N_4444);
xor U11524 (N_11524,N_7395,N_5681);
or U11525 (N_11525,N_4283,N_4704);
and U11526 (N_11526,N_4067,N_6007);
nand U11527 (N_11527,N_7881,N_5905);
and U11528 (N_11528,N_5445,N_6326);
nand U11529 (N_11529,N_6775,N_6768);
and U11530 (N_11530,N_7768,N_7947);
and U11531 (N_11531,N_7068,N_5831);
or U11532 (N_11532,N_6145,N_6827);
or U11533 (N_11533,N_6569,N_4003);
or U11534 (N_11534,N_7497,N_4775);
nand U11535 (N_11535,N_5322,N_7615);
nand U11536 (N_11536,N_7576,N_7288);
xnor U11537 (N_11537,N_5536,N_7381);
nor U11538 (N_11538,N_5135,N_6231);
xor U11539 (N_11539,N_4498,N_7324);
nor U11540 (N_11540,N_6529,N_5744);
xor U11541 (N_11541,N_6816,N_5311);
and U11542 (N_11542,N_7545,N_6094);
xnor U11543 (N_11543,N_4798,N_7095);
xnor U11544 (N_11544,N_4524,N_5525);
and U11545 (N_11545,N_7241,N_5809);
or U11546 (N_11546,N_7630,N_7827);
nand U11547 (N_11547,N_5598,N_4737);
nand U11548 (N_11548,N_4369,N_7448);
or U11549 (N_11549,N_6822,N_4399);
nand U11550 (N_11550,N_7646,N_5249);
and U11551 (N_11551,N_5230,N_7114);
nand U11552 (N_11552,N_6446,N_4813);
or U11553 (N_11553,N_7501,N_6555);
nor U11554 (N_11554,N_4835,N_7279);
nand U11555 (N_11555,N_7293,N_5293);
nor U11556 (N_11556,N_4858,N_7170);
nor U11557 (N_11557,N_7243,N_4100);
or U11558 (N_11558,N_4285,N_5198);
nand U11559 (N_11559,N_7925,N_6142);
or U11560 (N_11560,N_4431,N_5988);
nor U11561 (N_11561,N_6080,N_4747);
xnor U11562 (N_11562,N_6458,N_7287);
or U11563 (N_11563,N_7487,N_4164);
and U11564 (N_11564,N_6366,N_7597);
nor U11565 (N_11565,N_6282,N_4442);
xnor U11566 (N_11566,N_7738,N_6716);
or U11567 (N_11567,N_7428,N_6188);
and U11568 (N_11568,N_6531,N_7272);
nand U11569 (N_11569,N_7291,N_6790);
nor U11570 (N_11570,N_6305,N_6808);
nor U11571 (N_11571,N_5735,N_4768);
or U11572 (N_11572,N_4488,N_6942);
and U11573 (N_11573,N_6894,N_5983);
xnor U11574 (N_11574,N_6906,N_4423);
nand U11575 (N_11575,N_5041,N_6023);
or U11576 (N_11576,N_4167,N_4988);
and U11577 (N_11577,N_7321,N_7208);
and U11578 (N_11578,N_6445,N_4443);
xor U11579 (N_11579,N_5602,N_5196);
or U11580 (N_11580,N_4389,N_7397);
or U11581 (N_11581,N_4121,N_7302);
and U11582 (N_11582,N_4675,N_6749);
nand U11583 (N_11583,N_7062,N_7154);
nand U11584 (N_11584,N_7237,N_6513);
xor U11585 (N_11585,N_5939,N_6640);
nor U11586 (N_11586,N_5525,N_5307);
nand U11587 (N_11587,N_6939,N_5825);
nor U11588 (N_11588,N_7001,N_7321);
or U11589 (N_11589,N_6290,N_6234);
xor U11590 (N_11590,N_5048,N_6930);
or U11591 (N_11591,N_5049,N_7721);
and U11592 (N_11592,N_6097,N_5196);
nor U11593 (N_11593,N_4076,N_7018);
and U11594 (N_11594,N_5612,N_6706);
nor U11595 (N_11595,N_5003,N_4440);
xor U11596 (N_11596,N_5141,N_6349);
nor U11597 (N_11597,N_4014,N_7162);
xnor U11598 (N_11598,N_6409,N_5486);
xor U11599 (N_11599,N_7361,N_7751);
xnor U11600 (N_11600,N_5289,N_4106);
nor U11601 (N_11601,N_7567,N_5443);
or U11602 (N_11602,N_7476,N_6069);
or U11603 (N_11603,N_7608,N_7966);
nand U11604 (N_11604,N_6387,N_4144);
and U11605 (N_11605,N_4861,N_4250);
nor U11606 (N_11606,N_7406,N_7742);
nor U11607 (N_11607,N_4717,N_6217);
nor U11608 (N_11608,N_7120,N_5725);
or U11609 (N_11609,N_6889,N_7931);
xnor U11610 (N_11610,N_4915,N_4981);
and U11611 (N_11611,N_6391,N_6166);
nand U11612 (N_11612,N_7432,N_7691);
nor U11613 (N_11613,N_6098,N_4800);
nor U11614 (N_11614,N_5565,N_5691);
xor U11615 (N_11615,N_7232,N_4519);
or U11616 (N_11616,N_5272,N_6149);
nand U11617 (N_11617,N_5821,N_7369);
or U11618 (N_11618,N_5847,N_6941);
nand U11619 (N_11619,N_4440,N_5672);
xor U11620 (N_11620,N_6775,N_7357);
nand U11621 (N_11621,N_5201,N_6426);
xnor U11622 (N_11622,N_4391,N_5094);
nor U11623 (N_11623,N_5900,N_4392);
xor U11624 (N_11624,N_6343,N_7273);
nor U11625 (N_11625,N_5936,N_4742);
xor U11626 (N_11626,N_6528,N_4359);
nor U11627 (N_11627,N_6717,N_4524);
nor U11628 (N_11628,N_4698,N_7289);
nor U11629 (N_11629,N_4690,N_4785);
nor U11630 (N_11630,N_4745,N_6097);
nor U11631 (N_11631,N_7198,N_4330);
and U11632 (N_11632,N_6927,N_7074);
and U11633 (N_11633,N_4844,N_5458);
and U11634 (N_11634,N_5921,N_5671);
nor U11635 (N_11635,N_4794,N_4258);
nor U11636 (N_11636,N_5881,N_4718);
nor U11637 (N_11637,N_4623,N_4565);
nand U11638 (N_11638,N_5066,N_7218);
xnor U11639 (N_11639,N_4393,N_5534);
nor U11640 (N_11640,N_5083,N_5070);
and U11641 (N_11641,N_4602,N_5372);
and U11642 (N_11642,N_4870,N_4102);
xor U11643 (N_11643,N_5317,N_4526);
or U11644 (N_11644,N_5200,N_5441);
and U11645 (N_11645,N_4409,N_6833);
xnor U11646 (N_11646,N_6820,N_6097);
or U11647 (N_11647,N_7986,N_7008);
and U11648 (N_11648,N_4188,N_6749);
xor U11649 (N_11649,N_5534,N_7963);
nor U11650 (N_11650,N_6800,N_5877);
nand U11651 (N_11651,N_5855,N_6804);
xnor U11652 (N_11652,N_6021,N_5909);
or U11653 (N_11653,N_4916,N_6892);
nor U11654 (N_11654,N_4499,N_7376);
nand U11655 (N_11655,N_7929,N_5999);
and U11656 (N_11656,N_4747,N_6217);
nor U11657 (N_11657,N_5067,N_5082);
and U11658 (N_11658,N_7584,N_6872);
and U11659 (N_11659,N_5844,N_7503);
nand U11660 (N_11660,N_4896,N_7022);
or U11661 (N_11661,N_5827,N_6343);
nand U11662 (N_11662,N_6015,N_7602);
nand U11663 (N_11663,N_4731,N_7132);
or U11664 (N_11664,N_4733,N_7559);
and U11665 (N_11665,N_7268,N_4113);
nor U11666 (N_11666,N_4130,N_7534);
or U11667 (N_11667,N_4864,N_6686);
or U11668 (N_11668,N_6747,N_5856);
xnor U11669 (N_11669,N_7026,N_7638);
xor U11670 (N_11670,N_6488,N_5010);
or U11671 (N_11671,N_7319,N_5579);
nor U11672 (N_11672,N_4547,N_4315);
nor U11673 (N_11673,N_7980,N_5093);
and U11674 (N_11674,N_4533,N_5706);
nand U11675 (N_11675,N_7554,N_5995);
or U11676 (N_11676,N_7709,N_7740);
and U11677 (N_11677,N_5814,N_6733);
nor U11678 (N_11678,N_4962,N_7845);
xnor U11679 (N_11679,N_7121,N_7940);
nand U11680 (N_11680,N_7269,N_4866);
nor U11681 (N_11681,N_5018,N_4653);
or U11682 (N_11682,N_5620,N_5393);
and U11683 (N_11683,N_5753,N_7518);
nand U11684 (N_11684,N_7619,N_5876);
nand U11685 (N_11685,N_5017,N_5658);
and U11686 (N_11686,N_7526,N_4402);
nor U11687 (N_11687,N_6144,N_4812);
or U11688 (N_11688,N_4181,N_7032);
and U11689 (N_11689,N_5272,N_5847);
nand U11690 (N_11690,N_7825,N_4595);
xnor U11691 (N_11691,N_6155,N_5846);
or U11692 (N_11692,N_5863,N_5077);
xor U11693 (N_11693,N_4370,N_5744);
nand U11694 (N_11694,N_6503,N_6539);
nor U11695 (N_11695,N_5700,N_6742);
or U11696 (N_11696,N_4772,N_7982);
xor U11697 (N_11697,N_5990,N_5330);
nand U11698 (N_11698,N_5400,N_6944);
and U11699 (N_11699,N_4458,N_7541);
xnor U11700 (N_11700,N_4812,N_6031);
or U11701 (N_11701,N_7429,N_6915);
and U11702 (N_11702,N_7278,N_7257);
nand U11703 (N_11703,N_6670,N_4531);
xnor U11704 (N_11704,N_6669,N_5877);
or U11705 (N_11705,N_6086,N_6310);
and U11706 (N_11706,N_4176,N_6383);
and U11707 (N_11707,N_7347,N_4295);
nor U11708 (N_11708,N_7335,N_6929);
and U11709 (N_11709,N_5660,N_7203);
xor U11710 (N_11710,N_5580,N_5958);
nand U11711 (N_11711,N_5651,N_6275);
or U11712 (N_11712,N_6516,N_5239);
or U11713 (N_11713,N_7774,N_4938);
xnor U11714 (N_11714,N_5898,N_4564);
and U11715 (N_11715,N_4564,N_4837);
nand U11716 (N_11716,N_4328,N_5432);
nor U11717 (N_11717,N_4296,N_7984);
nor U11718 (N_11718,N_4921,N_6530);
or U11719 (N_11719,N_5548,N_6963);
nor U11720 (N_11720,N_6911,N_7784);
nand U11721 (N_11721,N_6955,N_7474);
xnor U11722 (N_11722,N_7524,N_7733);
nor U11723 (N_11723,N_6638,N_5722);
and U11724 (N_11724,N_6374,N_7173);
xor U11725 (N_11725,N_4584,N_7296);
nand U11726 (N_11726,N_6274,N_5635);
nand U11727 (N_11727,N_6652,N_4324);
nor U11728 (N_11728,N_6125,N_7249);
nor U11729 (N_11729,N_7278,N_4300);
nand U11730 (N_11730,N_7682,N_5176);
xor U11731 (N_11731,N_6816,N_4331);
nor U11732 (N_11732,N_6445,N_7291);
xor U11733 (N_11733,N_4566,N_7633);
xnor U11734 (N_11734,N_6739,N_6134);
nand U11735 (N_11735,N_4456,N_6989);
xnor U11736 (N_11736,N_4037,N_6782);
or U11737 (N_11737,N_5714,N_7889);
and U11738 (N_11738,N_4085,N_5540);
nand U11739 (N_11739,N_6375,N_6905);
or U11740 (N_11740,N_5446,N_5232);
nand U11741 (N_11741,N_7982,N_7249);
xnor U11742 (N_11742,N_7897,N_7968);
or U11743 (N_11743,N_4447,N_6224);
xor U11744 (N_11744,N_4872,N_4638);
or U11745 (N_11745,N_5179,N_6775);
nand U11746 (N_11746,N_4985,N_7627);
nor U11747 (N_11747,N_5231,N_7689);
xnor U11748 (N_11748,N_5799,N_4827);
nor U11749 (N_11749,N_4245,N_7377);
nand U11750 (N_11750,N_6652,N_6310);
and U11751 (N_11751,N_7348,N_5738);
or U11752 (N_11752,N_7478,N_5386);
or U11753 (N_11753,N_7477,N_5731);
and U11754 (N_11754,N_7793,N_4954);
nand U11755 (N_11755,N_6054,N_5822);
nand U11756 (N_11756,N_7433,N_6930);
nor U11757 (N_11757,N_6083,N_5515);
nor U11758 (N_11758,N_5004,N_5134);
or U11759 (N_11759,N_6960,N_6225);
xor U11760 (N_11760,N_7534,N_7416);
nor U11761 (N_11761,N_6065,N_7223);
xor U11762 (N_11762,N_7938,N_7210);
or U11763 (N_11763,N_5643,N_7740);
xnor U11764 (N_11764,N_5058,N_4616);
xnor U11765 (N_11765,N_6427,N_6599);
nand U11766 (N_11766,N_5400,N_6913);
nor U11767 (N_11767,N_6473,N_7422);
and U11768 (N_11768,N_7534,N_5019);
and U11769 (N_11769,N_5994,N_6114);
nor U11770 (N_11770,N_4626,N_4109);
nand U11771 (N_11771,N_7166,N_7348);
or U11772 (N_11772,N_5987,N_6167);
and U11773 (N_11773,N_6849,N_5899);
nor U11774 (N_11774,N_7125,N_4268);
and U11775 (N_11775,N_5552,N_4299);
nand U11776 (N_11776,N_6015,N_4882);
nor U11777 (N_11777,N_4769,N_6249);
nand U11778 (N_11778,N_5899,N_6956);
nor U11779 (N_11779,N_7278,N_4639);
nand U11780 (N_11780,N_6097,N_7405);
xnor U11781 (N_11781,N_6268,N_7730);
nor U11782 (N_11782,N_6063,N_6393);
or U11783 (N_11783,N_5488,N_7397);
xnor U11784 (N_11784,N_6808,N_5354);
and U11785 (N_11785,N_7347,N_7130);
xnor U11786 (N_11786,N_7402,N_5852);
xor U11787 (N_11787,N_7444,N_5601);
and U11788 (N_11788,N_7633,N_5829);
and U11789 (N_11789,N_5623,N_7663);
or U11790 (N_11790,N_6984,N_5152);
nor U11791 (N_11791,N_6476,N_5050);
nand U11792 (N_11792,N_5686,N_5253);
and U11793 (N_11793,N_5963,N_4139);
xor U11794 (N_11794,N_6537,N_5729);
nor U11795 (N_11795,N_5926,N_7653);
and U11796 (N_11796,N_7463,N_7802);
and U11797 (N_11797,N_4788,N_7497);
or U11798 (N_11798,N_6422,N_7263);
and U11799 (N_11799,N_6360,N_7058);
or U11800 (N_11800,N_7779,N_4822);
or U11801 (N_11801,N_7505,N_5606);
and U11802 (N_11802,N_7517,N_5792);
nor U11803 (N_11803,N_4700,N_6689);
and U11804 (N_11804,N_4578,N_4627);
and U11805 (N_11805,N_7185,N_5046);
xnor U11806 (N_11806,N_4845,N_7285);
nor U11807 (N_11807,N_7246,N_5913);
nor U11808 (N_11808,N_7086,N_5804);
and U11809 (N_11809,N_4492,N_7918);
and U11810 (N_11810,N_4146,N_7269);
nor U11811 (N_11811,N_5525,N_5083);
or U11812 (N_11812,N_7769,N_6637);
and U11813 (N_11813,N_4265,N_4462);
nand U11814 (N_11814,N_5107,N_6466);
xnor U11815 (N_11815,N_6662,N_6857);
and U11816 (N_11816,N_4516,N_5311);
xnor U11817 (N_11817,N_7956,N_4467);
or U11818 (N_11818,N_5944,N_6984);
nor U11819 (N_11819,N_5185,N_6595);
nand U11820 (N_11820,N_7979,N_7098);
or U11821 (N_11821,N_4532,N_5787);
and U11822 (N_11822,N_4654,N_7105);
or U11823 (N_11823,N_5749,N_5069);
or U11824 (N_11824,N_4291,N_5303);
nor U11825 (N_11825,N_4330,N_7074);
and U11826 (N_11826,N_4201,N_7015);
nor U11827 (N_11827,N_6750,N_7321);
or U11828 (N_11828,N_7436,N_4826);
or U11829 (N_11829,N_7427,N_4098);
nand U11830 (N_11830,N_7542,N_7807);
and U11831 (N_11831,N_4313,N_5958);
or U11832 (N_11832,N_4729,N_5575);
or U11833 (N_11833,N_5708,N_5254);
xor U11834 (N_11834,N_5767,N_6422);
nand U11835 (N_11835,N_5565,N_7613);
or U11836 (N_11836,N_4242,N_6338);
xor U11837 (N_11837,N_6865,N_5493);
xor U11838 (N_11838,N_7300,N_6755);
nor U11839 (N_11839,N_4377,N_5619);
xnor U11840 (N_11840,N_6561,N_6632);
nor U11841 (N_11841,N_6486,N_4635);
or U11842 (N_11842,N_6763,N_4243);
or U11843 (N_11843,N_5534,N_6782);
xor U11844 (N_11844,N_7686,N_6572);
nand U11845 (N_11845,N_7783,N_4694);
and U11846 (N_11846,N_4042,N_5242);
xnor U11847 (N_11847,N_4774,N_7225);
or U11848 (N_11848,N_6826,N_7987);
nand U11849 (N_11849,N_4897,N_7594);
nor U11850 (N_11850,N_6683,N_7375);
xnor U11851 (N_11851,N_7080,N_6560);
nor U11852 (N_11852,N_7719,N_5778);
or U11853 (N_11853,N_5807,N_7559);
and U11854 (N_11854,N_6067,N_7658);
xor U11855 (N_11855,N_4187,N_7734);
and U11856 (N_11856,N_6733,N_5959);
or U11857 (N_11857,N_7477,N_4929);
nor U11858 (N_11858,N_4579,N_5185);
or U11859 (N_11859,N_6373,N_6278);
xor U11860 (N_11860,N_5024,N_4117);
or U11861 (N_11861,N_4686,N_6543);
nand U11862 (N_11862,N_4744,N_6998);
nor U11863 (N_11863,N_5039,N_5857);
and U11864 (N_11864,N_5028,N_5819);
xor U11865 (N_11865,N_5729,N_7619);
nor U11866 (N_11866,N_6765,N_4594);
or U11867 (N_11867,N_5438,N_4931);
and U11868 (N_11868,N_5045,N_6535);
nor U11869 (N_11869,N_5430,N_5699);
or U11870 (N_11870,N_5773,N_5786);
nand U11871 (N_11871,N_5306,N_4659);
nor U11872 (N_11872,N_5555,N_7377);
nor U11873 (N_11873,N_5427,N_6930);
xnor U11874 (N_11874,N_5235,N_4939);
or U11875 (N_11875,N_6119,N_4874);
or U11876 (N_11876,N_5754,N_4322);
nor U11877 (N_11877,N_7495,N_7915);
and U11878 (N_11878,N_4507,N_7314);
xor U11879 (N_11879,N_5944,N_4043);
nand U11880 (N_11880,N_7721,N_6972);
nand U11881 (N_11881,N_7233,N_7067);
and U11882 (N_11882,N_4361,N_4828);
nor U11883 (N_11883,N_6161,N_5283);
nor U11884 (N_11884,N_4880,N_6838);
nand U11885 (N_11885,N_7305,N_7974);
nor U11886 (N_11886,N_4258,N_7666);
xor U11887 (N_11887,N_7311,N_4389);
and U11888 (N_11888,N_4979,N_6401);
and U11889 (N_11889,N_4388,N_5901);
or U11890 (N_11890,N_6543,N_6695);
nand U11891 (N_11891,N_7206,N_6540);
nor U11892 (N_11892,N_5263,N_6860);
nor U11893 (N_11893,N_7121,N_5480);
xnor U11894 (N_11894,N_4826,N_5994);
and U11895 (N_11895,N_7494,N_4934);
nor U11896 (N_11896,N_6208,N_6754);
nand U11897 (N_11897,N_4528,N_7938);
nor U11898 (N_11898,N_7982,N_6442);
xor U11899 (N_11899,N_5274,N_4719);
and U11900 (N_11900,N_6293,N_7521);
xnor U11901 (N_11901,N_7945,N_6511);
and U11902 (N_11902,N_7590,N_4177);
and U11903 (N_11903,N_5787,N_6782);
and U11904 (N_11904,N_6544,N_6951);
nor U11905 (N_11905,N_7852,N_5045);
xor U11906 (N_11906,N_5211,N_6160);
nor U11907 (N_11907,N_7889,N_6024);
and U11908 (N_11908,N_5974,N_7497);
and U11909 (N_11909,N_5280,N_6949);
and U11910 (N_11910,N_7314,N_5512);
and U11911 (N_11911,N_4202,N_4344);
nand U11912 (N_11912,N_7231,N_5764);
or U11913 (N_11913,N_7312,N_6644);
nor U11914 (N_11914,N_4719,N_5920);
xor U11915 (N_11915,N_4973,N_4344);
xnor U11916 (N_11916,N_4137,N_6225);
xnor U11917 (N_11917,N_6158,N_4380);
nor U11918 (N_11918,N_7190,N_6041);
xnor U11919 (N_11919,N_7561,N_7416);
nor U11920 (N_11920,N_7455,N_5491);
nor U11921 (N_11921,N_7240,N_7876);
nor U11922 (N_11922,N_5647,N_4908);
and U11923 (N_11923,N_5398,N_7882);
xor U11924 (N_11924,N_4138,N_4299);
nor U11925 (N_11925,N_5312,N_5921);
or U11926 (N_11926,N_7789,N_4977);
nand U11927 (N_11927,N_6589,N_6699);
xor U11928 (N_11928,N_7943,N_6446);
nor U11929 (N_11929,N_6567,N_5891);
xor U11930 (N_11930,N_5962,N_4489);
nand U11931 (N_11931,N_7422,N_7239);
nand U11932 (N_11932,N_5119,N_7837);
and U11933 (N_11933,N_4114,N_4183);
nand U11934 (N_11934,N_5012,N_5647);
xor U11935 (N_11935,N_7943,N_5284);
and U11936 (N_11936,N_6295,N_5932);
and U11937 (N_11937,N_6287,N_6684);
nand U11938 (N_11938,N_4768,N_7072);
nor U11939 (N_11939,N_7619,N_5117);
or U11940 (N_11940,N_6428,N_7825);
xnor U11941 (N_11941,N_4376,N_5659);
xor U11942 (N_11942,N_5760,N_6858);
nand U11943 (N_11943,N_6439,N_6072);
nand U11944 (N_11944,N_5324,N_6821);
xnor U11945 (N_11945,N_6518,N_5626);
and U11946 (N_11946,N_7617,N_7857);
or U11947 (N_11947,N_6009,N_4230);
nand U11948 (N_11948,N_7638,N_6815);
or U11949 (N_11949,N_4654,N_5044);
or U11950 (N_11950,N_7805,N_6095);
xnor U11951 (N_11951,N_5375,N_4418);
nand U11952 (N_11952,N_6350,N_4651);
xor U11953 (N_11953,N_5829,N_7716);
nand U11954 (N_11954,N_6813,N_7156);
nor U11955 (N_11955,N_4741,N_4124);
nand U11956 (N_11956,N_5714,N_6946);
or U11957 (N_11957,N_7306,N_6868);
or U11958 (N_11958,N_4184,N_6938);
and U11959 (N_11959,N_4313,N_4835);
and U11960 (N_11960,N_4908,N_7594);
nand U11961 (N_11961,N_6924,N_7981);
xnor U11962 (N_11962,N_5304,N_7304);
or U11963 (N_11963,N_5814,N_6419);
and U11964 (N_11964,N_5493,N_5853);
nand U11965 (N_11965,N_7998,N_7953);
xor U11966 (N_11966,N_4066,N_7501);
and U11967 (N_11967,N_4550,N_4440);
xnor U11968 (N_11968,N_6870,N_7761);
and U11969 (N_11969,N_4776,N_7188);
and U11970 (N_11970,N_7556,N_7011);
nor U11971 (N_11971,N_7620,N_5506);
nand U11972 (N_11972,N_7578,N_6591);
or U11973 (N_11973,N_5349,N_4136);
nor U11974 (N_11974,N_4056,N_6867);
or U11975 (N_11975,N_7613,N_4990);
and U11976 (N_11976,N_7518,N_7960);
xnor U11977 (N_11977,N_4734,N_5528);
or U11978 (N_11978,N_5334,N_5915);
or U11979 (N_11979,N_4144,N_5958);
and U11980 (N_11980,N_5944,N_7927);
or U11981 (N_11981,N_5589,N_7101);
nand U11982 (N_11982,N_7644,N_4176);
xnor U11983 (N_11983,N_4805,N_5258);
or U11984 (N_11984,N_7475,N_5387);
and U11985 (N_11985,N_4358,N_5876);
xor U11986 (N_11986,N_6974,N_5388);
or U11987 (N_11987,N_4332,N_4446);
nand U11988 (N_11988,N_5190,N_7614);
xor U11989 (N_11989,N_4115,N_6337);
and U11990 (N_11990,N_6913,N_5505);
and U11991 (N_11991,N_5096,N_7311);
nand U11992 (N_11992,N_5057,N_5337);
xnor U11993 (N_11993,N_5983,N_7437);
and U11994 (N_11994,N_5760,N_6294);
nor U11995 (N_11995,N_6397,N_4520);
xnor U11996 (N_11996,N_6949,N_5822);
nand U11997 (N_11997,N_5810,N_5716);
nor U11998 (N_11998,N_4239,N_7333);
nand U11999 (N_11999,N_4986,N_7655);
and U12000 (N_12000,N_10399,N_10851);
nor U12001 (N_12001,N_10903,N_10460);
xor U12002 (N_12002,N_9362,N_10975);
and U12003 (N_12003,N_10433,N_8510);
nand U12004 (N_12004,N_11929,N_8536);
and U12005 (N_12005,N_10067,N_11965);
or U12006 (N_12006,N_8334,N_10240);
nor U12007 (N_12007,N_9385,N_10722);
or U12008 (N_12008,N_8314,N_10747);
or U12009 (N_12009,N_10704,N_8262);
nor U12010 (N_12010,N_11981,N_11573);
nand U12011 (N_12011,N_10802,N_11888);
nand U12012 (N_12012,N_8843,N_9046);
nand U12013 (N_12013,N_8454,N_10138);
nand U12014 (N_12014,N_8156,N_9326);
nand U12015 (N_12015,N_10768,N_9800);
and U12016 (N_12016,N_9298,N_10529);
nand U12017 (N_12017,N_9043,N_11960);
nor U12018 (N_12018,N_11153,N_9719);
nor U12019 (N_12019,N_8374,N_10242);
nor U12020 (N_12020,N_11286,N_10264);
or U12021 (N_12021,N_11602,N_8324);
nor U12022 (N_12022,N_9579,N_8507);
nor U12023 (N_12023,N_11677,N_9999);
or U12024 (N_12024,N_11978,N_11575);
nor U12025 (N_12025,N_8500,N_9008);
xnor U12026 (N_12026,N_11473,N_11064);
or U12027 (N_12027,N_9885,N_10088);
and U12028 (N_12028,N_8357,N_9509);
xor U12029 (N_12029,N_8444,N_8355);
nand U12030 (N_12030,N_10835,N_11519);
and U12031 (N_12031,N_10760,N_10686);
and U12032 (N_12032,N_8197,N_8950);
xor U12033 (N_12033,N_9347,N_9744);
and U12034 (N_12034,N_11736,N_10350);
nand U12035 (N_12035,N_8328,N_8201);
or U12036 (N_12036,N_10480,N_9214);
xnor U12037 (N_12037,N_11379,N_11729);
nand U12038 (N_12038,N_8435,N_10390);
or U12039 (N_12039,N_9545,N_11662);
or U12040 (N_12040,N_8868,N_11100);
nand U12041 (N_12041,N_10905,N_10696);
nand U12042 (N_12042,N_10886,N_9196);
nor U12043 (N_12043,N_11655,N_11209);
and U12044 (N_12044,N_9118,N_11122);
and U12045 (N_12045,N_9612,N_9276);
nand U12046 (N_12046,N_10432,N_11325);
nand U12047 (N_12047,N_8647,N_8187);
nand U12048 (N_12048,N_8354,N_9714);
xnor U12049 (N_12049,N_10169,N_10007);
and U12050 (N_12050,N_9556,N_9845);
nand U12051 (N_12051,N_9132,N_11016);
nand U12052 (N_12052,N_8714,N_8504);
nor U12053 (N_12053,N_10537,N_11382);
xnor U12054 (N_12054,N_9318,N_11351);
xnor U12055 (N_12055,N_8017,N_9166);
or U12056 (N_12056,N_8805,N_11605);
nand U12057 (N_12057,N_8997,N_10613);
and U12058 (N_12058,N_9301,N_9954);
nor U12059 (N_12059,N_10646,N_11893);
or U12060 (N_12060,N_10134,N_10667);
or U12061 (N_12061,N_11048,N_9552);
and U12062 (N_12062,N_11322,N_10158);
nor U12063 (N_12063,N_8756,N_9128);
nand U12064 (N_12064,N_10687,N_11420);
and U12065 (N_12065,N_10873,N_9437);
or U12066 (N_12066,N_8616,N_8390);
nor U12067 (N_12067,N_10834,N_10622);
or U12068 (N_12068,N_8703,N_9784);
and U12069 (N_12069,N_8564,N_10643);
nand U12070 (N_12070,N_10414,N_10875);
nand U12071 (N_12071,N_9648,N_11020);
xnor U12072 (N_12072,N_9478,N_10235);
xor U12073 (N_12073,N_8109,N_9844);
xnor U12074 (N_12074,N_8934,N_11335);
nand U12075 (N_12075,N_10018,N_11009);
nor U12076 (N_12076,N_10694,N_11486);
or U12077 (N_12077,N_11877,N_8698);
xor U12078 (N_12078,N_10413,N_8654);
or U12079 (N_12079,N_9087,N_10815);
nor U12080 (N_12080,N_11703,N_11748);
nand U12081 (N_12081,N_10522,N_8863);
nand U12082 (N_12082,N_11727,N_11529);
or U12083 (N_12083,N_8169,N_8525);
nand U12084 (N_12084,N_8214,N_11433);
nand U12085 (N_12085,N_10459,N_9490);
nand U12086 (N_12086,N_9254,N_10231);
and U12087 (N_12087,N_9014,N_10910);
nand U12088 (N_12088,N_10915,N_10510);
and U12089 (N_12089,N_10317,N_8605);
and U12090 (N_12090,N_8825,N_8019);
and U12091 (N_12091,N_9164,N_8486);
and U12092 (N_12092,N_9642,N_8148);
xor U12093 (N_12093,N_10441,N_11266);
nand U12094 (N_12094,N_8153,N_10600);
and U12095 (N_12095,N_11264,N_11517);
and U12096 (N_12096,N_10650,N_9373);
nor U12097 (N_12097,N_8346,N_9617);
nand U12098 (N_12098,N_11394,N_10945);
or U12099 (N_12099,N_9093,N_10715);
nor U12100 (N_12100,N_9910,N_10526);
nand U12101 (N_12101,N_10409,N_8671);
and U12102 (N_12102,N_10482,N_10523);
nor U12103 (N_12103,N_10934,N_8502);
and U12104 (N_12104,N_9964,N_11767);
nand U12105 (N_12105,N_8277,N_8343);
nor U12106 (N_12106,N_9472,N_10926);
or U12107 (N_12107,N_8617,N_9782);
xnor U12108 (N_12108,N_8592,N_10228);
or U12109 (N_12109,N_10772,N_11706);
and U12110 (N_12110,N_11504,N_10415);
nor U12111 (N_12111,N_9045,N_9703);
xor U12112 (N_12112,N_10788,N_11721);
nor U12113 (N_12113,N_10180,N_11759);
and U12114 (N_12114,N_8327,N_9170);
nand U12115 (N_12115,N_11953,N_8437);
nor U12116 (N_12116,N_11024,N_8269);
nand U12117 (N_12117,N_11755,N_11537);
nand U12118 (N_12118,N_10006,N_9958);
xnor U12119 (N_12119,N_8035,N_8131);
and U12120 (N_12120,N_11352,N_10351);
nand U12121 (N_12121,N_9213,N_11171);
xor U12122 (N_12122,N_11902,N_10097);
nor U12123 (N_12123,N_10499,N_9313);
and U12124 (N_12124,N_11829,N_8348);
nor U12125 (N_12125,N_11788,N_11045);
or U12126 (N_12126,N_10695,N_11523);
nand U12127 (N_12127,N_11125,N_8782);
xnor U12128 (N_12128,N_10019,N_10394);
nand U12129 (N_12129,N_9914,N_10462);
xor U12130 (N_12130,N_8160,N_10367);
or U12131 (N_12131,N_10353,N_11040);
nand U12132 (N_12132,N_9309,N_9698);
nor U12133 (N_12133,N_9391,N_10592);
xor U12134 (N_12134,N_9572,N_8462);
xor U12135 (N_12135,N_9827,N_10133);
nor U12136 (N_12136,N_8886,N_10178);
xor U12137 (N_12137,N_8353,N_9027);
nand U12138 (N_12138,N_9908,N_9236);
nand U12139 (N_12139,N_11556,N_10001);
and U12140 (N_12140,N_11363,N_9248);
and U12141 (N_12141,N_8526,N_8810);
xnor U12142 (N_12142,N_10784,N_8340);
or U12143 (N_12143,N_8993,N_11050);
or U12144 (N_12144,N_9832,N_11852);
and U12145 (N_12145,N_8113,N_11320);
nor U12146 (N_12146,N_8759,N_9665);
nor U12147 (N_12147,N_10412,N_10253);
nand U12148 (N_12148,N_8761,N_10201);
or U12149 (N_12149,N_8967,N_10064);
xnor U12150 (N_12150,N_10058,N_11492);
and U12151 (N_12151,N_9032,N_11372);
or U12152 (N_12152,N_10050,N_8243);
xor U12153 (N_12153,N_10683,N_8827);
xnor U12154 (N_12154,N_11425,N_9191);
xnor U12155 (N_12155,N_11553,N_8920);
nand U12156 (N_12156,N_9283,N_11001);
nor U12157 (N_12157,N_9407,N_11114);
or U12158 (N_12158,N_9553,N_8938);
or U12159 (N_12159,N_9595,N_11306);
nor U12160 (N_12160,N_11479,N_11664);
nand U12161 (N_12161,N_11235,N_10444);
or U12162 (N_12162,N_9888,N_8190);
or U12163 (N_12163,N_8724,N_11448);
xor U12164 (N_12164,N_9245,N_10030);
xor U12165 (N_12165,N_11107,N_11327);
and U12166 (N_12166,N_8232,N_11735);
nand U12167 (N_12167,N_11871,N_10308);
nand U12168 (N_12168,N_11560,N_9621);
nor U12169 (N_12169,N_8414,N_9742);
nor U12170 (N_12170,N_11133,N_11915);
and U12171 (N_12171,N_8445,N_9447);
and U12172 (N_12172,N_10531,N_9038);
nor U12173 (N_12173,N_9105,N_8428);
xnor U12174 (N_12174,N_10419,N_10617);
nor U12175 (N_12175,N_10916,N_10188);
nor U12176 (N_12176,N_8817,N_10557);
or U12177 (N_12177,N_10345,N_8049);
nor U12178 (N_12178,N_11475,N_11731);
and U12179 (N_12179,N_10485,N_11079);
nor U12180 (N_12180,N_10372,N_9945);
nand U12181 (N_12181,N_8591,N_11857);
nand U12182 (N_12182,N_9411,N_8961);
or U12183 (N_12183,N_11521,N_10824);
nor U12184 (N_12184,N_8432,N_8167);
or U12185 (N_12185,N_8128,N_11797);
or U12186 (N_12186,N_10654,N_9293);
nor U12187 (N_12187,N_9146,N_10359);
nor U12188 (N_12188,N_10269,N_10319);
xnor U12189 (N_12189,N_8222,N_11751);
and U12190 (N_12190,N_10734,N_9836);
nor U12191 (N_12191,N_10864,N_9551);
xor U12192 (N_12192,N_10774,N_8323);
xnor U12193 (N_12193,N_9815,N_9876);
nor U12194 (N_12194,N_9348,N_9530);
nand U12195 (N_12195,N_9823,N_10422);
nand U12196 (N_12196,N_11691,N_11318);
nand U12197 (N_12197,N_8238,N_11455);
nand U12198 (N_12198,N_9991,N_11513);
nand U12199 (N_12199,N_8539,N_9272);
xor U12200 (N_12200,N_8272,N_11661);
and U12201 (N_12201,N_10487,N_10278);
nand U12202 (N_12202,N_11301,N_10465);
and U12203 (N_12203,N_10146,N_8072);
nor U12204 (N_12204,N_8776,N_8203);
nor U12205 (N_12205,N_9630,N_9417);
xnor U12206 (N_12206,N_11506,N_10985);
nor U12207 (N_12207,N_8608,N_11069);
nand U12208 (N_12208,N_8907,N_10380);
and U12209 (N_12209,N_10493,N_9380);
and U12210 (N_12210,N_11577,N_8080);
or U12211 (N_12211,N_11968,N_10120);
or U12212 (N_12212,N_10451,N_10026);
nand U12213 (N_12213,N_10448,N_8597);
nand U12214 (N_12214,N_9358,N_8003);
nand U12215 (N_12215,N_11890,N_11883);
and U12216 (N_12216,N_8789,N_10124);
nand U12217 (N_12217,N_9299,N_10859);
and U12218 (N_12218,N_9840,N_9103);
nor U12219 (N_12219,N_11592,N_11511);
nand U12220 (N_12220,N_10940,N_8958);
xor U12221 (N_12221,N_8060,N_9095);
and U12222 (N_12222,N_11637,N_9134);
and U12223 (N_12223,N_11572,N_9135);
and U12224 (N_12224,N_10321,N_10156);
nor U12225 (N_12225,N_8531,N_9178);
or U12226 (N_12226,N_11456,N_8086);
xnor U12227 (N_12227,N_9073,N_11060);
or U12228 (N_12228,N_11000,N_10434);
and U12229 (N_12229,N_9715,N_8151);
and U12230 (N_12230,N_10376,N_10805);
or U12231 (N_12231,N_8368,N_10628);
and U12232 (N_12232,N_9549,N_11167);
xnor U12233 (N_12233,N_10065,N_11168);
or U12234 (N_12234,N_10404,N_8016);
or U12235 (N_12235,N_8372,N_9382);
xnor U12236 (N_12236,N_8455,N_8794);
xnor U12237 (N_12237,N_8708,N_9446);
and U12238 (N_12238,N_10241,N_8037);
nand U12239 (N_12239,N_10852,N_8155);
xnor U12240 (N_12240,N_9930,N_11732);
and U12241 (N_12241,N_9247,N_10500);
or U12242 (N_12242,N_10816,N_10872);
and U12243 (N_12243,N_11381,N_9017);
nand U12244 (N_12244,N_9540,N_10458);
and U12245 (N_12245,N_8560,N_10958);
xor U12246 (N_12246,N_8484,N_8893);
and U12247 (N_12247,N_11940,N_8226);
xor U12248 (N_12248,N_8797,N_9675);
xnor U12249 (N_12249,N_9928,N_8194);
or U12250 (N_12250,N_8031,N_10825);
and U12251 (N_12251,N_8145,N_10103);
or U12252 (N_12252,N_10792,N_8304);
or U12253 (N_12253,N_8066,N_11354);
nor U12254 (N_12254,N_8528,N_10927);
and U12255 (N_12255,N_9237,N_10957);
and U12256 (N_12256,N_10749,N_11653);
xor U12257 (N_12257,N_9406,N_11061);
nor U12258 (N_12258,N_8733,N_10861);
nand U12259 (N_12259,N_8436,N_11065);
nand U12260 (N_12260,N_9314,N_8103);
or U12261 (N_12261,N_10011,N_8685);
xor U12262 (N_12262,N_11058,N_10648);
nand U12263 (N_12263,N_10143,N_10837);
nand U12264 (N_12264,N_8076,N_9106);
xor U12265 (N_12265,N_10371,N_10579);
and U12266 (N_12266,N_8318,N_10756);
xor U12267 (N_12267,N_9136,N_9275);
xor U12268 (N_12268,N_10899,N_10325);
or U12269 (N_12269,N_8609,N_11846);
or U12270 (N_12270,N_10265,N_10469);
xor U12271 (N_12271,N_8929,N_8281);
nand U12272 (N_12272,N_11823,N_9951);
nor U12273 (N_12273,N_10283,N_9671);
nand U12274 (N_12274,N_8866,N_10416);
or U12275 (N_12275,N_8063,N_9889);
nor U12276 (N_12276,N_10868,N_11076);
nor U12277 (N_12277,N_9709,N_11428);
and U12278 (N_12278,N_9229,N_9280);
nor U12279 (N_12279,N_10014,N_11142);
nor U12280 (N_12280,N_11358,N_9837);
nor U12281 (N_12281,N_8196,N_8569);
and U12282 (N_12282,N_8095,N_9850);
nor U12283 (N_12283,N_9831,N_9527);
and U12284 (N_12284,N_10437,N_9938);
nand U12285 (N_12285,N_11780,N_10970);
nand U12286 (N_12286,N_8449,N_9761);
and U12287 (N_12287,N_8315,N_11388);
nor U12288 (N_12288,N_8771,N_8847);
nand U12289 (N_12289,N_8468,N_11184);
xnor U12290 (N_12290,N_8081,N_8082);
or U12291 (N_12291,N_10125,N_11574);
and U12292 (N_12292,N_11265,N_10347);
xor U12293 (N_12293,N_11734,N_11546);
nor U12294 (N_12294,N_10769,N_10584);
or U12295 (N_12295,N_8573,N_9871);
nor U12296 (N_12296,N_10086,N_11545);
and U12297 (N_12297,N_9636,N_10327);
nand U12298 (N_12298,N_8820,N_9200);
nor U12299 (N_12299,N_10087,N_8188);
and U12300 (N_12300,N_11404,N_9581);
nand U12301 (N_12301,N_9244,N_10807);
and U12302 (N_12302,N_8699,N_9993);
nand U12303 (N_12303,N_8135,N_9585);
or U12304 (N_12304,N_9379,N_11740);
nand U12305 (N_12305,N_10583,N_11785);
nand U12306 (N_12306,N_11768,N_9408);
nand U12307 (N_12307,N_11175,N_10332);
and U12308 (N_12308,N_9000,N_8750);
nand U12309 (N_12309,N_10941,N_9234);
xor U12310 (N_12310,N_9687,N_11242);
and U12311 (N_12311,N_11134,N_8041);
and U12312 (N_12312,N_10753,N_9335);
nor U12313 (N_12313,N_8532,N_9352);
and U12314 (N_12314,N_9059,N_11961);
xnor U12315 (N_12315,N_8288,N_10168);
and U12316 (N_12316,N_10301,N_11126);
nor U12317 (N_12317,N_11702,N_10152);
nand U12318 (N_12318,N_9656,N_10547);
nor U12319 (N_12319,N_8168,N_8307);
nand U12320 (N_12320,N_10215,N_8199);
and U12321 (N_12321,N_10079,N_10318);
nand U12322 (N_12322,N_9153,N_9216);
or U12323 (N_12323,N_11928,N_10259);
nor U12324 (N_12324,N_10664,N_11904);
and U12325 (N_12325,N_10731,N_9026);
and U12326 (N_12326,N_9094,N_10291);
xor U12327 (N_12327,N_9481,N_8807);
nand U12328 (N_12328,N_8915,N_9693);
and U12329 (N_12329,N_8356,N_10644);
and U12330 (N_12330,N_9662,N_11195);
xnor U12331 (N_12331,N_10068,N_8464);
nand U12332 (N_12332,N_11089,N_9926);
nand U12333 (N_12333,N_11062,N_8630);
nand U12334 (N_12334,N_9565,N_8011);
and U12335 (N_12335,N_9536,N_9329);
nor U12336 (N_12336,N_11336,N_8032);
and U12337 (N_12337,N_9251,N_11399);
xor U12338 (N_12338,N_11021,N_11665);
and U12339 (N_12339,N_10368,N_9075);
xor U12340 (N_12340,N_11743,N_8611);
nand U12341 (N_12341,N_11027,N_10515);
nor U12342 (N_12342,N_11724,N_10032);
xor U12343 (N_12343,N_10727,N_11868);
nor U12344 (N_12344,N_10906,N_10285);
nand U12345 (N_12345,N_9913,N_11495);
nor U12346 (N_12346,N_10360,N_11243);
and U12347 (N_12347,N_9864,N_9249);
nand U12348 (N_12348,N_8955,N_8633);
nand U12349 (N_12349,N_8317,N_9496);
nor U12350 (N_12350,N_8692,N_10219);
or U12351 (N_12351,N_8702,N_9874);
nand U12352 (N_12352,N_9820,N_10542);
nor U12353 (N_12353,N_11843,N_10966);
nand U12354 (N_12354,N_8251,N_8036);
or U12355 (N_12355,N_10021,N_8244);
and U12356 (N_12356,N_9271,N_9351);
or U12357 (N_12357,N_8061,N_9525);
and U12358 (N_12358,N_11538,N_8954);
or U12359 (N_12359,N_10186,N_11332);
and U12360 (N_12360,N_11796,N_10268);
and U12361 (N_12361,N_9635,N_9706);
or U12362 (N_12362,N_8142,N_10436);
and U12363 (N_12363,N_11876,N_11183);
and U12364 (N_12364,N_8895,N_10733);
and U12365 (N_12365,N_10445,N_8697);
nand U12366 (N_12366,N_9848,N_10503);
or U12367 (N_12367,N_11112,N_8044);
xor U12368 (N_12368,N_10532,N_8496);
nor U12369 (N_12369,N_10209,N_8133);
or U12370 (N_12370,N_9450,N_9020);
or U12371 (N_12371,N_11109,N_11201);
xnor U12372 (N_12372,N_8575,N_10912);
and U12373 (N_12373,N_9495,N_9315);
and U12374 (N_12374,N_9033,N_10038);
nand U12375 (N_12375,N_10297,N_8839);
and U12376 (N_12376,N_10363,N_8914);
xor U12377 (N_12377,N_9976,N_8069);
or U12378 (N_12378,N_8921,N_10652);
nand U12379 (N_12379,N_9805,N_8010);
and U12380 (N_12380,N_10013,N_8758);
xnor U12381 (N_12381,N_9949,N_9183);
or U12382 (N_12382,N_9101,N_10177);
nor U12383 (N_12383,N_11726,N_11221);
xnor U12384 (N_12384,N_10044,N_11685);
nor U12385 (N_12385,N_11579,N_9988);
or U12386 (N_12386,N_10573,N_8034);
or U12387 (N_12387,N_8970,N_11692);
nor U12388 (N_12388,N_8184,N_8619);
or U12389 (N_12389,N_9503,N_8542);
or U12390 (N_12390,N_8058,N_11808);
or U12391 (N_12391,N_8298,N_10892);
xor U12392 (N_12392,N_11880,N_8881);
or U12393 (N_12393,N_8402,N_9802);
nand U12394 (N_12394,N_9907,N_10876);
nand U12395 (N_12395,N_11342,N_8163);
or U12396 (N_12396,N_8795,N_11710);
xor U12397 (N_12397,N_11279,N_8541);
or U12398 (N_12398,N_11870,N_9847);
nand U12399 (N_12399,N_10274,N_8102);
xor U12400 (N_12400,N_8140,N_9700);
xnor U12401 (N_12401,N_9232,N_11384);
nand U12402 (N_12402,N_10804,N_10216);
nor U12403 (N_12403,N_10881,N_11330);
nor U12404 (N_12404,N_11357,N_11131);
xnor U12405 (N_12405,N_11247,N_10314);
nor U12406 (N_12406,N_11362,N_10574);
nand U12407 (N_12407,N_8596,N_11348);
xnor U12408 (N_12408,N_9195,N_10238);
nor U12409 (N_12409,N_8865,N_10184);
or U12410 (N_12410,N_11924,N_11510);
or U12411 (N_12411,N_8514,N_8260);
xor U12412 (N_12412,N_10666,N_9594);
nor U12413 (N_12413,N_8770,N_11874);
or U12414 (N_12414,N_8373,N_11091);
or U12415 (N_12415,N_11493,N_9625);
nand U12416 (N_12416,N_9903,N_9520);
xnor U12417 (N_12417,N_9138,N_8803);
nand U12418 (N_12418,N_10511,N_9640);
nand U12419 (N_12419,N_8110,N_11887);
nor U12420 (N_12420,N_9062,N_9452);
or U12421 (N_12421,N_9300,N_9710);
and U12422 (N_12422,N_8589,N_11840);
xor U12423 (N_12423,N_11676,N_10386);
or U12424 (N_12424,N_8047,N_9535);
or U12425 (N_12425,N_9667,N_10928);
nor U12426 (N_12426,N_10635,N_11472);
or U12427 (N_12427,N_9219,N_10161);
nand U12428 (N_12428,N_8053,N_10496);
xnor U12429 (N_12429,N_8494,N_8090);
nor U12430 (N_12430,N_11291,N_11894);
and U12431 (N_12431,N_10535,N_10777);
or U12432 (N_12432,N_9977,N_10395);
xor U12433 (N_12433,N_11207,N_10832);
and U12434 (N_12434,N_8382,N_10095);
nor U12435 (N_12435,N_8008,N_8259);
or U12436 (N_12436,N_10456,N_10639);
or U12437 (N_12437,N_10427,N_10276);
xnor U12438 (N_12438,N_11194,N_11541);
xor U12439 (N_12439,N_8869,N_11187);
nand U12440 (N_12440,N_8711,N_8305);
or U12441 (N_12441,N_8185,N_11973);
nand U12442 (N_12442,N_11396,N_9738);
xor U12443 (N_12443,N_9370,N_11043);
nand U12444 (N_12444,N_8329,N_10625);
nor U12445 (N_12445,N_8115,N_11639);
and U12446 (N_12446,N_10385,N_9970);
and U12447 (N_12447,N_10763,N_8224);
and U12448 (N_12448,N_11347,N_10292);
xnor U12449 (N_12449,N_10411,N_8969);
nor U12450 (N_12450,N_11002,N_8079);
and U12451 (N_12451,N_8297,N_10937);
or U12452 (N_12452,N_8735,N_9317);
xor U12453 (N_12453,N_11841,N_8838);
nor U12454 (N_12454,N_9085,N_9978);
nor U12455 (N_12455,N_11427,N_11590);
and U12456 (N_12456,N_8129,N_10417);
xnor U12457 (N_12457,N_9186,N_9950);
xnor U12458 (N_12458,N_9076,N_8085);
or U12459 (N_12459,N_9401,N_9083);
xor U12460 (N_12460,N_8092,N_9395);
and U12461 (N_12461,N_11875,N_11720);
nor U12462 (N_12462,N_8883,N_10223);
and U12463 (N_12463,N_10726,N_9065);
nor U12464 (N_12464,N_11654,N_10155);
xnor U12465 (N_12465,N_9751,N_8279);
nor U12466 (N_12466,N_9797,N_9511);
or U12467 (N_12467,N_11786,N_11593);
or U12468 (N_12468,N_10010,N_9366);
xor U12469 (N_12469,N_10889,N_11143);
xor U12470 (N_12470,N_9946,N_11563);
xnor U12471 (N_12471,N_10481,N_8456);
nor U12472 (N_12472,N_8101,N_11791);
and U12473 (N_12473,N_8543,N_11006);
nor U12474 (N_12474,N_9338,N_8858);
nor U12475 (N_12475,N_11340,N_10682);
and U12476 (N_12476,N_9756,N_11343);
xor U12477 (N_12477,N_9460,N_11478);
nand U12478 (N_12478,N_8245,N_11825);
nand U12479 (N_12479,N_9957,N_11224);
nand U12480 (N_12480,N_8652,N_11552);
or U12481 (N_12481,N_8695,N_11837);
nor U12482 (N_12482,N_10978,N_9321);
xor U12483 (N_12483,N_11534,N_10962);
nand U12484 (N_12484,N_10530,N_11891);
or U12485 (N_12485,N_9754,N_9262);
nand U12486 (N_12486,N_10950,N_8848);
nand U12487 (N_12487,N_9499,N_10173);
or U12488 (N_12488,N_10587,N_9739);
nand U12489 (N_12489,N_11250,N_8585);
nand U12490 (N_12490,N_8694,N_10025);
nor U12491 (N_12491,N_11737,N_11094);
nor U12492 (N_12492,N_9097,N_11739);
nand U12493 (N_12493,N_9582,N_10426);
or U12494 (N_12494,N_11368,N_11858);
or U12495 (N_12495,N_8686,N_11672);
xor U12496 (N_12496,N_8242,N_11447);
nand U12497 (N_12497,N_9623,N_9597);
nor U12498 (N_12498,N_9505,N_8856);
and U12499 (N_12499,N_10714,N_11663);
nand U12500 (N_12500,N_9712,N_8553);
xor U12501 (N_12501,N_11297,N_8441);
or U12502 (N_12502,N_11567,N_10789);
and U12503 (N_12503,N_11338,N_9367);
or U12504 (N_12504,N_10245,N_10559);
nor U12505 (N_12505,N_10979,N_11622);
and U12506 (N_12506,N_11916,N_9985);
xor U12507 (N_12507,N_9398,N_8657);
and U12508 (N_12508,N_10720,N_9860);
and U12509 (N_12509,N_9807,N_9445);
nor U12510 (N_12510,N_9596,N_11765);
xor U12511 (N_12511,N_8459,N_9174);
nor U12512 (N_12512,N_8535,N_9857);
and U12513 (N_12513,N_9430,N_11263);
nor U12514 (N_12514,N_10597,N_9605);
nor U12515 (N_12515,N_10605,N_10247);
and U12516 (N_12516,N_10759,N_11008);
nor U12517 (N_12517,N_11569,N_11561);
nand U12518 (N_12518,N_10965,N_10939);
nand U12519 (N_12519,N_8179,N_8835);
or U12520 (N_12520,N_10953,N_11176);
xor U12521 (N_12521,N_8757,N_8120);
nor U12522 (N_12522,N_8829,N_9125);
nand U12523 (N_12523,N_11052,N_10121);
xnor U12524 (N_12524,N_8162,N_11121);
and U12525 (N_12525,N_9779,N_9331);
or U12526 (N_12526,N_11233,N_10907);
xnor U12527 (N_12527,N_10776,N_11943);
nor U12528 (N_12528,N_9728,N_11162);
nor U12529 (N_12529,N_10356,N_9965);
or U12530 (N_12530,N_10078,N_10000);
and U12531 (N_12531,N_10117,N_11019);
xor U12532 (N_12532,N_8980,N_9772);
or U12533 (N_12533,N_10885,N_8984);
or U12534 (N_12534,N_10042,N_8676);
xor U12535 (N_12535,N_9328,N_8554);
and U12536 (N_12536,N_10528,N_8784);
and U12537 (N_12537,N_9488,N_8139);
nand U12538 (N_12538,N_11208,N_9725);
xor U12539 (N_12539,N_9108,N_8798);
and U12540 (N_12540,N_11197,N_11776);
or U12541 (N_12541,N_11828,N_10634);
nor U12542 (N_12542,N_10140,N_8300);
nand U12543 (N_12543,N_11588,N_10170);
xnor U12544 (N_12544,N_8953,N_10183);
nor U12545 (N_12545,N_10670,N_9692);
and U12546 (N_12546,N_9184,N_11966);
or U12547 (N_12547,N_10867,N_9441);
and U12548 (N_12548,N_10663,N_10270);
xor U12549 (N_12549,N_11925,N_9281);
nor U12550 (N_12550,N_9901,N_11086);
xnor U12551 (N_12551,N_9483,N_8712);
xor U12552 (N_12552,N_8027,N_9102);
nand U12553 (N_12553,N_9168,N_8707);
xor U12554 (N_12554,N_10544,N_9852);
and U12555 (N_12555,N_11626,N_9632);
nor U12556 (N_12556,N_8475,N_11450);
nor U12557 (N_12557,N_11680,N_8285);
xor U12558 (N_12558,N_10735,N_9608);
nand U12559 (N_12559,N_11704,N_10397);
nor U12560 (N_12560,N_11296,N_11260);
nand U12561 (N_12561,N_9723,N_9758);
and U12562 (N_12562,N_11957,N_10827);
nand U12563 (N_12563,N_10781,N_9241);
and U12564 (N_12564,N_9266,N_11310);
or U12565 (N_12565,N_9131,N_10275);
and U12566 (N_12566,N_10562,N_10676);
nand U12567 (N_12567,N_9081,N_10651);
and U12568 (N_12568,N_11532,N_9804);
nor U12569 (N_12569,N_8202,N_11077);
xnor U12570 (N_12570,N_11502,N_10211);
xor U12571 (N_12571,N_9655,N_8715);
nand U12572 (N_12572,N_8957,N_8065);
nand U12573 (N_12573,N_11927,N_11930);
and U12574 (N_12574,N_9310,N_11584);
and U12575 (N_12575,N_9770,N_8273);
or U12576 (N_12576,N_11847,N_9663);
xnor U12577 (N_12577,N_11436,N_11611);
nor U12578 (N_12578,N_8990,N_10514);
xnor U12579 (N_12579,N_9258,N_10377);
xnor U12580 (N_12580,N_9619,N_9564);
or U12581 (N_12581,N_8204,N_9344);
nor U12582 (N_12582,N_11013,N_11860);
and U12583 (N_12583,N_9454,N_10576);
nand U12584 (N_12584,N_8067,N_11205);
nor U12585 (N_12585,N_11085,N_8342);
nand U12586 (N_12586,N_11778,N_9586);
nor U12587 (N_12587,N_10489,N_9649);
nor U12588 (N_12588,N_8389,N_10207);
and U12589 (N_12589,N_9487,N_8976);
nand U12590 (N_12590,N_8172,N_9826);
nand U12591 (N_12591,N_8641,N_8367);
nand U12592 (N_12592,N_9154,N_11512);
nand U12593 (N_12593,N_11146,N_10282);
nand U12594 (N_12594,N_11103,N_8130);
nor U12595 (N_12595,N_9084,N_9722);
nor U12596 (N_12596,N_8606,N_11919);
nor U12597 (N_12597,N_10083,N_11298);
nor U12598 (N_12598,N_9378,N_10076);
nand U12599 (N_12599,N_10396,N_8183);
and U12600 (N_12600,N_9975,N_10388);
nand U12601 (N_12601,N_8235,N_8239);
or U12602 (N_12602,N_10821,N_8351);
nor U12603 (N_12603,N_11658,N_8819);
or U12604 (N_12604,N_10632,N_10289);
or U12605 (N_12605,N_11635,N_10154);
or U12606 (N_12606,N_8256,N_10330);
or U12607 (N_12607,N_8599,N_8663);
nor U12608 (N_12608,N_9628,N_11232);
and U12609 (N_12609,N_8056,N_9233);
and U12610 (N_12610,N_10492,N_11449);
nand U12611 (N_12611,N_10681,N_10567);
xnor U12612 (N_12612,N_10135,N_11609);
xor U12613 (N_12613,N_11607,N_10619);
and U12614 (N_12614,N_11716,N_11903);
nor U12615 (N_12615,N_10595,N_8900);
or U12616 (N_12616,N_11944,N_10924);
nand U12617 (N_12617,N_8658,N_8176);
nor U12618 (N_12618,N_11813,N_10131);
nand U12619 (N_12619,N_9377,N_10599);
xor U12620 (N_12620,N_10384,N_8923);
xnor U12621 (N_12621,N_8653,N_8427);
nand U12622 (N_12622,N_9250,N_8816);
xnor U12623 (N_12623,N_8946,N_11256);
and U12624 (N_12624,N_11503,N_11317);
nor U12625 (N_12625,N_11218,N_9199);
xnor U12626 (N_12626,N_10988,N_11033);
xor U12627 (N_12627,N_10623,N_9403);
and U12628 (N_12628,N_9576,N_8623);
or U12629 (N_12629,N_9822,N_8089);
or U12630 (N_12630,N_10887,N_10972);
nand U12631 (N_12631,N_11989,N_9989);
and U12632 (N_12632,N_9522,N_10171);
and U12633 (N_12633,N_11423,N_8381);
or U12634 (N_12634,N_8062,N_9870);
or U12635 (N_12635,N_9531,N_10717);
nand U12636 (N_12636,N_9368,N_11276);
nor U12637 (N_12637,N_9255,N_11527);
xnor U12638 (N_12638,N_11206,N_8763);
and U12639 (N_12639,N_8563,N_10931);
xor U12640 (N_12640,N_10239,N_8191);
nor U12641 (N_12641,N_10842,N_10744);
nor U12642 (N_12642,N_8831,N_11366);
or U12643 (N_12643,N_11595,N_8739);
nand U12644 (N_12644,N_10254,N_8905);
or U12645 (N_12645,N_8005,N_8320);
or U12646 (N_12646,N_10799,N_11227);
or U12647 (N_12647,N_9861,N_10320);
nor U12648 (N_12648,N_8055,N_8439);
nand U12649 (N_12649,N_10474,N_11490);
xnor U12650 (N_12650,N_9175,N_8855);
nor U12651 (N_12651,N_11544,N_10336);
or U12652 (N_12652,N_8968,N_10826);
and U12653 (N_12653,N_11055,N_9547);
or U12654 (N_12654,N_10766,N_9799);
nand U12655 (N_12655,N_9918,N_11998);
or U12656 (N_12656,N_9830,N_8174);
nand U12657 (N_12657,N_9063,N_9602);
and U12658 (N_12658,N_10908,N_11525);
nand U12659 (N_12659,N_11316,N_11471);
nand U12660 (N_12660,N_10003,N_8769);
nor U12661 (N_12661,N_10812,N_11129);
and U12662 (N_12662,N_9171,N_8104);
xor U12663 (N_12663,N_10023,N_11023);
xor U12664 (N_12664,N_10871,N_10339);
xor U12665 (N_12665,N_9704,N_9028);
and U12666 (N_12666,N_10398,N_9737);
or U12667 (N_12667,N_9387,N_10961);
nor U12668 (N_12668,N_9528,N_10724);
xor U12669 (N_12669,N_9854,N_11747);
nor U12670 (N_12670,N_10582,N_9887);
xnor U12671 (N_12671,N_9645,N_10009);
or U12672 (N_12672,N_9031,N_8252);
or U12673 (N_12673,N_8296,N_11629);
nand U12674 (N_12674,N_11271,N_10938);
xnor U12675 (N_12675,N_11723,N_10218);
or U12676 (N_12676,N_11646,N_8826);
nor U12677 (N_12677,N_10935,N_8075);
or U12678 (N_12678,N_11942,N_11258);
xnor U12679 (N_12679,N_8401,N_10697);
or U12680 (N_12680,N_11700,N_9057);
nor U12681 (N_12681,N_10992,N_11565);
or U12682 (N_12682,N_8083,N_9676);
xor U12683 (N_12683,N_10642,N_8557);
nor U12684 (N_12684,N_8417,N_11025);
nand U12685 (N_12685,N_10693,N_9956);
xor U12686 (N_12686,N_10199,N_9090);
nand U12687 (N_12687,N_8524,N_9899);
nor U12688 (N_12688,N_11177,N_8595);
and U12689 (N_12689,N_10093,N_10475);
and U12690 (N_12690,N_10610,N_9862);
nor U12691 (N_12691,N_11365,N_9465);
and U12692 (N_12692,N_11483,N_10217);
xnor U12693 (N_12693,N_9192,N_10998);
nand U12694 (N_12694,N_10234,N_10328);
or U12695 (N_12695,N_9878,N_8755);
xor U12696 (N_12696,N_9194,N_10856);
xnor U12697 (N_12697,N_10607,N_9304);
or U12698 (N_12698,N_10062,N_10554);
and U12699 (N_12699,N_8180,N_9285);
or U12700 (N_12700,N_11757,N_8344);
nand U12701 (N_12701,N_8871,N_11155);
nand U12702 (N_12702,N_8540,N_9814);
nor U12703 (N_12703,N_9427,N_8675);
nand U12704 (N_12704,N_9732,N_8873);
and U12705 (N_12705,N_10921,N_11939);
nand U12706 (N_12706,N_11548,N_9631);
nor U12707 (N_12707,N_9100,N_9688);
or U12708 (N_12708,N_9187,N_11745);
nor U12709 (N_12709,N_8410,N_10206);
and U12710 (N_12710,N_11401,N_9268);
nor U12711 (N_12711,N_10406,N_11136);
nor U12712 (N_12712,N_10738,N_10703);
or U12713 (N_12713,N_8231,N_9121);
nand U12714 (N_12714,N_8257,N_8290);
nand U12715 (N_12715,N_11430,N_9474);
nor U12716 (N_12716,N_11977,N_11690);
nand U12717 (N_12717,N_8988,N_10723);
and U12718 (N_12718,N_10309,N_9176);
or U12719 (N_12719,N_9222,N_11044);
or U12720 (N_12720,N_8780,N_9777);
and U12721 (N_12721,N_11758,N_9932);
and U12722 (N_12722,N_8852,N_11409);
and U12723 (N_12723,N_11017,N_11497);
nor U12724 (N_12724,N_10151,N_11466);
and U12725 (N_12725,N_10572,N_9614);
nor U12726 (N_12726,N_8849,N_11926);
and U12727 (N_12727,N_8864,N_8098);
nor U12728 (N_12728,N_9127,N_8386);
and U12729 (N_12729,N_9555,N_11461);
or U12730 (N_12730,N_9792,N_9873);
xor U12731 (N_12731,N_11669,N_8161);
nor U12732 (N_12732,N_10479,N_11879);
nand U12733 (N_12733,N_11331,N_11108);
nand U12734 (N_12734,N_10039,N_10226);
nor U12735 (N_12735,N_8493,N_11738);
nor U12736 (N_12736,N_11432,N_9765);
and U12737 (N_12737,N_11299,N_9144);
or U12738 (N_12738,N_9064,N_9841);
and U12739 (N_12739,N_8149,N_10424);
and U12740 (N_12740,N_10260,N_11941);
and U12741 (N_12741,N_11705,N_9947);
or U12742 (N_12742,N_9780,N_9375);
xor U12743 (N_12743,N_9422,N_9086);
nor U12744 (N_12744,N_11711,N_9869);
or U12745 (N_12745,N_11328,N_10202);
xor U12746 (N_12746,N_8420,N_9801);
and U12747 (N_12747,N_9981,N_11859);
nor U12748 (N_12748,N_11810,N_8786);
and U12749 (N_12749,N_10895,N_11135);
and U12750 (N_12750,N_11564,N_11453);
and U12751 (N_12751,N_9316,N_9320);
or U12752 (N_12752,N_11636,N_11811);
nor U12753 (N_12753,N_11833,N_10302);
or U12754 (N_12754,N_9829,N_10830);
and U12755 (N_12755,N_9306,N_11979);
xnor U12756 (N_12756,N_9818,N_9995);
nor U12757 (N_12757,N_9931,N_10366);
nand U12758 (N_12758,N_10421,N_9610);
or U12759 (N_12759,N_9952,N_10818);
nand U12760 (N_12760,N_11460,N_10472);
or U12761 (N_12761,N_10981,N_11431);
nor U12762 (N_12762,N_11489,N_10316);
nand U12763 (N_12763,N_10112,N_10900);
nor U12764 (N_12764,N_8442,N_9240);
or U12765 (N_12765,N_11917,N_8398);
nand U12766 (N_12766,N_8537,N_10344);
nand U12767 (N_12767,N_11804,N_11610);
nor U12768 (N_12768,N_9116,N_11809);
or U12769 (N_12769,N_11733,N_8352);
nor U12770 (N_12770,N_8726,N_10943);
xnor U12771 (N_12771,N_9773,N_8477);
xnor U12772 (N_12772,N_10148,N_8792);
nand U12773 (N_12773,N_11390,N_11933);
and U12774 (N_12774,N_8777,N_8727);
nand U12775 (N_12775,N_11619,N_9669);
nand U12776 (N_12776,N_8705,N_11150);
xor U12777 (N_12777,N_10352,N_9653);
xor U12778 (N_12778,N_9983,N_8527);
xor U12779 (N_12779,N_9484,N_10049);
and U12780 (N_12780,N_10410,N_11402);
and U12781 (N_12781,N_9416,N_8364);
nand U12782 (N_12782,N_9616,N_8876);
and U12783 (N_12783,N_9592,N_10684);
or U12784 (N_12784,N_9159,N_11821);
nand U12785 (N_12785,N_10563,N_10431);
nor U12786 (N_12786,N_11624,N_8859);
nor U12787 (N_12787,N_11376,N_9162);
nor U12788 (N_12788,N_9668,N_8289);
nand U12789 (N_12789,N_9161,N_9322);
xor U12790 (N_12790,N_11528,N_10705);
or U12791 (N_12791,N_11954,N_11419);
and U12792 (N_12792,N_8478,N_8366);
xor U12793 (N_12793,N_11353,N_11374);
and U12794 (N_12794,N_8966,N_8013);
and U12795 (N_12795,N_9228,N_9235);
nand U12796 (N_12796,N_8460,N_11959);
nor U12797 (N_12797,N_11835,N_11170);
and U12798 (N_12798,N_9972,N_9816);
and U12799 (N_12799,N_10443,N_11949);
nor U12800 (N_12800,N_9265,N_9142);
or U12801 (N_12801,N_8078,N_10627);
and U12802 (N_12802,N_9126,N_11802);
xor U12803 (N_12803,N_10762,N_8361);
nor U12804 (N_12804,N_10608,N_11912);
nor U12805 (N_12805,N_10197,N_10438);
or U12806 (N_12806,N_11163,N_8469);
nand U12807 (N_12807,N_11585,N_11606);
nand U12808 (N_12808,N_9390,N_10338);
and U12809 (N_12809,N_8640,N_11225);
and U12810 (N_12810,N_10008,N_9350);
xor U12811 (N_12811,N_11464,N_8581);
nand U12812 (N_12812,N_11037,N_11935);
nor U12813 (N_12813,N_9433,N_11951);
and U12814 (N_12814,N_9225,N_11138);
nor U12815 (N_12815,N_8316,N_10122);
or U12816 (N_12816,N_11164,N_8523);
or U12817 (N_12817,N_8070,N_8116);
nand U12818 (N_12818,N_11531,N_11555);
nand U12819 (N_12819,N_8211,N_9603);
or U12820 (N_12820,N_9730,N_9400);
nor U12821 (N_12821,N_9110,N_10743);
nand U12822 (N_12822,N_9440,N_10603);
and U12823 (N_12823,N_9259,N_10976);
and U12824 (N_12824,N_8218,N_8960);
nand U12825 (N_12825,N_9882,N_9047);
xnor U12826 (N_12826,N_11216,N_11123);
or U12827 (N_12827,N_11172,N_10641);
or U12828 (N_12828,N_8717,N_9025);
or U12829 (N_12829,N_8963,N_8939);
or U12830 (N_12830,N_8051,N_9442);
nand U12831 (N_12831,N_9069,N_9542);
or U12832 (N_12832,N_10373,N_9664);
and U12833 (N_12833,N_11896,N_11687);
nor U12834 (N_12834,N_8582,N_11782);
and U12835 (N_12835,N_11906,N_8451);
or U12836 (N_12836,N_9567,N_11237);
nor U12837 (N_12837,N_11728,N_10956);
or U12838 (N_12838,N_8949,N_8143);
xnor U12839 (N_12839,N_11793,N_10942);
or U12840 (N_12840,N_10072,N_8952);
nor U12841 (N_12841,N_10611,N_10991);
nor U12842 (N_12842,N_11373,N_10849);
and U12843 (N_12843,N_8108,N_9537);
nand U12844 (N_12844,N_10266,N_11101);
nor U12845 (N_12845,N_9143,N_9923);
nor U12846 (N_12846,N_10116,N_10149);
nor U12847 (N_12847,N_9389,N_9699);
nor U12848 (N_12848,N_10449,N_10293);
nor U12849 (N_12849,N_10520,N_8376);
or U12850 (N_12850,N_9015,N_10237);
nand U12851 (N_12851,N_9810,N_10878);
xnor U12852 (N_12852,N_9179,N_9992);
xor U12853 (N_12853,N_11882,N_8925);
or U12854 (N_12854,N_8602,N_11068);
and U12855 (N_12855,N_9434,N_10286);
or U12856 (N_12856,N_10335,N_9070);
xor U12857 (N_12857,N_11559,N_9386);
xor U12858 (N_12858,N_10565,N_9423);
nor U12859 (N_12859,N_10963,N_8892);
or U12860 (N_12860,N_11272,N_9193);
and U12861 (N_12861,N_11038,N_10439);
nand U12862 (N_12862,N_11377,N_9269);
or U12863 (N_12863,N_8404,N_9402);
xor U12864 (N_12864,N_9284,N_11771);
or U12865 (N_12865,N_11246,N_8350);
and U12866 (N_12866,N_8228,N_8001);
xor U12867 (N_12867,N_8571,N_8562);
nand U12868 (N_12868,N_8265,N_10333);
nand U12869 (N_12869,N_11616,N_10990);
nand U12870 (N_12870,N_11007,N_11174);
xnor U12871 (N_12871,N_10017,N_10808);
xnor U12872 (N_12872,N_11371,N_11524);
xor U12873 (N_12873,N_9644,N_10288);
nor U12874 (N_12874,N_11976,N_8832);
xor U12875 (N_12875,N_11278,N_9577);
or U12876 (N_12876,N_8935,N_10690);
nor U12877 (N_12877,N_8877,N_10660);
or U12878 (N_12878,N_11526,N_10783);
and U12879 (N_12879,N_11898,N_9604);
nor U12880 (N_12880,N_8529,N_11712);
nor U12881 (N_12881,N_8250,N_9209);
nor U12882 (N_12882,N_10349,N_9296);
xor U12883 (N_12883,N_9959,N_9252);
nand U12884 (N_12884,N_10866,N_10596);
and U12885 (N_12885,N_8481,N_8588);
and U12886 (N_12886,N_9767,N_10699);
and U12887 (N_12887,N_9935,N_9332);
nand U12888 (N_12888,N_9998,N_9384);
nand U12889 (N_12889,N_8922,N_11360);
xor U12890 (N_12890,N_11270,N_9877);
and U12891 (N_12891,N_8635,N_9482);
nand U12892 (N_12892,N_8928,N_8105);
xnor U12893 (N_12893,N_8743,N_8802);
xnor U12894 (N_12894,N_9466,N_9034);
or U12895 (N_12895,N_9122,N_8506);
or U12896 (N_12896,N_10294,N_10797);
nand U12897 (N_12897,N_10615,N_11854);
and U12898 (N_12898,N_10389,N_10589);
nor U12899 (N_12899,N_8736,N_8088);
nor U12900 (N_12900,N_10082,N_11383);
or U12901 (N_12901,N_9279,N_8897);
nor U12902 (N_12902,N_11760,N_8380);
nand U12903 (N_12903,N_9342,N_9673);
and U12904 (N_12904,N_11681,N_8808);
xnor U12905 (N_12905,N_9415,N_10296);
nor U12906 (N_12906,N_8137,N_11416);
nand U12907 (N_12907,N_10793,N_9457);
or U12908 (N_12908,N_11719,N_9833);
nor U12909 (N_12909,N_10527,N_10877);
nor U12910 (N_12910,N_8258,N_11144);
or U12911 (N_12911,N_11165,N_9543);
and U12912 (N_12912,N_8747,N_8511);
and U12913 (N_12913,N_11920,N_10505);
nand U12914 (N_12914,N_8338,N_11424);
xor U12915 (N_12915,N_10591,N_8902);
nand U12916 (N_12916,N_9074,N_8962);
xor U12917 (N_12917,N_8830,N_8255);
nor U12918 (N_12918,N_10210,N_11132);
nand U12919 (N_12919,N_8731,N_8299);
or U12920 (N_12920,N_8627,N_11686);
nand U12921 (N_12921,N_8687,N_8713);
or U12922 (N_12922,N_11476,N_9418);
or U12923 (N_12923,N_8559,N_10343);
nand U12924 (N_12924,N_10263,N_11275);
xnor U12925 (N_12925,N_11190,N_8718);
nand U12926 (N_12926,N_10662,N_10200);
nor U12927 (N_12927,N_9507,N_11283);
and U12928 (N_12928,N_10689,N_8123);
xnor U12929 (N_12929,N_9785,N_11169);
xnor U12930 (N_12930,N_8870,N_11321);
xnor U12931 (N_12931,N_8042,N_9682);
and U12932 (N_12932,N_9896,N_11026);
and U12933 (N_12933,N_11307,N_10543);
and U12934 (N_12934,N_8490,N_10108);
or U12935 (N_12935,N_8046,N_9609);
or U12936 (N_12936,N_11761,N_11971);
and U12937 (N_12937,N_8930,N_11110);
nand U12938 (N_12938,N_9937,N_11158);
nor U12939 (N_12939,N_9588,N_10461);
nand U12940 (N_12940,N_9053,N_8396);
or U12941 (N_12941,N_11867,N_9421);
nand U12942 (N_12942,N_11011,N_11277);
or U12943 (N_12943,N_11800,N_11994);
xnor U12944 (N_12944,N_9180,N_9858);
nor U12945 (N_12945,N_10624,N_8467);
and U12946 (N_12946,N_10033,N_10823);
nand U12947 (N_12947,N_9217,N_8322);
and U12948 (N_12948,N_9618,N_9717);
and U12949 (N_12949,N_11620,N_10147);
or U12950 (N_12950,N_10012,N_9455);
or U12951 (N_12951,N_10775,N_11093);
or U12952 (N_12952,N_9456,N_8811);
and U12953 (N_12953,N_10740,N_11186);
xor U12954 (N_12954,N_9089,N_9641);
or U12955 (N_12955,N_10817,N_8360);
xor U12956 (N_12956,N_10679,N_10606);
nand U12957 (N_12957,N_11281,N_8394);
nand U12958 (N_12958,N_8601,N_10045);
xor U12959 (N_12959,N_8799,N_11230);
nor U12960 (N_12960,N_8546,N_9561);
nand U12961 (N_12961,N_11081,N_9601);
nor U12962 (N_12962,N_9763,N_11952);
nor U12963 (N_12963,N_11481,N_11648);
and U12964 (N_12964,N_10917,N_10920);
nor U12965 (N_12965,N_8783,N_10391);
and U12966 (N_12966,N_9502,N_10524);
or U12967 (N_12967,N_11262,N_10688);
xnor U12968 (N_12968,N_8800,N_8310);
nor U12969 (N_12969,N_10022,N_9695);
or U12970 (N_12970,N_11562,N_8022);
nor U12971 (N_12971,N_10174,N_11157);
and U12972 (N_12972,N_9292,N_8059);
and U12973 (N_12973,N_11118,N_11668);
nand U12974 (N_12974,N_8347,N_9109);
xnor U12975 (N_12975,N_10486,N_11947);
or U12976 (N_12976,N_8833,N_10501);
xor U12977 (N_12977,N_8662,N_10925);
xor U12978 (N_12978,N_11699,N_8806);
and U12979 (N_12979,N_11608,N_11443);
xor U12980 (N_12980,N_10027,N_10322);
nand U12981 (N_12981,N_10739,N_10874);
xor U12982 (N_12982,N_8937,N_11287);
and U12983 (N_12983,N_11991,N_9855);
nor U12984 (N_12984,N_9990,N_10034);
nor U12985 (N_12985,N_8207,N_8330);
xnor U12986 (N_12986,N_11397,N_10191);
and U12987 (N_12987,N_8522,N_8779);
and U12988 (N_12988,N_11128,N_10845);
nor U12989 (N_12989,N_11836,N_10809);
xor U12990 (N_12990,N_8217,N_9917);
nand U12991 (N_12991,N_9453,N_10841);
or U12992 (N_12992,N_8234,N_11408);
or U12993 (N_12993,N_10383,N_10273);
and U12994 (N_12994,N_8198,N_9757);
or U12995 (N_12995,N_10187,N_10393);
or U12996 (N_12996,N_9048,N_8884);
and U12997 (N_12997,N_10982,N_10803);
or U12998 (N_12998,N_11656,N_8480);
xnor U12999 (N_12999,N_11446,N_10497);
or U13000 (N_13000,N_10159,N_11439);
or U13001 (N_13001,N_10553,N_9766);
nor U13002 (N_13002,N_10674,N_10854);
nand U13003 (N_13003,N_11124,N_10106);
or U13004 (N_13004,N_11120,N_8045);
nand U13005 (N_13005,N_11028,N_11313);
nand U13006 (N_13006,N_8124,N_9124);
nand U13007 (N_13007,N_9485,N_8903);
or U13008 (N_13008,N_11709,N_9794);
xnor U13009 (N_13009,N_9012,N_9011);
and U13010 (N_13010,N_10773,N_10614);
or U13011 (N_13011,N_11934,N_9289);
or U13012 (N_13012,N_10080,N_10853);
or U13013 (N_13013,N_9469,N_11413);
nor U13014 (N_13014,N_9458,N_9040);
xor U13015 (N_13015,N_10716,N_10546);
nor U13016 (N_13016,N_10280,N_8248);
nand U13017 (N_13017,N_9264,N_9795);
nand U13018 (N_13018,N_11468,N_11491);
xor U13019 (N_13019,N_11909,N_11113);
and U13020 (N_13020,N_8488,N_10507);
nor U13021 (N_13021,N_9004,N_9117);
nor U13022 (N_13022,N_8132,N_11398);
and U13023 (N_13023,N_8753,N_8193);
xor U13024 (N_13024,N_9747,N_10659);
or U13025 (N_13025,N_11387,N_11644);
and U13026 (N_13026,N_8335,N_11406);
nor U13027 (N_13027,N_9745,N_8898);
and U13028 (N_13028,N_9997,N_11754);
nand U13029 (N_13029,N_9207,N_8371);
or U13030 (N_13030,N_9383,N_11566);
and U13031 (N_13031,N_8164,N_10675);
nor U13032 (N_13032,N_11203,N_11918);
nand U13033 (N_13033,N_11071,N_8225);
nand U13034 (N_13034,N_8578,N_8216);
nor U13035 (N_13035,N_9498,N_10440);
and U13036 (N_13036,N_10829,N_9253);
nor U13037 (N_13037,N_10262,N_9521);
xnor U13038 (N_13038,N_8422,N_9615);
and U13039 (N_13039,N_11805,N_10016);
nor U13040 (N_13040,N_8015,N_10779);
nor U13041 (N_13041,N_9140,N_9708);
or U13042 (N_13042,N_11803,N_10490);
xor U13043 (N_13043,N_11269,N_11215);
nor U13044 (N_13044,N_8333,N_9231);
or U13045 (N_13045,N_8696,N_9169);
or U13046 (N_13046,N_8052,N_11451);
and U13047 (N_13047,N_8851,N_9512);
and U13048 (N_13048,N_9376,N_9880);
nor U13049 (N_13049,N_9892,N_10787);
nor U13050 (N_13050,N_10473,N_8465);
or U13051 (N_13051,N_8730,N_11161);
xor U13052 (N_13052,N_8974,N_11744);
or U13053 (N_13053,N_9369,N_11993);
and U13054 (N_13054,N_8134,N_10712);
nor U13055 (N_13055,N_11580,N_11241);
and U13056 (N_13056,N_11617,N_8503);
or U13057 (N_13057,N_9133,N_10024);
nor U13058 (N_13058,N_9409,N_11034);
nand U13059 (N_13059,N_8762,N_8508);
xnor U13060 (N_13060,N_8620,N_8071);
and U13061 (N_13061,N_11477,N_10538);
nor U13062 (N_13062,N_8321,N_9001);
nor U13063 (N_13063,N_9287,N_11004);
or U13064 (N_13064,N_8186,N_9327);
and U13065 (N_13065,N_10403,N_11220);
or U13066 (N_13066,N_10629,N_8433);
xnor U13067 (N_13067,N_10190,N_11905);
xor U13068 (N_13068,N_8141,N_9912);
nand U13069 (N_13069,N_10160,N_8891);
xnor U13070 (N_13070,N_8219,N_11642);
xnor U13071 (N_13071,N_8412,N_8872);
nor U13072 (N_13072,N_11987,N_10028);
and U13073 (N_13073,N_10521,N_10061);
xnor U13074 (N_13074,N_8615,N_8021);
or U13075 (N_13075,N_9129,N_9414);
nand U13076 (N_13076,N_11795,N_10198);
nor U13077 (N_13077,N_11799,N_10453);
and U13078 (N_13078,N_10721,N_10464);
or U13079 (N_13079,N_11314,N_9500);
nand U13080 (N_13080,N_9731,N_9927);
xnor U13081 (N_13081,N_11293,N_11369);
and U13082 (N_13082,N_9463,N_11499);
and U13083 (N_13083,N_8483,N_9111);
or U13084 (N_13084,N_9030,N_9638);
nand U13085 (N_13085,N_9188,N_11982);
or U13086 (N_13086,N_8880,N_9971);
and U13087 (N_13087,N_11539,N_9846);
xnor U13088 (N_13088,N_9242,N_11238);
nor U13089 (N_13089,N_10858,N_10408);
nor U13090 (N_13090,N_10179,N_8948);
nor U13091 (N_13091,N_10882,N_8644);
or U13092 (N_13092,N_9686,N_10115);
nand U13093 (N_13093,N_11223,N_8492);
and U13094 (N_13094,N_11769,N_11741);
nor U13095 (N_13095,N_9746,N_10195);
nand U13096 (N_13096,N_9898,N_9412);
nor U13097 (N_13097,N_9571,N_11119);
nor U13098 (N_13098,N_8253,N_8068);
and U13099 (N_13099,N_11261,N_10698);
nor U13100 (N_13100,N_9021,N_11516);
nor U13101 (N_13101,N_10091,N_10983);
nor U13102 (N_13102,N_9943,N_10996);
nor U13103 (N_13103,N_11697,N_11104);
nor U13104 (N_13104,N_11411,N_8518);
nor U13105 (N_13105,N_11815,N_10548);
nor U13106 (N_13106,N_10831,N_8854);
and U13107 (N_13107,N_10692,N_10130);
nor U13108 (N_13108,N_8945,N_9019);
nand U13109 (N_13109,N_8998,N_11881);
and U13110 (N_13110,N_9221,N_9056);
nor U13111 (N_13111,N_9444,N_11140);
or U13112 (N_13112,N_10952,N_11282);
nor U13113 (N_13113,N_9018,N_11441);
or U13114 (N_13114,N_11660,N_8270);
nor U13115 (N_13115,N_8673,N_9881);
or U13116 (N_13116,N_10729,N_11095);
or U13117 (N_13117,N_11783,N_11781);
nand U13118 (N_13118,N_9337,N_8722);
or U13119 (N_13119,N_10303,N_9920);
xnor U13120 (N_13120,N_8639,N_10129);
nand U13121 (N_13121,N_11199,N_11219);
nand U13122 (N_13122,N_10801,N_9821);
or U13123 (N_13123,N_11444,N_9036);
and U13124 (N_13124,N_9578,N_10706);
nand U13125 (N_13125,N_9022,N_11507);
or U13126 (N_13126,N_11543,N_11536);
or U13127 (N_13127,N_10880,N_8583);
and U13128 (N_13128,N_9593,N_11863);
or U13129 (N_13129,N_11730,N_11087);
nand U13130 (N_13130,N_8613,N_9590);
xor U13131 (N_13131,N_8513,N_11253);
xor U13132 (N_13132,N_9519,N_9968);
or U13133 (N_13133,N_8020,N_9589);
xnor U13134 (N_13134,N_9107,N_10590);
and U13135 (N_13135,N_9055,N_10649);
nor U13136 (N_13136,N_8822,N_10750);
xor U13137 (N_13137,N_8122,N_9690);
xor U13138 (N_13138,N_11115,N_10621);
nor U13139 (N_13139,N_8975,N_11638);
or U13140 (N_13140,N_10348,N_10932);
and U13141 (N_13141,N_11907,N_11152);
xor U13142 (N_13142,N_9523,N_11214);
nand U13143 (N_13143,N_9149,N_10770);
and U13144 (N_13144,N_10094,N_9811);
and U13145 (N_13145,N_10890,N_8610);
nor U13146 (N_13146,N_11766,N_8889);
or U13147 (N_13147,N_11305,N_9883);
and U13148 (N_13148,N_8267,N_9334);
xor U13149 (N_13149,N_8586,N_10020);
and U13150 (N_13150,N_9459,N_10923);
nand U13151 (N_13151,N_9986,N_8278);
nand U13152 (N_13152,N_10153,N_11228);
nand U13153 (N_13153,N_8509,N_9683);
nand U13154 (N_13154,N_10290,N_8345);
nand U13155 (N_13155,N_9467,N_10236);
nand U13156 (N_13156,N_11586,N_8555);
xnor U13157 (N_13157,N_11185,N_8719);
nand U13158 (N_13158,N_10601,N_11613);
or U13159 (N_13159,N_10214,N_8230);
or U13160 (N_13160,N_8538,N_9839);
nand U13161 (N_13161,N_10598,N_8956);
xnor U13162 (N_13162,N_9652,N_11718);
nand U13163 (N_13163,N_8093,N_8774);
nand U13164 (N_13164,N_10227,N_10047);
nand U13165 (N_13165,N_10857,N_11239);
xnor U13166 (N_13166,N_10870,N_8916);
nor U13167 (N_13167,N_8941,N_9570);
nand U13168 (N_13168,N_11345,N_9919);
nor U13169 (N_13169,N_11213,N_11500);
nor U13170 (N_13170,N_9197,N_8728);
and U13171 (N_13171,N_9743,N_8397);
and U13172 (N_13172,N_11667,N_11774);
nor U13173 (N_13173,N_8530,N_9940);
or U13174 (N_13174,N_10454,N_9218);
nand U13175 (N_13175,N_9872,N_9607);
xor U13176 (N_13176,N_9534,N_9944);
nand U13177 (N_13177,N_9077,N_9573);
nor U13178 (N_13178,N_8742,N_10099);
or U13179 (N_13179,N_8693,N_8655);
xnor U13180 (N_13180,N_8408,N_8765);
and U13181 (N_13181,N_10267,N_9962);
and U13182 (N_13182,N_10418,N_11280);
nor U13183 (N_13183,N_8206,N_10884);
xnor U13184 (N_13184,N_9356,N_11355);
nor U13185 (N_13185,N_11173,N_10678);
nand U13186 (N_13186,N_10054,N_8418);
nand U13187 (N_13187,N_9925,N_11708);
or U13188 (N_13188,N_8862,N_10730);
or U13189 (N_13189,N_9404,N_8570);
nand U13190 (N_13190,N_11254,N_11075);
nor U13191 (N_13191,N_10631,N_9842);
and U13192 (N_13192,N_10863,N_11405);
and U13193 (N_13193,N_8919,N_8121);
or U13194 (N_13194,N_8025,N_9560);
nor U13195 (N_13195,N_8737,N_11599);
xor U13196 (N_13196,N_11222,N_10488);
or U13197 (N_13197,N_11958,N_9330);
or U13198 (N_13198,N_11817,N_8339);
nand U13199 (N_13199,N_8621,N_8393);
nand U13200 (N_13200,N_8943,N_8882);
nor U13201 (N_13201,N_8499,N_8241);
or U13202 (N_13202,N_10791,N_11193);
xor U13203 (N_13203,N_10164,N_10307);
nand U13204 (N_13204,N_10364,N_10819);
xor U13205 (N_13205,N_9468,N_11693);
nor U13206 (N_13206,N_8170,N_11621);
nor U13207 (N_13207,N_11356,N_8240);
or U13208 (N_13208,N_8438,N_8254);
xnor U13209 (N_13209,N_8788,N_8388);
xnor U13210 (N_13210,N_8415,N_8890);
or U13211 (N_13211,N_10279,N_8377);
xnor U13212 (N_13212,N_10162,N_8629);
nor U13213 (N_13213,N_9924,N_10442);
or U13214 (N_13214,N_9711,N_11679);
xnor U13215 (N_13215,N_8690,N_10556);
or U13216 (N_13216,N_8233,N_8561);
xnor U13217 (N_13217,N_9223,N_10914);
nand U13218 (N_13218,N_9145,N_8634);
or U13219 (N_13219,N_8048,N_11594);
or U13220 (N_13220,N_11252,N_11549);
nand U13221 (N_13221,N_8237,N_8672);
nand U13222 (N_13222,N_11049,N_11022);
nor U13223 (N_13223,N_10502,N_9230);
xor U13224 (N_13224,N_9824,N_9789);
xnor U13225 (N_13225,N_8643,N_10192);
nand U13226 (N_13226,N_9139,N_10100);
and U13227 (N_13227,N_8987,N_11827);
xnor U13228 (N_13228,N_9114,N_9591);
or U13229 (N_13229,N_11678,N_8751);
or U13230 (N_13230,N_11587,N_8729);
xor U13231 (N_13231,N_11312,N_8303);
nor U13232 (N_13232,N_11159,N_10114);
nor U13233 (N_13233,N_8760,N_10312);
or U13234 (N_13234,N_11137,N_8646);
or U13235 (N_13235,N_8618,N_9035);
nor U13236 (N_13236,N_10204,N_8453);
nor U13237 (N_13237,N_9868,N_10375);
xor U13238 (N_13238,N_9748,N_10755);
nor U13239 (N_13239,N_11059,N_9208);
and U13240 (N_13240,N_8282,N_9798);
nand U13241 (N_13241,N_10673,N_9494);
nand U13242 (N_13242,N_11713,N_8434);
nand U13243 (N_13243,N_11130,N_10796);
or U13244 (N_13244,N_9016,N_8999);
nor U13245 (N_13245,N_11311,N_9760);
and U13246 (N_13246,N_9246,N_11359);
xor U13247 (N_13247,N_8405,N_10902);
nor U13248 (N_13248,N_8824,N_9461);
nand U13249 (N_13249,N_8766,N_9227);
xor U13250 (N_13250,N_10069,N_8951);
and U13251 (N_13251,N_10295,N_9895);
xnor U13252 (N_13252,N_11410,N_11191);
nor U13253 (N_13253,N_9492,N_8487);
xnor U13254 (N_13254,N_8723,N_8407);
nor U13255 (N_13255,N_11612,N_8901);
nor U13256 (N_13256,N_11972,N_11469);
or U13257 (N_13257,N_8266,N_9546);
nor U13258 (N_13258,N_9096,N_9257);
nor U13259 (N_13259,N_8293,N_8649);
nand U13260 (N_13260,N_11459,N_8823);
and U13261 (N_13261,N_10476,N_11098);
nor U13262 (N_13262,N_10102,N_10533);
and U13263 (N_13263,N_11694,N_11300);
or U13264 (N_13264,N_11303,N_11673);
xor U13265 (N_13265,N_10564,N_11337);
xnor U13266 (N_13266,N_9311,N_9123);
or U13267 (N_13267,N_11627,N_8836);
xor U13268 (N_13268,N_10194,N_8861);
xnor U13269 (N_13269,N_10450,N_8359);
nor U13270 (N_13270,N_10181,N_8772);
nand U13271 (N_13271,N_9752,N_8192);
or U13272 (N_13272,N_8809,N_11647);
or U13273 (N_13273,N_11452,N_11180);
nor U13274 (N_13274,N_11488,N_9916);
nand U13275 (N_13275,N_9182,N_9204);
or U13276 (N_13276,N_11231,N_10566);
or U13277 (N_13277,N_11294,N_10331);
nor U13278 (N_13278,N_8166,N_11641);
nand U13279 (N_13279,N_10420,N_8458);
nor U13280 (N_13280,N_11391,N_11465);
and U13281 (N_13281,N_10936,N_11834);
or U13282 (N_13282,N_10362,N_8781);
xor U13283 (N_13283,N_9346,N_11474);
xnor U13284 (N_13284,N_10997,N_11454);
nand U13285 (N_13285,N_9270,N_11339);
and U13286 (N_13286,N_9051,N_8189);
xnor U13287 (N_13287,N_8926,N_11284);
and U13288 (N_13288,N_8741,N_8326);
and U13289 (N_13289,N_10137,N_11576);
nand U13290 (N_13290,N_9215,N_10092);
nand U13291 (N_13291,N_11480,N_9277);
and U13292 (N_13292,N_11386,N_8158);
xor U13293 (N_13293,N_9529,N_8384);
nor U13294 (N_13294,N_10761,N_11063);
or U13295 (N_13295,N_9600,N_8395);
xor U13296 (N_13296,N_10256,N_8857);
or U13297 (N_13297,N_10048,N_10329);
nand U13298 (N_13298,N_11866,N_9674);
nand U13299 (N_13299,N_9372,N_9774);
and U13300 (N_13300,N_8229,N_9897);
nor U13301 (N_13301,N_10665,N_11571);
or U13302 (N_13302,N_11787,N_9203);
xnor U13303 (N_13303,N_9691,N_9141);
xnor U13304 (N_13304,N_8651,N_8220);
nor U13305 (N_13305,N_10402,N_9464);
xor U13306 (N_13306,N_9023,N_10222);
and U13307 (N_13307,N_8472,N_11715);
and U13308 (N_13308,N_10758,N_10163);
or U13309 (N_13309,N_9749,N_11725);
nor U13310 (N_13310,N_8972,N_9718);
nor U13311 (N_13311,N_10742,N_10811);
and U13312 (N_13312,N_8519,N_10298);
xor U13313 (N_13313,N_10447,N_8896);
nand U13314 (N_13314,N_11403,N_9091);
or U13315 (N_13315,N_9666,N_9817);
and U13316 (N_13316,N_10229,N_10974);
or U13317 (N_13317,N_9974,N_11762);
or U13318 (N_13318,N_11792,N_11117);
nand U13319 (N_13319,N_10495,N_11166);
and U13320 (N_13320,N_8000,N_11508);
nand U13321 (N_13321,N_11671,N_9967);
nand U13322 (N_13322,N_9479,N_10568);
or U13323 (N_13323,N_9563,N_9806);
and U13324 (N_13324,N_10719,N_10732);
or U13325 (N_13325,N_10946,N_9532);
nor U13326 (N_13326,N_9198,N_10212);
nand U13327 (N_13327,N_8590,N_9424);
or U13328 (N_13328,N_11518,N_8813);
nand U13329 (N_13329,N_9933,N_10323);
nor U13330 (N_13330,N_9633,N_9911);
xnor U13331 (N_13331,N_10029,N_10136);
or U13332 (N_13332,N_8050,N_9428);
and U13333 (N_13333,N_10110,N_9768);
and U13334 (N_13334,N_10101,N_9288);
and U13335 (N_13335,N_10847,N_11039);
nor U13336 (N_13336,N_8227,N_9431);
or U13337 (N_13337,N_10090,N_11226);
and U13338 (N_13338,N_8684,N_9808);
or U13339 (N_13339,N_10999,N_11422);
and U13340 (N_13340,N_9489,N_9357);
or U13341 (N_13341,N_11400,N_10342);
or U13342 (N_13342,N_10306,N_9002);
and U13343 (N_13343,N_10512,N_10337);
or U13344 (N_13344,N_8894,N_8845);
and U13345 (N_13345,N_10980,N_11067);
nand U13346 (N_13346,N_10261,N_9120);
nand U13347 (N_13347,N_11643,N_8057);
nand U13348 (N_13348,N_11015,N_10244);
nand U13349 (N_13349,N_11820,N_8785);
or U13350 (N_13350,N_8677,N_11630);
or U13351 (N_13351,N_10516,N_10281);
nor U13352 (N_13352,N_9791,N_11211);
nand U13353 (N_13353,N_8014,N_8888);
and U13354 (N_13354,N_9082,N_11623);
and U13355 (N_13355,N_8400,N_11980);
or U13356 (N_13356,N_11600,N_8023);
or U13357 (N_13357,N_9735,N_10123);
xnor U13358 (N_13358,N_10782,N_10656);
xnor U13359 (N_13359,N_9303,N_8981);
nor U13360 (N_13360,N_11742,N_9539);
xor U13361 (N_13361,N_9172,N_9006);
xor U13362 (N_13362,N_10655,N_11181);
and U13363 (N_13363,N_11865,N_8024);
nand U13364 (N_13364,N_11984,N_11798);
and U13365 (N_13365,N_11707,N_8409);
nor U13366 (N_13366,N_8111,N_11897);
and U13367 (N_13367,N_9624,N_8043);
or U13368 (N_13368,N_11790,N_8645);
and U13369 (N_13369,N_10964,N_11603);
or U13370 (N_13370,N_8392,N_8146);
and U13371 (N_13371,N_10144,N_11445);
nor U13372 (N_13372,N_8791,N_9099);
nor U13373 (N_13373,N_9654,N_9973);
xnor U13374 (N_13374,N_11855,N_11849);
xnor U13375 (N_13375,N_11992,N_9803);
xor U13376 (N_13376,N_9813,N_11812);
and U13377 (N_13377,N_8313,N_11985);
nor U13378 (N_13378,N_8706,N_11234);
xor U13379 (N_13379,N_8495,N_10111);
and U13380 (N_13380,N_9282,N_8077);
and U13381 (N_13381,N_11777,N_11763);
nand U13382 (N_13382,N_11047,N_10653);
xnor U13383 (N_13383,N_11268,N_9113);
xnor U13384 (N_13384,N_10053,N_10357);
or U13385 (N_13385,N_9856,N_8801);
nand U13386 (N_13386,N_10545,N_8778);
nor U13387 (N_13387,N_8959,N_10041);
nor U13388 (N_13388,N_10378,N_9324);
or U13389 (N_13389,N_10879,N_9894);
xor U13390 (N_13390,N_8911,N_10233);
xor U13391 (N_13391,N_10208,N_8992);
or U13392 (N_13392,N_10536,N_8097);
nor U13393 (N_13393,N_9098,N_8125);
xnor U13394 (N_13394,N_10581,N_10040);
or U13395 (N_13395,N_10429,N_10494);
nor U13396 (N_13396,N_11964,N_11010);
or U13397 (N_13397,N_8474,N_10060);
nor U13398 (N_13398,N_9533,N_9295);
or U13399 (N_13399,N_11764,N_9960);
or U13400 (N_13400,N_11830,N_11872);
nor U13401 (N_13401,N_10075,N_11850);
nand U13402 (N_13402,N_10139,N_9759);
or U13403 (N_13403,N_10213,N_10513);
nor U13404 (N_13404,N_9104,N_8091);
nand U13405 (N_13405,N_8054,N_10630);
and U13406 (N_13406,N_10452,N_10984);
nor U13407 (N_13407,N_8263,N_10405);
or U13408 (N_13408,N_9392,N_11589);
xor U13409 (N_13409,N_9996,N_10571);
nand U13410 (N_13410,N_10392,N_11509);
xnor U13411 (N_13411,N_8626,N_10896);
nand U13412 (N_13412,N_9713,N_11041);
and U13413 (N_13413,N_8828,N_8875);
or U13414 (N_13414,N_8614,N_8700);
nor U13415 (N_13415,N_11701,N_8683);
nand U13416 (N_13416,N_9574,N_10534);
nor U13417 (N_13417,N_8463,N_8648);
and U13418 (N_13418,N_10304,N_8793);
and U13419 (N_13419,N_10865,N_8982);
and U13420 (N_13420,N_9514,N_9680);
nor U13421 (N_13421,N_10468,N_11435);
nor U13422 (N_13422,N_11463,N_8879);
nor U13423 (N_13423,N_10620,N_8917);
xor U13424 (N_13424,N_8283,N_10685);
xnor U13425 (N_13425,N_9448,N_8660);
and U13426 (N_13426,N_11842,N_8448);
nor U13427 (N_13427,N_9778,N_11099);
and U13428 (N_13428,N_8867,N_11392);
or U13429 (N_13429,N_10252,N_9697);
nand U13430 (N_13430,N_9694,N_10387);
xor U13431 (N_13431,N_8378,N_8178);
nor U13432 (N_13432,N_10484,N_9476);
xnor U13433 (N_13433,N_9622,N_8584);
and U13434 (N_13434,N_10225,N_8157);
nand U13435 (N_13435,N_11304,N_11012);
nor U13436 (N_13436,N_8208,N_9493);
and U13437 (N_13437,N_8385,N_9394);
xnor U13438 (N_13438,N_10725,N_9355);
nand U13439 (N_13439,N_9750,N_10994);
xor U13440 (N_13440,N_9439,N_8423);
or U13441 (N_13441,N_9477,N_9647);
nand U13442 (N_13442,N_10119,N_11082);
nor U13443 (N_13443,N_8018,N_9155);
nand U13444 (N_13444,N_8118,N_8009);
nand U13445 (N_13445,N_8973,N_10604);
nor U13446 (N_13446,N_9486,N_11097);
or U13447 (N_13447,N_8650,N_8138);
and U13448 (N_13448,N_10551,N_10506);
nor U13449 (N_13449,N_8028,N_11200);
nor U13450 (N_13450,N_8725,N_9361);
and U13451 (N_13451,N_10107,N_11688);
nor U13452 (N_13452,N_8275,N_10550);
and U13453 (N_13453,N_9510,N_10633);
or U13454 (N_13454,N_9853,N_9672);
xnor U13455 (N_13455,N_9626,N_11326);
or U13456 (N_13456,N_8642,N_11288);
nor U13457 (N_13457,N_8287,N_9961);
and U13458 (N_13458,N_10752,N_9982);
or U13459 (N_13459,N_9513,N_9156);
nand U13460 (N_13460,N_11395,N_11090);
nor U13461 (N_13461,N_11955,N_9307);
and U13462 (N_13462,N_10272,N_11030);
xnor U13463 (N_13463,N_10052,N_8247);
and U13464 (N_13464,N_10713,N_8574);
xor U13465 (N_13465,N_8594,N_9646);
and U13466 (N_13466,N_8096,N_8906);
and U13467 (N_13467,N_8213,N_11914);
or U13468 (N_13468,N_8979,N_9381);
nand U13469 (N_13469,N_11198,N_9491);
and U13470 (N_13470,N_8033,N_8844);
or U13471 (N_13471,N_9629,N_10968);
nor U13472 (N_13472,N_11634,N_9783);
nand U13473 (N_13473,N_10754,N_8552);
nor U13474 (N_13474,N_9684,N_8918);
and U13475 (N_13475,N_8112,N_11080);
nor U13476 (N_13476,N_8497,N_11329);
nor U13477 (N_13477,N_10778,N_11251);
and U13478 (N_13478,N_8182,N_9238);
or U13479 (N_13479,N_10109,N_8107);
xnor U13480 (N_13480,N_11102,N_11434);
and U13481 (N_13481,N_10374,N_10836);
nor U13482 (N_13482,N_10741,N_10002);
nand U13483 (N_13483,N_8637,N_9480);
nor U13484 (N_13484,N_9689,N_9042);
nand U13485 (N_13485,N_11794,N_11533);
xor U13486 (N_13486,N_9471,N_11775);
nor U13487 (N_13487,N_10299,N_10358);
xor U13488 (N_13488,N_8709,N_8271);
xnor U13489 (N_13489,N_11192,N_11615);
or U13490 (N_13490,N_10224,N_11822);
nor U13491 (N_13491,N_10771,N_9524);
nand U13492 (N_13492,N_11614,N_9068);
xnor U13493 (N_13493,N_10609,N_11784);
nor U13494 (N_13494,N_11309,N_8512);
and U13495 (N_13495,N_11248,N_10986);
xor U13496 (N_13496,N_9323,N_9130);
nor U13497 (N_13497,N_8087,N_10746);
or U13498 (N_13498,N_10189,N_9849);
nand U13499 (N_13499,N_11937,N_9443);
nand U13500 (N_13500,N_10015,N_8636);
nand U13501 (N_13501,N_8424,N_8038);
and U13502 (N_13502,N_10310,N_9226);
nor U13503 (N_13503,N_8567,N_11625);
nand U13504 (N_13504,N_8927,N_10989);
or U13505 (N_13505,N_9341,N_9256);
xnor U13506 (N_13506,N_8940,N_8908);
or U13507 (N_13507,N_11717,N_10555);
nand U13508 (N_13508,N_9007,N_11302);
nand U13509 (N_13509,N_8212,N_10324);
xnor U13510 (N_13510,N_10822,N_10063);
or U13511 (N_13511,N_11370,N_11649);
nor U13512 (N_13512,N_9984,N_11988);
nand U13513 (N_13513,N_8505,N_9538);
nand U13514 (N_13514,N_10118,N_8099);
or U13515 (N_13515,N_9575,N_10594);
and U13516 (N_13516,N_10346,N_8665);
nor U13517 (N_13517,N_10089,N_11873);
nand U13518 (N_13518,N_9239,N_9627);
xor U13519 (N_13519,N_9569,N_8947);
xnor U13520 (N_13520,N_9734,N_10059);
xnor U13521 (N_13521,N_8965,N_8430);
nand U13522 (N_13522,N_9435,N_11378);
nand U13523 (N_13523,N_9793,N_8030);
nand U13524 (N_13524,N_11913,N_11910);
or U13525 (N_13525,N_11962,N_10691);
nor U13526 (N_13526,N_8337,N_10230);
nor U13527 (N_13527,N_10113,N_11618);
nor U13528 (N_13528,N_8796,N_9753);
xnor U13529 (N_13529,N_10379,N_10561);
and U13530 (N_13530,N_8012,N_10205);
and U13531 (N_13531,N_10541,N_11196);
nand U13532 (N_13532,N_9286,N_8679);
xor U13533 (N_13533,N_9501,N_9205);
nor U13534 (N_13534,N_11899,N_10005);
nand U13535 (N_13535,N_8429,N_8910);
nand U13536 (N_13536,N_9202,N_11462);
and U13537 (N_13537,N_11308,N_9696);
nand U13538 (N_13538,N_8994,N_10737);
nor U13539 (N_13539,N_8341,N_8426);
or U13540 (N_13540,N_9966,N_11886);
xor U13541 (N_13541,N_8209,N_11494);
or U13542 (N_13542,N_9720,N_10518);
or U13543 (N_13543,N_10084,N_10365);
nor U13544 (N_13544,N_11035,N_9112);
nor U13545 (N_13545,N_10446,N_8548);
nor U13546 (N_13546,N_8482,N_9726);
and U13547 (N_13547,N_8308,N_9681);
nand U13548 (N_13548,N_11932,N_8274);
xor U13549 (N_13549,N_10677,N_8144);
nand U13550 (N_13550,N_8002,N_9294);
nand U13551 (N_13551,N_11147,N_10843);
nor U13552 (N_13552,N_8387,N_10255);
and U13553 (N_13553,N_11582,N_10718);
nor U13554 (N_13554,N_9013,N_8841);
or U13555 (N_13555,N_8084,N_10509);
xnor U13556 (N_13556,N_10736,N_9158);
nor U13557 (N_13557,N_11570,N_10400);
or U13558 (N_13558,N_9297,N_10810);
and U13559 (N_13559,N_11772,N_10166);
and U13560 (N_13560,N_9875,N_9891);
and U13561 (N_13561,N_8479,N_9061);
or U13562 (N_13562,N_11818,N_11496);
nand U13563 (N_13563,N_11969,N_8331);
nor U13564 (N_13564,N_11361,N_8425);
xor U13565 (N_13565,N_10246,N_8521);
and U13566 (N_13566,N_10326,N_9243);
or U13567 (N_13567,N_11996,N_9039);
nor U13568 (N_13568,N_11407,N_8117);
xnor U13569 (N_13569,N_11749,N_11632);
and U13570 (N_13570,N_8236,N_8040);
xnor U13571 (N_13571,N_11856,N_9637);
nor U13572 (N_13572,N_9729,N_8612);
nor U13573 (N_13573,N_8670,N_9634);
nand U13574 (N_13574,N_10455,N_8375);
xnor U13575 (N_13575,N_10425,N_9980);
and U13576 (N_13576,N_8565,N_11148);
nand U13577 (N_13577,N_11689,N_8996);
nor U13578 (N_13578,N_8210,N_10575);
or U13579 (N_13579,N_9506,N_10257);
nand U13580 (N_13580,N_11558,N_11520);
or U13581 (N_13581,N_11290,N_11018);
and U13582 (N_13582,N_10354,N_8878);
xnor U13583 (N_13583,N_8520,N_9953);
xor U13584 (N_13584,N_10071,N_11212);
nand U13585 (N_13585,N_11421,N_10891);
nor U13586 (N_13586,N_9902,N_9866);
nor U13587 (N_13587,N_11568,N_11557);
nand U13588 (N_13588,N_8362,N_10483);
and U13589 (N_13589,N_8572,N_10128);
and U13590 (N_13590,N_9024,N_11547);
nand U13591 (N_13591,N_8276,N_8195);
and U13592 (N_13592,N_11645,N_10913);
xnor U13593 (N_13593,N_10949,N_9396);
nor U13594 (N_13594,N_8306,N_11092);
xnor U13595 (N_13595,N_9410,N_9515);
or U13596 (N_13596,N_9969,N_9371);
and U13597 (N_13597,N_10077,N_9420);
nor U13598 (N_13598,N_10066,N_10800);
or U13599 (N_13599,N_9905,N_9835);
nand U13600 (N_13600,N_8607,N_11750);
and U13601 (N_13601,N_10277,N_10132);
nor U13602 (N_13602,N_11535,N_8312);
or U13603 (N_13603,N_10401,N_8545);
nor U13604 (N_13604,N_11990,N_11864);
nor U13605 (N_13605,N_9189,N_8603);
or U13606 (N_13606,N_10470,N_8470);
or U13607 (N_13607,N_11244,N_10141);
or U13608 (N_13608,N_9397,N_11078);
xnor U13609 (N_13609,N_11522,N_9825);
xnor U13610 (N_13610,N_8598,N_10334);
nor U13611 (N_13611,N_9419,N_8815);
xor U13612 (N_13612,N_11285,N_10085);
or U13613 (N_13613,N_11438,N_8749);
xor U13614 (N_13614,N_9921,N_10838);
nor U13615 (N_13615,N_8904,N_9071);
xnor U13616 (N_13616,N_9900,N_9851);
or U13617 (N_13617,N_8284,N_11650);
nand U13618 (N_13618,N_9963,N_8136);
and U13619 (N_13619,N_8787,N_8704);
xnor U13620 (N_13620,N_11578,N_11878);
or U13621 (N_13621,N_8991,N_9029);
xor U13622 (N_13622,N_10127,N_11844);
nor U13623 (N_13623,N_8294,N_9436);
nand U13624 (N_13624,N_9177,N_8498);
or U13625 (N_13625,N_8821,N_10820);
nand U13626 (N_13626,N_8744,N_8775);
nand U13627 (N_13627,N_8661,N_11853);
xor U13628 (N_13628,N_9834,N_8419);
nand U13629 (N_13629,N_8558,N_10894);
xor U13630 (N_13630,N_9724,N_11072);
nand U13631 (N_13631,N_10855,N_11542);
nand U13632 (N_13632,N_10560,N_10967);
nor U13633 (N_13633,N_9333,N_9041);
nand U13634 (N_13634,N_11861,N_8580);
nand U13635 (N_13635,N_9819,N_8150);
nor U13636 (N_13636,N_9058,N_11848);
nor U13637 (N_13637,N_8732,N_8600);
nor U13638 (N_13638,N_10850,N_8912);
and U13639 (N_13639,N_8995,N_11670);
and U13640 (N_13640,N_8666,N_9786);
nand U13641 (N_13641,N_11945,N_8773);
and U13642 (N_13642,N_10004,N_10618);
or U13643 (N_13643,N_9473,N_8688);
or U13644 (N_13644,N_8064,N_11257);
or U13645 (N_13645,N_8550,N_10435);
xor U13646 (N_13646,N_8721,N_10748);
nor U13647 (N_13647,N_10593,N_9702);
and U13648 (N_13648,N_9119,N_9657);
nand U13649 (N_13649,N_10142,N_10428);
or U13650 (N_13650,N_9599,N_9727);
nor U13651 (N_13651,N_8200,N_8159);
or U13652 (N_13652,N_9010,N_11467);
xnor U13653 (N_13653,N_11975,N_11073);
and U13654 (N_13654,N_11380,N_10221);
nand U13655 (N_13655,N_11141,N_9643);
and U13656 (N_13656,N_9388,N_10539);
nand U13657 (N_13657,N_10491,N_8173);
and U13658 (N_13658,N_8249,N_11323);
and U13659 (N_13659,N_8556,N_10182);
xnor U13660 (N_13660,N_10232,N_9994);
xor U13661 (N_13661,N_8678,N_11031);
nor U13662 (N_13662,N_11832,N_8476);
nand U13663 (N_13663,N_11505,N_9080);
nor U13664 (N_13664,N_11631,N_9429);
nor U13665 (N_13665,N_11900,N_11901);
or U13666 (N_13666,N_11684,N_10898);
and U13667 (N_13667,N_10193,N_8147);
nor U13668 (N_13668,N_11633,N_10767);
nand U13669 (N_13669,N_11983,N_9809);
or U13670 (N_13670,N_10909,N_10828);
and U13671 (N_13671,N_8336,N_10196);
nand U13672 (N_13672,N_9345,N_8154);
and U13673 (N_13673,N_10901,N_11145);
xnor U13674 (N_13674,N_8909,N_9865);
or U13675 (N_13675,N_9562,N_10765);
and U13676 (N_13676,N_10549,N_8450);
and U13677 (N_13677,N_11414,N_10911);
or U13678 (N_13678,N_9987,N_8246);
nand U13679 (N_13679,N_10814,N_10638);
or U13680 (N_13680,N_9210,N_8989);
or U13681 (N_13681,N_11950,N_8114);
or U13682 (N_13682,N_10569,N_11292);
xor U13683 (N_13683,N_11530,N_11003);
and U13684 (N_13684,N_8638,N_8874);
and U13685 (N_13685,N_11485,N_8440);
or U13686 (N_13686,N_11698,N_11889);
nor U13687 (N_13687,N_9449,N_8983);
nor U13688 (N_13688,N_8681,N_9828);
nand U13689 (N_13689,N_11417,N_11240);
and U13690 (N_13690,N_10929,N_11674);
nand U13691 (N_13691,N_9886,N_11259);
nor U13692 (N_13692,N_8860,N_9475);
xnor U13693 (N_13693,N_9611,N_9399);
xnor U13694 (N_13694,N_10145,N_10862);
xor U13695 (N_13695,N_10172,N_8624);
nor U13696 (N_13696,N_10300,N_11974);
nand U13697 (N_13697,N_10508,N_10954);
xnor U13698 (N_13698,N_8593,N_10709);
or U13699 (N_13699,N_10525,N_9598);
or U13700 (N_13700,N_9942,N_8551);
nor U13701 (N_13701,N_11429,N_11088);
nor U13702 (N_13702,N_9405,N_10046);
nor U13703 (N_13703,N_9037,N_10430);
and U13704 (N_13704,N_10457,N_10955);
nand U13705 (N_13705,N_10552,N_8669);
nor U13706 (N_13706,N_10602,N_8106);
or U13707 (N_13707,N_10150,N_9432);
nor U13708 (N_13708,N_11139,N_8931);
or U13709 (N_13709,N_9651,N_8215);
xor U13710 (N_13710,N_11814,N_11255);
xor U13711 (N_13711,N_10558,N_10930);
xor U13712 (N_13712,N_10504,N_9152);
and U13713 (N_13713,N_10933,N_9701);
and U13714 (N_13714,N_11597,N_9859);
and U13715 (N_13715,N_10918,N_11074);
nor U13716 (N_13716,N_11350,N_8171);
nand U13717 (N_13717,N_11415,N_9044);
nor U13718 (N_13718,N_9659,N_9557);
xor U13719 (N_13719,N_10616,N_9290);
nand U13720 (N_13720,N_9548,N_8632);
nor U13721 (N_13721,N_8319,N_9929);
or U13722 (N_13722,N_8489,N_8656);
nor U13723 (N_13723,N_11591,N_8399);
nand U13724 (N_13724,N_9160,N_11501);
xor U13725 (N_13725,N_9349,N_9079);
nor U13726 (N_13726,N_9812,N_9679);
and U13727 (N_13727,N_11696,N_11746);
xor U13728 (N_13728,N_8383,N_10626);
nand U13729 (N_13729,N_11756,N_8358);
nor U13730 (N_13730,N_11583,N_9078);
xor U13731 (N_13731,N_11070,N_11722);
or U13732 (N_13732,N_9893,N_9884);
and U13733 (N_13733,N_9904,N_8812);
xnor U13734 (N_13734,N_10341,N_10471);
nand U13735 (N_13735,N_8899,N_8302);
xor U13736 (N_13736,N_11682,N_8814);
xor U13737 (N_13737,N_9353,N_10126);
nand U13738 (N_13738,N_9741,N_10037);
and U13739 (N_13739,N_10519,N_9580);
or U13740 (N_13740,N_10960,N_11367);
xnor U13741 (N_13741,N_8533,N_8734);
xnor U13742 (N_13742,N_10795,N_9661);
nand U13743 (N_13743,N_9336,N_8680);
xor U13744 (N_13744,N_11845,N_9787);
and U13745 (N_13745,N_10848,N_8268);
nand U13746 (N_13746,N_8391,N_11178);
nor U13747 (N_13747,N_11484,N_8964);
or U13748 (N_13748,N_8834,N_11970);
nor U13749 (N_13749,N_8746,N_9771);
and U13750 (N_13750,N_10369,N_10165);
and U13751 (N_13751,N_11596,N_10407);
nor U13752 (N_13752,N_9052,N_9587);
or U13753 (N_13753,N_10846,N_8842);
nor U13754 (N_13754,N_10157,N_10284);
and U13755 (N_13755,N_10580,N_9639);
and U13756 (N_13756,N_8840,N_10167);
nor U13757 (N_13757,N_11273,N_11202);
and U13758 (N_13758,N_9363,N_8127);
and U13759 (N_13759,N_11838,N_11773);
nor U13760 (N_13760,N_11921,N_10540);
xor U13761 (N_13761,N_11458,N_11714);
xor U13762 (N_13762,N_10051,N_8073);
nand U13763 (N_13763,N_8379,N_11986);
and U13764 (N_13764,N_11540,N_8443);
nand U13765 (N_13765,N_9955,N_8026);
nor U13766 (N_13766,N_8978,N_8292);
and U13767 (N_13767,N_9273,N_8039);
nor U13768 (N_13768,N_11274,N_9206);
and U13769 (N_13769,N_8447,N_8286);
nor U13770 (N_13770,N_11581,N_8411);
xnor U13771 (N_13771,N_9359,N_8421);
and U13772 (N_13772,N_8309,N_9354);
and U13773 (N_13773,N_8205,N_9343);
or U13774 (N_13774,N_10708,N_10463);
nor U13775 (N_13775,N_10070,N_10971);
nand U13776 (N_13776,N_11801,N_8767);
or U13777 (N_13777,N_8295,N_8534);
nand U13778 (N_13778,N_11997,N_8790);
xnor U13779 (N_13779,N_11675,N_9049);
and U13780 (N_13780,N_9426,N_10248);
or U13781 (N_13781,N_10340,N_10897);
xor U13782 (N_13782,N_10647,N_10813);
or U13783 (N_13783,N_8325,N_10271);
or U13784 (N_13784,N_9566,N_10175);
xor U13785 (N_13785,N_10707,N_10869);
nor U13786 (N_13786,N_9775,N_8223);
nor U13787 (N_13787,N_11105,N_10382);
nor U13788 (N_13788,N_9451,N_9526);
or U13789 (N_13789,N_10893,N_9518);
xnor U13790 (N_13790,N_10969,N_10757);
nand U13791 (N_13791,N_11057,N_9261);
or U13792 (N_13792,N_11807,N_8413);
or U13793 (N_13793,N_9606,N_9733);
and U13794 (N_13794,N_9224,N_9190);
nor U13795 (N_13795,N_8221,N_9148);
nor U13796 (N_13796,N_10661,N_10073);
nor U13797 (N_13797,N_10035,N_9517);
or U13798 (N_13798,N_8074,N_10498);
xnor U13799 (N_13799,N_11182,N_11106);
nand U13800 (N_13800,N_10973,N_9705);
or U13801 (N_13801,N_10806,N_9438);
xnor U13802 (N_13802,N_10701,N_9838);
nand U13803 (N_13803,N_8887,N_11127);
nor U13804 (N_13804,N_11752,N_11160);
xnor U13805 (N_13805,N_9941,N_11770);
or U13806 (N_13806,N_11324,N_8846);
and U13807 (N_13807,N_9559,N_9906);
or U13808 (N_13808,N_8301,N_11657);
or U13809 (N_13809,N_11056,N_10577);
nor U13810 (N_13810,N_10423,N_11437);
xnor U13811 (N_13811,N_11046,N_10840);
xor U13812 (N_13812,N_11319,N_10657);
xnor U13813 (N_13813,N_11895,N_9762);
xor U13814 (N_13814,N_9568,N_11652);
nand U13815 (N_13815,N_8119,N_11393);
nor U13816 (N_13816,N_8007,N_10243);
nand U13817 (N_13817,N_9707,N_10786);
nor U13818 (N_13818,N_9260,N_8264);
or U13819 (N_13819,N_9201,N_9319);
nor U13820 (N_13820,N_11806,N_9948);
xnor U13821 (N_13821,N_9504,N_10315);
or U13822 (N_13822,N_10588,N_10098);
and U13823 (N_13823,N_8668,N_8544);
and U13824 (N_13824,N_11289,N_8853);
nand U13825 (N_13825,N_10764,N_10993);
xor U13826 (N_13826,N_9374,N_9393);
and U13827 (N_13827,N_8485,N_10844);
or U13828 (N_13828,N_10250,N_11236);
or U13829 (N_13829,N_10745,N_11346);
nor U13830 (N_13830,N_9764,N_10959);
and U13831 (N_13831,N_8701,N_8473);
nor U13832 (N_13832,N_11995,N_10711);
nand U13833 (N_13833,N_8501,N_8667);
and U13834 (N_13834,N_10220,N_11819);
and U13835 (N_13835,N_10780,N_11096);
and U13836 (N_13836,N_10785,N_11789);
and U13837 (N_13837,N_11948,N_11154);
nor U13838 (N_13838,N_8716,N_10586);
nand U13839 (N_13839,N_11885,N_8720);
xnor U13840 (N_13840,N_8406,N_11005);
nor U13841 (N_13841,N_8768,N_9470);
nand U13842 (N_13842,N_9658,N_8516);
or U13843 (N_13843,N_9554,N_10798);
xor U13844 (N_13844,N_10578,N_10258);
nand U13845 (N_13845,N_10313,N_8913);
nor U13846 (N_13846,N_11816,N_10096);
xnor U13847 (N_13847,N_11884,N_11922);
nand U13848 (N_13848,N_10947,N_10074);
nor U13849 (N_13849,N_10466,N_9776);
xor U13850 (N_13850,N_9979,N_8664);
nor U13851 (N_13851,N_11779,N_9934);
and U13852 (N_13852,N_10839,N_8689);
nor U13853 (N_13853,N_11923,N_9716);
nor U13854 (N_13854,N_11375,N_8452);
and U13855 (N_13855,N_11908,N_9165);
and U13856 (N_13856,N_8622,N_8933);
nor U13857 (N_13857,N_9670,N_11053);
nor U13858 (N_13858,N_11051,N_11179);
xnor U13859 (N_13859,N_11551,N_9613);
nor U13860 (N_13860,N_11457,N_8576);
nand U13861 (N_13861,N_8587,N_10669);
or U13862 (N_13862,N_8280,N_10904);
nor U13863 (N_13863,N_8924,N_9305);
or U13864 (N_13864,N_9541,N_11029);
nor U13865 (N_13865,N_8682,N_10056);
nor U13866 (N_13866,N_9005,N_8568);
or U13867 (N_13867,N_9660,N_10948);
or U13868 (N_13868,N_11229,N_11418);
nor U13869 (N_13869,N_9781,N_11956);
xor U13870 (N_13870,N_11604,N_8349);
xnor U13871 (N_13871,N_11938,N_10251);
or U13872 (N_13872,N_9274,N_9736);
xor U13873 (N_13873,N_10672,N_8818);
xor U13874 (N_13874,N_11683,N_9740);
or U13875 (N_13875,N_10203,N_10702);
and U13876 (N_13876,N_9009,N_11946);
or U13877 (N_13877,N_9147,N_11851);
nand U13878 (N_13878,N_9072,N_10381);
nor U13879 (N_13879,N_8126,N_8365);
nand U13880 (N_13880,N_10645,N_8332);
nand U13881 (N_13881,N_9879,N_9936);
or U13882 (N_13882,N_10977,N_10311);
and U13883 (N_13883,N_8566,N_8547);
nor U13884 (N_13884,N_8659,N_8579);
nand U13885 (N_13885,N_10043,N_10922);
or U13886 (N_13886,N_10995,N_11149);
nand U13887 (N_13887,N_8370,N_9339);
nor U13888 (N_13888,N_9325,N_8181);
nor U13889 (N_13889,N_9516,N_8986);
nand U13890 (N_13890,N_11267,N_11640);
xnor U13891 (N_13891,N_8748,N_9863);
nand U13892 (N_13892,N_9267,N_10305);
xor U13893 (N_13893,N_9211,N_9650);
xor U13894 (N_13894,N_10860,N_9115);
and U13895 (N_13895,N_10467,N_8471);
nor U13896 (N_13896,N_9312,N_11695);
xnor U13897 (N_13897,N_8944,N_9066);
and U13898 (N_13898,N_11204,N_9003);
and U13899 (N_13899,N_11333,N_8738);
or U13900 (N_13900,N_8029,N_11936);
and U13901 (N_13901,N_10919,N_8416);
or U13902 (N_13902,N_10105,N_10478);
nand U13903 (N_13903,N_8932,N_9163);
nor U13904 (N_13904,N_11442,N_8631);
nand U13905 (N_13905,N_11083,N_11659);
and U13906 (N_13906,N_11084,N_8004);
xor U13907 (N_13907,N_10637,N_11032);
or U13908 (N_13908,N_9151,N_9497);
xnor U13909 (N_13909,N_9413,N_11188);
nor U13910 (N_13910,N_11245,N_10668);
nand U13911 (N_13911,N_8674,N_11217);
xnor U13912 (N_13912,N_9462,N_8837);
nor U13913 (N_13913,N_8369,N_11967);
nand U13914 (N_13914,N_10176,N_9060);
xor U13915 (N_13915,N_10700,N_8261);
nand U13916 (N_13916,N_10680,N_10104);
xor U13917 (N_13917,N_8740,N_9092);
nand U13918 (N_13918,N_8745,N_9788);
nand U13919 (N_13919,N_10570,N_10081);
or U13920 (N_13920,N_11839,N_9088);
xor U13921 (N_13921,N_9544,N_9263);
nand U13922 (N_13922,N_9220,N_10751);
nand U13923 (N_13923,N_9620,N_8710);
or U13924 (N_13924,N_11911,N_10671);
nand U13925 (N_13925,N_9150,N_10057);
or U13926 (N_13926,N_9677,N_10640);
or U13927 (N_13927,N_8457,N_10055);
and U13928 (N_13928,N_9909,N_11156);
nand U13929 (N_13929,N_10944,N_11151);
or U13930 (N_13930,N_9790,N_8985);
or U13931 (N_13931,N_8515,N_8517);
nor U13932 (N_13932,N_11753,N_9939);
or U13933 (N_13933,N_8764,N_9054);
and U13934 (N_13934,N_11487,N_11826);
nand U13935 (N_13935,N_11892,N_11515);
nand U13936 (N_13936,N_9558,N_11862);
or U13937 (N_13937,N_8971,N_9867);
nand U13938 (N_13938,N_11036,N_9508);
and U13939 (N_13939,N_10794,N_9137);
or U13940 (N_13940,N_8754,N_9302);
or U13941 (N_13941,N_9157,N_8977);
nand U13942 (N_13942,N_9769,N_11440);
and U13943 (N_13943,N_8752,N_9583);
nor U13944 (N_13944,N_11831,N_8431);
xor U13945 (N_13945,N_10636,N_9364);
xnor U13946 (N_13946,N_8625,N_11666);
or U13947 (N_13947,N_10370,N_11315);
or U13948 (N_13948,N_8311,N_11824);
xor U13949 (N_13949,N_10951,N_11931);
and U13950 (N_13950,N_11364,N_11869);
or U13951 (N_13951,N_11554,N_9181);
and U13952 (N_13952,N_10361,N_8885);
nand U13953 (N_13953,N_8604,N_10355);
xor U13954 (N_13954,N_8850,N_8628);
and U13955 (N_13955,N_8006,N_11385);
nor U13956 (N_13956,N_9173,N_11341);
nand U13957 (N_13957,N_11470,N_9360);
or U13958 (N_13958,N_9915,N_10517);
or U13959 (N_13959,N_11426,N_9584);
and U13960 (N_13960,N_11249,N_11550);
nand U13961 (N_13961,N_11999,N_11111);
nor U13962 (N_13962,N_11189,N_8691);
xnor U13963 (N_13963,N_11295,N_9685);
nand U13964 (N_13964,N_10888,N_8363);
or U13965 (N_13965,N_9212,N_11066);
or U13966 (N_13966,N_9308,N_11651);
or U13967 (N_13967,N_11514,N_11042);
xnor U13968 (N_13968,N_11014,N_8491);
or U13969 (N_13969,N_9755,N_8461);
xor U13970 (N_13970,N_10658,N_8466);
nor U13971 (N_13971,N_8446,N_8549);
xor U13972 (N_13972,N_10585,N_9890);
nand U13973 (N_13973,N_8175,N_8094);
xor U13974 (N_13974,N_8804,N_8942);
xnor U13975 (N_13975,N_9721,N_9185);
nand U13976 (N_13976,N_10987,N_11598);
nor U13977 (N_13977,N_9278,N_8291);
nor U13978 (N_13978,N_10710,N_9340);
xor U13979 (N_13979,N_11334,N_8577);
or U13980 (N_13980,N_11412,N_8165);
nand U13981 (N_13981,N_10031,N_10477);
xor U13982 (N_13982,N_11389,N_10790);
nand U13983 (N_13983,N_8177,N_10728);
or U13984 (N_13984,N_9291,N_9678);
nand U13985 (N_13985,N_9843,N_10185);
and U13986 (N_13986,N_8100,N_8936);
and U13987 (N_13987,N_10833,N_11963);
nand U13988 (N_13988,N_9796,N_11210);
nand U13989 (N_13989,N_10883,N_11628);
nand U13990 (N_13990,N_11344,N_9425);
and U13991 (N_13991,N_9050,N_10249);
or U13992 (N_13992,N_10036,N_11498);
nor U13993 (N_13993,N_10287,N_11601);
nor U13994 (N_13994,N_11054,N_9550);
nand U13995 (N_13995,N_11349,N_8152);
and U13996 (N_13996,N_11116,N_9067);
nand U13997 (N_13997,N_8403,N_9167);
nor U13998 (N_13998,N_9922,N_9365);
nor U13999 (N_13999,N_11482,N_10612);
xor U14000 (N_14000,N_10450,N_9373);
and U14001 (N_14001,N_9770,N_8069);
xor U14002 (N_14002,N_10326,N_11637);
or U14003 (N_14003,N_11427,N_9875);
or U14004 (N_14004,N_11735,N_11449);
xnor U14005 (N_14005,N_9282,N_10177);
nor U14006 (N_14006,N_10290,N_8542);
nor U14007 (N_14007,N_11520,N_11316);
nand U14008 (N_14008,N_8659,N_11138);
nand U14009 (N_14009,N_11817,N_11513);
nor U14010 (N_14010,N_10916,N_11197);
xor U14011 (N_14011,N_11652,N_9179);
and U14012 (N_14012,N_11576,N_8409);
and U14013 (N_14013,N_11987,N_8732);
nor U14014 (N_14014,N_10384,N_9344);
or U14015 (N_14015,N_10690,N_11539);
or U14016 (N_14016,N_11249,N_11615);
or U14017 (N_14017,N_11038,N_9889);
or U14018 (N_14018,N_10126,N_11963);
xnor U14019 (N_14019,N_9775,N_11997);
xnor U14020 (N_14020,N_11294,N_10915);
and U14021 (N_14021,N_9434,N_8149);
xor U14022 (N_14022,N_10722,N_10090);
and U14023 (N_14023,N_11683,N_10738);
or U14024 (N_14024,N_10945,N_11175);
nand U14025 (N_14025,N_11807,N_9909);
or U14026 (N_14026,N_8711,N_10666);
nand U14027 (N_14027,N_8060,N_10565);
xnor U14028 (N_14028,N_10996,N_9249);
nor U14029 (N_14029,N_11257,N_8863);
nor U14030 (N_14030,N_11481,N_11403);
or U14031 (N_14031,N_9959,N_11994);
or U14032 (N_14032,N_11599,N_10986);
and U14033 (N_14033,N_9159,N_9240);
or U14034 (N_14034,N_8588,N_8806);
xor U14035 (N_14035,N_9170,N_10143);
nor U14036 (N_14036,N_8295,N_8259);
xor U14037 (N_14037,N_11001,N_11030);
nand U14038 (N_14038,N_8352,N_9220);
nand U14039 (N_14039,N_11077,N_8424);
or U14040 (N_14040,N_10025,N_10965);
nor U14041 (N_14041,N_11595,N_9066);
and U14042 (N_14042,N_11832,N_8543);
nor U14043 (N_14043,N_10844,N_8440);
nand U14044 (N_14044,N_8025,N_9699);
nor U14045 (N_14045,N_10429,N_10100);
nor U14046 (N_14046,N_8839,N_10984);
and U14047 (N_14047,N_8304,N_9129);
nor U14048 (N_14048,N_10690,N_11887);
nand U14049 (N_14049,N_8903,N_9635);
or U14050 (N_14050,N_8144,N_10410);
nand U14051 (N_14051,N_8322,N_10989);
nor U14052 (N_14052,N_11706,N_8029);
nand U14053 (N_14053,N_10417,N_10596);
xor U14054 (N_14054,N_9287,N_9354);
nand U14055 (N_14055,N_10827,N_8199);
nor U14056 (N_14056,N_10688,N_11364);
xnor U14057 (N_14057,N_9015,N_10335);
xor U14058 (N_14058,N_9236,N_8900);
and U14059 (N_14059,N_8641,N_10348);
xor U14060 (N_14060,N_9370,N_10512);
xnor U14061 (N_14061,N_10363,N_8897);
and U14062 (N_14062,N_8463,N_10265);
and U14063 (N_14063,N_9718,N_10241);
nand U14064 (N_14064,N_9608,N_11480);
and U14065 (N_14065,N_10836,N_8185);
nand U14066 (N_14066,N_11032,N_10275);
nor U14067 (N_14067,N_11586,N_11257);
and U14068 (N_14068,N_8694,N_9907);
or U14069 (N_14069,N_9455,N_8443);
and U14070 (N_14070,N_8234,N_10337);
and U14071 (N_14071,N_8541,N_8820);
xor U14072 (N_14072,N_10177,N_11614);
or U14073 (N_14073,N_9106,N_11115);
xor U14074 (N_14074,N_11032,N_8266);
nand U14075 (N_14075,N_11212,N_9262);
xnor U14076 (N_14076,N_8791,N_8615);
xnor U14077 (N_14077,N_10752,N_11499);
xor U14078 (N_14078,N_9451,N_9267);
xor U14079 (N_14079,N_11063,N_8333);
xnor U14080 (N_14080,N_11589,N_11737);
or U14081 (N_14081,N_10827,N_11757);
and U14082 (N_14082,N_11437,N_11945);
xor U14083 (N_14083,N_8292,N_8099);
or U14084 (N_14084,N_9263,N_9459);
nand U14085 (N_14085,N_9573,N_10357);
and U14086 (N_14086,N_11046,N_10485);
nor U14087 (N_14087,N_11111,N_11948);
and U14088 (N_14088,N_11352,N_10278);
or U14089 (N_14089,N_8507,N_8949);
and U14090 (N_14090,N_9258,N_8177);
or U14091 (N_14091,N_11531,N_9846);
nand U14092 (N_14092,N_10413,N_10947);
or U14093 (N_14093,N_8625,N_10286);
xor U14094 (N_14094,N_11764,N_8331);
or U14095 (N_14095,N_8370,N_9497);
xor U14096 (N_14096,N_11423,N_11016);
nor U14097 (N_14097,N_8457,N_8990);
or U14098 (N_14098,N_10456,N_8485);
and U14099 (N_14099,N_8866,N_8398);
xnor U14100 (N_14100,N_8509,N_10175);
or U14101 (N_14101,N_8318,N_11800);
xor U14102 (N_14102,N_8147,N_8796);
xor U14103 (N_14103,N_8979,N_8351);
nor U14104 (N_14104,N_10232,N_9044);
and U14105 (N_14105,N_10459,N_11898);
or U14106 (N_14106,N_8935,N_9473);
or U14107 (N_14107,N_11109,N_10535);
nand U14108 (N_14108,N_10724,N_10666);
or U14109 (N_14109,N_9994,N_11090);
nor U14110 (N_14110,N_9057,N_8852);
nor U14111 (N_14111,N_11463,N_10243);
or U14112 (N_14112,N_10374,N_8851);
nand U14113 (N_14113,N_10029,N_10591);
and U14114 (N_14114,N_9176,N_8605);
nand U14115 (N_14115,N_10272,N_8278);
and U14116 (N_14116,N_9938,N_8524);
nand U14117 (N_14117,N_10197,N_10830);
and U14118 (N_14118,N_9763,N_11361);
or U14119 (N_14119,N_9971,N_11916);
and U14120 (N_14120,N_10072,N_8296);
nor U14121 (N_14121,N_8160,N_9462);
xnor U14122 (N_14122,N_9828,N_9933);
nor U14123 (N_14123,N_10566,N_9702);
and U14124 (N_14124,N_11458,N_10908);
nand U14125 (N_14125,N_11793,N_10304);
xnor U14126 (N_14126,N_8610,N_10733);
nor U14127 (N_14127,N_9664,N_10061);
or U14128 (N_14128,N_9287,N_11247);
or U14129 (N_14129,N_8023,N_8381);
nand U14130 (N_14130,N_11299,N_9921);
and U14131 (N_14131,N_11121,N_8419);
nand U14132 (N_14132,N_8294,N_9283);
or U14133 (N_14133,N_10614,N_11438);
nand U14134 (N_14134,N_11506,N_11992);
and U14135 (N_14135,N_10854,N_11516);
nand U14136 (N_14136,N_10448,N_8013);
xnor U14137 (N_14137,N_11748,N_9015);
and U14138 (N_14138,N_9072,N_9235);
or U14139 (N_14139,N_10452,N_9200);
and U14140 (N_14140,N_8532,N_9363);
nand U14141 (N_14141,N_10653,N_11713);
nand U14142 (N_14142,N_10724,N_8527);
and U14143 (N_14143,N_9729,N_11203);
xnor U14144 (N_14144,N_8745,N_10495);
and U14145 (N_14145,N_9731,N_10312);
nand U14146 (N_14146,N_9155,N_10770);
xor U14147 (N_14147,N_8070,N_10323);
or U14148 (N_14148,N_8041,N_9701);
nand U14149 (N_14149,N_8776,N_11314);
or U14150 (N_14150,N_10716,N_8951);
xnor U14151 (N_14151,N_10300,N_11077);
xor U14152 (N_14152,N_9217,N_10635);
or U14153 (N_14153,N_10556,N_8814);
nor U14154 (N_14154,N_9454,N_10181);
and U14155 (N_14155,N_10672,N_10087);
and U14156 (N_14156,N_10572,N_8419);
and U14157 (N_14157,N_9586,N_11015);
nor U14158 (N_14158,N_11401,N_9378);
nor U14159 (N_14159,N_9569,N_8169);
nand U14160 (N_14160,N_10474,N_8452);
or U14161 (N_14161,N_11428,N_9473);
or U14162 (N_14162,N_11718,N_8798);
or U14163 (N_14163,N_11123,N_9494);
and U14164 (N_14164,N_11796,N_8270);
or U14165 (N_14165,N_8871,N_8056);
and U14166 (N_14166,N_9187,N_11110);
and U14167 (N_14167,N_9727,N_8725);
nor U14168 (N_14168,N_11687,N_9597);
or U14169 (N_14169,N_10468,N_10781);
xor U14170 (N_14170,N_11018,N_11553);
or U14171 (N_14171,N_8082,N_9936);
or U14172 (N_14172,N_9034,N_11545);
nand U14173 (N_14173,N_11300,N_11416);
xor U14174 (N_14174,N_10654,N_9970);
or U14175 (N_14175,N_10901,N_10943);
xor U14176 (N_14176,N_11892,N_8682);
nor U14177 (N_14177,N_8717,N_10109);
and U14178 (N_14178,N_10352,N_10039);
or U14179 (N_14179,N_11002,N_9172);
or U14180 (N_14180,N_10381,N_11315);
nor U14181 (N_14181,N_10178,N_11301);
or U14182 (N_14182,N_10080,N_10259);
nand U14183 (N_14183,N_8831,N_11756);
nor U14184 (N_14184,N_9768,N_9174);
or U14185 (N_14185,N_9782,N_8747);
and U14186 (N_14186,N_10223,N_9981);
nor U14187 (N_14187,N_11973,N_10541);
and U14188 (N_14188,N_9211,N_10725);
nand U14189 (N_14189,N_11579,N_11336);
nand U14190 (N_14190,N_8773,N_8008);
nor U14191 (N_14191,N_8064,N_10913);
xor U14192 (N_14192,N_9245,N_10478);
xor U14193 (N_14193,N_9167,N_8719);
or U14194 (N_14194,N_11287,N_10796);
nor U14195 (N_14195,N_9633,N_10474);
nand U14196 (N_14196,N_10165,N_8541);
or U14197 (N_14197,N_11298,N_11860);
xor U14198 (N_14198,N_8890,N_11551);
or U14199 (N_14199,N_9784,N_11680);
xnor U14200 (N_14200,N_9694,N_8191);
nand U14201 (N_14201,N_9214,N_9226);
and U14202 (N_14202,N_11533,N_10015);
nor U14203 (N_14203,N_8531,N_8827);
nand U14204 (N_14204,N_11602,N_8289);
nor U14205 (N_14205,N_8615,N_8997);
and U14206 (N_14206,N_9975,N_11278);
nand U14207 (N_14207,N_10072,N_8686);
or U14208 (N_14208,N_10804,N_8967);
nor U14209 (N_14209,N_10213,N_11532);
xor U14210 (N_14210,N_8624,N_9850);
nand U14211 (N_14211,N_10908,N_11664);
nand U14212 (N_14212,N_11250,N_9895);
xor U14213 (N_14213,N_11636,N_11970);
xnor U14214 (N_14214,N_10692,N_10589);
nand U14215 (N_14215,N_8988,N_10969);
xnor U14216 (N_14216,N_11739,N_11920);
or U14217 (N_14217,N_11296,N_8415);
nand U14218 (N_14218,N_11794,N_8289);
or U14219 (N_14219,N_8502,N_11359);
nand U14220 (N_14220,N_8931,N_10044);
nor U14221 (N_14221,N_8370,N_9472);
or U14222 (N_14222,N_8099,N_10067);
nand U14223 (N_14223,N_11555,N_8061);
nor U14224 (N_14224,N_10762,N_11061);
nor U14225 (N_14225,N_10976,N_10066);
or U14226 (N_14226,N_10831,N_8841);
nand U14227 (N_14227,N_8526,N_9058);
nor U14228 (N_14228,N_11645,N_11982);
or U14229 (N_14229,N_9622,N_11802);
nor U14230 (N_14230,N_11600,N_11118);
nor U14231 (N_14231,N_11669,N_11267);
nor U14232 (N_14232,N_8027,N_10118);
nor U14233 (N_14233,N_11310,N_10271);
and U14234 (N_14234,N_10148,N_8307);
xnor U14235 (N_14235,N_8820,N_10304);
nor U14236 (N_14236,N_10583,N_8424);
nor U14237 (N_14237,N_11383,N_11582);
or U14238 (N_14238,N_10648,N_9948);
nand U14239 (N_14239,N_10380,N_9635);
or U14240 (N_14240,N_10277,N_10335);
xor U14241 (N_14241,N_10319,N_10465);
or U14242 (N_14242,N_11320,N_8875);
nor U14243 (N_14243,N_10813,N_11619);
and U14244 (N_14244,N_9884,N_9433);
xnor U14245 (N_14245,N_8161,N_11302);
nor U14246 (N_14246,N_10993,N_8837);
and U14247 (N_14247,N_8834,N_10748);
nor U14248 (N_14248,N_11351,N_9649);
xor U14249 (N_14249,N_11189,N_11088);
xnor U14250 (N_14250,N_8640,N_11592);
nand U14251 (N_14251,N_10935,N_10073);
and U14252 (N_14252,N_8705,N_8318);
xor U14253 (N_14253,N_9520,N_8751);
and U14254 (N_14254,N_10144,N_10853);
nand U14255 (N_14255,N_8012,N_11991);
or U14256 (N_14256,N_10063,N_8677);
or U14257 (N_14257,N_9550,N_11463);
xor U14258 (N_14258,N_10938,N_10258);
nand U14259 (N_14259,N_10357,N_11860);
nand U14260 (N_14260,N_8404,N_8443);
nor U14261 (N_14261,N_11711,N_10310);
or U14262 (N_14262,N_8262,N_10309);
xnor U14263 (N_14263,N_8645,N_10208);
and U14264 (N_14264,N_8802,N_10757);
and U14265 (N_14265,N_8661,N_8069);
nor U14266 (N_14266,N_11790,N_11857);
and U14267 (N_14267,N_10613,N_8497);
nand U14268 (N_14268,N_11731,N_10947);
nor U14269 (N_14269,N_9899,N_9355);
nor U14270 (N_14270,N_9699,N_11660);
nand U14271 (N_14271,N_8465,N_10857);
nand U14272 (N_14272,N_10386,N_11118);
xnor U14273 (N_14273,N_9138,N_8047);
xor U14274 (N_14274,N_10382,N_10678);
or U14275 (N_14275,N_11477,N_8042);
or U14276 (N_14276,N_10910,N_9850);
xnor U14277 (N_14277,N_10750,N_9600);
nor U14278 (N_14278,N_9963,N_10312);
or U14279 (N_14279,N_9377,N_8304);
or U14280 (N_14280,N_10734,N_10492);
nor U14281 (N_14281,N_11774,N_8596);
xnor U14282 (N_14282,N_8785,N_10005);
nor U14283 (N_14283,N_11419,N_9856);
nor U14284 (N_14284,N_10957,N_9666);
and U14285 (N_14285,N_9883,N_9914);
nor U14286 (N_14286,N_10151,N_9143);
nor U14287 (N_14287,N_10588,N_10431);
nand U14288 (N_14288,N_11180,N_9439);
nand U14289 (N_14289,N_9704,N_8174);
and U14290 (N_14290,N_10889,N_11751);
nor U14291 (N_14291,N_10291,N_11861);
or U14292 (N_14292,N_8783,N_8003);
and U14293 (N_14293,N_9275,N_8112);
or U14294 (N_14294,N_9924,N_11361);
xor U14295 (N_14295,N_10878,N_10813);
or U14296 (N_14296,N_10053,N_11057);
xnor U14297 (N_14297,N_9724,N_9161);
or U14298 (N_14298,N_9354,N_10376);
nor U14299 (N_14299,N_9637,N_10601);
and U14300 (N_14300,N_10590,N_9894);
or U14301 (N_14301,N_9620,N_9846);
or U14302 (N_14302,N_11500,N_8952);
nor U14303 (N_14303,N_11513,N_9933);
and U14304 (N_14304,N_11712,N_8867);
nand U14305 (N_14305,N_8385,N_9718);
and U14306 (N_14306,N_8251,N_10499);
xnor U14307 (N_14307,N_9891,N_9048);
and U14308 (N_14308,N_9278,N_11314);
xor U14309 (N_14309,N_9823,N_11491);
nor U14310 (N_14310,N_11062,N_9080);
nor U14311 (N_14311,N_11109,N_9532);
and U14312 (N_14312,N_9650,N_11356);
xnor U14313 (N_14313,N_9767,N_9196);
xor U14314 (N_14314,N_9175,N_11319);
xnor U14315 (N_14315,N_11270,N_9915);
nor U14316 (N_14316,N_10276,N_10898);
or U14317 (N_14317,N_10977,N_8176);
nor U14318 (N_14318,N_8465,N_10680);
nor U14319 (N_14319,N_9787,N_10290);
nor U14320 (N_14320,N_9442,N_9232);
or U14321 (N_14321,N_11848,N_11735);
nand U14322 (N_14322,N_9715,N_8640);
nor U14323 (N_14323,N_8384,N_11025);
nand U14324 (N_14324,N_9034,N_11179);
nand U14325 (N_14325,N_11473,N_8051);
or U14326 (N_14326,N_10547,N_9992);
and U14327 (N_14327,N_9364,N_8991);
or U14328 (N_14328,N_10654,N_11773);
xor U14329 (N_14329,N_8677,N_9523);
nand U14330 (N_14330,N_10809,N_8229);
nand U14331 (N_14331,N_10808,N_9509);
and U14332 (N_14332,N_11784,N_10371);
or U14333 (N_14333,N_9320,N_9909);
and U14334 (N_14334,N_8095,N_9698);
and U14335 (N_14335,N_8560,N_9908);
and U14336 (N_14336,N_9732,N_9149);
nand U14337 (N_14337,N_10484,N_8988);
xnor U14338 (N_14338,N_9576,N_8201);
and U14339 (N_14339,N_10681,N_8925);
nand U14340 (N_14340,N_8070,N_11040);
xor U14341 (N_14341,N_9036,N_11572);
nor U14342 (N_14342,N_11475,N_9200);
and U14343 (N_14343,N_10082,N_10877);
xor U14344 (N_14344,N_11807,N_9555);
xor U14345 (N_14345,N_9889,N_10824);
xnor U14346 (N_14346,N_11867,N_8637);
nor U14347 (N_14347,N_10587,N_9023);
nand U14348 (N_14348,N_9713,N_10222);
xnor U14349 (N_14349,N_11337,N_11761);
nand U14350 (N_14350,N_9998,N_10937);
nor U14351 (N_14351,N_11147,N_11623);
and U14352 (N_14352,N_10749,N_10581);
and U14353 (N_14353,N_8684,N_10449);
or U14354 (N_14354,N_10609,N_11616);
nor U14355 (N_14355,N_11959,N_8436);
xnor U14356 (N_14356,N_9661,N_10241);
nor U14357 (N_14357,N_10505,N_10221);
nor U14358 (N_14358,N_8292,N_11935);
xor U14359 (N_14359,N_10370,N_9759);
nor U14360 (N_14360,N_11086,N_9459);
and U14361 (N_14361,N_10743,N_11554);
nor U14362 (N_14362,N_10728,N_10348);
xor U14363 (N_14363,N_9555,N_11347);
nand U14364 (N_14364,N_9338,N_8596);
and U14365 (N_14365,N_11094,N_11837);
nor U14366 (N_14366,N_8611,N_11721);
and U14367 (N_14367,N_11839,N_9821);
nand U14368 (N_14368,N_10184,N_8478);
xnor U14369 (N_14369,N_8200,N_9652);
xor U14370 (N_14370,N_11639,N_10189);
xnor U14371 (N_14371,N_8404,N_8743);
and U14372 (N_14372,N_8542,N_9470);
and U14373 (N_14373,N_9957,N_9827);
nand U14374 (N_14374,N_8069,N_10787);
nand U14375 (N_14375,N_9771,N_9740);
nor U14376 (N_14376,N_10589,N_8752);
or U14377 (N_14377,N_11867,N_8404);
nand U14378 (N_14378,N_8444,N_10711);
nand U14379 (N_14379,N_10469,N_9363);
nand U14380 (N_14380,N_10514,N_9392);
xnor U14381 (N_14381,N_9165,N_9807);
nand U14382 (N_14382,N_11804,N_10626);
and U14383 (N_14383,N_11610,N_11936);
and U14384 (N_14384,N_8482,N_8518);
and U14385 (N_14385,N_11616,N_11505);
xor U14386 (N_14386,N_8543,N_8580);
and U14387 (N_14387,N_8427,N_9355);
xnor U14388 (N_14388,N_8168,N_10004);
nand U14389 (N_14389,N_10371,N_8381);
and U14390 (N_14390,N_9004,N_8547);
nor U14391 (N_14391,N_8661,N_10605);
xnor U14392 (N_14392,N_8123,N_10172);
nor U14393 (N_14393,N_9956,N_8689);
nor U14394 (N_14394,N_11177,N_11376);
and U14395 (N_14395,N_11450,N_8578);
nor U14396 (N_14396,N_10798,N_9948);
and U14397 (N_14397,N_8538,N_9367);
and U14398 (N_14398,N_11418,N_8451);
xor U14399 (N_14399,N_8299,N_11335);
xor U14400 (N_14400,N_10016,N_10046);
or U14401 (N_14401,N_11574,N_8535);
or U14402 (N_14402,N_8967,N_8358);
nand U14403 (N_14403,N_10933,N_9360);
xnor U14404 (N_14404,N_9781,N_10904);
and U14405 (N_14405,N_8881,N_10313);
and U14406 (N_14406,N_10858,N_11232);
nand U14407 (N_14407,N_11751,N_11389);
nand U14408 (N_14408,N_9679,N_11340);
nand U14409 (N_14409,N_11043,N_10787);
or U14410 (N_14410,N_10844,N_9301);
or U14411 (N_14411,N_11840,N_10369);
nor U14412 (N_14412,N_10456,N_10735);
xor U14413 (N_14413,N_10439,N_11638);
and U14414 (N_14414,N_8740,N_9029);
or U14415 (N_14415,N_11258,N_10369);
and U14416 (N_14416,N_9265,N_8001);
or U14417 (N_14417,N_11840,N_11835);
xnor U14418 (N_14418,N_10214,N_10047);
nand U14419 (N_14419,N_10606,N_10189);
nand U14420 (N_14420,N_8815,N_11894);
nor U14421 (N_14421,N_10375,N_8490);
or U14422 (N_14422,N_10270,N_8255);
nand U14423 (N_14423,N_8710,N_8835);
nor U14424 (N_14424,N_9767,N_9135);
or U14425 (N_14425,N_9056,N_10988);
xor U14426 (N_14426,N_8419,N_11900);
nor U14427 (N_14427,N_11748,N_11028);
or U14428 (N_14428,N_8019,N_9301);
nor U14429 (N_14429,N_10015,N_9102);
xor U14430 (N_14430,N_11321,N_10502);
or U14431 (N_14431,N_11751,N_9980);
xnor U14432 (N_14432,N_8307,N_8225);
nand U14433 (N_14433,N_10938,N_11766);
nand U14434 (N_14434,N_10734,N_9739);
nand U14435 (N_14435,N_10701,N_9979);
nor U14436 (N_14436,N_10346,N_8501);
nand U14437 (N_14437,N_11361,N_11914);
nand U14438 (N_14438,N_11141,N_11734);
and U14439 (N_14439,N_8525,N_8448);
nor U14440 (N_14440,N_8381,N_9888);
xor U14441 (N_14441,N_10043,N_8395);
nand U14442 (N_14442,N_10748,N_10523);
nand U14443 (N_14443,N_9871,N_9580);
nor U14444 (N_14444,N_11106,N_9140);
nand U14445 (N_14445,N_11391,N_11147);
or U14446 (N_14446,N_11225,N_9025);
nor U14447 (N_14447,N_10943,N_10823);
or U14448 (N_14448,N_9694,N_10094);
nor U14449 (N_14449,N_10821,N_8479);
and U14450 (N_14450,N_11861,N_8869);
xnor U14451 (N_14451,N_11261,N_10155);
and U14452 (N_14452,N_10631,N_11178);
nor U14453 (N_14453,N_9317,N_10560);
nor U14454 (N_14454,N_9231,N_8777);
and U14455 (N_14455,N_9622,N_11744);
xnor U14456 (N_14456,N_9108,N_10542);
nand U14457 (N_14457,N_9926,N_11923);
nor U14458 (N_14458,N_9583,N_10379);
and U14459 (N_14459,N_8810,N_10606);
nor U14460 (N_14460,N_10854,N_11344);
or U14461 (N_14461,N_11196,N_10375);
nor U14462 (N_14462,N_8682,N_11666);
and U14463 (N_14463,N_8087,N_11887);
or U14464 (N_14464,N_10206,N_9226);
or U14465 (N_14465,N_10881,N_9420);
and U14466 (N_14466,N_10659,N_10148);
or U14467 (N_14467,N_11011,N_10389);
nand U14468 (N_14468,N_8048,N_9667);
nand U14469 (N_14469,N_10014,N_9559);
or U14470 (N_14470,N_10541,N_10930);
or U14471 (N_14471,N_10467,N_9261);
nor U14472 (N_14472,N_8623,N_9443);
nand U14473 (N_14473,N_8635,N_11451);
or U14474 (N_14474,N_8588,N_9267);
nor U14475 (N_14475,N_11698,N_10848);
xor U14476 (N_14476,N_10957,N_8137);
nor U14477 (N_14477,N_11197,N_11818);
nor U14478 (N_14478,N_8057,N_11349);
nand U14479 (N_14479,N_10903,N_8513);
nand U14480 (N_14480,N_10237,N_11465);
nand U14481 (N_14481,N_9142,N_8784);
nand U14482 (N_14482,N_9812,N_10380);
and U14483 (N_14483,N_10794,N_11402);
nor U14484 (N_14484,N_8979,N_11934);
nor U14485 (N_14485,N_9675,N_10981);
nand U14486 (N_14486,N_8857,N_9034);
xor U14487 (N_14487,N_9917,N_11098);
nand U14488 (N_14488,N_9672,N_10257);
xnor U14489 (N_14489,N_8650,N_8353);
xnor U14490 (N_14490,N_8672,N_9592);
or U14491 (N_14491,N_10837,N_11740);
nand U14492 (N_14492,N_8775,N_8377);
xor U14493 (N_14493,N_9299,N_11955);
or U14494 (N_14494,N_8464,N_10910);
nor U14495 (N_14495,N_8673,N_8220);
nand U14496 (N_14496,N_10759,N_11075);
and U14497 (N_14497,N_8838,N_10896);
or U14498 (N_14498,N_8138,N_8402);
xnor U14499 (N_14499,N_10189,N_10502);
or U14500 (N_14500,N_11759,N_10879);
and U14501 (N_14501,N_10845,N_11022);
xor U14502 (N_14502,N_9369,N_8784);
xor U14503 (N_14503,N_10053,N_8994);
nand U14504 (N_14504,N_10818,N_11241);
and U14505 (N_14505,N_11751,N_10388);
and U14506 (N_14506,N_8618,N_10180);
nand U14507 (N_14507,N_10908,N_9334);
nor U14508 (N_14508,N_9657,N_9918);
nand U14509 (N_14509,N_9312,N_9113);
nand U14510 (N_14510,N_9216,N_10088);
nand U14511 (N_14511,N_9196,N_11311);
and U14512 (N_14512,N_9608,N_9655);
and U14513 (N_14513,N_8129,N_10444);
nor U14514 (N_14514,N_11122,N_10077);
nand U14515 (N_14515,N_10572,N_8754);
nand U14516 (N_14516,N_11075,N_10819);
nor U14517 (N_14517,N_9525,N_9554);
or U14518 (N_14518,N_9485,N_10168);
xnor U14519 (N_14519,N_8752,N_8392);
or U14520 (N_14520,N_11445,N_8292);
nor U14521 (N_14521,N_8123,N_10079);
nor U14522 (N_14522,N_9657,N_10593);
nand U14523 (N_14523,N_11557,N_8119);
nand U14524 (N_14524,N_10115,N_11901);
xnor U14525 (N_14525,N_8654,N_8906);
xor U14526 (N_14526,N_10279,N_11224);
xor U14527 (N_14527,N_9422,N_8018);
and U14528 (N_14528,N_9251,N_10551);
or U14529 (N_14529,N_10819,N_10161);
xor U14530 (N_14530,N_8280,N_11769);
nand U14531 (N_14531,N_10217,N_9148);
nand U14532 (N_14532,N_8604,N_11771);
nor U14533 (N_14533,N_10731,N_10298);
xnor U14534 (N_14534,N_10261,N_11696);
and U14535 (N_14535,N_9065,N_11456);
xnor U14536 (N_14536,N_9083,N_11278);
nand U14537 (N_14537,N_10948,N_8011);
nor U14538 (N_14538,N_9432,N_8840);
and U14539 (N_14539,N_10879,N_10932);
or U14540 (N_14540,N_8789,N_10958);
or U14541 (N_14541,N_11121,N_11468);
or U14542 (N_14542,N_8900,N_9287);
xor U14543 (N_14543,N_11047,N_9385);
xnor U14544 (N_14544,N_8398,N_10905);
or U14545 (N_14545,N_9742,N_11427);
and U14546 (N_14546,N_11076,N_10722);
nand U14547 (N_14547,N_9202,N_9655);
and U14548 (N_14548,N_8899,N_9858);
and U14549 (N_14549,N_8485,N_10359);
nor U14550 (N_14550,N_8933,N_10460);
or U14551 (N_14551,N_9794,N_8003);
nand U14552 (N_14552,N_8366,N_11781);
nor U14553 (N_14553,N_11327,N_11815);
xnor U14554 (N_14554,N_9377,N_11018);
xnor U14555 (N_14555,N_8411,N_8285);
and U14556 (N_14556,N_10163,N_8043);
nor U14557 (N_14557,N_10006,N_8550);
xnor U14558 (N_14558,N_9345,N_11088);
xnor U14559 (N_14559,N_11532,N_8359);
nor U14560 (N_14560,N_9109,N_9670);
nor U14561 (N_14561,N_11753,N_10588);
nor U14562 (N_14562,N_8230,N_9598);
or U14563 (N_14563,N_10188,N_10250);
nor U14564 (N_14564,N_11921,N_8529);
or U14565 (N_14565,N_8165,N_10523);
and U14566 (N_14566,N_9899,N_11839);
nor U14567 (N_14567,N_8626,N_9602);
nand U14568 (N_14568,N_11550,N_11376);
xnor U14569 (N_14569,N_11366,N_11357);
or U14570 (N_14570,N_10872,N_10450);
xnor U14571 (N_14571,N_10563,N_10807);
and U14572 (N_14572,N_10514,N_11784);
or U14573 (N_14573,N_8727,N_9997);
xnor U14574 (N_14574,N_8650,N_10645);
and U14575 (N_14575,N_10331,N_9485);
xnor U14576 (N_14576,N_11386,N_8581);
or U14577 (N_14577,N_11146,N_11433);
xor U14578 (N_14578,N_8682,N_9000);
and U14579 (N_14579,N_11823,N_11767);
nand U14580 (N_14580,N_10676,N_8352);
or U14581 (N_14581,N_10232,N_10298);
and U14582 (N_14582,N_11432,N_11753);
xnor U14583 (N_14583,N_9646,N_9128);
nand U14584 (N_14584,N_8110,N_10124);
nand U14585 (N_14585,N_10968,N_10399);
or U14586 (N_14586,N_9858,N_9164);
and U14587 (N_14587,N_11938,N_9604);
xnor U14588 (N_14588,N_9857,N_9802);
or U14589 (N_14589,N_8094,N_8954);
xor U14590 (N_14590,N_9026,N_11221);
nand U14591 (N_14591,N_9597,N_10606);
or U14592 (N_14592,N_9310,N_10908);
and U14593 (N_14593,N_8781,N_9496);
and U14594 (N_14594,N_10288,N_11107);
and U14595 (N_14595,N_11066,N_11806);
and U14596 (N_14596,N_9752,N_11793);
and U14597 (N_14597,N_11738,N_11325);
and U14598 (N_14598,N_10339,N_8968);
xor U14599 (N_14599,N_11868,N_8027);
nor U14600 (N_14600,N_11676,N_11898);
xnor U14601 (N_14601,N_10244,N_10425);
or U14602 (N_14602,N_10231,N_9001);
nand U14603 (N_14603,N_11547,N_11383);
and U14604 (N_14604,N_11138,N_9244);
or U14605 (N_14605,N_9788,N_9106);
xor U14606 (N_14606,N_11474,N_11762);
xor U14607 (N_14607,N_11993,N_11780);
and U14608 (N_14608,N_9377,N_11285);
nor U14609 (N_14609,N_11379,N_8326);
or U14610 (N_14610,N_8007,N_8874);
xor U14611 (N_14611,N_11581,N_9771);
and U14612 (N_14612,N_10837,N_10730);
xor U14613 (N_14613,N_9127,N_11440);
nand U14614 (N_14614,N_8128,N_9241);
nor U14615 (N_14615,N_11455,N_8746);
or U14616 (N_14616,N_8324,N_10066);
or U14617 (N_14617,N_8625,N_11065);
nor U14618 (N_14618,N_11657,N_10074);
nand U14619 (N_14619,N_11074,N_9455);
nor U14620 (N_14620,N_9036,N_8509);
and U14621 (N_14621,N_10599,N_11049);
xnor U14622 (N_14622,N_10551,N_9984);
and U14623 (N_14623,N_9581,N_8658);
and U14624 (N_14624,N_11454,N_10193);
xor U14625 (N_14625,N_10500,N_9215);
and U14626 (N_14626,N_11976,N_8546);
nand U14627 (N_14627,N_9074,N_9564);
nand U14628 (N_14628,N_10873,N_10550);
nor U14629 (N_14629,N_8350,N_9577);
and U14630 (N_14630,N_11399,N_10016);
nand U14631 (N_14631,N_8107,N_8164);
xnor U14632 (N_14632,N_8342,N_8813);
or U14633 (N_14633,N_9548,N_9710);
or U14634 (N_14634,N_10105,N_11477);
nor U14635 (N_14635,N_10003,N_8634);
and U14636 (N_14636,N_11511,N_8650);
and U14637 (N_14637,N_9983,N_8542);
or U14638 (N_14638,N_11615,N_8528);
or U14639 (N_14639,N_10123,N_11690);
or U14640 (N_14640,N_9866,N_9849);
nor U14641 (N_14641,N_8930,N_11309);
xor U14642 (N_14642,N_8442,N_11971);
and U14643 (N_14643,N_9837,N_9714);
and U14644 (N_14644,N_10767,N_8165);
xor U14645 (N_14645,N_9504,N_10441);
xnor U14646 (N_14646,N_8287,N_8139);
or U14647 (N_14647,N_8482,N_8189);
or U14648 (N_14648,N_10517,N_10589);
or U14649 (N_14649,N_9224,N_11802);
nor U14650 (N_14650,N_11549,N_9882);
and U14651 (N_14651,N_8006,N_10962);
or U14652 (N_14652,N_11207,N_8405);
and U14653 (N_14653,N_11474,N_11512);
or U14654 (N_14654,N_11876,N_11473);
nor U14655 (N_14655,N_8544,N_9513);
and U14656 (N_14656,N_8583,N_9577);
nand U14657 (N_14657,N_10314,N_8625);
nor U14658 (N_14658,N_11245,N_8848);
and U14659 (N_14659,N_8719,N_8771);
or U14660 (N_14660,N_10245,N_11854);
or U14661 (N_14661,N_11898,N_9539);
nand U14662 (N_14662,N_8747,N_10092);
xor U14663 (N_14663,N_10520,N_9343);
and U14664 (N_14664,N_9513,N_9831);
nor U14665 (N_14665,N_9181,N_8014);
xnor U14666 (N_14666,N_8610,N_11351);
or U14667 (N_14667,N_8068,N_8906);
nor U14668 (N_14668,N_9730,N_11422);
or U14669 (N_14669,N_9774,N_8869);
nor U14670 (N_14670,N_8996,N_9110);
nand U14671 (N_14671,N_9326,N_10855);
and U14672 (N_14672,N_11840,N_9027);
and U14673 (N_14673,N_11901,N_11940);
and U14674 (N_14674,N_10889,N_10737);
nor U14675 (N_14675,N_10518,N_11744);
or U14676 (N_14676,N_9629,N_10412);
nand U14677 (N_14677,N_11744,N_10576);
and U14678 (N_14678,N_10438,N_8802);
xor U14679 (N_14679,N_9361,N_10674);
and U14680 (N_14680,N_8577,N_8962);
and U14681 (N_14681,N_11327,N_9008);
and U14682 (N_14682,N_9882,N_10466);
or U14683 (N_14683,N_10471,N_8277);
and U14684 (N_14684,N_8678,N_9811);
nand U14685 (N_14685,N_11153,N_9512);
or U14686 (N_14686,N_9764,N_8207);
and U14687 (N_14687,N_9902,N_8145);
and U14688 (N_14688,N_9382,N_11054);
and U14689 (N_14689,N_9659,N_11330);
nor U14690 (N_14690,N_11393,N_10959);
xor U14691 (N_14691,N_11852,N_11796);
and U14692 (N_14692,N_8059,N_9495);
or U14693 (N_14693,N_10480,N_8516);
xor U14694 (N_14694,N_11040,N_10454);
xnor U14695 (N_14695,N_10780,N_11107);
and U14696 (N_14696,N_8213,N_8836);
or U14697 (N_14697,N_11007,N_9840);
xnor U14698 (N_14698,N_9241,N_8866);
or U14699 (N_14699,N_9419,N_9623);
xor U14700 (N_14700,N_8918,N_8009);
and U14701 (N_14701,N_8215,N_8323);
nor U14702 (N_14702,N_11702,N_11042);
xor U14703 (N_14703,N_10526,N_8022);
and U14704 (N_14704,N_9389,N_9965);
or U14705 (N_14705,N_11551,N_8954);
xor U14706 (N_14706,N_9513,N_10462);
or U14707 (N_14707,N_8499,N_9342);
xor U14708 (N_14708,N_8522,N_11079);
nand U14709 (N_14709,N_10924,N_9920);
xor U14710 (N_14710,N_9070,N_10561);
xnor U14711 (N_14711,N_9146,N_9449);
nand U14712 (N_14712,N_9273,N_9622);
and U14713 (N_14713,N_9838,N_10240);
or U14714 (N_14714,N_9477,N_8756);
or U14715 (N_14715,N_11721,N_11372);
xor U14716 (N_14716,N_11700,N_11104);
or U14717 (N_14717,N_10166,N_10027);
and U14718 (N_14718,N_9622,N_9255);
xnor U14719 (N_14719,N_10972,N_8905);
xnor U14720 (N_14720,N_9598,N_11181);
and U14721 (N_14721,N_9970,N_8628);
xnor U14722 (N_14722,N_8973,N_11153);
xnor U14723 (N_14723,N_9841,N_11860);
nand U14724 (N_14724,N_8330,N_9631);
nor U14725 (N_14725,N_8430,N_11697);
nand U14726 (N_14726,N_9709,N_10551);
xor U14727 (N_14727,N_11926,N_9615);
nand U14728 (N_14728,N_11204,N_11334);
and U14729 (N_14729,N_10970,N_10886);
nor U14730 (N_14730,N_11992,N_10671);
nand U14731 (N_14731,N_11208,N_11838);
or U14732 (N_14732,N_10392,N_10248);
and U14733 (N_14733,N_8176,N_9604);
or U14734 (N_14734,N_11233,N_10219);
nand U14735 (N_14735,N_8574,N_8060);
nor U14736 (N_14736,N_10071,N_8879);
nor U14737 (N_14737,N_8305,N_8956);
or U14738 (N_14738,N_10907,N_10183);
nor U14739 (N_14739,N_9280,N_9628);
nand U14740 (N_14740,N_8132,N_10630);
and U14741 (N_14741,N_11184,N_10888);
xor U14742 (N_14742,N_9336,N_11538);
or U14743 (N_14743,N_9870,N_8693);
or U14744 (N_14744,N_10734,N_10915);
nor U14745 (N_14745,N_10582,N_11707);
and U14746 (N_14746,N_8515,N_11435);
and U14747 (N_14747,N_9124,N_9795);
xor U14748 (N_14748,N_11634,N_11511);
nand U14749 (N_14749,N_8954,N_10115);
and U14750 (N_14750,N_8525,N_11763);
nor U14751 (N_14751,N_9193,N_10214);
nor U14752 (N_14752,N_10350,N_10931);
xnor U14753 (N_14753,N_11394,N_8312);
nand U14754 (N_14754,N_10962,N_11312);
xor U14755 (N_14755,N_8510,N_11868);
nand U14756 (N_14756,N_9673,N_9224);
nor U14757 (N_14757,N_10795,N_8087);
nand U14758 (N_14758,N_9684,N_11776);
and U14759 (N_14759,N_9494,N_11552);
nand U14760 (N_14760,N_11241,N_11767);
nor U14761 (N_14761,N_8019,N_10658);
and U14762 (N_14762,N_11343,N_10176);
or U14763 (N_14763,N_10184,N_9365);
or U14764 (N_14764,N_8349,N_9797);
xor U14765 (N_14765,N_11554,N_9404);
and U14766 (N_14766,N_8883,N_11331);
xnor U14767 (N_14767,N_8748,N_11787);
nor U14768 (N_14768,N_11975,N_9181);
nor U14769 (N_14769,N_8149,N_11728);
nor U14770 (N_14770,N_11242,N_9862);
nor U14771 (N_14771,N_11340,N_11680);
and U14772 (N_14772,N_8296,N_8624);
xor U14773 (N_14773,N_9447,N_9616);
nor U14774 (N_14774,N_8852,N_11966);
nand U14775 (N_14775,N_9955,N_9268);
and U14776 (N_14776,N_11233,N_10234);
and U14777 (N_14777,N_8114,N_8843);
nand U14778 (N_14778,N_11370,N_8400);
nand U14779 (N_14779,N_8597,N_11755);
nor U14780 (N_14780,N_9250,N_11951);
and U14781 (N_14781,N_11993,N_8693);
and U14782 (N_14782,N_10842,N_11898);
and U14783 (N_14783,N_9353,N_11121);
or U14784 (N_14784,N_9824,N_8820);
nor U14785 (N_14785,N_9107,N_8124);
or U14786 (N_14786,N_8773,N_10362);
nand U14787 (N_14787,N_10951,N_10401);
or U14788 (N_14788,N_9037,N_8872);
and U14789 (N_14789,N_8356,N_8228);
xor U14790 (N_14790,N_11861,N_9483);
and U14791 (N_14791,N_8724,N_9721);
nor U14792 (N_14792,N_9556,N_11123);
xnor U14793 (N_14793,N_8787,N_9728);
xnor U14794 (N_14794,N_9446,N_9061);
or U14795 (N_14795,N_10844,N_10451);
nor U14796 (N_14796,N_8671,N_8265);
nor U14797 (N_14797,N_11638,N_8796);
and U14798 (N_14798,N_8147,N_11064);
xnor U14799 (N_14799,N_9131,N_8585);
xnor U14800 (N_14800,N_11135,N_9019);
and U14801 (N_14801,N_8193,N_10833);
nor U14802 (N_14802,N_8585,N_9309);
or U14803 (N_14803,N_9313,N_10573);
xnor U14804 (N_14804,N_10725,N_9807);
or U14805 (N_14805,N_10598,N_11655);
xor U14806 (N_14806,N_10484,N_11404);
and U14807 (N_14807,N_9082,N_9371);
xnor U14808 (N_14808,N_10282,N_11539);
nand U14809 (N_14809,N_10706,N_10208);
nor U14810 (N_14810,N_11273,N_9109);
or U14811 (N_14811,N_10558,N_10471);
or U14812 (N_14812,N_11143,N_9219);
nand U14813 (N_14813,N_9072,N_11538);
and U14814 (N_14814,N_9834,N_8463);
nor U14815 (N_14815,N_9838,N_9026);
and U14816 (N_14816,N_11509,N_10903);
nor U14817 (N_14817,N_10161,N_11472);
or U14818 (N_14818,N_11410,N_9709);
and U14819 (N_14819,N_10754,N_11844);
and U14820 (N_14820,N_11187,N_10785);
nand U14821 (N_14821,N_9725,N_8221);
and U14822 (N_14822,N_10369,N_11290);
and U14823 (N_14823,N_9106,N_11064);
nand U14824 (N_14824,N_8774,N_9015);
nor U14825 (N_14825,N_8324,N_9613);
nor U14826 (N_14826,N_11685,N_10118);
nand U14827 (N_14827,N_11153,N_10788);
xor U14828 (N_14828,N_11144,N_9726);
and U14829 (N_14829,N_9830,N_10964);
nand U14830 (N_14830,N_11656,N_11147);
or U14831 (N_14831,N_11934,N_11424);
and U14832 (N_14832,N_11350,N_8812);
or U14833 (N_14833,N_11688,N_11234);
nor U14834 (N_14834,N_11444,N_8687);
or U14835 (N_14835,N_9838,N_8816);
or U14836 (N_14836,N_9813,N_9100);
or U14837 (N_14837,N_9643,N_11103);
or U14838 (N_14838,N_10442,N_9942);
or U14839 (N_14839,N_10265,N_9300);
xnor U14840 (N_14840,N_8415,N_10449);
and U14841 (N_14841,N_11568,N_9231);
nand U14842 (N_14842,N_9009,N_8886);
nand U14843 (N_14843,N_11208,N_10329);
xor U14844 (N_14844,N_11548,N_10221);
nand U14845 (N_14845,N_11734,N_10298);
or U14846 (N_14846,N_11397,N_9464);
xnor U14847 (N_14847,N_10943,N_9597);
or U14848 (N_14848,N_9705,N_8412);
xnor U14849 (N_14849,N_8366,N_8177);
nand U14850 (N_14850,N_11299,N_9233);
xor U14851 (N_14851,N_11189,N_11843);
nand U14852 (N_14852,N_9448,N_11430);
or U14853 (N_14853,N_10163,N_9762);
nor U14854 (N_14854,N_9557,N_11024);
xnor U14855 (N_14855,N_11888,N_11541);
nand U14856 (N_14856,N_8189,N_9910);
nand U14857 (N_14857,N_10419,N_11936);
or U14858 (N_14858,N_9400,N_10923);
nor U14859 (N_14859,N_8875,N_8529);
nand U14860 (N_14860,N_10435,N_9302);
nor U14861 (N_14861,N_9072,N_10221);
nor U14862 (N_14862,N_8507,N_8808);
and U14863 (N_14863,N_11705,N_8563);
and U14864 (N_14864,N_8321,N_11251);
nor U14865 (N_14865,N_11674,N_9500);
or U14866 (N_14866,N_9659,N_11753);
or U14867 (N_14867,N_11513,N_9390);
nor U14868 (N_14868,N_11824,N_8887);
and U14869 (N_14869,N_8379,N_10344);
nor U14870 (N_14870,N_8936,N_8264);
and U14871 (N_14871,N_8174,N_10554);
nor U14872 (N_14872,N_8527,N_10820);
and U14873 (N_14873,N_10733,N_10379);
nand U14874 (N_14874,N_11608,N_10619);
nand U14875 (N_14875,N_8095,N_8112);
xnor U14876 (N_14876,N_9070,N_11289);
and U14877 (N_14877,N_11861,N_8912);
nand U14878 (N_14878,N_9638,N_9586);
nor U14879 (N_14879,N_10739,N_11179);
and U14880 (N_14880,N_10559,N_8007);
xnor U14881 (N_14881,N_11028,N_11413);
or U14882 (N_14882,N_10588,N_9779);
xnor U14883 (N_14883,N_11394,N_11581);
xor U14884 (N_14884,N_9513,N_10889);
xnor U14885 (N_14885,N_10088,N_10994);
and U14886 (N_14886,N_9990,N_8915);
nor U14887 (N_14887,N_9714,N_10740);
xor U14888 (N_14888,N_11304,N_11951);
xnor U14889 (N_14889,N_9094,N_9755);
xor U14890 (N_14890,N_11869,N_11608);
nor U14891 (N_14891,N_10329,N_11386);
nor U14892 (N_14892,N_9658,N_8781);
nor U14893 (N_14893,N_9697,N_9372);
nor U14894 (N_14894,N_8212,N_10901);
or U14895 (N_14895,N_10266,N_10871);
xor U14896 (N_14896,N_11066,N_10131);
and U14897 (N_14897,N_10371,N_11778);
nand U14898 (N_14898,N_10536,N_8484);
xor U14899 (N_14899,N_10892,N_10953);
and U14900 (N_14900,N_11952,N_8333);
xnor U14901 (N_14901,N_10527,N_9326);
or U14902 (N_14902,N_9055,N_10776);
xor U14903 (N_14903,N_9435,N_11469);
nor U14904 (N_14904,N_11631,N_8810);
nand U14905 (N_14905,N_8164,N_10523);
nor U14906 (N_14906,N_8661,N_9161);
or U14907 (N_14907,N_10891,N_9288);
nand U14908 (N_14908,N_8007,N_10616);
xor U14909 (N_14909,N_8398,N_9553);
nor U14910 (N_14910,N_9131,N_9347);
nand U14911 (N_14911,N_10924,N_8390);
xor U14912 (N_14912,N_8708,N_11870);
or U14913 (N_14913,N_9516,N_11780);
or U14914 (N_14914,N_8947,N_9172);
and U14915 (N_14915,N_11313,N_8490);
and U14916 (N_14916,N_8701,N_8648);
or U14917 (N_14917,N_11708,N_8879);
nor U14918 (N_14918,N_11067,N_8728);
or U14919 (N_14919,N_10549,N_11237);
nand U14920 (N_14920,N_9148,N_9193);
or U14921 (N_14921,N_11145,N_9706);
and U14922 (N_14922,N_11465,N_11475);
or U14923 (N_14923,N_11339,N_10446);
xor U14924 (N_14924,N_11388,N_8581);
xor U14925 (N_14925,N_8278,N_9937);
nand U14926 (N_14926,N_11147,N_11364);
or U14927 (N_14927,N_11452,N_9880);
or U14928 (N_14928,N_11349,N_11886);
or U14929 (N_14929,N_10922,N_10479);
nand U14930 (N_14930,N_9944,N_11226);
and U14931 (N_14931,N_8840,N_11591);
xnor U14932 (N_14932,N_11047,N_11979);
xor U14933 (N_14933,N_8215,N_9392);
or U14934 (N_14934,N_10739,N_10947);
and U14935 (N_14935,N_11361,N_9843);
nand U14936 (N_14936,N_11091,N_8567);
nand U14937 (N_14937,N_8523,N_11450);
nor U14938 (N_14938,N_10468,N_11372);
or U14939 (N_14939,N_10493,N_10878);
nor U14940 (N_14940,N_11908,N_9497);
nor U14941 (N_14941,N_8865,N_8926);
or U14942 (N_14942,N_10390,N_8655);
nand U14943 (N_14943,N_8513,N_8320);
nand U14944 (N_14944,N_10085,N_8383);
and U14945 (N_14945,N_10114,N_8293);
nor U14946 (N_14946,N_11539,N_8078);
xnor U14947 (N_14947,N_11930,N_10121);
nor U14948 (N_14948,N_8480,N_9890);
nor U14949 (N_14949,N_11104,N_9453);
nor U14950 (N_14950,N_8636,N_9597);
or U14951 (N_14951,N_8861,N_10865);
xnor U14952 (N_14952,N_10538,N_10422);
nand U14953 (N_14953,N_8139,N_9981);
nand U14954 (N_14954,N_11054,N_8914);
and U14955 (N_14955,N_10938,N_9836);
or U14956 (N_14956,N_11615,N_11484);
xnor U14957 (N_14957,N_8480,N_11216);
and U14958 (N_14958,N_11790,N_10368);
nor U14959 (N_14959,N_8658,N_9730);
or U14960 (N_14960,N_9047,N_8912);
xor U14961 (N_14961,N_10146,N_10554);
nor U14962 (N_14962,N_9764,N_8476);
nand U14963 (N_14963,N_8076,N_11308);
and U14964 (N_14964,N_10383,N_10938);
nand U14965 (N_14965,N_11118,N_9081);
and U14966 (N_14966,N_9142,N_11116);
nand U14967 (N_14967,N_8662,N_10322);
or U14968 (N_14968,N_9779,N_10999);
xnor U14969 (N_14969,N_10819,N_9443);
nand U14970 (N_14970,N_11236,N_10765);
nor U14971 (N_14971,N_10140,N_9124);
nor U14972 (N_14972,N_9416,N_9792);
or U14973 (N_14973,N_10724,N_8316);
nand U14974 (N_14974,N_11317,N_8888);
nand U14975 (N_14975,N_10842,N_11104);
nand U14976 (N_14976,N_10021,N_11764);
or U14977 (N_14977,N_9853,N_8322);
nor U14978 (N_14978,N_11265,N_8077);
nor U14979 (N_14979,N_11930,N_9052);
nand U14980 (N_14980,N_9063,N_11412);
nand U14981 (N_14981,N_9529,N_9416);
nor U14982 (N_14982,N_8065,N_10544);
nor U14983 (N_14983,N_9340,N_10285);
xor U14984 (N_14984,N_9244,N_10090);
or U14985 (N_14985,N_10897,N_9689);
nand U14986 (N_14986,N_10585,N_9415);
nor U14987 (N_14987,N_9867,N_10733);
or U14988 (N_14988,N_11086,N_8039);
nor U14989 (N_14989,N_10640,N_9258);
nor U14990 (N_14990,N_9044,N_10339);
xnor U14991 (N_14991,N_8962,N_8158);
nand U14992 (N_14992,N_10323,N_10863);
xnor U14993 (N_14993,N_11968,N_10037);
nor U14994 (N_14994,N_9128,N_10094);
xnor U14995 (N_14995,N_8014,N_10949);
nor U14996 (N_14996,N_10316,N_8325);
xnor U14997 (N_14997,N_11308,N_8888);
nor U14998 (N_14998,N_10946,N_10693);
nand U14999 (N_14999,N_9062,N_11273);
nand U15000 (N_15000,N_11622,N_9607);
nor U15001 (N_15001,N_11604,N_10513);
xnor U15002 (N_15002,N_8600,N_8143);
nor U15003 (N_15003,N_10336,N_10225);
or U15004 (N_15004,N_11054,N_10300);
nand U15005 (N_15005,N_11769,N_9695);
and U15006 (N_15006,N_9873,N_11367);
or U15007 (N_15007,N_9799,N_9249);
xor U15008 (N_15008,N_9227,N_8732);
xor U15009 (N_15009,N_10864,N_9151);
nand U15010 (N_15010,N_9929,N_8882);
and U15011 (N_15011,N_10299,N_11539);
nor U15012 (N_15012,N_11965,N_8884);
nor U15013 (N_15013,N_11806,N_10427);
nor U15014 (N_15014,N_9164,N_10431);
nand U15015 (N_15015,N_10373,N_9565);
and U15016 (N_15016,N_8531,N_11232);
xor U15017 (N_15017,N_8641,N_9696);
xnor U15018 (N_15018,N_9476,N_11023);
nand U15019 (N_15019,N_9799,N_11996);
or U15020 (N_15020,N_11671,N_10086);
and U15021 (N_15021,N_10763,N_8076);
nand U15022 (N_15022,N_10535,N_11106);
or U15023 (N_15023,N_11220,N_11059);
xor U15024 (N_15024,N_10894,N_9102);
nand U15025 (N_15025,N_9178,N_8258);
or U15026 (N_15026,N_11752,N_11553);
or U15027 (N_15027,N_8219,N_8894);
and U15028 (N_15028,N_11754,N_11664);
xnor U15029 (N_15029,N_11134,N_8193);
or U15030 (N_15030,N_11541,N_11240);
and U15031 (N_15031,N_8657,N_11792);
or U15032 (N_15032,N_10930,N_9135);
and U15033 (N_15033,N_8891,N_11560);
or U15034 (N_15034,N_11978,N_8215);
nor U15035 (N_15035,N_8408,N_10857);
xnor U15036 (N_15036,N_9750,N_9633);
nor U15037 (N_15037,N_11178,N_8508);
xnor U15038 (N_15038,N_8299,N_11920);
nand U15039 (N_15039,N_11381,N_9034);
xor U15040 (N_15040,N_11180,N_9048);
nand U15041 (N_15041,N_9798,N_10037);
or U15042 (N_15042,N_11808,N_9556);
nand U15043 (N_15043,N_11207,N_9322);
nor U15044 (N_15044,N_10639,N_10556);
xnor U15045 (N_15045,N_8208,N_8092);
nor U15046 (N_15046,N_8642,N_8014);
nand U15047 (N_15047,N_11189,N_9544);
nor U15048 (N_15048,N_9716,N_10799);
or U15049 (N_15049,N_8049,N_10352);
nor U15050 (N_15050,N_8421,N_11222);
nor U15051 (N_15051,N_8457,N_8981);
xnor U15052 (N_15052,N_10962,N_11341);
nor U15053 (N_15053,N_8364,N_10960);
nor U15054 (N_15054,N_8638,N_8827);
and U15055 (N_15055,N_11690,N_8429);
nand U15056 (N_15056,N_8575,N_9428);
xnor U15057 (N_15057,N_9061,N_10006);
and U15058 (N_15058,N_10692,N_9016);
nor U15059 (N_15059,N_9415,N_10403);
and U15060 (N_15060,N_11587,N_10879);
nor U15061 (N_15061,N_9993,N_9623);
nand U15062 (N_15062,N_10628,N_9092);
and U15063 (N_15063,N_9242,N_8925);
xor U15064 (N_15064,N_11102,N_10916);
nand U15065 (N_15065,N_9070,N_8927);
xnor U15066 (N_15066,N_10193,N_8598);
xor U15067 (N_15067,N_8656,N_10362);
nand U15068 (N_15068,N_9144,N_8523);
and U15069 (N_15069,N_9667,N_10914);
xnor U15070 (N_15070,N_11231,N_11065);
nor U15071 (N_15071,N_11435,N_8234);
nor U15072 (N_15072,N_9160,N_8852);
nand U15073 (N_15073,N_9463,N_8468);
xor U15074 (N_15074,N_11176,N_10957);
nor U15075 (N_15075,N_11238,N_8606);
nand U15076 (N_15076,N_10735,N_10872);
nor U15077 (N_15077,N_11727,N_8892);
xor U15078 (N_15078,N_10766,N_11127);
nor U15079 (N_15079,N_8997,N_10194);
xnor U15080 (N_15080,N_9061,N_10420);
or U15081 (N_15081,N_8303,N_8269);
nand U15082 (N_15082,N_11574,N_11236);
and U15083 (N_15083,N_8775,N_10787);
or U15084 (N_15084,N_11305,N_11376);
or U15085 (N_15085,N_10906,N_8312);
xor U15086 (N_15086,N_11213,N_10941);
and U15087 (N_15087,N_9175,N_10201);
and U15088 (N_15088,N_8664,N_11637);
xnor U15089 (N_15089,N_11326,N_9516);
and U15090 (N_15090,N_10463,N_8705);
xor U15091 (N_15091,N_9444,N_10438);
xnor U15092 (N_15092,N_8582,N_10582);
and U15093 (N_15093,N_10493,N_9714);
xnor U15094 (N_15094,N_9304,N_8966);
nand U15095 (N_15095,N_9473,N_9054);
or U15096 (N_15096,N_9141,N_9889);
xnor U15097 (N_15097,N_8165,N_10892);
nand U15098 (N_15098,N_9247,N_10448);
and U15099 (N_15099,N_10298,N_11367);
xor U15100 (N_15100,N_10714,N_8794);
nand U15101 (N_15101,N_9404,N_9894);
nor U15102 (N_15102,N_11997,N_10518);
nor U15103 (N_15103,N_9794,N_11726);
or U15104 (N_15104,N_8127,N_11679);
nand U15105 (N_15105,N_9857,N_11827);
nor U15106 (N_15106,N_9386,N_9394);
and U15107 (N_15107,N_10243,N_10172);
and U15108 (N_15108,N_10752,N_9630);
nand U15109 (N_15109,N_8219,N_11319);
and U15110 (N_15110,N_10463,N_11847);
nand U15111 (N_15111,N_10125,N_9298);
and U15112 (N_15112,N_8524,N_10674);
xnor U15113 (N_15113,N_8099,N_10318);
or U15114 (N_15114,N_10194,N_10129);
nor U15115 (N_15115,N_9543,N_11523);
and U15116 (N_15116,N_9867,N_10870);
nand U15117 (N_15117,N_10221,N_11343);
and U15118 (N_15118,N_9757,N_11137);
nand U15119 (N_15119,N_11280,N_9741);
nor U15120 (N_15120,N_10587,N_8990);
nand U15121 (N_15121,N_8010,N_9945);
and U15122 (N_15122,N_8338,N_11037);
nand U15123 (N_15123,N_11065,N_10393);
and U15124 (N_15124,N_9628,N_10098);
xnor U15125 (N_15125,N_11362,N_11842);
nor U15126 (N_15126,N_8882,N_11586);
nand U15127 (N_15127,N_11569,N_8206);
xor U15128 (N_15128,N_11292,N_9008);
xnor U15129 (N_15129,N_11496,N_9524);
nand U15130 (N_15130,N_10810,N_10759);
nand U15131 (N_15131,N_10348,N_9864);
and U15132 (N_15132,N_11258,N_11901);
and U15133 (N_15133,N_9693,N_11499);
and U15134 (N_15134,N_8202,N_10514);
nor U15135 (N_15135,N_11744,N_8790);
nor U15136 (N_15136,N_9351,N_10106);
xor U15137 (N_15137,N_9226,N_8064);
and U15138 (N_15138,N_11680,N_10160);
or U15139 (N_15139,N_11620,N_9464);
nand U15140 (N_15140,N_8726,N_11371);
and U15141 (N_15141,N_11428,N_9172);
or U15142 (N_15142,N_11694,N_11731);
or U15143 (N_15143,N_10351,N_9667);
nand U15144 (N_15144,N_10620,N_9786);
or U15145 (N_15145,N_11257,N_11686);
and U15146 (N_15146,N_8921,N_8430);
nor U15147 (N_15147,N_11041,N_11009);
nand U15148 (N_15148,N_8091,N_9745);
nor U15149 (N_15149,N_11949,N_10100);
xnor U15150 (N_15150,N_10132,N_8438);
and U15151 (N_15151,N_9825,N_8612);
nand U15152 (N_15152,N_11487,N_8059);
nand U15153 (N_15153,N_10103,N_8513);
and U15154 (N_15154,N_11066,N_8042);
and U15155 (N_15155,N_10210,N_9145);
nor U15156 (N_15156,N_10240,N_10322);
nor U15157 (N_15157,N_11653,N_8539);
xnor U15158 (N_15158,N_11550,N_11414);
nand U15159 (N_15159,N_10085,N_11015);
or U15160 (N_15160,N_8943,N_8435);
or U15161 (N_15161,N_9847,N_8657);
or U15162 (N_15162,N_8348,N_11025);
or U15163 (N_15163,N_8858,N_8459);
nor U15164 (N_15164,N_10627,N_9272);
nor U15165 (N_15165,N_11782,N_10976);
nand U15166 (N_15166,N_9316,N_9143);
xnor U15167 (N_15167,N_9804,N_11469);
and U15168 (N_15168,N_10745,N_8318);
and U15169 (N_15169,N_11471,N_9257);
or U15170 (N_15170,N_8037,N_11606);
or U15171 (N_15171,N_11607,N_11274);
xnor U15172 (N_15172,N_10324,N_11888);
or U15173 (N_15173,N_11147,N_9107);
and U15174 (N_15174,N_11784,N_10887);
or U15175 (N_15175,N_9438,N_8501);
and U15176 (N_15176,N_8107,N_8724);
xnor U15177 (N_15177,N_9402,N_9194);
and U15178 (N_15178,N_10953,N_10825);
nor U15179 (N_15179,N_9499,N_8104);
xnor U15180 (N_15180,N_10691,N_8205);
nor U15181 (N_15181,N_11994,N_8840);
nand U15182 (N_15182,N_11935,N_11930);
nor U15183 (N_15183,N_9299,N_10963);
nor U15184 (N_15184,N_11454,N_10423);
nand U15185 (N_15185,N_8050,N_9470);
nor U15186 (N_15186,N_8061,N_11512);
or U15187 (N_15187,N_9002,N_9399);
xor U15188 (N_15188,N_9146,N_10527);
nand U15189 (N_15189,N_9145,N_10753);
nor U15190 (N_15190,N_11340,N_8459);
and U15191 (N_15191,N_11092,N_9215);
nand U15192 (N_15192,N_8977,N_11270);
and U15193 (N_15193,N_8196,N_9094);
xor U15194 (N_15194,N_11120,N_10192);
and U15195 (N_15195,N_9382,N_11890);
nand U15196 (N_15196,N_8876,N_8071);
and U15197 (N_15197,N_11282,N_8398);
and U15198 (N_15198,N_10957,N_10387);
and U15199 (N_15199,N_11536,N_11670);
and U15200 (N_15200,N_11249,N_9072);
xor U15201 (N_15201,N_8486,N_10933);
or U15202 (N_15202,N_10709,N_10941);
nor U15203 (N_15203,N_9002,N_10722);
or U15204 (N_15204,N_10064,N_10603);
or U15205 (N_15205,N_11213,N_10406);
nor U15206 (N_15206,N_11833,N_8525);
nor U15207 (N_15207,N_10400,N_10079);
and U15208 (N_15208,N_10155,N_8038);
nor U15209 (N_15209,N_10260,N_11684);
nand U15210 (N_15210,N_11230,N_10327);
xor U15211 (N_15211,N_10540,N_10906);
or U15212 (N_15212,N_11808,N_9435);
xnor U15213 (N_15213,N_8062,N_9762);
and U15214 (N_15214,N_8725,N_9492);
or U15215 (N_15215,N_10704,N_11188);
nor U15216 (N_15216,N_8726,N_10396);
and U15217 (N_15217,N_8118,N_9319);
nor U15218 (N_15218,N_8021,N_11763);
nor U15219 (N_15219,N_8787,N_9386);
nor U15220 (N_15220,N_8053,N_8409);
and U15221 (N_15221,N_8839,N_9410);
nand U15222 (N_15222,N_10120,N_10242);
nand U15223 (N_15223,N_10344,N_8336);
or U15224 (N_15224,N_11419,N_9413);
nand U15225 (N_15225,N_10750,N_8497);
or U15226 (N_15226,N_8629,N_8015);
nand U15227 (N_15227,N_11055,N_8372);
or U15228 (N_15228,N_9964,N_11829);
nor U15229 (N_15229,N_8037,N_8936);
and U15230 (N_15230,N_8551,N_10169);
nand U15231 (N_15231,N_10458,N_9542);
nor U15232 (N_15232,N_10046,N_10577);
nor U15233 (N_15233,N_8038,N_10098);
or U15234 (N_15234,N_9792,N_11411);
nand U15235 (N_15235,N_11458,N_8250);
nand U15236 (N_15236,N_9817,N_8070);
nor U15237 (N_15237,N_10920,N_8600);
and U15238 (N_15238,N_8989,N_11639);
nand U15239 (N_15239,N_11043,N_10316);
xor U15240 (N_15240,N_10664,N_11826);
nand U15241 (N_15241,N_8859,N_11598);
xor U15242 (N_15242,N_11708,N_9823);
nand U15243 (N_15243,N_8294,N_9911);
nand U15244 (N_15244,N_10814,N_11672);
xor U15245 (N_15245,N_10962,N_8299);
xnor U15246 (N_15246,N_8316,N_8581);
nor U15247 (N_15247,N_11033,N_8177);
and U15248 (N_15248,N_11096,N_10218);
and U15249 (N_15249,N_11816,N_9664);
nor U15250 (N_15250,N_8132,N_11278);
nor U15251 (N_15251,N_8479,N_10042);
nand U15252 (N_15252,N_8464,N_8419);
nor U15253 (N_15253,N_11232,N_11854);
and U15254 (N_15254,N_11662,N_10162);
and U15255 (N_15255,N_10594,N_11651);
nand U15256 (N_15256,N_8167,N_9130);
and U15257 (N_15257,N_10357,N_11592);
and U15258 (N_15258,N_9753,N_9826);
nand U15259 (N_15259,N_9392,N_8034);
and U15260 (N_15260,N_11006,N_10240);
nor U15261 (N_15261,N_8089,N_9948);
and U15262 (N_15262,N_11552,N_9350);
and U15263 (N_15263,N_8189,N_8725);
xnor U15264 (N_15264,N_9153,N_10028);
or U15265 (N_15265,N_10531,N_11119);
and U15266 (N_15266,N_8774,N_11102);
nand U15267 (N_15267,N_9036,N_8550);
xor U15268 (N_15268,N_10453,N_8051);
xor U15269 (N_15269,N_8042,N_8681);
or U15270 (N_15270,N_9334,N_9030);
nor U15271 (N_15271,N_11665,N_10626);
nand U15272 (N_15272,N_8454,N_10684);
or U15273 (N_15273,N_8044,N_10058);
xor U15274 (N_15274,N_8802,N_10279);
xnor U15275 (N_15275,N_10226,N_9179);
nand U15276 (N_15276,N_10195,N_9902);
nor U15277 (N_15277,N_10383,N_10496);
or U15278 (N_15278,N_10226,N_8072);
or U15279 (N_15279,N_9236,N_8573);
or U15280 (N_15280,N_9046,N_9454);
and U15281 (N_15281,N_9711,N_11855);
or U15282 (N_15282,N_10284,N_10589);
xnor U15283 (N_15283,N_9767,N_9478);
xor U15284 (N_15284,N_8026,N_11571);
nor U15285 (N_15285,N_9884,N_11720);
and U15286 (N_15286,N_9068,N_10529);
or U15287 (N_15287,N_8433,N_10018);
nand U15288 (N_15288,N_8934,N_10927);
or U15289 (N_15289,N_9060,N_9985);
or U15290 (N_15290,N_8576,N_10074);
and U15291 (N_15291,N_10893,N_8466);
xnor U15292 (N_15292,N_9699,N_9569);
and U15293 (N_15293,N_10669,N_9146);
xnor U15294 (N_15294,N_9310,N_10386);
or U15295 (N_15295,N_10593,N_9640);
xor U15296 (N_15296,N_9714,N_8585);
nor U15297 (N_15297,N_9934,N_8685);
nor U15298 (N_15298,N_11114,N_11768);
xor U15299 (N_15299,N_11899,N_8953);
nor U15300 (N_15300,N_11894,N_11358);
xor U15301 (N_15301,N_8271,N_11545);
nand U15302 (N_15302,N_8122,N_8919);
or U15303 (N_15303,N_10654,N_11960);
and U15304 (N_15304,N_9613,N_10609);
nand U15305 (N_15305,N_9126,N_10889);
and U15306 (N_15306,N_10251,N_8115);
and U15307 (N_15307,N_9429,N_11732);
xnor U15308 (N_15308,N_10870,N_10465);
or U15309 (N_15309,N_9256,N_11573);
and U15310 (N_15310,N_8816,N_11196);
xnor U15311 (N_15311,N_8958,N_11380);
nand U15312 (N_15312,N_8865,N_11720);
nand U15313 (N_15313,N_9921,N_10826);
and U15314 (N_15314,N_9314,N_10879);
nor U15315 (N_15315,N_11755,N_11011);
and U15316 (N_15316,N_10568,N_8154);
or U15317 (N_15317,N_10509,N_10244);
nor U15318 (N_15318,N_11892,N_10896);
or U15319 (N_15319,N_8995,N_10856);
or U15320 (N_15320,N_9414,N_9618);
xnor U15321 (N_15321,N_11495,N_9236);
xor U15322 (N_15322,N_11617,N_8513);
nand U15323 (N_15323,N_11361,N_9617);
nor U15324 (N_15324,N_9174,N_10238);
xnor U15325 (N_15325,N_9045,N_10957);
nand U15326 (N_15326,N_9827,N_9078);
xnor U15327 (N_15327,N_11842,N_8690);
nand U15328 (N_15328,N_11080,N_11807);
nor U15329 (N_15329,N_11211,N_11185);
or U15330 (N_15330,N_8902,N_9648);
or U15331 (N_15331,N_9413,N_8497);
xor U15332 (N_15332,N_10925,N_9951);
and U15333 (N_15333,N_8287,N_9034);
or U15334 (N_15334,N_11923,N_10043);
and U15335 (N_15335,N_10942,N_11535);
xor U15336 (N_15336,N_10561,N_10816);
and U15337 (N_15337,N_10953,N_9336);
and U15338 (N_15338,N_8182,N_8705);
nor U15339 (N_15339,N_8260,N_11569);
nor U15340 (N_15340,N_8011,N_9560);
or U15341 (N_15341,N_11255,N_9607);
or U15342 (N_15342,N_10818,N_10436);
xnor U15343 (N_15343,N_9249,N_10038);
nor U15344 (N_15344,N_11623,N_11324);
or U15345 (N_15345,N_11323,N_9211);
or U15346 (N_15346,N_8241,N_9973);
or U15347 (N_15347,N_11131,N_11626);
or U15348 (N_15348,N_10559,N_9104);
or U15349 (N_15349,N_11459,N_9566);
nor U15350 (N_15350,N_9943,N_8369);
and U15351 (N_15351,N_8234,N_10864);
nor U15352 (N_15352,N_8793,N_9730);
and U15353 (N_15353,N_10055,N_11520);
nor U15354 (N_15354,N_10121,N_8511);
and U15355 (N_15355,N_9099,N_9715);
nand U15356 (N_15356,N_8004,N_9533);
or U15357 (N_15357,N_11538,N_11012);
nor U15358 (N_15358,N_10623,N_11427);
xnor U15359 (N_15359,N_10123,N_11192);
xnor U15360 (N_15360,N_9638,N_11192);
and U15361 (N_15361,N_9860,N_11475);
and U15362 (N_15362,N_10506,N_11601);
and U15363 (N_15363,N_11943,N_11150);
nor U15364 (N_15364,N_10530,N_9518);
nand U15365 (N_15365,N_11686,N_10848);
xnor U15366 (N_15366,N_8534,N_9427);
or U15367 (N_15367,N_9717,N_9904);
and U15368 (N_15368,N_10116,N_11553);
and U15369 (N_15369,N_11380,N_9365);
xnor U15370 (N_15370,N_11387,N_8537);
nand U15371 (N_15371,N_9435,N_11361);
nor U15372 (N_15372,N_9842,N_8459);
xnor U15373 (N_15373,N_10844,N_10426);
xor U15374 (N_15374,N_8532,N_8275);
nand U15375 (N_15375,N_9354,N_9625);
or U15376 (N_15376,N_8834,N_9766);
xnor U15377 (N_15377,N_10993,N_9681);
nand U15378 (N_15378,N_10714,N_9089);
nor U15379 (N_15379,N_8965,N_8495);
xnor U15380 (N_15380,N_8297,N_11850);
or U15381 (N_15381,N_11810,N_9874);
or U15382 (N_15382,N_8671,N_10419);
xnor U15383 (N_15383,N_8303,N_9599);
xor U15384 (N_15384,N_8784,N_9917);
xor U15385 (N_15385,N_9483,N_10517);
xor U15386 (N_15386,N_10831,N_10851);
or U15387 (N_15387,N_10273,N_10479);
nand U15388 (N_15388,N_9029,N_9859);
nor U15389 (N_15389,N_10033,N_11205);
and U15390 (N_15390,N_8883,N_11976);
xnor U15391 (N_15391,N_8497,N_8513);
or U15392 (N_15392,N_10242,N_11278);
nor U15393 (N_15393,N_10915,N_8179);
nor U15394 (N_15394,N_10144,N_8533);
nand U15395 (N_15395,N_8744,N_10842);
and U15396 (N_15396,N_11208,N_9508);
xor U15397 (N_15397,N_10241,N_10275);
and U15398 (N_15398,N_10521,N_10800);
xor U15399 (N_15399,N_9575,N_11834);
nor U15400 (N_15400,N_10927,N_8948);
or U15401 (N_15401,N_11099,N_11444);
nand U15402 (N_15402,N_9896,N_11422);
nand U15403 (N_15403,N_9639,N_9536);
xnor U15404 (N_15404,N_9687,N_11682);
nor U15405 (N_15405,N_10495,N_9572);
or U15406 (N_15406,N_11404,N_11599);
nor U15407 (N_15407,N_9348,N_9904);
xnor U15408 (N_15408,N_9108,N_10807);
xnor U15409 (N_15409,N_11935,N_11937);
or U15410 (N_15410,N_8032,N_11198);
or U15411 (N_15411,N_11949,N_11643);
nand U15412 (N_15412,N_9819,N_9731);
or U15413 (N_15413,N_8233,N_9022);
xor U15414 (N_15414,N_11348,N_9981);
and U15415 (N_15415,N_8223,N_11263);
or U15416 (N_15416,N_10246,N_10697);
or U15417 (N_15417,N_10379,N_10940);
nor U15418 (N_15418,N_10722,N_9220);
and U15419 (N_15419,N_10971,N_11963);
or U15420 (N_15420,N_8562,N_9236);
or U15421 (N_15421,N_9869,N_10471);
nor U15422 (N_15422,N_8506,N_9238);
or U15423 (N_15423,N_10886,N_10829);
and U15424 (N_15424,N_10592,N_8069);
nor U15425 (N_15425,N_8200,N_9461);
nor U15426 (N_15426,N_10147,N_9321);
nor U15427 (N_15427,N_11469,N_9810);
nor U15428 (N_15428,N_11929,N_8143);
and U15429 (N_15429,N_9818,N_8089);
nand U15430 (N_15430,N_11150,N_10123);
or U15431 (N_15431,N_11510,N_9986);
and U15432 (N_15432,N_8342,N_11790);
nor U15433 (N_15433,N_11846,N_8217);
nor U15434 (N_15434,N_11286,N_8569);
and U15435 (N_15435,N_9756,N_11696);
nand U15436 (N_15436,N_8400,N_10455);
and U15437 (N_15437,N_10156,N_11859);
nand U15438 (N_15438,N_10918,N_8500);
xnor U15439 (N_15439,N_9492,N_8896);
nor U15440 (N_15440,N_11627,N_9298);
nand U15441 (N_15441,N_8699,N_11499);
nor U15442 (N_15442,N_11568,N_9296);
or U15443 (N_15443,N_9085,N_11799);
or U15444 (N_15444,N_9367,N_9906);
xnor U15445 (N_15445,N_11152,N_11030);
nand U15446 (N_15446,N_8722,N_9109);
xor U15447 (N_15447,N_11377,N_9088);
and U15448 (N_15448,N_11588,N_11438);
nand U15449 (N_15449,N_8080,N_8809);
nand U15450 (N_15450,N_10959,N_11749);
nand U15451 (N_15451,N_9318,N_9228);
xor U15452 (N_15452,N_8777,N_10001);
or U15453 (N_15453,N_9724,N_10755);
nand U15454 (N_15454,N_9176,N_10673);
and U15455 (N_15455,N_11259,N_9941);
nand U15456 (N_15456,N_8667,N_9099);
xnor U15457 (N_15457,N_10605,N_11979);
or U15458 (N_15458,N_10630,N_9099);
xnor U15459 (N_15459,N_10592,N_10542);
or U15460 (N_15460,N_8497,N_9796);
or U15461 (N_15461,N_8348,N_11584);
nand U15462 (N_15462,N_9041,N_11990);
or U15463 (N_15463,N_11907,N_10730);
nor U15464 (N_15464,N_9324,N_10257);
xnor U15465 (N_15465,N_9842,N_10275);
or U15466 (N_15466,N_11149,N_11957);
nor U15467 (N_15467,N_8903,N_10692);
xor U15468 (N_15468,N_11651,N_9431);
nand U15469 (N_15469,N_10965,N_10305);
nand U15470 (N_15470,N_8052,N_8071);
nor U15471 (N_15471,N_8599,N_10292);
and U15472 (N_15472,N_10110,N_11504);
or U15473 (N_15473,N_8399,N_8831);
nand U15474 (N_15474,N_10015,N_10616);
nand U15475 (N_15475,N_11877,N_9940);
xor U15476 (N_15476,N_10895,N_11150);
or U15477 (N_15477,N_9268,N_11114);
nor U15478 (N_15478,N_8934,N_8462);
xor U15479 (N_15479,N_10699,N_8742);
or U15480 (N_15480,N_11037,N_11478);
and U15481 (N_15481,N_9665,N_11619);
nor U15482 (N_15482,N_10573,N_10626);
and U15483 (N_15483,N_10597,N_9142);
or U15484 (N_15484,N_11239,N_11391);
nor U15485 (N_15485,N_8893,N_8712);
or U15486 (N_15486,N_8867,N_11476);
or U15487 (N_15487,N_8063,N_11023);
nand U15488 (N_15488,N_9695,N_9521);
and U15489 (N_15489,N_11543,N_10714);
nor U15490 (N_15490,N_11749,N_11888);
xor U15491 (N_15491,N_9621,N_8453);
or U15492 (N_15492,N_10699,N_10008);
or U15493 (N_15493,N_11428,N_11710);
and U15494 (N_15494,N_11861,N_10701);
nand U15495 (N_15495,N_8392,N_9840);
nor U15496 (N_15496,N_10202,N_11683);
and U15497 (N_15497,N_9494,N_9557);
and U15498 (N_15498,N_8228,N_10096);
xnor U15499 (N_15499,N_10086,N_8201);
or U15500 (N_15500,N_8142,N_10851);
xnor U15501 (N_15501,N_9162,N_9936);
and U15502 (N_15502,N_11206,N_9055);
xnor U15503 (N_15503,N_10563,N_8139);
or U15504 (N_15504,N_11248,N_11482);
and U15505 (N_15505,N_8447,N_10300);
and U15506 (N_15506,N_8021,N_9044);
xnor U15507 (N_15507,N_9419,N_10996);
and U15508 (N_15508,N_8645,N_8602);
nor U15509 (N_15509,N_10632,N_10825);
and U15510 (N_15510,N_9075,N_10360);
nor U15511 (N_15511,N_11836,N_9454);
nand U15512 (N_15512,N_11665,N_9806);
or U15513 (N_15513,N_8703,N_9389);
or U15514 (N_15514,N_10629,N_9164);
or U15515 (N_15515,N_11634,N_9297);
and U15516 (N_15516,N_8131,N_11431);
and U15517 (N_15517,N_9410,N_8079);
and U15518 (N_15518,N_9806,N_9922);
or U15519 (N_15519,N_9569,N_8892);
xnor U15520 (N_15520,N_10635,N_9359);
and U15521 (N_15521,N_8439,N_10755);
or U15522 (N_15522,N_8292,N_9012);
nor U15523 (N_15523,N_9564,N_11936);
nor U15524 (N_15524,N_10723,N_11745);
nand U15525 (N_15525,N_9728,N_8945);
nand U15526 (N_15526,N_10407,N_9021);
nor U15527 (N_15527,N_11941,N_8694);
and U15528 (N_15528,N_10136,N_9577);
or U15529 (N_15529,N_9288,N_10890);
xnor U15530 (N_15530,N_9655,N_11760);
and U15531 (N_15531,N_11545,N_8243);
or U15532 (N_15532,N_9874,N_8225);
xor U15533 (N_15533,N_10773,N_8062);
nor U15534 (N_15534,N_11882,N_10632);
nand U15535 (N_15535,N_8998,N_10394);
nand U15536 (N_15536,N_10480,N_10831);
or U15537 (N_15537,N_8143,N_10019);
nor U15538 (N_15538,N_10008,N_9262);
nor U15539 (N_15539,N_10880,N_11704);
or U15540 (N_15540,N_8900,N_10275);
xnor U15541 (N_15541,N_11460,N_10058);
and U15542 (N_15542,N_10315,N_11884);
or U15543 (N_15543,N_8462,N_11126);
and U15544 (N_15544,N_8543,N_10095);
or U15545 (N_15545,N_11347,N_8450);
nor U15546 (N_15546,N_10175,N_9624);
or U15547 (N_15547,N_9442,N_9735);
and U15548 (N_15548,N_11098,N_10600);
and U15549 (N_15549,N_8322,N_9267);
and U15550 (N_15550,N_11965,N_8716);
nand U15551 (N_15551,N_10994,N_10512);
nand U15552 (N_15552,N_9670,N_11161);
and U15553 (N_15553,N_9502,N_8509);
nand U15554 (N_15554,N_8081,N_11838);
xor U15555 (N_15555,N_11653,N_11043);
nor U15556 (N_15556,N_9971,N_9691);
xor U15557 (N_15557,N_8895,N_10865);
nor U15558 (N_15558,N_9294,N_11693);
and U15559 (N_15559,N_10579,N_11592);
nand U15560 (N_15560,N_11662,N_11975);
xnor U15561 (N_15561,N_10167,N_11632);
and U15562 (N_15562,N_8719,N_8260);
nand U15563 (N_15563,N_8503,N_8731);
nor U15564 (N_15564,N_10013,N_10926);
or U15565 (N_15565,N_9528,N_10524);
nor U15566 (N_15566,N_10913,N_10986);
xnor U15567 (N_15567,N_8528,N_9076);
nor U15568 (N_15568,N_9133,N_9083);
nor U15569 (N_15569,N_9820,N_9535);
nand U15570 (N_15570,N_8977,N_10740);
or U15571 (N_15571,N_10121,N_10018);
nand U15572 (N_15572,N_8204,N_8191);
or U15573 (N_15573,N_11106,N_11667);
and U15574 (N_15574,N_9054,N_9105);
and U15575 (N_15575,N_10224,N_11788);
xnor U15576 (N_15576,N_8101,N_8153);
nor U15577 (N_15577,N_10080,N_11139);
or U15578 (N_15578,N_11900,N_9156);
and U15579 (N_15579,N_8997,N_10669);
xnor U15580 (N_15580,N_11716,N_9134);
xor U15581 (N_15581,N_11091,N_9093);
and U15582 (N_15582,N_9642,N_10984);
and U15583 (N_15583,N_9207,N_10654);
or U15584 (N_15584,N_11101,N_8853);
or U15585 (N_15585,N_10808,N_10364);
and U15586 (N_15586,N_8663,N_8445);
nand U15587 (N_15587,N_8617,N_10421);
and U15588 (N_15588,N_11680,N_11269);
nand U15589 (N_15589,N_9883,N_11173);
xnor U15590 (N_15590,N_8039,N_9892);
and U15591 (N_15591,N_11269,N_9069);
xnor U15592 (N_15592,N_11990,N_11834);
or U15593 (N_15593,N_8053,N_9414);
nor U15594 (N_15594,N_11092,N_9864);
or U15595 (N_15595,N_11961,N_10393);
and U15596 (N_15596,N_11016,N_9804);
and U15597 (N_15597,N_11499,N_9409);
nor U15598 (N_15598,N_9427,N_10273);
or U15599 (N_15599,N_10201,N_11038);
nor U15600 (N_15600,N_11962,N_9688);
nor U15601 (N_15601,N_9379,N_9704);
nor U15602 (N_15602,N_11429,N_8693);
xnor U15603 (N_15603,N_8687,N_8877);
xor U15604 (N_15604,N_9421,N_8498);
xor U15605 (N_15605,N_8740,N_11973);
xnor U15606 (N_15606,N_9797,N_11147);
nand U15607 (N_15607,N_8841,N_9027);
nor U15608 (N_15608,N_10092,N_9563);
nor U15609 (N_15609,N_9894,N_9663);
nand U15610 (N_15610,N_10195,N_9021);
or U15611 (N_15611,N_8290,N_11414);
nor U15612 (N_15612,N_11775,N_9925);
nor U15613 (N_15613,N_10392,N_11396);
and U15614 (N_15614,N_9939,N_8413);
nand U15615 (N_15615,N_9307,N_9978);
nor U15616 (N_15616,N_10815,N_8178);
nor U15617 (N_15617,N_10258,N_9447);
xnor U15618 (N_15618,N_10212,N_8897);
xnor U15619 (N_15619,N_10767,N_8820);
xnor U15620 (N_15620,N_10093,N_11643);
and U15621 (N_15621,N_8460,N_11712);
nor U15622 (N_15622,N_8681,N_11077);
nor U15623 (N_15623,N_11122,N_9769);
nand U15624 (N_15624,N_9599,N_10257);
nand U15625 (N_15625,N_9021,N_10478);
or U15626 (N_15626,N_9573,N_8444);
or U15627 (N_15627,N_8022,N_9284);
and U15628 (N_15628,N_11269,N_11710);
xor U15629 (N_15629,N_10659,N_8152);
xnor U15630 (N_15630,N_10751,N_10985);
and U15631 (N_15631,N_11103,N_10935);
and U15632 (N_15632,N_10356,N_10446);
xor U15633 (N_15633,N_10708,N_11095);
xor U15634 (N_15634,N_8841,N_11159);
and U15635 (N_15635,N_9517,N_8349);
nand U15636 (N_15636,N_11477,N_11142);
and U15637 (N_15637,N_9788,N_8460);
nor U15638 (N_15638,N_9907,N_9674);
and U15639 (N_15639,N_9111,N_9752);
nand U15640 (N_15640,N_11793,N_10438);
xor U15641 (N_15641,N_9808,N_11805);
nor U15642 (N_15642,N_11892,N_10923);
nand U15643 (N_15643,N_8343,N_8595);
nand U15644 (N_15644,N_10659,N_9212);
nor U15645 (N_15645,N_8549,N_9155);
nand U15646 (N_15646,N_8955,N_10836);
nand U15647 (N_15647,N_10219,N_8347);
and U15648 (N_15648,N_8065,N_11686);
xor U15649 (N_15649,N_10822,N_8209);
or U15650 (N_15650,N_11302,N_9806);
nor U15651 (N_15651,N_8215,N_11206);
and U15652 (N_15652,N_8456,N_9497);
xor U15653 (N_15653,N_10463,N_11552);
and U15654 (N_15654,N_9667,N_9236);
nor U15655 (N_15655,N_11829,N_10186);
or U15656 (N_15656,N_11605,N_9602);
or U15657 (N_15657,N_9601,N_8206);
or U15658 (N_15658,N_8073,N_8689);
and U15659 (N_15659,N_8951,N_9566);
or U15660 (N_15660,N_10739,N_10291);
nor U15661 (N_15661,N_9514,N_10137);
nand U15662 (N_15662,N_10252,N_11595);
or U15663 (N_15663,N_10975,N_11532);
nand U15664 (N_15664,N_11676,N_9531);
nand U15665 (N_15665,N_10416,N_9275);
xnor U15666 (N_15666,N_9102,N_11423);
or U15667 (N_15667,N_10657,N_10242);
nand U15668 (N_15668,N_9523,N_8966);
nand U15669 (N_15669,N_9696,N_8493);
nor U15670 (N_15670,N_10753,N_11009);
and U15671 (N_15671,N_11483,N_10495);
nand U15672 (N_15672,N_10230,N_10088);
or U15673 (N_15673,N_9416,N_10790);
and U15674 (N_15674,N_8677,N_9492);
or U15675 (N_15675,N_11940,N_9831);
nor U15676 (N_15676,N_8501,N_10791);
or U15677 (N_15677,N_10659,N_8728);
nand U15678 (N_15678,N_10209,N_10537);
nor U15679 (N_15679,N_9074,N_9508);
or U15680 (N_15680,N_9828,N_8124);
nor U15681 (N_15681,N_10039,N_11645);
nand U15682 (N_15682,N_9657,N_9591);
nor U15683 (N_15683,N_9975,N_10023);
xor U15684 (N_15684,N_10347,N_11140);
or U15685 (N_15685,N_10997,N_10156);
or U15686 (N_15686,N_8129,N_9835);
or U15687 (N_15687,N_9103,N_10427);
and U15688 (N_15688,N_11899,N_11519);
nor U15689 (N_15689,N_10328,N_9702);
xnor U15690 (N_15690,N_10037,N_9556);
xor U15691 (N_15691,N_11455,N_11772);
and U15692 (N_15692,N_11222,N_10011);
nand U15693 (N_15693,N_11610,N_11057);
nand U15694 (N_15694,N_10371,N_9408);
xor U15695 (N_15695,N_8832,N_11136);
nand U15696 (N_15696,N_11537,N_9848);
nor U15697 (N_15697,N_10497,N_11959);
or U15698 (N_15698,N_10040,N_8325);
nor U15699 (N_15699,N_8394,N_8265);
or U15700 (N_15700,N_10285,N_9619);
nor U15701 (N_15701,N_8063,N_8433);
or U15702 (N_15702,N_10446,N_10351);
xor U15703 (N_15703,N_8534,N_11564);
nor U15704 (N_15704,N_8337,N_8640);
or U15705 (N_15705,N_11953,N_10532);
nor U15706 (N_15706,N_10719,N_11079);
nor U15707 (N_15707,N_9151,N_8074);
nand U15708 (N_15708,N_11681,N_11433);
xnor U15709 (N_15709,N_11777,N_11532);
nor U15710 (N_15710,N_8913,N_11593);
or U15711 (N_15711,N_11114,N_9100);
nor U15712 (N_15712,N_11223,N_8949);
and U15713 (N_15713,N_8127,N_8727);
nand U15714 (N_15714,N_10565,N_8044);
or U15715 (N_15715,N_10796,N_11280);
and U15716 (N_15716,N_8100,N_11661);
or U15717 (N_15717,N_9028,N_10239);
nand U15718 (N_15718,N_8863,N_11639);
or U15719 (N_15719,N_9241,N_11371);
and U15720 (N_15720,N_11005,N_10530);
nand U15721 (N_15721,N_8534,N_8603);
nand U15722 (N_15722,N_10760,N_9693);
and U15723 (N_15723,N_9827,N_8907);
and U15724 (N_15724,N_8008,N_8915);
and U15725 (N_15725,N_11782,N_8053);
and U15726 (N_15726,N_9231,N_11502);
or U15727 (N_15727,N_10190,N_9820);
xor U15728 (N_15728,N_9738,N_11068);
and U15729 (N_15729,N_9256,N_10640);
xnor U15730 (N_15730,N_11870,N_11555);
nor U15731 (N_15731,N_9903,N_11118);
and U15732 (N_15732,N_8966,N_10494);
nand U15733 (N_15733,N_11805,N_9400);
nor U15734 (N_15734,N_9047,N_8066);
nand U15735 (N_15735,N_11569,N_9129);
or U15736 (N_15736,N_10011,N_11651);
nand U15737 (N_15737,N_9502,N_10834);
nor U15738 (N_15738,N_9585,N_9282);
xnor U15739 (N_15739,N_9345,N_11386);
or U15740 (N_15740,N_10811,N_11384);
and U15741 (N_15741,N_9072,N_8055);
nand U15742 (N_15742,N_8780,N_9403);
nor U15743 (N_15743,N_8889,N_11668);
and U15744 (N_15744,N_10091,N_9620);
and U15745 (N_15745,N_8115,N_9182);
xnor U15746 (N_15746,N_10406,N_9641);
or U15747 (N_15747,N_10987,N_11611);
xnor U15748 (N_15748,N_9813,N_11906);
nand U15749 (N_15749,N_9980,N_8469);
xor U15750 (N_15750,N_10251,N_10072);
nand U15751 (N_15751,N_8396,N_8908);
or U15752 (N_15752,N_11144,N_8195);
nand U15753 (N_15753,N_11369,N_8625);
nand U15754 (N_15754,N_8390,N_11882);
nor U15755 (N_15755,N_9589,N_10545);
xor U15756 (N_15756,N_8340,N_8271);
xor U15757 (N_15757,N_8652,N_10268);
and U15758 (N_15758,N_11820,N_9168);
or U15759 (N_15759,N_8475,N_8170);
or U15760 (N_15760,N_9934,N_9370);
xnor U15761 (N_15761,N_10186,N_10995);
xor U15762 (N_15762,N_11222,N_11198);
nor U15763 (N_15763,N_8052,N_9571);
nor U15764 (N_15764,N_10513,N_8076);
or U15765 (N_15765,N_8522,N_8260);
or U15766 (N_15766,N_9589,N_8808);
and U15767 (N_15767,N_11497,N_11105);
and U15768 (N_15768,N_10264,N_11981);
nor U15769 (N_15769,N_10447,N_10063);
or U15770 (N_15770,N_9533,N_8018);
nor U15771 (N_15771,N_11399,N_10705);
xnor U15772 (N_15772,N_8022,N_9073);
nand U15773 (N_15773,N_8808,N_9370);
or U15774 (N_15774,N_9233,N_11203);
nor U15775 (N_15775,N_10492,N_8115);
and U15776 (N_15776,N_10239,N_9309);
nand U15777 (N_15777,N_9931,N_9425);
nor U15778 (N_15778,N_8574,N_8595);
xnor U15779 (N_15779,N_10167,N_9139);
nor U15780 (N_15780,N_8184,N_11635);
nand U15781 (N_15781,N_9860,N_10908);
nand U15782 (N_15782,N_11355,N_8987);
or U15783 (N_15783,N_9658,N_8062);
or U15784 (N_15784,N_11322,N_11523);
xnor U15785 (N_15785,N_10199,N_8148);
nand U15786 (N_15786,N_8358,N_10671);
or U15787 (N_15787,N_9652,N_8612);
and U15788 (N_15788,N_10103,N_9183);
or U15789 (N_15789,N_8697,N_8072);
nor U15790 (N_15790,N_9524,N_8331);
or U15791 (N_15791,N_11478,N_10922);
xor U15792 (N_15792,N_8479,N_10162);
xor U15793 (N_15793,N_9356,N_10566);
nand U15794 (N_15794,N_9658,N_8785);
or U15795 (N_15795,N_9517,N_9446);
and U15796 (N_15796,N_10219,N_10118);
nor U15797 (N_15797,N_10012,N_8468);
xor U15798 (N_15798,N_9292,N_9515);
and U15799 (N_15799,N_11005,N_8884);
nand U15800 (N_15800,N_9305,N_8065);
or U15801 (N_15801,N_9952,N_10297);
xnor U15802 (N_15802,N_8202,N_11387);
or U15803 (N_15803,N_8958,N_9967);
or U15804 (N_15804,N_11514,N_10192);
nor U15805 (N_15805,N_10759,N_11091);
nor U15806 (N_15806,N_11539,N_11916);
or U15807 (N_15807,N_10737,N_10783);
or U15808 (N_15808,N_11743,N_8442);
nand U15809 (N_15809,N_8589,N_8088);
or U15810 (N_15810,N_8939,N_9027);
or U15811 (N_15811,N_9916,N_8097);
and U15812 (N_15812,N_11960,N_10879);
and U15813 (N_15813,N_11603,N_10031);
nor U15814 (N_15814,N_11999,N_8912);
xor U15815 (N_15815,N_10378,N_11761);
or U15816 (N_15816,N_9261,N_9133);
and U15817 (N_15817,N_11892,N_11596);
or U15818 (N_15818,N_11917,N_11171);
or U15819 (N_15819,N_8324,N_11791);
and U15820 (N_15820,N_8119,N_11794);
xnor U15821 (N_15821,N_10399,N_9187);
xor U15822 (N_15822,N_11323,N_10044);
nor U15823 (N_15823,N_9909,N_11134);
and U15824 (N_15824,N_9199,N_8108);
or U15825 (N_15825,N_11862,N_10896);
xnor U15826 (N_15826,N_8271,N_9423);
nand U15827 (N_15827,N_11185,N_10415);
xor U15828 (N_15828,N_8816,N_11726);
and U15829 (N_15829,N_10648,N_9195);
xnor U15830 (N_15830,N_11481,N_11321);
nand U15831 (N_15831,N_10823,N_8767);
nor U15832 (N_15832,N_10325,N_9048);
and U15833 (N_15833,N_10868,N_8070);
or U15834 (N_15834,N_9887,N_11276);
and U15835 (N_15835,N_11778,N_9325);
xor U15836 (N_15836,N_8017,N_10188);
nor U15837 (N_15837,N_11525,N_10850);
and U15838 (N_15838,N_8666,N_9688);
and U15839 (N_15839,N_9253,N_11331);
nor U15840 (N_15840,N_11201,N_8960);
or U15841 (N_15841,N_10892,N_11992);
nand U15842 (N_15842,N_8826,N_8653);
or U15843 (N_15843,N_10834,N_9097);
nand U15844 (N_15844,N_9951,N_11912);
and U15845 (N_15845,N_9569,N_9603);
xnor U15846 (N_15846,N_9280,N_10368);
or U15847 (N_15847,N_8855,N_11743);
or U15848 (N_15848,N_10144,N_11121);
xnor U15849 (N_15849,N_10340,N_9353);
nand U15850 (N_15850,N_9271,N_10664);
and U15851 (N_15851,N_10227,N_10623);
nor U15852 (N_15852,N_9902,N_10077);
nor U15853 (N_15853,N_9956,N_11733);
nand U15854 (N_15854,N_11163,N_9765);
nor U15855 (N_15855,N_8865,N_9306);
and U15856 (N_15856,N_8024,N_9633);
nor U15857 (N_15857,N_8463,N_11688);
nand U15858 (N_15858,N_8884,N_10083);
nor U15859 (N_15859,N_9584,N_9212);
nand U15860 (N_15860,N_10654,N_10470);
and U15861 (N_15861,N_11516,N_8757);
xnor U15862 (N_15862,N_11848,N_11567);
nor U15863 (N_15863,N_9943,N_8399);
and U15864 (N_15864,N_10377,N_11533);
xor U15865 (N_15865,N_9081,N_8780);
nand U15866 (N_15866,N_8683,N_11017);
or U15867 (N_15867,N_10815,N_11542);
xor U15868 (N_15868,N_10874,N_9390);
or U15869 (N_15869,N_9406,N_11826);
and U15870 (N_15870,N_10228,N_8913);
nor U15871 (N_15871,N_11320,N_9333);
xnor U15872 (N_15872,N_9048,N_11611);
nor U15873 (N_15873,N_11392,N_9125);
nand U15874 (N_15874,N_10705,N_11731);
nand U15875 (N_15875,N_9379,N_11842);
and U15876 (N_15876,N_8841,N_9208);
nand U15877 (N_15877,N_9632,N_8578);
or U15878 (N_15878,N_10201,N_11827);
nand U15879 (N_15879,N_8928,N_8388);
and U15880 (N_15880,N_8187,N_10579);
or U15881 (N_15881,N_11030,N_10264);
or U15882 (N_15882,N_11161,N_11030);
nand U15883 (N_15883,N_8858,N_9431);
or U15884 (N_15884,N_9957,N_10386);
nand U15885 (N_15885,N_9767,N_10335);
nand U15886 (N_15886,N_11922,N_10996);
nand U15887 (N_15887,N_8241,N_11615);
nor U15888 (N_15888,N_11783,N_8851);
or U15889 (N_15889,N_11996,N_10051);
nand U15890 (N_15890,N_10224,N_8820);
nand U15891 (N_15891,N_11360,N_10853);
nor U15892 (N_15892,N_11638,N_9632);
and U15893 (N_15893,N_8045,N_8686);
xnor U15894 (N_15894,N_10824,N_9389);
and U15895 (N_15895,N_11279,N_9085);
and U15896 (N_15896,N_10169,N_9069);
nand U15897 (N_15897,N_9061,N_11804);
nor U15898 (N_15898,N_8605,N_8113);
nor U15899 (N_15899,N_11530,N_10846);
xor U15900 (N_15900,N_11632,N_9944);
and U15901 (N_15901,N_11701,N_10003);
nor U15902 (N_15902,N_8853,N_9219);
nor U15903 (N_15903,N_8262,N_9205);
xor U15904 (N_15904,N_8993,N_11762);
nor U15905 (N_15905,N_10802,N_8218);
and U15906 (N_15906,N_11851,N_11070);
and U15907 (N_15907,N_10434,N_9099);
xnor U15908 (N_15908,N_9206,N_11089);
nor U15909 (N_15909,N_10783,N_10781);
nand U15910 (N_15910,N_9471,N_10077);
and U15911 (N_15911,N_9361,N_11102);
or U15912 (N_15912,N_11939,N_11604);
nand U15913 (N_15913,N_11677,N_9175);
nand U15914 (N_15914,N_10255,N_9528);
xor U15915 (N_15915,N_11267,N_9041);
xnor U15916 (N_15916,N_11548,N_9022);
or U15917 (N_15917,N_11543,N_9558);
or U15918 (N_15918,N_10924,N_11950);
or U15919 (N_15919,N_9914,N_8429);
and U15920 (N_15920,N_10526,N_10388);
nor U15921 (N_15921,N_11354,N_10147);
and U15922 (N_15922,N_8035,N_10560);
and U15923 (N_15923,N_9141,N_11939);
nand U15924 (N_15924,N_11457,N_11662);
nand U15925 (N_15925,N_11176,N_10261);
and U15926 (N_15926,N_8175,N_11402);
nand U15927 (N_15927,N_10325,N_10686);
nand U15928 (N_15928,N_11657,N_9263);
xnor U15929 (N_15929,N_9529,N_8841);
nand U15930 (N_15930,N_11688,N_11312);
or U15931 (N_15931,N_10921,N_10179);
nand U15932 (N_15932,N_10599,N_9299);
nand U15933 (N_15933,N_9291,N_9540);
nor U15934 (N_15934,N_11697,N_11745);
xor U15935 (N_15935,N_10919,N_9503);
nor U15936 (N_15936,N_11639,N_9551);
or U15937 (N_15937,N_8509,N_11666);
xnor U15938 (N_15938,N_8512,N_11978);
nor U15939 (N_15939,N_8071,N_10703);
or U15940 (N_15940,N_11874,N_11848);
nand U15941 (N_15941,N_9882,N_10948);
nand U15942 (N_15942,N_10499,N_10776);
and U15943 (N_15943,N_10279,N_11536);
and U15944 (N_15944,N_9728,N_10873);
nor U15945 (N_15945,N_9651,N_10260);
nor U15946 (N_15946,N_11715,N_9646);
nor U15947 (N_15947,N_11965,N_11729);
and U15948 (N_15948,N_11120,N_11992);
and U15949 (N_15949,N_10533,N_10691);
or U15950 (N_15950,N_10926,N_9975);
or U15951 (N_15951,N_11827,N_8058);
nor U15952 (N_15952,N_8447,N_11409);
xor U15953 (N_15953,N_8862,N_10054);
or U15954 (N_15954,N_10075,N_9076);
xor U15955 (N_15955,N_9383,N_11756);
nand U15956 (N_15956,N_9132,N_10298);
xnor U15957 (N_15957,N_8466,N_11585);
or U15958 (N_15958,N_10468,N_9148);
xnor U15959 (N_15959,N_11628,N_10269);
nor U15960 (N_15960,N_11521,N_9908);
nand U15961 (N_15961,N_8287,N_10186);
nand U15962 (N_15962,N_10595,N_9600);
and U15963 (N_15963,N_8251,N_10664);
and U15964 (N_15964,N_9169,N_10015);
xor U15965 (N_15965,N_9219,N_9905);
nor U15966 (N_15966,N_9855,N_10703);
nand U15967 (N_15967,N_11025,N_8792);
or U15968 (N_15968,N_9211,N_10204);
or U15969 (N_15969,N_9644,N_11383);
and U15970 (N_15970,N_10121,N_10760);
or U15971 (N_15971,N_10698,N_10687);
or U15972 (N_15972,N_8374,N_11554);
or U15973 (N_15973,N_8660,N_9321);
nand U15974 (N_15974,N_10371,N_9764);
xor U15975 (N_15975,N_9621,N_10355);
or U15976 (N_15976,N_10018,N_10508);
xor U15977 (N_15977,N_8380,N_11993);
and U15978 (N_15978,N_11473,N_10185);
or U15979 (N_15979,N_11261,N_9319);
or U15980 (N_15980,N_8121,N_11199);
and U15981 (N_15981,N_11315,N_11000);
and U15982 (N_15982,N_11771,N_11550);
nand U15983 (N_15983,N_8346,N_9821);
nand U15984 (N_15984,N_9312,N_8687);
or U15985 (N_15985,N_9090,N_8610);
nor U15986 (N_15986,N_10258,N_9663);
or U15987 (N_15987,N_9743,N_10785);
nand U15988 (N_15988,N_8359,N_10056);
nand U15989 (N_15989,N_8886,N_10691);
and U15990 (N_15990,N_9679,N_10163);
nand U15991 (N_15991,N_9890,N_10764);
nor U15992 (N_15992,N_11568,N_9828);
nor U15993 (N_15993,N_11270,N_10822);
and U15994 (N_15994,N_10353,N_8222);
nand U15995 (N_15995,N_9494,N_10906);
and U15996 (N_15996,N_8180,N_9633);
nand U15997 (N_15997,N_8983,N_8460);
or U15998 (N_15998,N_8835,N_9299);
and U15999 (N_15999,N_10370,N_11638);
and U16000 (N_16000,N_13102,N_12366);
or U16001 (N_16001,N_14331,N_15043);
nand U16002 (N_16002,N_14046,N_14790);
nand U16003 (N_16003,N_14542,N_12479);
or U16004 (N_16004,N_13084,N_12017);
xnor U16005 (N_16005,N_13182,N_13960);
or U16006 (N_16006,N_14213,N_12820);
or U16007 (N_16007,N_13567,N_12877);
and U16008 (N_16008,N_14184,N_13258);
and U16009 (N_16009,N_12000,N_15965);
and U16010 (N_16010,N_14474,N_14422);
xnor U16011 (N_16011,N_15277,N_15023);
nand U16012 (N_16012,N_12764,N_12657);
nor U16013 (N_16013,N_12559,N_12093);
or U16014 (N_16014,N_12548,N_12429);
nand U16015 (N_16015,N_14693,N_12505);
xnor U16016 (N_16016,N_15552,N_15814);
or U16017 (N_16017,N_13251,N_15512);
nand U16018 (N_16018,N_15659,N_12907);
xnor U16019 (N_16019,N_13246,N_12159);
nand U16020 (N_16020,N_15346,N_15788);
xor U16021 (N_16021,N_13552,N_14214);
and U16022 (N_16022,N_12055,N_15977);
nor U16023 (N_16023,N_14522,N_12014);
xor U16024 (N_16024,N_12279,N_14098);
xor U16025 (N_16025,N_15707,N_12362);
nor U16026 (N_16026,N_13684,N_12135);
and U16027 (N_16027,N_12941,N_14351);
nand U16028 (N_16028,N_15418,N_15143);
xor U16029 (N_16029,N_14970,N_15596);
or U16030 (N_16030,N_12403,N_13000);
or U16031 (N_16031,N_15085,N_15913);
or U16032 (N_16032,N_13659,N_12805);
xnor U16033 (N_16033,N_15833,N_12164);
or U16034 (N_16034,N_12507,N_15310);
or U16035 (N_16035,N_13028,N_14961);
xnor U16036 (N_16036,N_12622,N_13024);
nor U16037 (N_16037,N_14062,N_15269);
and U16038 (N_16038,N_14118,N_12608);
nand U16039 (N_16039,N_12328,N_12220);
xnor U16040 (N_16040,N_14018,N_14910);
nor U16041 (N_16041,N_13771,N_13862);
or U16042 (N_16042,N_12564,N_13207);
or U16043 (N_16043,N_14303,N_12112);
or U16044 (N_16044,N_13350,N_14721);
or U16045 (N_16045,N_13139,N_15472);
and U16046 (N_16046,N_14334,N_14732);
or U16047 (N_16047,N_14060,N_15754);
and U16048 (N_16048,N_15199,N_14020);
nor U16049 (N_16049,N_12800,N_12817);
or U16050 (N_16050,N_13415,N_12294);
and U16051 (N_16051,N_14851,N_13098);
and U16052 (N_16052,N_15349,N_13388);
and U16053 (N_16053,N_14038,N_12193);
nand U16054 (N_16054,N_15654,N_15585);
xor U16055 (N_16055,N_14688,N_13205);
nand U16056 (N_16056,N_14800,N_15210);
nand U16057 (N_16057,N_14363,N_15226);
nor U16058 (N_16058,N_15846,N_12818);
xnor U16059 (N_16059,N_13829,N_15054);
or U16060 (N_16060,N_12659,N_15114);
or U16061 (N_16061,N_14051,N_12268);
and U16062 (N_16062,N_14504,N_12632);
or U16063 (N_16063,N_15302,N_13640);
nor U16064 (N_16064,N_14263,N_13790);
and U16065 (N_16065,N_14544,N_14737);
nor U16066 (N_16066,N_12644,N_13734);
and U16067 (N_16067,N_12188,N_12738);
or U16068 (N_16068,N_12183,N_15436);
and U16069 (N_16069,N_14899,N_14571);
nand U16070 (N_16070,N_13656,N_14487);
nand U16071 (N_16071,N_15159,N_13781);
xnor U16072 (N_16072,N_15448,N_15527);
nor U16073 (N_16073,N_15225,N_15459);
xor U16074 (N_16074,N_13772,N_14215);
xor U16075 (N_16075,N_15460,N_13166);
xnor U16076 (N_16076,N_13204,N_12934);
nand U16077 (N_16077,N_13530,N_12936);
or U16078 (N_16078,N_15799,N_15883);
nor U16079 (N_16079,N_15174,N_12672);
nand U16080 (N_16080,N_13389,N_15372);
nor U16081 (N_16081,N_13383,N_14228);
or U16082 (N_16082,N_15755,N_13067);
nand U16083 (N_16083,N_15781,N_15286);
and U16084 (N_16084,N_12256,N_14682);
or U16085 (N_16085,N_14364,N_14878);
nor U16086 (N_16086,N_14403,N_12955);
or U16087 (N_16087,N_12367,N_14901);
xor U16088 (N_16088,N_14005,N_14077);
or U16089 (N_16089,N_12722,N_12804);
or U16090 (N_16090,N_15762,N_14229);
nand U16091 (N_16091,N_15200,N_15075);
nand U16092 (N_16092,N_15865,N_15259);
nor U16093 (N_16093,N_12196,N_15874);
nor U16094 (N_16094,N_13343,N_14358);
nand U16095 (N_16095,N_13577,N_13932);
nand U16096 (N_16096,N_13517,N_13588);
xnor U16097 (N_16097,N_13587,N_15869);
nand U16098 (N_16098,N_13602,N_13606);
nand U16099 (N_16099,N_15780,N_12034);
nand U16100 (N_16100,N_15766,N_15104);
nand U16101 (N_16101,N_12139,N_12615);
nor U16102 (N_16102,N_14289,N_12058);
nand U16103 (N_16103,N_13228,N_12953);
and U16104 (N_16104,N_12359,N_13768);
and U16105 (N_16105,N_15936,N_13706);
nor U16106 (N_16106,N_14557,N_12788);
xnor U16107 (N_16107,N_13574,N_15001);
nand U16108 (N_16108,N_14012,N_13676);
and U16109 (N_16109,N_14521,N_15972);
and U16110 (N_16110,N_12070,N_14966);
and U16111 (N_16111,N_14026,N_12902);
nand U16112 (N_16112,N_12521,N_15169);
nor U16113 (N_16113,N_13441,N_14455);
nor U16114 (N_16114,N_15635,N_12660);
nand U16115 (N_16115,N_14669,N_13725);
and U16116 (N_16116,N_14711,N_15028);
nand U16117 (N_16117,N_14196,N_13490);
nand U16118 (N_16118,N_12218,N_13275);
and U16119 (N_16119,N_13624,N_15880);
and U16120 (N_16120,N_12869,N_13203);
or U16121 (N_16121,N_14868,N_12591);
or U16122 (N_16122,N_12501,N_12245);
or U16123 (N_16123,N_13793,N_12832);
nor U16124 (N_16124,N_14823,N_15440);
xnor U16125 (N_16125,N_13023,N_14153);
or U16126 (N_16126,N_15840,N_14843);
and U16127 (N_16127,N_12520,N_15040);
or U16128 (N_16128,N_14766,N_14404);
xor U16129 (N_16129,N_13831,N_15523);
and U16130 (N_16130,N_12449,N_15734);
nor U16131 (N_16131,N_13455,N_14607);
nand U16132 (N_16132,N_15951,N_12562);
or U16133 (N_16133,N_12233,N_13549);
and U16134 (N_16134,N_14925,N_12103);
nand U16135 (N_16135,N_15929,N_13578);
nor U16136 (N_16136,N_13679,N_12285);
nand U16137 (N_16137,N_12810,N_15580);
xor U16138 (N_16138,N_14939,N_15901);
or U16139 (N_16139,N_13525,N_13064);
or U16140 (N_16140,N_13945,N_12225);
nand U16141 (N_16141,N_12595,N_13833);
xnor U16142 (N_16142,N_15690,N_13425);
nand U16143 (N_16143,N_15307,N_15417);
or U16144 (N_16144,N_15565,N_12523);
nand U16145 (N_16145,N_14269,N_14142);
or U16146 (N_16146,N_13596,N_14643);
nor U16147 (N_16147,N_12172,N_12799);
or U16148 (N_16148,N_15910,N_12555);
nor U16149 (N_16149,N_15966,N_14202);
or U16150 (N_16150,N_13086,N_14774);
nor U16151 (N_16151,N_15052,N_14988);
and U16152 (N_16152,N_14420,N_14964);
nor U16153 (N_16153,N_14848,N_14382);
or U16154 (N_16154,N_15904,N_12690);
or U16155 (N_16155,N_12508,N_14628);
or U16156 (N_16156,N_14250,N_14494);
nand U16157 (N_16157,N_15557,N_15623);
nor U16158 (N_16158,N_14989,N_12254);
xnor U16159 (N_16159,N_15399,N_12387);
or U16160 (N_16160,N_13621,N_14284);
and U16161 (N_16161,N_14114,N_13159);
and U16162 (N_16162,N_14928,N_15794);
xor U16163 (N_16163,N_12516,N_14943);
nor U16164 (N_16164,N_13542,N_12852);
nor U16165 (N_16165,N_12857,N_15428);
or U16166 (N_16166,N_12336,N_12871);
nand U16167 (N_16167,N_15918,N_15341);
nand U16168 (N_16168,N_15894,N_15669);
or U16169 (N_16169,N_14389,N_14483);
nor U16170 (N_16170,N_13110,N_12179);
nand U16171 (N_16171,N_15497,N_13079);
xor U16172 (N_16172,N_14468,N_15204);
and U16173 (N_16173,N_13398,N_13215);
and U16174 (N_16174,N_15222,N_13052);
or U16175 (N_16175,N_12811,N_15037);
or U16176 (N_16176,N_12077,N_12781);
nand U16177 (N_16177,N_15937,N_13172);
xnor U16178 (N_16178,N_12209,N_15775);
nor U16179 (N_16179,N_13322,N_13677);
xnor U16180 (N_16180,N_13816,N_15208);
or U16181 (N_16181,N_14911,N_14211);
or U16182 (N_16182,N_12812,N_12942);
and U16183 (N_16183,N_12861,N_13360);
nor U16184 (N_16184,N_14563,N_15543);
and U16185 (N_16185,N_14958,N_14866);
nor U16186 (N_16186,N_12290,N_15240);
xor U16187 (N_16187,N_13265,N_14997);
or U16188 (N_16188,N_14112,N_13674);
or U16189 (N_16189,N_14700,N_13498);
or U16190 (N_16190,N_15335,N_13197);
xnor U16191 (N_16191,N_15671,N_13035);
xnor U16192 (N_16192,N_12709,N_12797);
nor U16193 (N_16193,N_14169,N_12249);
and U16194 (N_16194,N_12854,N_12281);
or U16195 (N_16195,N_15514,N_15297);
and U16196 (N_16196,N_12736,N_12594);
nand U16197 (N_16197,N_12727,N_14765);
nand U16198 (N_16198,N_13106,N_15742);
and U16199 (N_16199,N_15125,N_15357);
and U16200 (N_16200,N_12607,N_15116);
and U16201 (N_16201,N_13237,N_13927);
xor U16202 (N_16202,N_15246,N_12324);
xor U16203 (N_16203,N_15877,N_13280);
or U16204 (N_16204,N_12757,N_13128);
xnor U16205 (N_16205,N_12122,N_15267);
nand U16206 (N_16206,N_13984,N_14400);
xor U16207 (N_16207,N_14632,N_15684);
or U16208 (N_16208,N_15151,N_12908);
nand U16209 (N_16209,N_15279,N_13012);
and U16210 (N_16210,N_12025,N_12692);
xor U16211 (N_16211,N_12386,N_13925);
nor U16212 (N_16212,N_14820,N_12205);
or U16213 (N_16213,N_12938,N_12782);
and U16214 (N_16214,N_13737,N_15410);
and U16215 (N_16215,N_14406,N_14549);
nor U16216 (N_16216,N_12625,N_13896);
and U16217 (N_16217,N_15163,N_14443);
nand U16218 (N_16218,N_15491,N_15171);
xnor U16219 (N_16219,N_13309,N_13785);
or U16220 (N_16220,N_15607,N_12866);
xnor U16221 (N_16221,N_12089,N_13700);
and U16222 (N_16222,N_14094,N_14120);
nand U16223 (N_16223,N_13374,N_13008);
nor U16224 (N_16224,N_12851,N_13328);
nand U16225 (N_16225,N_13426,N_15262);
xnor U16226 (N_16226,N_13288,N_15393);
or U16227 (N_16227,N_12988,N_13773);
xor U16228 (N_16228,N_15138,N_12785);
and U16229 (N_16229,N_12105,N_12629);
nand U16230 (N_16230,N_12566,N_14985);
xor U16231 (N_16231,N_12539,N_12189);
xor U16232 (N_16232,N_15147,N_14084);
and U16233 (N_16233,N_12260,N_14712);
or U16234 (N_16234,N_12377,N_12044);
xnor U16235 (N_16235,N_15636,N_14762);
or U16236 (N_16236,N_14503,N_15048);
nor U16237 (N_16237,N_14893,N_15777);
nor U16238 (N_16238,N_15213,N_12911);
xor U16239 (N_16239,N_15017,N_15696);
or U16240 (N_16240,N_12012,N_12373);
xnor U16241 (N_16241,N_12943,N_14245);
nand U16242 (N_16242,N_14031,N_12028);
and U16243 (N_16243,N_13997,N_13715);
and U16244 (N_16244,N_14696,N_14687);
nor U16245 (N_16245,N_12976,N_13645);
or U16246 (N_16246,N_15935,N_13241);
or U16247 (N_16247,N_14496,N_12925);
nor U16248 (N_16248,N_14044,N_13034);
nand U16249 (N_16249,N_14424,N_15857);
or U16250 (N_16250,N_14772,N_15254);
nand U16251 (N_16251,N_13681,N_14828);
and U16252 (N_16252,N_14749,N_14923);
nor U16253 (N_16253,N_14539,N_14520);
nand U16254 (N_16254,N_13272,N_14663);
nor U16255 (N_16255,N_15375,N_13902);
or U16256 (N_16256,N_12470,N_14174);
nor U16257 (N_16257,N_12345,N_14755);
or U16258 (N_16258,N_13568,N_15748);
nand U16259 (N_16259,N_14075,N_14055);
nand U16260 (N_16260,N_15651,N_15887);
nand U16261 (N_16261,N_13652,N_13890);
or U16262 (N_16262,N_14336,N_12829);
nand U16263 (N_16263,N_12540,N_13999);
and U16264 (N_16264,N_14286,N_15729);
or U16265 (N_16265,N_13589,N_14897);
xnor U16266 (N_16266,N_14004,N_12212);
or U16267 (N_16267,N_15178,N_12675);
nand U16268 (N_16268,N_13148,N_15994);
nand U16269 (N_16269,N_12541,N_14518);
nand U16270 (N_16270,N_14282,N_15480);
nor U16271 (N_16271,N_12425,N_14953);
or U16272 (N_16272,N_12104,N_13256);
xor U16273 (N_16273,N_12261,N_15381);
xnor U16274 (N_16274,N_14740,N_14272);
nand U16275 (N_16275,N_14817,N_15987);
or U16276 (N_16276,N_14088,N_12990);
and U16277 (N_16277,N_15526,N_14109);
nand U16278 (N_16278,N_15212,N_15203);
and U16279 (N_16279,N_13779,N_13669);
or U16280 (N_16280,N_13184,N_15000);
or U16281 (N_16281,N_12513,N_13274);
and U16282 (N_16282,N_14163,N_13060);
nand U16283 (N_16283,N_12506,N_12614);
and U16284 (N_16284,N_12453,N_12570);
and U16285 (N_16285,N_14234,N_12211);
or U16286 (N_16286,N_14301,N_15946);
and U16287 (N_16287,N_12519,N_15458);
nand U16288 (N_16288,N_14507,N_14600);
nor U16289 (N_16289,N_13692,N_14512);
or U16290 (N_16290,N_13848,N_12219);
or U16291 (N_16291,N_13232,N_15377);
or U16292 (N_16292,N_14806,N_14847);
nor U16293 (N_16293,N_14147,N_14064);
or U16294 (N_16294,N_15640,N_14535);
xor U16295 (N_16295,N_12855,N_12201);
nand U16296 (N_16296,N_14572,N_13996);
nor U16297 (N_16297,N_14456,N_12300);
or U16298 (N_16298,N_14429,N_15678);
nor U16299 (N_16299,N_14954,N_14362);
nor U16300 (N_16300,N_12415,N_14484);
xor U16301 (N_16301,N_15049,N_12666);
xor U16302 (N_16302,N_12525,N_13056);
nor U16303 (N_16303,N_12119,N_13100);
xor U16304 (N_16304,N_13391,N_15942);
and U16305 (N_16305,N_12282,N_12627);
or U16306 (N_16306,N_14130,N_13860);
or U16307 (N_16307,N_15862,N_12503);
nor U16308 (N_16308,N_14172,N_12773);
nor U16309 (N_16309,N_13562,N_13013);
nor U16310 (N_16310,N_13564,N_15949);
nand U16311 (N_16311,N_15504,N_13193);
or U16312 (N_16312,N_12596,N_13963);
nand U16313 (N_16313,N_14872,N_12108);
xnor U16314 (N_16314,N_15677,N_15312);
nand U16315 (N_16315,N_13697,N_12983);
and U16316 (N_16316,N_12531,N_12224);
nor U16317 (N_16317,N_15627,N_14380);
nor U16318 (N_16318,N_14891,N_12668);
xnor U16319 (N_16319,N_15905,N_13017);
nand U16320 (N_16320,N_12320,N_12763);
nor U16321 (N_16321,N_13263,N_15193);
nand U16322 (N_16322,N_12749,N_12039);
and U16323 (N_16323,N_13137,N_12681);
nand U16324 (N_16324,N_15045,N_14168);
or U16325 (N_16325,N_13791,N_12963);
and U16326 (N_16326,N_12563,N_13775);
xnor U16327 (N_16327,N_12417,N_12534);
and U16328 (N_16328,N_15184,N_15321);
or U16329 (N_16329,N_13036,N_12447);
nand U16330 (N_16330,N_13906,N_14050);
nor U16331 (N_16331,N_14764,N_14701);
nor U16332 (N_16332,N_15231,N_12396);
xnor U16333 (N_16333,N_15265,N_12707);
xnor U16334 (N_16334,N_12400,N_14582);
and U16335 (N_16335,N_13381,N_12244);
and U16336 (N_16336,N_13230,N_12035);
or U16337 (N_16337,N_14857,N_14871);
xor U16338 (N_16338,N_12951,N_15120);
and U16339 (N_16339,N_12289,N_15939);
and U16340 (N_16340,N_13248,N_14041);
nand U16341 (N_16341,N_12654,N_14787);
nor U16342 (N_16342,N_12372,N_15584);
xor U16343 (N_16343,N_14792,N_13800);
or U16344 (N_16344,N_14782,N_14812);
nor U16345 (N_16345,N_15498,N_13423);
xnor U16346 (N_16346,N_13660,N_12361);
and U16347 (N_16347,N_14049,N_15340);
nor U16348 (N_16348,N_12128,N_13158);
xnor U16349 (N_16349,N_15986,N_12796);
nand U16350 (N_16350,N_14637,N_13937);
xnor U16351 (N_16351,N_13006,N_15071);
or U16352 (N_16352,N_15324,N_12806);
nand U16353 (N_16353,N_13134,N_12185);
xnor U16354 (N_16354,N_14569,N_12716);
and U16355 (N_16355,N_15257,N_12027);
and U16356 (N_16356,N_14809,N_15510);
nand U16357 (N_16357,N_15858,N_13912);
nand U16358 (N_16358,N_12498,N_15400);
xnor U16359 (N_16359,N_12755,N_15122);
or U16360 (N_16360,N_13186,N_14015);
or U16361 (N_16361,N_12008,N_14299);
and U16362 (N_16362,N_13142,N_12978);
or U16363 (N_16363,N_13119,N_14803);
nor U16364 (N_16364,N_15978,N_14073);
xor U16365 (N_16365,N_13929,N_12079);
or U16366 (N_16366,N_12216,N_12074);
xor U16367 (N_16367,N_13088,N_14306);
xnor U16368 (N_16368,N_14720,N_13598);
and U16369 (N_16369,N_13864,N_12643);
nor U16370 (N_16370,N_13620,N_12354);
and U16371 (N_16371,N_14208,N_12437);
xor U16372 (N_16372,N_13509,N_15087);
xnor U16373 (N_16373,N_12919,N_13846);
or U16374 (N_16374,N_15509,N_14070);
and U16375 (N_16375,N_13075,N_14635);
or U16376 (N_16376,N_12502,N_12231);
or U16377 (N_16377,N_13018,N_14345);
xnor U16378 (N_16378,N_14519,N_12426);
and U16379 (N_16379,N_14831,N_12792);
nor U16380 (N_16380,N_14279,N_12980);
xor U16381 (N_16381,N_14421,N_15061);
nor U16382 (N_16382,N_15318,N_14273);
xor U16383 (N_16383,N_15332,N_14531);
xor U16384 (N_16384,N_13515,N_13078);
nor U16385 (N_16385,N_13613,N_13866);
or U16386 (N_16386,N_12131,N_14541);
nand U16387 (N_16387,N_14763,N_13192);
nor U16388 (N_16388,N_15759,N_13767);
nand U16389 (N_16389,N_12137,N_12464);
nand U16390 (N_16390,N_12102,N_15772);
or U16391 (N_16391,N_14113,N_12038);
or U16392 (N_16392,N_15657,N_15642);
and U16393 (N_16393,N_15374,N_12752);
nor U16394 (N_16394,N_15035,N_15610);
or U16395 (N_16395,N_12630,N_14902);
and U16396 (N_16396,N_14952,N_13301);
nand U16397 (N_16397,N_12054,N_12868);
xnor U16398 (N_16398,N_15027,N_15360);
or U16399 (N_16399,N_13375,N_14019);
xor U16400 (N_16400,N_13962,N_15342);
xnor U16401 (N_16401,N_14668,N_13225);
and U16402 (N_16402,N_15508,N_14680);
xnor U16403 (N_16403,N_12132,N_15442);
nor U16404 (N_16404,N_14283,N_14853);
nor U16405 (N_16405,N_15959,N_14069);
nor U16406 (N_16406,N_15232,N_12473);
nor U16407 (N_16407,N_14573,N_14661);
nor U16408 (N_16408,N_13903,N_12650);
and U16409 (N_16409,N_13479,N_13751);
nand U16410 (N_16410,N_14210,N_12917);
nor U16411 (N_16411,N_13413,N_12306);
or U16412 (N_16412,N_13546,N_12445);
and U16413 (N_16413,N_14779,N_14167);
and U16414 (N_16414,N_14973,N_15366);
nor U16415 (N_16415,N_12891,N_14604);
and U16416 (N_16416,N_14955,N_14944);
xor U16417 (N_16417,N_13736,N_13691);
and U16418 (N_16418,N_14469,N_14488);
nand U16419 (N_16419,N_13130,N_13163);
nor U16420 (N_16420,N_14904,N_15033);
and U16421 (N_16421,N_15077,N_12247);
nand U16422 (N_16422,N_13117,N_14277);
and U16423 (N_16423,N_15823,N_15237);
xor U16424 (N_16424,N_12087,N_12766);
or U16425 (N_16425,N_13538,N_14021);
nand U16426 (N_16426,N_15485,N_12931);
or U16427 (N_16427,N_14960,N_14719);
nand U16428 (N_16428,N_13459,N_12830);
or U16429 (N_16429,N_12569,N_13276);
xor U16430 (N_16430,N_14558,N_14589);
nand U16431 (N_16431,N_14645,N_12542);
or U16432 (N_16432,N_14934,N_12465);
xor U16433 (N_16433,N_13714,N_13419);
or U16434 (N_16434,N_14880,N_14586);
nand U16435 (N_16435,N_12126,N_15817);
nand U16436 (N_16436,N_14583,N_15095);
xnor U16437 (N_16437,N_12063,N_14742);
nor U16438 (N_16438,N_15562,N_13814);
nor U16439 (N_16439,N_14735,N_13755);
xor U16440 (N_16440,N_12878,N_14935);
nand U16441 (N_16441,N_12845,N_12295);
or U16442 (N_16442,N_13852,N_12343);
nand U16443 (N_16443,N_14786,N_12318);
and U16444 (N_16444,N_13758,N_12839);
and U16445 (N_16445,N_12537,N_13626);
and U16446 (N_16446,N_12587,N_14625);
xor U16447 (N_16447,N_15551,N_15680);
nand U16448 (N_16448,N_14956,N_12822);
xor U16449 (N_16449,N_14833,N_12332);
nand U16450 (N_16450,N_15709,N_14007);
or U16451 (N_16451,N_14411,N_15970);
xor U16452 (N_16452,N_13238,N_12062);
nor U16453 (N_16453,N_14950,N_15743);
nor U16454 (N_16454,N_14894,N_13686);
nor U16455 (N_16455,N_12571,N_15922);
or U16456 (N_16456,N_15244,N_13721);
nor U16457 (N_16457,N_12157,N_15142);
nor U16458 (N_16458,N_13959,N_15423);
or U16459 (N_16459,N_15433,N_12151);
or U16460 (N_16460,N_12843,N_15047);
or U16461 (N_16461,N_14689,N_15801);
xor U16462 (N_16462,N_12037,N_14937);
and U16463 (N_16463,N_12357,N_13534);
or U16464 (N_16464,N_13292,N_12146);
xor U16465 (N_16465,N_12375,N_15747);
nor U16466 (N_16466,N_13654,N_12613);
nor U16467 (N_16467,N_13319,N_13311);
or U16468 (N_16468,N_13111,N_15656);
or U16469 (N_16469,N_12731,N_13540);
or U16470 (N_16470,N_14236,N_14825);
xnor U16471 (N_16471,N_15084,N_12085);
nand U16472 (N_16472,N_13742,N_13453);
nand U16473 (N_16473,N_15521,N_12379);
xor U16474 (N_16474,N_12748,N_15813);
or U16475 (N_16475,N_12069,N_13727);
nor U16476 (N_16476,N_14029,N_15720);
nand U16477 (N_16477,N_12674,N_12259);
nor U16478 (N_16478,N_13764,N_14481);
nand U16479 (N_16479,N_13298,N_15046);
or U16480 (N_16480,N_12952,N_13089);
xor U16481 (N_16481,N_12496,N_13002);
or U16482 (N_16482,N_14375,N_12005);
xor U16483 (N_16483,N_15735,N_13231);
and U16484 (N_16484,N_15566,N_14080);
nand U16485 (N_16485,N_14132,N_12251);
nor U16486 (N_16486,N_14854,N_13026);
nand U16487 (N_16487,N_12100,N_12700);
and U16488 (N_16488,N_14328,N_14649);
xor U16489 (N_16489,N_12200,N_13612);
or U16490 (N_16490,N_13061,N_13488);
and U16491 (N_16491,N_12348,N_15844);
nor U16492 (N_16492,N_15652,N_13302);
and U16493 (N_16493,N_15556,N_15141);
xnor U16494 (N_16494,N_12360,N_14315);
and U16495 (N_16495,N_15902,N_12967);
nand U16496 (N_16496,N_13745,N_15838);
xor U16497 (N_16497,N_14365,N_13443);
nand U16498 (N_16498,N_15295,N_14949);
xnor U16499 (N_16499,N_12895,N_13746);
xor U16500 (N_16500,N_14342,N_13502);
nand U16501 (N_16501,N_12402,N_14395);
and U16502 (N_16502,N_13405,N_13236);
nand U16503 (N_16503,N_12689,N_12779);
nor U16504 (N_16504,N_15317,N_12031);
and U16505 (N_16505,N_15675,N_15752);
xor U16506 (N_16506,N_14523,N_12580);
nor U16507 (N_16507,N_12664,N_13330);
nand U16508 (N_16508,N_13402,N_14619);
or U16509 (N_16509,N_15903,N_14292);
nand U16510 (N_16510,N_13065,N_13329);
nor U16511 (N_16511,N_12834,N_12616);
nor U16512 (N_16512,N_15909,N_15029);
xor U16513 (N_16513,N_12169,N_15378);
nor U16514 (N_16514,N_13429,N_13304);
and U16515 (N_16515,N_12962,N_13438);
or U16516 (N_16516,N_14023,N_12896);
nand U16517 (N_16517,N_12497,N_13390);
xnor U16518 (N_16518,N_13961,N_12984);
and U16519 (N_16519,N_12443,N_15558);
nor U16520 (N_16520,N_12686,N_15756);
and U16521 (N_16521,N_13487,N_13716);
and U16522 (N_16522,N_15135,N_15301);
nor U16523 (N_16523,N_14751,N_13323);
nor U16524 (N_16524,N_13603,N_13054);
nor U16525 (N_16525,N_14591,N_13440);
nand U16526 (N_16526,N_12057,N_14707);
nand U16527 (N_16527,N_12450,N_13969);
nand U16528 (N_16528,N_15326,N_15981);
xnor U16529 (N_16529,N_14577,N_13543);
and U16530 (N_16530,N_12095,N_14335);
or U16531 (N_16531,N_15383,N_15784);
nor U16532 (N_16532,N_15700,N_13009);
and U16533 (N_16533,N_14968,N_13257);
nor U16534 (N_16534,N_15351,N_14929);
xnor U16535 (N_16535,N_13261,N_14010);
xor U16536 (N_16536,N_15173,N_12499);
nor U16537 (N_16537,N_14884,N_13647);
nand U16538 (N_16538,N_15875,N_15518);
xnor U16539 (N_16539,N_12641,N_13795);
and U16540 (N_16540,N_15117,N_15189);
nor U16541 (N_16541,N_13282,N_13217);
or U16542 (N_16542,N_13956,N_13571);
nor U16543 (N_16543,N_13718,N_15167);
nor U16544 (N_16544,N_15396,N_12986);
and U16545 (N_16545,N_12026,N_14071);
nor U16546 (N_16546,N_13518,N_12459);
or U16547 (N_16547,N_15150,N_15331);
nand U16548 (N_16548,N_14810,N_13942);
xnor U16549 (N_16549,N_13713,N_15009);
nand U16550 (N_16550,N_14407,N_14595);
nand U16551 (N_16551,N_13638,N_12050);
or U16552 (N_16552,N_14150,N_13774);
and U16553 (N_16553,N_15258,N_15545);
nor U16554 (N_16554,N_15287,N_15586);
nand U16555 (N_16555,N_15571,N_13373);
nor U16556 (N_16556,N_13105,N_13930);
and U16557 (N_16557,N_14471,N_13869);
nor U16558 (N_16558,N_14994,N_12836);
xor U16559 (N_16559,N_15081,N_15461);
and U16560 (N_16560,N_15807,N_14511);
or U16561 (N_16561,N_12322,N_14316);
xor U16562 (N_16562,N_13467,N_12195);
and U16563 (N_16563,N_14660,N_14148);
and U16564 (N_16564,N_13566,N_15289);
nand U16565 (N_16565,N_14673,N_15736);
nor U16566 (N_16566,N_15890,N_15774);
xor U16567 (N_16567,N_12374,N_13899);
or U16568 (N_16568,N_13726,N_13722);
nor U16569 (N_16569,N_14408,N_14222);
and U16570 (N_16570,N_12161,N_13699);
xor U16571 (N_16571,N_13744,N_15737);
nand U16572 (N_16572,N_12724,N_14832);
nor U16573 (N_16573,N_12418,N_15127);
nor U16574 (N_16574,N_13152,N_15697);
nor U16575 (N_16575,N_13689,N_13448);
nand U16576 (N_16576,N_12859,N_13551);
xnor U16577 (N_16577,N_14295,N_15725);
and U16578 (N_16578,N_15648,N_15996);
nor U16579 (N_16579,N_14115,N_15506);
and U16580 (N_16580,N_15064,N_13879);
and U16581 (N_16581,N_14037,N_13802);
or U16582 (N_16582,N_14886,N_13908);
and U16583 (N_16583,N_15379,N_13711);
nand U16584 (N_16584,N_14611,N_12168);
nor U16585 (N_16585,N_15599,N_15495);
and U16586 (N_16586,N_15924,N_15305);
xnor U16587 (N_16587,N_13641,N_15102);
and U16588 (N_16588,N_12321,N_14137);
and U16589 (N_16589,N_15073,N_12267);
and U16590 (N_16590,N_14372,N_13407);
nor U16591 (N_16591,N_13695,N_13346);
or U16592 (N_16592,N_15646,N_14435);
nand U16593 (N_16593,N_13125,N_14233);
or U16594 (N_16594,N_13160,N_13213);
and U16595 (N_16595,N_12856,N_14042);
nand U16596 (N_16596,N_15422,N_14346);
nor U16597 (N_16597,N_12884,N_15316);
nor U16598 (N_16598,N_15835,N_15311);
and U16599 (N_16599,N_13476,N_12957);
or U16600 (N_16600,N_15170,N_14254);
nor U16601 (N_16601,N_15129,N_13041);
and U16602 (N_16602,N_13757,N_15507);
xor U16603 (N_16603,N_14072,N_13032);
or U16604 (N_16604,N_14624,N_13433);
nor U16605 (N_16605,N_12944,N_15502);
and U16606 (N_16606,N_15940,N_15053);
nor U16607 (N_16607,N_14501,N_14308);
or U16608 (N_16608,N_14561,N_12626);
and U16609 (N_16609,N_14243,N_12427);
nand U16610 (N_16610,N_13162,N_12030);
and U16611 (N_16611,N_14996,N_13850);
xor U16612 (N_16612,N_13395,N_13741);
and U16613 (N_16613,N_15960,N_12317);
nand U16614 (N_16614,N_12765,N_15811);
or U16615 (N_16615,N_14220,N_14467);
nor U16616 (N_16616,N_15567,N_13586);
xor U16617 (N_16617,N_13770,N_13364);
nand U16618 (N_16618,N_15411,N_14144);
and U16619 (N_16619,N_14553,N_13499);
and U16620 (N_16620,N_13151,N_14480);
xnor U16621 (N_16621,N_15796,N_14634);
nor U16622 (N_16622,N_14185,N_14057);
and U16623 (N_16623,N_14811,N_15416);
nand U16624 (N_16624,N_13359,N_12954);
xor U16625 (N_16625,N_14508,N_12148);
nor U16626 (N_16626,N_15180,N_14203);
nor U16627 (N_16627,N_14490,N_13868);
nand U16628 (N_16628,N_15055,N_14546);
nor U16629 (N_16629,N_14465,N_13820);
or U16630 (N_16630,N_13055,N_15338);
and U16631 (N_16631,N_15911,N_15106);
or U16632 (N_16632,N_13289,N_13437);
nor U16633 (N_16633,N_13226,N_14492);
and U16634 (N_16634,N_14580,N_12353);
nor U16635 (N_16635,N_12874,N_12873);
or U16636 (N_16636,N_13417,N_14417);
nand U16637 (N_16637,N_15455,N_14826);
and U16638 (N_16638,N_12847,N_15984);
xor U16639 (N_16639,N_14709,N_14366);
xnor U16640 (N_16640,N_14441,N_15194);
or U16641 (N_16641,N_14399,N_13553);
xnor U16642 (N_16642,N_15323,N_14390);
nand U16643 (N_16643,N_15609,N_14230);
xnor U16644 (N_16644,N_12789,N_12325);
or U16645 (N_16645,N_12365,N_13877);
xnor U16646 (N_16646,N_12706,N_15293);
or U16647 (N_16647,N_13762,N_15907);
nor U16648 (N_16648,N_15481,N_15109);
or U16649 (N_16649,N_12494,N_13687);
xnor U16650 (N_16650,N_13095,N_15224);
nand U16651 (N_16651,N_15661,N_15097);
and U16652 (N_16652,N_14699,N_13955);
xnor U16653 (N_16653,N_13030,N_14918);
or U16654 (N_16654,N_14242,N_12270);
xor U16655 (N_16655,N_12628,N_13842);
nand U16656 (N_16656,N_15309,N_12222);
or U16657 (N_16657,N_13609,N_15443);
nand U16658 (N_16658,N_15975,N_12786);
nand U16659 (N_16659,N_14337,N_15172);
xnor U16660 (N_16660,N_13325,N_13510);
nor U16661 (N_16661,N_14844,N_13031);
and U16662 (N_16662,N_15993,N_13732);
nand U16663 (N_16663,N_15275,N_15253);
nor U16664 (N_16664,N_15590,N_12113);
nor U16665 (N_16665,N_13817,N_12182);
xor U16666 (N_16666,N_13112,N_13680);
xor U16667 (N_16667,N_12890,N_13297);
xnor U16668 (N_16668,N_14175,N_14837);
or U16669 (N_16669,N_15804,N_15401);
and U16670 (N_16670,N_13941,N_14177);
nand U16671 (N_16671,N_12699,N_15574);
xor U16672 (N_16672,N_15820,N_14183);
and U16673 (N_16673,N_12680,N_15444);
and U16674 (N_16674,N_12198,N_15487);
nor U16675 (N_16675,N_13888,N_14081);
nand U16676 (N_16676,N_14313,N_14106);
nand U16677 (N_16677,N_13472,N_13505);
xnor U16678 (N_16678,N_14397,N_14355);
or U16679 (N_16679,N_13607,N_13704);
or U16680 (N_16680,N_13935,N_12229);
nor U16681 (N_16681,N_12326,N_15274);
and U16682 (N_16682,N_14703,N_15739);
nor U16683 (N_16683,N_15611,N_12914);
and U16684 (N_16684,N_15841,N_13029);
nand U16685 (N_16685,N_12439,N_14191);
nand U16686 (N_16686,N_12180,N_15067);
or U16687 (N_16687,N_13858,N_13622);
or U16688 (N_16688,N_14993,N_14223);
and U16689 (N_16689,N_13449,N_14193);
or U16690 (N_16690,N_13920,N_12682);
xor U16691 (N_16691,N_15930,N_13780);
nor U16692 (N_16692,N_15519,N_12802);
and U16693 (N_16693,N_14917,N_12213);
nand U16694 (N_16694,N_13165,N_15281);
nor U16695 (N_16695,N_15753,N_15414);
or U16696 (N_16696,N_14548,N_14017);
nand U16697 (N_16697,N_15927,N_15870);
and U16698 (N_16698,N_12485,N_13167);
and U16699 (N_16699,N_13457,N_15803);
xor U16700 (N_16700,N_13563,N_15291);
nand U16701 (N_16701,N_13880,N_15068);
nor U16702 (N_16702,N_15836,N_12546);
and U16703 (N_16703,N_12667,N_13174);
or U16704 (N_16704,N_12423,N_12922);
nand U16705 (N_16705,N_15439,N_15536);
and U16706 (N_16706,N_12844,N_14922);
or U16707 (N_16707,N_15831,N_15158);
nand U16708 (N_16708,N_12080,N_13044);
nand U16709 (N_16709,N_12140,N_14377);
nor U16710 (N_16710,N_15544,N_12734);
nor U16711 (N_16711,N_13458,N_15353);
nand U16712 (N_16712,N_12454,N_14097);
and U16713 (N_16713,N_14875,N_15146);
nand U16714 (N_16714,N_14659,N_13978);
xor U16715 (N_16715,N_13337,N_13815);
or U16716 (N_16716,N_12619,N_14438);
nand U16717 (N_16717,N_15062,N_15608);
nor U16718 (N_16718,N_12414,N_13657);
or U16719 (N_16719,N_13911,N_14805);
xnor U16720 (N_16720,N_13936,N_15576);
or U16721 (N_16721,N_13526,N_12471);
nor U16722 (N_16722,N_15348,N_15663);
and U16723 (N_16723,N_14227,N_15207);
and U16724 (N_16724,N_15496,N_12585);
and U16725 (N_16725,N_14451,N_14984);
and U16726 (N_16726,N_15021,N_15394);
nor U16727 (N_16727,N_14385,N_12767);
or U16728 (N_16728,N_13445,N_15474);
and U16729 (N_16729,N_15490,N_12864);
and U16730 (N_16730,N_14333,N_15828);
or U16731 (N_16731,N_13227,N_15888);
xnor U16732 (N_16732,N_12081,N_14592);
or U16733 (N_16733,N_12610,N_14281);
nand U16734 (N_16734,N_14027,N_14783);
nor U16735 (N_16735,N_14271,N_13336);
xor U16736 (N_16736,N_15637,N_15368);
and U16737 (N_16737,N_12665,N_14255);
or U16738 (N_16738,N_14338,N_12370);
and U16739 (N_16739,N_13211,N_14698);
nor U16740 (N_16740,N_15397,N_15407);
xnor U16741 (N_16741,N_14760,N_15082);
and U16742 (N_16742,N_13033,N_12947);
or U16743 (N_16743,N_14567,N_13572);
nand U16744 (N_16744,N_15738,N_12578);
and U16745 (N_16745,N_14753,N_13447);
and U16746 (N_16746,N_13792,N_12518);
nand U16747 (N_16747,N_15952,N_15183);
nand U16748 (N_16748,N_13164,N_12278);
or U16749 (N_16749,N_12824,N_12111);
xor U16750 (N_16750,N_13729,N_15466);
nand U16751 (N_16751,N_13341,N_14946);
and U16752 (N_16752,N_12973,N_12436);
or U16753 (N_16753,N_14510,N_15653);
xnor U16754 (N_16754,N_14009,N_14259);
nand U16755 (N_16755,N_13837,N_13210);
nor U16756 (N_16756,N_14264,N_12395);
or U16757 (N_16757,N_13957,N_15529);
nor U16758 (N_16758,N_15908,N_14850);
and U16759 (N_16759,N_13305,N_13819);
nor U16760 (N_16760,N_12551,N_12187);
or U16761 (N_16761,N_14127,N_12826);
nor U16762 (N_16762,N_13273,N_12138);
and U16763 (N_16763,N_12334,N_15492);
xor U16764 (N_16764,N_15850,N_13580);
or U16765 (N_16765,N_12088,N_15468);
or U16766 (N_16766,N_14116,N_13967);
nor U16767 (N_16767,N_13672,N_14076);
nor U16768 (N_16768,N_14139,N_13262);
nand U16769 (N_16769,N_12206,N_12549);
nor U16770 (N_16770,N_12795,N_13870);
and U16771 (N_16771,N_13508,N_12670);
and U16772 (N_16772,N_12648,N_12637);
nor U16773 (N_16773,N_12492,N_15221);
xnor U16774 (N_16774,N_13242,N_15845);
nor U16775 (N_16775,N_13315,N_12011);
nand U16776 (N_16776,N_14562,N_14574);
xnor U16777 (N_16777,N_13884,N_14348);
nand U16778 (N_16778,N_14319,N_13717);
nand U16779 (N_16779,N_13914,N_15517);
and U16780 (N_16780,N_13900,N_14339);
nor U16781 (N_16781,N_12683,N_12303);
nor U16782 (N_16782,N_14915,N_12053);
or U16783 (N_16783,N_12557,N_12049);
nand U16784 (N_16784,N_15819,N_14559);
xor U16785 (N_16785,N_13783,N_14555);
xor U16786 (N_16786,N_12833,N_14609);
nor U16787 (N_16787,N_15464,N_14194);
and U16788 (N_16788,N_12676,N_15878);
and U16789 (N_16789,N_15484,N_13735);
xor U16790 (N_16790,N_13421,N_15470);
or U16791 (N_16791,N_14726,N_12448);
or U16792 (N_16792,N_12430,N_14750);
xnor U16793 (N_16793,N_14138,N_15177);
nor U16794 (N_16794,N_15899,N_12215);
xor U16795 (N_16795,N_15145,N_15148);
or U16796 (N_16796,N_13981,N_14444);
or U16797 (N_16797,N_15079,N_14105);
nand U16798 (N_16798,N_13901,N_15101);
nand U16799 (N_16799,N_14368,N_13201);
nand U16800 (N_16800,N_14002,N_12441);
and U16801 (N_16801,N_15776,N_13295);
and U16802 (N_16802,N_13907,N_15815);
xnor U16803 (N_16803,N_12530,N_12171);
xor U16804 (N_16804,N_13474,N_15091);
and U16805 (N_16805,N_12226,N_15619);
xor U16806 (N_16806,N_12246,N_15779);
nor U16807 (N_16807,N_15670,N_12036);
nor U16808 (N_16808,N_14056,N_12433);
or U16809 (N_16809,N_15013,N_13759);
nor U16810 (N_16810,N_13522,N_13254);
nor U16811 (N_16811,N_15721,N_13332);
xor U16812 (N_16812,N_13823,N_15511);
xnor U16813 (N_16813,N_14815,N_13739);
and U16814 (N_16814,N_12356,N_15546);
nor U16815 (N_16815,N_12388,N_14477);
xor U16816 (N_16816,N_15283,N_15294);
and U16817 (N_16817,N_15818,N_12892);
and U16818 (N_16818,N_15218,N_14125);
or U16819 (N_16819,N_14111,N_12634);
nand U16820 (N_16820,N_12770,N_13799);
or U16821 (N_16821,N_12556,N_15060);
and U16822 (N_16822,N_12886,N_14458);
and U16823 (N_16823,N_13385,N_15629);
nor U16824 (N_16824,N_12581,N_15915);
xor U16825 (N_16825,N_15467,N_12186);
nand U16826 (N_16826,N_13648,N_14302);
or U16827 (N_16827,N_15974,N_15825);
or U16828 (N_16828,N_13849,N_14131);
nor U16829 (N_16829,N_15398,N_12611);
nand U16830 (N_16830,N_15044,N_14432);
or U16831 (N_16831,N_14158,N_14667);
and U16832 (N_16832,N_13895,N_13495);
and U16833 (N_16833,N_15731,N_13378);
nor U16834 (N_16834,N_13855,N_13356);
or U16835 (N_16835,N_14298,N_15728);
nor U16836 (N_16836,N_14614,N_12301);
nor U16837 (N_16837,N_13471,N_15765);
xnor U16838 (N_16838,N_12097,N_14226);
nor U16839 (N_16839,N_14892,N_14770);
or U16840 (N_16840,N_14594,N_12535);
or U16841 (N_16841,N_12655,N_14486);
nor U16842 (N_16842,N_13806,N_14398);
nand U16843 (N_16843,N_12725,N_13396);
or U16844 (N_16844,N_13094,N_14224);
nand U16845 (N_16845,N_13761,N_13342);
nand U16846 (N_16846,N_12582,N_15800);
xnor U16847 (N_16847,N_15961,N_13528);
nand U16848 (N_16848,N_15534,N_15991);
and U16849 (N_16849,N_15008,N_12828);
xnor U16850 (N_16850,N_13196,N_14793);
nor U16851 (N_16851,N_14967,N_12384);
nand U16852 (N_16852,N_12966,N_14171);
and U16853 (N_16853,N_14052,N_15769);
and U16854 (N_16854,N_15469,N_13853);
and U16855 (N_16855,N_13998,N_14882);
xnor U16856 (N_16856,N_15805,N_15185);
nand U16857 (N_16857,N_15750,N_12517);
nand U16858 (N_16858,N_15525,N_13214);
and U16859 (N_16859,N_15370,N_14525);
and U16860 (N_16860,N_14995,N_15356);
nand U16861 (N_16861,N_14895,N_13818);
and U16862 (N_16862,N_12703,N_12344);
or U16863 (N_16863,N_15941,N_14361);
xor U16864 (N_16864,N_13608,N_14907);
or U16865 (N_16865,N_15699,N_15718);
nand U16866 (N_16866,N_14849,N_12750);
or U16867 (N_16867,N_13170,N_14900);
nand U16868 (N_16868,N_12712,N_14291);
xor U16869 (N_16869,N_14597,N_12780);
nand U16870 (N_16870,N_13972,N_13581);
nand U16871 (N_16871,N_15555,N_12949);
and U16872 (N_16872,N_12879,N_13986);
and U16873 (N_16873,N_14708,N_14722);
xor U16874 (N_16874,N_13178,N_14889);
and U16875 (N_16875,N_14881,N_14462);
xnor U16876 (N_16876,N_12013,N_13314);
xnor U16877 (N_16877,N_14646,N_14506);
or U16878 (N_16878,N_12228,N_12153);
nor U16879 (N_16879,N_13670,N_14278);
xnor U16880 (N_16880,N_15912,N_12073);
nor U16881 (N_16881,N_14290,N_13442);
and U16882 (N_16882,N_14500,N_13338);
nor U16883 (N_16883,N_13921,N_15427);
or U16884 (N_16884,N_12653,N_12236);
or U16885 (N_16885,N_12145,N_12803);
or U16886 (N_16886,N_15672,N_15074);
or U16887 (N_16887,N_13512,N_14305);
nand U16888 (N_16888,N_12298,N_14482);
nand U16889 (N_16889,N_12658,N_15425);
xnor U16890 (N_16890,N_13284,N_14327);
xnor U16891 (N_16891,N_15465,N_15821);
nor U16892 (N_16892,N_13556,N_14216);
and U16893 (N_16893,N_13630,N_14983);
nand U16894 (N_16894,N_13682,N_14166);
xor U16895 (N_16895,N_13470,N_14489);
xor U16896 (N_16896,N_14627,N_13610);
or U16897 (N_16897,N_15271,N_15578);
nand U16898 (N_16898,N_13027,N_14391);
nor U16899 (N_16899,N_13627,N_13354);
and U16900 (N_16900,N_12612,N_14692);
and U16901 (N_16901,N_13268,N_13983);
and U16902 (N_16902,N_14440,N_14543);
and U16903 (N_16903,N_13583,N_14716);
nand U16904 (N_16904,N_15998,N_12477);
and U16905 (N_16905,N_13382,N_14387);
nand U16906 (N_16906,N_14665,N_14947);
or U16907 (N_16907,N_15285,N_12305);
xor U16908 (N_16908,N_12754,N_12422);
xor U16909 (N_16909,N_12243,N_14430);
and U16910 (N_16910,N_14258,N_15650);
nand U16911 (N_16911,N_15625,N_15687);
or U16912 (N_16912,N_13267,N_13794);
nor U16913 (N_16913,N_13386,N_13221);
nand U16914 (N_16914,N_14623,N_14916);
and U16915 (N_16915,N_12769,N_12894);
nor U16916 (N_16916,N_14268,N_13335);
or U16917 (N_16917,N_15808,N_13651);
or U16918 (N_16918,N_14287,N_12526);
nor U16919 (N_16919,N_13200,N_15454);
xor U16920 (N_16920,N_13889,N_13918);
nand U16921 (N_16921,N_15945,N_12482);
nor U16922 (N_16922,N_12837,N_14992);
and U16923 (N_16923,N_13331,N_13090);
xor U16924 (N_16924,N_13436,N_12617);
nand U16925 (N_16925,N_12092,N_15190);
nand U16926 (N_16926,N_14244,N_15693);
xnor U16927 (N_16927,N_12977,N_13401);
xor U16928 (N_16928,N_14423,N_12190);
and U16929 (N_16929,N_15715,N_15706);
nand U16930 (N_16930,N_14888,N_13951);
nor U16931 (N_16931,N_15473,N_14251);
and U16932 (N_16932,N_14353,N_12469);
nor U16933 (N_16933,N_12758,N_15531);
and U16934 (N_16934,N_12958,N_15438);
xor U16935 (N_16935,N_12969,N_14675);
and U16936 (N_16936,N_15111,N_13843);
nor U16937 (N_16937,N_15980,N_12144);
xor U16938 (N_16938,N_15215,N_14942);
or U16939 (N_16939,N_12253,N_13547);
and U16940 (N_16940,N_14957,N_15031);
or U16941 (N_16941,N_13422,N_14373);
nor U16942 (N_16942,N_12339,N_15216);
and U16943 (N_16943,N_13296,N_13693);
and U16944 (N_16944,N_15505,N_14674);
or U16945 (N_16945,N_15235,N_12056);
or U16946 (N_16946,N_12309,N_14022);
nor U16947 (N_16947,N_15322,N_14173);
nor U16948 (N_16948,N_15770,N_15005);
and U16949 (N_16949,N_15290,N_14110);
or U16950 (N_16950,N_14493,N_15579);
nand U16951 (N_16951,N_14606,N_13592);
xor U16952 (N_16952,N_14769,N_12720);
or U16953 (N_16953,N_14221,N_15092);
nand U16954 (N_16954,N_13042,N_14461);
nand U16955 (N_16955,N_13461,N_13570);
xor U16956 (N_16956,N_12858,N_15406);
xnor U16957 (N_16957,N_14434,N_15475);
or U16958 (N_16958,N_12673,N_12527);
nor U16959 (N_16959,N_14585,N_13266);
and U16960 (N_16960,N_15421,N_12819);
or U16961 (N_16961,N_12018,N_13253);
xor U16962 (N_16962,N_15515,N_13579);
xor U16963 (N_16963,N_14323,N_14354);
xnor U16964 (N_16964,N_15260,N_13826);
xnor U16965 (N_16965,N_15477,N_13392);
or U16966 (N_16966,N_12718,N_15757);
or U16967 (N_16967,N_13202,N_14074);
and U16968 (N_16968,N_15415,N_13939);
xnor U16969 (N_16969,N_13696,N_15682);
nor U16970 (N_16970,N_14867,N_12084);
or U16971 (N_16971,N_12419,N_13367);
nand U16972 (N_16972,N_13928,N_14515);
and U16973 (N_16973,N_15668,N_15488);
xor U16974 (N_16974,N_14320,N_13279);
nor U16975 (N_16975,N_12933,N_15810);
nor U16976 (N_16976,N_14513,N_13154);
nand U16977 (N_16977,N_12532,N_13135);
nand U16978 (N_16978,N_15824,N_15773);
or U16979 (N_16979,N_14045,N_12831);
xnor U16980 (N_16980,N_12487,N_12434);
nand U16981 (N_16981,N_14841,N_13821);
nand U16982 (N_16982,N_14813,N_12001);
nand U16983 (N_16983,N_14412,N_13077);
and U16984 (N_16984,N_13212,N_12511);
or U16985 (N_16985,N_12997,N_13694);
nor U16986 (N_16986,N_15039,N_14636);
and U16987 (N_16987,N_14584,N_14360);
or U16988 (N_16988,N_14788,N_14164);
and U16989 (N_16989,N_14656,N_13703);
nor U16990 (N_16990,N_14647,N_14478);
and U16991 (N_16991,N_14690,N_14101);
nand U16992 (N_16992,N_13824,N_15420);
nand U16993 (N_16993,N_14063,N_13177);
nor U16994 (N_16994,N_13787,N_12435);
xor U16995 (N_16995,N_14463,N_14846);
nand U16996 (N_16996,N_14626,N_15798);
nor U16997 (N_16997,N_13478,N_13555);
or U16998 (N_16998,N_13637,N_12099);
nor U16999 (N_16999,N_13051,N_15369);
nor U17000 (N_17000,N_15022,N_13025);
nor U17001 (N_17001,N_14066,N_13114);
nand U17002 (N_17002,N_12191,N_15026);
and U17003 (N_17003,N_12483,N_13371);
nand U17004 (N_17004,N_14165,N_15166);
or U17005 (N_17005,N_15860,N_14517);
xor U17006 (N_17006,N_12340,N_13968);
nand U17007 (N_17007,N_13882,N_12544);
xnor U17008 (N_17008,N_12959,N_13801);
and U17009 (N_17009,N_15230,N_15489);
and U17010 (N_17010,N_12042,N_13074);
nor U17011 (N_17011,N_12762,N_15367);
or U17012 (N_17012,N_12717,N_14802);
nand U17013 (N_17013,N_15679,N_15633);
nor U17014 (N_17014,N_14620,N_14083);
and U17015 (N_17015,N_13618,N_12047);
nor U17016 (N_17016,N_13784,N_14836);
and U17017 (N_17017,N_13840,N_14212);
nand U17018 (N_17018,N_14349,N_15115);
xor U17019 (N_17019,N_15299,N_15155);
or U17020 (N_17020,N_15921,N_15108);
and U17021 (N_17021,N_14460,N_14948);
nand U17022 (N_17022,N_13991,N_12114);
xor U17023 (N_17023,N_13140,N_15694);
nand U17024 (N_17024,N_13913,N_14207);
or U17025 (N_17025,N_12747,N_15947);
and U17026 (N_17026,N_12639,N_12380);
or U17027 (N_17027,N_13506,N_13688);
or U17028 (N_17028,N_12350,N_13789);
nor U17029 (N_17029,N_14479,N_15730);
or U17030 (N_17030,N_12438,N_12152);
and U17031 (N_17031,N_15196,N_14485);
and U17032 (N_17032,N_13650,N_12910);
xor U17033 (N_17033,N_15673,N_13904);
nand U17034 (N_17034,N_14807,N_13264);
nand U17035 (N_17035,N_13798,N_14310);
xor U17036 (N_17036,N_15667,N_12410);
and U17037 (N_17037,N_13068,N_13063);
xor U17038 (N_17038,N_13597,N_12825);
or U17039 (N_17039,N_12992,N_13625);
nor U17040 (N_17040,N_15128,N_13224);
xor U17041 (N_17041,N_14091,N_14261);
nand U17042 (N_17042,N_13786,N_15598);
nand U17043 (N_17043,N_14498,N_12394);
xnor U17044 (N_17044,N_13181,N_13685);
xor U17045 (N_17045,N_14777,N_14034);
xor U17046 (N_17046,N_12872,N_13005);
or U17047 (N_17047,N_13206,N_15856);
nor U17048 (N_17048,N_13811,N_13804);
nand U17049 (N_17049,N_12130,N_12642);
nor U17050 (N_17050,N_12173,N_14524);
nand U17051 (N_17051,N_12597,N_13109);
and U17052 (N_17052,N_15920,N_14861);
and U17053 (N_17053,N_13990,N_13875);
nand U17054 (N_17054,N_12291,N_15893);
or U17055 (N_17055,N_15691,N_15462);
and U17056 (N_17056,N_15333,N_13541);
nor U17057 (N_17057,N_12467,N_14653);
or U17058 (N_17058,N_15624,N_14006);
xor U17059 (N_17059,N_14340,N_13797);
nand U17060 (N_17060,N_12838,N_12889);
nand U17061 (N_17061,N_13287,N_14001);
or U17062 (N_17062,N_15499,N_12771);
and U17063 (N_17063,N_12784,N_12898);
nand U17064 (N_17064,N_12592,N_12136);
xnor U17065 (N_17065,N_13492,N_15198);
xor U17066 (N_17066,N_13414,N_12455);
nand U17067 (N_17067,N_14566,N_14154);
nand U17068 (N_17068,N_12903,N_14821);
or U17069 (N_17069,N_13194,N_12401);
and U17070 (N_17070,N_12848,N_14738);
or U17071 (N_17071,N_13473,N_13400);
xnor U17072 (N_17072,N_13216,N_15594);
nand U17073 (N_17073,N_15354,N_13532);
or U17074 (N_17074,N_14392,N_14367);
nand U17075 (N_17075,N_15989,N_14702);
nor U17076 (N_17076,N_13513,N_14795);
xor U17077 (N_17077,N_13584,N_14999);
xor U17078 (N_17078,N_12051,N_14776);
and U17079 (N_17079,N_14528,N_15003);
nand U17080 (N_17080,N_12331,N_12274);
nand U17081 (N_17081,N_13524,N_15390);
nor U17082 (N_17082,N_13836,N_12584);
and U17083 (N_17083,N_13131,N_13573);
nor U17084 (N_17084,N_14296,N_15853);
or U17085 (N_17085,N_13039,N_13318);
nand U17086 (N_17086,N_12404,N_12174);
nor U17087 (N_17087,N_15563,N_15152);
or U17088 (N_17088,N_13993,N_15139);
or U17089 (N_17089,N_15176,N_12273);
nand U17090 (N_17090,N_12939,N_15154);
and U17091 (N_17091,N_13501,N_12003);
or U17092 (N_17092,N_15588,N_15157);
or U17093 (N_17093,N_13738,N_14149);
and U17094 (N_17094,N_15861,N_12491);
nand U17095 (N_17095,N_12509,N_14396);
and U17096 (N_17096,N_12466,N_15243);
xnor U17097 (N_17097,N_12971,N_12964);
nand U17098 (N_17098,N_15925,N_15430);
and U17099 (N_17099,N_13320,N_14393);
nand U17100 (N_17100,N_12846,N_13291);
nor U17101 (N_17101,N_12409,N_14560);
xnor U17102 (N_17102,N_12257,N_12813);
and U17103 (N_17103,N_15329,N_13873);
nor U17104 (N_17104,N_15376,N_13484);
nor U17105 (N_17105,N_13776,N_12333);
nand U17106 (N_17106,N_12961,N_14318);
and U17107 (N_17107,N_13387,N_12905);
or U17108 (N_17108,N_13037,N_13046);
nand U17109 (N_17109,N_12979,N_13673);
or U17110 (N_17110,N_14780,N_12107);
xnor U17111 (N_17111,N_15429,N_12993);
nor U17112 (N_17112,N_12850,N_13944);
nor U17113 (N_17113,N_12116,N_15708);
and U17114 (N_17114,N_12876,N_15561);
xor U17115 (N_17115,N_12292,N_12007);
and U17116 (N_17116,N_12840,N_14329);
and U17117 (N_17117,N_14713,N_15121);
nor U17118 (N_17118,N_15655,N_14706);
or U17119 (N_17119,N_15098,N_13269);
or U17120 (N_17120,N_14744,N_13675);
xnor U17121 (N_17121,N_13439,N_12271);
xor U17122 (N_17122,N_14085,N_14965);
nand U17123 (N_17123,N_13497,N_14409);
and U17124 (N_17124,N_13316,N_14804);
or U17125 (N_17125,N_13559,N_13970);
xor U17126 (N_17126,N_15320,N_15564);
nand U17127 (N_17127,N_13977,N_12397);
nand U17128 (N_17128,N_12862,N_15315);
nand U17129 (N_17129,N_12381,N_14033);
nor U17130 (N_17130,N_12478,N_14347);
or U17131 (N_17131,N_14746,N_12090);
nor U17132 (N_17132,N_14547,N_13103);
xnor U17133 (N_17133,N_15879,N_14791);
or U17134 (N_17134,N_12827,N_14859);
nor U17135 (N_17135,N_14727,N_15569);
nor U17136 (N_17136,N_12694,N_13120);
nand U17137 (N_17137,N_14605,N_13639);
or U17138 (N_17138,N_12288,N_12791);
xor U17139 (N_17139,N_12783,N_15957);
nor U17140 (N_17140,N_12915,N_15292);
xor U17141 (N_17141,N_15783,N_15666);
and U17142 (N_17142,N_12475,N_12314);
nand U17143 (N_17143,N_13136,N_13872);
xnor U17144 (N_17144,N_15528,N_14343);
or U17145 (N_17145,N_15864,N_15100);
xnor U17146 (N_17146,N_14312,N_14728);
and U17147 (N_17147,N_13377,N_12950);
or U17148 (N_17148,N_13040,N_15188);
xnor U17149 (N_17149,N_13372,N_13529);
and U17150 (N_17150,N_15983,N_12184);
nand U17151 (N_17151,N_13728,N_12446);
and U17152 (N_17152,N_14596,N_14976);
and U17153 (N_17153,N_15539,N_13153);
or U17154 (N_17154,N_12661,N_13053);
nor U17155 (N_17155,N_15313,N_12533);
and U17156 (N_17156,N_12129,N_14533);
nand U17157 (N_17157,N_12141,N_14527);
nor U17158 (N_17158,N_13952,N_13520);
xnor U17159 (N_17159,N_15713,N_12646);
and U17160 (N_17160,N_12916,N_13115);
or U17161 (N_17161,N_15219,N_12937);
or U17162 (N_17162,N_14855,N_15501);
nand U17163 (N_17163,N_15943,N_15134);
or U17164 (N_17164,N_15405,N_15012);
nand U17165 (N_17165,N_15034,N_15149);
nor U17166 (N_17166,N_13462,N_14414);
or U17167 (N_17167,N_15568,N_15686);
nor U17168 (N_17168,N_12774,N_14725);
and U17169 (N_17169,N_12576,N_13809);
nand U17170 (N_17170,N_12468,N_15744);
and U17171 (N_17171,N_15852,N_14161);
xnor U17172 (N_17172,N_15789,N_15953);
xnor U17173 (N_17173,N_14819,N_15268);
nand U17174 (N_17174,N_12158,N_12529);
nor U17175 (N_17175,N_13940,N_15063);
and U17176 (N_17176,N_15024,N_14534);
nand U17177 (N_17177,N_12900,N_15424);
xnor U17178 (N_17178,N_14418,N_14198);
xnor U17179 (N_17179,N_12677,N_13133);
nand U17180 (N_17180,N_15136,N_14186);
xnor U17181 (N_17181,N_12264,N_14117);
xnor U17182 (N_17182,N_14179,N_15057);
nor U17183 (N_17183,N_15205,N_12849);
and U17184 (N_17184,N_15336,N_15479);
or U17185 (N_17185,N_12687,N_14695);
nor U17186 (N_17186,N_15892,N_14008);
nand U17187 (N_17187,N_14615,N_13185);
and U17188 (N_17188,N_14651,N_13561);
nand U17189 (N_17189,N_15156,N_15263);
nand U17190 (N_17190,N_13408,N_13069);
or U17191 (N_17191,N_13368,N_12086);
and U17192 (N_17192,N_12493,N_15404);
xor U17193 (N_17193,N_12065,N_13922);
xnor U17194 (N_17194,N_12302,N_13754);
and U17195 (N_17195,N_12458,N_13073);
nand U17196 (N_17196,N_13765,N_15191);
nand U17197 (N_17197,N_12082,N_13958);
or U17198 (N_17198,N_14192,N_13631);
nand U17199 (N_17199,N_12127,N_13712);
nor U17200 (N_17200,N_15162,N_14096);
nand U17201 (N_17201,N_14926,N_13004);
and U17202 (N_17202,N_12347,N_12552);
and U17203 (N_17203,N_13950,N_15483);
nand U17204 (N_17204,N_15601,N_12775);
nor U17205 (N_17205,N_12787,N_14102);
xnor U17206 (N_17206,N_14552,N_14322);
xnor U17207 (N_17207,N_13234,N_15343);
and U17208 (N_17208,N_15688,N_12920);
or U17209 (N_17209,N_13485,N_12072);
nor U17210 (N_17210,N_15002,N_15626);
nor U17211 (N_17211,N_14415,N_14919);
or U17212 (N_17212,N_15105,N_15992);
nor U17213 (N_17213,N_14959,N_13463);
xnor U17214 (N_17214,N_15616,N_13250);
nor U17215 (N_17215,N_13460,N_12567);
or U17216 (N_17216,N_12407,N_12476);
xnor U17217 (N_17217,N_12759,N_13521);
nand U17218 (N_17218,N_14209,N_14433);
xnor U17219 (N_17219,N_13468,N_12378);
nor U17220 (N_17220,N_13085,N_12853);
nand U17221 (N_17221,N_15645,N_15771);
nand U17222 (N_17222,N_14157,N_15391);
or U17223 (N_17223,N_14724,N_14003);
xnor U17224 (N_17224,N_15118,N_13841);
or U17225 (N_17225,N_14472,N_15632);
nor U17226 (N_17226,N_15701,N_15705);
nand U17227 (N_17227,N_15692,N_15967);
nor U17228 (N_17228,N_14495,N_12995);
nor U17229 (N_17229,N_15768,N_13491);
xor U17230 (N_17230,N_12500,N_14376);
nand U17231 (N_17231,N_15209,N_13157);
xnor U17232 (N_17232,N_12208,N_14187);
and U17233 (N_17233,N_12913,N_12726);
and U17234 (N_17234,N_13411,N_13452);
or U17235 (N_17235,N_12510,N_13658);
nand U17236 (N_17236,N_12561,N_13548);
nand U17237 (N_17237,N_12391,N_15938);
nor U17238 (N_17238,N_14602,N_13565);
nor U17239 (N_17239,N_15809,N_13365);
nor U17240 (N_17240,N_14827,N_12881);
and U17241 (N_17241,N_13176,N_14249);
or U17242 (N_17242,N_12155,N_14325);
or U17243 (N_17243,N_12210,N_15471);
nand U17244 (N_17244,N_15059,N_13854);
and U17245 (N_17245,N_12329,N_12960);
nor U17246 (N_17246,N_14464,N_12486);
nor U17247 (N_17247,N_15897,N_13635);
nor U17248 (N_17248,N_15958,N_12994);
nand U17249 (N_17249,N_14128,N_12166);
and U17250 (N_17250,N_12867,N_13535);
xor U17251 (N_17251,N_12461,N_14201);
xor U17252 (N_17252,N_13394,N_13428);
nand U17253 (N_17253,N_12999,N_15577);
and U17254 (N_17254,N_15249,N_13493);
nand U17255 (N_17255,N_12297,N_14475);
nor U17256 (N_17256,N_15639,N_15971);
xnor U17257 (N_17257,N_14428,N_13397);
nor U17258 (N_17258,N_15703,N_15344);
xnor U17259 (N_17259,N_14304,N_12710);
nand U17260 (N_17260,N_12284,N_12230);
xor U17261 (N_17261,N_13431,N_14141);
and U17262 (N_17262,N_14638,N_14579);
nand U17263 (N_17263,N_14838,N_13016);
nand U17264 (N_17264,N_14715,N_13519);
and U17265 (N_17265,N_13591,N_15822);
nand U17266 (N_17266,N_13668,N_15649);
xnor U17267 (N_17267,N_13412,N_13050);
or U17268 (N_17268,N_15080,N_15359);
xor U17269 (N_17269,N_15891,N_14032);
nand U17270 (N_17270,N_14439,N_13384);
xnor U17271 (N_17271,N_15593,N_15288);
nand U17272 (N_17272,N_12524,N_12283);
nand U17273 (N_17273,N_12390,N_13351);
or U17274 (N_17274,N_15119,N_12728);
xnor U17275 (N_17275,N_12776,N_12046);
nand U17276 (N_17276,N_12022,N_14047);
and U17277 (N_17277,N_13290,N_12021);
or U17278 (N_17278,N_12002,N_12369);
nor U17279 (N_17279,N_14054,N_15113);
xor U17280 (N_17280,N_15615,N_13277);
nor U17281 (N_17281,N_15793,N_12405);
or U17282 (N_17282,N_12968,N_14629);
xnor U17283 (N_17283,N_13477,N_13708);
xnor U17284 (N_17284,N_14598,N_15923);
nor U17285 (N_17285,N_13933,N_13788);
or U17286 (N_17286,N_14743,N_13171);
or U17287 (N_17287,N_15622,N_14570);
nand U17288 (N_17288,N_12928,N_13141);
nand U17289 (N_17289,N_14426,N_12413);
xor U17290 (N_17290,N_13340,N_12041);
nor U17291 (N_17291,N_12432,N_12560);
nand U17292 (N_17292,N_13601,N_15702);
nor U17293 (N_17293,N_12412,N_12296);
or U17294 (N_17294,N_14862,N_12250);
or U17295 (N_17295,N_13731,N_13093);
and U17296 (N_17296,N_14747,N_12732);
nor U17297 (N_17297,N_15842,N_15140);
nor U17298 (N_17298,N_14095,N_13891);
or U17299 (N_17299,N_13710,N_12312);
or U17300 (N_17300,N_12149,N_15782);
xor U17301 (N_17301,N_14431,N_12956);
nand U17302 (N_17302,N_13851,N_14317);
xor U17303 (N_17303,N_14981,N_15727);
or U17304 (N_17304,N_13070,N_12383);
xor U17305 (N_17305,N_13370,N_12574);
nor U17306 (N_17306,N_12382,N_14685);
and U17307 (N_17307,N_14068,N_14476);
nand U17308 (N_17308,N_15812,N_14218);
nand U17309 (N_17309,N_14924,N_14024);
and U17310 (N_17310,N_14025,N_14384);
nand U17311 (N_17311,N_12893,N_14252);
nor U17312 (N_17312,N_12921,N_15873);
and U17313 (N_17313,N_14785,N_13980);
nor U17314 (N_17314,N_12696,N_15165);
xor U17315 (N_17315,N_14974,N_14930);
nand U17316 (N_17316,N_14909,N_15581);
and U17317 (N_17317,N_12167,N_14876);
and U17318 (N_17318,N_15328,N_15238);
nor U17319 (N_17319,N_13649,N_12045);
or U17320 (N_17320,N_12420,N_15733);
nand U17321 (N_17321,N_12684,N_13636);
xnor U17322 (N_17322,N_14752,N_14568);
xor U17323 (N_17323,N_14450,N_14119);
and U17324 (N_17324,N_14134,N_15767);
xor U17325 (N_17325,N_13604,N_13910);
xnor U17326 (N_17326,N_12227,N_13623);
nand U17327 (N_17327,N_15954,N_13379);
nand U17328 (N_17328,N_15371,N_14650);
or U17329 (N_17329,N_14446,N_15634);
or U17330 (N_17330,N_15554,N_13435);
or U17331 (N_17331,N_13965,N_14758);
xnor U17332 (N_17332,N_15618,N_13092);
nor U17333 (N_17333,N_14156,N_14419);
nand U17334 (N_17334,N_14497,N_12835);
nor U17335 (N_17335,N_12156,N_12258);
xor U17336 (N_17336,N_14633,N_15790);
or U17337 (N_17337,N_12024,N_12816);
or U17338 (N_17338,N_12265,N_15717);
and U17339 (N_17339,N_14865,N_14979);
and U17340 (N_17340,N_13188,N_13614);
or U17341 (N_17341,N_14262,N_13664);
nand U17342 (N_17342,N_12355,N_12823);
nor U17343 (N_17343,N_13892,N_15712);
nand U17344 (N_17344,N_15107,N_13244);
and U17345 (N_17345,N_15535,N_15926);
and U17346 (N_17346,N_13450,N_15096);
xor U17347 (N_17347,N_14359,N_13539);
xor U17348 (N_17348,N_12313,N_13312);
or U17349 (N_17349,N_15976,N_12175);
nand U17350 (N_17350,N_13427,N_13504);
nor U17351 (N_17351,N_13058,N_12214);
nand U17352 (N_17352,N_14694,N_13724);
nand U17353 (N_17353,N_12760,N_14067);
xor U17354 (N_17354,N_15538,N_14454);
or U17355 (N_17355,N_15732,N_15038);
and U17356 (N_17356,N_14189,N_14556);
or U17357 (N_17357,N_12162,N_13352);
nor U17358 (N_17358,N_14352,N_14379);
xor U17359 (N_17359,N_15242,N_12647);
or U17360 (N_17360,N_12579,N_12411);
and U17361 (N_17361,N_15251,N_12165);
nor U17362 (N_17362,N_12652,N_14016);
or U17363 (N_17363,N_15330,N_12586);
and U17364 (N_17364,N_13835,N_14381);
nor U17365 (N_17365,N_12442,N_15660);
or U17366 (N_17366,N_12918,N_12504);
or U17367 (N_17367,N_13948,N_12392);
and U17368 (N_17368,N_12255,N_15441);
and U17369 (N_17369,N_15827,N_12906);
and U17370 (N_17370,N_15917,N_14369);
nand U17371 (N_17371,N_15296,N_13076);
and U17372 (N_17372,N_14545,N_15553);
nor U17373 (N_17373,N_14231,N_12841);
and U17374 (N_17374,N_13173,N_12899);
or U17375 (N_17375,N_13299,N_13189);
nand U17376 (N_17376,N_14135,N_15236);
xor U17377 (N_17377,N_13376,N_14816);
xor U17378 (N_17378,N_13500,N_12276);
or U17379 (N_17379,N_14297,N_13071);
xnor U17380 (N_17380,N_15628,N_15327);
or U17381 (N_17381,N_15956,N_14079);
or U17382 (N_17382,N_14311,N_15453);
xnor U17383 (N_17383,N_15493,N_12590);
or U17384 (N_17384,N_13834,N_12522);
or U17385 (N_17385,N_13665,N_13813);
and U17386 (N_17386,N_14873,N_15306);
or U17387 (N_17387,N_15447,N_15168);
nor U17388 (N_17388,N_13576,N_15137);
and U17389 (N_17389,N_15164,N_15944);
or U17390 (N_17390,N_12528,N_14280);
and U17391 (N_17391,N_13418,N_14276);
xor U17392 (N_17392,N_12319,N_14256);
xnor U17393 (N_17393,N_13344,N_14473);
or U17394 (N_17394,N_12719,N_13116);
or U17395 (N_17395,N_12221,N_13147);
nand U17396 (N_17396,N_15186,N_12636);
or U17397 (N_17397,N_13317,N_12932);
or U17398 (N_17398,N_15456,N_12393);
nand U17399 (N_17399,N_12408,N_13245);
and U17400 (N_17400,N_15380,N_12685);
xor U17401 (N_17401,N_15582,N_15602);
nand U17402 (N_17402,N_14679,N_12583);
xnor U17403 (N_17403,N_12424,N_12170);
nor U17404 (N_17404,N_15886,N_14036);
or U17405 (N_17405,N_13893,N_14912);
or U17406 (N_17406,N_14314,N_12512);
nor U17407 (N_17407,N_14410,N_14449);
and U17408 (N_17408,N_12101,N_15434);
nand U17409 (N_17409,N_15144,N_12337);
xor U17410 (N_17410,N_14178,N_13223);
xor U17411 (N_17411,N_12751,N_15895);
and U17412 (N_17412,N_13832,N_13750);
or U17413 (N_17413,N_14714,N_14288);
and U17414 (N_17414,N_13072,N_15612);
xnor U17415 (N_17415,N_15758,N_12744);
or U17416 (N_17416,N_13923,N_14394);
nor U17417 (N_17417,N_13348,N_15011);
xor U17418 (N_17418,N_15382,N_15051);
or U17419 (N_17419,N_14914,N_14225);
nor U17420 (N_17420,N_13511,N_12342);
nand U17421 (N_17421,N_14499,N_12019);
and U17422 (N_17422,N_12351,N_13420);
and U17423 (N_17423,N_14565,N_13629);
nand U17424 (N_17424,N_15403,N_13168);
and U17425 (N_17425,N_14445,N_13655);
xnor U17426 (N_17426,N_15597,N_15385);
or U17427 (N_17427,N_12280,N_15560);
nor U17428 (N_17428,N_15849,N_13796);
or U17429 (N_17429,N_12293,N_13326);
nand U17430 (N_17430,N_15234,N_15550);
nand U17431 (N_17431,N_15847,N_13778);
nand U17432 (N_17432,N_12352,N_13971);
nand U17433 (N_17433,N_15126,N_13015);
or U17434 (N_17434,N_12790,N_13179);
xor U17435 (N_17435,N_12772,N_15457);
nand U17436 (N_17436,N_15881,N_13558);
or U17437 (N_17437,N_12870,N_14058);
nor U17438 (N_17438,N_13104,N_12456);
and U17439 (N_17439,N_14124,N_14931);
and U17440 (N_17440,N_15058,N_14538);
xor U17441 (N_17441,N_13611,N_13594);
nand U17442 (N_17442,N_14905,N_15007);
and U17443 (N_17443,N_13975,N_15245);
nor U17444 (N_17444,N_15832,N_14136);
nor U17445 (N_17445,N_12735,N_14332);
nand U17446 (N_17446,N_12975,N_12266);
nand U17447 (N_17447,N_12651,N_12553);
and U17448 (N_17448,N_12094,N_13595);
nor U17449 (N_17449,N_13208,N_15264);
nand U17450 (N_17450,N_15334,N_15866);
nor U17451 (N_17451,N_12761,N_13507);
xnor U17452 (N_17452,N_13403,N_13730);
nor U17453 (N_17453,N_13994,N_14453);
xnor U17454 (N_17454,N_12745,N_12452);
nand U17455 (N_17455,N_14639,N_15674);
xor U17456 (N_17456,N_15778,N_15826);
nand U17457 (N_17457,N_15613,N_15195);
xor U17458 (N_17458,N_14122,N_14672);
or U17459 (N_17459,N_14863,N_12398);
xor U17460 (N_17460,N_14123,N_12600);
or U17461 (N_17461,N_14140,N_12358);
nand U17462 (N_17462,N_14927,N_14794);
nor U17463 (N_17463,N_13705,N_12064);
nand U17464 (N_17464,N_14205,N_14388);
and U17465 (N_17465,N_15006,N_15884);
nor U17466 (N_17466,N_15094,N_14550);
or U17467 (N_17467,N_14575,N_14858);
or U17468 (N_17468,N_15229,N_14717);
and U17469 (N_17469,N_14530,N_13560);
xor U17470 (N_17470,N_15386,N_12124);
and U17471 (N_17471,N_15710,N_13803);
xnor U17472 (N_17472,N_14932,N_13634);
nand U17473 (N_17473,N_15816,N_14082);
xor U17474 (N_17474,N_13536,N_12730);
xnor U17475 (N_17475,N_12484,N_13187);
nor U17476 (N_17476,N_14593,N_13180);
or U17477 (N_17477,N_15217,N_12713);
nand U17478 (N_17478,N_12363,N_14796);
and U17479 (N_17479,N_14232,N_12338);
xnor U17480 (N_17480,N_12577,N_14808);
and U17481 (N_17481,N_13294,N_12768);
nor U17482 (N_17482,N_14257,N_15575);
nor U17483 (N_17483,N_13324,N_15070);
or U17484 (N_17484,N_14437,N_14240);
nor U17485 (N_17485,N_12075,N_15522);
nand U17486 (N_17486,N_13617,N_13361);
or U17487 (N_17487,N_13127,N_15785);
nand U17488 (N_17488,N_14963,N_13537);
nor U17489 (N_17489,N_13369,N_15450);
xnor U17490 (N_17490,N_15124,N_12807);
xnor U17491 (N_17491,N_13766,N_13845);
nor U17492 (N_17492,N_14048,N_12029);
nand U17493 (N_17493,N_13156,N_12904);
xor U17494 (N_17494,N_12481,N_12926);
xor U17495 (N_17495,N_14655,N_12691);
xor U17496 (N_17496,N_13953,N_15020);
xnor U17497 (N_17497,N_13406,N_13451);
nor U17498 (N_17498,N_13898,N_15806);
nor U17499 (N_17499,N_13976,N_14648);
nand U17500 (N_17500,N_15494,N_13219);
xnor U17501 (N_17501,N_14285,N_15931);
nand U17502 (N_17502,N_12451,N_15631);
nor U17503 (N_17503,N_12821,N_15325);
nor U17504 (N_17504,N_13306,N_14529);
nor U17505 (N_17505,N_14683,N_12739);
xnor U17506 (N_17506,N_14705,N_12460);
nand U17507 (N_17507,N_13931,N_12160);
xnor U17508 (N_17508,N_12620,N_12176);
nand U17509 (N_17509,N_12327,N_12125);
nand U17510 (N_17510,N_14941,N_15932);
or U17511 (N_17511,N_14159,N_15583);
nand U17512 (N_17512,N_15256,N_14035);
xnor U17513 (N_17513,N_15500,N_14657);
nor U17514 (N_17514,N_15570,N_12880);
nand U17515 (N_17515,N_14447,N_14197);
nor U17516 (N_17516,N_14344,N_15437);
nand U17517 (N_17517,N_15228,N_15662);
nand U17518 (N_17518,N_13857,N_14686);
nor U17519 (N_17519,N_12462,N_15837);
xnor U17520 (N_17520,N_15103,N_13247);
and U17521 (N_17521,N_15999,N_14697);
and U17522 (N_17522,N_13229,N_15843);
and U17523 (N_17523,N_12307,N_14374);
nand U17524 (N_17524,N_12133,N_15559);
or U17525 (N_17525,N_13099,N_15928);
nor U17526 (N_17526,N_14761,N_12399);
or U17527 (N_17527,N_14180,N_12929);
and U17528 (N_17528,N_15617,N_13486);
nand U17529 (N_17529,N_13043,N_14129);
nor U17530 (N_17530,N_13707,N_15197);
or U17531 (N_17531,N_14401,N_14030);
and U17532 (N_17532,N_15950,N_14039);
and U17533 (N_17533,N_13339,N_12020);
xor U17534 (N_17534,N_14448,N_14739);
nand U17535 (N_17535,N_14885,N_15889);
nand U17536 (N_17536,N_15802,N_15019);
nand U17537 (N_17537,N_13454,N_12777);
nand U17538 (N_17538,N_14676,N_15969);
or U17539 (N_17539,N_12142,N_13057);
nor U17540 (N_17540,N_15078,N_13243);
or U17541 (N_17541,N_13974,N_14090);
and U17542 (N_17542,N_12697,N_15099);
or U17543 (N_17543,N_12096,N_13593);
and U17544 (N_17544,N_15933,N_13096);
or U17545 (N_17545,N_12711,N_13661);
nor U17546 (N_17546,N_14824,N_13308);
and U17547 (N_17547,N_14457,N_14143);
or U17548 (N_17548,N_13749,N_13839);
or U17549 (N_17549,N_15604,N_14321);
or U17550 (N_17550,N_14908,N_15123);
nand U17551 (N_17551,N_14514,N_14829);
nand U17552 (N_17552,N_13321,N_14921);
xnor U17553 (N_17553,N_13585,N_15711);
xor U17554 (N_17554,N_14842,N_15606);
nor U17555 (N_17555,N_14104,N_15065);
xor U17556 (N_17556,N_14107,N_14799);
xnor U17557 (N_17557,N_15036,N_15698);
or U17558 (N_17558,N_14920,N_13575);
xnor U17559 (N_17559,N_14887,N_14652);
nand U17560 (N_17560,N_12071,N_14869);
or U17561 (N_17561,N_12737,N_12004);
nand U17562 (N_17562,N_12946,N_14622);
nor U17563 (N_17563,N_12515,N_12701);
or U17564 (N_17564,N_12385,N_13045);
xnor U17565 (N_17565,N_14248,N_15179);
nor U17566 (N_17566,N_14078,N_14182);
nand U17567 (N_17567,N_13353,N_12974);
xnor U17568 (N_17568,N_12985,N_12695);
and U17569 (N_17569,N_14903,N_14704);
nand U17570 (N_17570,N_14767,N_15644);
nand U17571 (N_17571,N_13191,N_12573);
or U17572 (N_17572,N_15760,N_13327);
nand U17573 (N_17573,N_13523,N_13828);
xor U17574 (N_17574,N_14784,N_14987);
xnor U17575 (N_17575,N_15795,N_15934);
nor U17576 (N_17576,N_12202,N_14677);
nand U17577 (N_17577,N_12134,N_13489);
nand U17578 (N_17578,N_14938,N_15241);
or U17579 (N_17579,N_15304,N_12067);
nor U17580 (N_17580,N_12808,N_13934);
and U17581 (N_17581,N_13666,N_12605);
nor U17582 (N_17582,N_13527,N_13844);
nand U17583 (N_17583,N_13883,N_15681);
or U17584 (N_17584,N_13769,N_13480);
xnor U17585 (N_17585,N_13183,N_12568);
and U17586 (N_17586,N_15751,N_14835);
xnor U17587 (N_17587,N_13404,N_13456);
or U17588 (N_17588,N_13003,N_13357);
nand U17589 (N_17589,N_14564,N_14087);
nor U17590 (N_17590,N_12865,N_12640);
or U17591 (N_17591,N_13777,N_13349);
or U17592 (N_17592,N_14998,N_15995);
nand U17593 (N_17593,N_14986,N_14874);
nand U17594 (N_17594,N_12649,N_13010);
xor U17595 (N_17595,N_14247,N_14014);
and U17596 (N_17596,N_14757,N_13138);
and U17597 (N_17597,N_14991,N_13047);
xnor U17598 (N_17598,N_13220,N_13979);
nand U17599 (N_17599,N_13876,N_14237);
xnor U17600 (N_17600,N_13469,N_15963);
xnor U17601 (N_17601,N_14610,N_12996);
and U17602 (N_17602,N_14413,N_14266);
nand U17603 (N_17603,N_13885,N_15547);
nand U17604 (N_17604,N_14729,N_12269);
xor U17605 (N_17605,N_13671,N_12860);
nand U17606 (N_17606,N_15202,N_15066);
nor U17607 (N_17607,N_15486,N_13270);
nand U17608 (N_17608,N_14452,N_15854);
xnor U17609 (N_17609,N_14356,N_13175);
xnor U17610 (N_17610,N_12693,N_15355);
nand U17611 (N_17611,N_15968,N_14239);
nor U17612 (N_17612,N_13954,N_12368);
xor U17613 (N_17613,N_12040,N_12150);
nand U17614 (N_17614,N_12272,N_15964);
nand U17615 (N_17615,N_14612,N_12631);
nor U17616 (N_17616,N_13557,N_15452);
nor U17617 (N_17617,N_15010,N_12545);
nor U17618 (N_17618,N_12431,N_15723);
or U17619 (N_17619,N_13949,N_13444);
and U17620 (N_17620,N_14662,N_12927);
nor U17621 (N_17621,N_14099,N_12277);
and U17622 (N_17622,N_12678,N_14204);
and U17623 (N_17623,N_15463,N_15859);
xor U17624 (N_17624,N_12406,N_12756);
and U17625 (N_17625,N_12705,N_14951);
nand U17626 (N_17626,N_14152,N_15284);
or U17627 (N_17627,N_12715,N_15032);
and U17628 (N_17628,N_12110,N_12618);
nand U17629 (N_17629,N_12234,N_15016);
or U17630 (N_17630,N_12237,N_13430);
or U17631 (N_17631,N_13283,N_12721);
nor U17632 (N_17632,N_13947,N_14155);
nor U17633 (N_17633,N_13235,N_14133);
or U17634 (N_17634,N_14294,N_15248);
or U17635 (N_17635,N_15041,N_12203);
and U17636 (N_17636,N_15520,N_12076);
or U17637 (N_17637,N_14877,N_13989);
or U17638 (N_17638,N_14883,N_14933);
and U17639 (N_17639,N_13943,N_14896);
and U17640 (N_17640,N_14181,N_12742);
or U17641 (N_17641,N_15408,N_15181);
or U17642 (N_17642,N_13434,N_15069);
or U17643 (N_17643,N_12242,N_13916);
nand U17644 (N_17644,N_14459,N_13424);
and U17645 (N_17645,N_12163,N_14734);
and U17646 (N_17646,N_12671,N_14491);
nand U17647 (N_17647,N_15233,N_13007);
or U17648 (N_17648,N_14977,N_14146);
nor U17649 (N_17649,N_13049,N_12514);
and U17650 (N_17650,N_13599,N_15955);
nand U17651 (N_17651,N_15345,N_12554);
and U17652 (N_17652,N_13698,N_15214);
xor U17653 (N_17653,N_12349,N_13362);
nor U17654 (N_17654,N_12118,N_12472);
and U17655 (N_17655,N_13059,N_14978);
nor U17656 (N_17656,N_13123,N_13271);
nand U17657 (N_17657,N_12998,N_14293);
nand U17658 (N_17658,N_13161,N_15764);
and U17659 (N_17659,N_14086,N_12741);
nand U17660 (N_17660,N_12923,N_14972);
xnor U17661 (N_17661,N_15541,N_15714);
or U17662 (N_17662,N_13062,N_15413);
xor U17663 (N_17663,N_13861,N_12991);
xnor U17664 (N_17664,N_12316,N_15621);
or U17665 (N_17665,N_12323,N_15255);
xnor U17666 (N_17666,N_15638,N_14630);
or U17667 (N_17667,N_14945,N_15272);
nor U17668 (N_17668,N_15643,N_15358);
nand U17669 (N_17669,N_13709,N_15573);
or U17670 (N_17670,N_14618,N_14040);
nand U17671 (N_17671,N_15741,N_14536);
or U17672 (N_17672,N_14617,N_14616);
or U17673 (N_17673,N_15435,N_13020);
or U17674 (N_17674,N_15056,N_15513);
xor U17675 (N_17675,N_12308,N_14670);
and U17676 (N_17676,N_12010,N_13569);
nand U17677 (N_17677,N_14631,N_15829);
or U17678 (N_17678,N_14736,N_13366);
nand U17679 (N_17679,N_13743,N_13380);
or U17680 (N_17680,N_14731,N_13240);
and U17681 (N_17681,N_13363,N_12016);
or U17682 (N_17682,N_15160,N_13919);
and U17683 (N_17683,N_13678,N_14176);
and U17684 (N_17684,N_13097,N_12120);
and U17685 (N_17685,N_15426,N_14733);
and U17686 (N_17686,N_13605,N_12753);
nor U17687 (N_17687,N_14576,N_14350);
nand U17688 (N_17688,N_14206,N_14265);
nor U17689 (N_17689,N_14089,N_12679);
and U17690 (N_17690,N_13514,N_14818);
or U17691 (N_17691,N_14505,N_14898);
and U17692 (N_17692,N_15223,N_15303);
nor U17693 (N_17693,N_13782,N_13988);
and U17694 (N_17694,N_12729,N_13083);
nor U17695 (N_17695,N_14425,N_12299);
xor U17696 (N_17696,N_15851,N_13066);
nand U17697 (N_17697,N_14771,N_14860);
and U17698 (N_17698,N_15387,N_14275);
xor U17699 (N_17699,N_12315,N_12311);
nor U17700 (N_17700,N_14839,N_14330);
xnor U17701 (N_17701,N_13723,N_13143);
nand U17702 (N_17702,N_13683,N_12801);
nor U17703 (N_17703,N_15247,N_13087);
or U17704 (N_17704,N_13964,N_15614);
nand U17705 (N_17705,N_13014,N_15206);
nand U17706 (N_17706,N_13482,N_13432);
nor U17707 (N_17707,N_14341,N_14427);
and U17708 (N_17708,N_14267,N_15015);
and U17709 (N_17709,N_12633,N_13300);
or U17710 (N_17710,N_13260,N_15704);
nand U17711 (N_17711,N_15270,N_15916);
and U17712 (N_17712,N_15863,N_14870);
xor U17713 (N_17713,N_15839,N_15476);
or U17714 (N_17714,N_12197,N_13198);
nor U17715 (N_17715,N_13081,N_14371);
nand U17716 (N_17716,N_13122,N_14151);
nor U17717 (N_17717,N_12609,N_12972);
nor U17718 (N_17718,N_13048,N_12121);
nor U17719 (N_17719,N_15319,N_15503);
xor U17720 (N_17720,N_15175,N_15537);
and U17721 (N_17721,N_12897,N_14532);
nor U17722 (N_17722,N_13155,N_15308);
and U17723 (N_17723,N_12032,N_13662);
or U17724 (N_17724,N_13481,N_12480);
xor U17725 (N_17725,N_12793,N_15042);
or U17726 (N_17726,N_13995,N_14241);
nand U17727 (N_17727,N_13144,N_14121);
nand U17728 (N_17728,N_15445,N_15982);
or U17729 (N_17729,N_13249,N_13667);
or U17730 (N_17730,N_13303,N_12635);
or U17731 (N_17731,N_14509,N_15389);
nor U17732 (N_17732,N_12669,N_13494);
xnor U17733 (N_17733,N_14864,N_14789);
or U17734 (N_17734,N_14053,N_15763);
and U17735 (N_17735,N_14990,N_14100);
or U17736 (N_17736,N_12371,N_13132);
nor U17737 (N_17737,N_14442,N_12842);
nand U17738 (N_17738,N_15362,N_13874);
and U17739 (N_17739,N_14324,N_15014);
xor U17740 (N_17740,N_15605,N_15695);
xnor U17741 (N_17741,N_12009,N_14640);
xnor U17742 (N_17742,N_13702,N_14199);
nor U17743 (N_17743,N_12704,N_14681);
xor U17744 (N_17744,N_14270,N_12023);
nor U17745 (N_17745,N_13255,N_12115);
or U17746 (N_17746,N_12740,N_13825);
nand U17747 (N_17747,N_12723,N_12935);
nor U17748 (N_17748,N_12708,N_13516);
nor U17749 (N_17749,N_13021,N_13748);
nand U17750 (N_17750,N_12204,N_12794);
nand U17751 (N_17751,N_13169,N_15050);
or U17752 (N_17752,N_13129,N_13145);
xnor U17753 (N_17753,N_13867,N_12275);
or U17754 (N_17754,N_12194,N_14601);
nor U17755 (N_17755,N_12006,N_12989);
nand U17756 (N_17756,N_13808,N_15548);
and U17757 (N_17757,N_12463,N_15446);
nor U17758 (N_17758,N_15549,N_14238);
and U17759 (N_17759,N_13533,N_15848);
and U17760 (N_17760,N_12965,N_12488);
and U17761 (N_17761,N_15792,N_15030);
and U17762 (N_17762,N_12223,N_15834);
xnor U17763 (N_17763,N_13195,N_13838);
nor U17764 (N_17764,N_14436,N_15314);
xnor U17765 (N_17765,N_15018,N_12239);
and U17766 (N_17766,N_15088,N_12060);
or U17767 (N_17767,N_15689,N_15130);
and U17768 (N_17768,N_12663,N_12376);
or U17769 (N_17769,N_13756,N_14666);
xnor U17770 (N_17770,N_13209,N_12341);
and U17771 (N_17771,N_12623,N_13333);
nor U17772 (N_17772,N_15885,N_15298);
or U17773 (N_17773,N_12109,N_13278);
xnor U17774 (N_17774,N_12883,N_15676);
or U17775 (N_17775,N_12043,N_13810);
nor U17776 (N_17776,N_13259,N_13550);
or U17777 (N_17777,N_15591,N_15132);
xnor U17778 (N_17778,N_13409,N_13286);
xor U17779 (N_17779,N_12930,N_14678);
nor U17780 (N_17780,N_14526,N_12364);
xnor U17781 (N_17781,N_15530,N_13107);
xor U17782 (N_17782,N_13733,N_15131);
nand U17783 (N_17783,N_14748,N_14691);
nand U17784 (N_17784,N_13531,N_15868);
nor U17785 (N_17785,N_14200,N_15572);
and U17786 (N_17786,N_13827,N_14710);
nor U17787 (N_17787,N_13643,N_14059);
and U17788 (N_17788,N_13446,N_13938);
and U17789 (N_17789,N_15153,N_15542);
xor U17790 (N_17790,N_15589,N_13747);
or U17791 (N_17791,N_15110,N_13113);
xnor U17792 (N_17792,N_15252,N_13987);
nor U17793 (N_17793,N_13307,N_12888);
nor U17794 (N_17794,N_13199,N_15388);
nand U17795 (N_17795,N_14936,N_13871);
xnor U17796 (N_17796,N_15761,N_13805);
and U17797 (N_17797,N_12909,N_12536);
and U17798 (N_17798,N_15630,N_13545);
xor U17799 (N_17799,N_15337,N_14654);
and U17800 (N_17800,N_13080,N_13101);
xnor U17801 (N_17801,N_14581,N_14516);
or U17802 (N_17802,N_15365,N_12262);
or U17803 (N_17803,N_12588,N_13926);
nand U17804 (N_17804,N_14554,N_14195);
nor U17805 (N_17805,N_13345,N_15603);
and U17806 (N_17806,N_12885,N_14011);
nand U17807 (N_17807,N_12178,N_15478);
and U17808 (N_17808,N_15867,N_14162);
and U17809 (N_17809,N_12489,N_13355);
or U17810 (N_17810,N_13830,N_12241);
nor U17811 (N_17811,N_13720,N_12310);
or U17812 (N_17812,N_13644,N_12091);
and U17813 (N_17813,N_15300,N_14814);
and U17814 (N_17814,N_15595,N_13859);
or U17815 (N_17815,N_12688,N_12940);
xor U17816 (N_17816,N_13149,N_12606);
or U17817 (N_17817,N_14599,N_15025);
and U17818 (N_17818,N_14969,N_14587);
nand U17819 (N_17819,N_13807,N_15997);
and U17820 (N_17820,N_15740,N_14253);
nor U17821 (N_17821,N_15524,N_13239);
xnor U17822 (N_17822,N_15089,N_12901);
or U17823 (N_17823,N_12389,N_12232);
nand U17824 (N_17824,N_14642,N_13856);
nand U17825 (N_17825,N_15451,N_12602);
nand U17826 (N_17826,N_14126,N_12814);
xnor U17827 (N_17827,N_13190,N_14797);
and U17828 (N_17828,N_13281,N_15914);
and U17829 (N_17829,N_13399,N_15919);
or U17830 (N_17830,N_14537,N_15280);
xor U17831 (N_17831,N_14775,N_15220);
xnor U17832 (N_17832,N_12428,N_14309);
and U17833 (N_17833,N_15882,N_14405);
xnor U17834 (N_17834,N_12199,N_13752);
nor U17835 (N_17835,N_12662,N_15187);
or U17836 (N_17836,N_14801,N_15664);
nand U17837 (N_17837,N_14590,N_15278);
nand U17838 (N_17838,N_13690,N_14684);
nand U17839 (N_17839,N_12287,N_13293);
xnor U17840 (N_17840,N_13628,N_12033);
or U17841 (N_17841,N_13150,N_13915);
nor U17842 (N_17842,N_13897,N_13822);
and U17843 (N_17843,N_15685,N_15533);
nor U17844 (N_17844,N_12048,N_15373);
nor U17845 (N_17845,N_13753,N_12656);
and U17846 (N_17846,N_14890,N_12981);
nand U17847 (N_17847,N_13554,N_12330);
nor U17848 (N_17848,N_12778,N_14402);
and U17849 (N_17849,N_14745,N_14975);
nor U17850 (N_17850,N_12078,N_15620);
nand U17851 (N_17851,N_14781,N_14962);
or U17852 (N_17852,N_15665,N_12809);
and U17853 (N_17853,N_15133,N_14578);
xnor U17854 (N_17854,N_15540,N_12702);
nor U17855 (N_17855,N_14093,N_14502);
nand U17856 (N_17856,N_12181,N_12154);
nand U17857 (N_17857,N_15161,N_14378);
and U17858 (N_17858,N_12733,N_15419);
xor U17859 (N_17859,N_12068,N_14671);
xor U17860 (N_17860,N_14759,N_15797);
and U17861 (N_17861,N_14416,N_14613);
xnor U17862 (N_17862,N_12621,N_15658);
nand U17863 (N_17863,N_12882,N_12550);
and U17864 (N_17864,N_15726,N_13483);
and U17865 (N_17865,N_13465,N_12543);
and U17866 (N_17866,N_15339,N_13886);
and U17867 (N_17867,N_13310,N_12982);
nand U17868 (N_17868,N_13632,N_14466);
or U17869 (N_17869,N_15948,N_12421);
xnor U17870 (N_17870,N_15093,N_13966);
or U17871 (N_17871,N_12059,N_13011);
xor U17872 (N_17872,N_13812,N_12217);
and U17873 (N_17873,N_14840,N_15072);
or U17874 (N_17874,N_13701,N_15361);
nand U17875 (N_17875,N_12106,N_13222);
nand U17876 (N_17876,N_12083,N_14940);
xor U17877 (N_17877,N_13973,N_15431);
nand U17878 (N_17878,N_13887,N_12970);
or U17879 (N_17879,N_15090,N_14307);
and U17880 (N_17880,N_13285,N_15516);
nand U17881 (N_17881,N_12638,N_15830);
nand U17882 (N_17882,N_12887,N_14608);
and U17883 (N_17883,N_12743,N_15749);
nand U17884 (N_17884,N_13760,N_14246);
xor U17885 (N_17885,N_15083,N_15282);
nand U17886 (N_17886,N_15250,N_12238);
nand U17887 (N_17887,N_13252,N_14043);
or U17888 (N_17888,N_13865,N_12457);
and U17889 (N_17889,N_12286,N_15988);
nand U17890 (N_17890,N_14830,N_13590);
or U17891 (N_17891,N_12601,N_12066);
nand U17892 (N_17892,N_15973,N_14982);
and U17893 (N_17893,N_15722,N_14906);
or U17894 (N_17894,N_14741,N_14260);
xnor U17895 (N_17895,N_13905,N_15872);
or U17896 (N_17896,N_14000,N_15076);
nand U17897 (N_17897,N_15600,N_15855);
and U17898 (N_17898,N_14664,N_15276);
nor U17899 (N_17899,N_14145,N_14658);
nand U17900 (N_17900,N_13653,N_12538);
and U17901 (N_17901,N_15004,N_14370);
or U17902 (N_17902,N_15979,N_15112);
nand U17903 (N_17903,N_12263,N_14723);
nand U17904 (N_17904,N_12593,N_15985);
xnor U17905 (N_17905,N_14386,N_13992);
nand U17906 (N_17906,N_12912,N_15896);
xor U17907 (N_17907,N_15898,N_14170);
xnor U17908 (N_17908,N_14190,N_15384);
nor U17909 (N_17909,N_12416,N_12645);
or U17910 (N_17910,N_15746,N_15900);
nor U17911 (N_17911,N_12948,N_12346);
nor U17912 (N_17912,N_13091,N_15787);
and U17913 (N_17913,N_15432,N_15724);
xnor U17914 (N_17914,N_14913,N_15273);
xnor U17915 (N_17915,N_12052,N_12604);
or U17916 (N_17916,N_13924,N_13108);
nor U17917 (N_17917,N_15192,N_12698);
xnor U17918 (N_17918,N_12714,N_15962);
nor U17919 (N_17919,N_13663,N_14061);
nor U17920 (N_17920,N_12589,N_14822);
xor U17921 (N_17921,N_14641,N_12924);
nand U17922 (N_17922,N_13740,N_13982);
nor U17923 (N_17923,N_12863,N_13946);
nand U17924 (N_17924,N_13334,N_12235);
xnor U17925 (N_17925,N_15719,N_15392);
and U17926 (N_17926,N_15587,N_14551);
or U17927 (N_17927,N_12207,N_13881);
or U17928 (N_17928,N_13582,N_13146);
nand U17929 (N_17929,N_14845,N_14160);
xor U17930 (N_17930,N_13985,N_15395);
nor U17931 (N_17931,N_13863,N_12815);
nor U17932 (N_17932,N_13118,N_14326);
xnor U17933 (N_17933,N_15182,N_12147);
or U17934 (N_17934,N_14754,N_12304);
xor U17935 (N_17935,N_13082,N_13633);
xnor U17936 (N_17936,N_13466,N_12061);
xnor U17937 (N_17937,N_12177,N_15449);
nand U17938 (N_17938,N_14383,N_13019);
or U17939 (N_17939,N_15350,N_15641);
or U17940 (N_17940,N_14773,N_14730);
nand U17941 (N_17941,N_13496,N_15227);
xor U17942 (N_17942,N_15592,N_13022);
nor U17943 (N_17943,N_14588,N_12444);
nor U17944 (N_17944,N_14357,N_14798);
and U17945 (N_17945,N_15266,N_12440);
xnor U17946 (N_17946,N_14834,N_12474);
nand U17947 (N_17947,N_13410,N_13464);
xor U17948 (N_17948,N_13126,N_15086);
nand U17949 (N_17949,N_13124,N_15716);
xnor U17950 (N_17950,N_14092,N_12547);
nor U17951 (N_17951,N_14065,N_15647);
nor U17952 (N_17952,N_13001,N_14219);
or U17953 (N_17953,N_12575,N_12558);
nand U17954 (N_17954,N_13218,N_14603);
nand U17955 (N_17955,N_12599,N_13347);
nor U17956 (N_17956,N_15261,N_13038);
or U17957 (N_17957,N_15482,N_12252);
and U17958 (N_17958,N_12143,N_14856);
xnor U17959 (N_17959,N_15745,N_12192);
xnor U17960 (N_17960,N_13917,N_13393);
nand U17961 (N_17961,N_14028,N_14621);
nand U17962 (N_17962,N_15412,N_13909);
and U17963 (N_17963,N_12495,N_13894);
and U17964 (N_17964,N_14274,N_15352);
or U17965 (N_17965,N_15211,N_14470);
and U17966 (N_17966,N_14188,N_15990);
xor U17967 (N_17967,N_14768,N_13615);
xnor U17968 (N_17968,N_12240,N_13619);
nor U17969 (N_17969,N_13121,N_14852);
xor U17970 (N_17970,N_14879,N_12598);
xnor U17971 (N_17971,N_13719,N_15239);
or U17972 (N_17972,N_13878,N_12248);
xnor U17973 (N_17973,N_12798,N_15786);
nand U17974 (N_17974,N_15402,N_13847);
nand U17975 (N_17975,N_12117,N_15363);
or U17976 (N_17976,N_15364,N_12945);
nor U17977 (N_17977,N_12624,N_12875);
xor U17978 (N_17978,N_15532,N_12565);
nor U17979 (N_17979,N_13642,N_14778);
or U17980 (N_17980,N_13416,N_14718);
nand U17981 (N_17981,N_12123,N_12746);
xnor U17982 (N_17982,N_12603,N_12098);
and U17983 (N_17983,N_12335,N_13503);
xnor U17984 (N_17984,N_14971,N_13475);
nor U17985 (N_17985,N_15347,N_14644);
nand U17986 (N_17986,N_15791,N_14103);
and U17987 (N_17987,N_14217,N_12490);
nor U17988 (N_17988,N_13600,N_15876);
nand U17989 (N_17989,N_13646,N_15906);
and U17990 (N_17990,N_15201,N_13358);
or U17991 (N_17991,N_14108,N_14540);
or U17992 (N_17992,N_14980,N_12572);
and U17993 (N_17993,N_12015,N_13233);
nor U17994 (N_17994,N_13313,N_15871);
or U17995 (N_17995,N_14300,N_14013);
or U17996 (N_17996,N_15683,N_12987);
xnor U17997 (N_17997,N_14235,N_13763);
xnor U17998 (N_17998,N_13616,N_14756);
nand U17999 (N_17999,N_15409,N_13544);
xor U18000 (N_18000,N_15085,N_15263);
nor U18001 (N_18001,N_14150,N_14397);
nand U18002 (N_18002,N_12426,N_15125);
or U18003 (N_18003,N_15870,N_13529);
nand U18004 (N_18004,N_12458,N_15805);
and U18005 (N_18005,N_13992,N_12374);
nand U18006 (N_18006,N_12537,N_15316);
nor U18007 (N_18007,N_12946,N_15695);
nand U18008 (N_18008,N_14322,N_13846);
nand U18009 (N_18009,N_12218,N_13525);
and U18010 (N_18010,N_15651,N_13253);
xnor U18011 (N_18011,N_15498,N_12875);
xnor U18012 (N_18012,N_15045,N_13080);
or U18013 (N_18013,N_13447,N_15816);
or U18014 (N_18014,N_13204,N_13760);
xnor U18015 (N_18015,N_15904,N_12593);
xor U18016 (N_18016,N_14554,N_14175);
or U18017 (N_18017,N_14467,N_15775);
and U18018 (N_18018,N_14399,N_14162);
and U18019 (N_18019,N_15552,N_14665);
xnor U18020 (N_18020,N_13661,N_14176);
nand U18021 (N_18021,N_12489,N_14238);
xnor U18022 (N_18022,N_12956,N_15868);
and U18023 (N_18023,N_15348,N_15141);
nand U18024 (N_18024,N_12020,N_12968);
or U18025 (N_18025,N_14277,N_15158);
or U18026 (N_18026,N_14672,N_15328);
and U18027 (N_18027,N_15164,N_15134);
nor U18028 (N_18028,N_14596,N_12056);
nor U18029 (N_18029,N_13401,N_13297);
nor U18030 (N_18030,N_14031,N_15014);
nand U18031 (N_18031,N_13985,N_12220);
or U18032 (N_18032,N_12136,N_14863);
xor U18033 (N_18033,N_13519,N_13933);
xor U18034 (N_18034,N_14649,N_12145);
nor U18035 (N_18035,N_14921,N_14653);
and U18036 (N_18036,N_12448,N_14471);
xor U18037 (N_18037,N_13920,N_15963);
or U18038 (N_18038,N_13400,N_12728);
nand U18039 (N_18039,N_12188,N_14467);
nand U18040 (N_18040,N_15144,N_15692);
nand U18041 (N_18041,N_14949,N_14879);
nor U18042 (N_18042,N_12089,N_14587);
and U18043 (N_18043,N_15558,N_12207);
nor U18044 (N_18044,N_14843,N_13278);
xnor U18045 (N_18045,N_14006,N_14923);
nand U18046 (N_18046,N_12790,N_12475);
nand U18047 (N_18047,N_14250,N_15128);
xor U18048 (N_18048,N_13310,N_12127);
xnor U18049 (N_18049,N_12778,N_13365);
nor U18050 (N_18050,N_15577,N_15058);
nor U18051 (N_18051,N_13063,N_14411);
nand U18052 (N_18052,N_15355,N_12231);
or U18053 (N_18053,N_14372,N_15908);
xnor U18054 (N_18054,N_13212,N_12030);
nand U18055 (N_18055,N_12885,N_13915);
xor U18056 (N_18056,N_13122,N_14932);
and U18057 (N_18057,N_13814,N_14252);
nor U18058 (N_18058,N_12337,N_12886);
and U18059 (N_18059,N_13934,N_13442);
or U18060 (N_18060,N_12878,N_12244);
or U18061 (N_18061,N_12589,N_12782);
nand U18062 (N_18062,N_13144,N_13110);
nor U18063 (N_18063,N_12938,N_15838);
nand U18064 (N_18064,N_15147,N_13442);
or U18065 (N_18065,N_13402,N_14645);
nor U18066 (N_18066,N_14663,N_12039);
xor U18067 (N_18067,N_12785,N_15070);
or U18068 (N_18068,N_12994,N_12535);
nor U18069 (N_18069,N_14515,N_14317);
nor U18070 (N_18070,N_13383,N_12706);
nor U18071 (N_18071,N_14131,N_13250);
or U18072 (N_18072,N_12276,N_14017);
nor U18073 (N_18073,N_15588,N_12705);
nor U18074 (N_18074,N_14256,N_13820);
or U18075 (N_18075,N_12316,N_15298);
nand U18076 (N_18076,N_15978,N_15567);
nand U18077 (N_18077,N_12994,N_15155);
and U18078 (N_18078,N_14366,N_13557);
nor U18079 (N_18079,N_12314,N_14026);
nand U18080 (N_18080,N_12637,N_12058);
xnor U18081 (N_18081,N_13505,N_15543);
xnor U18082 (N_18082,N_14406,N_14254);
and U18083 (N_18083,N_13111,N_14652);
xor U18084 (N_18084,N_12472,N_15368);
and U18085 (N_18085,N_13199,N_13222);
and U18086 (N_18086,N_15390,N_14322);
xnor U18087 (N_18087,N_12601,N_13886);
nor U18088 (N_18088,N_14289,N_13392);
or U18089 (N_18089,N_13809,N_12925);
or U18090 (N_18090,N_13454,N_12782);
and U18091 (N_18091,N_12172,N_13275);
or U18092 (N_18092,N_12138,N_13891);
nor U18093 (N_18093,N_14134,N_14603);
xor U18094 (N_18094,N_14306,N_12157);
xor U18095 (N_18095,N_15411,N_15652);
nand U18096 (N_18096,N_13122,N_15143);
xor U18097 (N_18097,N_12921,N_13760);
or U18098 (N_18098,N_12639,N_13320);
and U18099 (N_18099,N_12156,N_13635);
nor U18100 (N_18100,N_13406,N_15588);
xnor U18101 (N_18101,N_15954,N_15019);
nor U18102 (N_18102,N_15506,N_14058);
and U18103 (N_18103,N_12961,N_12416);
nand U18104 (N_18104,N_12015,N_13395);
and U18105 (N_18105,N_13919,N_12740);
nor U18106 (N_18106,N_12391,N_13587);
nand U18107 (N_18107,N_13138,N_14156);
or U18108 (N_18108,N_13889,N_13802);
and U18109 (N_18109,N_15540,N_13051);
or U18110 (N_18110,N_12865,N_14313);
nor U18111 (N_18111,N_12745,N_12157);
or U18112 (N_18112,N_12250,N_14261);
nor U18113 (N_18113,N_13991,N_12161);
xnor U18114 (N_18114,N_12845,N_12091);
and U18115 (N_18115,N_14870,N_13098);
nand U18116 (N_18116,N_12890,N_12123);
nor U18117 (N_18117,N_15005,N_15023);
nand U18118 (N_18118,N_15444,N_14234);
nand U18119 (N_18119,N_14975,N_14987);
nand U18120 (N_18120,N_14744,N_15458);
or U18121 (N_18121,N_12611,N_14844);
xor U18122 (N_18122,N_14388,N_14732);
xor U18123 (N_18123,N_14820,N_13574);
nor U18124 (N_18124,N_14754,N_15440);
and U18125 (N_18125,N_14430,N_14403);
and U18126 (N_18126,N_15915,N_14193);
nor U18127 (N_18127,N_15792,N_15759);
and U18128 (N_18128,N_15109,N_15708);
nor U18129 (N_18129,N_12647,N_12846);
nor U18130 (N_18130,N_15061,N_12248);
or U18131 (N_18131,N_14302,N_13576);
nor U18132 (N_18132,N_15220,N_14792);
nand U18133 (N_18133,N_13253,N_14814);
or U18134 (N_18134,N_14773,N_12840);
and U18135 (N_18135,N_12748,N_13033);
nand U18136 (N_18136,N_15696,N_13538);
and U18137 (N_18137,N_15761,N_14390);
nand U18138 (N_18138,N_14655,N_15363);
and U18139 (N_18139,N_12470,N_15640);
and U18140 (N_18140,N_14358,N_12235);
nor U18141 (N_18141,N_15253,N_15591);
or U18142 (N_18142,N_14733,N_12495);
xor U18143 (N_18143,N_12250,N_13567);
nor U18144 (N_18144,N_15709,N_12035);
xor U18145 (N_18145,N_12861,N_12216);
nor U18146 (N_18146,N_14132,N_15734);
nand U18147 (N_18147,N_14220,N_13824);
nand U18148 (N_18148,N_14341,N_15136);
or U18149 (N_18149,N_13230,N_13329);
nor U18150 (N_18150,N_12344,N_14173);
xor U18151 (N_18151,N_14153,N_15005);
nand U18152 (N_18152,N_15886,N_15781);
and U18153 (N_18153,N_13366,N_13965);
xnor U18154 (N_18154,N_15243,N_14581);
or U18155 (N_18155,N_15148,N_13115);
nand U18156 (N_18156,N_15624,N_12442);
nor U18157 (N_18157,N_12343,N_14867);
nand U18158 (N_18158,N_15773,N_14622);
nand U18159 (N_18159,N_12064,N_15365);
or U18160 (N_18160,N_12434,N_14758);
xnor U18161 (N_18161,N_12465,N_14939);
and U18162 (N_18162,N_13707,N_12294);
xnor U18163 (N_18163,N_14515,N_15065);
and U18164 (N_18164,N_12172,N_14071);
nor U18165 (N_18165,N_12329,N_14268);
xnor U18166 (N_18166,N_14560,N_14542);
nand U18167 (N_18167,N_13951,N_15663);
and U18168 (N_18168,N_14310,N_15141);
nor U18169 (N_18169,N_14226,N_15224);
nor U18170 (N_18170,N_14610,N_15104);
nand U18171 (N_18171,N_15591,N_13290);
xnor U18172 (N_18172,N_15770,N_12841);
xnor U18173 (N_18173,N_12603,N_15962);
or U18174 (N_18174,N_13979,N_12024);
xor U18175 (N_18175,N_14931,N_13306);
and U18176 (N_18176,N_14535,N_12874);
or U18177 (N_18177,N_13792,N_14259);
or U18178 (N_18178,N_13911,N_13848);
xor U18179 (N_18179,N_14486,N_12951);
nand U18180 (N_18180,N_13535,N_12515);
and U18181 (N_18181,N_12150,N_12301);
and U18182 (N_18182,N_15275,N_15352);
nor U18183 (N_18183,N_15429,N_13034);
and U18184 (N_18184,N_12520,N_14321);
and U18185 (N_18185,N_15469,N_12391);
nor U18186 (N_18186,N_15132,N_13215);
or U18187 (N_18187,N_14684,N_15192);
nor U18188 (N_18188,N_14187,N_15600);
or U18189 (N_18189,N_12519,N_12415);
nand U18190 (N_18190,N_15234,N_12266);
or U18191 (N_18191,N_15800,N_13179);
nor U18192 (N_18192,N_13633,N_14575);
or U18193 (N_18193,N_13068,N_14131);
nand U18194 (N_18194,N_15810,N_14912);
and U18195 (N_18195,N_15423,N_15666);
xor U18196 (N_18196,N_13525,N_15103);
nor U18197 (N_18197,N_12005,N_13243);
nand U18198 (N_18198,N_13692,N_14266);
or U18199 (N_18199,N_14901,N_13558);
xor U18200 (N_18200,N_12816,N_15778);
xor U18201 (N_18201,N_15519,N_12482);
nor U18202 (N_18202,N_13386,N_15075);
nand U18203 (N_18203,N_14220,N_13992);
xor U18204 (N_18204,N_12162,N_13508);
nand U18205 (N_18205,N_13312,N_15507);
and U18206 (N_18206,N_12769,N_15919);
or U18207 (N_18207,N_14314,N_15994);
and U18208 (N_18208,N_14628,N_15269);
and U18209 (N_18209,N_15780,N_13583);
nor U18210 (N_18210,N_13082,N_13590);
nor U18211 (N_18211,N_12100,N_15329);
nor U18212 (N_18212,N_14733,N_13397);
or U18213 (N_18213,N_14420,N_12369);
and U18214 (N_18214,N_15781,N_14116);
nor U18215 (N_18215,N_14584,N_13018);
and U18216 (N_18216,N_13937,N_12003);
nor U18217 (N_18217,N_12900,N_14980);
or U18218 (N_18218,N_13272,N_14608);
and U18219 (N_18219,N_15784,N_15490);
nor U18220 (N_18220,N_13437,N_15819);
xnor U18221 (N_18221,N_13112,N_12273);
and U18222 (N_18222,N_12242,N_14787);
and U18223 (N_18223,N_12642,N_13039);
or U18224 (N_18224,N_13149,N_14569);
nand U18225 (N_18225,N_14273,N_12727);
nor U18226 (N_18226,N_13963,N_14518);
or U18227 (N_18227,N_15114,N_13590);
and U18228 (N_18228,N_13484,N_14322);
nand U18229 (N_18229,N_13198,N_12140);
nor U18230 (N_18230,N_15582,N_14289);
nand U18231 (N_18231,N_13278,N_13832);
or U18232 (N_18232,N_15555,N_14598);
nand U18233 (N_18233,N_14335,N_15828);
xnor U18234 (N_18234,N_14354,N_13115);
xor U18235 (N_18235,N_12373,N_12689);
nor U18236 (N_18236,N_13878,N_12324);
nand U18237 (N_18237,N_14890,N_14866);
or U18238 (N_18238,N_13297,N_12842);
xor U18239 (N_18239,N_12833,N_14943);
nor U18240 (N_18240,N_12913,N_12633);
nand U18241 (N_18241,N_12407,N_12061);
nor U18242 (N_18242,N_14223,N_14495);
xnor U18243 (N_18243,N_12173,N_13859);
nor U18244 (N_18244,N_13255,N_12139);
or U18245 (N_18245,N_14447,N_13950);
and U18246 (N_18246,N_15737,N_12424);
or U18247 (N_18247,N_15784,N_14763);
nor U18248 (N_18248,N_12691,N_15733);
nor U18249 (N_18249,N_12188,N_13880);
and U18250 (N_18250,N_15590,N_13106);
xor U18251 (N_18251,N_14873,N_15996);
or U18252 (N_18252,N_14017,N_13345);
nand U18253 (N_18253,N_13994,N_13032);
xor U18254 (N_18254,N_15829,N_15753);
nand U18255 (N_18255,N_12005,N_13179);
xor U18256 (N_18256,N_14112,N_12047);
or U18257 (N_18257,N_12230,N_13661);
and U18258 (N_18258,N_14159,N_15469);
xor U18259 (N_18259,N_12499,N_14813);
and U18260 (N_18260,N_13224,N_12046);
or U18261 (N_18261,N_14890,N_15462);
nor U18262 (N_18262,N_14932,N_13901);
xnor U18263 (N_18263,N_12048,N_14446);
nand U18264 (N_18264,N_14776,N_15336);
nand U18265 (N_18265,N_15362,N_13612);
or U18266 (N_18266,N_12972,N_14484);
or U18267 (N_18267,N_13716,N_13867);
xnor U18268 (N_18268,N_12227,N_13106);
nand U18269 (N_18269,N_12068,N_15018);
nor U18270 (N_18270,N_14885,N_15773);
or U18271 (N_18271,N_12659,N_14700);
xnor U18272 (N_18272,N_12141,N_14465);
and U18273 (N_18273,N_12064,N_14053);
or U18274 (N_18274,N_13174,N_14659);
nor U18275 (N_18275,N_13452,N_15102);
or U18276 (N_18276,N_15128,N_15075);
xor U18277 (N_18277,N_13032,N_14880);
and U18278 (N_18278,N_14980,N_13672);
nor U18279 (N_18279,N_13181,N_14575);
or U18280 (N_18280,N_13376,N_15972);
nor U18281 (N_18281,N_12450,N_13036);
nand U18282 (N_18282,N_12942,N_15216);
nand U18283 (N_18283,N_13934,N_12567);
and U18284 (N_18284,N_15211,N_12613);
nor U18285 (N_18285,N_15476,N_14489);
or U18286 (N_18286,N_15719,N_14747);
xnor U18287 (N_18287,N_12611,N_14377);
nor U18288 (N_18288,N_14233,N_15546);
and U18289 (N_18289,N_15094,N_12518);
nand U18290 (N_18290,N_14948,N_12945);
xor U18291 (N_18291,N_15983,N_14244);
nor U18292 (N_18292,N_13398,N_15094);
nor U18293 (N_18293,N_14811,N_12760);
and U18294 (N_18294,N_15297,N_13250);
and U18295 (N_18295,N_14290,N_14137);
nor U18296 (N_18296,N_13884,N_12037);
xor U18297 (N_18297,N_15220,N_12584);
xor U18298 (N_18298,N_13300,N_13541);
nand U18299 (N_18299,N_15052,N_12569);
xor U18300 (N_18300,N_15654,N_15173);
nor U18301 (N_18301,N_15745,N_12450);
or U18302 (N_18302,N_13700,N_12003);
or U18303 (N_18303,N_13134,N_13111);
nor U18304 (N_18304,N_15957,N_12222);
xor U18305 (N_18305,N_13018,N_14179);
nor U18306 (N_18306,N_12402,N_14706);
nor U18307 (N_18307,N_13503,N_14048);
or U18308 (N_18308,N_13066,N_12749);
nor U18309 (N_18309,N_15904,N_13828);
or U18310 (N_18310,N_12825,N_12543);
xor U18311 (N_18311,N_13360,N_15110);
xnor U18312 (N_18312,N_15648,N_14392);
or U18313 (N_18313,N_14384,N_14922);
xor U18314 (N_18314,N_13213,N_12668);
and U18315 (N_18315,N_13811,N_15142);
nor U18316 (N_18316,N_15638,N_14635);
or U18317 (N_18317,N_14733,N_15403);
and U18318 (N_18318,N_13000,N_12991);
and U18319 (N_18319,N_15822,N_14626);
nand U18320 (N_18320,N_13453,N_14743);
or U18321 (N_18321,N_15148,N_15416);
nor U18322 (N_18322,N_12875,N_13464);
xnor U18323 (N_18323,N_12090,N_14111);
or U18324 (N_18324,N_15870,N_12152);
or U18325 (N_18325,N_13822,N_13585);
nand U18326 (N_18326,N_12449,N_14599);
or U18327 (N_18327,N_12007,N_14178);
or U18328 (N_18328,N_15109,N_14527);
and U18329 (N_18329,N_12832,N_14438);
xor U18330 (N_18330,N_12680,N_15514);
nand U18331 (N_18331,N_13700,N_12165);
xor U18332 (N_18332,N_13300,N_14509);
xnor U18333 (N_18333,N_15228,N_14508);
nand U18334 (N_18334,N_12952,N_15411);
nand U18335 (N_18335,N_12714,N_12439);
or U18336 (N_18336,N_14484,N_14102);
xor U18337 (N_18337,N_15136,N_15840);
or U18338 (N_18338,N_12736,N_12352);
or U18339 (N_18339,N_14730,N_15732);
nand U18340 (N_18340,N_13425,N_13100);
nor U18341 (N_18341,N_15467,N_12278);
or U18342 (N_18342,N_12649,N_13187);
or U18343 (N_18343,N_12326,N_12064);
xor U18344 (N_18344,N_14184,N_15542);
and U18345 (N_18345,N_12408,N_14337);
or U18346 (N_18346,N_14933,N_14490);
or U18347 (N_18347,N_12898,N_15972);
nor U18348 (N_18348,N_12274,N_13978);
xor U18349 (N_18349,N_15198,N_14557);
nor U18350 (N_18350,N_12868,N_14323);
nand U18351 (N_18351,N_15715,N_15263);
nand U18352 (N_18352,N_12555,N_12156);
xor U18353 (N_18353,N_14941,N_13238);
and U18354 (N_18354,N_13547,N_12661);
xnor U18355 (N_18355,N_15104,N_12436);
or U18356 (N_18356,N_13287,N_12420);
nor U18357 (N_18357,N_14920,N_12378);
nand U18358 (N_18358,N_13660,N_12676);
nor U18359 (N_18359,N_13136,N_15352);
or U18360 (N_18360,N_13518,N_15159);
or U18361 (N_18361,N_14710,N_12878);
and U18362 (N_18362,N_13576,N_12976);
xnor U18363 (N_18363,N_12798,N_13497);
or U18364 (N_18364,N_12780,N_12593);
nand U18365 (N_18365,N_12678,N_14015);
nor U18366 (N_18366,N_12604,N_15904);
nor U18367 (N_18367,N_13894,N_14606);
and U18368 (N_18368,N_14295,N_15132);
nand U18369 (N_18369,N_14001,N_15012);
nor U18370 (N_18370,N_15824,N_15889);
and U18371 (N_18371,N_13569,N_12074);
nand U18372 (N_18372,N_15886,N_15815);
nor U18373 (N_18373,N_13536,N_13153);
nor U18374 (N_18374,N_14073,N_12741);
or U18375 (N_18375,N_14823,N_13835);
xor U18376 (N_18376,N_14896,N_12778);
or U18377 (N_18377,N_12260,N_13404);
xor U18378 (N_18378,N_14689,N_12792);
or U18379 (N_18379,N_15340,N_15198);
xor U18380 (N_18380,N_14215,N_15675);
xnor U18381 (N_18381,N_13385,N_13923);
nand U18382 (N_18382,N_14421,N_12221);
nor U18383 (N_18383,N_14524,N_13869);
xnor U18384 (N_18384,N_13559,N_15402);
nand U18385 (N_18385,N_13617,N_12516);
xnor U18386 (N_18386,N_13331,N_15219);
xor U18387 (N_18387,N_15927,N_12105);
xor U18388 (N_18388,N_15251,N_12333);
or U18389 (N_18389,N_15614,N_13809);
nand U18390 (N_18390,N_13081,N_15527);
xor U18391 (N_18391,N_15228,N_14929);
xor U18392 (N_18392,N_12530,N_15590);
or U18393 (N_18393,N_14252,N_12701);
xor U18394 (N_18394,N_12025,N_12072);
or U18395 (N_18395,N_15230,N_14948);
xnor U18396 (N_18396,N_15257,N_15076);
and U18397 (N_18397,N_12128,N_12874);
and U18398 (N_18398,N_14819,N_15748);
or U18399 (N_18399,N_14542,N_15298);
xnor U18400 (N_18400,N_15221,N_12731);
xor U18401 (N_18401,N_15162,N_13400);
xnor U18402 (N_18402,N_15152,N_15506);
nand U18403 (N_18403,N_12382,N_13705);
and U18404 (N_18404,N_15056,N_12219);
xor U18405 (N_18405,N_15439,N_14629);
nand U18406 (N_18406,N_15369,N_15525);
nor U18407 (N_18407,N_14086,N_13395);
and U18408 (N_18408,N_14653,N_12158);
xnor U18409 (N_18409,N_12464,N_12535);
and U18410 (N_18410,N_13670,N_14854);
nand U18411 (N_18411,N_13215,N_15841);
or U18412 (N_18412,N_14412,N_14517);
or U18413 (N_18413,N_15100,N_15872);
or U18414 (N_18414,N_14262,N_14970);
nor U18415 (N_18415,N_14233,N_15431);
nand U18416 (N_18416,N_14961,N_13205);
and U18417 (N_18417,N_15870,N_13201);
xnor U18418 (N_18418,N_15406,N_15224);
or U18419 (N_18419,N_13052,N_12840);
or U18420 (N_18420,N_14122,N_12210);
nand U18421 (N_18421,N_12617,N_15205);
xnor U18422 (N_18422,N_14774,N_13421);
xnor U18423 (N_18423,N_14303,N_15008);
or U18424 (N_18424,N_15663,N_13457);
nor U18425 (N_18425,N_12051,N_14520);
nand U18426 (N_18426,N_14172,N_14612);
nor U18427 (N_18427,N_12375,N_12019);
and U18428 (N_18428,N_15782,N_15176);
xor U18429 (N_18429,N_15748,N_14123);
nand U18430 (N_18430,N_12934,N_14977);
xnor U18431 (N_18431,N_15107,N_12335);
and U18432 (N_18432,N_12035,N_14742);
or U18433 (N_18433,N_15563,N_12998);
nand U18434 (N_18434,N_15341,N_15381);
or U18435 (N_18435,N_14219,N_15630);
nor U18436 (N_18436,N_14801,N_12718);
or U18437 (N_18437,N_14369,N_15518);
or U18438 (N_18438,N_12610,N_13531);
nor U18439 (N_18439,N_14588,N_12036);
nand U18440 (N_18440,N_15001,N_14828);
or U18441 (N_18441,N_15309,N_13173);
xnor U18442 (N_18442,N_14030,N_13320);
nand U18443 (N_18443,N_12996,N_14433);
and U18444 (N_18444,N_14737,N_12752);
or U18445 (N_18445,N_12957,N_15017);
xnor U18446 (N_18446,N_12749,N_13816);
nor U18447 (N_18447,N_13369,N_15591);
nand U18448 (N_18448,N_14453,N_13999);
nand U18449 (N_18449,N_14922,N_15728);
and U18450 (N_18450,N_12181,N_13404);
xnor U18451 (N_18451,N_15716,N_14377);
or U18452 (N_18452,N_12790,N_12183);
xnor U18453 (N_18453,N_14321,N_15075);
or U18454 (N_18454,N_14321,N_14621);
or U18455 (N_18455,N_14128,N_12003);
or U18456 (N_18456,N_14428,N_13545);
nand U18457 (N_18457,N_14261,N_13617);
and U18458 (N_18458,N_14483,N_14461);
nand U18459 (N_18459,N_12266,N_12448);
nand U18460 (N_18460,N_14060,N_13678);
nand U18461 (N_18461,N_13338,N_15552);
and U18462 (N_18462,N_15521,N_15832);
xor U18463 (N_18463,N_15362,N_14398);
or U18464 (N_18464,N_13571,N_12264);
and U18465 (N_18465,N_13323,N_14707);
nor U18466 (N_18466,N_15877,N_14687);
and U18467 (N_18467,N_12460,N_13483);
nand U18468 (N_18468,N_14955,N_13813);
or U18469 (N_18469,N_15745,N_13922);
nor U18470 (N_18470,N_12086,N_14498);
and U18471 (N_18471,N_13022,N_13076);
xor U18472 (N_18472,N_14210,N_13498);
xnor U18473 (N_18473,N_14956,N_14263);
nand U18474 (N_18474,N_13547,N_15627);
or U18475 (N_18475,N_13132,N_14041);
nor U18476 (N_18476,N_13943,N_12533);
and U18477 (N_18477,N_15940,N_13475);
xor U18478 (N_18478,N_12632,N_12485);
and U18479 (N_18479,N_14811,N_13881);
nand U18480 (N_18480,N_15733,N_15978);
nor U18481 (N_18481,N_14285,N_15308);
and U18482 (N_18482,N_12452,N_15731);
and U18483 (N_18483,N_15186,N_15979);
and U18484 (N_18484,N_13771,N_14804);
nand U18485 (N_18485,N_15513,N_15039);
nand U18486 (N_18486,N_13164,N_12312);
and U18487 (N_18487,N_12465,N_13460);
xor U18488 (N_18488,N_15816,N_14884);
nor U18489 (N_18489,N_13720,N_14922);
xor U18490 (N_18490,N_12739,N_15710);
nor U18491 (N_18491,N_15502,N_12616);
nand U18492 (N_18492,N_14529,N_13518);
xnor U18493 (N_18493,N_15633,N_13702);
xnor U18494 (N_18494,N_14177,N_13326);
and U18495 (N_18495,N_13956,N_12703);
nor U18496 (N_18496,N_14555,N_12056);
nand U18497 (N_18497,N_14041,N_15519);
xor U18498 (N_18498,N_14377,N_12151);
nand U18499 (N_18499,N_14838,N_12446);
nand U18500 (N_18500,N_14893,N_15160);
nor U18501 (N_18501,N_15769,N_15370);
or U18502 (N_18502,N_15736,N_15243);
or U18503 (N_18503,N_14684,N_15708);
or U18504 (N_18504,N_13547,N_12057);
nor U18505 (N_18505,N_13934,N_15425);
or U18506 (N_18506,N_14837,N_13518);
or U18507 (N_18507,N_13253,N_13153);
nor U18508 (N_18508,N_15978,N_15111);
or U18509 (N_18509,N_12958,N_13574);
nand U18510 (N_18510,N_12999,N_14227);
or U18511 (N_18511,N_13787,N_12923);
nand U18512 (N_18512,N_14060,N_15779);
nor U18513 (N_18513,N_12823,N_12179);
xor U18514 (N_18514,N_13801,N_12541);
nand U18515 (N_18515,N_15300,N_12562);
nor U18516 (N_18516,N_14777,N_15034);
nor U18517 (N_18517,N_12965,N_13945);
or U18518 (N_18518,N_14610,N_13030);
and U18519 (N_18519,N_15475,N_13093);
and U18520 (N_18520,N_14961,N_14221);
nor U18521 (N_18521,N_13940,N_14305);
xnor U18522 (N_18522,N_14240,N_15423);
nand U18523 (N_18523,N_15480,N_15487);
and U18524 (N_18524,N_12604,N_14310);
nand U18525 (N_18525,N_12042,N_14245);
nand U18526 (N_18526,N_12550,N_14321);
and U18527 (N_18527,N_13087,N_12503);
xor U18528 (N_18528,N_14520,N_12432);
nand U18529 (N_18529,N_13280,N_14801);
nor U18530 (N_18530,N_14536,N_15884);
nand U18531 (N_18531,N_12715,N_14963);
xnor U18532 (N_18532,N_14858,N_13154);
or U18533 (N_18533,N_13855,N_12172);
nor U18534 (N_18534,N_15282,N_13893);
nand U18535 (N_18535,N_14201,N_15187);
xnor U18536 (N_18536,N_14438,N_14730);
or U18537 (N_18537,N_12498,N_13872);
or U18538 (N_18538,N_15049,N_15014);
nand U18539 (N_18539,N_15809,N_14248);
nand U18540 (N_18540,N_12692,N_12897);
and U18541 (N_18541,N_13396,N_15359);
nor U18542 (N_18542,N_13770,N_14464);
and U18543 (N_18543,N_15560,N_13477);
or U18544 (N_18544,N_12346,N_14160);
or U18545 (N_18545,N_12651,N_14563);
xnor U18546 (N_18546,N_13974,N_13895);
nor U18547 (N_18547,N_12907,N_14904);
or U18548 (N_18548,N_14290,N_14260);
nand U18549 (N_18549,N_12158,N_12834);
xor U18550 (N_18550,N_13426,N_13393);
nand U18551 (N_18551,N_15643,N_14271);
nand U18552 (N_18552,N_12396,N_13956);
nor U18553 (N_18553,N_14377,N_15099);
xor U18554 (N_18554,N_12443,N_12613);
xor U18555 (N_18555,N_13220,N_12513);
or U18556 (N_18556,N_12752,N_13076);
nor U18557 (N_18557,N_13745,N_13611);
or U18558 (N_18558,N_14956,N_13529);
xor U18559 (N_18559,N_13141,N_12118);
nand U18560 (N_18560,N_14924,N_14968);
and U18561 (N_18561,N_12157,N_13898);
nand U18562 (N_18562,N_12175,N_14830);
nor U18563 (N_18563,N_12982,N_13688);
nor U18564 (N_18564,N_15341,N_14091);
and U18565 (N_18565,N_13930,N_15227);
nand U18566 (N_18566,N_14340,N_14627);
xor U18567 (N_18567,N_15182,N_14484);
nand U18568 (N_18568,N_12798,N_14409);
nand U18569 (N_18569,N_13198,N_12550);
xnor U18570 (N_18570,N_13730,N_12493);
xor U18571 (N_18571,N_12529,N_14336);
or U18572 (N_18572,N_12127,N_13449);
xor U18573 (N_18573,N_12311,N_14354);
nand U18574 (N_18574,N_14584,N_13287);
nor U18575 (N_18575,N_15419,N_15017);
nor U18576 (N_18576,N_14984,N_12417);
nand U18577 (N_18577,N_12459,N_12791);
xor U18578 (N_18578,N_14365,N_12332);
xor U18579 (N_18579,N_15857,N_14587);
and U18580 (N_18580,N_14846,N_15844);
or U18581 (N_18581,N_15122,N_13584);
or U18582 (N_18582,N_14604,N_14197);
xnor U18583 (N_18583,N_15452,N_12354);
and U18584 (N_18584,N_14966,N_14000);
xor U18585 (N_18585,N_13579,N_13250);
or U18586 (N_18586,N_14366,N_14640);
nand U18587 (N_18587,N_14789,N_13119);
nand U18588 (N_18588,N_15517,N_14862);
xor U18589 (N_18589,N_13639,N_15168);
nand U18590 (N_18590,N_14515,N_15076);
nand U18591 (N_18591,N_15802,N_12358);
nand U18592 (N_18592,N_14559,N_13025);
xnor U18593 (N_18593,N_13034,N_13297);
nand U18594 (N_18594,N_13344,N_15832);
nor U18595 (N_18595,N_14897,N_12791);
and U18596 (N_18596,N_14673,N_13088);
nor U18597 (N_18597,N_15427,N_15870);
or U18598 (N_18598,N_12355,N_15732);
and U18599 (N_18599,N_15130,N_15591);
and U18600 (N_18600,N_15900,N_15443);
and U18601 (N_18601,N_15387,N_13347);
nand U18602 (N_18602,N_15981,N_12119);
or U18603 (N_18603,N_13610,N_13912);
nor U18604 (N_18604,N_13342,N_13422);
nand U18605 (N_18605,N_12719,N_13241);
xor U18606 (N_18606,N_13964,N_15372);
nand U18607 (N_18607,N_13589,N_13492);
and U18608 (N_18608,N_13224,N_12313);
and U18609 (N_18609,N_12730,N_14872);
nand U18610 (N_18610,N_12282,N_12405);
and U18611 (N_18611,N_12779,N_14474);
nor U18612 (N_18612,N_14148,N_13135);
and U18613 (N_18613,N_12753,N_14265);
nor U18614 (N_18614,N_15251,N_13843);
or U18615 (N_18615,N_13788,N_12429);
and U18616 (N_18616,N_14204,N_12720);
nor U18617 (N_18617,N_15621,N_15716);
and U18618 (N_18618,N_12982,N_13864);
xnor U18619 (N_18619,N_15680,N_12627);
xor U18620 (N_18620,N_15073,N_15873);
nor U18621 (N_18621,N_14758,N_12461);
or U18622 (N_18622,N_12076,N_14919);
or U18623 (N_18623,N_14190,N_13951);
and U18624 (N_18624,N_13724,N_15660);
or U18625 (N_18625,N_13682,N_13574);
nor U18626 (N_18626,N_13127,N_12090);
and U18627 (N_18627,N_15905,N_12465);
or U18628 (N_18628,N_14140,N_15798);
nor U18629 (N_18629,N_14291,N_12959);
xor U18630 (N_18630,N_14139,N_13901);
or U18631 (N_18631,N_14264,N_13291);
xnor U18632 (N_18632,N_14392,N_13602);
or U18633 (N_18633,N_14916,N_14726);
xor U18634 (N_18634,N_14914,N_12394);
nand U18635 (N_18635,N_15332,N_13303);
xor U18636 (N_18636,N_14853,N_15169);
nor U18637 (N_18637,N_13832,N_14000);
nor U18638 (N_18638,N_15999,N_12624);
and U18639 (N_18639,N_14495,N_13674);
nor U18640 (N_18640,N_15846,N_15766);
or U18641 (N_18641,N_14906,N_12568);
xor U18642 (N_18642,N_13295,N_14962);
xnor U18643 (N_18643,N_12453,N_14508);
nand U18644 (N_18644,N_13966,N_14453);
nor U18645 (N_18645,N_14892,N_14543);
and U18646 (N_18646,N_12618,N_15437);
nand U18647 (N_18647,N_14924,N_13160);
and U18648 (N_18648,N_12186,N_14203);
xor U18649 (N_18649,N_14945,N_12283);
or U18650 (N_18650,N_13472,N_13427);
xor U18651 (N_18651,N_13444,N_15181);
and U18652 (N_18652,N_15638,N_14981);
or U18653 (N_18653,N_15366,N_12956);
xor U18654 (N_18654,N_12532,N_14956);
nand U18655 (N_18655,N_14892,N_13901);
nor U18656 (N_18656,N_15359,N_13513);
or U18657 (N_18657,N_13895,N_14813);
nor U18658 (N_18658,N_12518,N_15639);
nand U18659 (N_18659,N_15981,N_12957);
nand U18660 (N_18660,N_15151,N_13553);
nor U18661 (N_18661,N_15426,N_14531);
nand U18662 (N_18662,N_12150,N_14400);
xnor U18663 (N_18663,N_13470,N_13793);
nor U18664 (N_18664,N_14032,N_12148);
nor U18665 (N_18665,N_13973,N_15721);
nor U18666 (N_18666,N_13217,N_12808);
or U18667 (N_18667,N_13552,N_13049);
and U18668 (N_18668,N_15915,N_14000);
or U18669 (N_18669,N_14659,N_12848);
and U18670 (N_18670,N_13497,N_13567);
and U18671 (N_18671,N_12954,N_12238);
and U18672 (N_18672,N_14721,N_13519);
and U18673 (N_18673,N_12214,N_14072);
or U18674 (N_18674,N_13442,N_14666);
nand U18675 (N_18675,N_14938,N_14787);
or U18676 (N_18676,N_14300,N_14956);
nor U18677 (N_18677,N_15123,N_12758);
nor U18678 (N_18678,N_13347,N_15791);
xor U18679 (N_18679,N_12769,N_13832);
and U18680 (N_18680,N_14111,N_12165);
or U18681 (N_18681,N_12362,N_14227);
nand U18682 (N_18682,N_15358,N_14683);
xnor U18683 (N_18683,N_13070,N_13562);
nor U18684 (N_18684,N_13284,N_14862);
and U18685 (N_18685,N_13950,N_14968);
nor U18686 (N_18686,N_12516,N_14612);
xor U18687 (N_18687,N_13642,N_13197);
or U18688 (N_18688,N_14487,N_15787);
nand U18689 (N_18689,N_12855,N_14244);
or U18690 (N_18690,N_12641,N_13065);
xor U18691 (N_18691,N_15848,N_14872);
nand U18692 (N_18692,N_13910,N_13964);
nand U18693 (N_18693,N_12714,N_14234);
and U18694 (N_18694,N_13568,N_14283);
or U18695 (N_18695,N_14414,N_15782);
nor U18696 (N_18696,N_15091,N_13304);
or U18697 (N_18697,N_14875,N_15581);
nand U18698 (N_18698,N_13580,N_13047);
and U18699 (N_18699,N_12373,N_12516);
nand U18700 (N_18700,N_15790,N_12581);
nand U18701 (N_18701,N_14511,N_12995);
nor U18702 (N_18702,N_14298,N_14550);
or U18703 (N_18703,N_13850,N_14512);
nand U18704 (N_18704,N_15474,N_14742);
or U18705 (N_18705,N_12784,N_13231);
xnor U18706 (N_18706,N_14787,N_13674);
xor U18707 (N_18707,N_13042,N_13258);
nand U18708 (N_18708,N_15167,N_13078);
or U18709 (N_18709,N_12766,N_13143);
nor U18710 (N_18710,N_14162,N_14784);
nor U18711 (N_18711,N_12875,N_12429);
or U18712 (N_18712,N_13186,N_14550);
or U18713 (N_18713,N_14302,N_14532);
xor U18714 (N_18714,N_14230,N_15139);
nand U18715 (N_18715,N_14524,N_14455);
and U18716 (N_18716,N_14432,N_12418);
nor U18717 (N_18717,N_12444,N_14674);
xnor U18718 (N_18718,N_14106,N_12196);
and U18719 (N_18719,N_14227,N_13091);
nor U18720 (N_18720,N_15674,N_12237);
nor U18721 (N_18721,N_14028,N_12816);
and U18722 (N_18722,N_12765,N_13970);
or U18723 (N_18723,N_15379,N_15664);
xnor U18724 (N_18724,N_14965,N_15206);
nor U18725 (N_18725,N_12976,N_14811);
and U18726 (N_18726,N_14877,N_12113);
nand U18727 (N_18727,N_15211,N_12514);
nor U18728 (N_18728,N_13842,N_13527);
and U18729 (N_18729,N_12621,N_14525);
nor U18730 (N_18730,N_14059,N_12793);
nand U18731 (N_18731,N_13143,N_14139);
nor U18732 (N_18732,N_14567,N_13079);
nor U18733 (N_18733,N_13643,N_14806);
nand U18734 (N_18734,N_13956,N_12264);
or U18735 (N_18735,N_13422,N_13938);
nand U18736 (N_18736,N_15136,N_13921);
and U18737 (N_18737,N_12546,N_13029);
nor U18738 (N_18738,N_14583,N_14957);
nor U18739 (N_18739,N_15464,N_14787);
and U18740 (N_18740,N_13980,N_15616);
and U18741 (N_18741,N_13697,N_13935);
or U18742 (N_18742,N_14521,N_15588);
and U18743 (N_18743,N_13197,N_15491);
xor U18744 (N_18744,N_13037,N_14004);
xor U18745 (N_18745,N_13800,N_13628);
and U18746 (N_18746,N_14979,N_15304);
and U18747 (N_18747,N_15104,N_13363);
xor U18748 (N_18748,N_12130,N_12413);
nand U18749 (N_18749,N_14558,N_15333);
nand U18750 (N_18750,N_12005,N_14587);
and U18751 (N_18751,N_14503,N_13233);
nand U18752 (N_18752,N_12899,N_13376);
or U18753 (N_18753,N_13534,N_13528);
xor U18754 (N_18754,N_12576,N_12677);
nand U18755 (N_18755,N_14263,N_13022);
nor U18756 (N_18756,N_12322,N_12863);
or U18757 (N_18757,N_15919,N_15247);
nand U18758 (N_18758,N_13606,N_13252);
and U18759 (N_18759,N_12007,N_14535);
and U18760 (N_18760,N_14358,N_14138);
nor U18761 (N_18761,N_14718,N_14258);
xnor U18762 (N_18762,N_12286,N_12123);
xnor U18763 (N_18763,N_15495,N_12418);
xnor U18764 (N_18764,N_14206,N_13359);
or U18765 (N_18765,N_12933,N_14083);
nor U18766 (N_18766,N_13806,N_13729);
nand U18767 (N_18767,N_12818,N_13955);
or U18768 (N_18768,N_14469,N_15995);
or U18769 (N_18769,N_13653,N_15008);
and U18770 (N_18770,N_12653,N_14108);
nand U18771 (N_18771,N_15234,N_14132);
nor U18772 (N_18772,N_12291,N_14217);
or U18773 (N_18773,N_15200,N_15906);
or U18774 (N_18774,N_15172,N_15094);
nand U18775 (N_18775,N_14984,N_13882);
or U18776 (N_18776,N_12699,N_12474);
and U18777 (N_18777,N_14818,N_15783);
or U18778 (N_18778,N_12852,N_12217);
nand U18779 (N_18779,N_14776,N_15327);
or U18780 (N_18780,N_13636,N_12784);
or U18781 (N_18781,N_12753,N_12607);
nor U18782 (N_18782,N_14791,N_15539);
nand U18783 (N_18783,N_12026,N_14813);
nor U18784 (N_18784,N_14954,N_12463);
nand U18785 (N_18785,N_12357,N_14015);
or U18786 (N_18786,N_12464,N_15956);
and U18787 (N_18787,N_14535,N_12913);
or U18788 (N_18788,N_12082,N_12129);
xor U18789 (N_18789,N_14244,N_13723);
xor U18790 (N_18790,N_12088,N_13906);
nand U18791 (N_18791,N_12872,N_12756);
nand U18792 (N_18792,N_15229,N_13825);
nor U18793 (N_18793,N_14257,N_14372);
and U18794 (N_18794,N_12340,N_14416);
nor U18795 (N_18795,N_13271,N_12476);
or U18796 (N_18796,N_13326,N_12349);
and U18797 (N_18797,N_14133,N_13965);
or U18798 (N_18798,N_13024,N_14076);
or U18799 (N_18799,N_12399,N_13631);
nor U18800 (N_18800,N_14283,N_15497);
nor U18801 (N_18801,N_12956,N_12661);
and U18802 (N_18802,N_15953,N_15773);
or U18803 (N_18803,N_15261,N_14653);
xnor U18804 (N_18804,N_14665,N_14986);
or U18805 (N_18805,N_12894,N_15660);
nor U18806 (N_18806,N_14055,N_12771);
and U18807 (N_18807,N_13825,N_13916);
nand U18808 (N_18808,N_12974,N_12137);
xor U18809 (N_18809,N_13592,N_14449);
nand U18810 (N_18810,N_13823,N_12409);
nor U18811 (N_18811,N_14368,N_14978);
xnor U18812 (N_18812,N_13663,N_12046);
or U18813 (N_18813,N_14228,N_13092);
or U18814 (N_18814,N_12354,N_14785);
nor U18815 (N_18815,N_12325,N_13628);
and U18816 (N_18816,N_12930,N_13912);
or U18817 (N_18817,N_14260,N_13382);
and U18818 (N_18818,N_13789,N_14012);
or U18819 (N_18819,N_15948,N_15583);
xnor U18820 (N_18820,N_14191,N_15132);
and U18821 (N_18821,N_13587,N_15550);
or U18822 (N_18822,N_15355,N_15264);
and U18823 (N_18823,N_14281,N_14191);
or U18824 (N_18824,N_14491,N_14823);
or U18825 (N_18825,N_15255,N_15663);
nor U18826 (N_18826,N_15343,N_14066);
nor U18827 (N_18827,N_14399,N_12837);
nor U18828 (N_18828,N_14129,N_15623);
xor U18829 (N_18829,N_14786,N_13503);
nand U18830 (N_18830,N_12604,N_13843);
xor U18831 (N_18831,N_13210,N_14812);
nor U18832 (N_18832,N_13313,N_12020);
nand U18833 (N_18833,N_15501,N_12375);
nor U18834 (N_18834,N_13558,N_12346);
nand U18835 (N_18835,N_12018,N_13476);
or U18836 (N_18836,N_15524,N_14731);
or U18837 (N_18837,N_13734,N_15387);
or U18838 (N_18838,N_15043,N_15809);
nor U18839 (N_18839,N_12814,N_14972);
or U18840 (N_18840,N_13366,N_12711);
or U18841 (N_18841,N_15833,N_14007);
xor U18842 (N_18842,N_12933,N_12260);
nor U18843 (N_18843,N_14451,N_13845);
or U18844 (N_18844,N_14041,N_14380);
or U18845 (N_18845,N_14203,N_15269);
and U18846 (N_18846,N_12302,N_15703);
nor U18847 (N_18847,N_12743,N_14952);
nand U18848 (N_18848,N_12951,N_13734);
and U18849 (N_18849,N_12739,N_13035);
and U18850 (N_18850,N_15965,N_14654);
nor U18851 (N_18851,N_13851,N_12680);
xor U18852 (N_18852,N_14884,N_14309);
or U18853 (N_18853,N_14663,N_15479);
and U18854 (N_18854,N_12975,N_15516);
nor U18855 (N_18855,N_12196,N_15135);
nor U18856 (N_18856,N_12191,N_15084);
xnor U18857 (N_18857,N_15860,N_12827);
nor U18858 (N_18858,N_15924,N_12681);
nand U18859 (N_18859,N_14754,N_15217);
nor U18860 (N_18860,N_13368,N_14875);
and U18861 (N_18861,N_14138,N_13737);
nor U18862 (N_18862,N_12966,N_13293);
xor U18863 (N_18863,N_15213,N_13614);
or U18864 (N_18864,N_14119,N_14571);
nand U18865 (N_18865,N_15489,N_14899);
or U18866 (N_18866,N_14679,N_15143);
or U18867 (N_18867,N_12639,N_13395);
or U18868 (N_18868,N_15458,N_12928);
and U18869 (N_18869,N_15919,N_14589);
and U18870 (N_18870,N_13520,N_12380);
and U18871 (N_18871,N_13799,N_12340);
or U18872 (N_18872,N_15639,N_15684);
nor U18873 (N_18873,N_14293,N_14842);
nor U18874 (N_18874,N_15817,N_15325);
nand U18875 (N_18875,N_12891,N_14317);
xnor U18876 (N_18876,N_14664,N_13443);
xor U18877 (N_18877,N_15912,N_15512);
xnor U18878 (N_18878,N_12996,N_15500);
and U18879 (N_18879,N_14256,N_13195);
nand U18880 (N_18880,N_14833,N_13572);
or U18881 (N_18881,N_13413,N_15630);
and U18882 (N_18882,N_13655,N_12560);
and U18883 (N_18883,N_13165,N_12425);
and U18884 (N_18884,N_14050,N_15092);
nor U18885 (N_18885,N_15426,N_13018);
nor U18886 (N_18886,N_14918,N_15655);
and U18887 (N_18887,N_15050,N_15804);
and U18888 (N_18888,N_14190,N_12153);
nor U18889 (N_18889,N_12670,N_15818);
nand U18890 (N_18890,N_13197,N_12845);
and U18891 (N_18891,N_14730,N_15147);
or U18892 (N_18892,N_14184,N_13879);
and U18893 (N_18893,N_15717,N_13090);
and U18894 (N_18894,N_15367,N_14366);
xor U18895 (N_18895,N_12320,N_15602);
xnor U18896 (N_18896,N_13232,N_15427);
nor U18897 (N_18897,N_14546,N_14699);
nand U18898 (N_18898,N_14285,N_13070);
xor U18899 (N_18899,N_13945,N_13807);
xnor U18900 (N_18900,N_14233,N_12800);
nor U18901 (N_18901,N_13821,N_14358);
xnor U18902 (N_18902,N_12040,N_13361);
or U18903 (N_18903,N_12541,N_12400);
nand U18904 (N_18904,N_12601,N_12684);
or U18905 (N_18905,N_15767,N_13774);
and U18906 (N_18906,N_14940,N_14647);
nor U18907 (N_18907,N_13937,N_14916);
or U18908 (N_18908,N_13337,N_12232);
xor U18909 (N_18909,N_12955,N_13196);
and U18910 (N_18910,N_12501,N_15312);
xnor U18911 (N_18911,N_12630,N_15502);
and U18912 (N_18912,N_13985,N_15769);
and U18913 (N_18913,N_14364,N_15684);
nand U18914 (N_18914,N_13122,N_13762);
and U18915 (N_18915,N_13156,N_13445);
or U18916 (N_18916,N_13459,N_15262);
or U18917 (N_18917,N_12344,N_14862);
nor U18918 (N_18918,N_14814,N_14038);
or U18919 (N_18919,N_12585,N_13793);
or U18920 (N_18920,N_12808,N_14156);
xor U18921 (N_18921,N_12159,N_14883);
and U18922 (N_18922,N_14571,N_14731);
nand U18923 (N_18923,N_14731,N_15298);
and U18924 (N_18924,N_12985,N_13797);
xor U18925 (N_18925,N_15284,N_14250);
nor U18926 (N_18926,N_12514,N_12386);
xor U18927 (N_18927,N_12311,N_15866);
xnor U18928 (N_18928,N_14771,N_15456);
xor U18929 (N_18929,N_15195,N_15371);
nor U18930 (N_18930,N_13651,N_12001);
nand U18931 (N_18931,N_12994,N_12752);
nand U18932 (N_18932,N_13861,N_12880);
and U18933 (N_18933,N_12773,N_12809);
nor U18934 (N_18934,N_15709,N_14125);
nand U18935 (N_18935,N_14733,N_12627);
nand U18936 (N_18936,N_14223,N_15549);
nor U18937 (N_18937,N_15404,N_13944);
nand U18938 (N_18938,N_12472,N_15468);
nor U18939 (N_18939,N_13838,N_15430);
xnor U18940 (N_18940,N_12667,N_15684);
and U18941 (N_18941,N_12927,N_15964);
or U18942 (N_18942,N_15064,N_15212);
xnor U18943 (N_18943,N_13745,N_15849);
and U18944 (N_18944,N_14968,N_12746);
nand U18945 (N_18945,N_12767,N_14085);
xnor U18946 (N_18946,N_13412,N_13909);
and U18947 (N_18947,N_14662,N_15290);
xor U18948 (N_18948,N_14803,N_12376);
nand U18949 (N_18949,N_13927,N_15585);
or U18950 (N_18950,N_15657,N_12040);
and U18951 (N_18951,N_12317,N_12682);
and U18952 (N_18952,N_13323,N_13670);
nor U18953 (N_18953,N_12232,N_14711);
nand U18954 (N_18954,N_14861,N_14146);
nor U18955 (N_18955,N_14766,N_14320);
and U18956 (N_18956,N_12432,N_15393);
and U18957 (N_18957,N_12499,N_15158);
xnor U18958 (N_18958,N_12078,N_13741);
and U18959 (N_18959,N_15516,N_12826);
xnor U18960 (N_18960,N_13028,N_12518);
nand U18961 (N_18961,N_13506,N_12918);
xnor U18962 (N_18962,N_15748,N_15203);
nor U18963 (N_18963,N_14518,N_15062);
or U18964 (N_18964,N_12596,N_12845);
nand U18965 (N_18965,N_13395,N_15503);
nand U18966 (N_18966,N_12883,N_15067);
or U18967 (N_18967,N_13114,N_12655);
and U18968 (N_18968,N_14345,N_14698);
nor U18969 (N_18969,N_12055,N_13658);
nor U18970 (N_18970,N_14331,N_13687);
nor U18971 (N_18971,N_12303,N_14930);
or U18972 (N_18972,N_12124,N_12828);
nor U18973 (N_18973,N_15426,N_15058);
xor U18974 (N_18974,N_13414,N_14135);
nor U18975 (N_18975,N_15268,N_12564);
and U18976 (N_18976,N_12910,N_12997);
or U18977 (N_18977,N_13132,N_12387);
or U18978 (N_18978,N_13037,N_13904);
xnor U18979 (N_18979,N_14890,N_15033);
or U18980 (N_18980,N_14553,N_13005);
xor U18981 (N_18981,N_13476,N_13671);
and U18982 (N_18982,N_14595,N_13658);
and U18983 (N_18983,N_12673,N_14573);
or U18984 (N_18984,N_14296,N_14322);
or U18985 (N_18985,N_13649,N_13085);
and U18986 (N_18986,N_12285,N_14430);
and U18987 (N_18987,N_15280,N_12868);
or U18988 (N_18988,N_12016,N_14354);
nor U18989 (N_18989,N_13974,N_12241);
nand U18990 (N_18990,N_12749,N_13230);
or U18991 (N_18991,N_12480,N_13243);
and U18992 (N_18992,N_15351,N_12524);
nand U18993 (N_18993,N_15405,N_13947);
xor U18994 (N_18994,N_13133,N_15446);
nand U18995 (N_18995,N_13106,N_12157);
or U18996 (N_18996,N_15210,N_14188);
nand U18997 (N_18997,N_14856,N_14196);
and U18998 (N_18998,N_13979,N_14672);
nor U18999 (N_18999,N_14377,N_14106);
and U19000 (N_19000,N_12116,N_15186);
and U19001 (N_19001,N_14779,N_15080);
or U19002 (N_19002,N_13566,N_15917);
or U19003 (N_19003,N_14244,N_13951);
or U19004 (N_19004,N_15801,N_12448);
and U19005 (N_19005,N_12286,N_12940);
nor U19006 (N_19006,N_13762,N_14227);
and U19007 (N_19007,N_15111,N_15559);
nor U19008 (N_19008,N_13740,N_14583);
nand U19009 (N_19009,N_15897,N_13027);
xor U19010 (N_19010,N_14161,N_15656);
or U19011 (N_19011,N_13384,N_12622);
and U19012 (N_19012,N_15329,N_15925);
xnor U19013 (N_19013,N_14888,N_12986);
or U19014 (N_19014,N_13428,N_12530);
nand U19015 (N_19015,N_12328,N_15322);
xor U19016 (N_19016,N_13859,N_12442);
xor U19017 (N_19017,N_12925,N_13524);
nand U19018 (N_19018,N_14602,N_14695);
nand U19019 (N_19019,N_13215,N_12114);
and U19020 (N_19020,N_15715,N_13839);
nor U19021 (N_19021,N_15699,N_15885);
nor U19022 (N_19022,N_15518,N_13423);
nand U19023 (N_19023,N_15880,N_12118);
xnor U19024 (N_19024,N_14254,N_14594);
nand U19025 (N_19025,N_14478,N_14485);
nand U19026 (N_19026,N_14069,N_15002);
nand U19027 (N_19027,N_13065,N_15357);
or U19028 (N_19028,N_12186,N_12635);
nor U19029 (N_19029,N_15285,N_14071);
xnor U19030 (N_19030,N_14203,N_15599);
and U19031 (N_19031,N_14635,N_14007);
and U19032 (N_19032,N_14845,N_13969);
xnor U19033 (N_19033,N_14688,N_12297);
xor U19034 (N_19034,N_14426,N_12418);
nor U19035 (N_19035,N_14629,N_12070);
nor U19036 (N_19036,N_15873,N_13382);
nor U19037 (N_19037,N_13419,N_13347);
xor U19038 (N_19038,N_12966,N_13937);
or U19039 (N_19039,N_15180,N_15686);
nand U19040 (N_19040,N_15643,N_14695);
nand U19041 (N_19041,N_12470,N_12180);
nand U19042 (N_19042,N_14435,N_12366);
xnor U19043 (N_19043,N_13131,N_13104);
nor U19044 (N_19044,N_12064,N_15797);
or U19045 (N_19045,N_14635,N_15631);
xor U19046 (N_19046,N_14217,N_14813);
and U19047 (N_19047,N_13791,N_14052);
nand U19048 (N_19048,N_14800,N_13521);
xnor U19049 (N_19049,N_13135,N_13878);
xnor U19050 (N_19050,N_15553,N_12171);
nor U19051 (N_19051,N_12895,N_12662);
nor U19052 (N_19052,N_15534,N_13786);
or U19053 (N_19053,N_13615,N_15924);
xnor U19054 (N_19054,N_14197,N_13954);
nor U19055 (N_19055,N_12445,N_14500);
nand U19056 (N_19056,N_14694,N_13997);
xnor U19057 (N_19057,N_12851,N_15341);
xor U19058 (N_19058,N_12851,N_12319);
nand U19059 (N_19059,N_15784,N_12046);
nor U19060 (N_19060,N_14063,N_14045);
or U19061 (N_19061,N_13547,N_13132);
nand U19062 (N_19062,N_15870,N_15902);
and U19063 (N_19063,N_14684,N_15601);
nor U19064 (N_19064,N_12550,N_14334);
nand U19065 (N_19065,N_15921,N_15702);
xor U19066 (N_19066,N_14814,N_12485);
and U19067 (N_19067,N_13248,N_13082);
and U19068 (N_19068,N_13287,N_12857);
nor U19069 (N_19069,N_15016,N_12314);
nand U19070 (N_19070,N_15407,N_14596);
nor U19071 (N_19071,N_12222,N_12632);
and U19072 (N_19072,N_12563,N_13716);
nor U19073 (N_19073,N_12964,N_13030);
and U19074 (N_19074,N_14618,N_12218);
nand U19075 (N_19075,N_12666,N_14223);
or U19076 (N_19076,N_15647,N_14644);
and U19077 (N_19077,N_12255,N_15277);
nor U19078 (N_19078,N_15223,N_13702);
nor U19079 (N_19079,N_15167,N_12839);
and U19080 (N_19080,N_14183,N_14299);
nor U19081 (N_19081,N_15672,N_15863);
nand U19082 (N_19082,N_15209,N_13962);
nor U19083 (N_19083,N_15245,N_15392);
xor U19084 (N_19084,N_13000,N_15395);
xnor U19085 (N_19085,N_14608,N_15813);
xnor U19086 (N_19086,N_15171,N_14941);
nand U19087 (N_19087,N_15430,N_14686);
or U19088 (N_19088,N_15904,N_14373);
or U19089 (N_19089,N_14519,N_14963);
xor U19090 (N_19090,N_14566,N_15424);
and U19091 (N_19091,N_14149,N_13998);
nand U19092 (N_19092,N_12919,N_14829);
and U19093 (N_19093,N_12021,N_15208);
nand U19094 (N_19094,N_14163,N_14243);
nand U19095 (N_19095,N_15902,N_13434);
nor U19096 (N_19096,N_15573,N_13194);
and U19097 (N_19097,N_14131,N_15697);
nand U19098 (N_19098,N_15443,N_14076);
nand U19099 (N_19099,N_15279,N_15900);
nor U19100 (N_19100,N_13565,N_12920);
nor U19101 (N_19101,N_13494,N_12882);
nand U19102 (N_19102,N_12804,N_12271);
xnor U19103 (N_19103,N_14399,N_14659);
xnor U19104 (N_19104,N_15014,N_12426);
nand U19105 (N_19105,N_14394,N_13927);
xnor U19106 (N_19106,N_12260,N_12672);
xnor U19107 (N_19107,N_15879,N_13453);
xnor U19108 (N_19108,N_14669,N_15517);
or U19109 (N_19109,N_14180,N_15813);
and U19110 (N_19110,N_14046,N_13363);
and U19111 (N_19111,N_15328,N_15860);
nor U19112 (N_19112,N_13504,N_13070);
nand U19113 (N_19113,N_12557,N_12484);
xor U19114 (N_19114,N_14183,N_13651);
nor U19115 (N_19115,N_14800,N_14985);
xor U19116 (N_19116,N_14384,N_14841);
nand U19117 (N_19117,N_14535,N_13520);
nand U19118 (N_19118,N_14152,N_14712);
nand U19119 (N_19119,N_14507,N_15606);
nor U19120 (N_19120,N_12401,N_12020);
and U19121 (N_19121,N_12240,N_14002);
nor U19122 (N_19122,N_12856,N_14663);
and U19123 (N_19123,N_13900,N_14178);
or U19124 (N_19124,N_13739,N_14534);
or U19125 (N_19125,N_13019,N_14339);
and U19126 (N_19126,N_12538,N_12839);
or U19127 (N_19127,N_14052,N_12725);
xnor U19128 (N_19128,N_15062,N_14071);
and U19129 (N_19129,N_12583,N_15813);
nand U19130 (N_19130,N_12009,N_12395);
or U19131 (N_19131,N_12563,N_14073);
nor U19132 (N_19132,N_12110,N_15873);
xor U19133 (N_19133,N_15786,N_13402);
nor U19134 (N_19134,N_14073,N_13107);
and U19135 (N_19135,N_13221,N_15861);
or U19136 (N_19136,N_15030,N_15098);
and U19137 (N_19137,N_15301,N_12781);
or U19138 (N_19138,N_13025,N_15676);
or U19139 (N_19139,N_15001,N_15432);
nor U19140 (N_19140,N_14089,N_14763);
xor U19141 (N_19141,N_14334,N_13580);
nor U19142 (N_19142,N_13403,N_14345);
and U19143 (N_19143,N_14348,N_12318);
or U19144 (N_19144,N_14902,N_12855);
or U19145 (N_19145,N_13299,N_12510);
xnor U19146 (N_19146,N_14260,N_15574);
xor U19147 (N_19147,N_12923,N_14942);
nand U19148 (N_19148,N_13391,N_13380);
xnor U19149 (N_19149,N_12348,N_15840);
or U19150 (N_19150,N_15342,N_15792);
nor U19151 (N_19151,N_14995,N_12100);
nand U19152 (N_19152,N_12285,N_12700);
nor U19153 (N_19153,N_12076,N_15902);
and U19154 (N_19154,N_13953,N_15892);
xnor U19155 (N_19155,N_14592,N_14238);
nor U19156 (N_19156,N_15566,N_12636);
nand U19157 (N_19157,N_12211,N_14761);
or U19158 (N_19158,N_12721,N_13175);
nor U19159 (N_19159,N_14037,N_14923);
nor U19160 (N_19160,N_14045,N_13739);
xor U19161 (N_19161,N_12465,N_13095);
xor U19162 (N_19162,N_14986,N_14510);
nor U19163 (N_19163,N_15271,N_13299);
xor U19164 (N_19164,N_14820,N_13917);
xor U19165 (N_19165,N_15360,N_13016);
or U19166 (N_19166,N_12716,N_12883);
or U19167 (N_19167,N_15853,N_14657);
nor U19168 (N_19168,N_14028,N_13752);
xnor U19169 (N_19169,N_12825,N_13089);
nor U19170 (N_19170,N_15381,N_14109);
and U19171 (N_19171,N_13090,N_14337);
nand U19172 (N_19172,N_14416,N_12768);
or U19173 (N_19173,N_13099,N_13862);
and U19174 (N_19174,N_15021,N_14207);
or U19175 (N_19175,N_13652,N_12970);
nor U19176 (N_19176,N_13684,N_15609);
xnor U19177 (N_19177,N_14740,N_12462);
xor U19178 (N_19178,N_15090,N_15168);
and U19179 (N_19179,N_14317,N_15143);
xor U19180 (N_19180,N_12906,N_13938);
nand U19181 (N_19181,N_13552,N_15203);
xnor U19182 (N_19182,N_15784,N_15364);
nor U19183 (N_19183,N_14088,N_15440);
and U19184 (N_19184,N_13436,N_14425);
or U19185 (N_19185,N_14890,N_14445);
nor U19186 (N_19186,N_14512,N_14943);
and U19187 (N_19187,N_13893,N_14657);
and U19188 (N_19188,N_12324,N_12939);
nor U19189 (N_19189,N_12419,N_14606);
nor U19190 (N_19190,N_14100,N_12904);
and U19191 (N_19191,N_15853,N_15855);
nand U19192 (N_19192,N_12717,N_13182);
nand U19193 (N_19193,N_14376,N_15564);
xor U19194 (N_19194,N_13765,N_12831);
nor U19195 (N_19195,N_13737,N_13480);
and U19196 (N_19196,N_15870,N_14782);
or U19197 (N_19197,N_13062,N_13306);
nor U19198 (N_19198,N_12031,N_15884);
and U19199 (N_19199,N_12550,N_15873);
and U19200 (N_19200,N_14911,N_13544);
and U19201 (N_19201,N_14784,N_14602);
or U19202 (N_19202,N_14961,N_13373);
xor U19203 (N_19203,N_14022,N_13318);
xor U19204 (N_19204,N_15102,N_13400);
or U19205 (N_19205,N_14990,N_15070);
and U19206 (N_19206,N_15153,N_14482);
or U19207 (N_19207,N_15441,N_14675);
xor U19208 (N_19208,N_12308,N_12586);
xnor U19209 (N_19209,N_15596,N_15146);
or U19210 (N_19210,N_14094,N_14455);
nand U19211 (N_19211,N_15250,N_15290);
nor U19212 (N_19212,N_13258,N_15974);
nand U19213 (N_19213,N_12285,N_13042);
or U19214 (N_19214,N_14904,N_13191);
or U19215 (N_19215,N_14631,N_14403);
nor U19216 (N_19216,N_12722,N_15363);
or U19217 (N_19217,N_14664,N_14084);
nor U19218 (N_19218,N_15493,N_12974);
xnor U19219 (N_19219,N_15042,N_14029);
or U19220 (N_19220,N_13479,N_15387);
nor U19221 (N_19221,N_13482,N_13809);
nor U19222 (N_19222,N_12567,N_13299);
and U19223 (N_19223,N_13856,N_14768);
or U19224 (N_19224,N_14870,N_12151);
or U19225 (N_19225,N_12764,N_14088);
xor U19226 (N_19226,N_13824,N_12574);
nor U19227 (N_19227,N_12231,N_13015);
or U19228 (N_19228,N_15066,N_12871);
xor U19229 (N_19229,N_14029,N_14580);
xor U19230 (N_19230,N_15247,N_14928);
nor U19231 (N_19231,N_14421,N_15382);
xnor U19232 (N_19232,N_13289,N_15311);
xnor U19233 (N_19233,N_15931,N_13179);
and U19234 (N_19234,N_13694,N_13560);
nand U19235 (N_19235,N_15148,N_14545);
xor U19236 (N_19236,N_14884,N_15527);
nand U19237 (N_19237,N_12744,N_13959);
nor U19238 (N_19238,N_14924,N_12841);
nand U19239 (N_19239,N_14995,N_12751);
and U19240 (N_19240,N_14769,N_12834);
xor U19241 (N_19241,N_12953,N_12251);
nor U19242 (N_19242,N_12714,N_13224);
or U19243 (N_19243,N_13453,N_15997);
xnor U19244 (N_19244,N_13230,N_15119);
or U19245 (N_19245,N_13629,N_12659);
or U19246 (N_19246,N_13766,N_12092);
xor U19247 (N_19247,N_15594,N_13486);
xnor U19248 (N_19248,N_15212,N_12173);
and U19249 (N_19249,N_15803,N_12054);
xor U19250 (N_19250,N_12084,N_14519);
xnor U19251 (N_19251,N_13951,N_14722);
or U19252 (N_19252,N_12439,N_13937);
or U19253 (N_19253,N_15661,N_12660);
xor U19254 (N_19254,N_13017,N_13102);
xor U19255 (N_19255,N_12883,N_14023);
nand U19256 (N_19256,N_12236,N_15693);
nor U19257 (N_19257,N_12496,N_15021);
nor U19258 (N_19258,N_14731,N_13266);
xnor U19259 (N_19259,N_15124,N_12815);
xor U19260 (N_19260,N_15028,N_12470);
xor U19261 (N_19261,N_15930,N_15073);
xor U19262 (N_19262,N_14246,N_13796);
nor U19263 (N_19263,N_13099,N_15758);
nand U19264 (N_19264,N_14457,N_14930);
and U19265 (N_19265,N_12481,N_13541);
and U19266 (N_19266,N_13677,N_14566);
nand U19267 (N_19267,N_14324,N_13563);
nor U19268 (N_19268,N_15727,N_12608);
xor U19269 (N_19269,N_15790,N_13803);
or U19270 (N_19270,N_13944,N_13751);
nor U19271 (N_19271,N_13912,N_15573);
or U19272 (N_19272,N_15836,N_15751);
or U19273 (N_19273,N_13418,N_14923);
xor U19274 (N_19274,N_14692,N_12046);
or U19275 (N_19275,N_12587,N_15538);
xor U19276 (N_19276,N_12213,N_13558);
xor U19277 (N_19277,N_12704,N_15377);
nor U19278 (N_19278,N_13597,N_15960);
or U19279 (N_19279,N_15697,N_15385);
xor U19280 (N_19280,N_12913,N_15233);
or U19281 (N_19281,N_14503,N_15823);
nand U19282 (N_19282,N_14031,N_12933);
nand U19283 (N_19283,N_12165,N_14928);
xnor U19284 (N_19284,N_15315,N_12680);
nor U19285 (N_19285,N_14969,N_13427);
or U19286 (N_19286,N_12839,N_14707);
nand U19287 (N_19287,N_14325,N_15103);
xor U19288 (N_19288,N_14236,N_15766);
nand U19289 (N_19289,N_13008,N_12423);
nor U19290 (N_19290,N_13504,N_13847);
nor U19291 (N_19291,N_13106,N_13149);
nor U19292 (N_19292,N_15894,N_12425);
nand U19293 (N_19293,N_13265,N_14181);
or U19294 (N_19294,N_13218,N_15073);
and U19295 (N_19295,N_15063,N_14116);
xor U19296 (N_19296,N_13637,N_15549);
xnor U19297 (N_19297,N_13962,N_14525);
and U19298 (N_19298,N_13937,N_15285);
or U19299 (N_19299,N_14526,N_14646);
nand U19300 (N_19300,N_14983,N_12318);
nor U19301 (N_19301,N_15306,N_14307);
and U19302 (N_19302,N_14492,N_15165);
or U19303 (N_19303,N_13609,N_13069);
nor U19304 (N_19304,N_12685,N_14765);
nand U19305 (N_19305,N_13962,N_14659);
and U19306 (N_19306,N_12341,N_12551);
nor U19307 (N_19307,N_14825,N_13280);
and U19308 (N_19308,N_14001,N_15922);
or U19309 (N_19309,N_15659,N_14680);
or U19310 (N_19310,N_13912,N_15364);
xor U19311 (N_19311,N_15902,N_13457);
nand U19312 (N_19312,N_14495,N_12274);
xor U19313 (N_19313,N_14842,N_12790);
and U19314 (N_19314,N_14315,N_12763);
or U19315 (N_19315,N_12214,N_12565);
or U19316 (N_19316,N_12825,N_12056);
nand U19317 (N_19317,N_13079,N_15189);
or U19318 (N_19318,N_12975,N_15080);
and U19319 (N_19319,N_15031,N_12436);
or U19320 (N_19320,N_14301,N_13147);
nor U19321 (N_19321,N_15057,N_12435);
and U19322 (N_19322,N_12020,N_12675);
and U19323 (N_19323,N_12602,N_15111);
nand U19324 (N_19324,N_15082,N_15219);
and U19325 (N_19325,N_13502,N_14318);
or U19326 (N_19326,N_15311,N_12793);
xor U19327 (N_19327,N_14290,N_12040);
nor U19328 (N_19328,N_13179,N_12897);
or U19329 (N_19329,N_14980,N_13990);
nand U19330 (N_19330,N_14401,N_13153);
or U19331 (N_19331,N_13764,N_14828);
nor U19332 (N_19332,N_15026,N_15167);
xor U19333 (N_19333,N_13140,N_15037);
xor U19334 (N_19334,N_15820,N_13695);
nor U19335 (N_19335,N_14245,N_13788);
or U19336 (N_19336,N_12324,N_15151);
xor U19337 (N_19337,N_12549,N_14533);
nor U19338 (N_19338,N_13613,N_15589);
xor U19339 (N_19339,N_14955,N_15301);
nor U19340 (N_19340,N_13052,N_15326);
or U19341 (N_19341,N_15938,N_12170);
or U19342 (N_19342,N_15725,N_14518);
nand U19343 (N_19343,N_12035,N_14607);
or U19344 (N_19344,N_15921,N_14202);
nor U19345 (N_19345,N_15058,N_13078);
nor U19346 (N_19346,N_15378,N_15133);
nor U19347 (N_19347,N_15965,N_15855);
xnor U19348 (N_19348,N_13956,N_13264);
nand U19349 (N_19349,N_13538,N_13746);
nor U19350 (N_19350,N_15121,N_14743);
or U19351 (N_19351,N_14414,N_14353);
nand U19352 (N_19352,N_14155,N_14652);
or U19353 (N_19353,N_13970,N_14825);
xor U19354 (N_19354,N_15887,N_13060);
xnor U19355 (N_19355,N_12681,N_12348);
or U19356 (N_19356,N_14763,N_13391);
nor U19357 (N_19357,N_12309,N_13970);
and U19358 (N_19358,N_12254,N_13861);
xor U19359 (N_19359,N_12662,N_15399);
and U19360 (N_19360,N_14367,N_12699);
nand U19361 (N_19361,N_14389,N_13527);
or U19362 (N_19362,N_14559,N_12536);
xor U19363 (N_19363,N_13733,N_14026);
nand U19364 (N_19364,N_15439,N_14657);
xnor U19365 (N_19365,N_15639,N_14878);
nand U19366 (N_19366,N_13547,N_15158);
xor U19367 (N_19367,N_12857,N_14167);
or U19368 (N_19368,N_14629,N_15948);
and U19369 (N_19369,N_14181,N_13520);
and U19370 (N_19370,N_14644,N_14679);
nor U19371 (N_19371,N_13671,N_13941);
nor U19372 (N_19372,N_13999,N_15474);
xnor U19373 (N_19373,N_15430,N_13413);
nor U19374 (N_19374,N_15823,N_12333);
nand U19375 (N_19375,N_13430,N_14731);
nand U19376 (N_19376,N_12531,N_14331);
and U19377 (N_19377,N_12110,N_15688);
nor U19378 (N_19378,N_12939,N_12297);
nor U19379 (N_19379,N_15609,N_15840);
nor U19380 (N_19380,N_14018,N_13033);
nand U19381 (N_19381,N_13897,N_13034);
xor U19382 (N_19382,N_15314,N_13815);
xnor U19383 (N_19383,N_14213,N_12015);
or U19384 (N_19384,N_12270,N_15594);
nand U19385 (N_19385,N_15031,N_14177);
nor U19386 (N_19386,N_14048,N_13425);
and U19387 (N_19387,N_13248,N_12994);
or U19388 (N_19388,N_14420,N_13066);
nand U19389 (N_19389,N_13264,N_14540);
nor U19390 (N_19390,N_12123,N_15297);
and U19391 (N_19391,N_12643,N_15025);
and U19392 (N_19392,N_13030,N_15786);
and U19393 (N_19393,N_12224,N_14307);
or U19394 (N_19394,N_14780,N_13562);
nor U19395 (N_19395,N_13381,N_12368);
nand U19396 (N_19396,N_13512,N_13770);
nor U19397 (N_19397,N_13752,N_13709);
or U19398 (N_19398,N_13024,N_13198);
or U19399 (N_19399,N_15145,N_12400);
and U19400 (N_19400,N_13263,N_12150);
or U19401 (N_19401,N_13259,N_15242);
and U19402 (N_19402,N_13961,N_15015);
xnor U19403 (N_19403,N_13833,N_14435);
and U19404 (N_19404,N_12480,N_12859);
xor U19405 (N_19405,N_13347,N_15876);
and U19406 (N_19406,N_14698,N_12682);
xnor U19407 (N_19407,N_13140,N_15806);
or U19408 (N_19408,N_13272,N_15980);
nand U19409 (N_19409,N_15515,N_12319);
nor U19410 (N_19410,N_13590,N_12618);
and U19411 (N_19411,N_15675,N_12144);
or U19412 (N_19412,N_12524,N_13848);
or U19413 (N_19413,N_14107,N_15233);
nand U19414 (N_19414,N_14288,N_13066);
nand U19415 (N_19415,N_15836,N_14779);
or U19416 (N_19416,N_14385,N_15121);
xor U19417 (N_19417,N_14295,N_15454);
nor U19418 (N_19418,N_14518,N_12309);
nand U19419 (N_19419,N_13494,N_13849);
xnor U19420 (N_19420,N_12280,N_13629);
nand U19421 (N_19421,N_13432,N_14699);
nor U19422 (N_19422,N_12068,N_13846);
nor U19423 (N_19423,N_12122,N_13861);
nor U19424 (N_19424,N_13973,N_13518);
nand U19425 (N_19425,N_15173,N_15803);
or U19426 (N_19426,N_15721,N_14967);
nor U19427 (N_19427,N_13593,N_13251);
or U19428 (N_19428,N_13517,N_15291);
nand U19429 (N_19429,N_14100,N_12723);
and U19430 (N_19430,N_15578,N_15211);
and U19431 (N_19431,N_14412,N_15148);
nand U19432 (N_19432,N_14823,N_15038);
xnor U19433 (N_19433,N_12020,N_14135);
and U19434 (N_19434,N_12580,N_14153);
nor U19435 (N_19435,N_13779,N_13628);
nand U19436 (N_19436,N_13920,N_15601);
nor U19437 (N_19437,N_14165,N_13980);
or U19438 (N_19438,N_14966,N_14908);
or U19439 (N_19439,N_15284,N_14956);
and U19440 (N_19440,N_13232,N_12898);
nand U19441 (N_19441,N_15154,N_12422);
and U19442 (N_19442,N_14912,N_13877);
and U19443 (N_19443,N_15665,N_13180);
and U19444 (N_19444,N_15276,N_15868);
and U19445 (N_19445,N_13917,N_15779);
nor U19446 (N_19446,N_12823,N_15456);
and U19447 (N_19447,N_12878,N_15509);
nor U19448 (N_19448,N_13181,N_13290);
xnor U19449 (N_19449,N_14336,N_13728);
nand U19450 (N_19450,N_12656,N_13728);
nor U19451 (N_19451,N_15982,N_12736);
or U19452 (N_19452,N_12758,N_14424);
or U19453 (N_19453,N_15596,N_13538);
or U19454 (N_19454,N_13638,N_13916);
nor U19455 (N_19455,N_15246,N_12842);
nor U19456 (N_19456,N_15259,N_15427);
xor U19457 (N_19457,N_13570,N_14744);
or U19458 (N_19458,N_13585,N_14622);
and U19459 (N_19459,N_14119,N_12910);
nand U19460 (N_19460,N_12978,N_14348);
nand U19461 (N_19461,N_12845,N_13965);
or U19462 (N_19462,N_13311,N_14940);
nand U19463 (N_19463,N_14739,N_15356);
nor U19464 (N_19464,N_15503,N_13552);
and U19465 (N_19465,N_14693,N_13451);
and U19466 (N_19466,N_14849,N_15038);
or U19467 (N_19467,N_13669,N_14859);
and U19468 (N_19468,N_15740,N_14180);
or U19469 (N_19469,N_14846,N_14635);
nand U19470 (N_19470,N_13828,N_14981);
nor U19471 (N_19471,N_13678,N_15609);
and U19472 (N_19472,N_12414,N_14830);
nand U19473 (N_19473,N_15484,N_14454);
xnor U19474 (N_19474,N_13209,N_14706);
nand U19475 (N_19475,N_14161,N_12809);
nor U19476 (N_19476,N_12052,N_14961);
or U19477 (N_19477,N_13672,N_14114);
xnor U19478 (N_19478,N_13908,N_12544);
and U19479 (N_19479,N_14748,N_12227);
nand U19480 (N_19480,N_12866,N_15373);
or U19481 (N_19481,N_14844,N_14765);
nor U19482 (N_19482,N_12732,N_12443);
xor U19483 (N_19483,N_15402,N_15303);
nand U19484 (N_19484,N_15927,N_13399);
nor U19485 (N_19485,N_13143,N_14294);
and U19486 (N_19486,N_13412,N_13301);
and U19487 (N_19487,N_13978,N_13134);
xnor U19488 (N_19488,N_13109,N_13718);
xnor U19489 (N_19489,N_15978,N_15378);
xor U19490 (N_19490,N_12450,N_12422);
or U19491 (N_19491,N_13412,N_14745);
xor U19492 (N_19492,N_14442,N_12731);
or U19493 (N_19493,N_14636,N_13032);
or U19494 (N_19494,N_12117,N_15114);
xor U19495 (N_19495,N_15375,N_13966);
nor U19496 (N_19496,N_14758,N_14289);
nand U19497 (N_19497,N_12555,N_15960);
nand U19498 (N_19498,N_12259,N_14957);
xnor U19499 (N_19499,N_15944,N_12790);
nand U19500 (N_19500,N_13898,N_15191);
or U19501 (N_19501,N_13279,N_15860);
and U19502 (N_19502,N_13783,N_12491);
nand U19503 (N_19503,N_14589,N_13109);
xor U19504 (N_19504,N_12357,N_12107);
and U19505 (N_19505,N_13158,N_12448);
nand U19506 (N_19506,N_15015,N_13794);
nand U19507 (N_19507,N_13841,N_12460);
xnor U19508 (N_19508,N_14879,N_14521);
nand U19509 (N_19509,N_14086,N_15298);
xor U19510 (N_19510,N_13944,N_14536);
or U19511 (N_19511,N_12807,N_12833);
nand U19512 (N_19512,N_15244,N_14265);
or U19513 (N_19513,N_12708,N_12297);
nand U19514 (N_19514,N_13313,N_14335);
nand U19515 (N_19515,N_12424,N_15422);
and U19516 (N_19516,N_13134,N_14920);
or U19517 (N_19517,N_15076,N_14984);
or U19518 (N_19518,N_12911,N_14715);
xnor U19519 (N_19519,N_13195,N_13674);
xor U19520 (N_19520,N_14485,N_14578);
xnor U19521 (N_19521,N_14547,N_15338);
xnor U19522 (N_19522,N_12097,N_15001);
nor U19523 (N_19523,N_15510,N_12114);
nand U19524 (N_19524,N_12315,N_14155);
or U19525 (N_19525,N_14683,N_15032);
or U19526 (N_19526,N_15964,N_12335);
nor U19527 (N_19527,N_15237,N_15375);
xnor U19528 (N_19528,N_12968,N_13604);
nor U19529 (N_19529,N_14936,N_14724);
nor U19530 (N_19530,N_15538,N_15965);
or U19531 (N_19531,N_13901,N_12048);
nand U19532 (N_19532,N_14421,N_15995);
xnor U19533 (N_19533,N_14379,N_12110);
and U19534 (N_19534,N_15580,N_15607);
nor U19535 (N_19535,N_15571,N_12061);
or U19536 (N_19536,N_15079,N_15924);
nor U19537 (N_19537,N_15587,N_12044);
or U19538 (N_19538,N_13253,N_15644);
and U19539 (N_19539,N_15449,N_15259);
nor U19540 (N_19540,N_14288,N_14820);
and U19541 (N_19541,N_15056,N_13782);
or U19542 (N_19542,N_12587,N_14468);
nor U19543 (N_19543,N_15685,N_14723);
nor U19544 (N_19544,N_13331,N_15287);
nor U19545 (N_19545,N_15315,N_15578);
and U19546 (N_19546,N_13858,N_12671);
nand U19547 (N_19547,N_12047,N_13970);
xnor U19548 (N_19548,N_14727,N_15771);
and U19549 (N_19549,N_14154,N_15980);
and U19550 (N_19550,N_14293,N_14116);
and U19551 (N_19551,N_13952,N_15317);
nand U19552 (N_19552,N_12636,N_14093);
nand U19553 (N_19553,N_13913,N_15105);
nor U19554 (N_19554,N_14037,N_12592);
nor U19555 (N_19555,N_15678,N_15574);
nor U19556 (N_19556,N_12142,N_15246);
and U19557 (N_19557,N_15944,N_13481);
nor U19558 (N_19558,N_14190,N_15205);
or U19559 (N_19559,N_15828,N_15337);
nand U19560 (N_19560,N_14887,N_12520);
xnor U19561 (N_19561,N_15861,N_15123);
nand U19562 (N_19562,N_12249,N_12893);
or U19563 (N_19563,N_13331,N_12453);
xor U19564 (N_19564,N_13342,N_14504);
and U19565 (N_19565,N_12934,N_12853);
nand U19566 (N_19566,N_12465,N_15362);
or U19567 (N_19567,N_12096,N_13537);
nand U19568 (N_19568,N_15683,N_15361);
xor U19569 (N_19569,N_12876,N_14874);
xnor U19570 (N_19570,N_12566,N_12743);
nand U19571 (N_19571,N_13694,N_13516);
nand U19572 (N_19572,N_13079,N_13983);
or U19573 (N_19573,N_12661,N_14371);
and U19574 (N_19574,N_12401,N_15804);
nand U19575 (N_19575,N_12378,N_15471);
xnor U19576 (N_19576,N_15370,N_12492);
or U19577 (N_19577,N_12213,N_13287);
nor U19578 (N_19578,N_12376,N_14358);
and U19579 (N_19579,N_14539,N_12560);
nand U19580 (N_19580,N_13754,N_15137);
xnor U19581 (N_19581,N_12762,N_14997);
xnor U19582 (N_19582,N_15342,N_13244);
or U19583 (N_19583,N_14443,N_15538);
nand U19584 (N_19584,N_13474,N_14607);
nand U19585 (N_19585,N_14920,N_15195);
nor U19586 (N_19586,N_13187,N_12938);
or U19587 (N_19587,N_15255,N_13564);
nand U19588 (N_19588,N_13286,N_12518);
and U19589 (N_19589,N_14043,N_15618);
nor U19590 (N_19590,N_12210,N_13548);
nand U19591 (N_19591,N_13097,N_14444);
and U19592 (N_19592,N_15221,N_14923);
nand U19593 (N_19593,N_12876,N_15404);
xnor U19594 (N_19594,N_13946,N_12334);
xor U19595 (N_19595,N_13739,N_13403);
and U19596 (N_19596,N_12221,N_14126);
or U19597 (N_19597,N_13279,N_12972);
nor U19598 (N_19598,N_14275,N_13879);
nand U19599 (N_19599,N_15641,N_14273);
nor U19600 (N_19600,N_12195,N_13144);
and U19601 (N_19601,N_14749,N_15944);
nand U19602 (N_19602,N_12862,N_13082);
or U19603 (N_19603,N_12500,N_14978);
nand U19604 (N_19604,N_13591,N_14832);
xor U19605 (N_19605,N_15730,N_13876);
nor U19606 (N_19606,N_14913,N_15745);
xnor U19607 (N_19607,N_12329,N_14391);
xor U19608 (N_19608,N_15126,N_12271);
or U19609 (N_19609,N_12220,N_13866);
nor U19610 (N_19610,N_15268,N_14552);
nor U19611 (N_19611,N_12374,N_15045);
nand U19612 (N_19612,N_12719,N_15222);
and U19613 (N_19613,N_14178,N_14738);
or U19614 (N_19614,N_13275,N_12101);
and U19615 (N_19615,N_12516,N_12062);
or U19616 (N_19616,N_13923,N_15049);
or U19617 (N_19617,N_15711,N_14656);
and U19618 (N_19618,N_15075,N_13223);
nand U19619 (N_19619,N_14271,N_12819);
nand U19620 (N_19620,N_12094,N_14640);
nand U19621 (N_19621,N_14451,N_15196);
and U19622 (N_19622,N_15469,N_13957);
nand U19623 (N_19623,N_12727,N_14234);
and U19624 (N_19624,N_15351,N_13528);
nand U19625 (N_19625,N_15385,N_13412);
xor U19626 (N_19626,N_14549,N_13222);
and U19627 (N_19627,N_15798,N_14188);
nand U19628 (N_19628,N_13436,N_15368);
xor U19629 (N_19629,N_15096,N_12762);
xnor U19630 (N_19630,N_13924,N_12745);
nor U19631 (N_19631,N_15484,N_12146);
and U19632 (N_19632,N_13703,N_15989);
nand U19633 (N_19633,N_15581,N_12285);
or U19634 (N_19634,N_13315,N_15697);
nand U19635 (N_19635,N_14208,N_13414);
or U19636 (N_19636,N_12399,N_13637);
and U19637 (N_19637,N_15340,N_14150);
and U19638 (N_19638,N_14285,N_14142);
nor U19639 (N_19639,N_13454,N_15979);
or U19640 (N_19640,N_13013,N_13300);
nor U19641 (N_19641,N_12088,N_15027);
xnor U19642 (N_19642,N_15262,N_15549);
nor U19643 (N_19643,N_14054,N_15754);
nand U19644 (N_19644,N_12295,N_13998);
nor U19645 (N_19645,N_12959,N_14900);
nor U19646 (N_19646,N_12438,N_15939);
nand U19647 (N_19647,N_12910,N_14439);
nand U19648 (N_19648,N_12153,N_15413);
xor U19649 (N_19649,N_14425,N_13265);
xnor U19650 (N_19650,N_12633,N_12072);
xnor U19651 (N_19651,N_13856,N_15739);
or U19652 (N_19652,N_15119,N_13851);
nor U19653 (N_19653,N_12341,N_13059);
xnor U19654 (N_19654,N_12300,N_13011);
and U19655 (N_19655,N_14019,N_13809);
nand U19656 (N_19656,N_14051,N_12376);
nand U19657 (N_19657,N_14338,N_13429);
and U19658 (N_19658,N_12779,N_13062);
nand U19659 (N_19659,N_14394,N_14829);
xnor U19660 (N_19660,N_15506,N_12906);
xor U19661 (N_19661,N_12377,N_12071);
and U19662 (N_19662,N_13416,N_15904);
nand U19663 (N_19663,N_13379,N_14586);
nor U19664 (N_19664,N_12995,N_15344);
nor U19665 (N_19665,N_13935,N_15670);
xnor U19666 (N_19666,N_14225,N_12586);
nand U19667 (N_19667,N_14410,N_14294);
nand U19668 (N_19668,N_14949,N_15640);
and U19669 (N_19669,N_13342,N_13072);
and U19670 (N_19670,N_12572,N_15848);
nand U19671 (N_19671,N_15919,N_13424);
and U19672 (N_19672,N_14428,N_14258);
nand U19673 (N_19673,N_13359,N_15101);
and U19674 (N_19674,N_15781,N_14617);
or U19675 (N_19675,N_13462,N_15978);
nor U19676 (N_19676,N_13273,N_12176);
and U19677 (N_19677,N_13098,N_14722);
xnor U19678 (N_19678,N_12458,N_14294);
nor U19679 (N_19679,N_12231,N_14460);
nand U19680 (N_19680,N_13852,N_12689);
nand U19681 (N_19681,N_13823,N_13558);
nand U19682 (N_19682,N_14656,N_15660);
xor U19683 (N_19683,N_14597,N_12883);
nand U19684 (N_19684,N_15376,N_15588);
nand U19685 (N_19685,N_13725,N_13297);
and U19686 (N_19686,N_14563,N_15051);
and U19687 (N_19687,N_14727,N_12776);
or U19688 (N_19688,N_13531,N_12146);
nand U19689 (N_19689,N_13994,N_15515);
nand U19690 (N_19690,N_12163,N_13200);
nand U19691 (N_19691,N_12961,N_13249);
nand U19692 (N_19692,N_14393,N_15253);
and U19693 (N_19693,N_14266,N_14260);
or U19694 (N_19694,N_12620,N_14964);
and U19695 (N_19695,N_12128,N_15936);
nor U19696 (N_19696,N_15706,N_13208);
and U19697 (N_19697,N_15695,N_14701);
nand U19698 (N_19698,N_12186,N_14265);
or U19699 (N_19699,N_14974,N_14196);
xnor U19700 (N_19700,N_14128,N_14853);
and U19701 (N_19701,N_14549,N_15374);
nand U19702 (N_19702,N_14908,N_14116);
or U19703 (N_19703,N_13308,N_14630);
xor U19704 (N_19704,N_12229,N_13745);
nand U19705 (N_19705,N_15330,N_14054);
or U19706 (N_19706,N_12276,N_12559);
nor U19707 (N_19707,N_15484,N_14710);
or U19708 (N_19708,N_12575,N_13205);
nand U19709 (N_19709,N_13827,N_14626);
or U19710 (N_19710,N_14928,N_14657);
nand U19711 (N_19711,N_15881,N_15983);
and U19712 (N_19712,N_13420,N_14852);
xor U19713 (N_19713,N_15643,N_12877);
or U19714 (N_19714,N_12703,N_13211);
nor U19715 (N_19715,N_12621,N_12990);
xor U19716 (N_19716,N_15753,N_15361);
and U19717 (N_19717,N_14015,N_14646);
nand U19718 (N_19718,N_15916,N_15853);
nand U19719 (N_19719,N_13162,N_14964);
nor U19720 (N_19720,N_14247,N_14818);
and U19721 (N_19721,N_12983,N_13646);
xor U19722 (N_19722,N_13853,N_13994);
xnor U19723 (N_19723,N_13526,N_12618);
and U19724 (N_19724,N_13954,N_15858);
nor U19725 (N_19725,N_15517,N_13384);
and U19726 (N_19726,N_14370,N_13367);
xor U19727 (N_19727,N_12659,N_13005);
nand U19728 (N_19728,N_13334,N_13671);
nor U19729 (N_19729,N_13428,N_12786);
and U19730 (N_19730,N_15623,N_15321);
or U19731 (N_19731,N_15677,N_14909);
nor U19732 (N_19732,N_14897,N_13340);
or U19733 (N_19733,N_15964,N_14946);
or U19734 (N_19734,N_13521,N_14761);
nor U19735 (N_19735,N_13589,N_12851);
xnor U19736 (N_19736,N_15873,N_14654);
xor U19737 (N_19737,N_14299,N_14605);
xnor U19738 (N_19738,N_12824,N_15853);
and U19739 (N_19739,N_13259,N_14451);
and U19740 (N_19740,N_15045,N_15527);
nand U19741 (N_19741,N_13004,N_15267);
or U19742 (N_19742,N_14288,N_13411);
xnor U19743 (N_19743,N_15814,N_14226);
nor U19744 (N_19744,N_14903,N_15544);
or U19745 (N_19745,N_12710,N_12330);
nand U19746 (N_19746,N_14790,N_15601);
xnor U19747 (N_19747,N_13118,N_15216);
nand U19748 (N_19748,N_14450,N_12111);
and U19749 (N_19749,N_15103,N_13859);
xor U19750 (N_19750,N_12220,N_12932);
xnor U19751 (N_19751,N_13317,N_13915);
nor U19752 (N_19752,N_14733,N_14813);
nor U19753 (N_19753,N_13865,N_12560);
nand U19754 (N_19754,N_12468,N_12906);
nand U19755 (N_19755,N_14814,N_12775);
and U19756 (N_19756,N_14099,N_12392);
xnor U19757 (N_19757,N_14990,N_13033);
nor U19758 (N_19758,N_13674,N_12718);
nor U19759 (N_19759,N_13289,N_15030);
and U19760 (N_19760,N_12986,N_12833);
nor U19761 (N_19761,N_14385,N_15463);
nand U19762 (N_19762,N_12104,N_14699);
nand U19763 (N_19763,N_13239,N_12491);
or U19764 (N_19764,N_12152,N_13489);
and U19765 (N_19765,N_14267,N_15642);
nand U19766 (N_19766,N_15919,N_12282);
and U19767 (N_19767,N_12957,N_12847);
nor U19768 (N_19768,N_13326,N_12269);
and U19769 (N_19769,N_13753,N_12780);
nor U19770 (N_19770,N_15989,N_14442);
and U19771 (N_19771,N_12311,N_13273);
nand U19772 (N_19772,N_12571,N_14655);
and U19773 (N_19773,N_13074,N_12708);
nand U19774 (N_19774,N_13314,N_13622);
xnor U19775 (N_19775,N_15897,N_14948);
or U19776 (N_19776,N_15845,N_12619);
or U19777 (N_19777,N_15663,N_13918);
nand U19778 (N_19778,N_13909,N_12364);
xor U19779 (N_19779,N_12861,N_12807);
nor U19780 (N_19780,N_12992,N_13899);
and U19781 (N_19781,N_15533,N_13274);
nand U19782 (N_19782,N_14194,N_15952);
and U19783 (N_19783,N_12015,N_13696);
or U19784 (N_19784,N_15987,N_13900);
and U19785 (N_19785,N_14775,N_15699);
xor U19786 (N_19786,N_12054,N_12796);
nor U19787 (N_19787,N_13063,N_14962);
or U19788 (N_19788,N_13069,N_14916);
xnor U19789 (N_19789,N_12739,N_14638);
xor U19790 (N_19790,N_12263,N_12625);
or U19791 (N_19791,N_15144,N_14255);
nand U19792 (N_19792,N_14237,N_15530);
nor U19793 (N_19793,N_12235,N_14814);
nor U19794 (N_19794,N_13800,N_12206);
nor U19795 (N_19795,N_13703,N_13813);
xnor U19796 (N_19796,N_15183,N_13186);
nor U19797 (N_19797,N_14538,N_12235);
or U19798 (N_19798,N_12653,N_14425);
and U19799 (N_19799,N_14281,N_14240);
nand U19800 (N_19800,N_12016,N_15477);
xnor U19801 (N_19801,N_14135,N_14845);
xnor U19802 (N_19802,N_13667,N_12814);
nor U19803 (N_19803,N_15398,N_14890);
xor U19804 (N_19804,N_14825,N_14201);
or U19805 (N_19805,N_13023,N_14930);
and U19806 (N_19806,N_14290,N_14318);
nand U19807 (N_19807,N_14217,N_12292);
nor U19808 (N_19808,N_13785,N_15648);
or U19809 (N_19809,N_12047,N_15600);
or U19810 (N_19810,N_15363,N_13621);
or U19811 (N_19811,N_12756,N_15958);
xnor U19812 (N_19812,N_12138,N_15272);
or U19813 (N_19813,N_12275,N_13337);
or U19814 (N_19814,N_15469,N_13865);
xnor U19815 (N_19815,N_15530,N_12129);
xnor U19816 (N_19816,N_14583,N_15514);
and U19817 (N_19817,N_13129,N_13983);
or U19818 (N_19818,N_13204,N_13703);
xor U19819 (N_19819,N_15917,N_12609);
nor U19820 (N_19820,N_14331,N_15248);
nand U19821 (N_19821,N_13147,N_13057);
and U19822 (N_19822,N_14950,N_14702);
nor U19823 (N_19823,N_12081,N_14035);
xnor U19824 (N_19824,N_15376,N_15221);
nor U19825 (N_19825,N_12076,N_15416);
nor U19826 (N_19826,N_13234,N_15166);
nand U19827 (N_19827,N_12989,N_15604);
nor U19828 (N_19828,N_14594,N_13149);
nand U19829 (N_19829,N_14041,N_12848);
nand U19830 (N_19830,N_12486,N_12540);
nand U19831 (N_19831,N_12069,N_13259);
xnor U19832 (N_19832,N_13430,N_14898);
or U19833 (N_19833,N_15644,N_12494);
xor U19834 (N_19834,N_13462,N_14878);
nor U19835 (N_19835,N_13914,N_12796);
nor U19836 (N_19836,N_12491,N_12006);
xor U19837 (N_19837,N_15601,N_13654);
nand U19838 (N_19838,N_12713,N_14380);
nor U19839 (N_19839,N_13757,N_13658);
or U19840 (N_19840,N_12627,N_12286);
xnor U19841 (N_19841,N_14516,N_13842);
nor U19842 (N_19842,N_14465,N_13548);
and U19843 (N_19843,N_15587,N_12550);
nand U19844 (N_19844,N_15652,N_12927);
and U19845 (N_19845,N_14910,N_12055);
nand U19846 (N_19846,N_12101,N_15229);
xnor U19847 (N_19847,N_14403,N_13719);
nand U19848 (N_19848,N_14291,N_13345);
xnor U19849 (N_19849,N_12230,N_15113);
or U19850 (N_19850,N_12142,N_15357);
nor U19851 (N_19851,N_12177,N_14615);
xnor U19852 (N_19852,N_13057,N_14379);
and U19853 (N_19853,N_14633,N_15571);
nor U19854 (N_19854,N_12048,N_15558);
nor U19855 (N_19855,N_14945,N_14387);
or U19856 (N_19856,N_13995,N_15482);
and U19857 (N_19857,N_14425,N_14579);
and U19858 (N_19858,N_14657,N_15141);
or U19859 (N_19859,N_13894,N_14940);
nand U19860 (N_19860,N_15715,N_15721);
nor U19861 (N_19861,N_12652,N_15291);
and U19862 (N_19862,N_15712,N_13845);
nor U19863 (N_19863,N_12206,N_12096);
nand U19864 (N_19864,N_12933,N_14398);
nor U19865 (N_19865,N_14183,N_14202);
nand U19866 (N_19866,N_15569,N_13155);
nand U19867 (N_19867,N_14149,N_13791);
xnor U19868 (N_19868,N_12769,N_13416);
or U19869 (N_19869,N_13091,N_12886);
xnor U19870 (N_19870,N_13447,N_15527);
nor U19871 (N_19871,N_12003,N_15708);
nor U19872 (N_19872,N_15770,N_13301);
or U19873 (N_19873,N_15902,N_14191);
nor U19874 (N_19874,N_13258,N_13629);
nor U19875 (N_19875,N_14808,N_15270);
and U19876 (N_19876,N_13084,N_13256);
nor U19877 (N_19877,N_15278,N_14894);
or U19878 (N_19878,N_12194,N_13028);
nand U19879 (N_19879,N_13115,N_14461);
and U19880 (N_19880,N_12349,N_13680);
or U19881 (N_19881,N_12383,N_14020);
nand U19882 (N_19882,N_14822,N_12797);
or U19883 (N_19883,N_14699,N_12229);
nor U19884 (N_19884,N_14025,N_13494);
nor U19885 (N_19885,N_15986,N_15286);
xnor U19886 (N_19886,N_15348,N_13702);
and U19887 (N_19887,N_14752,N_12884);
and U19888 (N_19888,N_13093,N_12937);
nor U19889 (N_19889,N_15059,N_13628);
xnor U19890 (N_19890,N_15706,N_13783);
and U19891 (N_19891,N_15291,N_13598);
or U19892 (N_19892,N_15586,N_15973);
nand U19893 (N_19893,N_12101,N_12488);
xnor U19894 (N_19894,N_15082,N_12302);
xor U19895 (N_19895,N_13672,N_13865);
nand U19896 (N_19896,N_12326,N_12307);
xnor U19897 (N_19897,N_13177,N_14959);
xor U19898 (N_19898,N_14568,N_12841);
or U19899 (N_19899,N_12832,N_14379);
nor U19900 (N_19900,N_14952,N_12099);
nand U19901 (N_19901,N_14513,N_12292);
nor U19902 (N_19902,N_12932,N_14927);
xor U19903 (N_19903,N_14387,N_14028);
or U19904 (N_19904,N_12891,N_14031);
or U19905 (N_19905,N_14131,N_15187);
or U19906 (N_19906,N_13527,N_15688);
nand U19907 (N_19907,N_13178,N_12520);
or U19908 (N_19908,N_15381,N_12448);
nor U19909 (N_19909,N_15898,N_14829);
nor U19910 (N_19910,N_12139,N_12473);
or U19911 (N_19911,N_14606,N_14134);
and U19912 (N_19912,N_15927,N_13821);
or U19913 (N_19913,N_14726,N_14729);
or U19914 (N_19914,N_13968,N_13342);
xor U19915 (N_19915,N_14406,N_12230);
nand U19916 (N_19916,N_13324,N_14546);
and U19917 (N_19917,N_15412,N_14352);
xor U19918 (N_19918,N_12680,N_13357);
xor U19919 (N_19919,N_12362,N_13515);
xor U19920 (N_19920,N_14675,N_12313);
xnor U19921 (N_19921,N_13421,N_14551);
and U19922 (N_19922,N_15999,N_13795);
and U19923 (N_19923,N_14503,N_12588);
or U19924 (N_19924,N_13891,N_14558);
nand U19925 (N_19925,N_12089,N_15833);
and U19926 (N_19926,N_14146,N_15894);
xnor U19927 (N_19927,N_13686,N_15873);
xnor U19928 (N_19928,N_12412,N_14988);
and U19929 (N_19929,N_15905,N_14971);
or U19930 (N_19930,N_12956,N_12444);
and U19931 (N_19931,N_13071,N_12656);
xor U19932 (N_19932,N_15516,N_14659);
nor U19933 (N_19933,N_13995,N_12754);
nand U19934 (N_19934,N_14982,N_15404);
and U19935 (N_19935,N_13388,N_15968);
xnor U19936 (N_19936,N_15812,N_14366);
xor U19937 (N_19937,N_13615,N_15705);
nand U19938 (N_19938,N_15830,N_14932);
xor U19939 (N_19939,N_15081,N_14290);
nand U19940 (N_19940,N_14028,N_14515);
or U19941 (N_19941,N_14146,N_15612);
xor U19942 (N_19942,N_12230,N_13714);
or U19943 (N_19943,N_14177,N_12349);
and U19944 (N_19944,N_12861,N_13799);
nand U19945 (N_19945,N_14143,N_14527);
or U19946 (N_19946,N_13668,N_13638);
xnor U19947 (N_19947,N_14528,N_13192);
and U19948 (N_19948,N_13306,N_13859);
and U19949 (N_19949,N_15079,N_15988);
or U19950 (N_19950,N_12107,N_14775);
xnor U19951 (N_19951,N_14966,N_12874);
or U19952 (N_19952,N_14737,N_12802);
nand U19953 (N_19953,N_12651,N_14818);
nor U19954 (N_19954,N_13150,N_14328);
nor U19955 (N_19955,N_12893,N_15314);
and U19956 (N_19956,N_14203,N_12727);
or U19957 (N_19957,N_14179,N_14706);
nor U19958 (N_19958,N_14572,N_14695);
nand U19959 (N_19959,N_15340,N_13408);
nand U19960 (N_19960,N_12467,N_13454);
xnor U19961 (N_19961,N_13707,N_13975);
nand U19962 (N_19962,N_13051,N_12290);
nor U19963 (N_19963,N_13558,N_14275);
or U19964 (N_19964,N_14342,N_12675);
nand U19965 (N_19965,N_15299,N_12148);
and U19966 (N_19966,N_13219,N_14019);
or U19967 (N_19967,N_14086,N_13585);
nor U19968 (N_19968,N_13752,N_12428);
or U19969 (N_19969,N_15959,N_15990);
nor U19970 (N_19970,N_15443,N_12432);
xor U19971 (N_19971,N_14144,N_15965);
or U19972 (N_19972,N_14546,N_13345);
or U19973 (N_19973,N_13778,N_13528);
nand U19974 (N_19974,N_12102,N_12034);
nor U19975 (N_19975,N_12412,N_14474);
nand U19976 (N_19976,N_13701,N_14034);
nand U19977 (N_19977,N_12929,N_15016);
or U19978 (N_19978,N_15229,N_14942);
xnor U19979 (N_19979,N_14879,N_12965);
or U19980 (N_19980,N_12163,N_13921);
nand U19981 (N_19981,N_15376,N_15766);
or U19982 (N_19982,N_15850,N_15176);
xnor U19983 (N_19983,N_14292,N_13344);
or U19984 (N_19984,N_12955,N_14859);
nand U19985 (N_19985,N_13051,N_12196);
or U19986 (N_19986,N_13873,N_12671);
xnor U19987 (N_19987,N_15283,N_13842);
xor U19988 (N_19988,N_15100,N_15073);
nand U19989 (N_19989,N_13022,N_14020);
and U19990 (N_19990,N_15121,N_14691);
nor U19991 (N_19991,N_14851,N_14003);
xnor U19992 (N_19992,N_13789,N_14577);
or U19993 (N_19993,N_12432,N_12587);
xor U19994 (N_19994,N_13674,N_14610);
nor U19995 (N_19995,N_15806,N_13332);
and U19996 (N_19996,N_14671,N_15672);
and U19997 (N_19997,N_14191,N_15331);
xnor U19998 (N_19998,N_12518,N_14216);
xnor U19999 (N_19999,N_15043,N_12464);
nand UO_0 (O_0,N_17536,N_19735);
nand UO_1 (O_1,N_16947,N_16648);
or UO_2 (O_2,N_16328,N_18848);
or UO_3 (O_3,N_17084,N_17156);
nor UO_4 (O_4,N_16730,N_19216);
and UO_5 (O_5,N_16080,N_16229);
or UO_6 (O_6,N_17723,N_18030);
or UO_7 (O_7,N_16275,N_19814);
nor UO_8 (O_8,N_16764,N_18738);
or UO_9 (O_9,N_19780,N_18752);
or UO_10 (O_10,N_16912,N_17042);
nand UO_11 (O_11,N_16369,N_16627);
and UO_12 (O_12,N_16313,N_19956);
or UO_13 (O_13,N_17123,N_19120);
and UO_14 (O_14,N_17659,N_19922);
xnor UO_15 (O_15,N_18607,N_16495);
and UO_16 (O_16,N_18514,N_18882);
and UO_17 (O_17,N_19830,N_19247);
nor UO_18 (O_18,N_17622,N_17615);
xor UO_19 (O_19,N_19519,N_19740);
nor UO_20 (O_20,N_19777,N_16344);
and UO_21 (O_21,N_18739,N_17891);
and UO_22 (O_22,N_18491,N_19374);
nand UO_23 (O_23,N_19803,N_17550);
nor UO_24 (O_24,N_16476,N_17218);
nand UO_25 (O_25,N_16432,N_18944);
nand UO_26 (O_26,N_17837,N_18158);
nor UO_27 (O_27,N_16854,N_16415);
xnor UO_28 (O_28,N_17259,N_16645);
xor UO_29 (O_29,N_16786,N_17649);
or UO_30 (O_30,N_18255,N_16209);
or UO_31 (O_31,N_17476,N_16750);
nor UO_32 (O_32,N_19020,N_18400);
nor UO_33 (O_33,N_17966,N_16021);
and UO_34 (O_34,N_17117,N_17493);
nor UO_35 (O_35,N_19222,N_16761);
xor UO_36 (O_36,N_17444,N_19415);
nor UO_37 (O_37,N_18122,N_19187);
or UO_38 (O_38,N_18991,N_16383);
and UO_39 (O_39,N_19698,N_17355);
xor UO_40 (O_40,N_17288,N_19496);
nor UO_41 (O_41,N_17268,N_17680);
and UO_42 (O_42,N_18694,N_18317);
and UO_43 (O_43,N_19508,N_17544);
nor UO_44 (O_44,N_18090,N_18154);
nand UO_45 (O_45,N_17818,N_16309);
and UO_46 (O_46,N_19224,N_16636);
nor UO_47 (O_47,N_17691,N_18722);
xnor UO_48 (O_48,N_18675,N_17369);
nand UO_49 (O_49,N_17667,N_17749);
and UO_50 (O_50,N_18241,N_16715);
nand UO_51 (O_51,N_18532,N_19254);
nand UO_52 (O_52,N_17535,N_17471);
and UO_53 (O_53,N_16401,N_17020);
nand UO_54 (O_54,N_16898,N_18492);
nor UO_55 (O_55,N_16033,N_16791);
nor UO_56 (O_56,N_17154,N_16129);
nand UO_57 (O_57,N_18399,N_19458);
and UO_58 (O_58,N_17706,N_19536);
and UO_59 (O_59,N_16671,N_19255);
nor UO_60 (O_60,N_18684,N_16258);
nor UO_61 (O_61,N_16113,N_16219);
and UO_62 (O_62,N_19721,N_16953);
nor UO_63 (O_63,N_18434,N_16980);
or UO_64 (O_64,N_16701,N_19895);
nor UO_65 (O_65,N_17119,N_18656);
xor UO_66 (O_66,N_18669,N_17423);
or UO_67 (O_67,N_18717,N_16324);
xnor UO_68 (O_68,N_18188,N_19694);
and UO_69 (O_69,N_16649,N_16011);
nand UO_70 (O_70,N_18518,N_18334);
nand UO_71 (O_71,N_16540,N_17373);
nand UO_72 (O_72,N_18945,N_16558);
or UO_73 (O_73,N_17756,N_19589);
or UO_74 (O_74,N_17167,N_19165);
xnor UO_75 (O_75,N_16465,N_18998);
nor UO_76 (O_76,N_19543,N_17008);
xor UO_77 (O_77,N_16569,N_19034);
and UO_78 (O_78,N_17990,N_19979);
or UO_79 (O_79,N_18558,N_16420);
nor UO_80 (O_80,N_17063,N_18500);
and UO_81 (O_81,N_19520,N_17525);
xnor UO_82 (O_82,N_17334,N_19865);
and UO_83 (O_83,N_18825,N_19331);
nand UO_84 (O_84,N_18450,N_18353);
or UO_85 (O_85,N_17343,N_17301);
and UO_86 (O_86,N_18105,N_16363);
and UO_87 (O_87,N_16343,N_18925);
or UO_88 (O_88,N_19320,N_18615);
xor UO_89 (O_89,N_17552,N_19928);
nor UO_90 (O_90,N_18181,N_17974);
xor UO_91 (O_91,N_16721,N_18469);
xor UO_92 (O_92,N_16873,N_17512);
xor UO_93 (O_93,N_16990,N_19510);
nor UO_94 (O_94,N_19964,N_17505);
or UO_95 (O_95,N_18690,N_18053);
nand UO_96 (O_96,N_17932,N_17068);
and UO_97 (O_97,N_17260,N_19731);
or UO_98 (O_98,N_17572,N_17242);
or UO_99 (O_99,N_18905,N_17443);
and UO_100 (O_100,N_18594,N_19884);
or UO_101 (O_101,N_19432,N_18830);
nand UO_102 (O_102,N_19974,N_17037);
xnor UO_103 (O_103,N_18017,N_19491);
and UO_104 (O_104,N_16187,N_18600);
nand UO_105 (O_105,N_17366,N_18680);
xnor UO_106 (O_106,N_17888,N_18130);
nand UO_107 (O_107,N_19977,N_18039);
nand UO_108 (O_108,N_16417,N_17670);
xor UO_109 (O_109,N_17780,N_18929);
or UO_110 (O_110,N_19565,N_19976);
or UO_111 (O_111,N_18796,N_19801);
and UO_112 (O_112,N_17832,N_16793);
nor UO_113 (O_113,N_16632,N_19675);
or UO_114 (O_114,N_18901,N_17120);
nor UO_115 (O_115,N_19604,N_18100);
or UO_116 (O_116,N_18144,N_17652);
nand UO_117 (O_117,N_16712,N_17580);
nand UO_118 (O_118,N_16248,N_19837);
xor UO_119 (O_119,N_19072,N_19963);
nor UO_120 (O_120,N_17675,N_17470);
nor UO_121 (O_121,N_19016,N_17795);
or UO_122 (O_122,N_18716,N_17111);
nand UO_123 (O_123,N_17569,N_19620);
xnor UO_124 (O_124,N_19524,N_19853);
xnor UO_125 (O_125,N_19628,N_19443);
nand UO_126 (O_126,N_17308,N_19258);
nand UO_127 (O_127,N_17735,N_18545);
nor UO_128 (O_128,N_17897,N_16546);
nand UO_129 (O_129,N_18623,N_18183);
and UO_130 (O_130,N_19166,N_18390);
xnor UO_131 (O_131,N_19397,N_19419);
nand UO_132 (O_132,N_18613,N_19232);
xor UO_133 (O_133,N_16245,N_17968);
xnor UO_134 (O_134,N_16002,N_19587);
or UO_135 (O_135,N_18475,N_18233);
or UO_136 (O_136,N_17320,N_19344);
nand UO_137 (O_137,N_17657,N_16646);
and UO_138 (O_138,N_17029,N_17087);
xnor UO_139 (O_139,N_16463,N_17671);
nor UO_140 (O_140,N_18461,N_17710);
nor UO_141 (O_141,N_19681,N_19714);
or UO_142 (O_142,N_18422,N_18194);
nor UO_143 (O_143,N_17985,N_17781);
xor UO_144 (O_144,N_18869,N_19493);
nand UO_145 (O_145,N_17944,N_18969);
nor UO_146 (O_146,N_17703,N_16138);
or UO_147 (O_147,N_16823,N_19026);
or UO_148 (O_148,N_19109,N_16342);
or UO_149 (O_149,N_18187,N_17921);
or UO_150 (O_150,N_18298,N_19215);
nor UO_151 (O_151,N_18127,N_17739);
nand UO_152 (O_152,N_19993,N_18078);
nand UO_153 (O_153,N_18780,N_16973);
and UO_154 (O_154,N_16287,N_17053);
nand UO_155 (O_155,N_16616,N_16188);
and UO_156 (O_156,N_17618,N_19051);
and UO_157 (O_157,N_16181,N_16836);
and UO_158 (O_158,N_19229,N_19248);
xor UO_159 (O_159,N_16135,N_17656);
and UO_160 (O_160,N_17959,N_16154);
nor UO_161 (O_161,N_18795,N_18295);
or UO_162 (O_162,N_18849,N_16625);
nand UO_163 (O_163,N_16095,N_17549);
nor UO_164 (O_164,N_19386,N_16934);
nor UO_165 (O_165,N_17876,N_19365);
nor UO_166 (O_166,N_16565,N_19502);
and UO_167 (O_167,N_17193,N_19151);
nor UO_168 (O_168,N_19287,N_17174);
nor UO_169 (O_169,N_19618,N_18981);
nand UO_170 (O_170,N_17930,N_19114);
xor UO_171 (O_171,N_16201,N_18678);
or UO_172 (O_172,N_17681,N_19366);
nor UO_173 (O_173,N_17179,N_18136);
nor UO_174 (O_174,N_18993,N_19185);
xnor UO_175 (O_175,N_19065,N_19709);
xor UO_176 (O_176,N_16162,N_18530);
xor UO_177 (O_177,N_18425,N_16959);
and UO_178 (O_178,N_16957,N_16094);
or UO_179 (O_179,N_18201,N_19501);
and UO_180 (O_180,N_17770,N_19245);
or UO_181 (O_181,N_16326,N_18749);
or UO_182 (O_182,N_16874,N_16100);
nand UO_183 (O_183,N_16255,N_19302);
nand UO_184 (O_184,N_19242,N_18843);
nor UO_185 (O_185,N_19391,N_19991);
and UO_186 (O_186,N_17311,N_17012);
nor UO_187 (O_187,N_18856,N_17364);
and UO_188 (O_188,N_19095,N_18305);
nor UO_189 (O_189,N_16123,N_16566);
nor UO_190 (O_190,N_16259,N_19434);
nor UO_191 (O_191,N_17131,N_17603);
and UO_192 (O_192,N_19941,N_19122);
and UO_193 (O_193,N_16544,N_16121);
xnor UO_194 (O_194,N_16948,N_18604);
or UO_195 (O_195,N_18184,N_17965);
nand UO_196 (O_196,N_16865,N_19656);
and UO_197 (O_197,N_19676,N_16320);
nand UO_198 (O_198,N_19351,N_17816);
or UO_199 (O_199,N_17753,N_19539);
xor UO_200 (O_200,N_19113,N_18727);
nand UO_201 (O_201,N_19172,N_17298);
xor UO_202 (O_202,N_17892,N_18239);
and UO_203 (O_203,N_16532,N_16808);
nand UO_204 (O_204,N_18971,N_16530);
xor UO_205 (O_205,N_18495,N_19677);
and UO_206 (O_206,N_16088,N_17917);
xor UO_207 (O_207,N_19293,N_16766);
and UO_208 (O_208,N_16779,N_16059);
nand UO_209 (O_209,N_18876,N_16394);
and UO_210 (O_210,N_19097,N_16938);
and UO_211 (O_211,N_17941,N_16991);
and UO_212 (O_212,N_16429,N_18966);
and UO_213 (O_213,N_19096,N_19102);
xnor UO_214 (O_214,N_18003,N_18629);
nor UO_215 (O_215,N_19023,N_17445);
nor UO_216 (O_216,N_17190,N_18186);
and UO_217 (O_217,N_17506,N_16265);
xor UO_218 (O_218,N_19877,N_18857);
nor UO_219 (O_219,N_19862,N_16106);
or UO_220 (O_220,N_18433,N_16185);
and UO_221 (O_221,N_17644,N_18045);
nand UO_222 (O_222,N_18814,N_19094);
or UO_223 (O_223,N_17745,N_16992);
and UO_224 (O_224,N_19966,N_18406);
nand UO_225 (O_225,N_16391,N_19768);
xnor UO_226 (O_226,N_16748,N_17957);
xor UO_227 (O_227,N_17215,N_19449);
and UO_228 (O_228,N_17490,N_18279);
or UO_229 (O_229,N_17527,N_18855);
nor UO_230 (O_230,N_19890,N_17538);
nand UO_231 (O_231,N_19284,N_18670);
or UO_232 (O_232,N_18146,N_19047);
xor UO_233 (O_233,N_16200,N_19541);
nor UO_234 (O_234,N_19171,N_17494);
and UO_235 (O_235,N_19492,N_19068);
and UO_236 (O_236,N_16932,N_17664);
nor UO_237 (O_237,N_17827,N_19568);
nand UO_238 (O_238,N_16414,N_17294);
or UO_239 (O_239,N_17358,N_16334);
and UO_240 (O_240,N_16346,N_18887);
nand UO_241 (O_241,N_16619,N_16966);
and UO_242 (O_242,N_16778,N_17559);
xor UO_243 (O_243,N_16858,N_16849);
xor UO_244 (O_244,N_19153,N_19367);
and UO_245 (O_245,N_19152,N_18863);
nor UO_246 (O_246,N_17028,N_17991);
xnor UO_247 (O_247,N_17518,N_19116);
and UO_248 (O_248,N_18565,N_16289);
xnor UO_249 (O_249,N_18572,N_18633);
nor UO_250 (O_250,N_16662,N_19923);
or UO_251 (O_251,N_16924,N_19075);
and UO_252 (O_252,N_16117,N_19815);
or UO_253 (O_253,N_17593,N_16230);
nand UO_254 (O_254,N_16582,N_18986);
xnor UO_255 (O_255,N_16733,N_16499);
nor UO_256 (O_256,N_19515,N_19926);
nand UO_257 (O_257,N_16086,N_16968);
xnor UO_258 (O_258,N_18954,N_19357);
nor UO_259 (O_259,N_16588,N_16338);
nor UO_260 (O_260,N_16537,N_17069);
nand UO_261 (O_261,N_18810,N_19791);
xor UO_262 (O_262,N_16160,N_18286);
nand UO_263 (O_263,N_16677,N_17376);
xnor UO_264 (O_264,N_19355,N_18919);
nand UO_265 (O_265,N_16408,N_19108);
xnor UO_266 (O_266,N_16672,N_17189);
xor UO_267 (O_267,N_18647,N_19813);
or UO_268 (O_268,N_18683,N_18909);
and UO_269 (O_269,N_18180,N_16950);
or UO_270 (O_270,N_16030,N_17132);
xor UO_271 (O_271,N_16169,N_16776);
or UO_272 (O_272,N_17500,N_18413);
nand UO_273 (O_273,N_18515,N_18125);
nor UO_274 (O_274,N_19314,N_19826);
nand UO_275 (O_275,N_17509,N_19058);
and UO_276 (O_276,N_17249,N_17121);
xor UO_277 (O_277,N_17740,N_16863);
or UO_278 (O_278,N_17555,N_18902);
nand UO_279 (O_279,N_18124,N_19869);
or UO_280 (O_280,N_19856,N_19405);
nor UO_281 (O_281,N_17195,N_19004);
nor UO_282 (O_282,N_17379,N_16983);
nand UO_283 (O_283,N_17620,N_17803);
xor UO_284 (O_284,N_16813,N_18240);
and UO_285 (O_285,N_17949,N_19457);
xnor UO_286 (O_286,N_17980,N_18024);
nand UO_287 (O_287,N_17432,N_16635);
nand UO_288 (O_288,N_17255,N_16487);
nand UO_289 (O_289,N_16236,N_16075);
nand UO_290 (O_290,N_18736,N_17910);
nand UO_291 (O_291,N_16228,N_19666);
xnor UO_292 (O_292,N_16302,N_16099);
xnor UO_293 (O_293,N_18432,N_16962);
nor UO_294 (O_294,N_17116,N_16908);
xnor UO_295 (O_295,N_19767,N_17669);
or UO_296 (O_296,N_16152,N_17489);
and UO_297 (O_297,N_19358,N_19615);
and UO_298 (O_298,N_19505,N_18685);
xor UO_299 (O_299,N_17626,N_18521);
nand UO_300 (O_300,N_16238,N_16612);
nand UO_301 (O_301,N_17365,N_17808);
or UO_302 (O_302,N_17779,N_16015);
xor UO_303 (O_303,N_19894,N_17272);
nand UO_304 (O_304,N_19650,N_19876);
nand UO_305 (O_305,N_18336,N_18285);
nor UO_306 (O_306,N_18951,N_16914);
and UO_307 (O_307,N_18637,N_19530);
and UO_308 (O_308,N_16428,N_19617);
nand UO_309 (O_309,N_16988,N_16835);
nand UO_310 (O_310,N_17606,N_17429);
nor UO_311 (O_311,N_16697,N_18363);
nand UO_312 (O_312,N_17108,N_16191);
xor UO_313 (O_313,N_19784,N_17336);
nand UO_314 (O_314,N_16489,N_19962);
and UO_315 (O_315,N_18101,N_19646);
xor UO_316 (O_316,N_17233,N_17912);
nor UO_317 (O_317,N_17651,N_19957);
and UO_318 (O_318,N_16769,N_19427);
nand UO_319 (O_319,N_19817,N_19001);
nor UO_320 (O_320,N_19164,N_16424);
and UO_321 (O_321,N_18595,N_19563);
xnor UO_322 (O_322,N_19401,N_18628);
or UO_323 (O_323,N_16159,N_16239);
xor UO_324 (O_324,N_19318,N_18546);
and UO_325 (O_325,N_19269,N_17911);
xor UO_326 (O_326,N_17537,N_19517);
and UO_327 (O_327,N_19010,N_17598);
and UO_328 (O_328,N_16746,N_18332);
and UO_329 (O_329,N_16797,N_17252);
nand UO_330 (O_330,N_16919,N_17824);
or UO_331 (O_331,N_17788,N_17475);
xnor UO_332 (O_332,N_19345,N_17383);
xnor UO_333 (O_333,N_17374,N_16945);
or UO_334 (O_334,N_18569,N_16332);
or UO_335 (O_335,N_17051,N_17777);
nor UO_336 (O_336,N_16585,N_18331);
nand UO_337 (O_337,N_18081,N_17258);
nor UO_338 (O_338,N_19661,N_18131);
or UO_339 (O_339,N_19073,N_17755);
xor UO_340 (O_340,N_17579,N_17043);
nand UO_341 (O_341,N_19041,N_17405);
xnor UO_342 (O_342,N_17672,N_18815);
or UO_343 (O_343,N_18196,N_17142);
nand UO_344 (O_344,N_19230,N_16350);
xnor UO_345 (O_345,N_16433,N_19796);
nor UO_346 (O_346,N_17953,N_18965);
and UO_347 (O_347,N_18952,N_17950);
nand UO_348 (O_348,N_19087,N_19907);
nor UO_349 (O_349,N_18946,N_19208);
nand UO_350 (O_350,N_19728,N_19867);
xor UO_351 (O_351,N_18947,N_16976);
and UO_352 (O_352,N_18330,N_18310);
xnor UO_353 (O_353,N_16150,N_17804);
xnor UO_354 (O_354,N_16400,N_17835);
or UO_355 (O_355,N_17278,N_18104);
nor UO_356 (O_356,N_16523,N_18593);
nor UO_357 (O_357,N_19175,N_17561);
xnor UO_358 (O_358,N_16122,N_17531);
nor UO_359 (O_359,N_18907,N_17751);
nand UO_360 (O_360,N_18702,N_16067);
nor UO_361 (O_361,N_18931,N_16944);
nand UO_362 (O_362,N_19454,N_16074);
nor UO_363 (O_363,N_18525,N_17660);
nand UO_364 (O_364,N_19018,N_16032);
xor UO_365 (O_365,N_19084,N_17165);
nand UO_366 (O_366,N_16385,N_16574);
or UO_367 (O_367,N_16213,N_18304);
or UO_368 (O_368,N_16581,N_19969);
xor UO_369 (O_369,N_17585,N_17833);
nor UO_370 (O_370,N_17474,N_16843);
nor UO_371 (O_371,N_18282,N_18973);
nor UO_372 (O_372,N_18010,N_19037);
nor UO_373 (O_373,N_16799,N_17674);
and UO_374 (O_374,N_16354,N_17945);
nand UO_375 (O_375,N_17164,N_17304);
nand UO_376 (O_376,N_18047,N_17420);
nand UO_377 (O_377,N_18044,N_17217);
or UO_378 (O_378,N_17858,N_19537);
or UO_379 (O_379,N_19573,N_17864);
or UO_380 (O_380,N_17934,N_19553);
nand UO_381 (O_381,N_16531,N_17662);
nand UO_382 (O_382,N_17642,N_17380);
and UO_383 (O_383,N_17079,N_18106);
or UO_384 (O_384,N_17629,N_19370);
xor UO_385 (O_385,N_19811,N_17351);
and UO_386 (O_386,N_19627,N_19158);
and UO_387 (O_387,N_18256,N_17315);
or UO_388 (O_388,N_19081,N_16457);
nand UO_389 (O_389,N_18687,N_16687);
or UO_390 (O_390,N_19375,N_18020);
nand UO_391 (O_391,N_19868,N_19659);
nand UO_392 (O_392,N_18155,N_19903);
or UO_393 (O_393,N_17138,N_16016);
and UO_394 (O_394,N_17451,N_17821);
nand UO_395 (O_395,N_16351,N_17316);
nor UO_396 (O_396,N_19836,N_18894);
xnor UO_397 (O_397,N_17234,N_19069);
nand UO_398 (O_398,N_18224,N_18174);
nand UO_399 (O_399,N_18387,N_17488);
and UO_400 (O_400,N_18189,N_16096);
and UO_401 (O_401,N_18803,N_19942);
xnor UO_402 (O_402,N_19256,N_19110);
or UO_403 (O_403,N_16456,N_17350);
nand UO_404 (O_404,N_17594,N_16058);
xnor UO_405 (O_405,N_18686,N_16753);
or UO_406 (O_406,N_19368,N_17963);
nor UO_407 (O_407,N_16707,N_18837);
nor UO_408 (O_408,N_16008,N_18471);
and UO_409 (O_409,N_17180,N_18964);
or UO_410 (O_410,N_17267,N_18041);
xnor UO_411 (O_411,N_16506,N_18524);
xnor UO_412 (O_412,N_17846,N_16089);
xnor UO_413 (O_413,N_18605,N_19022);
nor UO_414 (O_414,N_17246,N_18297);
xnor UO_415 (O_415,N_18776,N_17560);
or UO_416 (O_416,N_19693,N_18556);
and UO_417 (O_417,N_17446,N_17903);
xnor UO_418 (O_418,N_16374,N_18322);
nor UO_419 (O_419,N_19105,N_17162);
nand UO_420 (O_420,N_18200,N_18164);
nand UO_421 (O_421,N_19042,N_18488);
nor UO_422 (O_422,N_19897,N_17140);
nand UO_423 (O_423,N_19461,N_17501);
nand UO_424 (O_424,N_19495,N_19300);
and UO_425 (O_425,N_19762,N_19556);
nor UO_426 (O_426,N_17533,N_19481);
or UO_427 (O_427,N_16494,N_17746);
or UO_428 (O_428,N_16469,N_16832);
nor UO_429 (O_429,N_17842,N_19283);
and UO_430 (O_430,N_19755,N_17005);
nand UO_431 (O_431,N_19985,N_17955);
xnor UO_432 (O_432,N_18329,N_16744);
and UO_433 (O_433,N_16904,N_18542);
or UO_434 (O_434,N_17450,N_19115);
nand UO_435 (O_435,N_17307,N_17806);
xor UO_436 (O_436,N_18065,N_18376);
nand UO_437 (O_437,N_16987,N_16941);
nand UO_438 (O_438,N_19652,N_17113);
nand UO_439 (O_439,N_16997,N_17836);
and UO_440 (O_440,N_19795,N_17654);
or UO_441 (O_441,N_17168,N_19234);
and UO_442 (O_442,N_18232,N_17198);
nand UO_443 (O_443,N_16246,N_17922);
xnor UO_444 (O_444,N_18975,N_16994);
or UO_445 (O_445,N_19490,N_18316);
nor UO_446 (O_446,N_18482,N_17697);
and UO_447 (O_447,N_17573,N_18935);
xnor UO_448 (O_448,N_16247,N_16304);
xnor UO_449 (O_449,N_18624,N_17033);
and UO_450 (O_450,N_18753,N_17981);
nand UO_451 (O_451,N_16027,N_16130);
or UO_452 (O_452,N_17541,N_16599);
nand UO_453 (O_453,N_19612,N_17631);
xor UO_454 (O_454,N_17394,N_16807);
and UO_455 (O_455,N_18038,N_19819);
nor UO_456 (O_456,N_16528,N_18416);
nor UO_457 (O_457,N_16551,N_18910);
nor UO_458 (O_458,N_19289,N_17898);
nand UO_459 (O_459,N_19346,N_19267);
and UO_460 (O_460,N_18431,N_18342);
nand UO_461 (O_461,N_16192,N_16315);
nand UO_462 (O_462,N_16051,N_18484);
nor UO_463 (O_463,N_16846,N_18568);
xnor UO_464 (O_464,N_18289,N_19841);
nor UO_465 (O_465,N_18859,N_19040);
nand UO_466 (O_466,N_16855,N_17584);
and UO_467 (O_467,N_19719,N_16727);
nand UO_468 (O_468,N_19450,N_19686);
nand UO_469 (O_469,N_17270,N_16490);
and UO_470 (O_470,N_19438,N_16847);
nand UO_471 (O_471,N_18267,N_16686);
xnor UO_472 (O_472,N_16708,N_16844);
nor UO_473 (O_473,N_16892,N_16220);
xor UO_474 (O_474,N_18819,N_18867);
and UO_475 (O_475,N_18582,N_16597);
nor UO_476 (O_476,N_16867,N_18693);
or UO_477 (O_477,N_16440,N_19548);
nand UO_478 (O_478,N_19790,N_16911);
and UO_479 (O_479,N_16203,N_18323);
xor UO_480 (O_480,N_16584,N_19717);
nand UO_481 (O_481,N_16986,N_19905);
nand UO_482 (O_482,N_19732,N_16057);
xnor UO_483 (O_483,N_19244,N_17988);
nor UO_484 (O_484,N_16163,N_19141);
and UO_485 (O_485,N_17952,N_16436);
xnor UO_486 (O_486,N_18209,N_18040);
xor UO_487 (O_487,N_18563,N_18409);
nand UO_488 (O_488,N_18309,N_18747);
and UO_489 (O_489,N_16250,N_18745);
or UO_490 (O_490,N_17359,N_18149);
or UO_491 (O_491,N_19130,N_18713);
nor UO_492 (O_492,N_19882,N_17325);
or UO_493 (O_493,N_19581,N_16411);
xnor UO_494 (O_494,N_17763,N_17139);
and UO_495 (O_495,N_18735,N_19812);
xor UO_496 (O_496,N_19316,N_18025);
xnor UO_497 (O_497,N_17625,N_19625);
nor UO_498 (O_498,N_19007,N_18333);
nand UO_499 (O_499,N_18886,N_19015);
nor UO_500 (O_500,N_18562,N_19820);
nor UO_501 (O_501,N_16337,N_16970);
xor UO_502 (O_502,N_18625,N_19547);
and UO_503 (O_503,N_19685,N_18940);
nand UO_504 (O_504,N_18117,N_19270);
or UO_505 (O_505,N_17175,N_16549);
nand UO_506 (O_506,N_19468,N_19264);
nand UO_507 (O_507,N_18982,N_18494);
nand UO_508 (O_508,N_18222,N_17010);
nand UO_509 (O_509,N_16511,N_18429);
nand UO_510 (O_510,N_17129,N_18835);
or UO_511 (O_511,N_18630,N_17926);
nor UO_512 (O_512,N_17360,N_17613);
and UO_513 (O_513,N_17461,N_17347);
and UO_514 (O_514,N_16380,N_17464);
or UO_515 (O_515,N_18704,N_18699);
nor UO_516 (O_516,N_19742,N_19385);
xnor UO_517 (O_517,N_16056,N_16071);
and UO_518 (O_518,N_18248,N_19880);
nor UO_519 (O_519,N_18328,N_16331);
nor UO_520 (O_520,N_18300,N_19967);
or UO_521 (O_521,N_19525,N_19861);
and UO_522 (O_522,N_17466,N_17434);
nand UO_523 (O_523,N_18138,N_18707);
nor UO_524 (O_524,N_17595,N_16368);
and UO_525 (O_525,N_19067,N_19599);
xor UO_526 (O_526,N_16366,N_16996);
xor UO_527 (O_527,N_18371,N_16283);
and UO_528 (O_528,N_19399,N_19340);
nor UO_529 (O_529,N_16044,N_18436);
nor UO_530 (O_530,N_19570,N_17604);
nor UO_531 (O_531,N_17586,N_16404);
nor UO_532 (O_532,N_19915,N_17802);
nand UO_533 (O_533,N_16298,N_17924);
xor UO_534 (O_534,N_19843,N_17760);
nor UO_535 (O_535,N_18696,N_16470);
nor UO_536 (O_536,N_17236,N_19431);
or UO_537 (O_537,N_19045,N_16774);
nor UO_538 (O_538,N_18933,N_16652);
or UO_539 (O_539,N_19632,N_16809);
xor UO_540 (O_540,N_17194,N_16960);
or UO_541 (O_541,N_17157,N_18172);
xnor UO_542 (O_542,N_18895,N_17732);
nor UO_543 (O_543,N_16022,N_16198);
nor UO_544 (O_544,N_16745,N_18538);
and UO_545 (O_545,N_16647,N_19031);
or UO_546 (O_546,N_18591,N_16830);
xnor UO_547 (O_547,N_17805,N_19420);
nand UO_548 (O_548,N_19280,N_18058);
xnor UO_549 (O_549,N_17900,N_16093);
nand UO_550 (O_550,N_17378,N_19129);
xor UO_551 (O_551,N_16402,N_19460);
nand UO_552 (O_552,N_17507,N_17112);
xnor UO_553 (O_553,N_18864,N_18726);
nor UO_554 (O_554,N_18541,N_17729);
nand UO_555 (O_555,N_16762,N_18950);
nand UO_556 (O_556,N_16611,N_18207);
nand UO_557 (O_557,N_16111,N_19716);
nor UO_558 (O_558,N_17915,N_17820);
and UO_559 (O_559,N_18681,N_19008);
nor UO_560 (O_560,N_17575,N_18914);
and UO_561 (O_561,N_18543,N_19943);
or UO_562 (O_562,N_18778,N_16617);
nor UO_563 (O_563,N_18448,N_16949);
nand UO_564 (O_564,N_18299,N_17271);
nand UO_565 (O_565,N_19298,N_16000);
and UO_566 (O_566,N_18173,N_19860);
or UO_567 (O_567,N_18119,N_19463);
nor UO_568 (O_568,N_18344,N_18551);
xnor UO_569 (O_569,N_16055,N_19921);
nand UO_570 (O_570,N_17210,N_17863);
nand UO_571 (O_571,N_17040,N_17929);
nor UO_572 (O_572,N_18665,N_17693);
and UO_573 (O_573,N_16137,N_17630);
nor UO_574 (O_574,N_19692,N_17747);
or UO_575 (O_575,N_18664,N_16609);
and UO_576 (O_576,N_18401,N_16869);
or UO_577 (O_577,N_16232,N_17412);
xor UO_578 (O_578,N_19012,N_16365);
nor UO_579 (O_579,N_17721,N_18706);
nand UO_580 (O_580,N_19664,N_16703);
or UO_581 (O_581,N_18249,N_17150);
and UO_582 (O_582,N_17719,N_18638);
nor UO_583 (O_583,N_18160,N_16935);
nor UO_584 (O_584,N_18134,N_17279);
or UO_585 (O_585,N_19809,N_16743);
or UO_586 (O_586,N_19080,N_17689);
nor UO_587 (O_587,N_19464,N_16110);
nor UO_588 (O_588,N_16272,N_17022);
and UO_589 (O_589,N_17877,N_17971);
xnor UO_590 (O_590,N_17341,N_16426);
and UO_591 (O_591,N_16660,N_17744);
xnor UO_592 (O_592,N_19124,N_19873);
nand UO_593 (O_593,N_19718,N_17716);
nand UO_594 (O_594,N_17332,N_17172);
and UO_595 (O_595,N_19465,N_17483);
xor UO_596 (O_596,N_17510,N_18755);
nand UO_597 (O_597,N_16318,N_17639);
or UO_598 (O_598,N_19747,N_18846);
or UO_599 (O_599,N_18660,N_19326);
or UO_600 (O_600,N_16831,N_19177);
xnor UO_601 (O_601,N_16508,N_17056);
or UO_602 (O_602,N_17828,N_18705);
or UO_603 (O_603,N_17013,N_16208);
and UO_604 (O_604,N_16852,N_19064);
nand UO_605 (O_605,N_16918,N_16951);
nand UO_606 (O_606,N_17801,N_19690);
nand UO_607 (O_607,N_17727,N_19863);
nand UO_608 (O_608,N_16622,N_16507);
nor UO_609 (O_609,N_19272,N_16202);
nor UO_610 (O_610,N_19783,N_16965);
or UO_611 (O_611,N_16702,N_18728);
and UO_612 (O_612,N_18836,N_17522);
xnor UO_613 (O_613,N_17547,N_19341);
or UO_614 (O_614,N_19605,N_16425);
nor UO_615 (O_615,N_16593,N_18468);
xnor UO_616 (O_616,N_16468,N_18352);
nor UO_617 (O_617,N_17385,N_16692);
nand UO_618 (O_618,N_17076,N_19965);
or UO_619 (O_619,N_16422,N_19053);
or UO_620 (O_620,N_17503,N_17568);
or UO_621 (O_621,N_16041,N_18743);
nor UO_622 (O_622,N_17468,N_17460);
or UO_623 (O_623,N_18643,N_19844);
xor UO_624 (O_624,N_18979,N_16534);
or UO_625 (O_625,N_19428,N_19477);
nor UO_626 (O_626,N_17030,N_18567);
xor UO_627 (O_627,N_18888,N_16445);
and UO_628 (O_628,N_16126,N_16109);
nand UO_629 (O_629,N_17589,N_19754);
and UO_630 (O_630,N_19778,N_16262);
xor UO_631 (O_631,N_17617,N_18989);
and UO_632 (O_632,N_19315,N_16329);
or UO_633 (O_633,N_19059,N_18571);
and UO_634 (O_634,N_18767,N_18631);
xnor UO_635 (O_635,N_18465,N_17421);
and UO_636 (O_636,N_18682,N_16925);
xnor UO_637 (O_637,N_16413,N_19486);
nor UO_638 (O_638,N_16484,N_18251);
nor UO_639 (O_639,N_18817,N_16518);
nand UO_640 (O_640,N_19723,N_19975);
or UO_641 (O_641,N_16211,N_18012);
nor UO_642 (O_642,N_18768,N_16688);
and UO_643 (O_643,N_16801,N_18023);
nor UO_644 (O_644,N_16340,N_17548);
nor UO_645 (O_645,N_19898,N_18828);
nor UO_646 (O_646,N_18862,N_18573);
or UO_647 (O_647,N_17001,N_16166);
nand UO_648 (O_648,N_17003,N_17794);
nand UO_649 (O_649,N_19651,N_19196);
xnor UO_650 (O_650,N_18009,N_19142);
nor UO_651 (O_651,N_18800,N_19236);
nor UO_652 (O_652,N_19494,N_16943);
nor UO_653 (O_653,N_16971,N_19061);
or UO_654 (O_654,N_18636,N_18386);
nor UO_655 (O_655,N_19214,N_17713);
and UO_656 (O_656,N_17273,N_16290);
xor UO_657 (O_657,N_16336,N_19774);
and UO_658 (O_658,N_19237,N_18620);
xor UO_659 (O_659,N_17847,N_17170);
nor UO_660 (O_660,N_17853,N_19002);
or UO_661 (O_661,N_18396,N_19769);
or UO_662 (O_662,N_18640,N_18614);
and UO_663 (O_663,N_17484,N_18349);
and UO_664 (O_664,N_18446,N_18437);
xnor UO_665 (O_665,N_17070,N_18868);
xor UO_666 (O_666,N_16509,N_19441);
nor UO_667 (O_667,N_17435,N_18419);
nor UO_668 (O_668,N_19295,N_18792);
nor UO_669 (O_669,N_16389,N_19090);
nand UO_670 (O_670,N_18759,N_19902);
and UO_671 (O_671,N_19136,N_18114);
or UO_672 (O_672,N_19429,N_17878);
and UO_673 (O_673,N_18698,N_17021);
nor UO_674 (O_674,N_19235,N_17987);
and UO_675 (O_675,N_16267,N_17206);
or UO_676 (O_676,N_19889,N_16767);
and UO_677 (O_677,N_18765,N_19528);
nor UO_678 (O_678,N_19246,N_18063);
nand UO_679 (O_679,N_19776,N_19066);
or UO_680 (O_680,N_16734,N_18430);
nand UO_681 (O_681,N_16291,N_16127);
and UO_682 (O_682,N_18892,N_18708);
nand UO_683 (O_683,N_18340,N_19336);
and UO_684 (O_684,N_16442,N_18754);
and UO_685 (O_685,N_16438,N_18719);
and UO_686 (O_686,N_17807,N_18008);
xnor UO_687 (O_687,N_17994,N_17624);
xnor UO_688 (O_688,N_19402,N_17486);
or UO_689 (O_689,N_17829,N_16164);
nand UO_690 (O_690,N_17302,N_16643);
nand UO_691 (O_691,N_18477,N_17571);
xnor UO_692 (O_692,N_18626,N_18650);
and UO_693 (O_693,N_18639,N_17967);
nand UO_694 (O_694,N_17718,N_17809);
and UO_695 (O_695,N_19038,N_18715);
xor UO_696 (O_696,N_16177,N_17995);
or UO_697 (O_697,N_18746,N_18337);
xnor UO_698 (O_698,N_19071,N_18480);
or UO_699 (O_699,N_19184,N_17838);
or UO_700 (O_700,N_18958,N_18794);
and UO_701 (O_701,N_16501,N_19265);
nor UO_702 (O_702,N_16705,N_17019);
nor UO_703 (O_703,N_16513,N_18193);
or UO_704 (O_704,N_18262,N_17576);
and UO_705 (O_705,N_16307,N_17597);
nor UO_706 (O_706,N_16517,N_19466);
or UO_707 (O_707,N_17224,N_17783);
nand UO_708 (O_708,N_18899,N_19745);
nand UO_709 (O_709,N_16760,N_19197);
or UO_710 (O_710,N_16128,N_16077);
or UO_711 (O_711,N_16548,N_17024);
xor UO_712 (O_712,N_16765,N_18073);
or UO_713 (O_713,N_19091,N_16666);
nand UO_714 (O_714,N_17044,N_19440);
nand UO_715 (O_715,N_19734,N_18335);
and UO_716 (O_716,N_19533,N_19700);
nand UO_717 (O_717,N_16060,N_19883);
nor UO_718 (O_718,N_17239,N_19211);
xnor UO_719 (O_719,N_18393,N_17319);
nand UO_720 (O_720,N_17938,N_19984);
xnor UO_721 (O_721,N_18086,N_18917);
and UO_722 (O_722,N_16479,N_16757);
xor UO_723 (O_723,N_19304,N_17855);
nand UO_724 (O_724,N_19822,N_19487);
or UO_725 (O_725,N_19583,N_18466);
xor UO_726 (O_726,N_18564,N_19126);
and UO_727 (O_727,N_18143,N_16184);
or UO_728 (O_728,N_16978,N_17199);
nand UO_729 (O_729,N_18536,N_18381);
xnor UO_730 (O_730,N_18121,N_17293);
nand UO_731 (O_731,N_17738,N_18402);
and UO_732 (O_732,N_16043,N_18182);
nand UO_733 (O_733,N_18303,N_16136);
or UO_734 (O_734,N_18513,N_17313);
nor UO_735 (O_735,N_19810,N_19593);
xor UO_736 (O_736,N_18382,N_19892);
xor UO_737 (O_737,N_18062,N_18878);
and UO_738 (O_738,N_19833,N_18635);
xnor UO_739 (O_739,N_19194,N_16661);
nand UO_740 (O_740,N_17914,N_19891);
xor UO_741 (O_741,N_18539,N_18418);
or UO_742 (O_742,N_19027,N_19444);
and UO_743 (O_743,N_19866,N_18588);
nor UO_744 (O_744,N_17439,N_18355);
xor UO_745 (O_745,N_18254,N_19424);
nand UO_746 (O_746,N_17482,N_17391);
or UO_747 (O_747,N_17978,N_16591);
nand UO_748 (O_748,N_19488,N_18766);
xor UO_749 (O_749,N_18076,N_17283);
nand UO_750 (O_750,N_19855,N_19123);
or UO_751 (O_751,N_17227,N_16274);
xnor UO_752 (O_752,N_18597,N_18881);
and UO_753 (O_753,N_16142,N_16349);
or UO_754 (O_754,N_19789,N_18646);
and UO_755 (O_755,N_16386,N_19614);
xor UO_756 (O_756,N_16118,N_19162);
xor UO_757 (O_757,N_19117,N_18723);
and UO_758 (O_758,N_17523,N_19945);
xor UO_759 (O_759,N_18325,N_17904);
nand UO_760 (O_760,N_16460,N_16396);
nor UO_761 (O_761,N_16726,N_19174);
xnor UO_762 (O_762,N_19644,N_17377);
xnor UO_763 (O_763,N_19696,N_17769);
and UO_764 (O_764,N_19221,N_17993);
nand UO_765 (O_765,N_16023,N_17250);
nand UO_766 (O_766,N_19940,N_17430);
xor UO_767 (O_767,N_19392,N_16370);
nor UO_768 (O_768,N_18153,N_16025);
or UO_769 (O_769,N_16263,N_18061);
nor UO_770 (O_770,N_17996,N_19056);
or UO_771 (O_771,N_18609,N_18223);
or UO_772 (O_772,N_19220,N_17705);
or UO_773 (O_773,N_18374,N_19509);
or UO_774 (O_774,N_16675,N_18351);
and UO_775 (O_775,N_16300,N_19238);
and UO_776 (O_776,N_17811,N_18443);
and UO_777 (O_777,N_17059,N_16875);
nor UO_778 (O_778,N_16942,N_18213);
nand UO_779 (O_779,N_18663,N_18760);
nor UO_780 (O_780,N_19452,N_18007);
nor UO_781 (O_781,N_16592,N_19217);
nand UO_782 (O_782,N_18953,N_17975);
or UO_783 (O_783,N_17153,N_17025);
nand UO_784 (O_784,N_17321,N_19821);
nand UO_785 (O_785,N_17848,N_16552);
xnor UO_786 (O_786,N_18272,N_16268);
or UO_787 (O_787,N_17235,N_16223);
and UO_788 (O_788,N_18566,N_17124);
or UO_789 (O_789,N_17759,N_16606);
nor UO_790 (O_790,N_19695,N_19950);
and UO_791 (O_791,N_18897,N_17089);
and UO_792 (O_792,N_19920,N_19752);
or UO_793 (O_793,N_16270,N_18645);
nor UO_794 (O_794,N_16859,N_19137);
xor UO_795 (O_795,N_19078,N_19433);
and UO_796 (O_796,N_18851,N_19497);
xnor UO_797 (O_797,N_17055,N_18997);
xnor UO_798 (O_798,N_16804,N_18927);
nand UO_799 (O_799,N_19832,N_18270);
and UO_800 (O_800,N_19133,N_17031);
nand UO_801 (O_801,N_19846,N_16048);
or UO_802 (O_802,N_19055,N_18098);
or UO_803 (O_803,N_16073,N_17441);
nor UO_804 (O_804,N_17145,N_17086);
xor UO_805 (O_805,N_18424,N_17887);
and UO_806 (O_806,N_19377,N_18570);
or UO_807 (O_807,N_16153,N_17229);
nand UO_808 (O_808,N_18956,N_16480);
xnor UO_809 (O_809,N_16999,N_17411);
nand UO_810 (O_810,N_19911,N_17823);
nor UO_811 (O_811,N_19485,N_17621);
nand UO_812 (O_812,N_19000,N_17128);
xnor UO_813 (O_813,N_18102,N_17075);
nor UO_814 (O_814,N_18697,N_19572);
nand UO_815 (O_815,N_17885,N_17513);
and UO_816 (O_816,N_18055,N_19191);
nand UO_817 (O_817,N_18540,N_17372);
or UO_818 (O_818,N_16158,N_18816);
xnor UO_819 (O_819,N_17819,N_17186);
and UO_820 (O_820,N_16277,N_16963);
xnor UO_821 (O_821,N_16180,N_16335);
and UO_822 (O_822,N_19190,N_16634);
and UO_823 (O_823,N_19030,N_18490);
nand UO_824 (O_824,N_16222,N_17009);
xnor UO_825 (O_825,N_19608,N_19613);
nor UO_826 (O_826,N_17986,N_17638);
nand UO_827 (O_827,N_18666,N_17375);
xnor UO_828 (O_828,N_19291,N_19785);
and UO_829 (O_829,N_17731,N_18202);
nand UO_830 (O_830,N_18577,N_16435);
and UO_831 (O_831,N_19474,N_16157);
or UO_832 (O_832,N_19390,N_17976);
and UO_833 (O_833,N_19549,N_16282);
xnor UO_834 (O_834,N_17073,N_17454);
or UO_835 (O_835,N_16434,N_19702);
or UO_836 (O_836,N_17326,N_19688);
xnor UO_837 (O_837,N_17016,N_18912);
nor UO_838 (O_838,N_19623,N_16819);
or UO_839 (O_839,N_19321,N_19011);
nand UO_840 (O_840,N_17406,N_17134);
or UO_841 (O_841,N_18421,N_17141);
xnor UO_842 (O_842,N_19672,N_16231);
or UO_843 (O_843,N_16610,N_19986);
or UO_844 (O_844,N_17403,N_16148);
nor UO_845 (O_845,N_16824,N_19727);
xnor UO_846 (O_846,N_16311,N_16639);
nand UO_847 (O_847,N_18087,N_18291);
nor UO_848 (O_848,N_17353,N_17707);
xor UO_849 (O_849,N_18756,N_18343);
or UO_850 (O_850,N_19729,N_16718);
nor UO_851 (O_851,N_19683,N_18891);
nor UO_852 (O_852,N_16278,N_18311);
or UO_853 (O_853,N_16197,N_19766);
nand UO_854 (O_854,N_17477,N_16464);
xor UO_855 (O_855,N_19409,N_16174);
nand UO_856 (O_856,N_17363,N_16013);
or UO_857 (O_857,N_16860,N_16104);
nand UO_858 (O_858,N_19806,N_16958);
or UO_859 (O_859,N_17539,N_16235);
nor UO_860 (O_860,N_18671,N_16827);
nor UO_861 (O_861,N_18720,N_19338);
or UO_862 (O_862,N_18140,N_16078);
nand UO_863 (O_863,N_19679,N_16439);
nor UO_864 (O_864,N_17856,N_19250);
and UO_865 (O_865,N_18592,N_19626);
or UO_866 (O_866,N_16740,N_19179);
xnor UO_867 (O_867,N_19764,N_19206);
nand UO_868 (O_868,N_17045,N_16498);
or UO_869 (O_869,N_17792,N_17956);
or UO_870 (O_870,N_16781,N_17225);
or UO_871 (O_871,N_18084,N_19990);
nand UO_872 (O_872,N_18372,N_16141);
nor UO_873 (O_873,N_17826,N_19388);
and UO_874 (O_874,N_16946,N_19192);
and UO_875 (O_875,N_17558,N_19749);
nor UO_876 (O_876,N_16969,N_19479);
nand UO_877 (O_877,N_16885,N_16777);
xor UO_878 (O_878,N_16782,N_17698);
xnor UO_879 (O_879,N_17262,N_19978);
nand UO_880 (O_880,N_16503,N_19482);
or UO_881 (O_881,N_17151,N_19871);
xnor UO_882 (O_882,N_19426,N_19099);
and UO_883 (O_883,N_16995,N_18428);
or UO_884 (O_884,N_17782,N_16279);
nor UO_885 (O_885,N_16325,N_18955);
or UO_886 (O_886,N_17565,N_16107);
or UO_887 (O_887,N_17428,N_16049);
or UO_888 (O_888,N_19595,N_18779);
nand UO_889 (O_889,N_16024,N_17345);
xnor UO_890 (O_890,N_16216,N_17184);
xnor UO_891 (O_891,N_19266,N_16395);
or UO_892 (O_892,N_17305,N_16710);
xor UO_893 (O_893,N_16533,N_18733);
xnor UO_894 (O_894,N_16732,N_19119);
nor UO_895 (O_895,N_16237,N_17778);
xnor UO_896 (O_896,N_19908,N_19893);
nor UO_897 (O_897,N_19077,N_18266);
xor UO_898 (O_898,N_19958,N_18970);
xor UO_899 (O_899,N_17992,N_17508);
nand UO_900 (O_900,N_18939,N_18247);
xnor UO_901 (O_901,N_19057,N_16066);
nand UO_902 (O_902,N_16085,N_16529);
nand UO_903 (O_903,N_19112,N_16009);
nor UO_904 (O_904,N_18283,N_19363);
or UO_905 (O_905,N_19981,N_17264);
nand UO_906 (O_906,N_19887,N_17203);
or UO_907 (O_907,N_17469,N_18345);
nor UO_908 (O_908,N_16775,N_16155);
or UO_909 (O_909,N_16462,N_18218);
or UO_910 (O_910,N_16314,N_17327);
xnor UO_911 (O_911,N_18258,N_17187);
and UO_912 (O_912,N_16020,N_17202);
or UO_913 (O_913,N_18990,N_17143);
xor UO_914 (O_914,N_18085,N_19937);
nor UO_915 (O_915,N_17608,N_17125);
and UO_916 (O_916,N_19014,N_16909);
and UO_917 (O_917,N_19261,N_17136);
or UO_918 (O_918,N_18644,N_16522);
nand UO_919 (O_919,N_19063,N_19143);
xnor UO_920 (O_920,N_16728,N_17545);
nand UO_921 (O_921,N_17906,N_17958);
or UO_922 (O_922,N_18320,N_17787);
nand UO_923 (O_923,N_18928,N_16179);
nand UO_924 (O_924,N_16485,N_16261);
and UO_925 (O_925,N_19074,N_17999);
and UO_926 (O_926,N_19949,N_17607);
xnor UO_927 (O_927,N_18082,N_19279);
xor UO_928 (O_928,N_17256,N_16172);
and UO_929 (O_929,N_17567,N_16550);
or UO_930 (O_930,N_19313,N_17773);
and UO_931 (O_931,N_19673,N_17291);
xor UO_932 (O_932,N_18548,N_16711);
xnor UO_933 (O_933,N_16288,N_16031);
or UO_934 (O_934,N_19200,N_16837);
xor UO_935 (O_935,N_19665,N_18019);
nand UO_936 (O_936,N_17730,N_17467);
nand UO_937 (O_937,N_17408,N_18099);
nand UO_938 (O_938,N_19360,N_17704);
and UO_939 (O_939,N_19655,N_17743);
nor UO_940 (O_940,N_17018,N_16691);
or UO_941 (O_941,N_16838,N_19854);
nor UO_942 (O_942,N_16398,N_19052);
nand UO_943 (O_943,N_19551,N_17682);
nor UO_944 (O_944,N_16798,N_16562);
nor UO_945 (O_945,N_17916,N_19103);
xor UO_946 (O_946,N_18692,N_18301);
or UO_947 (O_947,N_16251,N_19689);
nor UO_948 (O_948,N_16783,N_19309);
nand UO_949 (O_949,N_16889,N_18520);
or UO_950 (O_950,N_17296,N_19334);
nor UO_951 (O_951,N_17335,N_16817);
xor UO_952 (O_952,N_18067,N_16967);
xnor UO_953 (O_953,N_17318,N_16596);
nand UO_954 (O_954,N_17962,N_19350);
nor UO_955 (O_955,N_19919,N_17741);
xnor UO_956 (O_956,N_17054,N_18516);
xnor UO_957 (O_957,N_18271,N_16629);
nor UO_958 (O_958,N_16496,N_16557);
nand UO_959 (O_959,N_18014,N_17839);
nand UO_960 (O_960,N_16280,N_16210);
nand UO_961 (O_961,N_18890,N_19403);
or UO_962 (O_962,N_16642,N_18763);
nand UO_963 (O_963,N_19181,N_17722);
nor UO_964 (O_964,N_18388,N_19807);
xor UO_965 (O_965,N_19342,N_16249);
nand UO_966 (O_966,N_16638,N_19389);
xor UO_967 (O_967,N_19252,N_18227);
nor UO_968 (O_968,N_17762,N_17207);
and UO_969 (O_969,N_17663,N_16825);
and UO_970 (O_970,N_16853,N_16448);
xor UO_971 (O_971,N_16284,N_17169);
nor UO_972 (O_972,N_19532,N_18263);
nor UO_973 (O_973,N_18877,N_18854);
nor UO_974 (O_974,N_18033,N_17280);
nand UO_975 (O_975,N_19202,N_19048);
nand UO_976 (O_976,N_17881,N_16035);
and UO_977 (O_977,N_17182,N_18415);
nor UO_978 (O_978,N_19249,N_17596);
nor UO_979 (O_979,N_19629,N_17869);
or UO_980 (O_980,N_18811,N_19147);
nor UO_981 (O_981,N_17640,N_18290);
nand UO_982 (O_982,N_16794,N_16952);
xnor UO_983 (O_983,N_17551,N_16316);
nand UO_984 (O_984,N_16937,N_19404);
or UO_985 (O_985,N_17458,N_18170);
nand UO_986 (O_986,N_16356,N_16676);
and UO_987 (O_987,N_17306,N_16930);
or UO_988 (O_988,N_18027,N_16176);
and UO_989 (O_989,N_18809,N_17257);
and UO_990 (O_990,N_18995,N_17504);
nand UO_991 (O_991,N_16119,N_16700);
and UO_992 (O_992,N_19961,N_18949);
nor UO_993 (O_993,N_19382,N_17879);
nor UO_994 (O_994,N_19413,N_16478);
nand UO_995 (O_995,N_18463,N_16173);
nor UO_996 (O_996,N_16193,N_16573);
nor UO_997 (O_997,N_16872,N_17582);
xor UO_998 (O_998,N_17865,N_19183);
or UO_999 (O_999,N_18603,N_18700);
nor UO_1000 (O_1000,N_16054,N_16927);
nand UO_1001 (O_1001,N_19725,N_16444);
nor UO_1002 (O_1002,N_18985,N_17297);
and UO_1003 (O_1003,N_17285,N_19711);
or UO_1004 (O_1004,N_18834,N_16524);
nor UO_1005 (O_1005,N_18555,N_19455);
nor UO_1006 (O_1006,N_18420,N_16387);
xor UO_1007 (O_1007,N_17083,N_18235);
and UO_1008 (O_1008,N_19006,N_19788);
xor UO_1009 (O_1009,N_16880,N_19564);
and UO_1010 (O_1010,N_19268,N_19864);
xor UO_1011 (O_1011,N_19559,N_17591);
xnor UO_1012 (O_1012,N_19135,N_16520);
nand UO_1013 (O_1013,N_18938,N_19332);
or UO_1014 (O_1014,N_17082,N_17696);
or UO_1015 (O_1015,N_18191,N_19442);
nor UO_1016 (O_1016,N_18403,N_19988);
and UO_1017 (O_1017,N_19827,N_16741);
and UO_1018 (O_1018,N_17158,N_18889);
xor UO_1019 (O_1019,N_18011,N_17641);
or UO_1020 (O_1020,N_16899,N_18557);
nor UO_1021 (O_1021,N_18865,N_16327);
xor UO_1022 (O_1022,N_19682,N_19294);
nand UO_1023 (O_1023,N_16876,N_17919);
or UO_1024 (O_1024,N_17231,N_17417);
nand UO_1025 (O_1025,N_18177,N_16323);
and UO_1026 (O_1026,N_16805,N_16678);
nor UO_1027 (O_1027,N_19726,N_18205);
nand UO_1028 (O_1028,N_17799,N_19590);
xnor UO_1029 (O_1029,N_17884,N_18206);
nor UO_1030 (O_1030,N_16598,N_16620);
nor UO_1031 (O_1031,N_18504,N_18994);
and UO_1032 (O_1032,N_18900,N_17678);
xor UO_1033 (O_1033,N_18253,N_18489);
or UO_1034 (O_1034,N_18712,N_18709);
nor UO_1035 (O_1035,N_18195,N_16091);
nand UO_1036 (O_1036,N_19750,N_18972);
and UO_1037 (O_1037,N_16372,N_16881);
xnor UO_1038 (O_1038,N_18587,N_19227);
or UO_1039 (O_1039,N_16771,N_17098);
and UO_1040 (O_1040,N_18366,N_16579);
and UO_1041 (O_1041,N_18051,N_19507);
nor UO_1042 (O_1042,N_18662,N_17392);
nor UO_1043 (O_1043,N_16841,N_18244);
nand UO_1044 (O_1044,N_18875,N_19858);
nor UO_1045 (O_1045,N_16984,N_19707);
and UO_1046 (O_1046,N_17232,N_19243);
xnor UO_1047 (O_1047,N_18074,N_17931);
xor UO_1048 (O_1048,N_18210,N_17882);
nor UO_1049 (O_1049,N_19448,N_18711);
nand UO_1050 (O_1050,N_17014,N_19601);
or UO_1051 (O_1051,N_16670,N_16403);
nor UO_1052 (O_1052,N_17209,N_16098);
or UO_1053 (O_1053,N_19231,N_19944);
nor UO_1054 (O_1054,N_18872,N_18225);
or UO_1055 (O_1055,N_17331,N_19310);
or UO_1056 (O_1056,N_16630,N_16568);
xnor UO_1057 (O_1057,N_17367,N_18508);
nor UO_1058 (O_1058,N_19838,N_18822);
and UO_1059 (O_1059,N_16621,N_17570);
and UO_1060 (O_1060,N_18391,N_19544);
or UO_1061 (O_1061,N_16348,N_19337);
xnor UO_1062 (O_1062,N_16317,N_18511);
nand UO_1063 (O_1063,N_17413,N_18580);
nand UO_1064 (O_1064,N_18350,N_17388);
or UO_1065 (O_1065,N_16253,N_18148);
nand UO_1066 (O_1066,N_18553,N_19534);
nor UO_1067 (O_1067,N_18652,N_16903);
nor UO_1068 (O_1068,N_17000,N_18807);
nor UO_1069 (O_1069,N_19361,N_19263);
and UO_1070 (O_1070,N_17447,N_19800);
nor UO_1071 (O_1071,N_16803,N_18841);
xor UO_1072 (O_1072,N_18159,N_16190);
and UO_1073 (O_1073,N_18932,N_19954);
and UO_1074 (O_1074,N_17039,N_16600);
xor UO_1075 (O_1075,N_18398,N_19408);
or UO_1076 (O_1076,N_18339,N_18068);
nand UO_1077 (O_1077,N_19744,N_19188);
nand UO_1078 (O_1078,N_18276,N_17902);
and UO_1079 (O_1079,N_19182,N_18916);
or UO_1080 (O_1080,N_18152,N_18487);
and UO_1081 (O_1081,N_16657,N_16665);
and UO_1082 (O_1082,N_18937,N_17973);
nand UO_1083 (O_1083,N_16483,N_17226);
nand UO_1084 (O_1084,N_17946,N_17893);
nand UO_1085 (O_1085,N_17400,N_18132);
nand UO_1086 (O_1086,N_16933,N_18037);
nand UO_1087 (O_1087,N_18440,N_17874);
or UO_1088 (O_1088,N_16547,N_18028);
nor UO_1089 (O_1089,N_19526,N_16896);
nor UO_1090 (O_1090,N_18397,N_16412);
and UO_1091 (O_1091,N_17314,N_16850);
xor UO_1092 (O_1092,N_18619,N_16907);
and UO_1093 (O_1093,N_16845,N_18963);
and UO_1094 (O_1094,N_18576,N_19929);
xnor UO_1095 (O_1095,N_17700,N_18214);
nor UO_1096 (O_1096,N_18744,N_17243);
and UO_1097 (O_1097,N_17797,N_19271);
or UO_1098 (O_1098,N_18231,N_17422);
xor UO_1099 (O_1099,N_17205,N_16633);
xor UO_1100 (O_1100,N_19180,N_16500);
nand UO_1101 (O_1101,N_16042,N_17754);
and UO_1102 (O_1102,N_16493,N_19925);
nand UO_1103 (O_1103,N_18474,N_18092);
nor UO_1104 (O_1104,N_18166,N_17942);
xnor UO_1105 (O_1105,N_19622,N_17066);
nand UO_1106 (O_1106,N_17173,N_19411);
nor UO_1107 (O_1107,N_18284,N_16306);
xor UO_1108 (O_1108,N_19118,N_18658);
xor UO_1109 (O_1109,N_17036,N_18264);
xor UO_1110 (O_1110,N_16735,N_18107);
nand UO_1111 (O_1111,N_18731,N_16312);
or UO_1112 (O_1112,N_18974,N_19879);
xor UO_1113 (O_1113,N_17543,N_18460);
xor UO_1114 (O_1114,N_17309,N_17849);
nand UO_1115 (O_1115,N_18013,N_19881);
or UO_1116 (O_1116,N_19557,N_19003);
or UO_1117 (O_1117,N_17317,N_17396);
or UO_1118 (O_1118,N_17312,N_17733);
nor UO_1119 (O_1119,N_19013,N_17485);
nor UO_1120 (O_1120,N_19878,N_19835);
and UO_1121 (O_1121,N_17085,N_16281);
nand UO_1122 (O_1122,N_17935,N_18341);
or UO_1123 (O_1123,N_16580,N_18220);
nand UO_1124 (O_1124,N_18364,N_18197);
nor UO_1125 (O_1125,N_16297,N_16006);
or UO_1126 (O_1126,N_16101,N_18083);
or UO_1127 (O_1127,N_16144,N_18307);
nor UO_1128 (O_1128,N_16243,N_19483);
nand UO_1129 (O_1129,N_16956,N_18554);
and UO_1130 (O_1130,N_17768,N_17287);
xnor UO_1131 (O_1131,N_17708,N_16604);
xor UO_1132 (O_1132,N_18049,N_16358);
xnor UO_1133 (O_1133,N_16681,N_17163);
nor UO_1134 (O_1134,N_16419,N_17118);
nand UO_1135 (O_1135,N_16382,N_18229);
xnor UO_1136 (O_1136,N_16816,N_18354);
nor UO_1137 (O_1137,N_16516,N_18449);
or UO_1138 (O_1138,N_19607,N_18034);
nor UO_1139 (O_1139,N_19657,N_18943);
nand UO_1140 (O_1140,N_16189,N_17046);
xnor UO_1141 (O_1141,N_19009,N_17023);
nor UO_1142 (O_1142,N_16003,N_17599);
xnor UO_1143 (O_1143,N_18077,N_18924);
nand UO_1144 (O_1144,N_17786,N_18838);
and UO_1145 (O_1145,N_17647,N_19430);
and UO_1146 (O_1146,N_19722,N_16802);
nor UO_1147 (O_1147,N_17761,N_18075);
nor UO_1148 (O_1148,N_19277,N_17983);
nand UO_1149 (O_1149,N_16818,N_19278);
nand UO_1150 (O_1150,N_16345,N_16273);
nand UO_1151 (O_1151,N_16682,N_17972);
or UO_1152 (O_1152,N_16614,N_18596);
and UO_1153 (O_1153,N_18930,N_16626);
nor UO_1154 (O_1154,N_18141,N_18632);
and UO_1155 (O_1155,N_17265,N_17937);
xnor UO_1156 (O_1156,N_19580,N_16305);
and UO_1157 (O_1157,N_16171,N_16052);
and UO_1158 (O_1158,N_18478,N_17936);
or UO_1159 (O_1159,N_18384,N_18379);
xor UO_1160 (O_1160,N_16587,N_18531);
nand UO_1161 (O_1161,N_16575,N_19369);
or UO_1162 (O_1162,N_18190,N_18793);
xor UO_1163 (O_1163,N_19204,N_17448);
nor UO_1164 (O_1164,N_18832,N_16698);
nor UO_1165 (O_1165,N_19394,N_17857);
xnor UO_1166 (O_1166,N_17238,N_17810);
nand UO_1167 (O_1167,N_19343,N_19218);
and UO_1168 (O_1168,N_17524,N_18550);
or UO_1169 (O_1169,N_18544,N_17883);
or UO_1170 (O_1170,N_18043,N_18259);
xor UO_1171 (O_1171,N_19330,N_16308);
nor UO_1172 (O_1172,N_18395,N_16578);
or UO_1173 (O_1173,N_19471,N_19610);
nor UO_1174 (O_1174,N_18641,N_18896);
and UO_1175 (O_1175,N_19226,N_16301);
and UO_1176 (O_1176,N_19955,N_16266);
xor UO_1177 (O_1177,N_19751,N_18111);
and UO_1178 (O_1178,N_19076,N_16921);
nand UO_1179 (O_1179,N_17135,N_19328);
and UO_1180 (O_1180,N_18860,N_17093);
and UO_1181 (O_1181,N_17071,N_18942);
nand UO_1182 (O_1182,N_19475,N_17765);
nor UO_1183 (O_1183,N_16423,N_16696);
xnor UO_1184 (O_1184,N_19098,N_19904);
nor UO_1185 (O_1185,N_16062,N_19720);
or UO_1186 (O_1186,N_19478,N_17913);
or UO_1187 (O_1187,N_18479,N_17303);
nor UO_1188 (O_1188,N_18103,N_17147);
or UO_1189 (O_1189,N_19571,N_16360);
nand UO_1190 (O_1190,N_17390,N_18360);
and UO_1191 (O_1191,N_19624,N_17692);
xnor UO_1192 (O_1192,N_16655,N_18066);
or UO_1193 (O_1193,N_17177,N_18048);
nand UO_1194 (O_1194,N_18870,N_16286);
or UO_1195 (O_1195,N_16224,N_16955);
or UO_1196 (O_1196,N_19422,N_16659);
nand UO_1197 (O_1197,N_17440,N_19209);
nor UO_1198 (O_1198,N_18378,N_16038);
nor UO_1199 (O_1199,N_17349,N_19319);
xnor UO_1200 (O_1200,N_19874,N_18357);
and UO_1201 (O_1201,N_16504,N_19849);
and UO_1202 (O_1202,N_19641,N_16563);
xor UO_1203 (O_1203,N_18326,N_17775);
xor UO_1204 (O_1204,N_17683,N_19980);
nand UO_1205 (O_1205,N_18022,N_19566);
nand UO_1206 (O_1206,N_18599,N_18506);
or UO_1207 (O_1207,N_16212,N_17602);
or UO_1208 (O_1208,N_17758,N_19970);
nor UO_1209 (O_1209,N_18688,N_17346);
or UO_1210 (O_1210,N_19602,N_18823);
xor UO_1211 (O_1211,N_17633,N_19674);
and UO_1212 (O_1212,N_19085,N_18423);
nand UO_1213 (O_1213,N_19913,N_16981);
or UO_1214 (O_1214,N_18977,N_16628);
nor UO_1215 (O_1215,N_16640,N_16264);
nor UO_1216 (O_1216,N_18534,N_17263);
nand UO_1217 (O_1217,N_18842,N_18483);
nor UO_1218 (O_1218,N_17666,N_19851);
or UO_1219 (O_1219,N_18622,N_16070);
nand UO_1220 (O_1220,N_17219,N_16114);
nand UO_1221 (O_1221,N_17637,N_18162);
nand UO_1222 (O_1222,N_19706,N_16482);
or UO_1223 (O_1223,N_19603,N_19467);
nor UO_1224 (O_1224,N_19947,N_17338);
and UO_1225 (O_1225,N_19825,N_18677);
and UO_1226 (O_1226,N_17286,N_17456);
and UO_1227 (O_1227,N_17300,N_16742);
xor UO_1228 (O_1228,N_18893,N_18741);
xnor UO_1229 (O_1229,N_16879,N_17648);
xnor UO_1230 (O_1230,N_19354,N_19353);
nor UO_1231 (O_1231,N_18230,N_19396);
nand UO_1232 (O_1232,N_17687,N_17840);
nand UO_1233 (O_1233,N_18537,N_18216);
xnor UO_1234 (O_1234,N_18913,N_16227);
or UO_1235 (O_1235,N_18414,N_18847);
nand UO_1236 (O_1236,N_16608,N_17094);
or UO_1237 (O_1237,N_17583,N_18523);
or UO_1238 (O_1238,N_17065,N_16406);
and UO_1239 (O_1239,N_16151,N_16010);
and UO_1240 (O_1240,N_18659,N_17382);
nor UO_1241 (O_1241,N_16359,N_18655);
nand UO_1242 (O_1242,N_17984,N_19484);
and UO_1243 (O_1243,N_17062,N_17867);
and UO_1244 (O_1244,N_19888,N_19393);
nand UO_1245 (O_1245,N_18445,N_18126);
xnor UO_1246 (O_1246,N_17702,N_17766);
nand UO_1247 (O_1247,N_16567,N_18962);
nand UO_1248 (O_1248,N_18091,N_19535);
nor UO_1249 (O_1249,N_18179,N_16427);
nor UO_1250 (O_1250,N_16352,N_16871);
and UO_1251 (O_1251,N_17127,N_16124);
and UO_1252 (O_1252,N_19914,N_17564);
nand UO_1253 (O_1253,N_16145,N_19645);
or UO_1254 (O_1254,N_18112,N_17480);
nor UO_1255 (O_1255,N_17077,N_18120);
nor UO_1256 (O_1256,N_18653,N_18404);
or UO_1257 (O_1257,N_17886,N_18742);
nor UO_1258 (O_1258,N_16577,N_19469);
xnor UO_1259 (O_1259,N_18281,N_18552);
nor UO_1260 (O_1260,N_16758,N_18961);
or UO_1261 (O_1261,N_16076,N_18052);
and UO_1262 (O_1262,N_19529,N_16393);
nor UO_1263 (O_1263,N_17519,N_19538);
and UO_1264 (O_1264,N_17587,N_18476);
and UO_1265 (O_1265,N_16221,N_16560);
or UO_1266 (O_1266,N_17299,N_19301);
nand UO_1267 (O_1267,N_16367,N_18142);
xor UO_1268 (O_1268,N_17554,N_19567);
and UO_1269 (O_1269,N_16466,N_19660);
xnor UO_1270 (O_1270,N_18627,N_19918);
and UO_1271 (O_1271,N_16954,N_19470);
nor UO_1272 (O_1272,N_17927,N_16755);
nor UO_1273 (O_1273,N_17516,N_19697);
xnor UO_1274 (O_1274,N_17960,N_19952);
or UO_1275 (O_1275,N_16473,N_17027);
xnor UO_1276 (O_1276,N_19705,N_18827);
nor UO_1277 (O_1277,N_17368,N_18497);
nor UO_1278 (O_1278,N_17577,N_17614);
or UO_1279 (O_1279,N_16542,N_16257);
nand UO_1280 (O_1280,N_16505,N_16723);
and UO_1281 (O_1281,N_17455,N_17436);
nor UO_1282 (O_1282,N_17923,N_16886);
and UO_1283 (O_1283,N_19901,N_19782);
or UO_1284 (O_1284,N_17688,N_19092);
nand UO_1285 (O_1285,N_18748,N_18296);
and UO_1286 (O_1286,N_17130,N_18237);
nor UO_1287 (O_1287,N_19356,N_18968);
xor UO_1288 (O_1288,N_18046,N_18586);
nor UO_1289 (O_1289,N_17026,N_16453);
and UO_1290 (O_1290,N_18221,N_19834);
or UO_1291 (O_1291,N_18261,N_17414);
and UO_1292 (O_1292,N_16512,N_19746);
and UO_1293 (O_1293,N_17679,N_19049);
and UO_1294 (O_1294,N_17771,N_16650);
xnor UO_1295 (O_1295,N_18115,N_18701);
or UO_1296 (O_1296,N_19306,N_16206);
or UO_1297 (O_1297,N_18858,N_17686);
nand UO_1298 (O_1298,N_17352,N_19323);
nand UO_1299 (O_1299,N_16641,N_19219);
nand UO_1300 (O_1300,N_19439,N_19924);
nor UO_1301 (O_1301,N_18657,N_17514);
nand UO_1302 (O_1302,N_18579,N_18021);
xnor UO_1303 (O_1303,N_18499,N_18649);
nor UO_1304 (O_1304,N_19670,N_19691);
and UO_1305 (O_1305,N_17650,N_19193);
nor UO_1306 (O_1306,N_18002,N_17861);
xnor UO_1307 (O_1307,N_18383,N_18999);
and UO_1308 (O_1308,N_18472,N_18526);
and UO_1309 (O_1309,N_17834,N_17213);
xnor UO_1310 (O_1310,N_19824,N_17908);
or UO_1311 (O_1311,N_17340,N_18691);
or UO_1312 (O_1312,N_18250,N_19043);
and UO_1313 (O_1313,N_18375,N_16704);
nand UO_1314 (O_1314,N_16256,N_17137);
nor UO_1315 (O_1315,N_16553,N_19818);
and UO_1316 (O_1316,N_17357,N_19349);
nand UO_1317 (O_1317,N_16502,N_18486);
xor UO_1318 (O_1318,N_18485,N_18467);
nand UO_1319 (O_1319,N_16656,N_16082);
nor UO_1320 (O_1320,N_17222,N_18714);
or UO_1321 (O_1321,N_18137,N_19592);
nor UO_1322 (O_1322,N_16736,N_16295);
and UO_1323 (O_1323,N_18761,N_16102);
nand UO_1324 (O_1324,N_16012,N_19195);
and UO_1325 (O_1325,N_17032,N_19106);
and UO_1326 (O_1326,N_17498,N_19577);
and UO_1327 (O_1327,N_16602,N_19156);
nor UO_1328 (O_1328,N_16450,N_19086);
and UO_1329 (O_1329,N_17457,N_19773);
xnor UO_1330 (O_1330,N_17067,N_17748);
nor UO_1331 (O_1331,N_17427,N_17115);
nand UO_1332 (O_1332,N_16796,N_17517);
and UO_1333 (O_1333,N_18787,N_17099);
or UO_1334 (O_1334,N_16371,N_19017);
nand UO_1335 (O_1335,N_19761,N_17695);
xnor UO_1336 (O_1336,N_18410,N_18089);
nand UO_1337 (O_1337,N_16631,N_19753);
nor UO_1338 (O_1338,N_19398,N_18439);
nand UO_1339 (O_1339,N_16866,N_18056);
nor UO_1340 (O_1340,N_17875,N_17371);
and UO_1341 (O_1341,N_19708,N_16083);
or UO_1342 (O_1342,N_16780,N_19558);
nor UO_1343 (O_1343,N_16993,N_18338);
nor UO_1344 (O_1344,N_17845,N_18236);
nand UO_1345 (O_1345,N_18575,N_17868);
or UO_1346 (O_1346,N_17616,N_18150);
and UO_1347 (O_1347,N_19435,N_19648);
nor UO_1348 (O_1348,N_19715,N_19447);
or UO_1349 (O_1349,N_16161,N_17854);
or UO_1350 (O_1350,N_19554,N_16471);
and UO_1351 (O_1351,N_18452,N_16361);
or UO_1352 (O_1352,N_17909,N_16821);
nor UO_1353 (O_1353,N_19591,N_18018);
xnor UO_1354 (O_1354,N_18829,N_18175);
nor UO_1355 (O_1355,N_19619,N_17767);
nor UO_1356 (O_1356,N_16001,N_18151);
and UO_1357 (O_1357,N_16377,N_17872);
or UO_1358 (O_1358,N_19875,N_17284);
and UO_1359 (O_1359,N_18584,N_17977);
nor UO_1360 (O_1360,N_18362,N_19634);
or UO_1361 (O_1361,N_17553,N_16679);
or UO_1362 (O_1362,N_18211,N_19453);
and UO_1363 (O_1363,N_18444,N_19500);
nand UO_1364 (O_1364,N_18108,N_18585);
xnor UO_1365 (O_1365,N_17725,N_16149);
xnor UO_1366 (O_1366,N_16624,N_16814);
or UO_1367 (O_1367,N_16064,N_18941);
nor UO_1368 (O_1368,N_17948,N_16922);
nor UO_1369 (O_1369,N_16857,N_16472);
nand UO_1370 (O_1370,N_17188,N_17452);
or UO_1371 (O_1371,N_19802,N_17361);
nand UO_1372 (O_1372,N_18411,N_18770);
nor UO_1373 (O_1373,N_18789,N_18804);
xor UO_1374 (O_1374,N_19938,N_19417);
or UO_1375 (O_1375,N_19146,N_16690);
or UO_1376 (O_1376,N_18734,N_16977);
or UO_1377 (O_1377,N_17133,N_16538);
xnor UO_1378 (O_1378,N_16720,N_19395);
nand UO_1379 (O_1379,N_16693,N_17734);
xor UO_1380 (O_1380,N_16481,N_18510);
or UO_1381 (O_1381,N_17701,N_16069);
nor UO_1382 (O_1382,N_19207,N_19569);
nand UO_1383 (O_1383,N_18774,N_16792);
xor UO_1384 (O_1384,N_16651,N_17041);
xor UO_1385 (O_1385,N_19205,N_17814);
and UO_1386 (O_1386,N_19831,N_18840);
xor UO_1387 (O_1387,N_18319,N_19736);
or UO_1388 (O_1388,N_16928,N_16005);
nand UO_1389 (O_1389,N_16384,N_17419);
nand UO_1390 (O_1390,N_19808,N_19414);
nand UO_1391 (O_1391,N_19083,N_16416);
or UO_1392 (O_1392,N_16895,N_18006);
or UO_1393 (O_1393,N_18004,N_19786);
nor UO_1394 (O_1394,N_19948,N_18059);
xor UO_1395 (O_1395,N_19703,N_18407);
or UO_1396 (O_1396,N_18773,N_17473);
xnor UO_1397 (O_1397,N_16644,N_17511);
or UO_1398 (O_1398,N_17237,N_18833);
nand UO_1399 (O_1399,N_19145,N_16165);
or UO_1400 (O_1400,N_18031,N_17635);
nor UO_1401 (O_1401,N_18788,N_19446);
and UO_1402 (O_1402,N_19596,N_19609);
xor UO_1403 (O_1403,N_19327,N_17431);
or UO_1404 (O_1404,N_16618,N_17694);
nand UO_1405 (O_1405,N_16979,N_16092);
or UO_1406 (O_1406,N_19292,N_17462);
xor UO_1407 (O_1407,N_17101,N_18885);
nor UO_1408 (O_1408,N_19829,N_16240);
and UO_1409 (O_1409,N_19312,N_18908);
xnor UO_1410 (O_1410,N_18960,N_19149);
nor UO_1411 (O_1411,N_19512,N_17901);
nor UO_1412 (O_1412,N_17532,N_19044);
nand UO_1413 (O_1413,N_18408,N_17442);
nand UO_1414 (O_1414,N_18093,N_18654);
nand UO_1415 (O_1415,N_18880,N_17556);
xor UO_1416 (O_1416,N_18934,N_16390);
nor UO_1417 (O_1417,N_17951,N_19325);
and UO_1418 (O_1418,N_19667,N_19912);
nor UO_1419 (O_1419,N_18616,N_16294);
nor UO_1420 (O_1420,N_19576,N_18821);
and UO_1421 (O_1421,N_16998,N_16029);
xnor UO_1422 (O_1422,N_18060,N_19939);
xor UO_1423 (O_1423,N_16545,N_19201);
and UO_1424 (O_1424,N_19384,N_16037);
and UO_1425 (O_1425,N_16842,N_17499);
or UO_1426 (O_1426,N_18676,N_17342);
and UO_1427 (O_1427,N_16207,N_19730);
or UO_1428 (O_1428,N_19847,N_19372);
nand UO_1429 (O_1429,N_18535,N_18367);
and UO_1430 (O_1430,N_17880,N_19712);
xnor UO_1431 (O_1431,N_18470,N_19588);
or UO_1432 (O_1432,N_16050,N_19418);
xor UO_1433 (O_1433,N_16680,N_16559);
nor UO_1434 (O_1434,N_16806,N_18957);
nand UO_1435 (O_1435,N_17104,N_16525);
and UO_1436 (O_1436,N_16014,N_16964);
nand UO_1437 (O_1437,N_18921,N_16039);
or UO_1438 (O_1438,N_19359,N_19060);
and UO_1439 (O_1439,N_17290,N_17627);
and UO_1440 (O_1440,N_17389,N_18128);
nand UO_1441 (O_1441,N_18094,N_16182);
nor UO_1442 (O_1442,N_16214,N_19225);
xor UO_1443 (O_1443,N_19311,N_17109);
xor UO_1444 (O_1444,N_18312,N_19684);
and UO_1445 (O_1445,N_17665,N_18757);
or UO_1446 (O_1446,N_18903,N_18392);
xnor UO_1447 (O_1447,N_19303,N_17728);
xnor UO_1448 (O_1448,N_19383,N_16437);
and UO_1449 (O_1449,N_19989,N_18456);
nand UO_1450 (O_1450,N_19699,N_16829);
nand UO_1451 (O_1451,N_18561,N_17791);
or UO_1452 (O_1452,N_17677,N_19131);
nand UO_1453 (O_1453,N_19253,N_19499);
or UO_1454 (O_1454,N_17402,N_19032);
or UO_1455 (O_1455,N_19994,N_16084);
nand UO_1456 (O_1456,N_16375,N_18071);
nor UO_1457 (O_1457,N_18808,N_16285);
nand UO_1458 (O_1458,N_16669,N_17673);
and UO_1459 (O_1459,N_16884,N_19260);
nor UO_1460 (O_1460,N_17397,N_17989);
or UO_1461 (O_1461,N_18178,N_18365);
nor UO_1462 (O_1462,N_19035,N_16594);
nor UO_1463 (O_1463,N_19870,N_19574);
xor UO_1464 (O_1464,N_16475,N_17105);
or UO_1465 (O_1465,N_18212,N_17928);
or UO_1466 (O_1466,N_17348,N_19203);
nand UO_1467 (O_1467,N_18918,N_17002);
xor UO_1468 (O_1468,N_17601,N_16810);
xor UO_1469 (O_1469,N_16940,N_16910);
xnor UO_1470 (O_1470,N_16583,N_16081);
nor UO_1471 (O_1471,N_17011,N_19987);
or UO_1472 (O_1472,N_19630,N_17918);
nor UO_1473 (O_1473,N_17896,N_17078);
nor UO_1474 (O_1474,N_18412,N_19036);
and UO_1475 (O_1475,N_18185,N_17050);
and UO_1476 (O_1476,N_18204,N_18724);
nor UO_1477 (O_1477,N_18238,N_16763);
xor UO_1478 (O_1478,N_19472,N_16392);
nor UO_1479 (O_1479,N_19169,N_19852);
nand UO_1480 (O_1480,N_18029,N_16906);
and UO_1481 (O_1481,N_19953,N_17492);
nand UO_1482 (O_1482,N_18243,N_16293);
nand UO_1483 (O_1483,N_18215,N_19376);
xnor UO_1484 (O_1484,N_19998,N_19241);
nand UO_1485 (O_1485,N_16694,N_17661);
and UO_1486 (O_1486,N_18547,N_17581);
and UO_1487 (O_1487,N_19960,N_17081);
xnor UO_1488 (O_1488,N_19959,N_18451);
nand UO_1489 (O_1489,N_16917,N_18069);
nor UO_1490 (O_1490,N_19932,N_19111);
nand UO_1491 (O_1491,N_16722,N_16936);
xor UO_1492 (O_1492,N_17254,N_16007);
xor UO_1493 (O_1493,N_19513,N_17726);
xnor UO_1494 (O_1494,N_16046,N_16749);
nand UO_1495 (O_1495,N_18509,N_16430);
and UO_1496 (O_1496,N_18519,N_18464);
nand UO_1497 (O_1497,N_17690,N_18294);
nand UO_1498 (O_1498,N_16168,N_17546);
nor UO_1499 (O_1499,N_19935,N_18503);
nand UO_1500 (O_1500,N_19550,N_16787);
nor UO_1501 (O_1501,N_17757,N_16554);
nand UO_1502 (O_1502,N_18777,N_16752);
nand UO_1503 (O_1503,N_17244,N_16120);
nor UO_1504 (O_1504,N_19934,N_19545);
nand UO_1505 (O_1505,N_16116,N_19597);
xor UO_1506 (O_1506,N_17772,N_17496);
and UO_1507 (O_1507,N_19823,N_18820);
or UO_1508 (O_1508,N_17529,N_19307);
and UO_1509 (O_1509,N_17230,N_19757);
nand UO_1510 (O_1510,N_16388,N_18831);
nand UO_1511 (O_1511,N_19400,N_18368);
and UO_1512 (O_1512,N_17813,N_18133);
and UO_1513 (O_1513,N_18050,N_17969);
and UO_1514 (O_1514,N_18324,N_16087);
nor UO_1515 (O_1515,N_16601,N_19412);
or UO_1516 (O_1516,N_18710,N_19296);
nand UO_1517 (O_1517,N_17201,N_18984);
nor UO_1518 (O_1518,N_16409,N_17223);
nor UO_1519 (O_1519,N_17851,N_16923);
xnor UO_1520 (O_1520,N_18668,N_17424);
xnor UO_1521 (O_1521,N_17645,N_16410);
xor UO_1522 (O_1522,N_18198,N_19104);
or UO_1523 (O_1523,N_19606,N_17709);
and UO_1524 (O_1524,N_17634,N_19968);
and UO_1525 (O_1525,N_16916,N_19805);
xor UO_1526 (O_1526,N_19910,N_18442);
nor UO_1527 (O_1527,N_17737,N_17323);
or UO_1528 (O_1528,N_16754,N_17240);
nand UO_1529 (O_1529,N_18109,N_17487);
or UO_1530 (O_1530,N_16459,N_17961);
nor UO_1531 (O_1531,N_16747,N_17074);
and UO_1532 (O_1532,N_19159,N_18802);
xnor UO_1533 (O_1533,N_16848,N_19362);
and UO_1534 (O_1534,N_16488,N_16901);
nor UO_1535 (O_1535,N_19154,N_19333);
or UO_1536 (O_1536,N_17592,N_17106);
xnor UO_1537 (O_1537,N_18097,N_16491);
or UO_1538 (O_1538,N_18911,N_16800);
and UO_1539 (O_1539,N_17197,N_19189);
and UO_1540 (O_1540,N_16713,N_16714);
nor UO_1541 (O_1541,N_18288,N_16486);
nor UO_1542 (O_1542,N_16772,N_19552);
xnor UO_1543 (O_1543,N_19741,N_16785);
xor UO_1544 (O_1544,N_18234,N_17557);
nor UO_1545 (O_1545,N_18861,N_17970);
and UO_1546 (O_1546,N_16205,N_18116);
or UO_1547 (O_1547,N_17144,N_18560);
nor UO_1548 (O_1548,N_16637,N_16576);
or UO_1549 (O_1549,N_19759,N_18762);
nor UO_1550 (O_1550,N_17038,N_17736);
and UO_1551 (O_1551,N_17178,N_18080);
nand UO_1552 (O_1552,N_16047,N_19839);
nor UO_1553 (O_1553,N_18246,N_18781);
xor UO_1554 (O_1554,N_17997,N_16133);
nand UO_1555 (O_1555,N_16897,N_18529);
and UO_1556 (O_1556,N_16299,N_17724);
nor UO_1557 (O_1557,N_19170,N_16882);
xor UO_1558 (O_1558,N_18274,N_17600);
and UO_1559 (O_1559,N_18042,N_19079);
and UO_1560 (O_1560,N_17472,N_18265);
xnor UO_1561 (O_1561,N_19381,N_18000);
nor UO_1562 (O_1562,N_17612,N_18369);
nand UO_1563 (O_1563,N_16362,N_19899);
xor UO_1564 (O_1564,N_18072,N_16737);
nor UO_1565 (O_1565,N_19669,N_18517);
xnor UO_1566 (O_1566,N_18457,N_17668);
nand UO_1567 (O_1567,N_19909,N_18167);
xnor UO_1568 (O_1568,N_19107,N_19025);
nor UO_1569 (O_1569,N_19371,N_19579);
nand UO_1570 (O_1570,N_16521,N_16773);
xnor UO_1571 (O_1571,N_17789,N_18695);
nor UO_1572 (O_1572,N_19916,N_16515);
xor UO_1573 (O_1573,N_18785,N_17655);
or UO_1574 (O_1574,N_18873,N_16132);
nand UO_1575 (O_1575,N_16905,N_16467);
and UO_1576 (O_1576,N_17841,N_18679);
and UO_1577 (O_1577,N_17520,N_18992);
xnor UO_1578 (O_1578,N_19504,N_18740);
nand UO_1579 (O_1579,N_16455,N_19373);
xor UO_1580 (O_1580,N_17699,N_19560);
xnor UO_1581 (O_1581,N_18926,N_16036);
nand UO_1582 (O_1582,N_17393,N_19062);
or UO_1583 (O_1583,N_19540,N_17870);
xor UO_1584 (O_1584,N_17588,N_19678);
and UO_1585 (O_1585,N_18269,N_18750);
or UO_1586 (O_1586,N_19771,N_19459);
or UO_1587 (O_1587,N_19668,N_19364);
nor UO_1588 (O_1588,N_19134,N_17061);
nor UO_1589 (O_1589,N_19506,N_19531);
or UO_1590 (O_1590,N_19643,N_19546);
and UO_1591 (O_1591,N_16613,N_16739);
and UO_1592 (O_1592,N_19748,N_17574);
and UO_1593 (O_1593,N_19816,N_17211);
nand UO_1594 (O_1594,N_18168,N_17103);
or UO_1595 (O_1595,N_16405,N_19616);
and UO_1596 (O_1596,N_19456,N_19339);
and UO_1597 (O_1597,N_18601,N_17566);
nand UO_1598 (O_1598,N_16381,N_16572);
xnor UO_1599 (O_1599,N_16170,N_18725);
nand UO_1600 (O_1600,N_16045,N_18361);
nand UO_1601 (O_1601,N_17798,N_18203);
xor UO_1602 (O_1602,N_17685,N_19514);
nor UO_1603 (O_1603,N_17212,N_16862);
and UO_1604 (O_1604,N_17822,N_16571);
xnor UO_1605 (O_1605,N_18462,N_19503);
or UO_1606 (O_1606,N_17866,N_19687);
nand UO_1607 (O_1607,N_18703,N_17785);
or UO_1608 (O_1608,N_17515,N_16134);
xor UO_1609 (O_1609,N_16667,N_17711);
nand UO_1610 (O_1610,N_16929,N_16974);
xor UO_1611 (O_1611,N_16795,N_19251);
and UO_1612 (O_1612,N_19896,N_18813);
nand UO_1613 (O_1613,N_17292,N_17295);
and UO_1614 (O_1614,N_18784,N_19756);
or UO_1615 (O_1615,N_18118,N_17890);
nand UO_1616 (O_1616,N_16178,N_17007);
or UO_1617 (O_1617,N_18327,N_16461);
xnor UO_1618 (O_1618,N_17720,N_19997);
xnor UO_1619 (O_1619,N_17459,N_19210);
nor UO_1620 (O_1620,N_19642,N_19763);
or UO_1621 (O_1621,N_18161,N_17015);
nand UO_1622 (O_1622,N_16241,N_19324);
nor UO_1623 (O_1623,N_16564,N_17354);
nor UO_1624 (O_1624,N_18522,N_18453);
xor UO_1625 (O_1625,N_18380,N_16878);
nor UO_1626 (O_1626,N_17281,N_19798);
xor UO_1627 (O_1627,N_17221,N_17410);
nand UO_1628 (O_1628,N_17282,N_16421);
xnor UO_1629 (O_1629,N_19842,N_16443);
nand UO_1630 (O_1630,N_16447,N_19132);
xor UO_1631 (O_1631,N_18598,N_17160);
nor UO_1632 (O_1632,N_16861,N_16079);
or UO_1633 (O_1633,N_18219,N_19649);
xnor UO_1634 (O_1634,N_17401,N_17220);
nor UO_1635 (O_1635,N_18257,N_17940);
nand UO_1636 (O_1636,N_18602,N_16731);
nor UO_1637 (O_1637,N_17241,N_18359);
nor UO_1638 (O_1638,N_17530,N_18447);
or UO_1639 (O_1639,N_18347,N_18313);
and UO_1640 (O_1640,N_19840,N_16982);
nor UO_1641 (O_1641,N_16868,N_17609);
nand UO_1642 (O_1642,N_17047,N_18139);
or UO_1643 (O_1643,N_16840,N_17370);
nand UO_1644 (O_1644,N_16674,N_17048);
nand UO_1645 (O_1645,N_16654,N_16090);
xnor UO_1646 (O_1646,N_17562,N_16770);
nor UO_1647 (O_1647,N_18826,N_19653);
xor UO_1648 (O_1648,N_16589,N_16851);
and UO_1649 (O_1649,N_16607,N_18435);
xor UO_1650 (O_1650,N_19281,N_19173);
and UO_1651 (O_1651,N_17426,N_18583);
nand UO_1652 (O_1652,N_16199,N_16738);
nor UO_1653 (O_1653,N_16397,N_19239);
and UO_1654 (O_1654,N_17925,N_18481);
or UO_1655 (O_1655,N_18824,N_19562);
xor UO_1656 (O_1656,N_18217,N_17636);
xnor UO_1657 (O_1657,N_19410,N_17251);
or UO_1658 (O_1658,N_17253,N_18527);
xor UO_1659 (O_1659,N_19039,N_16822);
nand UO_1660 (O_1660,N_17228,N_16004);
xor UO_1661 (O_1661,N_16233,N_19421);
xnor UO_1662 (O_1662,N_19160,N_17330);
or UO_1663 (O_1663,N_18242,N_16541);
nand UO_1664 (O_1664,N_17774,N_18610);
xnor UO_1665 (O_1665,N_16768,N_18839);
and UO_1666 (O_1666,N_18370,N_17096);
nor UO_1667 (O_1667,N_17717,N_19380);
nand UO_1668 (O_1668,N_16407,N_19286);
nand UO_1669 (O_1669,N_18199,N_18923);
and UO_1670 (O_1670,N_17899,N_19933);
and UO_1671 (O_1671,N_16931,N_19093);
or UO_1672 (O_1672,N_19845,N_16653);
nor UO_1673 (O_1673,N_17146,N_19637);
or UO_1674 (O_1674,N_17356,N_18095);
and UO_1675 (O_1675,N_19781,N_19335);
or UO_1676 (O_1676,N_19437,N_17563);
or UO_1677 (O_1677,N_19779,N_19527);
nand UO_1678 (O_1678,N_17416,N_19900);
nor UO_1679 (O_1679,N_19743,N_17479);
nor UO_1680 (O_1680,N_19021,N_17183);
xnor UO_1681 (O_1681,N_18528,N_18001);
nand UO_1682 (O_1682,N_19662,N_18226);
nand UO_1683 (O_1683,N_17049,N_17715);
or UO_1684 (O_1684,N_16915,N_18634);
and UO_1685 (O_1685,N_18922,N_18805);
or UO_1686 (O_1686,N_17862,N_19019);
and UO_1687 (O_1687,N_18157,N_19611);
xnor UO_1688 (O_1688,N_17610,N_17860);
and UO_1689 (O_1689,N_19917,N_19347);
nand UO_1690 (O_1690,N_18915,N_18618);
xnor UO_1691 (O_1691,N_18642,N_17628);
or UO_1692 (O_1692,N_17276,N_17275);
or UO_1693 (O_1693,N_16195,N_19787);
nor UO_1694 (O_1694,N_17920,N_19100);
or UO_1695 (O_1695,N_17052,N_19996);
nand UO_1696 (O_1696,N_16458,N_16451);
xor UO_1697 (O_1697,N_17844,N_16590);
or UO_1698 (O_1698,N_17632,N_19647);
or UO_1699 (O_1699,N_18501,N_17676);
nand UO_1700 (O_1700,N_18268,N_17248);
nand UO_1701 (O_1701,N_19046,N_18280);
nand UO_1702 (O_1702,N_16833,N_16811);
xor UO_1703 (O_1703,N_17712,N_16826);
nor UO_1704 (O_1704,N_17939,N_17894);
nor UO_1705 (O_1705,N_16373,N_17611);
nor UO_1706 (O_1706,N_17247,N_19054);
and UO_1707 (O_1707,N_16788,N_18302);
or UO_1708 (O_1708,N_18252,N_17398);
and UO_1709 (O_1709,N_16218,N_16555);
or UO_1710 (O_1710,N_19416,N_16112);
or UO_1711 (O_1711,N_18608,N_16514);
and UO_1712 (O_1712,N_19555,N_19462);
nand UO_1713 (O_1713,N_17161,N_18498);
nand UO_1714 (O_1714,N_18496,N_19223);
and UO_1715 (O_1715,N_19498,N_17004);
nor UO_1716 (O_1716,N_18228,N_18356);
xor UO_1717 (O_1717,N_18156,N_17216);
nand UO_1718 (O_1718,N_17776,N_17064);
or UO_1719 (O_1719,N_18171,N_18764);
xor UO_1720 (O_1720,N_16539,N_18790);
xor UO_1721 (O_1721,N_19906,N_16839);
nor UO_1722 (O_1722,N_19598,N_18978);
nor UO_1723 (O_1723,N_16913,N_19282);
and UO_1724 (O_1724,N_19992,N_19600);
nand UO_1725 (O_1725,N_18389,N_18996);
xor UO_1726 (O_1726,N_18438,N_19511);
and UO_1727 (O_1727,N_16330,N_18306);
or UO_1728 (O_1728,N_17684,N_16789);
nand UO_1729 (O_1729,N_17269,N_17578);
xor UO_1730 (O_1730,N_17006,N_16605);
xor UO_1731 (O_1731,N_18611,N_17261);
and UO_1732 (O_1732,N_18559,N_19516);
nor UO_1733 (O_1733,N_16097,N_16269);
or UO_1734 (O_1734,N_16143,N_19005);
or UO_1735 (O_1735,N_16364,N_18275);
and UO_1736 (O_1736,N_17034,N_18798);
or UO_1737 (O_1737,N_17092,N_18581);
or UO_1738 (O_1738,N_16217,N_16815);
nand UO_1739 (O_1739,N_16902,N_19828);
xor UO_1740 (O_1740,N_16900,N_18801);
and UO_1741 (O_1741,N_19436,N_18054);
nand UO_1742 (O_1742,N_19639,N_16683);
and UO_1743 (O_1743,N_17339,N_18455);
or UO_1744 (O_1744,N_19724,N_17200);
or UO_1745 (O_1745,N_17871,N_17166);
nor UO_1746 (O_1746,N_19297,N_18208);
nor UO_1747 (O_1747,N_18287,N_18812);
nor UO_1748 (O_1748,N_16888,N_16535);
nand UO_1749 (O_1749,N_18015,N_16147);
nor UO_1750 (O_1750,N_19138,N_18454);
xor UO_1751 (O_1751,N_16828,N_17155);
nor UO_1752 (O_1752,N_16139,N_16105);
nor UO_1753 (O_1753,N_19285,N_17171);
xnor UO_1754 (O_1754,N_19273,N_18405);
xor UO_1755 (O_1755,N_17329,N_19799);
xor UO_1756 (O_1756,N_16244,N_16864);
nor UO_1757 (O_1757,N_19521,N_18026);
nor UO_1758 (O_1758,N_18036,N_16856);
or UO_1759 (O_1759,N_17107,N_17590);
and UO_1760 (O_1760,N_19317,N_17905);
nand UO_1761 (O_1761,N_19178,N_16603);
xor UO_1762 (O_1762,N_17859,N_18845);
and UO_1763 (O_1763,N_18987,N_16561);
nor UO_1764 (O_1764,N_16452,N_17148);
and UO_1765 (O_1765,N_18129,N_17122);
nand UO_1766 (O_1766,N_16065,N_19982);
xor UO_1767 (O_1767,N_19999,N_17100);
or UO_1768 (O_1768,N_16663,N_18786);
or UO_1769 (O_1769,N_18016,N_19518);
nand UO_1770 (O_1770,N_16454,N_16355);
nand UO_1771 (O_1771,N_17328,N_16115);
nand UO_1772 (O_1772,N_17478,N_18394);
nand UO_1773 (O_1773,N_16890,N_17214);
and UO_1774 (O_1774,N_19050,N_16378);
or UO_1775 (O_1775,N_16751,N_17463);
or UO_1776 (O_1776,N_17812,N_16260);
or UO_1777 (O_1777,N_18612,N_19407);
nand UO_1778 (O_1778,N_18769,N_18385);
nand UO_1779 (O_1779,N_18729,N_18976);
nand UO_1780 (O_1780,N_17542,N_18879);
or UO_1781 (O_1781,N_19290,N_19140);
nor UO_1782 (O_1782,N_16543,N_19995);
nand UO_1783 (O_1783,N_16474,N_16357);
and UO_1784 (O_1784,N_16972,N_18852);
and UO_1785 (O_1785,N_16673,N_18775);
nor UO_1786 (O_1786,N_17850,N_19794);
or UO_1787 (O_1787,N_17449,N_17815);
or UO_1788 (O_1788,N_18980,N_17752);
or UO_1789 (O_1789,N_16019,N_16699);
xnor UO_1790 (O_1790,N_16870,N_17409);
xnor UO_1791 (O_1791,N_17159,N_16431);
xor UO_1792 (O_1792,N_19671,N_16891);
nand UO_1793 (O_1793,N_18427,N_19155);
xnor UO_1794 (O_1794,N_17274,N_19275);
and UO_1795 (O_1795,N_19739,N_16725);
or UO_1796 (O_1796,N_19029,N_18318);
or UO_1797 (O_1797,N_16376,N_17204);
xnor UO_1798 (O_1798,N_17465,N_17395);
xnor UO_1799 (O_1799,N_17060,N_17873);
nor UO_1800 (O_1800,N_16961,N_19322);
or UO_1801 (O_1801,N_16719,N_17528);
or UO_1802 (O_1802,N_17947,N_17521);
or UO_1803 (O_1803,N_19082,N_16204);
xnor UO_1804 (O_1804,N_19972,N_19257);
nor UO_1805 (O_1805,N_19168,N_19582);
or UO_1806 (O_1806,N_17035,N_16353);
xor UO_1807 (O_1807,N_19489,N_17830);
or UO_1808 (O_1808,N_18292,N_17017);
nor UO_1809 (O_1809,N_16225,N_19770);
or UO_1810 (O_1810,N_16322,N_18871);
nor UO_1811 (O_1811,N_16536,N_17495);
nand UO_1812 (O_1812,N_18493,N_18797);
xor UO_1813 (O_1813,N_17646,N_19262);
xnor UO_1814 (O_1814,N_19233,N_19951);
nand UO_1815 (O_1815,N_17907,N_19305);
nand UO_1816 (O_1816,N_18782,N_18245);
nor UO_1817 (O_1817,N_19737,N_16303);
nor UO_1818 (O_1818,N_19542,N_17399);
and UO_1819 (O_1819,N_16570,N_17502);
or UO_1820 (O_1820,N_16108,N_19480);
nor UO_1821 (O_1821,N_17322,N_18621);
and UO_1822 (O_1822,N_16497,N_16615);
nor UO_1823 (O_1823,N_19640,N_18617);
or UO_1824 (O_1824,N_17534,N_16276);
nor UO_1825 (O_1825,N_18674,N_19585);
or UO_1826 (O_1826,N_16418,N_18771);
and UO_1827 (O_1827,N_16729,N_16989);
nor UO_1828 (O_1828,N_16333,N_16140);
and UO_1829 (O_1829,N_17072,N_19561);
and UO_1830 (O_1830,N_17895,N_18502);
nand UO_1831 (O_1831,N_16820,N_17742);
and UO_1832 (O_1832,N_16053,N_17114);
nand UO_1833 (O_1833,N_16684,N_19635);
nand UO_1834 (O_1834,N_18732,N_19121);
nor UO_1835 (O_1835,N_18315,N_16724);
nand UO_1836 (O_1836,N_18672,N_17643);
or UO_1837 (O_1837,N_17149,N_17889);
xor UO_1838 (O_1838,N_17266,N_18032);
nand UO_1839 (O_1839,N_16028,N_18321);
nand UO_1840 (O_1840,N_18273,N_19176);
and UO_1841 (O_1841,N_16492,N_18667);
nor UO_1842 (O_1842,N_19406,N_19101);
nor UO_1843 (O_1843,N_18772,N_18988);
nor UO_1844 (O_1844,N_17333,N_16175);
and UO_1845 (O_1845,N_16668,N_16226);
and UO_1846 (O_1846,N_17208,N_18590);
and UO_1847 (O_1847,N_16920,N_18673);
nor UO_1848 (O_1848,N_18512,N_19308);
nand UO_1849 (O_1849,N_19161,N_19578);
and UO_1850 (O_1850,N_16341,N_18904);
nand UO_1851 (O_1851,N_18123,N_16321);
nand UO_1852 (O_1852,N_18589,N_17437);
or UO_1853 (O_1853,N_19765,N_19128);
xnor UO_1854 (O_1854,N_19425,N_18920);
and UO_1855 (O_1855,N_16449,N_18818);
xor UO_1856 (O_1856,N_17191,N_17362);
or UO_1857 (O_1857,N_16784,N_17418);
nor UO_1858 (O_1858,N_16131,N_18806);
and UO_1859 (O_1859,N_18799,N_18441);
nor UO_1860 (O_1860,N_17057,N_18661);
and UO_1861 (O_1861,N_17176,N_16034);
xor UO_1862 (O_1862,N_18147,N_18507);
xnor UO_1863 (O_1863,N_17943,N_19793);
or UO_1864 (O_1864,N_18113,N_16063);
nor UO_1865 (O_1865,N_18606,N_19198);
xnor UO_1866 (O_1866,N_19276,N_17605);
xnor UO_1867 (O_1867,N_19701,N_18718);
nor UO_1868 (O_1868,N_16706,N_19586);
and UO_1869 (O_1869,N_17095,N_19522);
or UO_1870 (O_1870,N_17800,N_19240);
or UO_1871 (O_1871,N_18850,N_16477);
nand UO_1872 (O_1872,N_19850,N_19886);
or UO_1873 (O_1873,N_16883,N_16040);
and UO_1874 (O_1874,N_18005,N_16146);
nor UO_1875 (O_1875,N_18088,N_19575);
nand UO_1876 (O_1876,N_19872,N_19930);
xnor UO_1877 (O_1877,N_16441,N_19971);
nand UO_1878 (O_1878,N_16812,N_17097);
or UO_1879 (O_1879,N_17852,N_16017);
or UO_1880 (O_1880,N_18758,N_19476);
nand UO_1881 (O_1881,N_18948,N_18967);
and UO_1882 (O_1882,N_17058,N_19621);
nor UO_1883 (O_1883,N_18751,N_18417);
xor UO_1884 (O_1884,N_16985,N_16689);
and UO_1885 (O_1885,N_18866,N_18035);
xnor UO_1886 (O_1886,N_16018,N_16194);
nor UO_1887 (O_1887,N_17933,N_17152);
and UO_1888 (O_1888,N_17425,N_18791);
nand UO_1889 (O_1889,N_19125,N_17404);
and UO_1890 (O_1890,N_18473,N_18574);
or UO_1891 (O_1891,N_17790,N_18358);
and UO_1892 (O_1892,N_19638,N_17497);
xnor UO_1893 (O_1893,N_17192,N_17245);
xor UO_1894 (O_1894,N_19704,N_16215);
nor UO_1895 (O_1895,N_19033,N_16716);
nand UO_1896 (O_1896,N_19088,N_19654);
and UO_1897 (O_1897,N_18874,N_19983);
nand UO_1898 (O_1898,N_16234,N_19348);
nor UO_1899 (O_1899,N_19636,N_19144);
nor UO_1900 (O_1900,N_17784,N_17415);
and UO_1901 (O_1901,N_18260,N_18308);
nand UO_1902 (O_1902,N_18549,N_16252);
nor UO_1903 (O_1903,N_19070,N_16310);
nor UO_1904 (O_1904,N_19212,N_16887);
nor UO_1905 (O_1905,N_17386,N_19804);
xnor UO_1906 (O_1906,N_19946,N_19028);
xor UO_1907 (O_1907,N_16510,N_18079);
or UO_1908 (O_1908,N_16526,N_17091);
nor UO_1909 (O_1909,N_19228,N_19797);
nor UO_1910 (O_1910,N_18426,N_18853);
xnor UO_1911 (O_1911,N_18314,N_17653);
nor UO_1912 (O_1912,N_17181,N_19167);
nor UO_1913 (O_1913,N_19150,N_17825);
and UO_1914 (O_1914,N_16061,N_17196);
nand UO_1915 (O_1915,N_16595,N_17310);
nand UO_1916 (O_1916,N_17658,N_16254);
and UO_1917 (O_1917,N_19148,N_17954);
xnor UO_1918 (O_1918,N_18165,N_16877);
or UO_1919 (O_1919,N_19710,N_16347);
xnor UO_1920 (O_1920,N_18277,N_18176);
nor UO_1921 (O_1921,N_19885,N_18169);
and UO_1922 (O_1922,N_19927,N_19663);
xnor UO_1923 (O_1923,N_18459,N_17381);
and UO_1924 (O_1924,N_17793,N_18898);
xnor UO_1925 (O_1925,N_18884,N_19631);
and UO_1926 (O_1926,N_18377,N_17102);
and UO_1927 (O_1927,N_18648,N_18737);
nand UO_1928 (O_1928,N_18458,N_18096);
xor UO_1929 (O_1929,N_16446,N_17324);
nor UO_1930 (O_1930,N_16975,N_17384);
and UO_1931 (O_1931,N_17481,N_16759);
xor UO_1932 (O_1932,N_19931,N_16196);
nand UO_1933 (O_1933,N_18373,N_19772);
nand UO_1934 (O_1934,N_17289,N_18057);
nor UO_1935 (O_1935,N_16319,N_17619);
nor UO_1936 (O_1936,N_17438,N_17126);
nand UO_1937 (O_1937,N_18346,N_19936);
or UO_1938 (O_1938,N_16068,N_19186);
xor UO_1939 (O_1939,N_19157,N_17623);
xor UO_1940 (O_1940,N_19584,N_16939);
nor UO_1941 (O_1941,N_19792,N_16790);
nand UO_1942 (O_1942,N_18730,N_16399);
or UO_1943 (O_1943,N_17090,N_19259);
nand UO_1944 (O_1944,N_17185,N_16271);
and UO_1945 (O_1945,N_19163,N_17764);
nand UO_1946 (O_1946,N_18689,N_16926);
or UO_1947 (O_1947,N_19274,N_18070);
nand UO_1948 (O_1948,N_17453,N_16527);
nand UO_1949 (O_1949,N_16623,N_17277);
xor UO_1950 (O_1950,N_18505,N_18348);
or UO_1951 (O_1951,N_16834,N_17817);
xnor UO_1952 (O_1952,N_16026,N_18844);
or UO_1953 (O_1953,N_19288,N_17433);
and UO_1954 (O_1954,N_17387,N_16556);
nor UO_1955 (O_1955,N_19379,N_17979);
or UO_1956 (O_1956,N_16664,N_19713);
nand UO_1957 (O_1957,N_18135,N_19758);
and UO_1958 (O_1958,N_17337,N_17491);
nor UO_1959 (O_1959,N_17796,N_17080);
nor UO_1960 (O_1960,N_19848,N_19378);
or UO_1961 (O_1961,N_19738,N_19973);
nor UO_1962 (O_1962,N_17843,N_19127);
xnor UO_1963 (O_1963,N_18959,N_19299);
nor UO_1964 (O_1964,N_19760,N_16072);
nor UO_1965 (O_1965,N_17110,N_16242);
nand UO_1966 (O_1966,N_17540,N_19213);
or UO_1967 (O_1967,N_18064,N_17982);
xnor UO_1968 (O_1968,N_17714,N_16519);
xor UO_1969 (O_1969,N_18533,N_16183);
nor UO_1970 (O_1970,N_16296,N_18906);
nand UO_1971 (O_1971,N_19775,N_18721);
nand UO_1972 (O_1972,N_18936,N_19733);
nor UO_1973 (O_1973,N_16167,N_19680);
nor UO_1974 (O_1974,N_18192,N_16186);
and UO_1975 (O_1975,N_16156,N_19594);
nand UO_1976 (O_1976,N_19024,N_17088);
nor UO_1977 (O_1977,N_19857,N_17407);
or UO_1978 (O_1978,N_16695,N_16339);
and UO_1979 (O_1979,N_17750,N_17831);
nand UO_1980 (O_1980,N_16658,N_18651);
nor UO_1981 (O_1981,N_19199,N_19473);
nor UO_1982 (O_1982,N_18278,N_17964);
nand UO_1983 (O_1983,N_19423,N_18145);
nor UO_1984 (O_1984,N_16125,N_16717);
xor UO_1985 (O_1985,N_17998,N_19352);
and UO_1986 (O_1986,N_18293,N_18163);
nand UO_1987 (O_1987,N_16709,N_19387);
and UO_1988 (O_1988,N_19859,N_16379);
xnor UO_1989 (O_1989,N_19139,N_19445);
nor UO_1990 (O_1990,N_16756,N_18983);
nor UO_1991 (O_1991,N_16586,N_16103);
nor UO_1992 (O_1992,N_18783,N_18110);
or UO_1993 (O_1993,N_19329,N_19658);
and UO_1994 (O_1994,N_19523,N_16894);
xnor UO_1995 (O_1995,N_18883,N_16893);
or UO_1996 (O_1996,N_17344,N_19089);
and UO_1997 (O_1997,N_19451,N_18578);
and UO_1998 (O_1998,N_16685,N_16292);
xor UO_1999 (O_1999,N_17526,N_19633);
and UO_2000 (O_2000,N_17271,N_17463);
and UO_2001 (O_2001,N_19018,N_18531);
and UO_2002 (O_2002,N_19698,N_18127);
and UO_2003 (O_2003,N_16830,N_19705);
nand UO_2004 (O_2004,N_18253,N_17212);
and UO_2005 (O_2005,N_18527,N_19967);
nand UO_2006 (O_2006,N_19707,N_16291);
nand UO_2007 (O_2007,N_16314,N_17762);
nand UO_2008 (O_2008,N_19568,N_19295);
nand UO_2009 (O_2009,N_19813,N_18277);
or UO_2010 (O_2010,N_16482,N_17519);
xor UO_2011 (O_2011,N_18387,N_18161);
xnor UO_2012 (O_2012,N_16327,N_18268);
and UO_2013 (O_2013,N_19966,N_19504);
nand UO_2014 (O_2014,N_18020,N_16110);
or UO_2015 (O_2015,N_16623,N_16552);
and UO_2016 (O_2016,N_18628,N_19337);
nor UO_2017 (O_2017,N_19771,N_17903);
nor UO_2018 (O_2018,N_18507,N_19090);
or UO_2019 (O_2019,N_16589,N_18418);
and UO_2020 (O_2020,N_16126,N_19828);
nor UO_2021 (O_2021,N_19536,N_19239);
xnor UO_2022 (O_2022,N_16706,N_17828);
or UO_2023 (O_2023,N_16642,N_17879);
xnor UO_2024 (O_2024,N_17815,N_18880);
and UO_2025 (O_2025,N_18084,N_17875);
nor UO_2026 (O_2026,N_19717,N_19530);
xnor UO_2027 (O_2027,N_19011,N_17378);
and UO_2028 (O_2028,N_17054,N_16273);
nor UO_2029 (O_2029,N_18657,N_16843);
nor UO_2030 (O_2030,N_18651,N_16784);
and UO_2031 (O_2031,N_19863,N_18230);
xor UO_2032 (O_2032,N_19607,N_18150);
xnor UO_2033 (O_2033,N_17051,N_16039);
nor UO_2034 (O_2034,N_17628,N_16664);
nand UO_2035 (O_2035,N_18747,N_17468);
xnor UO_2036 (O_2036,N_19109,N_16764);
or UO_2037 (O_2037,N_17294,N_16942);
and UO_2038 (O_2038,N_17800,N_17288);
nor UO_2039 (O_2039,N_19346,N_17335);
and UO_2040 (O_2040,N_17887,N_16325);
nand UO_2041 (O_2041,N_19231,N_16833);
nand UO_2042 (O_2042,N_17045,N_17496);
nor UO_2043 (O_2043,N_18336,N_17123);
and UO_2044 (O_2044,N_19045,N_18856);
nand UO_2045 (O_2045,N_16232,N_16078);
xnor UO_2046 (O_2046,N_18120,N_17127);
or UO_2047 (O_2047,N_18224,N_17661);
or UO_2048 (O_2048,N_16907,N_18982);
or UO_2049 (O_2049,N_19869,N_17032);
xor UO_2050 (O_2050,N_17948,N_18877);
and UO_2051 (O_2051,N_19971,N_18670);
nor UO_2052 (O_2052,N_19362,N_19522);
nand UO_2053 (O_2053,N_17116,N_17528);
or UO_2054 (O_2054,N_19851,N_19467);
nand UO_2055 (O_2055,N_18338,N_19794);
nor UO_2056 (O_2056,N_17520,N_18921);
and UO_2057 (O_2057,N_16679,N_17025);
nand UO_2058 (O_2058,N_16441,N_16832);
or UO_2059 (O_2059,N_18096,N_19978);
xor UO_2060 (O_2060,N_18278,N_16192);
nand UO_2061 (O_2061,N_18299,N_19785);
xnor UO_2062 (O_2062,N_18996,N_19294);
nand UO_2063 (O_2063,N_16449,N_18096);
nand UO_2064 (O_2064,N_19945,N_16434);
or UO_2065 (O_2065,N_18853,N_17175);
or UO_2066 (O_2066,N_19257,N_19607);
nor UO_2067 (O_2067,N_16641,N_16203);
nor UO_2068 (O_2068,N_16386,N_18217);
nor UO_2069 (O_2069,N_17615,N_16723);
and UO_2070 (O_2070,N_18752,N_16498);
xor UO_2071 (O_2071,N_16111,N_17340);
and UO_2072 (O_2072,N_19144,N_16890);
or UO_2073 (O_2073,N_16096,N_18456);
xnor UO_2074 (O_2074,N_17862,N_18865);
xnor UO_2075 (O_2075,N_18534,N_18633);
nand UO_2076 (O_2076,N_16093,N_17303);
and UO_2077 (O_2077,N_19086,N_17063);
or UO_2078 (O_2078,N_19576,N_16329);
xor UO_2079 (O_2079,N_16274,N_16139);
nor UO_2080 (O_2080,N_17261,N_17934);
xor UO_2081 (O_2081,N_16852,N_17529);
or UO_2082 (O_2082,N_19751,N_18918);
and UO_2083 (O_2083,N_19848,N_19774);
and UO_2084 (O_2084,N_16739,N_17932);
nor UO_2085 (O_2085,N_17531,N_17088);
and UO_2086 (O_2086,N_18832,N_18174);
xor UO_2087 (O_2087,N_17026,N_18527);
nand UO_2088 (O_2088,N_19290,N_16011);
or UO_2089 (O_2089,N_19993,N_17013);
nor UO_2090 (O_2090,N_16113,N_16856);
and UO_2091 (O_2091,N_17380,N_16534);
xnor UO_2092 (O_2092,N_17318,N_19741);
nand UO_2093 (O_2093,N_16703,N_19503);
nand UO_2094 (O_2094,N_19889,N_17447);
nand UO_2095 (O_2095,N_16738,N_18977);
and UO_2096 (O_2096,N_16412,N_19473);
xor UO_2097 (O_2097,N_17962,N_18223);
xor UO_2098 (O_2098,N_16579,N_17644);
and UO_2099 (O_2099,N_16156,N_16390);
xor UO_2100 (O_2100,N_17781,N_18955);
or UO_2101 (O_2101,N_18315,N_17801);
nand UO_2102 (O_2102,N_16044,N_17004);
xor UO_2103 (O_2103,N_17951,N_19700);
or UO_2104 (O_2104,N_17116,N_19722);
xnor UO_2105 (O_2105,N_17571,N_18228);
nor UO_2106 (O_2106,N_16756,N_19635);
and UO_2107 (O_2107,N_19527,N_17734);
nand UO_2108 (O_2108,N_18776,N_16700);
or UO_2109 (O_2109,N_16538,N_18810);
nor UO_2110 (O_2110,N_16289,N_19261);
xor UO_2111 (O_2111,N_18636,N_18562);
nand UO_2112 (O_2112,N_19149,N_16458);
nor UO_2113 (O_2113,N_17576,N_19360);
nand UO_2114 (O_2114,N_17115,N_17465);
nand UO_2115 (O_2115,N_19726,N_16393);
nand UO_2116 (O_2116,N_16951,N_16655);
or UO_2117 (O_2117,N_19138,N_16305);
nand UO_2118 (O_2118,N_19175,N_19044);
xnor UO_2119 (O_2119,N_19686,N_19280);
and UO_2120 (O_2120,N_17008,N_16952);
and UO_2121 (O_2121,N_17212,N_19273);
or UO_2122 (O_2122,N_18747,N_17524);
xnor UO_2123 (O_2123,N_16027,N_17278);
nor UO_2124 (O_2124,N_16445,N_17601);
nand UO_2125 (O_2125,N_19032,N_18018);
nand UO_2126 (O_2126,N_16643,N_18541);
and UO_2127 (O_2127,N_16534,N_17546);
nor UO_2128 (O_2128,N_16427,N_19564);
and UO_2129 (O_2129,N_19322,N_17104);
and UO_2130 (O_2130,N_16830,N_17530);
xnor UO_2131 (O_2131,N_18878,N_18964);
and UO_2132 (O_2132,N_18419,N_17589);
or UO_2133 (O_2133,N_16070,N_17963);
nor UO_2134 (O_2134,N_17560,N_17091);
or UO_2135 (O_2135,N_16741,N_17864);
or UO_2136 (O_2136,N_18277,N_19368);
xor UO_2137 (O_2137,N_17824,N_18712);
nand UO_2138 (O_2138,N_19844,N_19185);
xnor UO_2139 (O_2139,N_18036,N_18247);
or UO_2140 (O_2140,N_16010,N_17649);
xnor UO_2141 (O_2141,N_17815,N_17235);
and UO_2142 (O_2142,N_18596,N_18447);
or UO_2143 (O_2143,N_18561,N_18029);
nand UO_2144 (O_2144,N_16071,N_19715);
and UO_2145 (O_2145,N_17117,N_16855);
xor UO_2146 (O_2146,N_16448,N_19881);
nor UO_2147 (O_2147,N_19521,N_16340);
and UO_2148 (O_2148,N_18838,N_17112);
nor UO_2149 (O_2149,N_16697,N_19774);
xor UO_2150 (O_2150,N_19157,N_16619);
nand UO_2151 (O_2151,N_17980,N_19977);
xnor UO_2152 (O_2152,N_19052,N_19293);
or UO_2153 (O_2153,N_17331,N_18809);
nor UO_2154 (O_2154,N_17591,N_17330);
xnor UO_2155 (O_2155,N_19567,N_19925);
nor UO_2156 (O_2156,N_17665,N_17654);
nor UO_2157 (O_2157,N_16575,N_16135);
and UO_2158 (O_2158,N_19228,N_16608);
xor UO_2159 (O_2159,N_17344,N_19374);
or UO_2160 (O_2160,N_19701,N_16198);
and UO_2161 (O_2161,N_16123,N_18452);
nand UO_2162 (O_2162,N_17693,N_17601);
xor UO_2163 (O_2163,N_16432,N_17896);
nand UO_2164 (O_2164,N_19655,N_17864);
and UO_2165 (O_2165,N_16615,N_16039);
and UO_2166 (O_2166,N_16586,N_18336);
or UO_2167 (O_2167,N_19861,N_17862);
nor UO_2168 (O_2168,N_16380,N_17000);
nand UO_2169 (O_2169,N_18877,N_18611);
and UO_2170 (O_2170,N_16942,N_18943);
xor UO_2171 (O_2171,N_18105,N_18155);
xor UO_2172 (O_2172,N_16259,N_19132);
and UO_2173 (O_2173,N_19958,N_17601);
xor UO_2174 (O_2174,N_16595,N_16430);
or UO_2175 (O_2175,N_18653,N_18368);
xnor UO_2176 (O_2176,N_19969,N_16048);
xnor UO_2177 (O_2177,N_19370,N_19789);
and UO_2178 (O_2178,N_16548,N_18007);
or UO_2179 (O_2179,N_18625,N_16581);
xor UO_2180 (O_2180,N_18988,N_19766);
or UO_2181 (O_2181,N_18344,N_17560);
xnor UO_2182 (O_2182,N_17017,N_16689);
nor UO_2183 (O_2183,N_19782,N_18142);
nor UO_2184 (O_2184,N_17273,N_19422);
nand UO_2185 (O_2185,N_19150,N_18424);
nor UO_2186 (O_2186,N_18041,N_18951);
nand UO_2187 (O_2187,N_19588,N_16264);
nand UO_2188 (O_2188,N_16725,N_18753);
nor UO_2189 (O_2189,N_17689,N_17046);
nor UO_2190 (O_2190,N_17443,N_18040);
xor UO_2191 (O_2191,N_16238,N_16388);
or UO_2192 (O_2192,N_18648,N_18255);
nand UO_2193 (O_2193,N_16549,N_18961);
nand UO_2194 (O_2194,N_18218,N_16702);
nor UO_2195 (O_2195,N_18505,N_19232);
nand UO_2196 (O_2196,N_16220,N_16249);
or UO_2197 (O_2197,N_16709,N_19276);
xor UO_2198 (O_2198,N_16231,N_16649);
xnor UO_2199 (O_2199,N_18177,N_19691);
nor UO_2200 (O_2200,N_19370,N_18152);
and UO_2201 (O_2201,N_18172,N_16723);
nor UO_2202 (O_2202,N_17744,N_19027);
xor UO_2203 (O_2203,N_18188,N_19414);
xnor UO_2204 (O_2204,N_18443,N_19082);
or UO_2205 (O_2205,N_18097,N_19556);
and UO_2206 (O_2206,N_18664,N_16162);
nand UO_2207 (O_2207,N_16876,N_17355);
nor UO_2208 (O_2208,N_16715,N_19853);
nand UO_2209 (O_2209,N_17386,N_18199);
nor UO_2210 (O_2210,N_19120,N_18746);
and UO_2211 (O_2211,N_16757,N_16280);
nand UO_2212 (O_2212,N_17209,N_18357);
nand UO_2213 (O_2213,N_18716,N_17727);
xnor UO_2214 (O_2214,N_17151,N_19163);
xor UO_2215 (O_2215,N_17143,N_19321);
nor UO_2216 (O_2216,N_16179,N_17010);
and UO_2217 (O_2217,N_16707,N_17963);
xnor UO_2218 (O_2218,N_19287,N_19579);
nor UO_2219 (O_2219,N_18511,N_16516);
nor UO_2220 (O_2220,N_17630,N_16864);
nor UO_2221 (O_2221,N_16530,N_19640);
and UO_2222 (O_2222,N_18408,N_17227);
and UO_2223 (O_2223,N_19371,N_16772);
xor UO_2224 (O_2224,N_16124,N_16352);
nand UO_2225 (O_2225,N_16683,N_17428);
nand UO_2226 (O_2226,N_17092,N_19437);
xor UO_2227 (O_2227,N_19129,N_19551);
or UO_2228 (O_2228,N_18276,N_17183);
and UO_2229 (O_2229,N_17915,N_18753);
and UO_2230 (O_2230,N_16175,N_18478);
xnor UO_2231 (O_2231,N_18669,N_19266);
or UO_2232 (O_2232,N_19872,N_16023);
nor UO_2233 (O_2233,N_18661,N_19636);
and UO_2234 (O_2234,N_17242,N_18311);
xor UO_2235 (O_2235,N_19294,N_18072);
nor UO_2236 (O_2236,N_18701,N_19654);
nand UO_2237 (O_2237,N_18121,N_18410);
xor UO_2238 (O_2238,N_16663,N_18955);
or UO_2239 (O_2239,N_16012,N_19547);
nor UO_2240 (O_2240,N_19583,N_16188);
nand UO_2241 (O_2241,N_17971,N_19531);
and UO_2242 (O_2242,N_17911,N_16105);
xor UO_2243 (O_2243,N_16165,N_17562);
nor UO_2244 (O_2244,N_17865,N_17984);
nand UO_2245 (O_2245,N_18321,N_19371);
or UO_2246 (O_2246,N_17058,N_18830);
xnor UO_2247 (O_2247,N_19151,N_18153);
or UO_2248 (O_2248,N_19538,N_18707);
and UO_2249 (O_2249,N_16609,N_16263);
nand UO_2250 (O_2250,N_17015,N_19293);
nor UO_2251 (O_2251,N_16064,N_16067);
nand UO_2252 (O_2252,N_19666,N_18526);
or UO_2253 (O_2253,N_17561,N_19237);
or UO_2254 (O_2254,N_18765,N_17470);
and UO_2255 (O_2255,N_17376,N_16417);
and UO_2256 (O_2256,N_16178,N_19969);
nand UO_2257 (O_2257,N_19669,N_16344);
xor UO_2258 (O_2258,N_19343,N_18160);
or UO_2259 (O_2259,N_19516,N_19397);
nand UO_2260 (O_2260,N_16022,N_16448);
nor UO_2261 (O_2261,N_17802,N_16543);
or UO_2262 (O_2262,N_16156,N_19836);
nand UO_2263 (O_2263,N_18418,N_16965);
nor UO_2264 (O_2264,N_18286,N_17589);
xnor UO_2265 (O_2265,N_16869,N_17508);
nor UO_2266 (O_2266,N_18693,N_17251);
and UO_2267 (O_2267,N_19543,N_19551);
or UO_2268 (O_2268,N_18494,N_18617);
and UO_2269 (O_2269,N_17271,N_17426);
xnor UO_2270 (O_2270,N_16263,N_18202);
xnor UO_2271 (O_2271,N_19693,N_18266);
and UO_2272 (O_2272,N_19596,N_17698);
and UO_2273 (O_2273,N_16939,N_17226);
nand UO_2274 (O_2274,N_18495,N_18251);
or UO_2275 (O_2275,N_18595,N_17271);
and UO_2276 (O_2276,N_19742,N_17809);
nor UO_2277 (O_2277,N_17563,N_18889);
xnor UO_2278 (O_2278,N_16672,N_18882);
and UO_2279 (O_2279,N_19943,N_18986);
or UO_2280 (O_2280,N_16842,N_17799);
nor UO_2281 (O_2281,N_18676,N_17053);
and UO_2282 (O_2282,N_18866,N_16938);
and UO_2283 (O_2283,N_18921,N_16855);
or UO_2284 (O_2284,N_17438,N_19752);
xor UO_2285 (O_2285,N_17096,N_17276);
nand UO_2286 (O_2286,N_19515,N_18178);
and UO_2287 (O_2287,N_18408,N_17669);
and UO_2288 (O_2288,N_19444,N_18841);
nor UO_2289 (O_2289,N_16487,N_19424);
nor UO_2290 (O_2290,N_17149,N_18470);
xor UO_2291 (O_2291,N_19495,N_16135);
nand UO_2292 (O_2292,N_19733,N_19872);
nor UO_2293 (O_2293,N_16265,N_19325);
nor UO_2294 (O_2294,N_17285,N_19324);
nand UO_2295 (O_2295,N_17919,N_19684);
nor UO_2296 (O_2296,N_19830,N_19083);
xnor UO_2297 (O_2297,N_16411,N_16284);
or UO_2298 (O_2298,N_18403,N_17386);
or UO_2299 (O_2299,N_19341,N_16419);
and UO_2300 (O_2300,N_19785,N_16809);
or UO_2301 (O_2301,N_19627,N_18765);
and UO_2302 (O_2302,N_16846,N_19773);
nor UO_2303 (O_2303,N_18403,N_17134);
nor UO_2304 (O_2304,N_16632,N_18950);
or UO_2305 (O_2305,N_16491,N_17985);
nor UO_2306 (O_2306,N_18285,N_16009);
nand UO_2307 (O_2307,N_16039,N_17956);
and UO_2308 (O_2308,N_16886,N_19414);
and UO_2309 (O_2309,N_16955,N_17711);
nand UO_2310 (O_2310,N_19610,N_19059);
nor UO_2311 (O_2311,N_18895,N_18822);
or UO_2312 (O_2312,N_18131,N_17106);
or UO_2313 (O_2313,N_16165,N_16382);
and UO_2314 (O_2314,N_18127,N_16338);
or UO_2315 (O_2315,N_17923,N_18065);
or UO_2316 (O_2316,N_17799,N_17372);
xor UO_2317 (O_2317,N_16694,N_17149);
nand UO_2318 (O_2318,N_17750,N_19919);
xnor UO_2319 (O_2319,N_17271,N_18856);
nor UO_2320 (O_2320,N_18963,N_16638);
xor UO_2321 (O_2321,N_16665,N_16439);
nor UO_2322 (O_2322,N_16126,N_19781);
or UO_2323 (O_2323,N_19169,N_19375);
xor UO_2324 (O_2324,N_19527,N_19113);
nand UO_2325 (O_2325,N_18452,N_16116);
xor UO_2326 (O_2326,N_18547,N_16781);
nor UO_2327 (O_2327,N_19186,N_16187);
xnor UO_2328 (O_2328,N_16847,N_17081);
nor UO_2329 (O_2329,N_16780,N_19963);
or UO_2330 (O_2330,N_16547,N_17999);
nor UO_2331 (O_2331,N_19521,N_19177);
nor UO_2332 (O_2332,N_18555,N_19771);
nor UO_2333 (O_2333,N_19525,N_16947);
nor UO_2334 (O_2334,N_17346,N_18100);
and UO_2335 (O_2335,N_16091,N_17523);
nor UO_2336 (O_2336,N_18741,N_16320);
nand UO_2337 (O_2337,N_18569,N_18438);
nor UO_2338 (O_2338,N_18782,N_19596);
nor UO_2339 (O_2339,N_18341,N_16879);
or UO_2340 (O_2340,N_16895,N_19316);
and UO_2341 (O_2341,N_16180,N_17386);
nand UO_2342 (O_2342,N_16929,N_19174);
nand UO_2343 (O_2343,N_18079,N_19263);
xor UO_2344 (O_2344,N_17018,N_19783);
nand UO_2345 (O_2345,N_19531,N_18076);
nor UO_2346 (O_2346,N_17305,N_17272);
nand UO_2347 (O_2347,N_19651,N_19729);
or UO_2348 (O_2348,N_19822,N_19591);
nand UO_2349 (O_2349,N_18455,N_16344);
and UO_2350 (O_2350,N_18061,N_18140);
and UO_2351 (O_2351,N_17141,N_17396);
nor UO_2352 (O_2352,N_17140,N_17672);
or UO_2353 (O_2353,N_17046,N_19973);
xor UO_2354 (O_2354,N_19766,N_17290);
and UO_2355 (O_2355,N_16278,N_17179);
nor UO_2356 (O_2356,N_16986,N_19799);
nand UO_2357 (O_2357,N_18712,N_19853);
or UO_2358 (O_2358,N_18746,N_17722);
nand UO_2359 (O_2359,N_19704,N_17427);
or UO_2360 (O_2360,N_17657,N_16330);
or UO_2361 (O_2361,N_18828,N_18991);
nand UO_2362 (O_2362,N_19491,N_19603);
nor UO_2363 (O_2363,N_18013,N_16240);
nand UO_2364 (O_2364,N_18026,N_18428);
nor UO_2365 (O_2365,N_16358,N_18079);
and UO_2366 (O_2366,N_16819,N_18544);
nor UO_2367 (O_2367,N_18036,N_18655);
xnor UO_2368 (O_2368,N_18908,N_18712);
or UO_2369 (O_2369,N_17895,N_16156);
nand UO_2370 (O_2370,N_18844,N_18560);
nand UO_2371 (O_2371,N_19772,N_18133);
xor UO_2372 (O_2372,N_17031,N_16488);
xor UO_2373 (O_2373,N_17564,N_18457);
or UO_2374 (O_2374,N_17129,N_19826);
nor UO_2375 (O_2375,N_19157,N_18360);
and UO_2376 (O_2376,N_18525,N_19486);
and UO_2377 (O_2377,N_17870,N_17705);
nand UO_2378 (O_2378,N_16543,N_19514);
and UO_2379 (O_2379,N_18568,N_16061);
or UO_2380 (O_2380,N_18765,N_16015);
and UO_2381 (O_2381,N_16742,N_18191);
xor UO_2382 (O_2382,N_19031,N_16736);
and UO_2383 (O_2383,N_16913,N_18580);
and UO_2384 (O_2384,N_16772,N_19137);
and UO_2385 (O_2385,N_16602,N_16737);
nor UO_2386 (O_2386,N_19480,N_17021);
xor UO_2387 (O_2387,N_16381,N_16779);
nand UO_2388 (O_2388,N_18172,N_18710);
or UO_2389 (O_2389,N_19141,N_19090);
and UO_2390 (O_2390,N_18192,N_19909);
or UO_2391 (O_2391,N_16586,N_19216);
nand UO_2392 (O_2392,N_16829,N_17487);
xor UO_2393 (O_2393,N_18349,N_19444);
and UO_2394 (O_2394,N_18283,N_16171);
and UO_2395 (O_2395,N_18737,N_16555);
nand UO_2396 (O_2396,N_19424,N_19856);
xnor UO_2397 (O_2397,N_18599,N_17827);
and UO_2398 (O_2398,N_19547,N_18373);
xnor UO_2399 (O_2399,N_17252,N_19427);
nand UO_2400 (O_2400,N_19101,N_18140);
or UO_2401 (O_2401,N_17535,N_17401);
and UO_2402 (O_2402,N_18750,N_17594);
nand UO_2403 (O_2403,N_18443,N_16460);
xnor UO_2404 (O_2404,N_18578,N_16131);
or UO_2405 (O_2405,N_16442,N_16803);
nand UO_2406 (O_2406,N_16775,N_16085);
nor UO_2407 (O_2407,N_18848,N_16193);
nor UO_2408 (O_2408,N_18365,N_18875);
xor UO_2409 (O_2409,N_16640,N_18931);
nand UO_2410 (O_2410,N_18828,N_19282);
or UO_2411 (O_2411,N_19192,N_17349);
nand UO_2412 (O_2412,N_18735,N_19465);
or UO_2413 (O_2413,N_19746,N_18606);
or UO_2414 (O_2414,N_18284,N_18163);
and UO_2415 (O_2415,N_19824,N_16950);
nor UO_2416 (O_2416,N_16624,N_18629);
xor UO_2417 (O_2417,N_18661,N_16219);
and UO_2418 (O_2418,N_17116,N_18980);
or UO_2419 (O_2419,N_17029,N_18494);
xor UO_2420 (O_2420,N_18938,N_17158);
xnor UO_2421 (O_2421,N_19361,N_18097);
nand UO_2422 (O_2422,N_18841,N_19824);
or UO_2423 (O_2423,N_17834,N_17423);
nor UO_2424 (O_2424,N_18339,N_19233);
nor UO_2425 (O_2425,N_18599,N_16932);
nor UO_2426 (O_2426,N_18999,N_17024);
xnor UO_2427 (O_2427,N_19310,N_17988);
nand UO_2428 (O_2428,N_17327,N_19065);
or UO_2429 (O_2429,N_19215,N_19004);
and UO_2430 (O_2430,N_17081,N_18618);
or UO_2431 (O_2431,N_16808,N_19359);
or UO_2432 (O_2432,N_19168,N_18584);
nor UO_2433 (O_2433,N_16454,N_18911);
or UO_2434 (O_2434,N_16493,N_19698);
nand UO_2435 (O_2435,N_18523,N_18812);
and UO_2436 (O_2436,N_16879,N_19773);
and UO_2437 (O_2437,N_16056,N_16130);
nand UO_2438 (O_2438,N_19666,N_16154);
or UO_2439 (O_2439,N_17144,N_18617);
xnor UO_2440 (O_2440,N_16587,N_16966);
nand UO_2441 (O_2441,N_18095,N_19351);
nor UO_2442 (O_2442,N_17399,N_16399);
or UO_2443 (O_2443,N_16819,N_17426);
nor UO_2444 (O_2444,N_17032,N_19403);
xor UO_2445 (O_2445,N_19189,N_18070);
xnor UO_2446 (O_2446,N_19330,N_19246);
xnor UO_2447 (O_2447,N_17930,N_17695);
nor UO_2448 (O_2448,N_18563,N_17157);
or UO_2449 (O_2449,N_16505,N_18988);
and UO_2450 (O_2450,N_16615,N_16843);
or UO_2451 (O_2451,N_17382,N_19342);
xnor UO_2452 (O_2452,N_17067,N_17815);
and UO_2453 (O_2453,N_19146,N_16106);
xor UO_2454 (O_2454,N_17093,N_17849);
nor UO_2455 (O_2455,N_18388,N_16286);
xnor UO_2456 (O_2456,N_19635,N_17138);
or UO_2457 (O_2457,N_19016,N_17623);
nor UO_2458 (O_2458,N_19164,N_18776);
nor UO_2459 (O_2459,N_19000,N_18785);
xor UO_2460 (O_2460,N_16456,N_16002);
nor UO_2461 (O_2461,N_17935,N_16925);
or UO_2462 (O_2462,N_16611,N_19886);
nand UO_2463 (O_2463,N_17623,N_18260);
or UO_2464 (O_2464,N_18599,N_17395);
xnor UO_2465 (O_2465,N_19526,N_18194);
nor UO_2466 (O_2466,N_19169,N_16142);
xor UO_2467 (O_2467,N_17474,N_19221);
nor UO_2468 (O_2468,N_18071,N_18953);
and UO_2469 (O_2469,N_18855,N_18131);
xnor UO_2470 (O_2470,N_16383,N_17489);
and UO_2471 (O_2471,N_18571,N_18779);
or UO_2472 (O_2472,N_18106,N_18713);
and UO_2473 (O_2473,N_19497,N_16269);
nor UO_2474 (O_2474,N_19505,N_16112);
nor UO_2475 (O_2475,N_17769,N_19070);
nor UO_2476 (O_2476,N_16361,N_16060);
and UO_2477 (O_2477,N_19514,N_18415);
nand UO_2478 (O_2478,N_17953,N_17413);
or UO_2479 (O_2479,N_16801,N_19148);
and UO_2480 (O_2480,N_18026,N_17425);
and UO_2481 (O_2481,N_17524,N_17714);
or UO_2482 (O_2482,N_19283,N_17477);
or UO_2483 (O_2483,N_19980,N_16071);
nand UO_2484 (O_2484,N_17913,N_18988);
xnor UO_2485 (O_2485,N_16912,N_16037);
nand UO_2486 (O_2486,N_17190,N_18867);
and UO_2487 (O_2487,N_16118,N_17088);
xnor UO_2488 (O_2488,N_17576,N_17836);
xor UO_2489 (O_2489,N_17891,N_16032);
nor UO_2490 (O_2490,N_19679,N_18723);
or UO_2491 (O_2491,N_16553,N_16557);
xor UO_2492 (O_2492,N_19339,N_16022);
or UO_2493 (O_2493,N_19803,N_17125);
or UO_2494 (O_2494,N_17894,N_18995);
nand UO_2495 (O_2495,N_18605,N_18742);
and UO_2496 (O_2496,N_17655,N_18577);
xnor UO_2497 (O_2497,N_19452,N_18089);
or UO_2498 (O_2498,N_17959,N_17518);
or UO_2499 (O_2499,N_18234,N_17234);
endmodule