module basic_1500_15000_2000_60_levels_5xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
xor U0 (N_0,In_532,In_101);
nor U1 (N_1,In_607,In_1011);
nor U2 (N_2,In_522,In_370);
or U3 (N_3,In_1410,In_476);
and U4 (N_4,In_9,In_1302);
nand U5 (N_5,In_499,In_821);
xor U6 (N_6,In_356,In_599);
nand U7 (N_7,In_295,In_791);
or U8 (N_8,In_7,In_335);
xor U9 (N_9,In_741,In_94);
and U10 (N_10,In_763,In_865);
nand U11 (N_11,In_41,In_1223);
nor U12 (N_12,In_758,In_1133);
or U13 (N_13,In_1009,In_1010);
nand U14 (N_14,In_1016,In_606);
and U15 (N_15,In_185,In_677);
and U16 (N_16,In_942,In_1353);
and U17 (N_17,In_771,In_627);
nor U18 (N_18,In_266,In_750);
nand U19 (N_19,In_330,In_353);
xor U20 (N_20,In_51,In_1293);
and U21 (N_21,In_938,In_176);
nor U22 (N_22,In_565,In_1460);
nand U23 (N_23,In_731,In_492);
xnor U24 (N_24,In_90,In_1144);
and U25 (N_25,In_40,In_316);
or U26 (N_26,In_1207,In_389);
and U27 (N_27,In_275,In_911);
or U28 (N_28,In_1475,In_475);
xor U29 (N_29,In_31,In_318);
or U30 (N_30,In_177,In_551);
and U31 (N_31,In_1152,In_1156);
nor U32 (N_32,In_840,In_1147);
nor U33 (N_33,In_50,In_996);
or U34 (N_34,In_161,In_935);
xor U35 (N_35,In_1192,In_1168);
or U36 (N_36,In_766,In_1245);
nor U37 (N_37,In_450,In_512);
xor U38 (N_38,In_16,In_500);
nor U39 (N_39,In_716,In_798);
and U40 (N_40,In_1237,In_901);
or U41 (N_41,In_296,In_1306);
nand U42 (N_42,In_703,In_1195);
and U43 (N_43,In_253,In_976);
and U44 (N_44,In_718,In_642);
nand U45 (N_45,In_1014,In_579);
and U46 (N_46,In_320,In_645);
or U47 (N_47,In_472,In_454);
nor U48 (N_48,In_1116,In_993);
or U49 (N_49,In_625,In_1413);
nand U50 (N_50,In_770,In_644);
nand U51 (N_51,In_156,In_270);
and U52 (N_52,In_534,In_464);
or U53 (N_53,In_560,In_1139);
nor U54 (N_54,In_1498,In_847);
and U55 (N_55,In_1231,In_406);
xnor U56 (N_56,In_381,In_197);
nand U57 (N_57,In_635,In_785);
and U58 (N_58,In_822,In_224);
nor U59 (N_59,In_649,In_819);
or U60 (N_60,In_113,In_291);
nand U61 (N_61,In_285,In_234);
nor U62 (N_62,In_1338,In_251);
nor U63 (N_63,In_337,In_1472);
or U64 (N_64,In_844,In_1111);
nor U65 (N_65,In_1126,In_636);
or U66 (N_66,In_114,In_870);
and U67 (N_67,In_298,In_1070);
or U68 (N_68,In_547,In_45);
nand U69 (N_69,In_1027,In_1076);
nand U70 (N_70,In_1469,In_1436);
xor U71 (N_71,In_792,In_1154);
nor U72 (N_72,In_1159,In_1491);
nand U73 (N_73,In_67,In_116);
nand U74 (N_74,In_438,In_546);
nand U75 (N_75,In_1290,In_1361);
nand U76 (N_76,In_658,In_1467);
nor U77 (N_77,In_1319,In_46);
nand U78 (N_78,In_1104,In_172);
nand U79 (N_79,In_1142,In_962);
nor U80 (N_80,In_768,In_199);
and U81 (N_81,In_308,In_539);
nor U82 (N_82,In_437,In_524);
nor U83 (N_83,In_707,In_66);
and U84 (N_84,In_1103,In_1050);
and U85 (N_85,In_1158,In_783);
and U86 (N_86,In_687,In_478);
and U87 (N_87,In_1176,In_1360);
nand U88 (N_88,In_1217,In_417);
xnor U89 (N_89,In_1199,In_98);
or U90 (N_90,In_991,In_926);
and U91 (N_91,In_32,In_773);
or U92 (N_92,In_214,In_357);
and U93 (N_93,In_733,In_1257);
nand U94 (N_94,In_132,In_812);
and U95 (N_95,In_1375,In_659);
and U96 (N_96,In_252,In_30);
xnor U97 (N_97,In_691,In_588);
and U98 (N_98,In_611,In_860);
nand U99 (N_99,In_1214,In_1187);
nor U100 (N_100,In_520,In_340);
nand U101 (N_101,In_1004,In_1330);
and U102 (N_102,In_927,In_790);
xnor U103 (N_103,In_853,In_401);
and U104 (N_104,In_299,In_1119);
nand U105 (N_105,In_441,In_345);
or U106 (N_106,In_1053,In_838);
and U107 (N_107,In_630,In_324);
nor U108 (N_108,In_972,In_1327);
nor U109 (N_109,In_1239,In_100);
or U110 (N_110,In_1412,In_816);
xor U111 (N_111,In_1107,In_728);
nor U112 (N_112,In_1493,In_1040);
nor U113 (N_113,In_1459,In_958);
and U114 (N_114,In_1274,In_1387);
nand U115 (N_115,In_814,In_681);
nand U116 (N_116,In_313,In_1457);
nor U117 (N_117,In_535,In_894);
nand U118 (N_118,In_1454,In_196);
and U119 (N_119,In_1465,In_79);
nor U120 (N_120,In_756,In_1072);
xnor U121 (N_121,In_457,In_694);
nor U122 (N_122,In_1186,In_754);
nor U123 (N_123,In_173,In_829);
or U124 (N_124,In_143,In_980);
nor U125 (N_125,In_123,In_257);
nand U126 (N_126,In_1316,In_1197);
nor U127 (N_127,In_474,In_28);
nor U128 (N_128,In_1440,In_1099);
and U129 (N_129,In_1148,In_201);
or U130 (N_130,In_88,In_307);
and U131 (N_131,In_1028,In_297);
nand U132 (N_132,In_777,In_76);
nor U133 (N_133,In_559,In_1419);
and U134 (N_134,In_724,In_775);
and U135 (N_135,In_1025,In_1437);
nor U136 (N_136,In_1259,In_1249);
and U137 (N_137,In_426,In_1313);
nand U138 (N_138,In_761,In_831);
nand U139 (N_139,In_1458,In_633);
or U140 (N_140,In_1281,In_1370);
nand U141 (N_141,In_405,In_698);
or U142 (N_142,In_710,In_797);
and U143 (N_143,In_315,In_849);
nand U144 (N_144,In_973,In_498);
xor U145 (N_145,In_13,In_84);
or U146 (N_146,In_1446,In_1059);
and U147 (N_147,In_1426,In_1150);
nor U148 (N_148,In_566,In_1321);
or U149 (N_149,In_1496,In_1096);
nand U150 (N_150,In_47,In_10);
and U151 (N_151,In_517,In_671);
or U152 (N_152,In_455,In_637);
nand U153 (N_153,In_704,In_1389);
nor U154 (N_154,In_1391,In_378);
nand U155 (N_155,In_826,In_1211);
and U156 (N_156,In_19,In_836);
or U157 (N_157,In_825,In_1282);
or U158 (N_158,In_834,In_892);
or U159 (N_159,In_24,In_1265);
or U160 (N_160,In_530,In_721);
or U161 (N_161,In_227,In_105);
nand U162 (N_162,In_815,In_941);
nand U163 (N_163,In_439,In_1435);
nand U164 (N_164,In_1057,In_1242);
or U165 (N_165,In_321,In_646);
and U166 (N_166,In_1205,In_1487);
and U167 (N_167,In_1155,In_923);
nand U168 (N_168,In_1185,In_471);
and U169 (N_169,In_384,In_909);
nor U170 (N_170,In_1171,In_578);
nor U171 (N_171,In_392,In_540);
or U172 (N_172,In_194,In_857);
and U173 (N_173,In_638,In_218);
nand U174 (N_174,In_985,In_1210);
or U175 (N_175,In_1055,In_1042);
and U176 (N_176,In_835,In_33);
nor U177 (N_177,In_1453,In_1429);
nor U178 (N_178,In_1007,In_695);
or U179 (N_179,In_582,In_626);
nand U180 (N_180,In_443,In_372);
and U181 (N_181,In_348,In_216);
xor U182 (N_182,In_1444,In_984);
xor U183 (N_183,In_130,In_709);
or U184 (N_184,In_928,In_1234);
xnor U185 (N_185,In_706,In_1203);
or U186 (N_186,In_1374,In_977);
and U187 (N_187,In_311,In_288);
nor U188 (N_188,In_1029,In_1071);
or U189 (N_189,In_1143,In_619);
nand U190 (N_190,In_1189,In_1318);
nand U191 (N_191,In_518,In_1013);
nand U192 (N_192,In_513,In_1032);
and U193 (N_193,In_869,In_1052);
or U194 (N_194,In_422,In_212);
nand U195 (N_195,In_52,In_360);
nand U196 (N_196,In_749,In_845);
nand U197 (N_197,In_1173,In_1329);
nor U198 (N_198,In_782,In_477);
and U199 (N_199,In_1235,In_1124);
nor U200 (N_200,In_715,In_887);
nand U201 (N_201,In_1178,In_598);
nor U202 (N_202,In_1082,In_423);
and U203 (N_203,In_1091,In_59);
and U204 (N_204,In_590,In_1035);
or U205 (N_205,In_364,In_1325);
and U206 (N_206,In_362,In_1320);
xor U207 (N_207,In_541,In_1431);
and U208 (N_208,In_1196,In_511);
or U209 (N_209,In_789,In_117);
nand U210 (N_210,In_466,In_469);
nand U211 (N_211,In_974,In_97);
nor U212 (N_212,In_317,In_618);
and U213 (N_213,In_289,In_239);
or U214 (N_214,In_661,In_26);
nor U215 (N_215,In_460,In_495);
nand U216 (N_216,In_602,In_1074);
or U217 (N_217,In_178,In_752);
nor U218 (N_218,In_14,In_329);
and U219 (N_219,In_886,In_519);
or U220 (N_220,In_209,In_846);
and U221 (N_221,In_413,In_391);
xor U222 (N_222,In_503,In_440);
nand U223 (N_223,In_1344,In_878);
or U224 (N_224,In_331,In_230);
and U225 (N_225,In_434,In_429);
nor U226 (N_226,In_1106,In_1191);
and U227 (N_227,In_960,In_956);
nand U228 (N_228,In_605,In_1001);
nor U229 (N_229,In_78,In_1153);
and U230 (N_230,In_122,In_15);
nor U231 (N_231,In_436,In_482);
nand U232 (N_232,In_1180,In_425);
nor U233 (N_233,In_427,In_1182);
and U234 (N_234,In_641,In_508);
nand U235 (N_235,In_501,In_1296);
and U236 (N_236,In_505,In_608);
xor U237 (N_237,In_1455,In_139);
or U238 (N_238,In_1347,In_1031);
nand U239 (N_239,In_278,In_202);
nand U240 (N_240,In_759,In_463);
nor U241 (N_241,In_62,In_86);
nand U242 (N_242,In_119,In_686);
nor U243 (N_243,In_1462,In_1289);
xor U244 (N_244,In_850,In_528);
nor U245 (N_245,In_903,In_1381);
and U246 (N_246,In_494,In_366);
or U247 (N_247,In_747,In_667);
nand U248 (N_248,In_1228,In_355);
and U249 (N_249,In_967,In_806);
xnor U250 (N_250,In_1030,In_981);
xnor U251 (N_251,In_1405,N_172);
and U252 (N_252,In_1271,In_730);
nand U253 (N_253,In_91,In_1408);
nand U254 (N_254,N_184,In_1258);
nand U255 (N_255,N_111,In_720);
xnor U256 (N_256,In_322,In_1084);
or U257 (N_257,In_1006,In_924);
nand U258 (N_258,In_964,N_114);
or U259 (N_259,In_1129,In_1273);
and U260 (N_260,In_548,In_53);
xnor U261 (N_261,In_109,In_1005);
nor U262 (N_262,In_653,In_190);
nand U263 (N_263,In_1450,N_16);
or U264 (N_264,In_1300,N_55);
nor U265 (N_265,In_1489,In_1218);
and U266 (N_266,In_688,In_930);
xor U267 (N_267,In_3,In_265);
nand U268 (N_268,N_21,In_171);
nor U269 (N_269,In_226,In_260);
nor U270 (N_270,In_553,In_371);
nor U271 (N_271,In_778,In_481);
and U272 (N_272,In_1400,In_760);
nor U273 (N_273,N_164,In_1415);
nor U274 (N_274,In_244,In_1366);
nand U275 (N_275,In_148,In_556);
nand U276 (N_276,In_134,In_660);
and U277 (N_277,In_568,In_700);
or U278 (N_278,In_1219,In_138);
or U279 (N_279,In_1089,In_533);
or U280 (N_280,In_1067,In_449);
and U281 (N_281,In_25,In_1401);
nand U282 (N_282,In_342,N_62);
nand U283 (N_283,N_189,In_1399);
and U284 (N_284,In_562,In_841);
and U285 (N_285,In_622,In_170);
xor U286 (N_286,N_162,N_141);
and U287 (N_287,In_81,In_612);
nand U288 (N_288,In_314,In_839);
xor U289 (N_289,In_49,N_70);
nand U290 (N_290,N_147,N_187);
or U291 (N_291,In_920,In_1221);
nand U292 (N_292,In_153,N_7);
and U293 (N_293,In_1065,In_1238);
or U294 (N_294,In_651,N_13);
nor U295 (N_295,In_1132,In_685);
nand U296 (N_296,In_1179,N_158);
nand U297 (N_297,In_305,In_419);
nor U298 (N_298,In_830,N_130);
or U299 (N_299,In_1108,N_245);
or U300 (N_300,N_12,In_22);
nor U301 (N_301,In_36,N_188);
or U302 (N_302,In_988,N_122);
nor U303 (N_303,In_8,In_263);
or U304 (N_304,In_430,In_420);
nor U305 (N_305,N_40,In_793);
nand U306 (N_306,In_1363,In_751);
or U307 (N_307,N_210,In_282);
nor U308 (N_308,In_280,In_369);
or U309 (N_309,N_170,In_757);
nand U310 (N_310,In_1086,In_1220);
and U311 (N_311,In_21,In_325);
or U312 (N_312,In_365,In_1247);
nor U313 (N_313,N_103,In_396);
or U314 (N_314,N_222,In_1166);
nand U315 (N_315,In_1000,In_874);
nor U316 (N_316,In_1488,In_950);
nand U317 (N_317,In_1127,In_1101);
nor U318 (N_318,In_665,In_854);
xnor U319 (N_319,In_167,In_828);
xnor U320 (N_320,In_1310,In_1463);
and U321 (N_321,In_1388,In_943);
and U322 (N_322,In_1085,In_693);
nand U323 (N_323,In_744,In_1334);
nor U324 (N_324,N_175,In_1349);
nand U325 (N_325,In_650,In_276);
nand U326 (N_326,N_209,In_719);
or U327 (N_327,In_1317,In_587);
nor U328 (N_328,In_428,N_26);
xor U329 (N_329,In_743,In_875);
nand U330 (N_330,In_393,In_444);
or U331 (N_331,In_1193,In_1174);
or U332 (N_332,N_97,N_127);
nand U333 (N_333,In_452,In_1277);
xor U334 (N_334,In_1226,In_1145);
or U335 (N_335,In_294,N_56);
and U336 (N_336,N_243,In_852);
xor U337 (N_337,In_1486,In_1246);
nand U338 (N_338,In_737,In_833);
or U339 (N_339,In_1439,N_43);
nor U340 (N_340,N_159,In_390);
nor U341 (N_341,In_899,N_144);
nand U342 (N_342,N_54,N_205);
nor U343 (N_343,In_292,N_106);
nor U344 (N_344,In_1054,In_584);
xor U345 (N_345,In_347,N_173);
nor U346 (N_346,In_616,In_410);
nor U347 (N_347,In_205,In_794);
or U348 (N_348,In_168,In_732);
or U349 (N_349,In_545,In_1015);
and U350 (N_350,In_1432,In_151);
or U351 (N_351,N_33,N_190);
nand U352 (N_352,In_1115,N_161);
and U353 (N_353,In_1441,In_1324);
xnor U354 (N_354,In_604,In_497);
nand U355 (N_355,N_213,N_211);
nand U356 (N_356,N_206,In_147);
and U357 (N_357,In_851,In_863);
xor U358 (N_358,In_1141,In_895);
nand U359 (N_359,In_1190,In_407);
nor U360 (N_360,In_787,In_917);
nand U361 (N_361,In_1364,In_774);
or U362 (N_362,In_893,In_504);
nor U363 (N_363,In_187,In_388);
nand U364 (N_364,In_191,In_488);
or U365 (N_365,N_143,In_986);
and U366 (N_366,In_1240,N_75);
or U367 (N_367,In_326,In_1477);
or U368 (N_368,In_1088,In_1418);
or U369 (N_369,In_722,N_34);
nor U370 (N_370,In_250,In_807);
nor U371 (N_371,In_1309,In_264);
or U372 (N_372,In_888,In_1270);
nand U373 (N_373,In_764,N_214);
or U374 (N_374,In_217,N_38);
nand U375 (N_375,In_692,In_1254);
nand U376 (N_376,In_735,In_827);
or U377 (N_377,In_1402,In_456);
or U378 (N_378,In_154,In_955);
and U379 (N_379,In_537,In_418);
and U380 (N_380,In_966,In_73);
nand U381 (N_381,In_445,In_940);
nor U382 (N_382,In_1200,In_281);
or U383 (N_383,In_1297,In_1298);
nor U384 (N_384,In_1024,N_140);
or U385 (N_385,In_103,In_593);
or U386 (N_386,In_1339,N_228);
nand U387 (N_387,In_699,In_652);
nor U388 (N_388,In_610,In_1411);
or U389 (N_389,In_1177,In_1326);
nor U390 (N_390,In_906,In_195);
nor U391 (N_391,In_183,In_1280);
or U392 (N_392,N_29,N_112);
nand U393 (N_393,N_18,In_344);
and U394 (N_394,In_83,In_1102);
nor U395 (N_395,In_166,N_71);
nor U396 (N_396,In_1022,In_261);
nor U397 (N_397,N_107,In_748);
nor U398 (N_398,In_1314,In_1379);
or U399 (N_399,In_1002,N_79);
nor U400 (N_400,N_238,In_1351);
or U401 (N_401,In_502,In_363);
or U402 (N_402,N_195,In_269);
nor U403 (N_403,In_1083,In_1064);
xnor U404 (N_404,In_1380,In_1003);
and U405 (N_405,In_395,In_465);
nor U406 (N_406,In_1073,In_1134);
or U407 (N_407,N_248,N_63);
nor U408 (N_408,In_550,In_256);
nand U409 (N_409,In_39,In_1383);
and U410 (N_410,In_323,In_601);
or U411 (N_411,In_1340,In_1255);
nor U412 (N_412,In_279,In_1406);
nor U413 (N_413,N_6,In_979);
nor U414 (N_414,In_961,In_1068);
nand U415 (N_415,In_377,In_1213);
or U416 (N_416,In_859,N_113);
nor U417 (N_417,In_1036,In_780);
or U418 (N_418,In_769,In_87);
nand U419 (N_419,In_1058,N_39);
and U420 (N_420,In_969,N_247);
or U421 (N_421,N_128,In_1322);
and U422 (N_422,In_664,In_343);
or U423 (N_423,N_48,In_957);
nor U424 (N_424,In_1276,In_1224);
nor U425 (N_425,N_30,In_1470);
or U426 (N_426,In_421,In_398);
nor U427 (N_427,In_1110,In_223);
nor U428 (N_428,In_600,In_1136);
nand U429 (N_429,In_576,In_583);
nor U430 (N_430,In_312,N_100);
xor U431 (N_431,In_678,In_952);
and U432 (N_432,In_319,In_301);
or U433 (N_433,In_394,In_1372);
nand U434 (N_434,In_542,In_192);
nor U435 (N_435,In_1393,In_1260);
and U436 (N_436,In_1362,N_249);
nand U437 (N_437,In_862,In_1263);
or U438 (N_438,In_403,N_207);
and U439 (N_439,In_1230,In_1033);
or U440 (N_440,In_801,N_36);
nand U441 (N_441,In_1384,In_634);
and U442 (N_442,In_27,In_34);
nor U443 (N_443,N_9,N_120);
or U444 (N_444,In_679,In_1464);
or U445 (N_445,In_1098,In_293);
nor U446 (N_446,N_84,In_1355);
nor U447 (N_447,In_200,In_1161);
and U448 (N_448,In_824,In_231);
and U449 (N_449,N_168,In_872);
nor U450 (N_450,In_1471,In_781);
nand U451 (N_451,In_225,In_561);
nand U452 (N_452,In_93,In_682);
and U453 (N_453,In_141,In_1252);
or U454 (N_454,In_697,In_543);
or U455 (N_455,In_146,In_246);
xnor U456 (N_456,In_573,In_1473);
nor U457 (N_457,In_746,N_5);
xnor U458 (N_458,In_108,N_155);
nand U459 (N_459,In_842,In_975);
nor U460 (N_460,In_1378,In_1288);
xnor U461 (N_461,In_60,In_64);
nor U462 (N_462,In_152,In_1371);
nor U463 (N_463,In_1202,In_617);
nor U464 (N_464,In_125,In_1241);
nor U465 (N_465,N_105,In_92);
nor U466 (N_466,In_1275,In_1283);
or U467 (N_467,In_914,N_41);
nand U468 (N_468,In_1109,In_998);
or U469 (N_469,In_1165,In_11);
xnor U470 (N_470,N_178,In_1476);
xnor U471 (N_471,In_1485,In_668);
nor U472 (N_472,In_591,In_944);
nand U473 (N_473,In_273,In_1294);
and U474 (N_474,In_12,In_529);
nor U475 (N_475,In_1430,In_690);
or U476 (N_476,In_925,N_177);
nor U477 (N_477,N_227,In_1392);
nand U478 (N_478,In_55,In_965);
or U479 (N_479,In_259,In_1093);
and U480 (N_480,In_1365,In_411);
or U481 (N_481,In_1377,In_1012);
and U482 (N_482,In_1066,N_201);
xor U483 (N_483,In_72,In_949);
or U484 (N_484,In_990,N_93);
nor U485 (N_485,In_409,In_1301);
and U486 (N_486,In_1081,N_47);
nand U487 (N_487,In_572,In_629);
xnor U488 (N_488,In_1345,In_586);
or U489 (N_489,In_557,N_85);
nand U490 (N_490,In_527,In_1201);
nand U491 (N_491,In_1368,In_376);
nand U492 (N_492,In_919,In_95);
and U493 (N_493,N_116,In_309);
nor U494 (N_494,In_354,In_563);
or U495 (N_495,In_1308,In_898);
nand U496 (N_496,In_1079,In_1272);
nand U497 (N_497,In_1090,N_80);
and U498 (N_498,N_11,N_233);
nand U499 (N_499,In_631,N_154);
nand U500 (N_500,In_1354,In_776);
and U501 (N_501,In_558,N_354);
nand U502 (N_502,In_1452,N_412);
nand U503 (N_503,N_419,In_467);
or U504 (N_504,In_1481,In_1350);
or U505 (N_505,In_414,In_753);
and U506 (N_506,In_435,In_1284);
or U507 (N_507,In_883,N_199);
xnor U508 (N_508,N_407,N_69);
nand U509 (N_509,N_102,In_702);
and U510 (N_510,N_439,N_250);
nor U511 (N_511,In_1461,In_1404);
nor U512 (N_512,In_585,In_983);
or U513 (N_513,N_367,In_788);
nor U514 (N_514,In_352,In_1047);
and U515 (N_515,N_194,In_803);
nor U516 (N_516,In_442,In_1261);
nor U517 (N_517,N_397,In_666);
nand U518 (N_518,N_20,In_336);
and U519 (N_519,In_876,In_184);
or U520 (N_520,N_495,In_711);
nor U521 (N_521,N_453,In_932);
xnor U522 (N_522,In_229,In_1140);
nor U523 (N_523,N_132,In_1037);
or U524 (N_524,In_206,N_322);
and U525 (N_525,In_1390,In_684);
and U526 (N_526,N_253,N_202);
nand U527 (N_527,In_399,In_861);
nand U528 (N_528,N_362,In_462);
nand U529 (N_529,In_254,In_779);
and U530 (N_530,N_426,N_160);
nand U531 (N_531,N_477,N_212);
or U532 (N_532,In_639,N_292);
xnor U533 (N_533,In_385,In_328);
and U534 (N_534,In_589,In_864);
nor U535 (N_535,In_1499,In_987);
and U536 (N_536,In_121,In_655);
nor U537 (N_537,In_286,N_196);
xor U538 (N_538,In_208,N_387);
nor U539 (N_539,In_662,In_71);
or U540 (N_540,In_163,In_1121);
and U541 (N_541,In_203,In_921);
nand U542 (N_542,N_139,N_276);
or U543 (N_543,N_208,In_705);
and U544 (N_544,N_185,In_663);
and U545 (N_545,In_982,N_437);
nor U546 (N_546,In_889,In_1336);
nor U547 (N_547,In_63,In_20);
nand U548 (N_548,N_423,In_516);
or U549 (N_549,N_115,N_98);
and U550 (N_550,In_484,In_912);
nor U551 (N_551,N_491,In_102);
and U552 (N_552,In_729,N_379);
or U553 (N_553,N_458,In_1039);
nor U554 (N_554,In_4,In_228);
and U555 (N_555,In_5,N_396);
or U556 (N_556,In_1311,In_211);
or U557 (N_557,In_37,N_220);
or U558 (N_558,In_900,N_288);
xor U559 (N_559,In_1474,In_1020);
and U560 (N_560,N_96,N_497);
and U561 (N_561,In_181,In_723);
or U562 (N_562,In_243,N_347);
nand U563 (N_563,N_408,In_1026);
or U564 (N_564,N_270,N_231);
or U565 (N_565,N_429,N_335);
or U566 (N_566,N_23,N_390);
nand U567 (N_567,In_1333,In_762);
or U568 (N_568,N_94,N_434);
nand U569 (N_569,N_417,In_1376);
nand U570 (N_570,In_300,In_866);
nand U571 (N_571,In_1172,N_312);
or U572 (N_572,In_908,In_1092);
xnor U573 (N_573,In_544,In_1112);
nor U574 (N_574,N_358,N_443);
nand U575 (N_575,N_24,N_255);
and U576 (N_576,N_370,In_341);
xnor U577 (N_577,In_1216,N_265);
and U578 (N_578,In_1125,N_267);
nor U579 (N_579,In_1342,In_215);
nor U580 (N_580,In_1157,N_361);
nand U581 (N_581,In_1279,N_395);
nand U582 (N_582,N_323,N_151);
nand U583 (N_583,N_319,In_609);
or U584 (N_584,In_82,In_727);
nand U585 (N_585,N_331,In_1286);
or U586 (N_586,In_954,In_6);
nor U587 (N_587,In_290,In_971);
or U588 (N_588,N_92,In_509);
nor U589 (N_589,N_149,N_488);
or U590 (N_590,In_1422,In_174);
nor U591 (N_591,N_404,In_1358);
nand U592 (N_592,N_371,In_904);
nor U593 (N_593,N_37,In_525);
nor U594 (N_594,In_1212,In_220);
and U595 (N_595,In_137,N_317);
nor U596 (N_596,N_285,In_338);
and U597 (N_597,In_1448,N_389);
nand U598 (N_598,N_340,In_740);
or U599 (N_599,In_470,In_717);
nor U600 (N_600,In_708,In_506);
nor U601 (N_601,In_447,N_448);
or U602 (N_602,In_643,N_333);
xnor U603 (N_603,N_350,In_128);
nor U604 (N_604,In_858,In_734);
and U605 (N_605,In_1122,In_538);
nand U606 (N_606,In_43,N_492);
and U607 (N_607,In_1105,N_46);
nor U608 (N_608,N_383,N_64);
and U609 (N_609,In_1304,N_215);
or U610 (N_610,N_480,In_56);
nor U611 (N_611,In_1443,In_327);
nor U612 (N_612,N_60,In_222);
nor U613 (N_613,In_913,In_933);
nor U614 (N_614,N_136,In_233);
and U615 (N_615,In_349,N_165);
nor U616 (N_616,In_271,N_313);
or U617 (N_617,N_82,N_123);
or U618 (N_618,N_193,In_567);
nor U619 (N_619,In_978,In_881);
nor U620 (N_620,N_254,N_17);
and U621 (N_621,In_160,In_284);
nand U622 (N_622,N_342,In_963);
and U623 (N_623,N_300,N_341);
and U624 (N_624,In_1256,N_451);
nor U625 (N_625,N_261,In_810);
nor U626 (N_626,In_453,N_237);
nand U627 (N_627,N_275,In_1236);
nand U628 (N_628,N_31,N_355);
nand U629 (N_629,In_1395,N_446);
nand U630 (N_630,N_171,In_880);
nor U631 (N_631,N_422,In_575);
nand U632 (N_632,In_877,N_2);
and U633 (N_633,N_66,In_1267);
or U634 (N_634,In_614,In_796);
and U635 (N_635,In_673,N_240);
and U636 (N_636,N_330,In_603);
and U637 (N_637,N_471,N_157);
nor U638 (N_638,In_42,In_169);
and U639 (N_639,In_902,N_459);
nor U640 (N_640,N_148,In_189);
xor U641 (N_641,In_931,In_951);
nor U642 (N_642,N_131,N_372);
nor U643 (N_643,In_1421,N_436);
or U644 (N_644,In_17,In_670);
nor U645 (N_645,In_1018,In_1046);
or U646 (N_646,In_817,In_683);
or U647 (N_647,N_182,N_51);
or U648 (N_648,In_873,In_1341);
and U649 (N_649,In_574,N_295);
or U650 (N_650,In_1382,N_262);
nand U651 (N_651,N_125,In_552);
nand U652 (N_652,In_1445,N_452);
and U653 (N_653,N_420,N_234);
nor U654 (N_654,In_536,In_188);
and U655 (N_655,N_427,N_298);
nand U656 (N_656,In_242,In_448);
and U657 (N_657,In_150,N_402);
and U658 (N_658,In_1130,In_44);
nand U659 (N_659,N_278,In_657);
or U660 (N_660,In_1248,In_1479);
or U661 (N_661,In_1038,In_1100);
and U662 (N_662,In_1097,N_235);
or U663 (N_663,In_910,N_388);
and U664 (N_664,In_656,In_1120);
nor U665 (N_665,N_61,In_848);
or U666 (N_666,In_433,N_462);
nor U667 (N_667,N_456,In_248);
nand U668 (N_668,N_134,N_356);
xor U669 (N_669,In_432,In_713);
nor U670 (N_670,N_413,N_186);
and U671 (N_671,In_1307,In_1373);
or U672 (N_672,N_183,In_35);
and U673 (N_673,N_83,N_307);
nand U674 (N_674,In_939,In_140);
nand U675 (N_675,N_391,In_592);
nor U676 (N_676,In_89,In_175);
xnor U677 (N_677,In_1397,N_418);
and U678 (N_678,N_481,In_1328);
xor U679 (N_679,In_54,N_325);
nor U680 (N_680,In_38,In_1069);
and U681 (N_681,In_304,N_192);
and U682 (N_682,N_81,In_1295);
and U683 (N_683,In_48,In_891);
nand U684 (N_684,In_1356,In_2);
and U685 (N_685,N_266,In_232);
nand U686 (N_686,In_1209,N_430);
or U687 (N_687,In_124,In_654);
and U688 (N_688,N_303,In_1117);
nand U689 (N_689,N_174,N_339);
nand U690 (N_690,N_53,In_1080);
xnor U691 (N_691,In_1434,In_1268);
or U692 (N_692,In_1428,In_1056);
nor U693 (N_693,In_1433,N_470);
nand U694 (N_694,N_95,In_131);
or U695 (N_695,N_204,In_531);
or U696 (N_696,N_400,In_386);
nand U697 (N_697,N_324,In_1227);
and U698 (N_698,N_163,In_283);
or U699 (N_699,In_287,In_1051);
or U700 (N_700,N_499,In_918);
xor U701 (N_701,N_138,N_251);
or U702 (N_702,In_767,N_284);
nor U703 (N_703,In_1420,In_491);
nor U704 (N_704,N_447,In_104);
nand U705 (N_705,In_1492,In_245);
nand U706 (N_706,In_339,In_358);
xnor U707 (N_707,N_428,N_25);
and U708 (N_708,N_398,In_1305);
and U709 (N_709,In_68,In_268);
nand U710 (N_710,In_361,In_58);
nor U711 (N_711,N_119,N_344);
nand U712 (N_712,N_380,N_191);
nand U713 (N_713,In_805,In_1215);
nand U714 (N_714,In_1335,In_1253);
nand U715 (N_715,In_1034,N_246);
and U716 (N_716,In_946,N_289);
and U717 (N_717,N_121,N_455);
nor U718 (N_718,In_1170,In_110);
and U719 (N_719,N_76,In_468);
nor U720 (N_720,In_1331,N_304);
and U721 (N_721,N_42,In_523);
nand U722 (N_722,N_281,N_65);
nand U723 (N_723,In_745,In_1222);
and U724 (N_724,In_367,N_454);
nor U725 (N_725,N_259,N_345);
xnor U726 (N_726,N_135,N_386);
nand U727 (N_727,In_784,N_241);
nand U728 (N_728,N_472,N_438);
or U729 (N_729,In_75,In_1343);
xor U730 (N_730,In_632,In_916);
and U731 (N_731,In_571,N_226);
nand U732 (N_732,In_1423,N_376);
nor U733 (N_733,N_118,In_489);
nand U734 (N_734,In_142,In_947);
nand U735 (N_735,In_1244,In_129);
nand U736 (N_736,N_137,In_1447);
and U737 (N_737,In_879,In_374);
nor U738 (N_738,In_1352,N_293);
nor U739 (N_739,N_10,N_320);
or U740 (N_740,In_867,In_922);
nor U741 (N_741,N_269,N_353);
and U742 (N_742,N_296,In_1151);
nand U743 (N_743,In_526,In_1483);
or U744 (N_744,N_308,In_479);
and U745 (N_745,N_406,In_1466);
or U746 (N_746,N_282,In_306);
and U747 (N_747,In_714,N_19);
and U748 (N_748,In_379,In_1497);
xnor U749 (N_749,In_310,In_193);
nand U750 (N_750,N_473,In_997);
and U751 (N_751,N_264,In_1044);
nand U752 (N_752,N_727,N_476);
or U753 (N_753,In_1332,N_373);
and U754 (N_754,In_255,N_582);
or U755 (N_755,N_618,In_621);
xnor U756 (N_756,N_363,N_747);
or U757 (N_757,In_70,In_29);
and U758 (N_758,N_634,N_283);
nand U759 (N_759,N_603,In_258);
and U760 (N_760,N_657,N_672);
xor U761 (N_761,In_213,N_494);
nor U762 (N_762,N_578,N_636);
nand U763 (N_763,In_905,In_1063);
xnor U764 (N_764,In_989,N_552);
and U765 (N_765,N_432,N_302);
nor U766 (N_766,N_167,In_267);
xnor U767 (N_767,N_604,In_382);
xor U768 (N_768,N_644,N_216);
or U769 (N_769,In_1194,N_587);
nand U770 (N_770,N_385,In_674);
nor U771 (N_771,In_1060,In_272);
nand U772 (N_772,N_653,In_1113);
and U773 (N_773,In_934,N_498);
or U774 (N_774,In_179,N_503);
or U775 (N_775,N_433,In_1451);
nand U776 (N_776,In_1398,N_501);
nor U777 (N_777,In_240,In_1206);
or U778 (N_778,N_217,N_545);
and U779 (N_779,In_1494,In_487);
nand U780 (N_780,N_365,In_1043);
and U781 (N_781,N_507,In_1480);
or U782 (N_782,In_1225,N_508);
or U783 (N_783,In_164,N_109);
nor U784 (N_784,In_80,In_594);
xor U785 (N_785,N_328,In_577);
nand U786 (N_786,N_424,N_534);
or U787 (N_787,N_124,N_461);
nand U788 (N_788,In_897,N_533);
nor U789 (N_789,N_725,In_380);
or U790 (N_790,N_695,N_381);
nand U791 (N_791,N_702,In_804);
or U792 (N_792,In_1232,In_249);
xor U793 (N_793,In_795,N_502);
nand U794 (N_794,In_1438,N_153);
and U795 (N_795,In_157,N_518);
nor U796 (N_796,N_542,N_748);
nor U797 (N_797,N_274,N_639);
or U798 (N_798,N_572,N_463);
nor U799 (N_799,In_628,N_180);
and U800 (N_800,N_57,In_1424);
nand U801 (N_801,N_532,N_525);
xor U802 (N_802,N_263,N_585);
nor U803 (N_803,In_597,N_3);
xnor U804 (N_804,N_647,N_431);
and U805 (N_805,N_628,N_297);
nand U806 (N_806,N_425,N_660);
and U807 (N_807,N_357,In_431);
nand U808 (N_808,In_115,N_611);
or U809 (N_809,In_1278,In_404);
or U810 (N_810,N_466,N_527);
and U811 (N_811,N_489,N_50);
nand U812 (N_812,In_818,In_1094);
and U813 (N_813,In_1017,N_150);
nand U814 (N_814,In_736,In_1285);
nor U815 (N_815,In_1175,N_720);
xnor U816 (N_816,In_800,In_1169);
or U817 (N_817,N_91,N_244);
or U818 (N_818,N_599,In_1149);
nand U819 (N_819,N_515,In_581);
nand U820 (N_820,In_995,N_682);
and U821 (N_821,N_715,N_32);
nor U822 (N_822,N_712,N_600);
nor U823 (N_823,In_959,In_1299);
or U824 (N_824,In_885,N_181);
nand U825 (N_825,N_286,In_554);
or U826 (N_826,N_537,In_57);
nand U827 (N_827,N_737,N_743);
and U828 (N_828,N_74,In_274);
and U829 (N_829,In_277,N_625);
nor U830 (N_830,N_576,N_593);
and U831 (N_831,N_15,N_359);
nand U832 (N_832,N_384,In_118);
or U833 (N_833,In_1045,In_112);
xor U834 (N_834,In_1128,N_169);
nand U835 (N_835,In_77,In_303);
xnor U836 (N_836,N_531,N_718);
nand U837 (N_837,N_726,N_334);
nand U838 (N_838,In_813,N_72);
nor U839 (N_839,N_351,N_592);
or U840 (N_840,N_692,In_675);
and U841 (N_841,N_590,In_884);
or U842 (N_842,N_613,N_393);
nor U843 (N_843,N_684,N_101);
or U844 (N_844,In_1442,In_1484);
or U845 (N_845,In_373,N_553);
or U846 (N_846,In_133,N_530);
nor U847 (N_847,N_557,In_1041);
nand U848 (N_848,N_675,N_687);
or U849 (N_849,N_729,N_375);
and U850 (N_850,N_619,N_724);
nor U851 (N_851,In_1061,In_640);
nor U852 (N_852,N_719,N_457);
or U853 (N_853,In_1367,In_368);
or U854 (N_854,N_126,In_61);
nor U855 (N_855,N_280,In_1049);
nor U856 (N_856,N_674,N_364);
nor U857 (N_857,N_560,N_326);
and U858 (N_858,In_739,N_668);
or U859 (N_859,In_823,In_415);
nand U860 (N_860,N_554,N_224);
or U861 (N_861,N_669,N_732);
nor U862 (N_862,N_479,In_375);
xnor U863 (N_863,N_221,N_708);
or U864 (N_864,In_480,N_610);
nand U865 (N_865,In_929,N_705);
nand U866 (N_866,In_1385,N_623);
xor U867 (N_867,In_992,N_617);
and U868 (N_868,In_855,In_221);
nor U869 (N_869,In_69,In_490);
or U870 (N_870,In_1208,In_408);
nand U871 (N_871,In_755,N_291);
or U872 (N_872,N_703,N_701);
nand U873 (N_873,N_549,In_96);
nor U874 (N_874,N_577,N_573);
or U875 (N_875,In_1062,N_602);
or U876 (N_876,N_706,N_166);
or U877 (N_877,N_49,N_689);
or U878 (N_878,N_67,N_277);
nand U879 (N_879,In_580,N_467);
and U880 (N_880,N_273,N_627);
or U881 (N_881,In_461,In_1);
and U882 (N_882,In_1369,N_176);
nor U883 (N_883,N_671,In_999);
or U884 (N_884,In_451,N_440);
or U885 (N_885,In_1167,N_487);
and U886 (N_886,N_409,In_564);
and U887 (N_887,In_595,In_1048);
or U888 (N_888,N_474,N_567);
nand U889 (N_889,N_315,In_1198);
and U890 (N_890,N_523,In_165);
and U891 (N_891,N_609,In_332);
or U892 (N_892,N_117,In_446);
or U893 (N_893,N_252,In_521);
xnor U894 (N_894,N_667,N_294);
nor U895 (N_895,In_809,N_655);
nand U896 (N_896,N_722,N_691);
and U897 (N_897,N_646,N_318);
nand U898 (N_898,N_562,N_486);
or U899 (N_899,N_435,N_654);
nor U900 (N_900,N_329,N_239);
or U901 (N_901,N_574,N_526);
nand U902 (N_902,N_519,N_225);
nand U903 (N_903,N_377,In_890);
or U904 (N_904,N_641,N_58);
or U905 (N_905,In_871,N_343);
nand U906 (N_906,N_699,N_460);
nor U907 (N_907,N_598,N_561);
and U908 (N_908,N_45,In_689);
nand U909 (N_909,In_907,N_568);
nand U910 (N_910,In_149,N_739);
nand U911 (N_911,N_78,N_89);
or U912 (N_912,N_374,N_612);
and U913 (N_913,N_99,N_694);
nand U914 (N_914,N_493,In_459);
nand U915 (N_915,N_368,N_607);
nand U916 (N_916,N_632,In_1262);
xor U917 (N_917,In_458,N_110);
xor U918 (N_918,In_1414,N_524);
xnor U919 (N_919,N_622,N_505);
xor U920 (N_920,N_392,In_23);
nand U921 (N_921,N_643,In_1287);
nor U922 (N_922,N_22,N_414);
xnor U923 (N_923,In_1348,N_544);
or U924 (N_924,N_449,In_569);
or U925 (N_925,N_490,In_837);
xor U926 (N_926,N_90,N_640);
and U927 (N_927,N_538,In_74);
and U928 (N_928,N_536,N_741);
nand U929 (N_929,N_348,In_210);
or U930 (N_930,N_711,In_1490);
and U931 (N_931,N_145,N_366);
and U932 (N_932,N_749,In_994);
nand U933 (N_933,In_483,N_575);
nor U934 (N_934,In_843,In_1396);
nor U935 (N_935,N_475,N_521);
or U936 (N_936,In_1403,In_247);
and U937 (N_937,N_745,In_400);
nor U938 (N_938,N_734,N_258);
and U939 (N_939,In_936,N_735);
xnor U940 (N_940,In_507,N_88);
nor U941 (N_941,In_0,In_555);
and U942 (N_942,N_679,In_1251);
nor U943 (N_943,N_620,In_158);
nand U944 (N_944,In_1468,N_676);
or U945 (N_945,N_401,N_416);
nand U946 (N_946,In_159,N_730);
and U947 (N_947,N_198,In_126);
or U948 (N_948,In_808,N_223);
nand U949 (N_949,In_1075,N_257);
nand U950 (N_950,N_104,N_511);
or U951 (N_951,In_412,In_424);
or U952 (N_952,N_744,In_738);
and U953 (N_953,In_726,N_44);
nor U954 (N_954,N_415,N_638);
nor U955 (N_955,In_1163,N_59);
nor U956 (N_956,N_648,N_77);
and U957 (N_957,N_290,N_268);
and U958 (N_958,N_586,In_186);
nand U959 (N_959,In_106,N_529);
xnor U960 (N_960,N_547,In_120);
and U961 (N_961,N_68,N_595);
or U962 (N_962,In_485,N_652);
nor U963 (N_963,N_483,In_945);
or U964 (N_964,N_665,N_710);
nand U965 (N_965,N_465,N_232);
or U966 (N_966,In_772,In_198);
or U967 (N_967,N_555,N_73);
nand U968 (N_968,N_442,In_896);
nor U969 (N_969,N_129,N_566);
nand U970 (N_970,N_738,In_1204);
nor U971 (N_971,N_709,In_346);
nor U972 (N_972,N_571,In_1417);
xor U973 (N_973,In_1250,N_594);
nor U974 (N_974,N_133,In_624);
nor U975 (N_975,N_27,N_405);
and U976 (N_976,N_642,In_1409);
nor U977 (N_977,N_673,N_338);
or U978 (N_978,N_704,In_334);
nand U979 (N_979,N_677,N_740);
nand U980 (N_980,N_218,N_535);
nand U981 (N_981,N_651,N_219);
xor U982 (N_982,In_1123,In_1291);
nand U983 (N_983,In_145,N_608);
or U984 (N_984,In_712,In_514);
and U985 (N_985,N_152,N_661);
and U986 (N_986,N_321,N_504);
or U987 (N_987,N_87,N_444);
or U988 (N_988,N_565,In_1359);
nor U989 (N_989,N_633,In_1023);
and U990 (N_990,N_450,N_346);
nand U991 (N_991,N_746,In_359);
xnor U992 (N_992,N_514,N_314);
xor U993 (N_993,N_229,N_614);
and U994 (N_994,In_1138,N_394);
nor U995 (N_995,N_696,In_1229);
nand U996 (N_996,N_678,In_1078);
nand U997 (N_997,In_99,N_399);
nand U998 (N_998,In_1077,In_387);
or U999 (N_999,In_136,N_601);
nor U1000 (N_1000,In_1323,In_970);
nand U1001 (N_1001,N_976,N_811);
and U1002 (N_1002,N_581,N_605);
nor U1003 (N_1003,In_1233,N_787);
or U1004 (N_1004,N_336,In_786);
xnor U1005 (N_1005,N_752,N_774);
xor U1006 (N_1006,N_893,N_775);
and U1007 (N_1007,N_516,N_813);
or U1008 (N_1008,N_803,N_543);
nor U1009 (N_1009,N_945,N_635);
or U1010 (N_1010,N_770,N_802);
nor U1011 (N_1011,In_180,N_597);
xnor U1012 (N_1012,N_751,N_658);
and U1013 (N_1013,In_676,N_841);
nor U1014 (N_1014,N_310,N_306);
nand U1015 (N_1015,N_861,In_1131);
xnor U1016 (N_1016,N_287,N_685);
nor U1017 (N_1017,N_925,In_135);
nand U1018 (N_1018,N_659,N_823);
and U1019 (N_1019,N_776,In_241);
nand U1020 (N_1020,N_421,N_753);
and U1021 (N_1021,N_954,In_1087);
and U1022 (N_1022,N_580,N_0);
or U1023 (N_1023,N_860,N_889);
or U1024 (N_1024,N_795,N_798);
nor U1025 (N_1025,N_990,In_799);
xor U1026 (N_1026,N_790,N_822);
nand U1027 (N_1027,N_271,In_953);
and U1028 (N_1028,In_162,N_924);
and U1029 (N_1029,N_839,In_1337);
and U1030 (N_1030,N_736,In_672);
nor U1031 (N_1031,N_875,N_700);
nor U1032 (N_1032,N_937,In_1407);
nand U1033 (N_1033,N_833,In_820);
nor U1034 (N_1034,N_482,N_907);
or U1035 (N_1035,N_936,In_868);
and U1036 (N_1036,N_940,N_804);
nor U1037 (N_1037,N_917,In_1386);
nor U1038 (N_1038,In_493,In_1346);
or U1039 (N_1039,N_984,In_1495);
xor U1040 (N_1040,In_620,N_894);
xor U1041 (N_1041,N_949,N_539);
or U1042 (N_1042,In_182,In_219);
nor U1043 (N_1043,N_817,N_688);
nor U1044 (N_1044,In_473,N_563);
or U1045 (N_1045,N_332,N_903);
xor U1046 (N_1046,N_550,N_978);
xor U1047 (N_1047,N_403,N_510);
nor U1048 (N_1048,N_809,N_849);
nand U1049 (N_1049,In_648,N_878);
nand U1050 (N_1050,N_716,N_974);
nand U1051 (N_1051,N_807,In_570);
and U1052 (N_1052,N_411,N_961);
nand U1053 (N_1053,In_596,N_584);
nand U1054 (N_1054,N_360,N_828);
and U1055 (N_1055,N_800,N_956);
or U1056 (N_1056,N_801,N_793);
or U1057 (N_1057,N_588,N_970);
and U1058 (N_1058,In_1118,N_955);
xor U1059 (N_1059,In_1160,N_980);
nand U1060 (N_1060,N_950,N_272);
nor U1061 (N_1061,N_832,N_884);
or U1062 (N_1062,N_666,N_964);
nor U1063 (N_1063,In_1019,In_1292);
nand U1064 (N_1064,N_818,N_819);
or U1065 (N_1065,N_886,N_926);
and U1066 (N_1066,N_898,N_778);
xnor U1067 (N_1067,N_777,N_142);
nor U1068 (N_1068,N_656,N_680);
and U1069 (N_1069,N_830,N_847);
and U1070 (N_1070,N_757,N_988);
and U1071 (N_1071,N_768,In_402);
nor U1072 (N_1072,In_107,N_836);
nand U1073 (N_1073,N_857,N_873);
or U1074 (N_1074,N_966,N_859);
and U1075 (N_1075,N_8,N_897);
and U1076 (N_1076,In_1425,N_957);
nor U1077 (N_1077,In_302,N_838);
nor U1078 (N_1078,In_238,N_868);
or U1079 (N_1079,N_352,N_179);
nor U1080 (N_1080,N_681,N_1);
nand U1081 (N_1081,N_879,N_520);
or U1082 (N_1082,N_570,N_779);
or U1083 (N_1083,N_14,N_944);
and U1084 (N_1084,N_871,N_969);
and U1085 (N_1085,N_305,N_971);
nand U1086 (N_1086,N_880,N_626);
and U1087 (N_1087,N_981,N_693);
nor U1088 (N_1088,In_613,N_837);
xnor U1089 (N_1089,In_236,N_987);
or U1090 (N_1090,N_992,N_781);
and U1091 (N_1091,In_1135,N_670);
and U1092 (N_1092,N_901,N_522);
or U1093 (N_1093,In_1183,N_763);
or U1094 (N_1094,N_941,N_853);
nor U1095 (N_1095,N_200,In_397);
nor U1096 (N_1096,N_918,N_864);
or U1097 (N_1097,N_929,N_863);
and U1098 (N_1098,N_756,N_707);
and U1099 (N_1099,N_517,N_441);
and U1100 (N_1100,In_1269,N_690);
or U1101 (N_1101,N_848,In_882);
xnor U1102 (N_1102,In_948,In_515);
nor U1103 (N_1103,In_1266,N_887);
or U1104 (N_1104,N_606,In_1095);
and U1105 (N_1105,In_1312,N_596);
nand U1106 (N_1106,N_892,N_994);
and U1107 (N_1107,N_899,N_629);
or U1108 (N_1108,N_108,N_927);
nand U1109 (N_1109,N_662,N_855);
nor U1110 (N_1110,In_696,N_378);
nand U1111 (N_1111,N_891,N_714);
nand U1112 (N_1112,N_900,N_904);
nand U1113 (N_1113,N_867,N_989);
or U1114 (N_1114,N_279,N_713);
xnor U1115 (N_1115,N_946,N_834);
nor U1116 (N_1116,N_888,In_832);
nor U1117 (N_1117,N_983,In_1188);
xnor U1118 (N_1118,N_915,In_1478);
nor U1119 (N_1119,In_765,N_920);
and U1120 (N_1120,In_1243,N_242);
or U1121 (N_1121,N_808,N_769);
nand U1122 (N_1122,In_615,N_569);
nor U1123 (N_1123,N_876,N_464);
xnor U1124 (N_1124,In_1021,N_968);
or U1125 (N_1125,N_870,N_951);
xor U1126 (N_1126,N_869,N_995);
or U1127 (N_1127,In_207,N_979);
and U1128 (N_1128,N_548,N_916);
and U1129 (N_1129,N_615,In_144);
nor U1130 (N_1130,N_723,In_937);
nor U1131 (N_1131,N_999,In_1181);
and U1132 (N_1132,N_509,N_773);
xor U1133 (N_1133,In_1303,N_967);
or U1134 (N_1134,N_928,N_299);
nand U1135 (N_1135,In_155,In_968);
xnor U1136 (N_1136,N_882,N_759);
nand U1137 (N_1137,N_972,N_883);
and U1138 (N_1138,N_986,In_351);
or U1139 (N_1139,In_1264,N_842);
nand U1140 (N_1140,N_28,N_663);
and U1141 (N_1141,In_669,In_856);
and U1142 (N_1142,N_827,N_923);
nand U1143 (N_1143,N_934,N_513);
and U1144 (N_1144,N_500,N_579);
xnor U1145 (N_1145,N_975,N_156);
and U1146 (N_1146,In_623,N_794);
nor U1147 (N_1147,N_496,In_1456);
nand U1148 (N_1148,In_1184,N_260);
and U1149 (N_1149,N_821,N_624);
or U1150 (N_1150,In_416,In_204);
xor U1151 (N_1151,N_858,In_725);
xor U1152 (N_1152,N_960,N_846);
nor U1153 (N_1153,In_1146,In_1162);
and U1154 (N_1154,N_829,In_111);
nand U1155 (N_1155,N_885,N_754);
and U1156 (N_1156,In_1394,N_559);
and U1157 (N_1157,N_469,N_784);
and U1158 (N_1158,In_65,N_558);
xor U1159 (N_1159,N_616,N_997);
nor U1160 (N_1160,N_783,N_445);
nand U1161 (N_1161,N_799,N_309);
nand U1162 (N_1162,N_850,N_985);
xnor U1163 (N_1163,N_788,N_812);
or U1164 (N_1164,N_311,N_906);
and U1165 (N_1165,N_506,N_301);
nor U1166 (N_1166,N_650,N_721);
and U1167 (N_1167,N_780,In_85);
or U1168 (N_1168,N_913,N_468);
nand U1169 (N_1169,N_912,N_792);
nand U1170 (N_1170,In_1315,N_478);
nand U1171 (N_1171,N_814,N_910);
or U1172 (N_1172,N_583,In_742);
nand U1173 (N_1173,N_905,In_647);
nor U1174 (N_1174,N_909,N_872);
xor U1175 (N_1175,N_919,In_1357);
nor U1176 (N_1176,N_782,N_844);
nor U1177 (N_1177,In_510,N_764);
xor U1178 (N_1178,N_728,N_541);
and U1179 (N_1179,N_645,N_824);
and U1180 (N_1180,In_811,In_235);
nor U1181 (N_1181,N_742,N_835);
nand U1182 (N_1182,N_933,N_820);
and U1183 (N_1183,N_922,N_998);
and U1184 (N_1184,N_786,N_826);
or U1185 (N_1185,N_958,N_942);
or U1186 (N_1186,N_758,N_698);
xor U1187 (N_1187,N_760,In_237);
and U1188 (N_1188,N_750,N_816);
and U1189 (N_1189,N_825,N_935);
nand U1190 (N_1190,N_591,N_256);
and U1191 (N_1191,N_512,N_664);
nand U1192 (N_1192,In_701,N_902);
or U1193 (N_1193,N_948,N_952);
and U1194 (N_1194,In_802,N_914);
and U1195 (N_1195,N_649,N_852);
nor U1196 (N_1196,N_731,N_35);
nand U1197 (N_1197,N_890,N_996);
nand U1198 (N_1198,In_350,In_915);
xor U1199 (N_1199,N_349,N_963);
nand U1200 (N_1200,N_197,N_546);
and U1201 (N_1201,N_556,N_791);
nand U1202 (N_1202,In_1164,N_410);
nand U1203 (N_1203,N_717,N_686);
nand U1204 (N_1204,In_383,N_856);
nand U1205 (N_1205,N_840,N_86);
nor U1206 (N_1206,N_785,N_843);
nor U1207 (N_1207,In_333,In_1449);
nor U1208 (N_1208,N_874,N_369);
nand U1209 (N_1209,N_564,N_865);
or U1210 (N_1210,N_762,N_797);
nor U1211 (N_1211,N_845,N_796);
or U1212 (N_1212,N_789,N_881);
nand U1213 (N_1213,N_203,N_528);
and U1214 (N_1214,N_683,N_805);
nand U1215 (N_1215,N_993,N_772);
nor U1216 (N_1216,N_962,N_982);
xor U1217 (N_1217,N_932,N_877);
nand U1218 (N_1218,N_911,N_959);
and U1219 (N_1219,N_965,N_4);
nor U1220 (N_1220,N_540,N_896);
or U1221 (N_1221,N_767,In_262);
nand U1222 (N_1222,N_895,N_146);
or U1223 (N_1223,N_765,In_1427);
or U1224 (N_1224,N_931,N_973);
and U1225 (N_1225,N_851,N_755);
nor U1226 (N_1226,N_908,N_930);
nand U1227 (N_1227,N_337,N_327);
and U1228 (N_1228,In_496,N_815);
and U1229 (N_1229,N_939,In_549);
or U1230 (N_1230,N_697,N_977);
nand U1231 (N_1231,N_806,N_637);
nand U1232 (N_1232,N_943,N_854);
or U1233 (N_1233,In_1482,N_766);
or U1234 (N_1234,N_52,N_938);
and U1235 (N_1235,N_921,N_862);
and U1236 (N_1236,In_680,N_953);
nor U1237 (N_1237,N_831,N_631);
xor U1238 (N_1238,N_316,N_771);
nand U1239 (N_1239,N_866,N_810);
nand U1240 (N_1240,N_236,N_589);
or U1241 (N_1241,In_127,N_621);
nand U1242 (N_1242,In_18,N_761);
nor U1243 (N_1243,N_991,N_630);
nand U1244 (N_1244,N_551,N_485);
nor U1245 (N_1245,N_382,N_733);
nor U1246 (N_1246,In_1137,In_1114);
nor U1247 (N_1247,N_230,In_1416);
nor U1248 (N_1248,In_486,N_947);
nand U1249 (N_1249,N_484,In_1008);
and U1250 (N_1250,N_1144,N_1186);
nor U1251 (N_1251,N_1002,N_1006);
or U1252 (N_1252,N_1185,N_1188);
and U1253 (N_1253,N_1178,N_1001);
nor U1254 (N_1254,N_1096,N_1079);
nand U1255 (N_1255,N_1154,N_1242);
nand U1256 (N_1256,N_1100,N_1166);
nand U1257 (N_1257,N_1072,N_1080);
nor U1258 (N_1258,N_1011,N_1152);
nor U1259 (N_1259,N_1134,N_1123);
xor U1260 (N_1260,N_1076,N_1075);
nor U1261 (N_1261,N_1232,N_1170);
and U1262 (N_1262,N_1004,N_1065);
nor U1263 (N_1263,N_1095,N_1026);
or U1264 (N_1264,N_1235,N_1051);
nand U1265 (N_1265,N_1248,N_1088);
and U1266 (N_1266,N_1056,N_1145);
xor U1267 (N_1267,N_1191,N_1227);
nor U1268 (N_1268,N_1219,N_1163);
xor U1269 (N_1269,N_1125,N_1069);
and U1270 (N_1270,N_1031,N_1119);
xor U1271 (N_1271,N_1244,N_1218);
nor U1272 (N_1272,N_1099,N_1043);
or U1273 (N_1273,N_1038,N_1087);
or U1274 (N_1274,N_1236,N_1239);
nand U1275 (N_1275,N_1103,N_1193);
nor U1276 (N_1276,N_1113,N_1046);
nand U1277 (N_1277,N_1211,N_1008);
nor U1278 (N_1278,N_1199,N_1161);
or U1279 (N_1279,N_1019,N_1128);
nand U1280 (N_1280,N_1139,N_1068);
or U1281 (N_1281,N_1210,N_1017);
or U1282 (N_1282,N_1212,N_1115);
and U1283 (N_1283,N_1053,N_1034);
nand U1284 (N_1284,N_1222,N_1184);
and U1285 (N_1285,N_1246,N_1045);
or U1286 (N_1286,N_1054,N_1165);
nand U1287 (N_1287,N_1225,N_1141);
nand U1288 (N_1288,N_1206,N_1195);
and U1289 (N_1289,N_1176,N_1122);
nand U1290 (N_1290,N_1117,N_1175);
or U1291 (N_1291,N_1209,N_1084);
and U1292 (N_1292,N_1149,N_1156);
and U1293 (N_1293,N_1021,N_1231);
xnor U1294 (N_1294,N_1097,N_1120);
and U1295 (N_1295,N_1090,N_1005);
nand U1296 (N_1296,N_1171,N_1027);
nor U1297 (N_1297,N_1007,N_1058);
nand U1298 (N_1298,N_1140,N_1180);
nor U1299 (N_1299,N_1025,N_1213);
or U1300 (N_1300,N_1245,N_1015);
nand U1301 (N_1301,N_1229,N_1063);
xor U1302 (N_1302,N_1077,N_1224);
nor U1303 (N_1303,N_1055,N_1190);
nor U1304 (N_1304,N_1086,N_1220);
nand U1305 (N_1305,N_1057,N_1143);
or U1306 (N_1306,N_1137,N_1040);
and U1307 (N_1307,N_1108,N_1129);
or U1308 (N_1308,N_1150,N_1221);
or U1309 (N_1309,N_1033,N_1121);
nand U1310 (N_1310,N_1030,N_1216);
nand U1311 (N_1311,N_1238,N_1164);
and U1312 (N_1312,N_1203,N_1240);
nor U1313 (N_1313,N_1059,N_1102);
nand U1314 (N_1314,N_1182,N_1196);
or U1315 (N_1315,N_1064,N_1228);
or U1316 (N_1316,N_1052,N_1130);
nand U1317 (N_1317,N_1142,N_1197);
or U1318 (N_1318,N_1172,N_1024);
nand U1319 (N_1319,N_1094,N_1157);
and U1320 (N_1320,N_1018,N_1158);
nor U1321 (N_1321,N_1060,N_1013);
or U1322 (N_1322,N_1237,N_1020);
and U1323 (N_1323,N_1230,N_1135);
and U1324 (N_1324,N_1133,N_1214);
xor U1325 (N_1325,N_1151,N_1061);
nand U1326 (N_1326,N_1098,N_1116);
nor U1327 (N_1327,N_1041,N_1029);
and U1328 (N_1328,N_1010,N_1067);
nor U1329 (N_1329,N_1155,N_1204);
nand U1330 (N_1330,N_1162,N_1070);
xnor U1331 (N_1331,N_1153,N_1009);
and U1332 (N_1332,N_1249,N_1168);
or U1333 (N_1333,N_1016,N_1159);
and U1334 (N_1334,N_1234,N_1181);
or U1335 (N_1335,N_1147,N_1071);
nand U1336 (N_1336,N_1187,N_1112);
and U1337 (N_1337,N_1091,N_1243);
xor U1338 (N_1338,N_1192,N_1014);
nor U1339 (N_1339,N_1132,N_1201);
nor U1340 (N_1340,N_1124,N_1082);
nand U1341 (N_1341,N_1114,N_1101);
nand U1342 (N_1342,N_1198,N_1160);
or U1343 (N_1343,N_1223,N_1208);
nor U1344 (N_1344,N_1173,N_1194);
or U1345 (N_1345,N_1105,N_1032);
and U1346 (N_1346,N_1022,N_1215);
nor U1347 (N_1347,N_1174,N_1044);
nand U1348 (N_1348,N_1036,N_1189);
nand U1349 (N_1349,N_1217,N_1138);
or U1350 (N_1350,N_1118,N_1126);
nand U1351 (N_1351,N_1106,N_1247);
nor U1352 (N_1352,N_1066,N_1104);
nor U1353 (N_1353,N_1028,N_1131);
and U1354 (N_1354,N_1148,N_1035);
and U1355 (N_1355,N_1167,N_1241);
nor U1356 (N_1356,N_1136,N_1000);
nor U1357 (N_1357,N_1089,N_1042);
nand U1358 (N_1358,N_1233,N_1107);
xor U1359 (N_1359,N_1177,N_1023);
nor U1360 (N_1360,N_1093,N_1085);
or U1361 (N_1361,N_1207,N_1078);
and U1362 (N_1362,N_1012,N_1092);
or U1363 (N_1363,N_1083,N_1074);
nor U1364 (N_1364,N_1081,N_1146);
or U1365 (N_1365,N_1205,N_1062);
and U1366 (N_1366,N_1226,N_1169);
nor U1367 (N_1367,N_1039,N_1202);
nor U1368 (N_1368,N_1109,N_1003);
or U1369 (N_1369,N_1111,N_1200);
or U1370 (N_1370,N_1048,N_1037);
or U1371 (N_1371,N_1049,N_1073);
nand U1372 (N_1372,N_1127,N_1050);
or U1373 (N_1373,N_1183,N_1047);
xnor U1374 (N_1374,N_1110,N_1179);
nand U1375 (N_1375,N_1126,N_1029);
nand U1376 (N_1376,N_1020,N_1001);
xor U1377 (N_1377,N_1183,N_1232);
nand U1378 (N_1378,N_1072,N_1091);
and U1379 (N_1379,N_1013,N_1102);
nor U1380 (N_1380,N_1059,N_1243);
and U1381 (N_1381,N_1246,N_1161);
or U1382 (N_1382,N_1046,N_1145);
or U1383 (N_1383,N_1009,N_1202);
or U1384 (N_1384,N_1116,N_1234);
nand U1385 (N_1385,N_1014,N_1005);
nor U1386 (N_1386,N_1234,N_1045);
and U1387 (N_1387,N_1052,N_1011);
xnor U1388 (N_1388,N_1162,N_1047);
and U1389 (N_1389,N_1133,N_1095);
nor U1390 (N_1390,N_1188,N_1085);
nor U1391 (N_1391,N_1199,N_1096);
nand U1392 (N_1392,N_1230,N_1244);
nand U1393 (N_1393,N_1244,N_1152);
or U1394 (N_1394,N_1102,N_1099);
nor U1395 (N_1395,N_1119,N_1187);
xor U1396 (N_1396,N_1194,N_1178);
and U1397 (N_1397,N_1225,N_1001);
nand U1398 (N_1398,N_1058,N_1086);
and U1399 (N_1399,N_1099,N_1187);
nand U1400 (N_1400,N_1217,N_1154);
or U1401 (N_1401,N_1027,N_1090);
and U1402 (N_1402,N_1002,N_1017);
nor U1403 (N_1403,N_1150,N_1074);
and U1404 (N_1404,N_1098,N_1071);
nor U1405 (N_1405,N_1147,N_1068);
nor U1406 (N_1406,N_1015,N_1013);
or U1407 (N_1407,N_1007,N_1106);
nand U1408 (N_1408,N_1139,N_1183);
nand U1409 (N_1409,N_1029,N_1025);
nor U1410 (N_1410,N_1061,N_1085);
nand U1411 (N_1411,N_1193,N_1209);
nor U1412 (N_1412,N_1136,N_1178);
nand U1413 (N_1413,N_1167,N_1090);
nor U1414 (N_1414,N_1179,N_1133);
nor U1415 (N_1415,N_1060,N_1075);
nand U1416 (N_1416,N_1176,N_1077);
or U1417 (N_1417,N_1227,N_1070);
nand U1418 (N_1418,N_1226,N_1172);
and U1419 (N_1419,N_1221,N_1006);
or U1420 (N_1420,N_1090,N_1191);
nand U1421 (N_1421,N_1111,N_1088);
nor U1422 (N_1422,N_1043,N_1157);
nand U1423 (N_1423,N_1149,N_1051);
nand U1424 (N_1424,N_1197,N_1207);
or U1425 (N_1425,N_1135,N_1195);
or U1426 (N_1426,N_1002,N_1248);
nor U1427 (N_1427,N_1045,N_1031);
and U1428 (N_1428,N_1045,N_1161);
or U1429 (N_1429,N_1011,N_1119);
nor U1430 (N_1430,N_1007,N_1186);
or U1431 (N_1431,N_1039,N_1215);
or U1432 (N_1432,N_1006,N_1141);
nand U1433 (N_1433,N_1053,N_1140);
nand U1434 (N_1434,N_1107,N_1227);
or U1435 (N_1435,N_1170,N_1161);
or U1436 (N_1436,N_1208,N_1014);
nor U1437 (N_1437,N_1160,N_1126);
xnor U1438 (N_1438,N_1051,N_1136);
nor U1439 (N_1439,N_1039,N_1154);
nand U1440 (N_1440,N_1024,N_1163);
nand U1441 (N_1441,N_1007,N_1236);
xnor U1442 (N_1442,N_1101,N_1194);
and U1443 (N_1443,N_1215,N_1047);
or U1444 (N_1444,N_1171,N_1186);
nor U1445 (N_1445,N_1111,N_1065);
and U1446 (N_1446,N_1210,N_1074);
nand U1447 (N_1447,N_1049,N_1132);
nand U1448 (N_1448,N_1021,N_1181);
xor U1449 (N_1449,N_1173,N_1066);
nor U1450 (N_1450,N_1245,N_1186);
or U1451 (N_1451,N_1149,N_1082);
xor U1452 (N_1452,N_1087,N_1216);
nor U1453 (N_1453,N_1223,N_1171);
nand U1454 (N_1454,N_1015,N_1042);
nand U1455 (N_1455,N_1070,N_1164);
nor U1456 (N_1456,N_1174,N_1223);
nor U1457 (N_1457,N_1158,N_1036);
and U1458 (N_1458,N_1169,N_1215);
nor U1459 (N_1459,N_1126,N_1083);
and U1460 (N_1460,N_1007,N_1044);
or U1461 (N_1461,N_1231,N_1109);
or U1462 (N_1462,N_1127,N_1088);
nand U1463 (N_1463,N_1082,N_1044);
or U1464 (N_1464,N_1215,N_1076);
and U1465 (N_1465,N_1033,N_1013);
or U1466 (N_1466,N_1079,N_1143);
and U1467 (N_1467,N_1030,N_1231);
and U1468 (N_1468,N_1158,N_1015);
xnor U1469 (N_1469,N_1240,N_1175);
nor U1470 (N_1470,N_1061,N_1087);
nor U1471 (N_1471,N_1216,N_1003);
and U1472 (N_1472,N_1166,N_1213);
nor U1473 (N_1473,N_1070,N_1031);
or U1474 (N_1474,N_1075,N_1081);
nor U1475 (N_1475,N_1143,N_1146);
nand U1476 (N_1476,N_1070,N_1101);
nor U1477 (N_1477,N_1220,N_1227);
and U1478 (N_1478,N_1167,N_1154);
and U1479 (N_1479,N_1075,N_1171);
xnor U1480 (N_1480,N_1090,N_1069);
nand U1481 (N_1481,N_1033,N_1135);
and U1482 (N_1482,N_1202,N_1182);
or U1483 (N_1483,N_1183,N_1013);
nand U1484 (N_1484,N_1221,N_1101);
and U1485 (N_1485,N_1144,N_1115);
nand U1486 (N_1486,N_1095,N_1244);
nor U1487 (N_1487,N_1168,N_1052);
xor U1488 (N_1488,N_1191,N_1228);
or U1489 (N_1489,N_1006,N_1043);
and U1490 (N_1490,N_1192,N_1162);
or U1491 (N_1491,N_1192,N_1153);
and U1492 (N_1492,N_1078,N_1184);
and U1493 (N_1493,N_1034,N_1096);
and U1494 (N_1494,N_1084,N_1165);
or U1495 (N_1495,N_1087,N_1011);
xnor U1496 (N_1496,N_1169,N_1107);
nand U1497 (N_1497,N_1244,N_1249);
and U1498 (N_1498,N_1112,N_1018);
nand U1499 (N_1499,N_1227,N_1076);
or U1500 (N_1500,N_1293,N_1435);
xor U1501 (N_1501,N_1420,N_1391);
nand U1502 (N_1502,N_1408,N_1275);
nand U1503 (N_1503,N_1307,N_1333);
nor U1504 (N_1504,N_1447,N_1319);
nand U1505 (N_1505,N_1364,N_1350);
nand U1506 (N_1506,N_1268,N_1273);
nand U1507 (N_1507,N_1424,N_1394);
or U1508 (N_1508,N_1474,N_1372);
or U1509 (N_1509,N_1277,N_1462);
and U1510 (N_1510,N_1499,N_1310);
or U1511 (N_1511,N_1254,N_1423);
nand U1512 (N_1512,N_1495,N_1317);
nand U1513 (N_1513,N_1450,N_1296);
or U1514 (N_1514,N_1329,N_1303);
nor U1515 (N_1515,N_1363,N_1376);
or U1516 (N_1516,N_1266,N_1458);
or U1517 (N_1517,N_1430,N_1467);
nor U1518 (N_1518,N_1460,N_1416);
and U1519 (N_1519,N_1417,N_1475);
and U1520 (N_1520,N_1481,N_1491);
nor U1521 (N_1521,N_1308,N_1335);
and U1522 (N_1522,N_1353,N_1461);
or U1523 (N_1523,N_1356,N_1494);
and U1524 (N_1524,N_1334,N_1316);
and U1525 (N_1525,N_1401,N_1337);
xor U1526 (N_1526,N_1385,N_1397);
and U1527 (N_1527,N_1471,N_1270);
and U1528 (N_1528,N_1252,N_1441);
or U1529 (N_1529,N_1330,N_1369);
or U1530 (N_1530,N_1428,N_1290);
and U1531 (N_1531,N_1298,N_1351);
nor U1532 (N_1532,N_1287,N_1341);
nor U1533 (N_1533,N_1285,N_1378);
nand U1534 (N_1534,N_1406,N_1279);
nor U1535 (N_1535,N_1263,N_1429);
nor U1536 (N_1536,N_1312,N_1257);
xnor U1537 (N_1537,N_1325,N_1414);
nor U1538 (N_1538,N_1465,N_1468);
and U1539 (N_1539,N_1473,N_1343);
or U1540 (N_1540,N_1313,N_1269);
nor U1541 (N_1541,N_1304,N_1284);
and U1542 (N_1542,N_1448,N_1379);
and U1543 (N_1543,N_1432,N_1340);
xnor U1544 (N_1544,N_1410,N_1311);
nor U1545 (N_1545,N_1281,N_1452);
nand U1546 (N_1546,N_1360,N_1347);
or U1547 (N_1547,N_1256,N_1455);
or U1548 (N_1548,N_1274,N_1265);
nor U1549 (N_1549,N_1282,N_1342);
nor U1550 (N_1550,N_1404,N_1331);
and U1551 (N_1551,N_1492,N_1396);
xor U1552 (N_1552,N_1482,N_1431);
nand U1553 (N_1553,N_1449,N_1453);
nor U1554 (N_1554,N_1288,N_1487);
nor U1555 (N_1555,N_1361,N_1387);
nor U1556 (N_1556,N_1426,N_1476);
and U1557 (N_1557,N_1382,N_1253);
nand U1558 (N_1558,N_1365,N_1358);
and U1559 (N_1559,N_1301,N_1261);
xnor U1560 (N_1560,N_1264,N_1291);
or U1561 (N_1561,N_1402,N_1255);
nor U1562 (N_1562,N_1251,N_1367);
nand U1563 (N_1563,N_1464,N_1392);
nand U1564 (N_1564,N_1393,N_1366);
or U1565 (N_1565,N_1444,N_1490);
nand U1566 (N_1566,N_1403,N_1456);
and U1567 (N_1567,N_1442,N_1496);
nand U1568 (N_1568,N_1321,N_1434);
and U1569 (N_1569,N_1322,N_1383);
xnor U1570 (N_1570,N_1346,N_1297);
or U1571 (N_1571,N_1348,N_1418);
nor U1572 (N_1572,N_1259,N_1271);
nand U1573 (N_1573,N_1286,N_1421);
nand U1574 (N_1574,N_1498,N_1489);
nand U1575 (N_1575,N_1479,N_1381);
nand U1576 (N_1576,N_1294,N_1370);
or U1577 (N_1577,N_1437,N_1422);
and U1578 (N_1578,N_1445,N_1354);
nor U1579 (N_1579,N_1493,N_1440);
nand U1580 (N_1580,N_1446,N_1349);
nand U1581 (N_1581,N_1338,N_1405);
xnor U1582 (N_1582,N_1413,N_1332);
xor U1583 (N_1583,N_1438,N_1262);
or U1584 (N_1584,N_1436,N_1357);
and U1585 (N_1585,N_1400,N_1485);
and U1586 (N_1586,N_1427,N_1336);
nand U1587 (N_1587,N_1466,N_1272);
nor U1588 (N_1588,N_1425,N_1314);
or U1589 (N_1589,N_1362,N_1457);
nor U1590 (N_1590,N_1386,N_1326);
or U1591 (N_1591,N_1368,N_1384);
or U1592 (N_1592,N_1483,N_1486);
or U1593 (N_1593,N_1407,N_1480);
or U1594 (N_1594,N_1377,N_1345);
nand U1595 (N_1595,N_1451,N_1328);
or U1596 (N_1596,N_1389,N_1344);
nand U1597 (N_1597,N_1470,N_1339);
nand U1598 (N_1598,N_1373,N_1419);
xor U1599 (N_1599,N_1409,N_1412);
and U1600 (N_1600,N_1250,N_1305);
nand U1601 (N_1601,N_1497,N_1359);
xor U1602 (N_1602,N_1463,N_1380);
nand U1603 (N_1603,N_1260,N_1478);
nand U1604 (N_1604,N_1472,N_1374);
nor U1605 (N_1605,N_1302,N_1267);
or U1606 (N_1606,N_1280,N_1283);
and U1607 (N_1607,N_1390,N_1411);
xnor U1608 (N_1608,N_1352,N_1299);
and U1609 (N_1609,N_1318,N_1433);
nand U1610 (N_1610,N_1323,N_1324);
or U1611 (N_1611,N_1309,N_1399);
or U1612 (N_1612,N_1477,N_1375);
and U1613 (N_1613,N_1300,N_1355);
nor U1614 (N_1614,N_1315,N_1398);
or U1615 (N_1615,N_1295,N_1258);
xor U1616 (N_1616,N_1289,N_1292);
and U1617 (N_1617,N_1454,N_1439);
nand U1618 (N_1618,N_1327,N_1388);
or U1619 (N_1619,N_1371,N_1469);
and U1620 (N_1620,N_1278,N_1415);
and U1621 (N_1621,N_1276,N_1459);
and U1622 (N_1622,N_1395,N_1484);
nand U1623 (N_1623,N_1443,N_1320);
and U1624 (N_1624,N_1306,N_1488);
nor U1625 (N_1625,N_1324,N_1489);
nand U1626 (N_1626,N_1436,N_1301);
nand U1627 (N_1627,N_1279,N_1487);
or U1628 (N_1628,N_1384,N_1408);
and U1629 (N_1629,N_1392,N_1356);
nand U1630 (N_1630,N_1414,N_1317);
nand U1631 (N_1631,N_1371,N_1432);
or U1632 (N_1632,N_1412,N_1408);
or U1633 (N_1633,N_1320,N_1264);
or U1634 (N_1634,N_1455,N_1435);
nor U1635 (N_1635,N_1415,N_1462);
or U1636 (N_1636,N_1286,N_1352);
nand U1637 (N_1637,N_1255,N_1269);
and U1638 (N_1638,N_1289,N_1474);
nand U1639 (N_1639,N_1284,N_1476);
nor U1640 (N_1640,N_1326,N_1413);
nand U1641 (N_1641,N_1296,N_1323);
nor U1642 (N_1642,N_1333,N_1448);
and U1643 (N_1643,N_1488,N_1391);
and U1644 (N_1644,N_1342,N_1269);
nor U1645 (N_1645,N_1362,N_1435);
or U1646 (N_1646,N_1374,N_1417);
nand U1647 (N_1647,N_1256,N_1420);
or U1648 (N_1648,N_1339,N_1420);
xnor U1649 (N_1649,N_1444,N_1466);
or U1650 (N_1650,N_1387,N_1381);
nor U1651 (N_1651,N_1361,N_1438);
nand U1652 (N_1652,N_1395,N_1341);
and U1653 (N_1653,N_1309,N_1331);
xnor U1654 (N_1654,N_1271,N_1276);
nor U1655 (N_1655,N_1259,N_1474);
or U1656 (N_1656,N_1413,N_1433);
and U1657 (N_1657,N_1394,N_1311);
and U1658 (N_1658,N_1291,N_1306);
nor U1659 (N_1659,N_1261,N_1365);
nor U1660 (N_1660,N_1448,N_1490);
nor U1661 (N_1661,N_1467,N_1282);
or U1662 (N_1662,N_1445,N_1417);
nor U1663 (N_1663,N_1300,N_1354);
or U1664 (N_1664,N_1287,N_1397);
nor U1665 (N_1665,N_1471,N_1399);
nor U1666 (N_1666,N_1458,N_1281);
or U1667 (N_1667,N_1295,N_1366);
and U1668 (N_1668,N_1493,N_1403);
or U1669 (N_1669,N_1438,N_1314);
and U1670 (N_1670,N_1395,N_1467);
nor U1671 (N_1671,N_1352,N_1450);
nand U1672 (N_1672,N_1315,N_1444);
nand U1673 (N_1673,N_1297,N_1381);
nand U1674 (N_1674,N_1337,N_1378);
or U1675 (N_1675,N_1309,N_1420);
or U1676 (N_1676,N_1405,N_1445);
nor U1677 (N_1677,N_1358,N_1272);
nand U1678 (N_1678,N_1480,N_1351);
nand U1679 (N_1679,N_1277,N_1499);
nor U1680 (N_1680,N_1438,N_1380);
nand U1681 (N_1681,N_1286,N_1314);
nand U1682 (N_1682,N_1481,N_1288);
xnor U1683 (N_1683,N_1330,N_1340);
or U1684 (N_1684,N_1299,N_1486);
nor U1685 (N_1685,N_1323,N_1368);
and U1686 (N_1686,N_1315,N_1272);
nor U1687 (N_1687,N_1439,N_1448);
and U1688 (N_1688,N_1426,N_1367);
nor U1689 (N_1689,N_1453,N_1330);
nor U1690 (N_1690,N_1298,N_1255);
and U1691 (N_1691,N_1282,N_1357);
nand U1692 (N_1692,N_1330,N_1423);
nand U1693 (N_1693,N_1370,N_1345);
or U1694 (N_1694,N_1370,N_1469);
nor U1695 (N_1695,N_1363,N_1408);
nor U1696 (N_1696,N_1357,N_1368);
xor U1697 (N_1697,N_1268,N_1480);
and U1698 (N_1698,N_1300,N_1399);
nor U1699 (N_1699,N_1288,N_1252);
or U1700 (N_1700,N_1276,N_1283);
or U1701 (N_1701,N_1283,N_1474);
nor U1702 (N_1702,N_1256,N_1396);
or U1703 (N_1703,N_1491,N_1447);
xor U1704 (N_1704,N_1374,N_1428);
nand U1705 (N_1705,N_1331,N_1365);
or U1706 (N_1706,N_1361,N_1318);
nand U1707 (N_1707,N_1289,N_1443);
or U1708 (N_1708,N_1333,N_1499);
or U1709 (N_1709,N_1353,N_1291);
and U1710 (N_1710,N_1486,N_1325);
xor U1711 (N_1711,N_1328,N_1353);
and U1712 (N_1712,N_1331,N_1440);
xnor U1713 (N_1713,N_1338,N_1394);
and U1714 (N_1714,N_1421,N_1471);
and U1715 (N_1715,N_1301,N_1351);
nand U1716 (N_1716,N_1384,N_1366);
and U1717 (N_1717,N_1496,N_1484);
and U1718 (N_1718,N_1482,N_1310);
or U1719 (N_1719,N_1291,N_1315);
or U1720 (N_1720,N_1469,N_1428);
nor U1721 (N_1721,N_1384,N_1397);
and U1722 (N_1722,N_1274,N_1257);
or U1723 (N_1723,N_1334,N_1359);
or U1724 (N_1724,N_1495,N_1309);
or U1725 (N_1725,N_1404,N_1327);
nor U1726 (N_1726,N_1406,N_1395);
or U1727 (N_1727,N_1294,N_1490);
or U1728 (N_1728,N_1459,N_1429);
nor U1729 (N_1729,N_1466,N_1454);
or U1730 (N_1730,N_1458,N_1252);
nand U1731 (N_1731,N_1490,N_1461);
xor U1732 (N_1732,N_1250,N_1257);
nand U1733 (N_1733,N_1402,N_1373);
nor U1734 (N_1734,N_1317,N_1310);
and U1735 (N_1735,N_1353,N_1336);
and U1736 (N_1736,N_1494,N_1368);
and U1737 (N_1737,N_1447,N_1480);
nand U1738 (N_1738,N_1446,N_1318);
or U1739 (N_1739,N_1349,N_1357);
or U1740 (N_1740,N_1396,N_1411);
nor U1741 (N_1741,N_1420,N_1492);
nand U1742 (N_1742,N_1411,N_1296);
nand U1743 (N_1743,N_1458,N_1342);
and U1744 (N_1744,N_1304,N_1407);
nand U1745 (N_1745,N_1391,N_1442);
and U1746 (N_1746,N_1334,N_1366);
nor U1747 (N_1747,N_1395,N_1460);
nor U1748 (N_1748,N_1342,N_1316);
or U1749 (N_1749,N_1400,N_1429);
nor U1750 (N_1750,N_1685,N_1740);
nor U1751 (N_1751,N_1733,N_1594);
nor U1752 (N_1752,N_1708,N_1659);
nand U1753 (N_1753,N_1695,N_1686);
or U1754 (N_1754,N_1619,N_1622);
nor U1755 (N_1755,N_1613,N_1720);
nor U1756 (N_1756,N_1543,N_1743);
or U1757 (N_1757,N_1724,N_1616);
nand U1758 (N_1758,N_1649,N_1610);
nand U1759 (N_1759,N_1676,N_1634);
or U1760 (N_1760,N_1564,N_1711);
and U1761 (N_1761,N_1520,N_1660);
or U1762 (N_1762,N_1651,N_1555);
nor U1763 (N_1763,N_1525,N_1705);
nand U1764 (N_1764,N_1746,N_1575);
and U1765 (N_1765,N_1584,N_1748);
nor U1766 (N_1766,N_1508,N_1742);
and U1767 (N_1767,N_1657,N_1745);
and U1768 (N_1768,N_1551,N_1603);
nor U1769 (N_1769,N_1547,N_1532);
or U1770 (N_1770,N_1704,N_1537);
nand U1771 (N_1771,N_1557,N_1702);
xnor U1772 (N_1772,N_1553,N_1572);
xor U1773 (N_1773,N_1739,N_1530);
nor U1774 (N_1774,N_1735,N_1672);
or U1775 (N_1775,N_1527,N_1599);
nand U1776 (N_1776,N_1524,N_1573);
and U1777 (N_1777,N_1630,N_1717);
xor U1778 (N_1778,N_1697,N_1500);
nor U1779 (N_1779,N_1747,N_1604);
or U1780 (N_1780,N_1552,N_1533);
or U1781 (N_1781,N_1511,N_1669);
or U1782 (N_1782,N_1693,N_1648);
nor U1783 (N_1783,N_1519,N_1692);
and U1784 (N_1784,N_1698,N_1640);
nand U1785 (N_1785,N_1600,N_1545);
nand U1786 (N_1786,N_1618,N_1569);
xnor U1787 (N_1787,N_1558,N_1510);
xor U1788 (N_1788,N_1606,N_1609);
nand U1789 (N_1789,N_1621,N_1503);
and U1790 (N_1790,N_1658,N_1666);
nor U1791 (N_1791,N_1561,N_1540);
nor U1792 (N_1792,N_1614,N_1699);
and U1793 (N_1793,N_1712,N_1586);
nand U1794 (N_1794,N_1624,N_1568);
or U1795 (N_1795,N_1722,N_1576);
or U1796 (N_1796,N_1738,N_1516);
nand U1797 (N_1797,N_1668,N_1680);
and U1798 (N_1798,N_1522,N_1515);
and U1799 (N_1799,N_1591,N_1637);
nand U1800 (N_1800,N_1579,N_1694);
xnor U1801 (N_1801,N_1647,N_1571);
or U1802 (N_1802,N_1662,N_1677);
and U1803 (N_1803,N_1546,N_1736);
or U1804 (N_1804,N_1653,N_1675);
and U1805 (N_1805,N_1732,N_1727);
nor U1806 (N_1806,N_1534,N_1631);
nor U1807 (N_1807,N_1663,N_1531);
or U1808 (N_1808,N_1679,N_1623);
nand U1809 (N_1809,N_1521,N_1731);
and U1810 (N_1810,N_1726,N_1718);
xnor U1811 (N_1811,N_1517,N_1501);
and U1812 (N_1812,N_1667,N_1544);
nor U1813 (N_1813,N_1581,N_1707);
and U1814 (N_1814,N_1741,N_1556);
xor U1815 (N_1815,N_1696,N_1691);
nand U1816 (N_1816,N_1504,N_1636);
and U1817 (N_1817,N_1585,N_1681);
and U1818 (N_1818,N_1567,N_1593);
nand U1819 (N_1819,N_1639,N_1628);
or U1820 (N_1820,N_1719,N_1526);
nor U1821 (N_1821,N_1749,N_1563);
and U1822 (N_1822,N_1588,N_1554);
nand U1823 (N_1823,N_1528,N_1656);
nor U1824 (N_1824,N_1661,N_1690);
and U1825 (N_1825,N_1505,N_1645);
or U1826 (N_1826,N_1578,N_1629);
and U1827 (N_1827,N_1674,N_1678);
nor U1828 (N_1828,N_1650,N_1611);
and U1829 (N_1829,N_1509,N_1713);
and U1830 (N_1830,N_1598,N_1744);
or U1831 (N_1831,N_1632,N_1596);
and U1832 (N_1832,N_1577,N_1580);
nand U1833 (N_1833,N_1550,N_1682);
nor U1834 (N_1834,N_1587,N_1597);
nand U1835 (N_1835,N_1644,N_1673);
and U1836 (N_1836,N_1560,N_1723);
xnor U1837 (N_1837,N_1683,N_1626);
nand U1838 (N_1838,N_1684,N_1541);
and U1839 (N_1839,N_1716,N_1523);
nand U1840 (N_1840,N_1607,N_1565);
and U1841 (N_1841,N_1595,N_1592);
nand U1842 (N_1842,N_1700,N_1703);
or U1843 (N_1843,N_1714,N_1506);
and U1844 (N_1844,N_1687,N_1670);
or U1845 (N_1845,N_1542,N_1652);
and U1846 (N_1846,N_1620,N_1518);
nand U1847 (N_1847,N_1734,N_1688);
or U1848 (N_1848,N_1548,N_1725);
xnor U1849 (N_1849,N_1602,N_1665);
nand U1850 (N_1850,N_1709,N_1538);
nor U1851 (N_1851,N_1605,N_1589);
nor U1852 (N_1852,N_1625,N_1617);
or U1853 (N_1853,N_1549,N_1706);
nor U1854 (N_1854,N_1721,N_1701);
nor U1855 (N_1855,N_1566,N_1627);
or U1856 (N_1856,N_1562,N_1671);
and U1857 (N_1857,N_1583,N_1514);
nor U1858 (N_1858,N_1582,N_1728);
nor U1859 (N_1859,N_1633,N_1737);
nor U1860 (N_1860,N_1641,N_1729);
and U1861 (N_1861,N_1730,N_1502);
nor U1862 (N_1862,N_1643,N_1536);
nand U1863 (N_1863,N_1512,N_1715);
xnor U1864 (N_1864,N_1601,N_1590);
and U1865 (N_1865,N_1529,N_1638);
nor U1866 (N_1866,N_1642,N_1612);
nand U1867 (N_1867,N_1635,N_1539);
or U1868 (N_1868,N_1570,N_1655);
and U1869 (N_1869,N_1654,N_1535);
and U1870 (N_1870,N_1664,N_1513);
nand U1871 (N_1871,N_1689,N_1574);
nand U1872 (N_1872,N_1615,N_1608);
and U1873 (N_1873,N_1710,N_1646);
or U1874 (N_1874,N_1559,N_1507);
and U1875 (N_1875,N_1678,N_1625);
nand U1876 (N_1876,N_1707,N_1508);
xor U1877 (N_1877,N_1646,N_1601);
or U1878 (N_1878,N_1625,N_1662);
or U1879 (N_1879,N_1562,N_1527);
or U1880 (N_1880,N_1660,N_1746);
nand U1881 (N_1881,N_1737,N_1553);
or U1882 (N_1882,N_1674,N_1724);
and U1883 (N_1883,N_1593,N_1639);
nand U1884 (N_1884,N_1745,N_1524);
or U1885 (N_1885,N_1712,N_1572);
nand U1886 (N_1886,N_1625,N_1594);
or U1887 (N_1887,N_1739,N_1596);
or U1888 (N_1888,N_1723,N_1543);
and U1889 (N_1889,N_1593,N_1535);
and U1890 (N_1890,N_1692,N_1689);
nor U1891 (N_1891,N_1558,N_1612);
nand U1892 (N_1892,N_1692,N_1503);
or U1893 (N_1893,N_1634,N_1603);
xnor U1894 (N_1894,N_1601,N_1700);
or U1895 (N_1895,N_1701,N_1723);
nor U1896 (N_1896,N_1749,N_1738);
nand U1897 (N_1897,N_1654,N_1716);
xor U1898 (N_1898,N_1747,N_1570);
or U1899 (N_1899,N_1581,N_1702);
and U1900 (N_1900,N_1748,N_1736);
xnor U1901 (N_1901,N_1528,N_1705);
and U1902 (N_1902,N_1690,N_1509);
or U1903 (N_1903,N_1664,N_1702);
nor U1904 (N_1904,N_1612,N_1702);
nand U1905 (N_1905,N_1658,N_1586);
nand U1906 (N_1906,N_1594,N_1612);
and U1907 (N_1907,N_1724,N_1667);
nor U1908 (N_1908,N_1509,N_1595);
nand U1909 (N_1909,N_1668,N_1622);
nor U1910 (N_1910,N_1590,N_1562);
nand U1911 (N_1911,N_1684,N_1688);
and U1912 (N_1912,N_1704,N_1688);
nor U1913 (N_1913,N_1725,N_1563);
nand U1914 (N_1914,N_1518,N_1562);
or U1915 (N_1915,N_1673,N_1523);
and U1916 (N_1916,N_1672,N_1597);
nand U1917 (N_1917,N_1603,N_1591);
nand U1918 (N_1918,N_1650,N_1636);
and U1919 (N_1919,N_1613,N_1623);
nand U1920 (N_1920,N_1727,N_1578);
nor U1921 (N_1921,N_1593,N_1671);
nand U1922 (N_1922,N_1678,N_1655);
or U1923 (N_1923,N_1527,N_1583);
or U1924 (N_1924,N_1575,N_1727);
nor U1925 (N_1925,N_1725,N_1732);
nor U1926 (N_1926,N_1710,N_1614);
nor U1927 (N_1927,N_1642,N_1631);
or U1928 (N_1928,N_1539,N_1722);
nand U1929 (N_1929,N_1683,N_1706);
nand U1930 (N_1930,N_1721,N_1707);
nor U1931 (N_1931,N_1583,N_1651);
xor U1932 (N_1932,N_1607,N_1559);
nand U1933 (N_1933,N_1705,N_1520);
and U1934 (N_1934,N_1732,N_1684);
xor U1935 (N_1935,N_1506,N_1699);
or U1936 (N_1936,N_1691,N_1563);
and U1937 (N_1937,N_1537,N_1547);
and U1938 (N_1938,N_1653,N_1656);
nor U1939 (N_1939,N_1624,N_1704);
nor U1940 (N_1940,N_1705,N_1652);
or U1941 (N_1941,N_1706,N_1558);
and U1942 (N_1942,N_1518,N_1741);
nand U1943 (N_1943,N_1749,N_1621);
nor U1944 (N_1944,N_1529,N_1583);
and U1945 (N_1945,N_1713,N_1661);
nor U1946 (N_1946,N_1610,N_1709);
and U1947 (N_1947,N_1635,N_1595);
nand U1948 (N_1948,N_1605,N_1730);
or U1949 (N_1949,N_1635,N_1515);
xnor U1950 (N_1950,N_1658,N_1623);
and U1951 (N_1951,N_1676,N_1586);
nor U1952 (N_1952,N_1714,N_1533);
nor U1953 (N_1953,N_1533,N_1549);
nor U1954 (N_1954,N_1518,N_1632);
nand U1955 (N_1955,N_1551,N_1724);
and U1956 (N_1956,N_1677,N_1521);
and U1957 (N_1957,N_1667,N_1524);
and U1958 (N_1958,N_1619,N_1692);
or U1959 (N_1959,N_1698,N_1537);
nor U1960 (N_1960,N_1685,N_1627);
nor U1961 (N_1961,N_1741,N_1662);
or U1962 (N_1962,N_1697,N_1730);
or U1963 (N_1963,N_1669,N_1528);
nor U1964 (N_1964,N_1736,N_1596);
and U1965 (N_1965,N_1524,N_1673);
nand U1966 (N_1966,N_1514,N_1591);
xnor U1967 (N_1967,N_1694,N_1710);
nor U1968 (N_1968,N_1594,N_1646);
and U1969 (N_1969,N_1666,N_1660);
xnor U1970 (N_1970,N_1607,N_1537);
and U1971 (N_1971,N_1632,N_1507);
xnor U1972 (N_1972,N_1558,N_1712);
and U1973 (N_1973,N_1701,N_1747);
xor U1974 (N_1974,N_1543,N_1691);
nor U1975 (N_1975,N_1548,N_1554);
or U1976 (N_1976,N_1715,N_1500);
nand U1977 (N_1977,N_1576,N_1716);
nand U1978 (N_1978,N_1516,N_1611);
nand U1979 (N_1979,N_1671,N_1640);
and U1980 (N_1980,N_1671,N_1745);
xor U1981 (N_1981,N_1707,N_1596);
nand U1982 (N_1982,N_1515,N_1736);
xnor U1983 (N_1983,N_1661,N_1554);
or U1984 (N_1984,N_1573,N_1727);
and U1985 (N_1985,N_1523,N_1607);
nand U1986 (N_1986,N_1544,N_1523);
nand U1987 (N_1987,N_1678,N_1518);
and U1988 (N_1988,N_1747,N_1510);
or U1989 (N_1989,N_1647,N_1589);
xnor U1990 (N_1990,N_1673,N_1742);
or U1991 (N_1991,N_1635,N_1656);
and U1992 (N_1992,N_1561,N_1710);
nand U1993 (N_1993,N_1718,N_1639);
or U1994 (N_1994,N_1690,N_1601);
or U1995 (N_1995,N_1640,N_1572);
nor U1996 (N_1996,N_1663,N_1677);
nor U1997 (N_1997,N_1699,N_1552);
nand U1998 (N_1998,N_1709,N_1735);
and U1999 (N_1999,N_1552,N_1702);
or U2000 (N_2000,N_1916,N_1866);
or U2001 (N_2001,N_1774,N_1845);
nand U2002 (N_2002,N_1940,N_1964);
and U2003 (N_2003,N_1911,N_1891);
or U2004 (N_2004,N_1989,N_1987);
nand U2005 (N_2005,N_1763,N_1859);
nand U2006 (N_2006,N_1840,N_1848);
nor U2007 (N_2007,N_1949,N_1929);
or U2008 (N_2008,N_1927,N_1833);
nand U2009 (N_2009,N_1938,N_1985);
and U2010 (N_2010,N_1800,N_1978);
nand U2011 (N_2011,N_1808,N_1956);
and U2012 (N_2012,N_1856,N_1770);
or U2013 (N_2013,N_1829,N_1977);
nand U2014 (N_2014,N_1996,N_1967);
or U2015 (N_2015,N_1832,N_1971);
xor U2016 (N_2016,N_1999,N_1926);
xnor U2017 (N_2017,N_1823,N_1753);
nor U2018 (N_2018,N_1993,N_1904);
or U2019 (N_2019,N_1819,N_1909);
nand U2020 (N_2020,N_1941,N_1895);
nand U2021 (N_2021,N_1902,N_1947);
xnor U2022 (N_2022,N_1908,N_1882);
nor U2023 (N_2023,N_1771,N_1836);
nand U2024 (N_2024,N_1750,N_1870);
and U2025 (N_2025,N_1953,N_1806);
nand U2026 (N_2026,N_1835,N_1874);
nor U2027 (N_2027,N_1849,N_1959);
nand U2028 (N_2028,N_1883,N_1915);
xnor U2029 (N_2029,N_1762,N_1755);
nand U2030 (N_2030,N_1852,N_1963);
or U2031 (N_2031,N_1888,N_1944);
and U2032 (N_2032,N_1983,N_1863);
or U2033 (N_2033,N_1919,N_1776);
nand U2034 (N_2034,N_1816,N_1864);
nand U2035 (N_2035,N_1758,N_1751);
or U2036 (N_2036,N_1943,N_1799);
and U2037 (N_2037,N_1998,N_1962);
nor U2038 (N_2038,N_1754,N_1934);
nor U2039 (N_2039,N_1980,N_1855);
or U2040 (N_2040,N_1769,N_1752);
or U2041 (N_2041,N_1905,N_1767);
nand U2042 (N_2042,N_1955,N_1928);
and U2043 (N_2043,N_1844,N_1890);
or U2044 (N_2044,N_1778,N_1777);
and U2045 (N_2045,N_1913,N_1860);
xor U2046 (N_2046,N_1906,N_1981);
xor U2047 (N_2047,N_1807,N_1781);
and U2048 (N_2048,N_1881,N_1923);
nand U2049 (N_2049,N_1968,N_1954);
nor U2050 (N_2050,N_1804,N_1990);
and U2051 (N_2051,N_1847,N_1970);
nor U2052 (N_2052,N_1851,N_1825);
nand U2053 (N_2053,N_1957,N_1795);
and U2054 (N_2054,N_1810,N_1939);
nand U2055 (N_2055,N_1850,N_1995);
and U2056 (N_2056,N_1988,N_1910);
nand U2057 (N_2057,N_1924,N_1885);
nand U2058 (N_2058,N_1986,N_1871);
and U2059 (N_2059,N_1936,N_1805);
and U2060 (N_2060,N_1787,N_1812);
or U2061 (N_2061,N_1857,N_1876);
nand U2062 (N_2062,N_1868,N_1821);
xor U2063 (N_2063,N_1946,N_1893);
nand U2064 (N_2064,N_1786,N_1764);
nand U2065 (N_2065,N_1775,N_1780);
nor U2066 (N_2066,N_1950,N_1854);
nor U2067 (N_2067,N_1896,N_1969);
or U2068 (N_2068,N_1912,N_1958);
nor U2069 (N_2069,N_1965,N_1788);
nor U2070 (N_2070,N_1772,N_1984);
and U2071 (N_2071,N_1793,N_1921);
and U2072 (N_2072,N_1820,N_1900);
nor U2073 (N_2073,N_1817,N_1815);
xor U2074 (N_2074,N_1875,N_1973);
xnor U2075 (N_2075,N_1846,N_1801);
and U2076 (N_2076,N_1917,N_1994);
nand U2077 (N_2077,N_1878,N_1975);
nand U2078 (N_2078,N_1794,N_1858);
or U2079 (N_2079,N_1822,N_1879);
or U2080 (N_2080,N_1797,N_1757);
nand U2081 (N_2081,N_1952,N_1861);
nor U2082 (N_2082,N_1897,N_1785);
nor U2083 (N_2083,N_1792,N_1789);
or U2084 (N_2084,N_1831,N_1841);
xor U2085 (N_2085,N_1997,N_1782);
nand U2086 (N_2086,N_1826,N_1925);
nor U2087 (N_2087,N_1843,N_1880);
and U2088 (N_2088,N_1894,N_1867);
nor U2089 (N_2089,N_1920,N_1982);
and U2090 (N_2090,N_1948,N_1979);
nor U2091 (N_2091,N_1760,N_1872);
nand U2092 (N_2092,N_1828,N_1813);
and U2093 (N_2093,N_1937,N_1930);
or U2094 (N_2094,N_1759,N_1803);
nor U2095 (N_2095,N_1898,N_1918);
nand U2096 (N_2096,N_1837,N_1842);
nand U2097 (N_2097,N_1884,N_1756);
xnor U2098 (N_2098,N_1922,N_1818);
nand U2099 (N_2099,N_1935,N_1853);
nand U2100 (N_2100,N_1903,N_1783);
and U2101 (N_2101,N_1838,N_1877);
nand U2102 (N_2102,N_1830,N_1886);
and U2103 (N_2103,N_1972,N_1798);
and U2104 (N_2104,N_1889,N_1765);
nor U2105 (N_2105,N_1768,N_1761);
nand U2106 (N_2106,N_1892,N_1960);
xnor U2107 (N_2107,N_1991,N_1976);
xnor U2108 (N_2108,N_1961,N_1796);
nor U2109 (N_2109,N_1824,N_1790);
nor U2110 (N_2110,N_1933,N_1784);
and U2111 (N_2111,N_1814,N_1773);
xor U2112 (N_2112,N_1899,N_1914);
or U2113 (N_2113,N_1827,N_1945);
nand U2114 (N_2114,N_1809,N_1931);
or U2115 (N_2115,N_1873,N_1869);
or U2116 (N_2116,N_1865,N_1802);
nor U2117 (N_2117,N_1942,N_1839);
nand U2118 (N_2118,N_1966,N_1834);
nand U2119 (N_2119,N_1974,N_1811);
or U2120 (N_2120,N_1887,N_1901);
or U2121 (N_2121,N_1992,N_1932);
nand U2122 (N_2122,N_1779,N_1862);
or U2123 (N_2123,N_1907,N_1766);
nand U2124 (N_2124,N_1791,N_1951);
xor U2125 (N_2125,N_1979,N_1905);
nor U2126 (N_2126,N_1828,N_1877);
nor U2127 (N_2127,N_1842,N_1812);
xor U2128 (N_2128,N_1792,N_1825);
nand U2129 (N_2129,N_1985,N_1875);
nand U2130 (N_2130,N_1931,N_1805);
and U2131 (N_2131,N_1851,N_1786);
nand U2132 (N_2132,N_1993,N_1767);
nand U2133 (N_2133,N_1982,N_1973);
nand U2134 (N_2134,N_1883,N_1770);
and U2135 (N_2135,N_1920,N_1932);
nor U2136 (N_2136,N_1797,N_1998);
or U2137 (N_2137,N_1886,N_1776);
nor U2138 (N_2138,N_1754,N_1971);
nor U2139 (N_2139,N_1801,N_1900);
or U2140 (N_2140,N_1977,N_1763);
xor U2141 (N_2141,N_1934,N_1933);
nor U2142 (N_2142,N_1759,N_1964);
nand U2143 (N_2143,N_1905,N_1930);
and U2144 (N_2144,N_1934,N_1889);
nand U2145 (N_2145,N_1813,N_1873);
nor U2146 (N_2146,N_1753,N_1992);
nand U2147 (N_2147,N_1826,N_1995);
xnor U2148 (N_2148,N_1839,N_1890);
nor U2149 (N_2149,N_1871,N_1940);
or U2150 (N_2150,N_1847,N_1885);
nor U2151 (N_2151,N_1771,N_1892);
nand U2152 (N_2152,N_1834,N_1816);
xnor U2153 (N_2153,N_1932,N_1769);
nor U2154 (N_2154,N_1826,N_1768);
or U2155 (N_2155,N_1968,N_1782);
nor U2156 (N_2156,N_1901,N_1912);
xor U2157 (N_2157,N_1970,N_1894);
xor U2158 (N_2158,N_1752,N_1845);
nand U2159 (N_2159,N_1973,N_1933);
and U2160 (N_2160,N_1875,N_1900);
and U2161 (N_2161,N_1991,N_1982);
xnor U2162 (N_2162,N_1849,N_1762);
or U2163 (N_2163,N_1956,N_1992);
nand U2164 (N_2164,N_1833,N_1785);
xnor U2165 (N_2165,N_1957,N_1881);
xnor U2166 (N_2166,N_1862,N_1789);
and U2167 (N_2167,N_1962,N_1791);
nand U2168 (N_2168,N_1789,N_1807);
and U2169 (N_2169,N_1939,N_1797);
or U2170 (N_2170,N_1951,N_1974);
nor U2171 (N_2171,N_1960,N_1897);
nand U2172 (N_2172,N_1818,N_1905);
nand U2173 (N_2173,N_1880,N_1997);
or U2174 (N_2174,N_1806,N_1908);
nor U2175 (N_2175,N_1863,N_1962);
nor U2176 (N_2176,N_1869,N_1962);
and U2177 (N_2177,N_1965,N_1899);
nor U2178 (N_2178,N_1771,N_1891);
nor U2179 (N_2179,N_1967,N_1757);
or U2180 (N_2180,N_1855,N_1974);
nor U2181 (N_2181,N_1795,N_1806);
and U2182 (N_2182,N_1884,N_1893);
and U2183 (N_2183,N_1929,N_1809);
nand U2184 (N_2184,N_1984,N_1945);
xnor U2185 (N_2185,N_1879,N_1804);
nand U2186 (N_2186,N_1782,N_1897);
nand U2187 (N_2187,N_1816,N_1805);
nand U2188 (N_2188,N_1917,N_1940);
nand U2189 (N_2189,N_1815,N_1799);
nand U2190 (N_2190,N_1774,N_1854);
or U2191 (N_2191,N_1818,N_1877);
nand U2192 (N_2192,N_1979,N_1989);
or U2193 (N_2193,N_1842,N_1906);
or U2194 (N_2194,N_1774,N_1998);
nand U2195 (N_2195,N_1958,N_1927);
and U2196 (N_2196,N_1917,N_1944);
and U2197 (N_2197,N_1804,N_1943);
or U2198 (N_2198,N_1994,N_1784);
or U2199 (N_2199,N_1819,N_1817);
nand U2200 (N_2200,N_1797,N_1793);
nor U2201 (N_2201,N_1845,N_1884);
nand U2202 (N_2202,N_1829,N_1808);
and U2203 (N_2203,N_1814,N_1921);
nand U2204 (N_2204,N_1910,N_1857);
or U2205 (N_2205,N_1841,N_1797);
and U2206 (N_2206,N_1923,N_1911);
xnor U2207 (N_2207,N_1810,N_1906);
nand U2208 (N_2208,N_1842,N_1877);
and U2209 (N_2209,N_1991,N_1902);
nor U2210 (N_2210,N_1868,N_1808);
xor U2211 (N_2211,N_1846,N_1754);
and U2212 (N_2212,N_1947,N_1841);
and U2213 (N_2213,N_1874,N_1901);
nor U2214 (N_2214,N_1969,N_1895);
or U2215 (N_2215,N_1838,N_1804);
xnor U2216 (N_2216,N_1969,N_1848);
or U2217 (N_2217,N_1818,N_1970);
or U2218 (N_2218,N_1852,N_1967);
nor U2219 (N_2219,N_1768,N_1833);
or U2220 (N_2220,N_1794,N_1855);
xor U2221 (N_2221,N_1879,N_1779);
nand U2222 (N_2222,N_1780,N_1863);
xor U2223 (N_2223,N_1975,N_1804);
nor U2224 (N_2224,N_1949,N_1763);
or U2225 (N_2225,N_1793,N_1821);
and U2226 (N_2226,N_1761,N_1811);
nand U2227 (N_2227,N_1874,N_1999);
nor U2228 (N_2228,N_1825,N_1819);
nand U2229 (N_2229,N_1942,N_1830);
or U2230 (N_2230,N_1963,N_1817);
xnor U2231 (N_2231,N_1806,N_1901);
nor U2232 (N_2232,N_1817,N_1821);
or U2233 (N_2233,N_1885,N_1978);
xor U2234 (N_2234,N_1930,N_1754);
xor U2235 (N_2235,N_1921,N_1774);
and U2236 (N_2236,N_1916,N_1925);
nand U2237 (N_2237,N_1961,N_1791);
and U2238 (N_2238,N_1890,N_1919);
or U2239 (N_2239,N_1965,N_1874);
and U2240 (N_2240,N_1887,N_1998);
nand U2241 (N_2241,N_1962,N_1803);
and U2242 (N_2242,N_1924,N_1919);
xor U2243 (N_2243,N_1972,N_1996);
xnor U2244 (N_2244,N_1919,N_1953);
and U2245 (N_2245,N_1922,N_1973);
and U2246 (N_2246,N_1917,N_1999);
and U2247 (N_2247,N_1793,N_1829);
and U2248 (N_2248,N_1971,N_1884);
nor U2249 (N_2249,N_1906,N_1830);
xor U2250 (N_2250,N_2048,N_2060);
or U2251 (N_2251,N_2021,N_2025);
and U2252 (N_2252,N_2099,N_2180);
nand U2253 (N_2253,N_2136,N_2115);
nand U2254 (N_2254,N_2174,N_2065);
xnor U2255 (N_2255,N_2061,N_2028);
nand U2256 (N_2256,N_2244,N_2124);
or U2257 (N_2257,N_2153,N_2245);
nand U2258 (N_2258,N_2204,N_2077);
and U2259 (N_2259,N_2074,N_2046);
nor U2260 (N_2260,N_2004,N_2148);
nand U2261 (N_2261,N_2139,N_2181);
and U2262 (N_2262,N_2164,N_2083);
and U2263 (N_2263,N_2167,N_2135);
and U2264 (N_2264,N_2126,N_2159);
nor U2265 (N_2265,N_2178,N_2230);
nor U2266 (N_2266,N_2017,N_2149);
nor U2267 (N_2267,N_2201,N_2087);
nand U2268 (N_2268,N_2018,N_2224);
or U2269 (N_2269,N_2128,N_2014);
and U2270 (N_2270,N_2089,N_2005);
xor U2271 (N_2271,N_2160,N_2179);
and U2272 (N_2272,N_2214,N_2080);
and U2273 (N_2273,N_2229,N_2103);
xor U2274 (N_2274,N_2078,N_2073);
and U2275 (N_2275,N_2091,N_2225);
or U2276 (N_2276,N_2055,N_2098);
nand U2277 (N_2277,N_2079,N_2033);
or U2278 (N_2278,N_2234,N_2039);
and U2279 (N_2279,N_2247,N_2192);
xor U2280 (N_2280,N_2205,N_2050);
nand U2281 (N_2281,N_2209,N_2026);
nor U2282 (N_2282,N_2112,N_2152);
nand U2283 (N_2283,N_2047,N_2238);
nor U2284 (N_2284,N_2165,N_2030);
or U2285 (N_2285,N_2249,N_2236);
and U2286 (N_2286,N_2085,N_2027);
nor U2287 (N_2287,N_2000,N_2095);
xor U2288 (N_2288,N_2031,N_2189);
nand U2289 (N_2289,N_2243,N_2022);
nor U2290 (N_2290,N_2151,N_2187);
xor U2291 (N_2291,N_2125,N_2184);
nand U2292 (N_2292,N_2138,N_2067);
and U2293 (N_2293,N_2043,N_2196);
xor U2294 (N_2294,N_2239,N_2104);
and U2295 (N_2295,N_2131,N_2155);
nand U2296 (N_2296,N_2008,N_2037);
xor U2297 (N_2297,N_2010,N_2215);
or U2298 (N_2298,N_2158,N_2141);
and U2299 (N_2299,N_2146,N_2101);
nand U2300 (N_2300,N_2094,N_2009);
nand U2301 (N_2301,N_2032,N_2162);
or U2302 (N_2302,N_2070,N_2097);
and U2303 (N_2303,N_2102,N_2075);
nand U2304 (N_2304,N_2117,N_2210);
nand U2305 (N_2305,N_2202,N_2071);
and U2306 (N_2306,N_2206,N_2185);
or U2307 (N_2307,N_2182,N_2216);
nor U2308 (N_2308,N_2090,N_2049);
nand U2309 (N_2309,N_2203,N_2169);
xnor U2310 (N_2310,N_2121,N_2036);
xnor U2311 (N_2311,N_2110,N_2109);
or U2312 (N_2312,N_2147,N_2154);
or U2313 (N_2313,N_2093,N_2076);
nand U2314 (N_2314,N_2183,N_2016);
and U2315 (N_2315,N_2217,N_2198);
and U2316 (N_2316,N_2052,N_2246);
and U2317 (N_2317,N_2231,N_2233);
and U2318 (N_2318,N_2193,N_2173);
nor U2319 (N_2319,N_2175,N_2056);
or U2320 (N_2320,N_2199,N_2129);
nor U2321 (N_2321,N_2150,N_2156);
and U2322 (N_2322,N_2086,N_2140);
nor U2323 (N_2323,N_2145,N_2228);
and U2324 (N_2324,N_2059,N_2120);
nand U2325 (N_2325,N_2081,N_2096);
nand U2326 (N_2326,N_2044,N_2133);
or U2327 (N_2327,N_2134,N_2208);
or U2328 (N_2328,N_2137,N_2054);
nor U2329 (N_2329,N_2100,N_2114);
xnor U2330 (N_2330,N_2066,N_2069);
xnor U2331 (N_2331,N_2188,N_2132);
or U2332 (N_2332,N_2123,N_2002);
nand U2333 (N_2333,N_2003,N_2212);
nor U2334 (N_2334,N_2144,N_2237);
nand U2335 (N_2335,N_2088,N_2105);
nor U2336 (N_2336,N_2053,N_2219);
nand U2337 (N_2337,N_2045,N_2106);
nand U2338 (N_2338,N_2063,N_2040);
and U2339 (N_2339,N_2171,N_2191);
nor U2340 (N_2340,N_2057,N_2108);
nor U2341 (N_2341,N_2068,N_2197);
and U2342 (N_2342,N_2235,N_2242);
nand U2343 (N_2343,N_2195,N_2127);
and U2344 (N_2344,N_2023,N_2213);
xor U2345 (N_2345,N_2001,N_2062);
or U2346 (N_2346,N_2200,N_2220);
nor U2347 (N_2347,N_2051,N_2176);
and U2348 (N_2348,N_2006,N_2222);
or U2349 (N_2349,N_2194,N_2142);
or U2350 (N_2350,N_2227,N_2020);
xor U2351 (N_2351,N_2072,N_2107);
nand U2352 (N_2352,N_2172,N_2143);
or U2353 (N_2353,N_2011,N_2019);
and U2354 (N_2354,N_2012,N_2232);
nand U2355 (N_2355,N_2226,N_2240);
nor U2356 (N_2356,N_2161,N_2211);
or U2357 (N_2357,N_2118,N_2035);
or U2358 (N_2358,N_2163,N_2207);
or U2359 (N_2359,N_2166,N_2092);
or U2360 (N_2360,N_2058,N_2084);
xor U2361 (N_2361,N_2034,N_2015);
nand U2362 (N_2362,N_2130,N_2190);
or U2363 (N_2363,N_2218,N_2024);
xor U2364 (N_2364,N_2186,N_2241);
and U2365 (N_2365,N_2177,N_2038);
xor U2366 (N_2366,N_2157,N_2113);
or U2367 (N_2367,N_2064,N_2007);
or U2368 (N_2368,N_2029,N_2248);
nor U2369 (N_2369,N_2168,N_2042);
nand U2370 (N_2370,N_2119,N_2223);
and U2371 (N_2371,N_2170,N_2111);
nor U2372 (N_2372,N_2041,N_2082);
and U2373 (N_2373,N_2116,N_2013);
nor U2374 (N_2374,N_2122,N_2221);
or U2375 (N_2375,N_2150,N_2033);
nor U2376 (N_2376,N_2128,N_2045);
nor U2377 (N_2377,N_2082,N_2203);
nand U2378 (N_2378,N_2195,N_2188);
nand U2379 (N_2379,N_2010,N_2039);
and U2380 (N_2380,N_2216,N_2135);
xnor U2381 (N_2381,N_2036,N_2159);
and U2382 (N_2382,N_2010,N_2044);
or U2383 (N_2383,N_2032,N_2006);
xor U2384 (N_2384,N_2012,N_2024);
or U2385 (N_2385,N_2170,N_2032);
nand U2386 (N_2386,N_2053,N_2241);
nand U2387 (N_2387,N_2032,N_2187);
or U2388 (N_2388,N_2229,N_2243);
or U2389 (N_2389,N_2174,N_2090);
or U2390 (N_2390,N_2155,N_2161);
and U2391 (N_2391,N_2004,N_2131);
nor U2392 (N_2392,N_2208,N_2066);
or U2393 (N_2393,N_2123,N_2228);
nand U2394 (N_2394,N_2047,N_2148);
nor U2395 (N_2395,N_2217,N_2083);
nor U2396 (N_2396,N_2027,N_2019);
nor U2397 (N_2397,N_2085,N_2194);
nand U2398 (N_2398,N_2124,N_2206);
nand U2399 (N_2399,N_2169,N_2065);
nand U2400 (N_2400,N_2047,N_2034);
nor U2401 (N_2401,N_2118,N_2187);
nor U2402 (N_2402,N_2248,N_2067);
or U2403 (N_2403,N_2095,N_2033);
or U2404 (N_2404,N_2028,N_2071);
and U2405 (N_2405,N_2112,N_2059);
xor U2406 (N_2406,N_2149,N_2109);
and U2407 (N_2407,N_2078,N_2238);
or U2408 (N_2408,N_2148,N_2201);
nor U2409 (N_2409,N_2060,N_2155);
xor U2410 (N_2410,N_2027,N_2080);
xor U2411 (N_2411,N_2226,N_2113);
nor U2412 (N_2412,N_2228,N_2080);
and U2413 (N_2413,N_2247,N_2070);
nor U2414 (N_2414,N_2139,N_2125);
nor U2415 (N_2415,N_2123,N_2097);
nand U2416 (N_2416,N_2206,N_2014);
nor U2417 (N_2417,N_2146,N_2241);
or U2418 (N_2418,N_2183,N_2055);
nor U2419 (N_2419,N_2232,N_2216);
or U2420 (N_2420,N_2088,N_2033);
nand U2421 (N_2421,N_2018,N_2017);
nor U2422 (N_2422,N_2162,N_2046);
or U2423 (N_2423,N_2075,N_2100);
xor U2424 (N_2424,N_2066,N_2027);
and U2425 (N_2425,N_2138,N_2212);
and U2426 (N_2426,N_2174,N_2059);
or U2427 (N_2427,N_2078,N_2013);
and U2428 (N_2428,N_2175,N_2011);
xor U2429 (N_2429,N_2004,N_2169);
nor U2430 (N_2430,N_2247,N_2116);
nand U2431 (N_2431,N_2241,N_2205);
xnor U2432 (N_2432,N_2068,N_2180);
nor U2433 (N_2433,N_2049,N_2084);
nand U2434 (N_2434,N_2025,N_2148);
or U2435 (N_2435,N_2053,N_2000);
xor U2436 (N_2436,N_2009,N_2031);
xor U2437 (N_2437,N_2127,N_2062);
and U2438 (N_2438,N_2141,N_2049);
or U2439 (N_2439,N_2137,N_2123);
nand U2440 (N_2440,N_2167,N_2245);
xor U2441 (N_2441,N_2117,N_2229);
nand U2442 (N_2442,N_2125,N_2124);
nor U2443 (N_2443,N_2237,N_2108);
and U2444 (N_2444,N_2008,N_2124);
nor U2445 (N_2445,N_2031,N_2044);
nand U2446 (N_2446,N_2103,N_2110);
nand U2447 (N_2447,N_2171,N_2129);
or U2448 (N_2448,N_2182,N_2095);
or U2449 (N_2449,N_2178,N_2170);
nor U2450 (N_2450,N_2153,N_2143);
and U2451 (N_2451,N_2184,N_2105);
nand U2452 (N_2452,N_2011,N_2142);
nand U2453 (N_2453,N_2031,N_2242);
nand U2454 (N_2454,N_2149,N_2131);
and U2455 (N_2455,N_2207,N_2205);
nor U2456 (N_2456,N_2062,N_2081);
or U2457 (N_2457,N_2155,N_2040);
nand U2458 (N_2458,N_2195,N_2076);
and U2459 (N_2459,N_2171,N_2126);
and U2460 (N_2460,N_2142,N_2064);
or U2461 (N_2461,N_2227,N_2228);
or U2462 (N_2462,N_2173,N_2170);
nand U2463 (N_2463,N_2220,N_2232);
nand U2464 (N_2464,N_2006,N_2149);
xnor U2465 (N_2465,N_2144,N_2060);
nand U2466 (N_2466,N_2166,N_2206);
or U2467 (N_2467,N_2208,N_2228);
and U2468 (N_2468,N_2109,N_2234);
nor U2469 (N_2469,N_2094,N_2122);
or U2470 (N_2470,N_2127,N_2233);
or U2471 (N_2471,N_2185,N_2047);
and U2472 (N_2472,N_2161,N_2131);
nor U2473 (N_2473,N_2093,N_2236);
or U2474 (N_2474,N_2188,N_2005);
or U2475 (N_2475,N_2222,N_2147);
nand U2476 (N_2476,N_2072,N_2238);
nand U2477 (N_2477,N_2050,N_2137);
or U2478 (N_2478,N_2193,N_2218);
nor U2479 (N_2479,N_2114,N_2248);
xnor U2480 (N_2480,N_2009,N_2013);
or U2481 (N_2481,N_2050,N_2081);
or U2482 (N_2482,N_2221,N_2016);
and U2483 (N_2483,N_2197,N_2015);
or U2484 (N_2484,N_2190,N_2202);
nand U2485 (N_2485,N_2220,N_2105);
or U2486 (N_2486,N_2238,N_2097);
xor U2487 (N_2487,N_2091,N_2129);
or U2488 (N_2488,N_2069,N_2088);
nor U2489 (N_2489,N_2117,N_2035);
or U2490 (N_2490,N_2204,N_2015);
or U2491 (N_2491,N_2082,N_2139);
nor U2492 (N_2492,N_2197,N_2059);
xor U2493 (N_2493,N_2076,N_2109);
xnor U2494 (N_2494,N_2114,N_2198);
nand U2495 (N_2495,N_2044,N_2112);
or U2496 (N_2496,N_2069,N_2047);
nor U2497 (N_2497,N_2118,N_2071);
nand U2498 (N_2498,N_2172,N_2198);
nand U2499 (N_2499,N_2224,N_2244);
or U2500 (N_2500,N_2373,N_2259);
nor U2501 (N_2501,N_2411,N_2418);
and U2502 (N_2502,N_2399,N_2365);
or U2503 (N_2503,N_2293,N_2298);
nand U2504 (N_2504,N_2367,N_2296);
nand U2505 (N_2505,N_2398,N_2271);
nand U2506 (N_2506,N_2467,N_2308);
nand U2507 (N_2507,N_2316,N_2310);
nor U2508 (N_2508,N_2301,N_2360);
nand U2509 (N_2509,N_2427,N_2265);
and U2510 (N_2510,N_2452,N_2317);
nand U2511 (N_2511,N_2392,N_2419);
and U2512 (N_2512,N_2486,N_2483);
and U2513 (N_2513,N_2309,N_2498);
nor U2514 (N_2514,N_2257,N_2304);
nor U2515 (N_2515,N_2458,N_2376);
nor U2516 (N_2516,N_2444,N_2258);
xor U2517 (N_2517,N_2445,N_2457);
nand U2518 (N_2518,N_2253,N_2328);
nor U2519 (N_2519,N_2449,N_2471);
or U2520 (N_2520,N_2480,N_2269);
and U2521 (N_2521,N_2279,N_2340);
nor U2522 (N_2522,N_2432,N_2366);
nor U2523 (N_2523,N_2330,N_2435);
and U2524 (N_2524,N_2393,N_2312);
and U2525 (N_2525,N_2266,N_2256);
or U2526 (N_2526,N_2433,N_2277);
nor U2527 (N_2527,N_2369,N_2268);
nand U2528 (N_2528,N_2437,N_2494);
and U2529 (N_2529,N_2351,N_2254);
nand U2530 (N_2530,N_2335,N_2270);
xnor U2531 (N_2531,N_2421,N_2276);
and U2532 (N_2532,N_2462,N_2417);
nand U2533 (N_2533,N_2350,N_2288);
nand U2534 (N_2534,N_2464,N_2405);
or U2535 (N_2535,N_2368,N_2286);
nor U2536 (N_2536,N_2453,N_2447);
nor U2537 (N_2537,N_2319,N_2281);
nor U2538 (N_2538,N_2386,N_2451);
nor U2539 (N_2539,N_2388,N_2374);
or U2540 (N_2540,N_2285,N_2396);
nand U2541 (N_2541,N_2429,N_2355);
or U2542 (N_2542,N_2323,N_2381);
and U2543 (N_2543,N_2280,N_2278);
xor U2544 (N_2544,N_2315,N_2482);
nand U2545 (N_2545,N_2290,N_2299);
nand U2546 (N_2546,N_2476,N_2272);
and U2547 (N_2547,N_2463,N_2345);
and U2548 (N_2548,N_2456,N_2371);
xor U2549 (N_2549,N_2481,N_2260);
or U2550 (N_2550,N_2251,N_2460);
nand U2551 (N_2551,N_2344,N_2338);
nor U2552 (N_2552,N_2391,N_2375);
and U2553 (N_2553,N_2414,N_2384);
or U2554 (N_2554,N_2475,N_2262);
nand U2555 (N_2555,N_2305,N_2336);
nand U2556 (N_2556,N_2496,N_2264);
nand U2557 (N_2557,N_2383,N_2287);
xor U2558 (N_2558,N_2415,N_2466);
nand U2559 (N_2559,N_2422,N_2359);
nor U2560 (N_2560,N_2354,N_2321);
nor U2561 (N_2561,N_2306,N_2461);
nand U2562 (N_2562,N_2473,N_2395);
or U2563 (N_2563,N_2292,N_2313);
nor U2564 (N_2564,N_2250,N_2492);
and U2565 (N_2565,N_2283,N_2442);
nor U2566 (N_2566,N_2311,N_2327);
nand U2567 (N_2567,N_2361,N_2479);
and U2568 (N_2568,N_2425,N_2289);
and U2569 (N_2569,N_2346,N_2337);
or U2570 (N_2570,N_2294,N_2300);
nand U2571 (N_2571,N_2497,N_2389);
or U2572 (N_2572,N_2412,N_2404);
nor U2573 (N_2573,N_2379,N_2434);
xnor U2574 (N_2574,N_2485,N_2341);
nor U2575 (N_2575,N_2487,N_2261);
nor U2576 (N_2576,N_2339,N_2291);
nand U2577 (N_2577,N_2499,N_2401);
nor U2578 (N_2578,N_2358,N_2402);
and U2579 (N_2579,N_2380,N_2267);
or U2580 (N_2580,N_2420,N_2318);
nand U2581 (N_2581,N_2349,N_2430);
xnor U2582 (N_2582,N_2275,N_2416);
and U2583 (N_2583,N_2477,N_2438);
nor U2584 (N_2584,N_2363,N_2295);
nand U2585 (N_2585,N_2474,N_2390);
xor U2586 (N_2586,N_2413,N_2297);
nor U2587 (N_2587,N_2274,N_2441);
or U2588 (N_2588,N_2353,N_2439);
or U2589 (N_2589,N_2394,N_2364);
or U2590 (N_2590,N_2284,N_2331);
xnor U2591 (N_2591,N_2409,N_2408);
or U2592 (N_2592,N_2455,N_2490);
and U2593 (N_2593,N_2493,N_2465);
and U2594 (N_2594,N_2356,N_2469);
and U2595 (N_2595,N_2428,N_2282);
nor U2596 (N_2596,N_2377,N_2370);
and U2597 (N_2597,N_2378,N_2488);
xor U2598 (N_2598,N_2326,N_2329);
nor U2599 (N_2599,N_2252,N_2324);
nor U2600 (N_2600,N_2357,N_2382);
or U2601 (N_2601,N_2454,N_2440);
and U2602 (N_2602,N_2325,N_2424);
or U2603 (N_2603,N_2362,N_2431);
nor U2604 (N_2604,N_2255,N_2484);
and U2605 (N_2605,N_2478,N_2307);
nor U2606 (N_2606,N_2320,N_2342);
and U2607 (N_2607,N_2343,N_2436);
nor U2608 (N_2608,N_2410,N_2489);
nand U2609 (N_2609,N_2443,N_2372);
and U2610 (N_2610,N_2472,N_2273);
or U2611 (N_2611,N_2446,N_2385);
nor U2612 (N_2612,N_2426,N_2303);
nand U2613 (N_2613,N_2352,N_2423);
nand U2614 (N_2614,N_2263,N_2397);
nand U2615 (N_2615,N_2314,N_2403);
nor U2616 (N_2616,N_2387,N_2332);
xor U2617 (N_2617,N_2459,N_2333);
and U2618 (N_2618,N_2470,N_2491);
and U2619 (N_2619,N_2302,N_2406);
nand U2620 (N_2620,N_2347,N_2400);
or U2621 (N_2621,N_2348,N_2450);
nor U2622 (N_2622,N_2334,N_2407);
nand U2623 (N_2623,N_2468,N_2495);
or U2624 (N_2624,N_2448,N_2322);
nor U2625 (N_2625,N_2484,N_2445);
or U2626 (N_2626,N_2328,N_2315);
nor U2627 (N_2627,N_2496,N_2299);
or U2628 (N_2628,N_2377,N_2367);
nand U2629 (N_2629,N_2328,N_2329);
nand U2630 (N_2630,N_2316,N_2328);
or U2631 (N_2631,N_2355,N_2349);
nor U2632 (N_2632,N_2476,N_2482);
nand U2633 (N_2633,N_2444,N_2459);
or U2634 (N_2634,N_2428,N_2474);
or U2635 (N_2635,N_2479,N_2273);
or U2636 (N_2636,N_2298,N_2323);
nor U2637 (N_2637,N_2331,N_2434);
and U2638 (N_2638,N_2289,N_2450);
or U2639 (N_2639,N_2298,N_2455);
or U2640 (N_2640,N_2329,N_2499);
and U2641 (N_2641,N_2292,N_2317);
nor U2642 (N_2642,N_2441,N_2420);
nor U2643 (N_2643,N_2331,N_2499);
nor U2644 (N_2644,N_2282,N_2255);
nor U2645 (N_2645,N_2319,N_2474);
xor U2646 (N_2646,N_2319,N_2346);
or U2647 (N_2647,N_2284,N_2364);
xor U2648 (N_2648,N_2354,N_2475);
and U2649 (N_2649,N_2465,N_2270);
xor U2650 (N_2650,N_2265,N_2349);
nor U2651 (N_2651,N_2406,N_2427);
or U2652 (N_2652,N_2303,N_2468);
nor U2653 (N_2653,N_2429,N_2343);
or U2654 (N_2654,N_2491,N_2270);
or U2655 (N_2655,N_2435,N_2319);
or U2656 (N_2656,N_2456,N_2254);
nand U2657 (N_2657,N_2466,N_2316);
and U2658 (N_2658,N_2428,N_2327);
nor U2659 (N_2659,N_2378,N_2476);
and U2660 (N_2660,N_2324,N_2474);
or U2661 (N_2661,N_2488,N_2271);
and U2662 (N_2662,N_2351,N_2310);
xor U2663 (N_2663,N_2451,N_2430);
or U2664 (N_2664,N_2424,N_2441);
nor U2665 (N_2665,N_2311,N_2272);
nand U2666 (N_2666,N_2353,N_2488);
xor U2667 (N_2667,N_2398,N_2294);
or U2668 (N_2668,N_2278,N_2268);
nand U2669 (N_2669,N_2424,N_2300);
xnor U2670 (N_2670,N_2328,N_2317);
and U2671 (N_2671,N_2300,N_2456);
nand U2672 (N_2672,N_2376,N_2468);
or U2673 (N_2673,N_2450,N_2281);
or U2674 (N_2674,N_2252,N_2410);
nand U2675 (N_2675,N_2445,N_2479);
and U2676 (N_2676,N_2486,N_2434);
or U2677 (N_2677,N_2300,N_2358);
and U2678 (N_2678,N_2351,N_2409);
nor U2679 (N_2679,N_2394,N_2374);
and U2680 (N_2680,N_2442,N_2464);
and U2681 (N_2681,N_2407,N_2428);
or U2682 (N_2682,N_2287,N_2404);
nor U2683 (N_2683,N_2494,N_2360);
or U2684 (N_2684,N_2477,N_2453);
and U2685 (N_2685,N_2286,N_2251);
and U2686 (N_2686,N_2261,N_2343);
nor U2687 (N_2687,N_2405,N_2292);
nor U2688 (N_2688,N_2315,N_2255);
nand U2689 (N_2689,N_2459,N_2485);
nand U2690 (N_2690,N_2367,N_2485);
xnor U2691 (N_2691,N_2361,N_2498);
nor U2692 (N_2692,N_2267,N_2297);
or U2693 (N_2693,N_2427,N_2283);
xnor U2694 (N_2694,N_2391,N_2331);
or U2695 (N_2695,N_2326,N_2277);
xor U2696 (N_2696,N_2345,N_2270);
nand U2697 (N_2697,N_2338,N_2425);
or U2698 (N_2698,N_2467,N_2449);
nand U2699 (N_2699,N_2420,N_2429);
nand U2700 (N_2700,N_2255,N_2300);
and U2701 (N_2701,N_2293,N_2261);
nor U2702 (N_2702,N_2344,N_2288);
xnor U2703 (N_2703,N_2367,N_2341);
or U2704 (N_2704,N_2476,N_2399);
and U2705 (N_2705,N_2464,N_2373);
xor U2706 (N_2706,N_2252,N_2292);
and U2707 (N_2707,N_2361,N_2353);
and U2708 (N_2708,N_2459,N_2442);
nand U2709 (N_2709,N_2348,N_2392);
nor U2710 (N_2710,N_2285,N_2352);
and U2711 (N_2711,N_2411,N_2250);
nand U2712 (N_2712,N_2388,N_2359);
or U2713 (N_2713,N_2380,N_2422);
or U2714 (N_2714,N_2352,N_2498);
or U2715 (N_2715,N_2312,N_2380);
and U2716 (N_2716,N_2398,N_2362);
and U2717 (N_2717,N_2462,N_2446);
nor U2718 (N_2718,N_2362,N_2357);
nand U2719 (N_2719,N_2302,N_2389);
or U2720 (N_2720,N_2250,N_2285);
nand U2721 (N_2721,N_2483,N_2305);
nor U2722 (N_2722,N_2313,N_2311);
and U2723 (N_2723,N_2433,N_2311);
nand U2724 (N_2724,N_2450,N_2315);
nor U2725 (N_2725,N_2443,N_2393);
nand U2726 (N_2726,N_2446,N_2331);
nor U2727 (N_2727,N_2449,N_2325);
or U2728 (N_2728,N_2464,N_2316);
nand U2729 (N_2729,N_2254,N_2318);
or U2730 (N_2730,N_2352,N_2324);
and U2731 (N_2731,N_2447,N_2365);
and U2732 (N_2732,N_2378,N_2393);
nor U2733 (N_2733,N_2316,N_2418);
nor U2734 (N_2734,N_2474,N_2277);
and U2735 (N_2735,N_2447,N_2451);
nor U2736 (N_2736,N_2497,N_2443);
nand U2737 (N_2737,N_2480,N_2418);
and U2738 (N_2738,N_2340,N_2404);
nor U2739 (N_2739,N_2483,N_2312);
nand U2740 (N_2740,N_2468,N_2447);
or U2741 (N_2741,N_2456,N_2280);
and U2742 (N_2742,N_2449,N_2446);
or U2743 (N_2743,N_2486,N_2424);
and U2744 (N_2744,N_2330,N_2436);
nor U2745 (N_2745,N_2409,N_2253);
nand U2746 (N_2746,N_2418,N_2309);
or U2747 (N_2747,N_2251,N_2329);
nand U2748 (N_2748,N_2252,N_2282);
nand U2749 (N_2749,N_2389,N_2264);
nand U2750 (N_2750,N_2742,N_2583);
and U2751 (N_2751,N_2700,N_2521);
or U2752 (N_2752,N_2601,N_2565);
and U2753 (N_2753,N_2658,N_2524);
nand U2754 (N_2754,N_2647,N_2645);
and U2755 (N_2755,N_2589,N_2523);
xnor U2756 (N_2756,N_2689,N_2615);
and U2757 (N_2757,N_2690,N_2640);
nor U2758 (N_2758,N_2596,N_2633);
nor U2759 (N_2759,N_2665,N_2699);
nand U2760 (N_2760,N_2519,N_2528);
nand U2761 (N_2761,N_2575,N_2676);
or U2762 (N_2762,N_2569,N_2574);
nand U2763 (N_2763,N_2624,N_2610);
nand U2764 (N_2764,N_2622,N_2616);
nor U2765 (N_2765,N_2543,N_2687);
nor U2766 (N_2766,N_2570,N_2571);
nand U2767 (N_2767,N_2560,N_2515);
nor U2768 (N_2768,N_2664,N_2539);
nand U2769 (N_2769,N_2732,N_2558);
or U2770 (N_2770,N_2654,N_2582);
and U2771 (N_2771,N_2723,N_2627);
nand U2772 (N_2772,N_2604,N_2661);
and U2773 (N_2773,N_2675,N_2577);
or U2774 (N_2774,N_2729,N_2554);
nand U2775 (N_2775,N_2737,N_2681);
nor U2776 (N_2776,N_2709,N_2697);
or U2777 (N_2777,N_2608,N_2638);
nor U2778 (N_2778,N_2717,N_2694);
nand U2779 (N_2779,N_2708,N_2567);
nor U2780 (N_2780,N_2719,N_2642);
nand U2781 (N_2781,N_2650,N_2688);
nand U2782 (N_2782,N_2634,N_2651);
nand U2783 (N_2783,N_2612,N_2573);
or U2784 (N_2784,N_2630,N_2532);
nor U2785 (N_2785,N_2621,N_2551);
and U2786 (N_2786,N_2686,N_2663);
nand U2787 (N_2787,N_2679,N_2692);
nand U2788 (N_2788,N_2727,N_2656);
xnor U2789 (N_2789,N_2667,N_2741);
nor U2790 (N_2790,N_2525,N_2730);
and U2791 (N_2791,N_2516,N_2562);
nor U2792 (N_2792,N_2598,N_2626);
nor U2793 (N_2793,N_2710,N_2643);
nor U2794 (N_2794,N_2550,N_2628);
nand U2795 (N_2795,N_2619,N_2535);
and U2796 (N_2796,N_2597,N_2629);
or U2797 (N_2797,N_2715,N_2504);
nand U2798 (N_2798,N_2648,N_2544);
xor U2799 (N_2799,N_2744,N_2685);
nand U2800 (N_2800,N_2536,N_2733);
or U2801 (N_2801,N_2542,N_2579);
and U2802 (N_2802,N_2605,N_2631);
or U2803 (N_2803,N_2618,N_2509);
nor U2804 (N_2804,N_2713,N_2514);
xnor U2805 (N_2805,N_2563,N_2555);
and U2806 (N_2806,N_2572,N_2586);
or U2807 (N_2807,N_2607,N_2557);
and U2808 (N_2808,N_2540,N_2617);
and U2809 (N_2809,N_2644,N_2641);
or U2810 (N_2810,N_2613,N_2545);
nor U2811 (N_2811,N_2533,N_2623);
or U2812 (N_2812,N_2748,N_2501);
or U2813 (N_2813,N_2541,N_2507);
and U2814 (N_2814,N_2749,N_2672);
and U2815 (N_2815,N_2746,N_2502);
nor U2816 (N_2816,N_2506,N_2703);
nor U2817 (N_2817,N_2520,N_2736);
or U2818 (N_2818,N_2635,N_2691);
nor U2819 (N_2819,N_2718,N_2701);
and U2820 (N_2820,N_2580,N_2659);
xor U2821 (N_2821,N_2602,N_2743);
nor U2822 (N_2822,N_2548,N_2711);
nand U2823 (N_2823,N_2531,N_2720);
nand U2824 (N_2824,N_2518,N_2603);
or U2825 (N_2825,N_2508,N_2632);
nor U2826 (N_2826,N_2677,N_2553);
nand U2827 (N_2827,N_2725,N_2646);
and U2828 (N_2828,N_2660,N_2592);
or U2829 (N_2829,N_2588,N_2682);
or U2830 (N_2830,N_2581,N_2614);
nand U2831 (N_2831,N_2706,N_2747);
nor U2832 (N_2832,N_2561,N_2505);
nor U2833 (N_2833,N_2714,N_2513);
nor U2834 (N_2834,N_2500,N_2662);
or U2835 (N_2835,N_2716,N_2620);
or U2836 (N_2836,N_2704,N_2671);
or U2837 (N_2837,N_2693,N_2584);
nand U2838 (N_2838,N_2611,N_2740);
and U2839 (N_2839,N_2625,N_2670);
or U2840 (N_2840,N_2568,N_2546);
nand U2841 (N_2841,N_2657,N_2652);
nand U2842 (N_2842,N_2695,N_2739);
and U2843 (N_2843,N_2526,N_2530);
or U2844 (N_2844,N_2552,N_2722);
nand U2845 (N_2845,N_2517,N_2559);
xnor U2846 (N_2846,N_2698,N_2680);
and U2847 (N_2847,N_2609,N_2636);
and U2848 (N_2848,N_2594,N_2639);
nor U2849 (N_2849,N_2529,N_2578);
nor U2850 (N_2850,N_2538,N_2599);
nor U2851 (N_2851,N_2684,N_2734);
xor U2852 (N_2852,N_2591,N_2731);
and U2853 (N_2853,N_2745,N_2547);
xnor U2854 (N_2854,N_2585,N_2705);
nand U2855 (N_2855,N_2726,N_2537);
nor U2856 (N_2856,N_2721,N_2590);
nand U2857 (N_2857,N_2724,N_2600);
nand U2858 (N_2858,N_2668,N_2593);
or U2859 (N_2859,N_2649,N_2738);
nand U2860 (N_2860,N_2549,N_2707);
nand U2861 (N_2861,N_2673,N_2683);
nand U2862 (N_2862,N_2503,N_2712);
or U2863 (N_2863,N_2674,N_2564);
or U2864 (N_2864,N_2510,N_2696);
nand U2865 (N_2865,N_2702,N_2669);
nand U2866 (N_2866,N_2606,N_2595);
nor U2867 (N_2867,N_2522,N_2587);
nor U2868 (N_2868,N_2527,N_2735);
nor U2869 (N_2869,N_2511,N_2678);
nand U2870 (N_2870,N_2576,N_2655);
nand U2871 (N_2871,N_2566,N_2653);
nor U2872 (N_2872,N_2512,N_2556);
nor U2873 (N_2873,N_2666,N_2728);
xor U2874 (N_2874,N_2637,N_2534);
nand U2875 (N_2875,N_2581,N_2553);
or U2876 (N_2876,N_2525,N_2571);
or U2877 (N_2877,N_2618,N_2706);
nor U2878 (N_2878,N_2588,N_2552);
and U2879 (N_2879,N_2653,N_2655);
nand U2880 (N_2880,N_2536,N_2545);
xnor U2881 (N_2881,N_2672,N_2715);
xor U2882 (N_2882,N_2502,N_2546);
nor U2883 (N_2883,N_2516,N_2522);
nor U2884 (N_2884,N_2652,N_2609);
and U2885 (N_2885,N_2595,N_2737);
and U2886 (N_2886,N_2673,N_2712);
and U2887 (N_2887,N_2659,N_2692);
nand U2888 (N_2888,N_2679,N_2506);
xor U2889 (N_2889,N_2596,N_2628);
nor U2890 (N_2890,N_2607,N_2662);
nor U2891 (N_2891,N_2698,N_2690);
nor U2892 (N_2892,N_2622,N_2542);
nand U2893 (N_2893,N_2670,N_2544);
nand U2894 (N_2894,N_2721,N_2609);
xor U2895 (N_2895,N_2640,N_2599);
or U2896 (N_2896,N_2510,N_2570);
or U2897 (N_2897,N_2553,N_2624);
and U2898 (N_2898,N_2675,N_2698);
nor U2899 (N_2899,N_2688,N_2514);
and U2900 (N_2900,N_2633,N_2710);
nor U2901 (N_2901,N_2618,N_2571);
nor U2902 (N_2902,N_2503,N_2748);
or U2903 (N_2903,N_2542,N_2540);
nor U2904 (N_2904,N_2664,N_2698);
or U2905 (N_2905,N_2546,N_2586);
or U2906 (N_2906,N_2683,N_2677);
and U2907 (N_2907,N_2714,N_2623);
nand U2908 (N_2908,N_2746,N_2616);
nand U2909 (N_2909,N_2556,N_2644);
or U2910 (N_2910,N_2665,N_2615);
nand U2911 (N_2911,N_2558,N_2643);
nor U2912 (N_2912,N_2726,N_2521);
nor U2913 (N_2913,N_2695,N_2504);
or U2914 (N_2914,N_2658,N_2578);
nand U2915 (N_2915,N_2584,N_2573);
or U2916 (N_2916,N_2588,N_2607);
or U2917 (N_2917,N_2687,N_2660);
or U2918 (N_2918,N_2718,N_2731);
or U2919 (N_2919,N_2612,N_2593);
or U2920 (N_2920,N_2589,N_2678);
and U2921 (N_2921,N_2559,N_2653);
and U2922 (N_2922,N_2681,N_2676);
and U2923 (N_2923,N_2535,N_2569);
and U2924 (N_2924,N_2697,N_2526);
or U2925 (N_2925,N_2644,N_2618);
nand U2926 (N_2926,N_2621,N_2558);
or U2927 (N_2927,N_2645,N_2591);
xnor U2928 (N_2928,N_2602,N_2706);
or U2929 (N_2929,N_2587,N_2536);
or U2930 (N_2930,N_2556,N_2514);
and U2931 (N_2931,N_2681,N_2520);
or U2932 (N_2932,N_2642,N_2623);
nand U2933 (N_2933,N_2604,N_2737);
nand U2934 (N_2934,N_2528,N_2610);
and U2935 (N_2935,N_2610,N_2733);
and U2936 (N_2936,N_2683,N_2535);
or U2937 (N_2937,N_2560,N_2516);
or U2938 (N_2938,N_2583,N_2629);
nor U2939 (N_2939,N_2662,N_2569);
xnor U2940 (N_2940,N_2526,N_2723);
and U2941 (N_2941,N_2727,N_2539);
or U2942 (N_2942,N_2743,N_2567);
nand U2943 (N_2943,N_2692,N_2559);
or U2944 (N_2944,N_2635,N_2507);
nor U2945 (N_2945,N_2623,N_2573);
nand U2946 (N_2946,N_2662,N_2601);
nor U2947 (N_2947,N_2627,N_2606);
nand U2948 (N_2948,N_2652,N_2556);
nor U2949 (N_2949,N_2620,N_2698);
and U2950 (N_2950,N_2688,N_2518);
nand U2951 (N_2951,N_2662,N_2563);
or U2952 (N_2952,N_2706,N_2682);
and U2953 (N_2953,N_2700,N_2619);
and U2954 (N_2954,N_2718,N_2671);
nand U2955 (N_2955,N_2504,N_2745);
nand U2956 (N_2956,N_2694,N_2538);
and U2957 (N_2957,N_2746,N_2658);
nand U2958 (N_2958,N_2648,N_2511);
xor U2959 (N_2959,N_2590,N_2599);
and U2960 (N_2960,N_2687,N_2534);
or U2961 (N_2961,N_2721,N_2612);
or U2962 (N_2962,N_2727,N_2735);
and U2963 (N_2963,N_2744,N_2715);
and U2964 (N_2964,N_2610,N_2694);
and U2965 (N_2965,N_2608,N_2503);
or U2966 (N_2966,N_2577,N_2689);
and U2967 (N_2967,N_2613,N_2694);
nor U2968 (N_2968,N_2686,N_2695);
and U2969 (N_2969,N_2707,N_2685);
or U2970 (N_2970,N_2652,N_2688);
or U2971 (N_2971,N_2575,N_2554);
nand U2972 (N_2972,N_2535,N_2641);
or U2973 (N_2973,N_2693,N_2646);
nor U2974 (N_2974,N_2578,N_2590);
and U2975 (N_2975,N_2529,N_2547);
nand U2976 (N_2976,N_2554,N_2612);
nor U2977 (N_2977,N_2529,N_2648);
nor U2978 (N_2978,N_2700,N_2703);
and U2979 (N_2979,N_2679,N_2538);
or U2980 (N_2980,N_2642,N_2708);
nand U2981 (N_2981,N_2725,N_2583);
and U2982 (N_2982,N_2658,N_2661);
and U2983 (N_2983,N_2632,N_2603);
xnor U2984 (N_2984,N_2525,N_2642);
or U2985 (N_2985,N_2662,N_2595);
nand U2986 (N_2986,N_2738,N_2598);
or U2987 (N_2987,N_2587,N_2734);
and U2988 (N_2988,N_2700,N_2661);
or U2989 (N_2989,N_2741,N_2548);
xor U2990 (N_2990,N_2558,N_2733);
xnor U2991 (N_2991,N_2738,N_2533);
or U2992 (N_2992,N_2509,N_2655);
nand U2993 (N_2993,N_2618,N_2668);
nor U2994 (N_2994,N_2570,N_2549);
and U2995 (N_2995,N_2573,N_2613);
and U2996 (N_2996,N_2739,N_2713);
or U2997 (N_2997,N_2684,N_2575);
nand U2998 (N_2998,N_2680,N_2541);
nand U2999 (N_2999,N_2559,N_2508);
and U3000 (N_3000,N_2783,N_2842);
nor U3001 (N_3001,N_2894,N_2849);
nor U3002 (N_3002,N_2833,N_2765);
and U3003 (N_3003,N_2802,N_2846);
or U3004 (N_3004,N_2979,N_2975);
nor U3005 (N_3005,N_2836,N_2829);
and U3006 (N_3006,N_2798,N_2936);
and U3007 (N_3007,N_2834,N_2855);
and U3008 (N_3008,N_2985,N_2808);
or U3009 (N_3009,N_2954,N_2789);
or U3010 (N_3010,N_2790,N_2993);
xor U3011 (N_3011,N_2948,N_2759);
or U3012 (N_3012,N_2882,N_2897);
nor U3013 (N_3013,N_2949,N_2881);
nand U3014 (N_3014,N_2967,N_2776);
or U3015 (N_3015,N_2838,N_2786);
nand U3016 (N_3016,N_2755,N_2876);
or U3017 (N_3017,N_2792,N_2767);
or U3018 (N_3018,N_2856,N_2950);
nor U3019 (N_3019,N_2911,N_2885);
or U3020 (N_3020,N_2952,N_2983);
nor U3021 (N_3021,N_2916,N_2866);
or U3022 (N_3022,N_2957,N_2895);
and U3023 (N_3023,N_2915,N_2840);
nand U3024 (N_3024,N_2880,N_2988);
or U3025 (N_3025,N_2997,N_2977);
or U3026 (N_3026,N_2922,N_2784);
nand U3027 (N_3027,N_2809,N_2926);
or U3028 (N_3028,N_2814,N_2945);
or U3029 (N_3029,N_2843,N_2906);
nand U3030 (N_3030,N_2812,N_2837);
nand U3031 (N_3031,N_2995,N_2799);
or U3032 (N_3032,N_2861,N_2818);
nand U3033 (N_3033,N_2944,N_2811);
nor U3034 (N_3034,N_2779,N_2921);
nand U3035 (N_3035,N_2955,N_2807);
nor U3036 (N_3036,N_2850,N_2930);
nand U3037 (N_3037,N_2934,N_2782);
nor U3038 (N_3038,N_2973,N_2963);
or U3039 (N_3039,N_2788,N_2970);
or U3040 (N_3040,N_2974,N_2825);
xor U3041 (N_3041,N_2946,N_2870);
xnor U3042 (N_3042,N_2868,N_2819);
nor U3043 (N_3043,N_2907,N_2780);
nand U3044 (N_3044,N_2873,N_2901);
and U3045 (N_3045,N_2864,N_2917);
nand U3046 (N_3046,N_2800,N_2925);
and U3047 (N_3047,N_2938,N_2877);
or U3048 (N_3048,N_2933,N_2787);
nand U3049 (N_3049,N_2773,N_2998);
nor U3050 (N_3050,N_2832,N_2891);
nor U3051 (N_3051,N_2960,N_2781);
nand U3052 (N_3052,N_2888,N_2871);
xor U3053 (N_3053,N_2844,N_2953);
or U3054 (N_3054,N_2813,N_2968);
nand U3055 (N_3055,N_2791,N_2991);
and U3056 (N_3056,N_2996,N_2965);
or U3057 (N_3057,N_2956,N_2887);
xnor U3058 (N_3058,N_2869,N_2980);
or U3059 (N_3059,N_2939,N_2890);
and U3060 (N_3060,N_2865,N_2803);
xnor U3061 (N_3061,N_2824,N_2878);
nand U3062 (N_3062,N_2937,N_2879);
or U3063 (N_3063,N_2909,N_2893);
and U3064 (N_3064,N_2750,N_2794);
or U3065 (N_3065,N_2902,N_2986);
nor U3066 (N_3066,N_2820,N_2839);
or U3067 (N_3067,N_2999,N_2775);
nor U3068 (N_3068,N_2962,N_2827);
or U3069 (N_3069,N_2912,N_2896);
nor U3070 (N_3070,N_2947,N_2920);
xor U3071 (N_3071,N_2935,N_2994);
nor U3072 (N_3072,N_2772,N_2828);
nor U3073 (N_3073,N_2778,N_2845);
xnor U3074 (N_3074,N_2969,N_2764);
and U3075 (N_3075,N_2966,N_2931);
nor U3076 (N_3076,N_2910,N_2908);
xnor U3077 (N_3077,N_2984,N_2990);
and U3078 (N_3078,N_2805,N_2810);
nand U3079 (N_3079,N_2905,N_2981);
nor U3080 (N_3080,N_2927,N_2872);
or U3081 (N_3081,N_2900,N_2768);
or U3082 (N_3082,N_2929,N_2958);
and U3083 (N_3083,N_2961,N_2815);
and U3084 (N_3084,N_2848,N_2889);
or U3085 (N_3085,N_2806,N_2989);
nor U3086 (N_3086,N_2752,N_2756);
or U3087 (N_3087,N_2831,N_2854);
nand U3088 (N_3088,N_2817,N_2851);
nand U3089 (N_3089,N_2801,N_2987);
xor U3090 (N_3090,N_2821,N_2853);
and U3091 (N_3091,N_2785,N_2771);
nor U3092 (N_3092,N_2903,N_2835);
nor U3093 (N_3093,N_2830,N_2976);
or U3094 (N_3094,N_2884,N_2761);
and U3095 (N_3095,N_2860,N_2932);
nor U3096 (N_3096,N_2859,N_2923);
nor U3097 (N_3097,N_2892,N_2918);
nand U3098 (N_3098,N_2751,N_2857);
and U3099 (N_3099,N_2914,N_2795);
or U3100 (N_3100,N_2978,N_2886);
and U3101 (N_3101,N_2992,N_2758);
xor U3102 (N_3102,N_2847,N_2919);
xor U3103 (N_3103,N_2862,N_2982);
nand U3104 (N_3104,N_2972,N_2971);
and U3105 (N_3105,N_2763,N_2793);
nand U3106 (N_3106,N_2777,N_2823);
and U3107 (N_3107,N_2753,N_2762);
nand U3108 (N_3108,N_2904,N_2757);
and U3109 (N_3109,N_2760,N_2852);
nor U3110 (N_3110,N_2964,N_2875);
nand U3111 (N_3111,N_2913,N_2774);
nand U3112 (N_3112,N_2874,N_2841);
nor U3113 (N_3113,N_2766,N_2943);
or U3114 (N_3114,N_2928,N_2942);
xor U3115 (N_3115,N_2769,N_2883);
nor U3116 (N_3116,N_2804,N_2959);
nor U3117 (N_3117,N_2941,N_2867);
nor U3118 (N_3118,N_2796,N_2822);
xnor U3119 (N_3119,N_2826,N_2816);
nor U3120 (N_3120,N_2863,N_2754);
nor U3121 (N_3121,N_2924,N_2898);
and U3122 (N_3122,N_2951,N_2940);
and U3123 (N_3123,N_2858,N_2899);
nand U3124 (N_3124,N_2770,N_2797);
nor U3125 (N_3125,N_2803,N_2947);
nor U3126 (N_3126,N_2832,N_2787);
nand U3127 (N_3127,N_2903,N_2857);
or U3128 (N_3128,N_2961,N_2887);
nor U3129 (N_3129,N_2917,N_2775);
nor U3130 (N_3130,N_2777,N_2974);
xnor U3131 (N_3131,N_2935,N_2913);
nand U3132 (N_3132,N_2793,N_2772);
or U3133 (N_3133,N_2943,N_2942);
or U3134 (N_3134,N_2943,N_2775);
nor U3135 (N_3135,N_2888,N_2969);
and U3136 (N_3136,N_2770,N_2942);
or U3137 (N_3137,N_2937,N_2975);
and U3138 (N_3138,N_2983,N_2858);
nor U3139 (N_3139,N_2792,N_2833);
and U3140 (N_3140,N_2998,N_2789);
nand U3141 (N_3141,N_2790,N_2894);
and U3142 (N_3142,N_2828,N_2867);
and U3143 (N_3143,N_2811,N_2927);
and U3144 (N_3144,N_2810,N_2945);
and U3145 (N_3145,N_2819,N_2950);
and U3146 (N_3146,N_2961,N_2840);
or U3147 (N_3147,N_2755,N_2904);
nand U3148 (N_3148,N_2979,N_2980);
nor U3149 (N_3149,N_2782,N_2916);
nor U3150 (N_3150,N_2904,N_2964);
and U3151 (N_3151,N_2990,N_2789);
or U3152 (N_3152,N_2964,N_2946);
nor U3153 (N_3153,N_2816,N_2778);
nand U3154 (N_3154,N_2896,N_2998);
and U3155 (N_3155,N_2848,N_2837);
nor U3156 (N_3156,N_2793,N_2870);
nor U3157 (N_3157,N_2933,N_2986);
nor U3158 (N_3158,N_2867,N_2907);
xor U3159 (N_3159,N_2964,N_2818);
nor U3160 (N_3160,N_2862,N_2858);
nor U3161 (N_3161,N_2820,N_2875);
or U3162 (N_3162,N_2963,N_2910);
or U3163 (N_3163,N_2951,N_2837);
nor U3164 (N_3164,N_2965,N_2974);
and U3165 (N_3165,N_2942,N_2759);
or U3166 (N_3166,N_2844,N_2859);
or U3167 (N_3167,N_2945,N_2889);
and U3168 (N_3168,N_2989,N_2753);
nor U3169 (N_3169,N_2754,N_2973);
nand U3170 (N_3170,N_2802,N_2833);
xnor U3171 (N_3171,N_2782,N_2829);
and U3172 (N_3172,N_2925,N_2798);
nor U3173 (N_3173,N_2946,N_2976);
and U3174 (N_3174,N_2894,N_2757);
nor U3175 (N_3175,N_2784,N_2761);
and U3176 (N_3176,N_2825,N_2939);
nor U3177 (N_3177,N_2833,N_2995);
nor U3178 (N_3178,N_2765,N_2752);
nor U3179 (N_3179,N_2911,N_2847);
or U3180 (N_3180,N_2856,N_2865);
nor U3181 (N_3181,N_2882,N_2988);
xor U3182 (N_3182,N_2845,N_2905);
and U3183 (N_3183,N_2817,N_2825);
and U3184 (N_3184,N_2767,N_2768);
nand U3185 (N_3185,N_2990,N_2774);
and U3186 (N_3186,N_2781,N_2944);
or U3187 (N_3187,N_2917,N_2844);
nor U3188 (N_3188,N_2968,N_2970);
nand U3189 (N_3189,N_2989,N_2891);
xnor U3190 (N_3190,N_2989,N_2954);
and U3191 (N_3191,N_2817,N_2756);
and U3192 (N_3192,N_2863,N_2989);
and U3193 (N_3193,N_2998,N_2870);
or U3194 (N_3194,N_2871,N_2890);
or U3195 (N_3195,N_2757,N_2998);
and U3196 (N_3196,N_2954,N_2986);
nand U3197 (N_3197,N_2751,N_2900);
nor U3198 (N_3198,N_2752,N_2960);
nor U3199 (N_3199,N_2773,N_2866);
or U3200 (N_3200,N_2865,N_2890);
and U3201 (N_3201,N_2911,N_2792);
nor U3202 (N_3202,N_2841,N_2906);
and U3203 (N_3203,N_2861,N_2759);
xor U3204 (N_3204,N_2925,N_2955);
or U3205 (N_3205,N_2890,N_2928);
nor U3206 (N_3206,N_2971,N_2786);
nor U3207 (N_3207,N_2864,N_2815);
nand U3208 (N_3208,N_2821,N_2825);
and U3209 (N_3209,N_2901,N_2927);
or U3210 (N_3210,N_2929,N_2823);
or U3211 (N_3211,N_2930,N_2922);
and U3212 (N_3212,N_2841,N_2800);
or U3213 (N_3213,N_2919,N_2889);
nor U3214 (N_3214,N_2961,N_2830);
nor U3215 (N_3215,N_2877,N_2900);
or U3216 (N_3216,N_2891,N_2864);
xnor U3217 (N_3217,N_2936,N_2963);
or U3218 (N_3218,N_2901,N_2787);
and U3219 (N_3219,N_2777,N_2760);
and U3220 (N_3220,N_2785,N_2826);
nor U3221 (N_3221,N_2779,N_2911);
and U3222 (N_3222,N_2796,N_2753);
or U3223 (N_3223,N_2885,N_2868);
xnor U3224 (N_3224,N_2795,N_2765);
nand U3225 (N_3225,N_2970,N_2803);
nand U3226 (N_3226,N_2764,N_2985);
and U3227 (N_3227,N_2780,N_2985);
and U3228 (N_3228,N_2766,N_2966);
or U3229 (N_3229,N_2964,N_2792);
or U3230 (N_3230,N_2751,N_2811);
nand U3231 (N_3231,N_2880,N_2982);
xnor U3232 (N_3232,N_2967,N_2924);
xnor U3233 (N_3233,N_2858,N_2845);
nand U3234 (N_3234,N_2930,N_2782);
and U3235 (N_3235,N_2766,N_2774);
nand U3236 (N_3236,N_2776,N_2893);
or U3237 (N_3237,N_2897,N_2800);
nand U3238 (N_3238,N_2968,N_2931);
nand U3239 (N_3239,N_2998,N_2990);
and U3240 (N_3240,N_2987,N_2900);
nor U3241 (N_3241,N_2941,N_2939);
nor U3242 (N_3242,N_2879,N_2915);
nand U3243 (N_3243,N_2975,N_2974);
nand U3244 (N_3244,N_2943,N_2829);
or U3245 (N_3245,N_2869,N_2793);
nand U3246 (N_3246,N_2769,N_2922);
nor U3247 (N_3247,N_2793,N_2788);
xnor U3248 (N_3248,N_2930,N_2815);
and U3249 (N_3249,N_2876,N_2937);
or U3250 (N_3250,N_3101,N_3018);
or U3251 (N_3251,N_3016,N_3045);
or U3252 (N_3252,N_3079,N_3173);
nand U3253 (N_3253,N_3144,N_3139);
or U3254 (N_3254,N_3196,N_3064);
nor U3255 (N_3255,N_3058,N_3230);
nand U3256 (N_3256,N_3061,N_3067);
xnor U3257 (N_3257,N_3108,N_3096);
or U3258 (N_3258,N_3050,N_3154);
and U3259 (N_3259,N_3161,N_3080);
nor U3260 (N_3260,N_3219,N_3147);
nor U3261 (N_3261,N_3125,N_3231);
xor U3262 (N_3262,N_3035,N_3094);
nor U3263 (N_3263,N_3047,N_3142);
and U3264 (N_3264,N_3100,N_3241);
and U3265 (N_3265,N_3111,N_3178);
nor U3266 (N_3266,N_3185,N_3207);
and U3267 (N_3267,N_3148,N_3118);
nand U3268 (N_3268,N_3209,N_3056);
or U3269 (N_3269,N_3120,N_3038);
xnor U3270 (N_3270,N_3183,N_3040);
and U3271 (N_3271,N_3223,N_3075);
nor U3272 (N_3272,N_3098,N_3189);
nand U3273 (N_3273,N_3221,N_3232);
nor U3274 (N_3274,N_3205,N_3225);
and U3275 (N_3275,N_3062,N_3169);
and U3276 (N_3276,N_3210,N_3179);
nor U3277 (N_3277,N_3030,N_3171);
and U3278 (N_3278,N_3106,N_3182);
nand U3279 (N_3279,N_3107,N_3020);
nand U3280 (N_3280,N_3136,N_3117);
or U3281 (N_3281,N_3034,N_3188);
or U3282 (N_3282,N_3156,N_3002);
nor U3283 (N_3283,N_3175,N_3124);
xnor U3284 (N_3284,N_3194,N_3163);
and U3285 (N_3285,N_3087,N_3127);
or U3286 (N_3286,N_3095,N_3217);
or U3287 (N_3287,N_3190,N_3104);
nand U3288 (N_3288,N_3160,N_3081);
and U3289 (N_3289,N_3206,N_3119);
or U3290 (N_3290,N_3017,N_3074);
xnor U3291 (N_3291,N_3009,N_3069);
or U3292 (N_3292,N_3245,N_3170);
nor U3293 (N_3293,N_3110,N_3021);
nand U3294 (N_3294,N_3236,N_3138);
nor U3295 (N_3295,N_3141,N_3208);
nor U3296 (N_3296,N_3083,N_3114);
nand U3297 (N_3297,N_3229,N_3036);
nor U3298 (N_3298,N_3072,N_3088);
and U3299 (N_3299,N_3240,N_3049);
and U3300 (N_3300,N_3168,N_3105);
nor U3301 (N_3301,N_3073,N_3126);
xnor U3302 (N_3302,N_3066,N_3243);
or U3303 (N_3303,N_3023,N_3186);
xnor U3304 (N_3304,N_3068,N_3115);
nand U3305 (N_3305,N_3005,N_3197);
or U3306 (N_3306,N_3007,N_3137);
and U3307 (N_3307,N_3248,N_3015);
or U3308 (N_3308,N_3203,N_3130);
and U3309 (N_3309,N_3011,N_3247);
nand U3310 (N_3310,N_3006,N_3218);
nand U3311 (N_3311,N_3180,N_3084);
nand U3312 (N_3312,N_3140,N_3019);
nand U3313 (N_3313,N_3102,N_3165);
and U3314 (N_3314,N_3151,N_3202);
nand U3315 (N_3315,N_3085,N_3042);
and U3316 (N_3316,N_3060,N_3063);
or U3317 (N_3317,N_3046,N_3199);
nand U3318 (N_3318,N_3043,N_3145);
nor U3319 (N_3319,N_3132,N_3033);
and U3320 (N_3320,N_3028,N_3013);
nand U3321 (N_3321,N_3158,N_3135);
or U3322 (N_3322,N_3201,N_3224);
xor U3323 (N_3323,N_3044,N_3014);
or U3324 (N_3324,N_3071,N_3131);
or U3325 (N_3325,N_3109,N_3192);
nor U3326 (N_3326,N_3001,N_3200);
xnor U3327 (N_3327,N_3057,N_3143);
and U3328 (N_3328,N_3012,N_3093);
or U3329 (N_3329,N_3181,N_3249);
or U3330 (N_3330,N_3238,N_3198);
nor U3331 (N_3331,N_3193,N_3025);
or U3332 (N_3332,N_3032,N_3082);
nand U3333 (N_3333,N_3176,N_3022);
or U3334 (N_3334,N_3157,N_3055);
or U3335 (N_3335,N_3152,N_3213);
or U3336 (N_3336,N_3133,N_3214);
or U3337 (N_3337,N_3123,N_3031);
and U3338 (N_3338,N_3053,N_3167);
or U3339 (N_3339,N_3146,N_3091);
and U3340 (N_3340,N_3010,N_3177);
or U3341 (N_3341,N_3195,N_3166);
and U3342 (N_3342,N_3065,N_3164);
nand U3343 (N_3343,N_3078,N_3116);
or U3344 (N_3344,N_3204,N_3041);
and U3345 (N_3345,N_3051,N_3172);
nand U3346 (N_3346,N_3003,N_3244);
nor U3347 (N_3347,N_3070,N_3246);
nor U3348 (N_3348,N_3159,N_3187);
and U3349 (N_3349,N_3024,N_3155);
and U3350 (N_3350,N_3099,N_3048);
and U3351 (N_3351,N_3162,N_3026);
nor U3352 (N_3352,N_3128,N_3228);
xnor U3353 (N_3353,N_3122,N_3134);
nor U3354 (N_3354,N_3077,N_3097);
nand U3355 (N_3355,N_3027,N_3234);
and U3356 (N_3356,N_3092,N_3000);
and U3357 (N_3357,N_3184,N_3076);
and U3358 (N_3358,N_3215,N_3129);
and U3359 (N_3359,N_3090,N_3008);
and U3360 (N_3360,N_3212,N_3191);
nand U3361 (N_3361,N_3059,N_3242);
nor U3362 (N_3362,N_3239,N_3211);
and U3363 (N_3363,N_3226,N_3103);
nor U3364 (N_3364,N_3037,N_3039);
nor U3365 (N_3365,N_3004,N_3235);
xor U3366 (N_3366,N_3216,N_3113);
and U3367 (N_3367,N_3029,N_3227);
nand U3368 (N_3368,N_3086,N_3174);
and U3369 (N_3369,N_3233,N_3089);
nand U3370 (N_3370,N_3222,N_3220);
and U3371 (N_3371,N_3052,N_3149);
or U3372 (N_3372,N_3237,N_3153);
xnor U3373 (N_3373,N_3112,N_3121);
nand U3374 (N_3374,N_3054,N_3150);
nand U3375 (N_3375,N_3249,N_3140);
xor U3376 (N_3376,N_3089,N_3235);
xor U3377 (N_3377,N_3240,N_3144);
and U3378 (N_3378,N_3051,N_3042);
or U3379 (N_3379,N_3196,N_3141);
or U3380 (N_3380,N_3191,N_3137);
nand U3381 (N_3381,N_3108,N_3141);
nor U3382 (N_3382,N_3053,N_3076);
nor U3383 (N_3383,N_3211,N_3126);
or U3384 (N_3384,N_3227,N_3180);
nand U3385 (N_3385,N_3185,N_3046);
or U3386 (N_3386,N_3210,N_3008);
and U3387 (N_3387,N_3102,N_3028);
nand U3388 (N_3388,N_3076,N_3095);
nand U3389 (N_3389,N_3226,N_3133);
and U3390 (N_3390,N_3139,N_3231);
nand U3391 (N_3391,N_3199,N_3110);
and U3392 (N_3392,N_3155,N_3211);
xnor U3393 (N_3393,N_3248,N_3236);
and U3394 (N_3394,N_3090,N_3246);
and U3395 (N_3395,N_3005,N_3069);
or U3396 (N_3396,N_3110,N_3023);
and U3397 (N_3397,N_3139,N_3200);
or U3398 (N_3398,N_3121,N_3017);
or U3399 (N_3399,N_3193,N_3124);
nor U3400 (N_3400,N_3217,N_3086);
and U3401 (N_3401,N_3078,N_3142);
and U3402 (N_3402,N_3194,N_3010);
and U3403 (N_3403,N_3105,N_3172);
xnor U3404 (N_3404,N_3109,N_3063);
nor U3405 (N_3405,N_3004,N_3019);
or U3406 (N_3406,N_3072,N_3194);
or U3407 (N_3407,N_3249,N_3014);
or U3408 (N_3408,N_3047,N_3005);
nor U3409 (N_3409,N_3015,N_3061);
and U3410 (N_3410,N_3027,N_3154);
and U3411 (N_3411,N_3195,N_3005);
nand U3412 (N_3412,N_3040,N_3101);
xnor U3413 (N_3413,N_3189,N_3033);
and U3414 (N_3414,N_3109,N_3102);
nand U3415 (N_3415,N_3136,N_3218);
nand U3416 (N_3416,N_3047,N_3008);
nor U3417 (N_3417,N_3056,N_3005);
nand U3418 (N_3418,N_3049,N_3129);
nand U3419 (N_3419,N_3020,N_3132);
and U3420 (N_3420,N_3030,N_3223);
or U3421 (N_3421,N_3230,N_3226);
nor U3422 (N_3422,N_3032,N_3165);
and U3423 (N_3423,N_3091,N_3024);
xnor U3424 (N_3424,N_3146,N_3206);
nor U3425 (N_3425,N_3207,N_3145);
xnor U3426 (N_3426,N_3126,N_3179);
and U3427 (N_3427,N_3045,N_3138);
nand U3428 (N_3428,N_3169,N_3008);
xnor U3429 (N_3429,N_3194,N_3061);
nor U3430 (N_3430,N_3046,N_3061);
nor U3431 (N_3431,N_3058,N_3052);
xnor U3432 (N_3432,N_3232,N_3084);
nor U3433 (N_3433,N_3197,N_3059);
nor U3434 (N_3434,N_3055,N_3249);
nand U3435 (N_3435,N_3083,N_3187);
and U3436 (N_3436,N_3131,N_3188);
or U3437 (N_3437,N_3213,N_3208);
or U3438 (N_3438,N_3123,N_3102);
nand U3439 (N_3439,N_3014,N_3209);
or U3440 (N_3440,N_3112,N_3079);
nand U3441 (N_3441,N_3125,N_3037);
xor U3442 (N_3442,N_3185,N_3173);
or U3443 (N_3443,N_3165,N_3066);
xnor U3444 (N_3444,N_3082,N_3200);
and U3445 (N_3445,N_3155,N_3097);
nand U3446 (N_3446,N_3199,N_3045);
nand U3447 (N_3447,N_3108,N_3241);
nand U3448 (N_3448,N_3075,N_3211);
and U3449 (N_3449,N_3039,N_3004);
nand U3450 (N_3450,N_3040,N_3082);
nor U3451 (N_3451,N_3119,N_3162);
or U3452 (N_3452,N_3011,N_3105);
or U3453 (N_3453,N_3078,N_3162);
nor U3454 (N_3454,N_3049,N_3152);
or U3455 (N_3455,N_3221,N_3090);
xor U3456 (N_3456,N_3247,N_3027);
and U3457 (N_3457,N_3075,N_3245);
or U3458 (N_3458,N_3125,N_3009);
or U3459 (N_3459,N_3131,N_3078);
nand U3460 (N_3460,N_3236,N_3249);
nand U3461 (N_3461,N_3232,N_3226);
and U3462 (N_3462,N_3058,N_3154);
or U3463 (N_3463,N_3016,N_3069);
nand U3464 (N_3464,N_3058,N_3006);
xnor U3465 (N_3465,N_3199,N_3188);
and U3466 (N_3466,N_3048,N_3111);
and U3467 (N_3467,N_3246,N_3117);
nand U3468 (N_3468,N_3009,N_3060);
nor U3469 (N_3469,N_3222,N_3070);
nor U3470 (N_3470,N_3247,N_3141);
nor U3471 (N_3471,N_3063,N_3091);
and U3472 (N_3472,N_3025,N_3035);
or U3473 (N_3473,N_3088,N_3041);
nor U3474 (N_3474,N_3063,N_3094);
or U3475 (N_3475,N_3201,N_3056);
nor U3476 (N_3476,N_3126,N_3223);
or U3477 (N_3477,N_3206,N_3238);
and U3478 (N_3478,N_3185,N_3023);
or U3479 (N_3479,N_3178,N_3004);
nand U3480 (N_3480,N_3134,N_3125);
nand U3481 (N_3481,N_3191,N_3173);
and U3482 (N_3482,N_3016,N_3033);
nand U3483 (N_3483,N_3236,N_3103);
and U3484 (N_3484,N_3120,N_3227);
and U3485 (N_3485,N_3222,N_3029);
nor U3486 (N_3486,N_3032,N_3109);
and U3487 (N_3487,N_3192,N_3096);
nand U3488 (N_3488,N_3098,N_3106);
or U3489 (N_3489,N_3040,N_3036);
or U3490 (N_3490,N_3072,N_3245);
xor U3491 (N_3491,N_3089,N_3192);
or U3492 (N_3492,N_3088,N_3091);
and U3493 (N_3493,N_3194,N_3210);
and U3494 (N_3494,N_3057,N_3249);
or U3495 (N_3495,N_3083,N_3084);
nor U3496 (N_3496,N_3085,N_3000);
nor U3497 (N_3497,N_3135,N_3035);
nor U3498 (N_3498,N_3126,N_3040);
nand U3499 (N_3499,N_3208,N_3097);
and U3500 (N_3500,N_3486,N_3355);
or U3501 (N_3501,N_3328,N_3427);
and U3502 (N_3502,N_3269,N_3430);
or U3503 (N_3503,N_3481,N_3408);
nor U3504 (N_3504,N_3395,N_3267);
and U3505 (N_3505,N_3346,N_3413);
nand U3506 (N_3506,N_3389,N_3354);
nand U3507 (N_3507,N_3420,N_3336);
or U3508 (N_3508,N_3313,N_3296);
nor U3509 (N_3509,N_3251,N_3468);
and U3510 (N_3510,N_3320,N_3387);
or U3511 (N_3511,N_3291,N_3488);
and U3512 (N_3512,N_3283,N_3286);
or U3513 (N_3513,N_3396,N_3435);
nand U3514 (N_3514,N_3268,N_3423);
or U3515 (N_3515,N_3479,N_3455);
xnor U3516 (N_3516,N_3311,N_3397);
or U3517 (N_3517,N_3298,N_3460);
nor U3518 (N_3518,N_3330,N_3329);
nand U3519 (N_3519,N_3318,N_3492);
nor U3520 (N_3520,N_3357,N_3288);
and U3521 (N_3521,N_3327,N_3418);
or U3522 (N_3522,N_3446,N_3258);
and U3523 (N_3523,N_3473,N_3294);
xnor U3524 (N_3524,N_3301,N_3458);
nand U3525 (N_3525,N_3487,N_3347);
and U3526 (N_3526,N_3266,N_3381);
nor U3527 (N_3527,N_3363,N_3367);
and U3528 (N_3528,N_3308,N_3404);
nand U3529 (N_3529,N_3449,N_3332);
and U3530 (N_3530,N_3457,N_3314);
nor U3531 (N_3531,N_3276,N_3338);
nand U3532 (N_3532,N_3401,N_3317);
xor U3533 (N_3533,N_3371,N_3364);
nor U3534 (N_3534,N_3254,N_3358);
nor U3535 (N_3535,N_3461,N_3496);
nand U3536 (N_3536,N_3337,N_3440);
nand U3537 (N_3537,N_3275,N_3482);
or U3538 (N_3538,N_3256,N_3421);
nor U3539 (N_3539,N_3369,N_3334);
nor U3540 (N_3540,N_3265,N_3277);
nor U3541 (N_3541,N_3469,N_3433);
or U3542 (N_3542,N_3478,N_3491);
or U3543 (N_3543,N_3304,N_3339);
nand U3544 (N_3544,N_3352,N_3426);
or U3545 (N_3545,N_3470,N_3459);
nand U3546 (N_3546,N_3490,N_3303);
nand U3547 (N_3547,N_3350,N_3484);
nand U3548 (N_3548,N_3333,N_3359);
or U3549 (N_3549,N_3410,N_3305);
or U3550 (N_3550,N_3432,N_3343);
nand U3551 (N_3551,N_3411,N_3263);
and U3552 (N_3552,N_3429,N_3417);
and U3553 (N_3553,N_3422,N_3377);
nand U3554 (N_3554,N_3253,N_3451);
nor U3555 (N_3555,N_3365,N_3398);
or U3556 (N_3556,N_3462,N_3340);
nand U3557 (N_3557,N_3374,N_3274);
nor U3558 (N_3558,N_3375,N_3450);
and U3559 (N_3559,N_3316,N_3376);
nor U3560 (N_3560,N_3373,N_3448);
nand U3561 (N_3561,N_3441,N_3424);
xnor U3562 (N_3562,N_3349,N_3498);
or U3563 (N_3563,N_3271,N_3425);
and U3564 (N_3564,N_3467,N_3335);
nor U3565 (N_3565,N_3285,N_3264);
or U3566 (N_3566,N_3259,N_3439);
and U3567 (N_3567,N_3443,N_3326);
or U3568 (N_3568,N_3345,N_3250);
and U3569 (N_3569,N_3454,N_3366);
nand U3570 (N_3570,N_3279,N_3261);
nand U3571 (N_3571,N_3436,N_3306);
nor U3572 (N_3572,N_3483,N_3257);
and U3573 (N_3573,N_3262,N_3452);
and U3574 (N_3574,N_3463,N_3287);
nor U3575 (N_3575,N_3322,N_3400);
nand U3576 (N_3576,N_3447,N_3284);
or U3577 (N_3577,N_3407,N_3475);
xor U3578 (N_3578,N_3499,N_3270);
xnor U3579 (N_3579,N_3370,N_3412);
nand U3580 (N_3580,N_3278,N_3299);
nor U3581 (N_3581,N_3403,N_3466);
nand U3582 (N_3582,N_3379,N_3471);
and U3583 (N_3583,N_3321,N_3344);
and U3584 (N_3584,N_3319,N_3282);
or U3585 (N_3585,N_3356,N_3391);
and U3586 (N_3586,N_3260,N_3480);
and U3587 (N_3587,N_3297,N_3292);
or U3588 (N_3588,N_3378,N_3315);
or U3589 (N_3589,N_3353,N_3409);
nand U3590 (N_3590,N_3309,N_3302);
and U3591 (N_3591,N_3384,N_3348);
and U3592 (N_3592,N_3392,N_3431);
nand U3593 (N_3593,N_3293,N_3489);
or U3594 (N_3594,N_3399,N_3341);
nor U3595 (N_3595,N_3405,N_3402);
or U3596 (N_3596,N_3485,N_3494);
xnor U3597 (N_3597,N_3289,N_3428);
and U3598 (N_3598,N_3324,N_3255);
or U3599 (N_3599,N_3497,N_3493);
nor U3600 (N_3600,N_3437,N_3453);
nor U3601 (N_3601,N_3273,N_3290);
nor U3602 (N_3602,N_3414,N_3464);
xor U3603 (N_3603,N_3307,N_3361);
and U3604 (N_3604,N_3360,N_3456);
nand U3605 (N_3605,N_3442,N_3444);
or U3606 (N_3606,N_3362,N_3382);
and U3607 (N_3607,N_3252,N_3394);
and U3608 (N_3608,N_3415,N_3393);
nor U3609 (N_3609,N_3477,N_3434);
or U3610 (N_3610,N_3295,N_3383);
and U3611 (N_3611,N_3472,N_3419);
and U3612 (N_3612,N_3476,N_3465);
and U3613 (N_3613,N_3281,N_3323);
nand U3614 (N_3614,N_3300,N_3312);
and U3615 (N_3615,N_3390,N_3325);
and U3616 (N_3616,N_3386,N_3445);
nand U3617 (N_3617,N_3474,N_3406);
nor U3618 (N_3618,N_3280,N_3331);
and U3619 (N_3619,N_3351,N_3272);
nand U3620 (N_3620,N_3385,N_3495);
nor U3621 (N_3621,N_3342,N_3380);
nand U3622 (N_3622,N_3388,N_3372);
or U3623 (N_3623,N_3310,N_3438);
nor U3624 (N_3624,N_3368,N_3416);
nand U3625 (N_3625,N_3300,N_3276);
nand U3626 (N_3626,N_3365,N_3264);
and U3627 (N_3627,N_3350,N_3492);
and U3628 (N_3628,N_3383,N_3326);
nand U3629 (N_3629,N_3488,N_3499);
nor U3630 (N_3630,N_3435,N_3290);
or U3631 (N_3631,N_3253,N_3320);
xnor U3632 (N_3632,N_3288,N_3489);
or U3633 (N_3633,N_3441,N_3339);
xor U3634 (N_3634,N_3292,N_3364);
xnor U3635 (N_3635,N_3282,N_3305);
or U3636 (N_3636,N_3395,N_3320);
or U3637 (N_3637,N_3316,N_3262);
nor U3638 (N_3638,N_3441,N_3288);
nand U3639 (N_3639,N_3423,N_3251);
nor U3640 (N_3640,N_3315,N_3421);
xnor U3641 (N_3641,N_3269,N_3371);
nand U3642 (N_3642,N_3277,N_3330);
xor U3643 (N_3643,N_3296,N_3261);
nand U3644 (N_3644,N_3323,N_3495);
and U3645 (N_3645,N_3397,N_3319);
or U3646 (N_3646,N_3312,N_3395);
or U3647 (N_3647,N_3263,N_3369);
nor U3648 (N_3648,N_3375,N_3478);
xor U3649 (N_3649,N_3262,N_3311);
or U3650 (N_3650,N_3254,N_3346);
nand U3651 (N_3651,N_3275,N_3460);
xor U3652 (N_3652,N_3406,N_3342);
nand U3653 (N_3653,N_3292,N_3496);
xnor U3654 (N_3654,N_3307,N_3494);
nor U3655 (N_3655,N_3278,N_3322);
or U3656 (N_3656,N_3301,N_3484);
xnor U3657 (N_3657,N_3342,N_3480);
and U3658 (N_3658,N_3325,N_3345);
and U3659 (N_3659,N_3330,N_3351);
nor U3660 (N_3660,N_3451,N_3424);
nor U3661 (N_3661,N_3269,N_3485);
and U3662 (N_3662,N_3381,N_3272);
xor U3663 (N_3663,N_3476,N_3275);
xnor U3664 (N_3664,N_3416,N_3403);
or U3665 (N_3665,N_3457,N_3345);
nand U3666 (N_3666,N_3390,N_3298);
nand U3667 (N_3667,N_3418,N_3355);
and U3668 (N_3668,N_3400,N_3473);
and U3669 (N_3669,N_3422,N_3269);
nand U3670 (N_3670,N_3388,N_3280);
or U3671 (N_3671,N_3401,N_3306);
nor U3672 (N_3672,N_3467,N_3305);
nand U3673 (N_3673,N_3485,N_3430);
nor U3674 (N_3674,N_3353,N_3453);
nor U3675 (N_3675,N_3275,N_3471);
nor U3676 (N_3676,N_3405,N_3342);
xnor U3677 (N_3677,N_3443,N_3439);
nor U3678 (N_3678,N_3463,N_3289);
nor U3679 (N_3679,N_3351,N_3461);
nand U3680 (N_3680,N_3394,N_3473);
or U3681 (N_3681,N_3389,N_3311);
nor U3682 (N_3682,N_3402,N_3337);
nand U3683 (N_3683,N_3474,N_3400);
and U3684 (N_3684,N_3360,N_3311);
nor U3685 (N_3685,N_3321,N_3273);
and U3686 (N_3686,N_3302,N_3401);
or U3687 (N_3687,N_3437,N_3311);
nor U3688 (N_3688,N_3366,N_3358);
xor U3689 (N_3689,N_3370,N_3292);
or U3690 (N_3690,N_3444,N_3274);
and U3691 (N_3691,N_3296,N_3302);
or U3692 (N_3692,N_3463,N_3471);
or U3693 (N_3693,N_3444,N_3478);
nand U3694 (N_3694,N_3252,N_3382);
nor U3695 (N_3695,N_3271,N_3296);
nor U3696 (N_3696,N_3366,N_3435);
nand U3697 (N_3697,N_3460,N_3323);
and U3698 (N_3698,N_3260,N_3279);
and U3699 (N_3699,N_3395,N_3341);
nor U3700 (N_3700,N_3381,N_3369);
or U3701 (N_3701,N_3341,N_3387);
and U3702 (N_3702,N_3362,N_3406);
or U3703 (N_3703,N_3333,N_3275);
or U3704 (N_3704,N_3393,N_3304);
nor U3705 (N_3705,N_3315,N_3428);
xor U3706 (N_3706,N_3346,N_3459);
nand U3707 (N_3707,N_3304,N_3381);
nand U3708 (N_3708,N_3404,N_3368);
nor U3709 (N_3709,N_3367,N_3354);
xnor U3710 (N_3710,N_3321,N_3258);
or U3711 (N_3711,N_3335,N_3304);
nand U3712 (N_3712,N_3373,N_3411);
and U3713 (N_3713,N_3488,N_3375);
or U3714 (N_3714,N_3265,N_3451);
nor U3715 (N_3715,N_3487,N_3396);
or U3716 (N_3716,N_3389,N_3265);
nor U3717 (N_3717,N_3305,N_3266);
nand U3718 (N_3718,N_3378,N_3474);
xnor U3719 (N_3719,N_3426,N_3481);
or U3720 (N_3720,N_3336,N_3402);
and U3721 (N_3721,N_3340,N_3327);
and U3722 (N_3722,N_3405,N_3435);
nor U3723 (N_3723,N_3436,N_3314);
nand U3724 (N_3724,N_3463,N_3402);
nand U3725 (N_3725,N_3432,N_3444);
nor U3726 (N_3726,N_3392,N_3408);
and U3727 (N_3727,N_3283,N_3499);
and U3728 (N_3728,N_3291,N_3478);
or U3729 (N_3729,N_3353,N_3482);
or U3730 (N_3730,N_3294,N_3384);
nand U3731 (N_3731,N_3374,N_3423);
and U3732 (N_3732,N_3464,N_3391);
nor U3733 (N_3733,N_3460,N_3402);
xor U3734 (N_3734,N_3254,N_3259);
and U3735 (N_3735,N_3251,N_3382);
nand U3736 (N_3736,N_3353,N_3276);
or U3737 (N_3737,N_3493,N_3409);
nand U3738 (N_3738,N_3342,N_3353);
nand U3739 (N_3739,N_3337,N_3356);
nor U3740 (N_3740,N_3297,N_3382);
nor U3741 (N_3741,N_3318,N_3399);
nor U3742 (N_3742,N_3457,N_3469);
nor U3743 (N_3743,N_3429,N_3398);
or U3744 (N_3744,N_3315,N_3348);
and U3745 (N_3745,N_3411,N_3319);
or U3746 (N_3746,N_3405,N_3459);
xor U3747 (N_3747,N_3369,N_3457);
and U3748 (N_3748,N_3281,N_3367);
or U3749 (N_3749,N_3367,N_3456);
and U3750 (N_3750,N_3569,N_3521);
xor U3751 (N_3751,N_3597,N_3552);
and U3752 (N_3752,N_3726,N_3631);
or U3753 (N_3753,N_3624,N_3604);
or U3754 (N_3754,N_3553,N_3584);
xor U3755 (N_3755,N_3705,N_3572);
nor U3756 (N_3756,N_3534,N_3635);
nand U3757 (N_3757,N_3731,N_3659);
xor U3758 (N_3758,N_3746,N_3643);
nor U3759 (N_3759,N_3570,N_3587);
and U3760 (N_3760,N_3546,N_3540);
nand U3761 (N_3761,N_3713,N_3551);
xor U3762 (N_3762,N_3628,N_3532);
nand U3763 (N_3763,N_3655,N_3711);
nor U3764 (N_3764,N_3725,N_3562);
nand U3765 (N_3765,N_3594,N_3672);
and U3766 (N_3766,N_3614,N_3695);
and U3767 (N_3767,N_3727,N_3742);
or U3768 (N_3768,N_3622,N_3679);
and U3769 (N_3769,N_3652,N_3689);
and U3770 (N_3770,N_3688,N_3583);
nor U3771 (N_3771,N_3682,N_3548);
nor U3772 (N_3772,N_3722,N_3729);
or U3773 (N_3773,N_3674,N_3704);
xnor U3774 (N_3774,N_3706,N_3737);
and U3775 (N_3775,N_3611,N_3636);
nor U3776 (N_3776,N_3524,N_3623);
xnor U3777 (N_3777,N_3681,N_3707);
nand U3778 (N_3778,N_3627,N_3533);
nor U3779 (N_3779,N_3686,N_3618);
or U3780 (N_3780,N_3596,N_3621);
nand U3781 (N_3781,N_3511,N_3609);
nor U3782 (N_3782,N_3660,N_3512);
nand U3783 (N_3783,N_3745,N_3556);
or U3784 (N_3784,N_3749,N_3560);
and U3785 (N_3785,N_3700,N_3566);
nand U3786 (N_3786,N_3554,N_3542);
and U3787 (N_3787,N_3740,N_3589);
nor U3788 (N_3788,N_3634,N_3510);
or U3789 (N_3789,N_3644,N_3559);
nand U3790 (N_3790,N_3603,N_3503);
or U3791 (N_3791,N_3638,N_3717);
nor U3792 (N_3792,N_3739,N_3580);
and U3793 (N_3793,N_3616,N_3646);
or U3794 (N_3794,N_3654,N_3502);
and U3795 (N_3795,N_3549,N_3574);
nand U3796 (N_3796,N_3598,N_3736);
or U3797 (N_3797,N_3592,N_3687);
nand U3798 (N_3798,N_3645,N_3617);
and U3799 (N_3799,N_3509,N_3661);
nor U3800 (N_3800,N_3613,N_3665);
nor U3801 (N_3801,N_3642,N_3504);
nand U3802 (N_3802,N_3565,N_3507);
xor U3803 (N_3803,N_3678,N_3667);
nor U3804 (N_3804,N_3730,N_3668);
or U3805 (N_3805,N_3732,N_3670);
or U3806 (N_3806,N_3577,N_3578);
and U3807 (N_3807,N_3608,N_3581);
or U3808 (N_3808,N_3520,N_3639);
nor U3809 (N_3809,N_3517,N_3538);
or U3810 (N_3810,N_3610,N_3514);
nand U3811 (N_3811,N_3516,N_3649);
or U3812 (N_3812,N_3664,N_3710);
nand U3813 (N_3813,N_3677,N_3691);
xnor U3814 (N_3814,N_3747,N_3696);
nand U3815 (N_3815,N_3709,N_3666);
or U3816 (N_3816,N_3724,N_3653);
nor U3817 (N_3817,N_3723,N_3568);
nor U3818 (N_3818,N_3573,N_3586);
nand U3819 (N_3819,N_3536,N_3529);
nand U3820 (N_3820,N_3637,N_3715);
and U3821 (N_3821,N_3515,N_3721);
xor U3822 (N_3822,N_3625,N_3530);
xnor U3823 (N_3823,N_3694,N_3734);
and U3824 (N_3824,N_3693,N_3523);
nor U3825 (N_3825,N_3685,N_3738);
xor U3826 (N_3826,N_3571,N_3720);
or U3827 (N_3827,N_3605,N_3513);
or U3828 (N_3828,N_3719,N_3733);
nor U3829 (N_3829,N_3541,N_3663);
or U3830 (N_3830,N_3683,N_3545);
xor U3831 (N_3831,N_3590,N_3528);
nand U3832 (N_3832,N_3650,N_3599);
xnor U3833 (N_3833,N_3575,N_3714);
xnor U3834 (N_3834,N_3595,N_3676);
nand U3835 (N_3835,N_3585,N_3718);
or U3836 (N_3836,N_3539,N_3647);
nor U3837 (N_3837,N_3632,N_3531);
or U3838 (N_3838,N_3684,N_3601);
nor U3839 (N_3839,N_3582,N_3669);
nor U3840 (N_3840,N_3527,N_3630);
or U3841 (N_3841,N_3612,N_3716);
or U3842 (N_3842,N_3526,N_3748);
nand U3843 (N_3843,N_3697,N_3712);
and U3844 (N_3844,N_3544,N_3550);
or U3845 (N_3845,N_3519,N_3701);
and U3846 (N_3846,N_3626,N_3558);
or U3847 (N_3847,N_3698,N_3563);
nor U3848 (N_3848,N_3702,N_3699);
or U3849 (N_3849,N_3620,N_3588);
and U3850 (N_3850,N_3567,N_3657);
and U3851 (N_3851,N_3607,N_3506);
nor U3852 (N_3852,N_3651,N_3537);
nand U3853 (N_3853,N_3505,N_3535);
nand U3854 (N_3854,N_3576,N_3675);
and U3855 (N_3855,N_3602,N_3518);
nand U3856 (N_3856,N_3640,N_3547);
nand U3857 (N_3857,N_3615,N_3692);
or U3858 (N_3858,N_3593,N_3600);
or U3859 (N_3859,N_3508,N_3501);
nand U3860 (N_3860,N_3591,N_3579);
nor U3861 (N_3861,N_3561,N_3671);
or U3862 (N_3862,N_3633,N_3662);
or U3863 (N_3863,N_3690,N_3656);
nor U3864 (N_3864,N_3743,N_3564);
or U3865 (N_3865,N_3522,N_3741);
and U3866 (N_3866,N_3500,N_3703);
and U3867 (N_3867,N_3680,N_3658);
nand U3868 (N_3868,N_3555,N_3744);
nor U3869 (N_3869,N_3641,N_3648);
and U3870 (N_3870,N_3543,N_3708);
and U3871 (N_3871,N_3728,N_3619);
nand U3872 (N_3872,N_3735,N_3673);
nand U3873 (N_3873,N_3557,N_3629);
nand U3874 (N_3874,N_3525,N_3606);
and U3875 (N_3875,N_3522,N_3633);
or U3876 (N_3876,N_3716,N_3579);
and U3877 (N_3877,N_3509,N_3701);
or U3878 (N_3878,N_3672,N_3659);
and U3879 (N_3879,N_3726,N_3573);
nand U3880 (N_3880,N_3703,N_3675);
nor U3881 (N_3881,N_3667,N_3657);
nor U3882 (N_3882,N_3595,N_3594);
xor U3883 (N_3883,N_3693,N_3712);
xor U3884 (N_3884,N_3605,N_3717);
or U3885 (N_3885,N_3553,N_3587);
nand U3886 (N_3886,N_3666,N_3534);
or U3887 (N_3887,N_3696,N_3649);
and U3888 (N_3888,N_3678,N_3564);
nor U3889 (N_3889,N_3663,N_3565);
and U3890 (N_3890,N_3609,N_3729);
nor U3891 (N_3891,N_3720,N_3575);
and U3892 (N_3892,N_3545,N_3738);
nor U3893 (N_3893,N_3602,N_3624);
xnor U3894 (N_3894,N_3623,N_3631);
and U3895 (N_3895,N_3506,N_3620);
or U3896 (N_3896,N_3568,N_3744);
or U3897 (N_3897,N_3526,N_3749);
nand U3898 (N_3898,N_3634,N_3549);
nand U3899 (N_3899,N_3638,N_3541);
nor U3900 (N_3900,N_3553,N_3695);
and U3901 (N_3901,N_3723,N_3735);
and U3902 (N_3902,N_3617,N_3565);
nor U3903 (N_3903,N_3627,N_3654);
nand U3904 (N_3904,N_3588,N_3554);
nor U3905 (N_3905,N_3553,N_3562);
and U3906 (N_3906,N_3728,N_3729);
nor U3907 (N_3907,N_3601,N_3673);
nand U3908 (N_3908,N_3683,N_3563);
nor U3909 (N_3909,N_3673,N_3606);
nor U3910 (N_3910,N_3543,N_3679);
nor U3911 (N_3911,N_3614,N_3512);
and U3912 (N_3912,N_3725,N_3584);
nand U3913 (N_3913,N_3591,N_3745);
nand U3914 (N_3914,N_3542,N_3560);
xor U3915 (N_3915,N_3677,N_3580);
nor U3916 (N_3916,N_3539,N_3526);
or U3917 (N_3917,N_3553,N_3697);
and U3918 (N_3918,N_3563,N_3700);
or U3919 (N_3919,N_3675,N_3628);
and U3920 (N_3920,N_3591,N_3644);
and U3921 (N_3921,N_3524,N_3520);
nand U3922 (N_3922,N_3562,N_3561);
or U3923 (N_3923,N_3563,N_3733);
nand U3924 (N_3924,N_3620,N_3563);
or U3925 (N_3925,N_3709,N_3600);
nor U3926 (N_3926,N_3672,N_3611);
and U3927 (N_3927,N_3631,N_3716);
nand U3928 (N_3928,N_3639,N_3637);
or U3929 (N_3929,N_3742,N_3652);
xor U3930 (N_3930,N_3589,N_3704);
nand U3931 (N_3931,N_3632,N_3511);
and U3932 (N_3932,N_3512,N_3609);
or U3933 (N_3933,N_3521,N_3559);
and U3934 (N_3934,N_3514,N_3619);
or U3935 (N_3935,N_3697,N_3534);
or U3936 (N_3936,N_3658,N_3707);
and U3937 (N_3937,N_3733,N_3523);
xnor U3938 (N_3938,N_3583,N_3599);
nand U3939 (N_3939,N_3639,N_3601);
or U3940 (N_3940,N_3746,N_3543);
nor U3941 (N_3941,N_3685,N_3736);
nand U3942 (N_3942,N_3671,N_3508);
nor U3943 (N_3943,N_3543,N_3706);
nor U3944 (N_3944,N_3659,N_3704);
nand U3945 (N_3945,N_3503,N_3615);
or U3946 (N_3946,N_3713,N_3637);
xor U3947 (N_3947,N_3511,N_3655);
nor U3948 (N_3948,N_3570,N_3689);
and U3949 (N_3949,N_3526,N_3655);
or U3950 (N_3950,N_3690,N_3632);
and U3951 (N_3951,N_3625,N_3626);
and U3952 (N_3952,N_3635,N_3741);
and U3953 (N_3953,N_3707,N_3573);
nor U3954 (N_3954,N_3508,N_3611);
or U3955 (N_3955,N_3731,N_3730);
nand U3956 (N_3956,N_3593,N_3738);
nor U3957 (N_3957,N_3561,N_3739);
nor U3958 (N_3958,N_3736,N_3623);
nor U3959 (N_3959,N_3531,N_3568);
nor U3960 (N_3960,N_3519,N_3625);
xor U3961 (N_3961,N_3570,N_3584);
and U3962 (N_3962,N_3565,N_3722);
xor U3963 (N_3963,N_3666,N_3547);
and U3964 (N_3964,N_3746,N_3610);
and U3965 (N_3965,N_3624,N_3730);
nand U3966 (N_3966,N_3737,N_3597);
or U3967 (N_3967,N_3673,N_3745);
nor U3968 (N_3968,N_3662,N_3542);
or U3969 (N_3969,N_3686,N_3733);
nor U3970 (N_3970,N_3690,N_3695);
nand U3971 (N_3971,N_3583,N_3586);
and U3972 (N_3972,N_3530,N_3721);
nand U3973 (N_3973,N_3531,N_3661);
and U3974 (N_3974,N_3593,N_3584);
or U3975 (N_3975,N_3514,N_3729);
and U3976 (N_3976,N_3662,N_3522);
or U3977 (N_3977,N_3633,N_3692);
or U3978 (N_3978,N_3693,N_3727);
nor U3979 (N_3979,N_3567,N_3708);
nand U3980 (N_3980,N_3709,N_3570);
or U3981 (N_3981,N_3675,N_3695);
nor U3982 (N_3982,N_3657,N_3597);
and U3983 (N_3983,N_3521,N_3607);
nand U3984 (N_3984,N_3582,N_3634);
or U3985 (N_3985,N_3606,N_3517);
or U3986 (N_3986,N_3572,N_3742);
and U3987 (N_3987,N_3610,N_3555);
nand U3988 (N_3988,N_3629,N_3534);
or U3989 (N_3989,N_3689,N_3657);
and U3990 (N_3990,N_3534,N_3700);
or U3991 (N_3991,N_3600,N_3741);
nor U3992 (N_3992,N_3537,N_3504);
or U3993 (N_3993,N_3740,N_3528);
and U3994 (N_3994,N_3716,N_3707);
nor U3995 (N_3995,N_3558,N_3529);
xor U3996 (N_3996,N_3728,N_3627);
nand U3997 (N_3997,N_3521,N_3640);
or U3998 (N_3998,N_3533,N_3561);
or U3999 (N_3999,N_3523,N_3644);
nand U4000 (N_4000,N_3911,N_3872);
and U4001 (N_4001,N_3853,N_3752);
and U4002 (N_4002,N_3836,N_3763);
nor U4003 (N_4003,N_3985,N_3941);
nor U4004 (N_4004,N_3901,N_3775);
and U4005 (N_4005,N_3935,N_3999);
nand U4006 (N_4006,N_3802,N_3788);
or U4007 (N_4007,N_3975,N_3857);
nor U4008 (N_4008,N_3793,N_3767);
and U4009 (N_4009,N_3869,N_3914);
or U4010 (N_4010,N_3990,N_3821);
nor U4011 (N_4011,N_3844,N_3795);
nor U4012 (N_4012,N_3863,N_3895);
nor U4013 (N_4013,N_3867,N_3979);
or U4014 (N_4014,N_3851,N_3965);
nor U4015 (N_4015,N_3797,N_3826);
xor U4016 (N_4016,N_3924,N_3960);
nor U4017 (N_4017,N_3873,N_3774);
nor U4018 (N_4018,N_3839,N_3982);
and U4019 (N_4019,N_3959,N_3784);
and U4020 (N_4020,N_3886,N_3879);
and U4021 (N_4021,N_3799,N_3884);
xor U4022 (N_4022,N_3829,N_3903);
nand U4023 (N_4023,N_3807,N_3991);
and U4024 (N_4024,N_3865,N_3974);
nor U4025 (N_4025,N_3871,N_3880);
nor U4026 (N_4026,N_3943,N_3904);
nor U4027 (N_4027,N_3925,N_3921);
nand U4028 (N_4028,N_3846,N_3868);
or U4029 (N_4029,N_3824,N_3957);
nand U4030 (N_4030,N_3980,N_3930);
nor U4031 (N_4031,N_3951,N_3874);
nor U4032 (N_4032,N_3781,N_3801);
nand U4033 (N_4033,N_3971,N_3758);
and U4034 (N_4034,N_3998,N_3968);
nor U4035 (N_4035,N_3885,N_3918);
nor U4036 (N_4036,N_3814,N_3757);
and U4037 (N_4037,N_3907,N_3997);
nor U4038 (N_4038,N_3789,N_3768);
xnor U4039 (N_4039,N_3771,N_3927);
and U4040 (N_4040,N_3843,N_3913);
nand U4041 (N_4041,N_3803,N_3915);
or U4042 (N_4042,N_3820,N_3887);
or U4043 (N_4043,N_3861,N_3766);
xor U4044 (N_4044,N_3894,N_3977);
xor U4045 (N_4045,N_3806,N_3950);
and U4046 (N_4046,N_3779,N_3899);
nand U4047 (N_4047,N_3883,N_3892);
nand U4048 (N_4048,N_3944,N_3772);
nor U4049 (N_4049,N_3856,N_3852);
and U4050 (N_4050,N_3822,N_3841);
and U4051 (N_4051,N_3833,N_3966);
or U4052 (N_4052,N_3945,N_3791);
nand U4053 (N_4053,N_3770,N_3931);
xnor U4054 (N_4054,N_3818,N_3860);
or U4055 (N_4055,N_3922,N_3961);
or U4056 (N_4056,N_3900,N_3854);
nand U4057 (N_4057,N_3858,N_3984);
nand U4058 (N_4058,N_3993,N_3926);
nor U4059 (N_4059,N_3783,N_3923);
and U4060 (N_4060,N_3952,N_3988);
nor U4061 (N_4061,N_3849,N_3798);
nand U4062 (N_4062,N_3811,N_3905);
nand U4063 (N_4063,N_3896,N_3889);
nand U4064 (N_4064,N_3987,N_3906);
nand U4065 (N_4065,N_3762,N_3756);
and U4066 (N_4066,N_3837,N_3759);
nand U4067 (N_4067,N_3776,N_3850);
and U4068 (N_4068,N_3996,N_3992);
or U4069 (N_4069,N_3765,N_3898);
or U4070 (N_4070,N_3875,N_3912);
and U4071 (N_4071,N_3817,N_3809);
nand U4072 (N_4072,N_3981,N_3815);
or U4073 (N_4073,N_3840,N_3755);
nand U4074 (N_4074,N_3787,N_3964);
xnor U4075 (N_4075,N_3972,N_3777);
and U4076 (N_4076,N_3835,N_3902);
or U4077 (N_4077,N_3859,N_3819);
or U4078 (N_4078,N_3893,N_3928);
nand U4079 (N_4079,N_3954,N_3995);
xor U4080 (N_4080,N_3769,N_3751);
xor U4081 (N_4081,N_3816,N_3813);
xnor U4082 (N_4082,N_3761,N_3862);
nand U4083 (N_4083,N_3848,N_3949);
or U4084 (N_4084,N_3866,N_3828);
nand U4085 (N_4085,N_3780,N_3934);
nor U4086 (N_4086,N_3804,N_3973);
nor U4087 (N_4087,N_3908,N_3834);
or U4088 (N_4088,N_3963,N_3754);
xor U4089 (N_4089,N_3897,N_3986);
nand U4090 (N_4090,N_3842,N_3810);
nand U4091 (N_4091,N_3882,N_3823);
nor U4092 (N_4092,N_3870,N_3792);
nor U4093 (N_4093,N_3910,N_3794);
nor U4094 (N_4094,N_3929,N_3920);
and U4095 (N_4095,N_3778,N_3946);
nor U4096 (N_4096,N_3845,N_3962);
nor U4097 (N_4097,N_3838,N_3937);
nand U4098 (N_4098,N_3994,N_3936);
nor U4099 (N_4099,N_3890,N_3948);
nand U4100 (N_4100,N_3933,N_3753);
or U4101 (N_4101,N_3881,N_3891);
and U4102 (N_4102,N_3967,N_3938);
nor U4103 (N_4103,N_3983,N_3830);
nand U4104 (N_4104,N_3953,N_3760);
nor U4105 (N_4105,N_3947,N_3989);
nor U4106 (N_4106,N_3969,N_3825);
or U4107 (N_4107,N_3909,N_3878);
nor U4108 (N_4108,N_3831,N_3976);
or U4109 (N_4109,N_3796,N_3855);
nand U4110 (N_4110,N_3773,N_3764);
nand U4111 (N_4111,N_3955,N_3942);
xor U4112 (N_4112,N_3940,N_3919);
and U4113 (N_4113,N_3970,N_3876);
nor U4114 (N_4114,N_3808,N_3958);
nand U4115 (N_4115,N_3785,N_3750);
or U4116 (N_4116,N_3864,N_3782);
nor U4117 (N_4117,N_3790,N_3978);
and U4118 (N_4118,N_3917,N_3847);
nand U4119 (N_4119,N_3832,N_3786);
nor U4120 (N_4120,N_3888,N_3877);
nor U4121 (N_4121,N_3805,N_3956);
or U4122 (N_4122,N_3827,N_3800);
xnor U4123 (N_4123,N_3939,N_3812);
and U4124 (N_4124,N_3932,N_3916);
and U4125 (N_4125,N_3916,N_3853);
nand U4126 (N_4126,N_3834,N_3989);
or U4127 (N_4127,N_3933,N_3839);
or U4128 (N_4128,N_3934,N_3871);
and U4129 (N_4129,N_3778,N_3804);
nand U4130 (N_4130,N_3941,N_3752);
or U4131 (N_4131,N_3953,N_3979);
or U4132 (N_4132,N_3949,N_3893);
and U4133 (N_4133,N_3917,N_3923);
and U4134 (N_4134,N_3998,N_3938);
or U4135 (N_4135,N_3808,N_3842);
nor U4136 (N_4136,N_3816,N_3764);
nor U4137 (N_4137,N_3942,N_3958);
or U4138 (N_4138,N_3752,N_3816);
nor U4139 (N_4139,N_3978,N_3898);
xnor U4140 (N_4140,N_3841,N_3750);
or U4141 (N_4141,N_3922,N_3987);
nand U4142 (N_4142,N_3884,N_3984);
nand U4143 (N_4143,N_3958,N_3907);
and U4144 (N_4144,N_3850,N_3894);
nand U4145 (N_4145,N_3882,N_3921);
nor U4146 (N_4146,N_3911,N_3975);
and U4147 (N_4147,N_3768,N_3890);
or U4148 (N_4148,N_3924,N_3889);
nand U4149 (N_4149,N_3815,N_3974);
nor U4150 (N_4150,N_3850,N_3751);
nand U4151 (N_4151,N_3912,N_3804);
nand U4152 (N_4152,N_3944,N_3851);
xor U4153 (N_4153,N_3962,N_3763);
nand U4154 (N_4154,N_3940,N_3917);
nor U4155 (N_4155,N_3801,N_3778);
and U4156 (N_4156,N_3791,N_3897);
and U4157 (N_4157,N_3765,N_3999);
nand U4158 (N_4158,N_3855,N_3902);
and U4159 (N_4159,N_3975,N_3791);
nand U4160 (N_4160,N_3994,N_3784);
nor U4161 (N_4161,N_3781,N_3939);
nor U4162 (N_4162,N_3756,N_3967);
nand U4163 (N_4163,N_3870,N_3969);
xor U4164 (N_4164,N_3784,N_3848);
and U4165 (N_4165,N_3781,N_3965);
nand U4166 (N_4166,N_3905,N_3886);
or U4167 (N_4167,N_3772,N_3948);
or U4168 (N_4168,N_3757,N_3790);
nor U4169 (N_4169,N_3853,N_3825);
nor U4170 (N_4170,N_3981,N_3971);
or U4171 (N_4171,N_3872,N_3821);
and U4172 (N_4172,N_3851,N_3834);
or U4173 (N_4173,N_3793,N_3835);
or U4174 (N_4174,N_3997,N_3862);
or U4175 (N_4175,N_3815,N_3792);
or U4176 (N_4176,N_3928,N_3975);
nand U4177 (N_4177,N_3952,N_3779);
nor U4178 (N_4178,N_3809,N_3770);
nand U4179 (N_4179,N_3787,N_3851);
and U4180 (N_4180,N_3810,N_3938);
nand U4181 (N_4181,N_3900,N_3752);
xor U4182 (N_4182,N_3752,N_3833);
or U4183 (N_4183,N_3859,N_3972);
xor U4184 (N_4184,N_3886,N_3977);
xnor U4185 (N_4185,N_3851,N_3991);
or U4186 (N_4186,N_3755,N_3939);
and U4187 (N_4187,N_3984,N_3792);
or U4188 (N_4188,N_3964,N_3907);
or U4189 (N_4189,N_3814,N_3798);
and U4190 (N_4190,N_3917,N_3778);
nor U4191 (N_4191,N_3868,N_3982);
nand U4192 (N_4192,N_3879,N_3866);
nand U4193 (N_4193,N_3826,N_3778);
and U4194 (N_4194,N_3866,N_3784);
nor U4195 (N_4195,N_3789,N_3872);
xnor U4196 (N_4196,N_3979,N_3986);
or U4197 (N_4197,N_3819,N_3928);
and U4198 (N_4198,N_3979,N_3933);
and U4199 (N_4199,N_3873,N_3843);
nor U4200 (N_4200,N_3826,N_3819);
nand U4201 (N_4201,N_3864,N_3784);
nand U4202 (N_4202,N_3903,N_3900);
and U4203 (N_4203,N_3798,N_3765);
nor U4204 (N_4204,N_3828,N_3802);
nor U4205 (N_4205,N_3856,N_3980);
or U4206 (N_4206,N_3840,N_3821);
nor U4207 (N_4207,N_3983,N_3986);
nor U4208 (N_4208,N_3792,N_3976);
nor U4209 (N_4209,N_3870,N_3785);
nand U4210 (N_4210,N_3968,N_3980);
or U4211 (N_4211,N_3867,N_3769);
and U4212 (N_4212,N_3981,N_3763);
or U4213 (N_4213,N_3865,N_3925);
or U4214 (N_4214,N_3983,N_3816);
and U4215 (N_4215,N_3967,N_3838);
nor U4216 (N_4216,N_3784,N_3787);
or U4217 (N_4217,N_3858,N_3811);
nand U4218 (N_4218,N_3754,N_3872);
or U4219 (N_4219,N_3773,N_3931);
nor U4220 (N_4220,N_3877,N_3751);
nor U4221 (N_4221,N_3879,N_3758);
nand U4222 (N_4222,N_3780,N_3879);
or U4223 (N_4223,N_3956,N_3757);
or U4224 (N_4224,N_3892,N_3797);
nand U4225 (N_4225,N_3979,N_3814);
or U4226 (N_4226,N_3999,N_3930);
nor U4227 (N_4227,N_3974,N_3789);
nand U4228 (N_4228,N_3826,N_3852);
and U4229 (N_4229,N_3932,N_3984);
nor U4230 (N_4230,N_3958,N_3906);
and U4231 (N_4231,N_3895,N_3969);
and U4232 (N_4232,N_3763,N_3786);
or U4233 (N_4233,N_3784,N_3883);
nand U4234 (N_4234,N_3803,N_3907);
xor U4235 (N_4235,N_3955,N_3793);
xnor U4236 (N_4236,N_3894,N_3777);
and U4237 (N_4237,N_3768,N_3829);
and U4238 (N_4238,N_3989,N_3899);
and U4239 (N_4239,N_3769,N_3907);
xnor U4240 (N_4240,N_3939,N_3918);
xor U4241 (N_4241,N_3963,N_3836);
and U4242 (N_4242,N_3977,N_3838);
nor U4243 (N_4243,N_3779,N_3949);
xnor U4244 (N_4244,N_3784,N_3804);
nand U4245 (N_4245,N_3881,N_3828);
nor U4246 (N_4246,N_3764,N_3762);
and U4247 (N_4247,N_3823,N_3954);
and U4248 (N_4248,N_3775,N_3790);
or U4249 (N_4249,N_3907,N_3974);
nand U4250 (N_4250,N_4187,N_4116);
nand U4251 (N_4251,N_4146,N_4021);
nor U4252 (N_4252,N_4121,N_4211);
nor U4253 (N_4253,N_4096,N_4230);
nand U4254 (N_4254,N_4088,N_4022);
and U4255 (N_4255,N_4157,N_4115);
nor U4256 (N_4256,N_4108,N_4225);
and U4257 (N_4257,N_4140,N_4165);
xnor U4258 (N_4258,N_4171,N_4052);
nor U4259 (N_4259,N_4010,N_4164);
or U4260 (N_4260,N_4085,N_4014);
nor U4261 (N_4261,N_4122,N_4217);
nand U4262 (N_4262,N_4200,N_4007);
nor U4263 (N_4263,N_4031,N_4128);
nand U4264 (N_4264,N_4219,N_4240);
or U4265 (N_4265,N_4023,N_4113);
nor U4266 (N_4266,N_4106,N_4220);
or U4267 (N_4267,N_4001,N_4068);
or U4268 (N_4268,N_4170,N_4124);
nor U4269 (N_4269,N_4098,N_4097);
nor U4270 (N_4270,N_4195,N_4210);
and U4271 (N_4271,N_4233,N_4125);
and U4272 (N_4272,N_4047,N_4180);
nor U4273 (N_4273,N_4107,N_4150);
nand U4274 (N_4274,N_4201,N_4119);
nor U4275 (N_4275,N_4015,N_4175);
or U4276 (N_4276,N_4109,N_4101);
nor U4277 (N_4277,N_4199,N_4186);
nor U4278 (N_4278,N_4004,N_4080);
nand U4279 (N_4279,N_4244,N_4030);
or U4280 (N_4280,N_4154,N_4159);
and U4281 (N_4281,N_4102,N_4167);
and U4282 (N_4282,N_4188,N_4087);
nor U4283 (N_4283,N_4055,N_4151);
or U4284 (N_4284,N_4215,N_4092);
xor U4285 (N_4285,N_4099,N_4218);
and U4286 (N_4286,N_4232,N_4148);
nand U4287 (N_4287,N_4060,N_4064);
and U4288 (N_4288,N_4105,N_4011);
nor U4289 (N_4289,N_4002,N_4174);
nor U4290 (N_4290,N_4071,N_4182);
nor U4291 (N_4291,N_4231,N_4212);
nand U4292 (N_4292,N_4197,N_4178);
and U4293 (N_4293,N_4156,N_4049);
and U4294 (N_4294,N_4062,N_4142);
nor U4295 (N_4295,N_4027,N_4053);
or U4296 (N_4296,N_4246,N_4091);
nand U4297 (N_4297,N_4050,N_4051);
and U4298 (N_4298,N_4003,N_4089);
nor U4299 (N_4299,N_4247,N_4183);
nand U4300 (N_4300,N_4249,N_4077);
and U4301 (N_4301,N_4192,N_4173);
nand U4302 (N_4302,N_4228,N_4054);
and U4303 (N_4303,N_4090,N_4082);
nor U4304 (N_4304,N_4118,N_4185);
nand U4305 (N_4305,N_4209,N_4086);
nor U4306 (N_4306,N_4202,N_4074);
nand U4307 (N_4307,N_4243,N_4226);
or U4308 (N_4308,N_4227,N_4206);
nor U4309 (N_4309,N_4069,N_4032);
or U4310 (N_4310,N_4073,N_4078);
or U4311 (N_4311,N_4234,N_4061);
and U4312 (N_4312,N_4149,N_4035);
or U4313 (N_4313,N_4045,N_4152);
nand U4314 (N_4314,N_4036,N_4133);
and U4315 (N_4315,N_4114,N_4057);
nor U4316 (N_4316,N_4044,N_4155);
or U4317 (N_4317,N_4039,N_4138);
and U4318 (N_4318,N_4163,N_4239);
nor U4319 (N_4319,N_4016,N_4205);
and U4320 (N_4320,N_4213,N_4093);
xnor U4321 (N_4321,N_4123,N_4241);
nor U4322 (N_4322,N_4132,N_4198);
nand U4323 (N_4323,N_4075,N_4141);
nor U4324 (N_4324,N_4134,N_4110);
xor U4325 (N_4325,N_4196,N_4166);
and U4326 (N_4326,N_4139,N_4059);
and U4327 (N_4327,N_4079,N_4177);
nor U4328 (N_4328,N_4029,N_4076);
or U4329 (N_4329,N_4037,N_4137);
or U4330 (N_4330,N_4147,N_4203);
xnor U4331 (N_4331,N_4019,N_4158);
nand U4332 (N_4332,N_4094,N_4190);
or U4333 (N_4333,N_4048,N_4103);
and U4334 (N_4334,N_4236,N_4008);
and U4335 (N_4335,N_4025,N_4081);
nor U4336 (N_4336,N_4120,N_4070);
or U4337 (N_4337,N_4006,N_4179);
and U4338 (N_4338,N_4130,N_4235);
or U4339 (N_4339,N_4018,N_4135);
and U4340 (N_4340,N_4204,N_4127);
xor U4341 (N_4341,N_4160,N_4034);
nand U4342 (N_4342,N_4012,N_4238);
nand U4343 (N_4343,N_4143,N_4013);
or U4344 (N_4344,N_4112,N_4066);
and U4345 (N_4345,N_4153,N_4028);
nand U4346 (N_4346,N_4193,N_4005);
nor U4347 (N_4347,N_4046,N_4020);
nor U4348 (N_4348,N_4168,N_4058);
and U4349 (N_4349,N_4009,N_4095);
nor U4350 (N_4350,N_4017,N_4026);
nand U4351 (N_4351,N_4056,N_4194);
nand U4352 (N_4352,N_4043,N_4131);
nand U4353 (N_4353,N_4136,N_4191);
nor U4354 (N_4354,N_4072,N_4224);
xnor U4355 (N_4355,N_4126,N_4214);
and U4356 (N_4356,N_4242,N_4000);
xnor U4357 (N_4357,N_4189,N_4222);
xnor U4358 (N_4358,N_4176,N_4162);
and U4359 (N_4359,N_4111,N_4229);
and U4360 (N_4360,N_4129,N_4223);
and U4361 (N_4361,N_4083,N_4207);
and U4362 (N_4362,N_4145,N_4038);
nand U4363 (N_4363,N_4245,N_4169);
xnor U4364 (N_4364,N_4067,N_4172);
and U4365 (N_4365,N_4181,N_4216);
xor U4366 (N_4366,N_4065,N_4184);
xnor U4367 (N_4367,N_4041,N_4024);
xnor U4368 (N_4368,N_4237,N_4161);
or U4369 (N_4369,N_4104,N_4033);
nor U4370 (N_4370,N_4117,N_4084);
xnor U4371 (N_4371,N_4208,N_4040);
xor U4372 (N_4372,N_4042,N_4248);
nor U4373 (N_4373,N_4100,N_4063);
xnor U4374 (N_4374,N_4221,N_4144);
nor U4375 (N_4375,N_4108,N_4150);
nand U4376 (N_4376,N_4208,N_4214);
and U4377 (N_4377,N_4015,N_4100);
or U4378 (N_4378,N_4152,N_4168);
nand U4379 (N_4379,N_4115,N_4201);
nor U4380 (N_4380,N_4202,N_4223);
and U4381 (N_4381,N_4103,N_4238);
nand U4382 (N_4382,N_4196,N_4126);
xor U4383 (N_4383,N_4131,N_4067);
and U4384 (N_4384,N_4067,N_4194);
nand U4385 (N_4385,N_4083,N_4179);
nor U4386 (N_4386,N_4126,N_4216);
or U4387 (N_4387,N_4082,N_4098);
xnor U4388 (N_4388,N_4058,N_4017);
nor U4389 (N_4389,N_4150,N_4075);
and U4390 (N_4390,N_4102,N_4141);
nand U4391 (N_4391,N_4236,N_4111);
and U4392 (N_4392,N_4177,N_4227);
xor U4393 (N_4393,N_4084,N_4180);
nand U4394 (N_4394,N_4244,N_4120);
or U4395 (N_4395,N_4090,N_4044);
and U4396 (N_4396,N_4153,N_4139);
nand U4397 (N_4397,N_4213,N_4001);
and U4398 (N_4398,N_4179,N_4227);
or U4399 (N_4399,N_4061,N_4238);
nand U4400 (N_4400,N_4055,N_4088);
nand U4401 (N_4401,N_4162,N_4167);
nor U4402 (N_4402,N_4192,N_4124);
or U4403 (N_4403,N_4161,N_4201);
and U4404 (N_4404,N_4177,N_4138);
nand U4405 (N_4405,N_4170,N_4043);
nand U4406 (N_4406,N_4008,N_4173);
nand U4407 (N_4407,N_4144,N_4117);
nand U4408 (N_4408,N_4183,N_4225);
or U4409 (N_4409,N_4143,N_4101);
or U4410 (N_4410,N_4204,N_4108);
or U4411 (N_4411,N_4045,N_4154);
and U4412 (N_4412,N_4093,N_4075);
and U4413 (N_4413,N_4112,N_4001);
or U4414 (N_4414,N_4015,N_4153);
nor U4415 (N_4415,N_4078,N_4197);
nand U4416 (N_4416,N_4190,N_4027);
and U4417 (N_4417,N_4248,N_4039);
and U4418 (N_4418,N_4078,N_4195);
nor U4419 (N_4419,N_4184,N_4168);
nand U4420 (N_4420,N_4166,N_4181);
nand U4421 (N_4421,N_4144,N_4235);
or U4422 (N_4422,N_4159,N_4202);
xnor U4423 (N_4423,N_4144,N_4028);
and U4424 (N_4424,N_4074,N_4234);
nor U4425 (N_4425,N_4230,N_4018);
nand U4426 (N_4426,N_4042,N_4125);
nand U4427 (N_4427,N_4106,N_4149);
nor U4428 (N_4428,N_4015,N_4209);
and U4429 (N_4429,N_4113,N_4000);
nor U4430 (N_4430,N_4247,N_4136);
nand U4431 (N_4431,N_4021,N_4196);
and U4432 (N_4432,N_4143,N_4165);
nand U4433 (N_4433,N_4157,N_4190);
or U4434 (N_4434,N_4122,N_4158);
and U4435 (N_4435,N_4084,N_4098);
and U4436 (N_4436,N_4129,N_4077);
nor U4437 (N_4437,N_4244,N_4164);
xnor U4438 (N_4438,N_4001,N_4212);
or U4439 (N_4439,N_4087,N_4054);
or U4440 (N_4440,N_4093,N_4131);
nand U4441 (N_4441,N_4095,N_4144);
nand U4442 (N_4442,N_4046,N_4160);
nor U4443 (N_4443,N_4028,N_4133);
nand U4444 (N_4444,N_4217,N_4099);
nor U4445 (N_4445,N_4107,N_4156);
xnor U4446 (N_4446,N_4071,N_4004);
nor U4447 (N_4447,N_4170,N_4207);
nor U4448 (N_4448,N_4164,N_4192);
and U4449 (N_4449,N_4106,N_4047);
nand U4450 (N_4450,N_4249,N_4216);
nor U4451 (N_4451,N_4200,N_4141);
nor U4452 (N_4452,N_4138,N_4097);
and U4453 (N_4453,N_4138,N_4223);
nor U4454 (N_4454,N_4013,N_4168);
xor U4455 (N_4455,N_4142,N_4207);
nor U4456 (N_4456,N_4111,N_4009);
nand U4457 (N_4457,N_4082,N_4065);
xor U4458 (N_4458,N_4116,N_4017);
or U4459 (N_4459,N_4206,N_4008);
or U4460 (N_4460,N_4037,N_4066);
xor U4461 (N_4461,N_4237,N_4132);
and U4462 (N_4462,N_4142,N_4064);
nor U4463 (N_4463,N_4170,N_4139);
and U4464 (N_4464,N_4181,N_4227);
or U4465 (N_4465,N_4201,N_4027);
nor U4466 (N_4466,N_4077,N_4237);
or U4467 (N_4467,N_4072,N_4060);
nor U4468 (N_4468,N_4121,N_4226);
nor U4469 (N_4469,N_4037,N_4176);
nand U4470 (N_4470,N_4025,N_4196);
nand U4471 (N_4471,N_4126,N_4042);
or U4472 (N_4472,N_4005,N_4039);
and U4473 (N_4473,N_4146,N_4190);
xnor U4474 (N_4474,N_4198,N_4206);
nor U4475 (N_4475,N_4010,N_4056);
or U4476 (N_4476,N_4181,N_4240);
nor U4477 (N_4477,N_4208,N_4050);
and U4478 (N_4478,N_4136,N_4057);
nor U4479 (N_4479,N_4054,N_4166);
nor U4480 (N_4480,N_4220,N_4024);
xnor U4481 (N_4481,N_4100,N_4212);
or U4482 (N_4482,N_4212,N_4144);
nor U4483 (N_4483,N_4216,N_4134);
nand U4484 (N_4484,N_4132,N_4077);
nand U4485 (N_4485,N_4203,N_4168);
nor U4486 (N_4486,N_4056,N_4162);
or U4487 (N_4487,N_4135,N_4026);
or U4488 (N_4488,N_4158,N_4200);
nor U4489 (N_4489,N_4104,N_4170);
and U4490 (N_4490,N_4071,N_4094);
or U4491 (N_4491,N_4153,N_4013);
or U4492 (N_4492,N_4097,N_4023);
nor U4493 (N_4493,N_4128,N_4190);
and U4494 (N_4494,N_4094,N_4237);
or U4495 (N_4495,N_4045,N_4218);
nand U4496 (N_4496,N_4026,N_4128);
nor U4497 (N_4497,N_4072,N_4226);
xor U4498 (N_4498,N_4132,N_4232);
and U4499 (N_4499,N_4070,N_4203);
or U4500 (N_4500,N_4325,N_4327);
or U4501 (N_4501,N_4320,N_4472);
nor U4502 (N_4502,N_4411,N_4297);
nand U4503 (N_4503,N_4289,N_4313);
nand U4504 (N_4504,N_4401,N_4268);
nor U4505 (N_4505,N_4453,N_4455);
and U4506 (N_4506,N_4326,N_4392);
nor U4507 (N_4507,N_4419,N_4408);
nand U4508 (N_4508,N_4266,N_4433);
and U4509 (N_4509,N_4280,N_4413);
nand U4510 (N_4510,N_4386,N_4436);
or U4511 (N_4511,N_4260,N_4349);
and U4512 (N_4512,N_4459,N_4442);
nand U4513 (N_4513,N_4415,N_4288);
nor U4514 (N_4514,N_4430,N_4254);
xnor U4515 (N_4515,N_4259,N_4375);
nand U4516 (N_4516,N_4283,N_4412);
or U4517 (N_4517,N_4370,N_4337);
nand U4518 (N_4518,N_4388,N_4402);
xnor U4519 (N_4519,N_4489,N_4305);
and U4520 (N_4520,N_4467,N_4323);
or U4521 (N_4521,N_4279,N_4286);
and U4522 (N_4522,N_4292,N_4443);
nor U4523 (N_4523,N_4319,N_4368);
or U4524 (N_4524,N_4485,N_4366);
nor U4525 (N_4525,N_4369,N_4397);
and U4526 (N_4526,N_4449,N_4380);
and U4527 (N_4527,N_4480,N_4348);
nand U4528 (N_4528,N_4376,N_4308);
and U4529 (N_4529,N_4252,N_4444);
xnor U4530 (N_4530,N_4322,N_4364);
nand U4531 (N_4531,N_4490,N_4422);
nand U4532 (N_4532,N_4361,N_4373);
and U4533 (N_4533,N_4309,N_4387);
and U4534 (N_4534,N_4466,N_4491);
nor U4535 (N_4535,N_4458,N_4451);
and U4536 (N_4536,N_4318,N_4351);
and U4537 (N_4537,N_4316,N_4333);
and U4538 (N_4538,N_4488,N_4476);
nor U4539 (N_4539,N_4416,N_4423);
or U4540 (N_4540,N_4394,N_4311);
nor U4541 (N_4541,N_4344,N_4383);
or U4542 (N_4542,N_4468,N_4493);
nand U4543 (N_4543,N_4438,N_4251);
and U4544 (N_4544,N_4456,N_4298);
and U4545 (N_4545,N_4331,N_4427);
nor U4546 (N_4546,N_4439,N_4463);
or U4547 (N_4547,N_4477,N_4400);
nor U4548 (N_4548,N_4473,N_4350);
nor U4549 (N_4549,N_4317,N_4482);
and U4550 (N_4550,N_4278,N_4446);
or U4551 (N_4551,N_4372,N_4474);
or U4552 (N_4552,N_4447,N_4478);
xor U4553 (N_4553,N_4374,N_4296);
and U4554 (N_4554,N_4354,N_4399);
and U4555 (N_4555,N_4267,N_4469);
and U4556 (N_4556,N_4441,N_4285);
nand U4557 (N_4557,N_4435,N_4434);
nand U4558 (N_4558,N_4410,N_4464);
nand U4559 (N_4559,N_4404,N_4276);
or U4560 (N_4560,N_4420,N_4271);
and U4561 (N_4561,N_4270,N_4258);
nor U4562 (N_4562,N_4290,N_4452);
xnor U4563 (N_4563,N_4315,N_4256);
and U4564 (N_4564,N_4498,N_4330);
or U4565 (N_4565,N_4407,N_4269);
and U4566 (N_4566,N_4346,N_4450);
and U4567 (N_4567,N_4377,N_4340);
nand U4568 (N_4568,N_4429,N_4409);
or U4569 (N_4569,N_4274,N_4303);
or U4570 (N_4570,N_4324,N_4355);
and U4571 (N_4571,N_4277,N_4462);
nand U4572 (N_4572,N_4424,N_4390);
nand U4573 (N_4573,N_4284,N_4481);
or U4574 (N_4574,N_4275,N_4367);
nand U4575 (N_4575,N_4460,N_4357);
or U4576 (N_4576,N_4250,N_4314);
xnor U4577 (N_4577,N_4263,N_4414);
nor U4578 (N_4578,N_4470,N_4282);
nand U4579 (N_4579,N_4253,N_4360);
and U4580 (N_4580,N_4483,N_4301);
and U4581 (N_4581,N_4353,N_4294);
and U4582 (N_4582,N_4454,N_4381);
or U4583 (N_4583,N_4356,N_4405);
nor U4584 (N_4584,N_4428,N_4461);
nor U4585 (N_4585,N_4479,N_4255);
and U4586 (N_4586,N_4291,N_4440);
and U4587 (N_4587,N_4273,N_4382);
and U4588 (N_4588,N_4261,N_4343);
and U4589 (N_4589,N_4300,N_4425);
nor U4590 (N_4590,N_4445,N_4395);
nor U4591 (N_4591,N_4471,N_4304);
or U4592 (N_4592,N_4406,N_4432);
and U4593 (N_4593,N_4338,N_4342);
or U4594 (N_4594,N_4345,N_4465);
nand U4595 (N_4595,N_4431,N_4293);
xor U4596 (N_4596,N_4495,N_4362);
nor U4597 (N_4597,N_4496,N_4457);
or U4598 (N_4598,N_4389,N_4287);
and U4599 (N_4599,N_4334,N_4295);
nor U4600 (N_4600,N_4299,N_4494);
nand U4601 (N_4601,N_4312,N_4336);
and U4602 (N_4602,N_4329,N_4332);
nand U4603 (N_4603,N_4484,N_4398);
nand U4604 (N_4604,N_4302,N_4307);
xor U4605 (N_4605,N_4257,N_4499);
nor U4606 (N_4606,N_4363,N_4426);
nand U4607 (N_4607,N_4487,N_4448);
nor U4608 (N_4608,N_4281,N_4264);
nand U4609 (N_4609,N_4396,N_4379);
and U4610 (N_4610,N_4475,N_4492);
and U4611 (N_4611,N_4437,N_4335);
and U4612 (N_4612,N_4359,N_4393);
or U4613 (N_4613,N_4497,N_4365);
and U4614 (N_4614,N_4421,N_4262);
nor U4615 (N_4615,N_4378,N_4358);
nand U4616 (N_4616,N_4328,N_4403);
nand U4617 (N_4617,N_4339,N_4265);
and U4618 (N_4618,N_4310,N_4371);
xor U4619 (N_4619,N_4418,N_4341);
and U4620 (N_4620,N_4391,N_4352);
and U4621 (N_4621,N_4321,N_4272);
and U4622 (N_4622,N_4385,N_4384);
nand U4623 (N_4623,N_4347,N_4486);
or U4624 (N_4624,N_4306,N_4417);
and U4625 (N_4625,N_4362,N_4379);
nand U4626 (N_4626,N_4426,N_4491);
and U4627 (N_4627,N_4307,N_4370);
and U4628 (N_4628,N_4371,N_4277);
nand U4629 (N_4629,N_4452,N_4373);
nand U4630 (N_4630,N_4443,N_4338);
and U4631 (N_4631,N_4261,N_4390);
or U4632 (N_4632,N_4438,N_4413);
xnor U4633 (N_4633,N_4272,N_4456);
and U4634 (N_4634,N_4396,N_4410);
xnor U4635 (N_4635,N_4287,N_4330);
nand U4636 (N_4636,N_4487,N_4377);
nor U4637 (N_4637,N_4322,N_4419);
nor U4638 (N_4638,N_4276,N_4452);
xnor U4639 (N_4639,N_4318,N_4389);
nor U4640 (N_4640,N_4473,N_4392);
nand U4641 (N_4641,N_4416,N_4497);
or U4642 (N_4642,N_4374,N_4299);
nor U4643 (N_4643,N_4393,N_4411);
nand U4644 (N_4644,N_4472,N_4385);
or U4645 (N_4645,N_4411,N_4350);
or U4646 (N_4646,N_4350,N_4323);
nor U4647 (N_4647,N_4394,N_4414);
and U4648 (N_4648,N_4410,N_4295);
and U4649 (N_4649,N_4376,N_4383);
and U4650 (N_4650,N_4399,N_4413);
nor U4651 (N_4651,N_4250,N_4288);
and U4652 (N_4652,N_4294,N_4375);
and U4653 (N_4653,N_4258,N_4382);
nand U4654 (N_4654,N_4421,N_4288);
nor U4655 (N_4655,N_4327,N_4356);
or U4656 (N_4656,N_4486,N_4413);
nand U4657 (N_4657,N_4491,N_4394);
or U4658 (N_4658,N_4381,N_4261);
or U4659 (N_4659,N_4269,N_4425);
nor U4660 (N_4660,N_4481,N_4480);
nor U4661 (N_4661,N_4353,N_4270);
and U4662 (N_4662,N_4388,N_4430);
nor U4663 (N_4663,N_4256,N_4278);
nand U4664 (N_4664,N_4496,N_4389);
nor U4665 (N_4665,N_4282,N_4452);
nand U4666 (N_4666,N_4371,N_4325);
xnor U4667 (N_4667,N_4441,N_4433);
or U4668 (N_4668,N_4455,N_4355);
or U4669 (N_4669,N_4377,N_4492);
nor U4670 (N_4670,N_4365,N_4308);
nand U4671 (N_4671,N_4363,N_4293);
nand U4672 (N_4672,N_4331,N_4481);
xnor U4673 (N_4673,N_4331,N_4333);
and U4674 (N_4674,N_4289,N_4450);
nand U4675 (N_4675,N_4476,N_4385);
xnor U4676 (N_4676,N_4461,N_4437);
nand U4677 (N_4677,N_4491,N_4344);
or U4678 (N_4678,N_4298,N_4398);
or U4679 (N_4679,N_4397,N_4344);
nor U4680 (N_4680,N_4488,N_4409);
and U4681 (N_4681,N_4285,N_4472);
or U4682 (N_4682,N_4350,N_4424);
nor U4683 (N_4683,N_4494,N_4278);
and U4684 (N_4684,N_4399,N_4297);
nand U4685 (N_4685,N_4380,N_4484);
nand U4686 (N_4686,N_4421,N_4468);
and U4687 (N_4687,N_4323,N_4304);
or U4688 (N_4688,N_4355,N_4432);
or U4689 (N_4689,N_4417,N_4250);
and U4690 (N_4690,N_4368,N_4452);
or U4691 (N_4691,N_4430,N_4296);
nor U4692 (N_4692,N_4317,N_4445);
nand U4693 (N_4693,N_4490,N_4328);
nor U4694 (N_4694,N_4373,N_4385);
nand U4695 (N_4695,N_4296,N_4396);
nand U4696 (N_4696,N_4328,N_4260);
xor U4697 (N_4697,N_4358,N_4496);
or U4698 (N_4698,N_4488,N_4433);
nor U4699 (N_4699,N_4392,N_4499);
or U4700 (N_4700,N_4300,N_4490);
or U4701 (N_4701,N_4348,N_4264);
or U4702 (N_4702,N_4341,N_4306);
or U4703 (N_4703,N_4437,N_4455);
nand U4704 (N_4704,N_4289,N_4461);
nor U4705 (N_4705,N_4273,N_4438);
xor U4706 (N_4706,N_4336,N_4254);
and U4707 (N_4707,N_4274,N_4282);
nor U4708 (N_4708,N_4419,N_4387);
or U4709 (N_4709,N_4293,N_4447);
nand U4710 (N_4710,N_4406,N_4286);
nor U4711 (N_4711,N_4289,N_4340);
xnor U4712 (N_4712,N_4263,N_4311);
and U4713 (N_4713,N_4271,N_4406);
xor U4714 (N_4714,N_4481,N_4291);
or U4715 (N_4715,N_4282,N_4297);
and U4716 (N_4716,N_4340,N_4451);
nor U4717 (N_4717,N_4415,N_4398);
nand U4718 (N_4718,N_4474,N_4295);
nand U4719 (N_4719,N_4367,N_4454);
or U4720 (N_4720,N_4250,N_4276);
or U4721 (N_4721,N_4293,N_4446);
xnor U4722 (N_4722,N_4276,N_4410);
or U4723 (N_4723,N_4296,N_4429);
nand U4724 (N_4724,N_4385,N_4449);
nand U4725 (N_4725,N_4451,N_4252);
or U4726 (N_4726,N_4366,N_4313);
and U4727 (N_4727,N_4428,N_4347);
nand U4728 (N_4728,N_4495,N_4357);
and U4729 (N_4729,N_4477,N_4371);
xnor U4730 (N_4730,N_4356,N_4353);
nor U4731 (N_4731,N_4483,N_4439);
nand U4732 (N_4732,N_4319,N_4335);
nand U4733 (N_4733,N_4482,N_4387);
and U4734 (N_4734,N_4438,N_4324);
nor U4735 (N_4735,N_4347,N_4296);
and U4736 (N_4736,N_4478,N_4437);
xnor U4737 (N_4737,N_4330,N_4465);
and U4738 (N_4738,N_4380,N_4389);
or U4739 (N_4739,N_4254,N_4424);
nor U4740 (N_4740,N_4273,N_4387);
xnor U4741 (N_4741,N_4272,N_4396);
nand U4742 (N_4742,N_4442,N_4307);
nor U4743 (N_4743,N_4486,N_4432);
nor U4744 (N_4744,N_4262,N_4342);
nand U4745 (N_4745,N_4324,N_4368);
nand U4746 (N_4746,N_4302,N_4303);
xor U4747 (N_4747,N_4314,N_4454);
xor U4748 (N_4748,N_4310,N_4291);
and U4749 (N_4749,N_4447,N_4357);
or U4750 (N_4750,N_4536,N_4647);
nor U4751 (N_4751,N_4643,N_4532);
or U4752 (N_4752,N_4605,N_4733);
or U4753 (N_4753,N_4575,N_4744);
or U4754 (N_4754,N_4644,N_4514);
nand U4755 (N_4755,N_4691,N_4638);
nand U4756 (N_4756,N_4746,N_4646);
nand U4757 (N_4757,N_4660,N_4731);
and U4758 (N_4758,N_4739,N_4736);
nand U4759 (N_4759,N_4601,N_4729);
or U4760 (N_4760,N_4672,N_4524);
and U4761 (N_4761,N_4577,N_4580);
nand U4762 (N_4762,N_4694,N_4718);
xor U4763 (N_4763,N_4604,N_4742);
and U4764 (N_4764,N_4700,N_4712);
nor U4765 (N_4765,N_4545,N_4500);
or U4766 (N_4766,N_4669,N_4619);
xor U4767 (N_4767,N_4664,N_4683);
nand U4768 (N_4768,N_4728,N_4556);
xnor U4769 (N_4769,N_4618,N_4745);
and U4770 (N_4770,N_4584,N_4651);
nor U4771 (N_4771,N_4547,N_4502);
nor U4772 (N_4772,N_4696,N_4697);
xnor U4773 (N_4773,N_4741,N_4549);
and U4774 (N_4774,N_4613,N_4709);
or U4775 (N_4775,N_4639,N_4698);
nor U4776 (N_4776,N_4705,N_4678);
nand U4777 (N_4777,N_4544,N_4603);
and U4778 (N_4778,N_4714,N_4525);
or U4779 (N_4779,N_4515,N_4535);
and U4780 (N_4780,N_4607,N_4609);
xnor U4781 (N_4781,N_4555,N_4567);
or U4782 (N_4782,N_4543,N_4716);
xnor U4783 (N_4783,N_4597,N_4551);
nor U4784 (N_4784,N_4677,N_4627);
or U4785 (N_4785,N_4570,N_4637);
nand U4786 (N_4786,N_4686,N_4610);
or U4787 (N_4787,N_4624,N_4702);
and U4788 (N_4788,N_4723,N_4732);
or U4789 (N_4789,N_4519,N_4717);
or U4790 (N_4790,N_4511,N_4722);
xor U4791 (N_4791,N_4558,N_4522);
and U4792 (N_4792,N_4665,N_4565);
nand U4793 (N_4793,N_4501,N_4743);
and U4794 (N_4794,N_4541,N_4670);
nor U4795 (N_4795,N_4526,N_4740);
or U4796 (N_4796,N_4685,N_4513);
or U4797 (N_4797,N_4621,N_4676);
nand U4798 (N_4798,N_4578,N_4630);
nand U4799 (N_4799,N_4560,N_4715);
or U4800 (N_4800,N_4747,N_4661);
nand U4801 (N_4801,N_4719,N_4616);
nand U4802 (N_4802,N_4680,N_4690);
and U4803 (N_4803,N_4615,N_4591);
nor U4804 (N_4804,N_4645,N_4582);
and U4805 (N_4805,N_4562,N_4521);
xnor U4806 (N_4806,N_4659,N_4509);
nor U4807 (N_4807,N_4730,N_4632);
nand U4808 (N_4808,N_4503,N_4512);
xor U4809 (N_4809,N_4623,N_4537);
or U4810 (N_4810,N_4612,N_4552);
and U4811 (N_4811,N_4738,N_4517);
or U4812 (N_4812,N_4735,N_4564);
or U4813 (N_4813,N_4546,N_4505);
nand U4814 (N_4814,N_4640,N_4726);
nand U4815 (N_4815,N_4542,N_4557);
and U4816 (N_4816,N_4574,N_4581);
nor U4817 (N_4817,N_4529,N_4625);
or U4818 (N_4818,N_4682,N_4679);
nand U4819 (N_4819,N_4510,N_4688);
xnor U4820 (N_4820,N_4720,N_4527);
nor U4821 (N_4821,N_4657,N_4654);
or U4822 (N_4822,N_4550,N_4649);
and U4823 (N_4823,N_4662,N_4569);
nor U4824 (N_4824,N_4590,N_4588);
nand U4825 (N_4825,N_4563,N_4622);
nor U4826 (N_4826,N_4703,N_4693);
nor U4827 (N_4827,N_4599,N_4583);
and U4828 (N_4828,N_4626,N_4533);
nand U4829 (N_4829,N_4506,N_4658);
nand U4830 (N_4830,N_4592,N_4674);
nand U4831 (N_4831,N_4595,N_4633);
or U4832 (N_4832,N_4508,N_4518);
and U4833 (N_4833,N_4681,N_4713);
nor U4834 (N_4834,N_4531,N_4606);
nand U4835 (N_4835,N_4673,N_4579);
xor U4836 (N_4836,N_4585,N_4699);
or U4837 (N_4837,N_4641,N_4652);
xnor U4838 (N_4838,N_4684,N_4568);
nor U4839 (N_4839,N_4655,N_4523);
or U4840 (N_4840,N_4663,N_4587);
or U4841 (N_4841,N_4553,N_4516);
or U4842 (N_4842,N_4721,N_4701);
or U4843 (N_4843,N_4636,N_4614);
nor U4844 (N_4844,N_4704,N_4648);
nor U4845 (N_4845,N_4561,N_4600);
nand U4846 (N_4846,N_4737,N_4617);
nand U4847 (N_4847,N_4692,N_4594);
or U4848 (N_4848,N_4724,N_4593);
nor U4849 (N_4849,N_4530,N_4586);
nor U4850 (N_4850,N_4540,N_4749);
or U4851 (N_4851,N_4711,N_4573);
nand U4852 (N_4852,N_4554,N_4653);
nand U4853 (N_4853,N_4608,N_4635);
nor U4854 (N_4854,N_4589,N_4707);
nor U4855 (N_4855,N_4710,N_4725);
nand U4856 (N_4856,N_4734,N_4566);
xor U4857 (N_4857,N_4727,N_4695);
nor U4858 (N_4858,N_4656,N_4611);
and U4859 (N_4859,N_4534,N_4666);
or U4860 (N_4860,N_4528,N_4687);
or U4861 (N_4861,N_4668,N_4559);
nor U4862 (N_4862,N_4708,N_4507);
nor U4863 (N_4863,N_4548,N_4596);
and U4864 (N_4864,N_4572,N_4539);
or U4865 (N_4865,N_4689,N_4667);
nor U4866 (N_4866,N_4671,N_4650);
nor U4867 (N_4867,N_4628,N_4602);
or U4868 (N_4868,N_4748,N_4571);
or U4869 (N_4869,N_4598,N_4576);
or U4870 (N_4870,N_4504,N_4706);
or U4871 (N_4871,N_4538,N_4629);
xor U4872 (N_4872,N_4631,N_4675);
nor U4873 (N_4873,N_4634,N_4620);
nor U4874 (N_4874,N_4642,N_4520);
or U4875 (N_4875,N_4645,N_4590);
or U4876 (N_4876,N_4730,N_4567);
or U4877 (N_4877,N_4534,N_4721);
nand U4878 (N_4878,N_4704,N_4666);
and U4879 (N_4879,N_4690,N_4604);
nor U4880 (N_4880,N_4524,N_4518);
or U4881 (N_4881,N_4744,N_4650);
xnor U4882 (N_4882,N_4536,N_4664);
nand U4883 (N_4883,N_4524,N_4720);
nand U4884 (N_4884,N_4570,N_4529);
nor U4885 (N_4885,N_4734,N_4642);
or U4886 (N_4886,N_4722,N_4705);
or U4887 (N_4887,N_4703,N_4577);
nor U4888 (N_4888,N_4653,N_4730);
or U4889 (N_4889,N_4707,N_4507);
nor U4890 (N_4890,N_4673,N_4663);
or U4891 (N_4891,N_4651,N_4745);
nand U4892 (N_4892,N_4519,N_4619);
nor U4893 (N_4893,N_4670,N_4569);
and U4894 (N_4894,N_4629,N_4611);
nor U4895 (N_4895,N_4564,N_4536);
nor U4896 (N_4896,N_4553,N_4526);
nand U4897 (N_4897,N_4529,N_4658);
or U4898 (N_4898,N_4716,N_4718);
nor U4899 (N_4899,N_4717,N_4558);
and U4900 (N_4900,N_4720,N_4702);
xnor U4901 (N_4901,N_4508,N_4699);
or U4902 (N_4902,N_4588,N_4609);
nor U4903 (N_4903,N_4520,N_4593);
xnor U4904 (N_4904,N_4628,N_4708);
or U4905 (N_4905,N_4536,N_4679);
xor U4906 (N_4906,N_4670,N_4504);
nor U4907 (N_4907,N_4520,N_4568);
xor U4908 (N_4908,N_4734,N_4698);
or U4909 (N_4909,N_4587,N_4644);
or U4910 (N_4910,N_4572,N_4528);
or U4911 (N_4911,N_4680,N_4581);
nor U4912 (N_4912,N_4547,N_4725);
nor U4913 (N_4913,N_4544,N_4649);
nor U4914 (N_4914,N_4690,N_4515);
nor U4915 (N_4915,N_4572,N_4716);
or U4916 (N_4916,N_4519,N_4573);
nand U4917 (N_4917,N_4518,N_4701);
nor U4918 (N_4918,N_4577,N_4565);
or U4919 (N_4919,N_4604,N_4663);
nand U4920 (N_4920,N_4568,N_4627);
nand U4921 (N_4921,N_4563,N_4738);
nand U4922 (N_4922,N_4656,N_4556);
nand U4923 (N_4923,N_4520,N_4727);
nor U4924 (N_4924,N_4513,N_4558);
nand U4925 (N_4925,N_4557,N_4638);
or U4926 (N_4926,N_4656,N_4500);
or U4927 (N_4927,N_4573,N_4551);
nor U4928 (N_4928,N_4581,N_4561);
or U4929 (N_4929,N_4586,N_4735);
xnor U4930 (N_4930,N_4615,N_4734);
or U4931 (N_4931,N_4709,N_4532);
nand U4932 (N_4932,N_4649,N_4611);
xnor U4933 (N_4933,N_4702,N_4632);
or U4934 (N_4934,N_4671,N_4699);
nor U4935 (N_4935,N_4732,N_4667);
nor U4936 (N_4936,N_4726,N_4540);
and U4937 (N_4937,N_4585,N_4550);
nand U4938 (N_4938,N_4703,N_4664);
and U4939 (N_4939,N_4530,N_4588);
or U4940 (N_4940,N_4545,N_4526);
nor U4941 (N_4941,N_4527,N_4718);
and U4942 (N_4942,N_4523,N_4536);
or U4943 (N_4943,N_4632,N_4672);
and U4944 (N_4944,N_4585,N_4734);
and U4945 (N_4945,N_4537,N_4584);
or U4946 (N_4946,N_4603,N_4604);
and U4947 (N_4947,N_4554,N_4552);
and U4948 (N_4948,N_4598,N_4532);
and U4949 (N_4949,N_4674,N_4680);
nor U4950 (N_4950,N_4726,N_4704);
nor U4951 (N_4951,N_4660,N_4608);
or U4952 (N_4952,N_4610,N_4722);
and U4953 (N_4953,N_4527,N_4635);
or U4954 (N_4954,N_4528,N_4701);
or U4955 (N_4955,N_4673,N_4624);
nand U4956 (N_4956,N_4618,N_4740);
nor U4957 (N_4957,N_4571,N_4663);
or U4958 (N_4958,N_4601,N_4739);
nand U4959 (N_4959,N_4738,N_4588);
nor U4960 (N_4960,N_4625,N_4606);
and U4961 (N_4961,N_4535,N_4617);
xor U4962 (N_4962,N_4637,N_4533);
nand U4963 (N_4963,N_4513,N_4630);
and U4964 (N_4964,N_4617,N_4571);
xor U4965 (N_4965,N_4605,N_4731);
and U4966 (N_4966,N_4550,N_4701);
and U4967 (N_4967,N_4737,N_4530);
or U4968 (N_4968,N_4747,N_4745);
and U4969 (N_4969,N_4661,N_4741);
or U4970 (N_4970,N_4527,N_4525);
nand U4971 (N_4971,N_4559,N_4516);
nor U4972 (N_4972,N_4532,N_4686);
and U4973 (N_4973,N_4506,N_4712);
or U4974 (N_4974,N_4681,N_4632);
nand U4975 (N_4975,N_4628,N_4729);
nor U4976 (N_4976,N_4505,N_4514);
or U4977 (N_4977,N_4658,N_4711);
xor U4978 (N_4978,N_4680,N_4676);
nor U4979 (N_4979,N_4543,N_4544);
or U4980 (N_4980,N_4580,N_4697);
or U4981 (N_4981,N_4539,N_4621);
nor U4982 (N_4982,N_4676,N_4702);
or U4983 (N_4983,N_4660,N_4585);
nor U4984 (N_4984,N_4626,N_4686);
or U4985 (N_4985,N_4577,N_4702);
or U4986 (N_4986,N_4504,N_4562);
nand U4987 (N_4987,N_4624,N_4734);
or U4988 (N_4988,N_4597,N_4582);
and U4989 (N_4989,N_4744,N_4631);
nand U4990 (N_4990,N_4682,N_4521);
nand U4991 (N_4991,N_4635,N_4705);
and U4992 (N_4992,N_4641,N_4587);
nand U4993 (N_4993,N_4632,N_4566);
nand U4994 (N_4994,N_4574,N_4634);
xnor U4995 (N_4995,N_4702,N_4674);
nor U4996 (N_4996,N_4564,N_4545);
and U4997 (N_4997,N_4573,N_4609);
nand U4998 (N_4998,N_4620,N_4682);
nand U4999 (N_4999,N_4713,N_4706);
nand U5000 (N_5000,N_4965,N_4894);
and U5001 (N_5001,N_4860,N_4834);
nand U5002 (N_5002,N_4836,N_4843);
nand U5003 (N_5003,N_4776,N_4941);
nor U5004 (N_5004,N_4900,N_4920);
and U5005 (N_5005,N_4958,N_4835);
nand U5006 (N_5006,N_4767,N_4787);
nor U5007 (N_5007,N_4858,N_4824);
or U5008 (N_5008,N_4773,N_4810);
and U5009 (N_5009,N_4873,N_4970);
or U5010 (N_5010,N_4959,N_4888);
nor U5011 (N_5011,N_4973,N_4798);
nor U5012 (N_5012,N_4809,N_4936);
and U5013 (N_5013,N_4874,N_4785);
or U5014 (N_5014,N_4772,N_4995);
or U5015 (N_5015,N_4831,N_4988);
and U5016 (N_5016,N_4823,N_4901);
and U5017 (N_5017,N_4851,N_4914);
and U5018 (N_5018,N_4840,N_4909);
nand U5019 (N_5019,N_4879,N_4911);
xor U5020 (N_5020,N_4897,N_4999);
nor U5021 (N_5021,N_4937,N_4980);
or U5022 (N_5022,N_4946,N_4786);
nand U5023 (N_5023,N_4863,N_4754);
nor U5024 (N_5024,N_4753,N_4885);
nand U5025 (N_5025,N_4949,N_4800);
nor U5026 (N_5026,N_4871,N_4876);
nand U5027 (N_5027,N_4804,N_4902);
nand U5028 (N_5028,N_4927,N_4945);
xnor U5029 (N_5029,N_4884,N_4757);
and U5030 (N_5030,N_4816,N_4813);
nor U5031 (N_5031,N_4947,N_4991);
and U5032 (N_5032,N_4916,N_4774);
and U5033 (N_5033,N_4982,N_4951);
and U5034 (N_5034,N_4953,N_4822);
nand U5035 (N_5035,N_4756,N_4933);
or U5036 (N_5036,N_4960,N_4938);
nand U5037 (N_5037,N_4790,N_4985);
nand U5038 (N_5038,N_4839,N_4907);
xnor U5039 (N_5039,N_4864,N_4921);
or U5040 (N_5040,N_4766,N_4848);
nand U5041 (N_5041,N_4811,N_4977);
and U5042 (N_5042,N_4849,N_4950);
and U5043 (N_5043,N_4775,N_4913);
xnor U5044 (N_5044,N_4881,N_4964);
nand U5045 (N_5045,N_4818,N_4758);
nand U5046 (N_5046,N_4918,N_4802);
or U5047 (N_5047,N_4861,N_4768);
xnor U5048 (N_5048,N_4877,N_4752);
or U5049 (N_5049,N_4865,N_4948);
nor U5050 (N_5050,N_4987,N_4764);
and U5051 (N_5051,N_4783,N_4975);
nand U5052 (N_5052,N_4917,N_4808);
nor U5053 (N_5053,N_4968,N_4910);
nand U5054 (N_5054,N_4967,N_4765);
nand U5055 (N_5055,N_4944,N_4782);
or U5056 (N_5056,N_4979,N_4912);
or U5057 (N_5057,N_4788,N_4781);
and U5058 (N_5058,N_4795,N_4929);
nand U5059 (N_5059,N_4963,N_4961);
nor U5060 (N_5060,N_4779,N_4807);
xor U5061 (N_5061,N_4784,N_4998);
or U5062 (N_5062,N_4990,N_4895);
and U5063 (N_5063,N_4854,N_4996);
or U5064 (N_5064,N_4883,N_4924);
and U5065 (N_5065,N_4815,N_4896);
nand U5066 (N_5066,N_4828,N_4966);
nor U5067 (N_5067,N_4750,N_4806);
nor U5068 (N_5068,N_4978,N_4797);
and U5069 (N_5069,N_4972,N_4763);
nor U5070 (N_5070,N_4777,N_4870);
nand U5071 (N_5071,N_4821,N_4827);
nand U5072 (N_5072,N_4867,N_4856);
nor U5073 (N_5073,N_4889,N_4762);
xnor U5074 (N_5074,N_4904,N_4915);
or U5075 (N_5075,N_4971,N_4832);
and U5076 (N_5076,N_4847,N_4923);
nand U5077 (N_5077,N_4983,N_4794);
xor U5078 (N_5078,N_4799,N_4986);
nor U5079 (N_5079,N_4844,N_4761);
and U5080 (N_5080,N_4837,N_4976);
nand U5081 (N_5081,N_4857,N_4819);
and U5082 (N_5082,N_4791,N_4957);
nand U5083 (N_5083,N_4887,N_4866);
nor U5084 (N_5084,N_4993,N_4825);
xnor U5085 (N_5085,N_4939,N_4789);
nor U5086 (N_5086,N_4931,N_4855);
and U5087 (N_5087,N_4922,N_4869);
nor U5088 (N_5088,N_4755,N_4955);
or U5089 (N_5089,N_4751,N_4845);
or U5090 (N_5090,N_4796,N_4899);
and U5091 (N_5091,N_4935,N_4956);
and U5092 (N_5092,N_4829,N_4940);
and U5093 (N_5093,N_4760,N_4997);
and U5094 (N_5094,N_4981,N_4830);
nor U5095 (N_5095,N_4759,N_4872);
or U5096 (N_5096,N_4994,N_4771);
xor U5097 (N_5097,N_4992,N_4850);
and U5098 (N_5098,N_4838,N_4928);
and U5099 (N_5099,N_4880,N_4793);
nor U5100 (N_5100,N_4934,N_4833);
or U5101 (N_5101,N_4892,N_4846);
nor U5102 (N_5102,N_4984,N_4778);
or U5103 (N_5103,N_4769,N_4925);
and U5104 (N_5104,N_4969,N_4954);
or U5105 (N_5105,N_4841,N_4820);
nor U5106 (N_5106,N_4908,N_4962);
or U5107 (N_5107,N_4878,N_4801);
xnor U5108 (N_5108,N_4906,N_4803);
or U5109 (N_5109,N_4882,N_4862);
nor U5110 (N_5110,N_4805,N_4817);
or U5111 (N_5111,N_4792,N_4859);
nor U5112 (N_5112,N_4905,N_4974);
or U5113 (N_5113,N_4890,N_4932);
and U5114 (N_5114,N_4891,N_4886);
or U5115 (N_5115,N_4770,N_4930);
nor U5116 (N_5116,N_4852,N_4989);
or U5117 (N_5117,N_4898,N_4812);
nor U5118 (N_5118,N_4842,N_4826);
and U5119 (N_5119,N_4926,N_4893);
nand U5120 (N_5120,N_4942,N_4952);
and U5121 (N_5121,N_4853,N_4919);
nor U5122 (N_5122,N_4903,N_4814);
xor U5123 (N_5123,N_4875,N_4780);
nand U5124 (N_5124,N_4868,N_4943);
and U5125 (N_5125,N_4974,N_4936);
nor U5126 (N_5126,N_4940,N_4930);
xor U5127 (N_5127,N_4767,N_4798);
nand U5128 (N_5128,N_4857,N_4759);
or U5129 (N_5129,N_4769,N_4980);
or U5130 (N_5130,N_4803,N_4804);
nor U5131 (N_5131,N_4883,N_4985);
nor U5132 (N_5132,N_4865,N_4888);
nand U5133 (N_5133,N_4875,N_4784);
nor U5134 (N_5134,N_4814,N_4762);
nand U5135 (N_5135,N_4838,N_4786);
and U5136 (N_5136,N_4799,N_4908);
xor U5137 (N_5137,N_4831,N_4887);
and U5138 (N_5138,N_4902,N_4865);
nor U5139 (N_5139,N_4941,N_4785);
nor U5140 (N_5140,N_4823,N_4965);
or U5141 (N_5141,N_4825,N_4835);
or U5142 (N_5142,N_4768,N_4752);
or U5143 (N_5143,N_4967,N_4847);
or U5144 (N_5144,N_4863,N_4883);
or U5145 (N_5145,N_4903,N_4911);
and U5146 (N_5146,N_4809,N_4967);
and U5147 (N_5147,N_4757,N_4786);
nand U5148 (N_5148,N_4801,N_4818);
or U5149 (N_5149,N_4889,N_4909);
nand U5150 (N_5150,N_4848,N_4852);
nor U5151 (N_5151,N_4989,N_4883);
nand U5152 (N_5152,N_4974,N_4810);
nor U5153 (N_5153,N_4967,N_4878);
or U5154 (N_5154,N_4851,N_4901);
or U5155 (N_5155,N_4767,N_4950);
nand U5156 (N_5156,N_4827,N_4947);
or U5157 (N_5157,N_4942,N_4779);
or U5158 (N_5158,N_4993,N_4896);
or U5159 (N_5159,N_4814,N_4999);
xnor U5160 (N_5160,N_4993,N_4981);
or U5161 (N_5161,N_4775,N_4974);
nand U5162 (N_5162,N_4882,N_4873);
nor U5163 (N_5163,N_4798,N_4871);
nand U5164 (N_5164,N_4800,N_4974);
nand U5165 (N_5165,N_4951,N_4841);
nor U5166 (N_5166,N_4988,N_4955);
and U5167 (N_5167,N_4784,N_4847);
nor U5168 (N_5168,N_4951,N_4825);
nand U5169 (N_5169,N_4877,N_4833);
nor U5170 (N_5170,N_4995,N_4947);
nor U5171 (N_5171,N_4955,N_4924);
or U5172 (N_5172,N_4867,N_4978);
or U5173 (N_5173,N_4869,N_4769);
and U5174 (N_5174,N_4904,N_4812);
nor U5175 (N_5175,N_4915,N_4861);
or U5176 (N_5176,N_4996,N_4813);
nor U5177 (N_5177,N_4846,N_4962);
nand U5178 (N_5178,N_4773,N_4824);
nand U5179 (N_5179,N_4955,N_4826);
and U5180 (N_5180,N_4797,N_4889);
nor U5181 (N_5181,N_4918,N_4917);
nor U5182 (N_5182,N_4808,N_4752);
or U5183 (N_5183,N_4792,N_4816);
nand U5184 (N_5184,N_4986,N_4823);
xnor U5185 (N_5185,N_4783,N_4821);
and U5186 (N_5186,N_4759,N_4922);
nand U5187 (N_5187,N_4840,N_4865);
nand U5188 (N_5188,N_4753,N_4754);
and U5189 (N_5189,N_4796,N_4841);
and U5190 (N_5190,N_4826,N_4789);
nor U5191 (N_5191,N_4936,N_4999);
and U5192 (N_5192,N_4890,N_4943);
nand U5193 (N_5193,N_4759,N_4771);
nor U5194 (N_5194,N_4852,N_4863);
xor U5195 (N_5195,N_4827,N_4857);
nand U5196 (N_5196,N_4871,N_4785);
or U5197 (N_5197,N_4978,N_4930);
xor U5198 (N_5198,N_4943,N_4858);
or U5199 (N_5199,N_4882,N_4779);
nand U5200 (N_5200,N_4823,N_4961);
nand U5201 (N_5201,N_4769,N_4758);
or U5202 (N_5202,N_4851,N_4869);
nor U5203 (N_5203,N_4808,N_4983);
and U5204 (N_5204,N_4800,N_4905);
and U5205 (N_5205,N_4981,N_4778);
nand U5206 (N_5206,N_4929,N_4893);
nand U5207 (N_5207,N_4999,N_4948);
nand U5208 (N_5208,N_4947,N_4842);
xnor U5209 (N_5209,N_4923,N_4905);
or U5210 (N_5210,N_4997,N_4866);
or U5211 (N_5211,N_4917,N_4984);
or U5212 (N_5212,N_4792,N_4794);
xor U5213 (N_5213,N_4815,N_4760);
xor U5214 (N_5214,N_4908,N_4818);
nor U5215 (N_5215,N_4890,N_4946);
xor U5216 (N_5216,N_4844,N_4752);
or U5217 (N_5217,N_4961,N_4764);
xnor U5218 (N_5218,N_4926,N_4896);
or U5219 (N_5219,N_4973,N_4990);
nor U5220 (N_5220,N_4926,N_4783);
or U5221 (N_5221,N_4900,N_4757);
nand U5222 (N_5222,N_4877,N_4881);
nor U5223 (N_5223,N_4914,N_4837);
and U5224 (N_5224,N_4841,N_4794);
and U5225 (N_5225,N_4806,N_4874);
and U5226 (N_5226,N_4751,N_4993);
xnor U5227 (N_5227,N_4825,N_4774);
and U5228 (N_5228,N_4844,N_4814);
or U5229 (N_5229,N_4753,N_4887);
or U5230 (N_5230,N_4780,N_4808);
and U5231 (N_5231,N_4846,N_4958);
nor U5232 (N_5232,N_4899,N_4997);
or U5233 (N_5233,N_4905,N_4912);
xnor U5234 (N_5234,N_4956,N_4851);
or U5235 (N_5235,N_4941,N_4822);
or U5236 (N_5236,N_4927,N_4797);
nor U5237 (N_5237,N_4767,N_4768);
or U5238 (N_5238,N_4973,N_4960);
and U5239 (N_5239,N_4801,N_4832);
xnor U5240 (N_5240,N_4836,N_4854);
nand U5241 (N_5241,N_4817,N_4852);
nor U5242 (N_5242,N_4824,N_4867);
and U5243 (N_5243,N_4757,N_4925);
and U5244 (N_5244,N_4796,N_4833);
nand U5245 (N_5245,N_4858,N_4841);
nor U5246 (N_5246,N_4751,N_4933);
nor U5247 (N_5247,N_4812,N_4852);
and U5248 (N_5248,N_4974,N_4812);
xnor U5249 (N_5249,N_4957,N_4880);
nor U5250 (N_5250,N_5007,N_5188);
nand U5251 (N_5251,N_5184,N_5003);
and U5252 (N_5252,N_5209,N_5066);
nand U5253 (N_5253,N_5070,N_5226);
and U5254 (N_5254,N_5020,N_5141);
xor U5255 (N_5255,N_5138,N_5163);
and U5256 (N_5256,N_5216,N_5104);
and U5257 (N_5257,N_5147,N_5248);
nor U5258 (N_5258,N_5123,N_5035);
nand U5259 (N_5259,N_5233,N_5051);
or U5260 (N_5260,N_5156,N_5182);
nand U5261 (N_5261,N_5203,N_5229);
nand U5262 (N_5262,N_5239,N_5024);
and U5263 (N_5263,N_5162,N_5149);
and U5264 (N_5264,N_5198,N_5140);
nor U5265 (N_5265,N_5037,N_5013);
nand U5266 (N_5266,N_5048,N_5175);
xnor U5267 (N_5267,N_5222,N_5113);
nor U5268 (N_5268,N_5179,N_5171);
and U5269 (N_5269,N_5073,N_5200);
and U5270 (N_5270,N_5206,N_5208);
and U5271 (N_5271,N_5089,N_5095);
and U5272 (N_5272,N_5106,N_5069);
or U5273 (N_5273,N_5168,N_5165);
or U5274 (N_5274,N_5065,N_5122);
nand U5275 (N_5275,N_5011,N_5078);
and U5276 (N_5276,N_5129,N_5185);
or U5277 (N_5277,N_5195,N_5067);
nand U5278 (N_5278,N_5231,N_5211);
nor U5279 (N_5279,N_5097,N_5120);
and U5280 (N_5280,N_5001,N_5083);
xnor U5281 (N_5281,N_5170,N_5006);
and U5282 (N_5282,N_5016,N_5192);
nor U5283 (N_5283,N_5029,N_5088);
and U5284 (N_5284,N_5143,N_5155);
or U5285 (N_5285,N_5101,N_5081);
nand U5286 (N_5286,N_5099,N_5042);
nor U5287 (N_5287,N_5121,N_5153);
or U5288 (N_5288,N_5093,N_5151);
nand U5289 (N_5289,N_5117,N_5018);
nor U5290 (N_5290,N_5112,N_5119);
or U5291 (N_5291,N_5193,N_5232);
nand U5292 (N_5292,N_5082,N_5098);
nand U5293 (N_5293,N_5044,N_5017);
and U5294 (N_5294,N_5105,N_5139);
nand U5295 (N_5295,N_5154,N_5027);
and U5296 (N_5296,N_5110,N_5009);
xnor U5297 (N_5297,N_5130,N_5199);
and U5298 (N_5298,N_5235,N_5166);
and U5299 (N_5299,N_5036,N_5126);
nor U5300 (N_5300,N_5012,N_5102);
and U5301 (N_5301,N_5189,N_5196);
nand U5302 (N_5302,N_5047,N_5063);
or U5303 (N_5303,N_5059,N_5079);
nor U5304 (N_5304,N_5023,N_5055);
or U5305 (N_5305,N_5215,N_5234);
xnor U5306 (N_5306,N_5076,N_5114);
or U5307 (N_5307,N_5243,N_5228);
nand U5308 (N_5308,N_5207,N_5186);
and U5309 (N_5309,N_5021,N_5237);
nand U5310 (N_5310,N_5157,N_5049);
nor U5311 (N_5311,N_5190,N_5212);
and U5312 (N_5312,N_5194,N_5052);
or U5313 (N_5313,N_5014,N_5085);
and U5314 (N_5314,N_5077,N_5022);
nand U5315 (N_5315,N_5075,N_5000);
and U5316 (N_5316,N_5238,N_5202);
nand U5317 (N_5317,N_5204,N_5004);
xor U5318 (N_5318,N_5136,N_5015);
nand U5319 (N_5319,N_5096,N_5100);
or U5320 (N_5320,N_5030,N_5010);
nor U5321 (N_5321,N_5084,N_5033);
nand U5322 (N_5322,N_5227,N_5174);
nand U5323 (N_5323,N_5127,N_5146);
nand U5324 (N_5324,N_5094,N_5178);
or U5325 (N_5325,N_5148,N_5158);
nor U5326 (N_5326,N_5080,N_5164);
nor U5327 (N_5327,N_5177,N_5150);
nor U5328 (N_5328,N_5135,N_5002);
nor U5329 (N_5329,N_5054,N_5005);
or U5330 (N_5330,N_5041,N_5214);
and U5331 (N_5331,N_5172,N_5245);
nor U5332 (N_5332,N_5092,N_5244);
nand U5333 (N_5333,N_5111,N_5125);
and U5334 (N_5334,N_5205,N_5038);
nand U5335 (N_5335,N_5220,N_5133);
nor U5336 (N_5336,N_5240,N_5062);
nand U5337 (N_5337,N_5103,N_5134);
nor U5338 (N_5338,N_5025,N_5064);
nand U5339 (N_5339,N_5223,N_5068);
nand U5340 (N_5340,N_5181,N_5180);
and U5341 (N_5341,N_5145,N_5210);
or U5342 (N_5342,N_5169,N_5053);
or U5343 (N_5343,N_5201,N_5241);
xor U5344 (N_5344,N_5167,N_5058);
and U5345 (N_5345,N_5225,N_5219);
nand U5346 (N_5346,N_5008,N_5173);
and U5347 (N_5347,N_5221,N_5213);
nor U5348 (N_5348,N_5247,N_5217);
xor U5349 (N_5349,N_5249,N_5090);
and U5350 (N_5350,N_5224,N_5132);
and U5351 (N_5351,N_5124,N_5031);
nand U5352 (N_5352,N_5074,N_5091);
nor U5353 (N_5353,N_5032,N_5028);
and U5354 (N_5354,N_5236,N_5131);
and U5355 (N_5355,N_5183,N_5109);
and U5356 (N_5356,N_5230,N_5108);
nor U5357 (N_5357,N_5039,N_5218);
nor U5358 (N_5358,N_5128,N_5242);
nand U5359 (N_5359,N_5072,N_5144);
and U5360 (N_5360,N_5060,N_5115);
nand U5361 (N_5361,N_5161,N_5046);
or U5362 (N_5362,N_5159,N_5034);
nor U5363 (N_5363,N_5191,N_5107);
nand U5364 (N_5364,N_5152,N_5142);
and U5365 (N_5365,N_5116,N_5071);
and U5366 (N_5366,N_5118,N_5057);
or U5367 (N_5367,N_5137,N_5050);
and U5368 (N_5368,N_5086,N_5061);
and U5369 (N_5369,N_5197,N_5160);
nand U5370 (N_5370,N_5043,N_5040);
xor U5371 (N_5371,N_5019,N_5176);
and U5372 (N_5372,N_5026,N_5056);
nand U5373 (N_5373,N_5246,N_5045);
nor U5374 (N_5374,N_5187,N_5087);
nor U5375 (N_5375,N_5228,N_5124);
xnor U5376 (N_5376,N_5212,N_5030);
nor U5377 (N_5377,N_5103,N_5070);
or U5378 (N_5378,N_5233,N_5006);
xor U5379 (N_5379,N_5046,N_5069);
nor U5380 (N_5380,N_5200,N_5202);
or U5381 (N_5381,N_5069,N_5125);
nand U5382 (N_5382,N_5045,N_5234);
and U5383 (N_5383,N_5073,N_5134);
or U5384 (N_5384,N_5149,N_5085);
and U5385 (N_5385,N_5088,N_5233);
nand U5386 (N_5386,N_5242,N_5232);
or U5387 (N_5387,N_5216,N_5178);
or U5388 (N_5388,N_5115,N_5047);
and U5389 (N_5389,N_5113,N_5008);
nand U5390 (N_5390,N_5176,N_5186);
nor U5391 (N_5391,N_5023,N_5073);
nand U5392 (N_5392,N_5200,N_5134);
and U5393 (N_5393,N_5193,N_5204);
nor U5394 (N_5394,N_5108,N_5097);
nand U5395 (N_5395,N_5225,N_5234);
or U5396 (N_5396,N_5166,N_5108);
xor U5397 (N_5397,N_5114,N_5016);
or U5398 (N_5398,N_5082,N_5022);
nor U5399 (N_5399,N_5161,N_5190);
nand U5400 (N_5400,N_5184,N_5158);
nor U5401 (N_5401,N_5041,N_5001);
and U5402 (N_5402,N_5141,N_5129);
nor U5403 (N_5403,N_5153,N_5110);
or U5404 (N_5404,N_5110,N_5248);
nand U5405 (N_5405,N_5215,N_5197);
or U5406 (N_5406,N_5187,N_5004);
and U5407 (N_5407,N_5212,N_5177);
or U5408 (N_5408,N_5059,N_5163);
and U5409 (N_5409,N_5170,N_5133);
or U5410 (N_5410,N_5167,N_5248);
xnor U5411 (N_5411,N_5106,N_5065);
or U5412 (N_5412,N_5042,N_5072);
nor U5413 (N_5413,N_5121,N_5148);
and U5414 (N_5414,N_5188,N_5053);
xor U5415 (N_5415,N_5225,N_5053);
xnor U5416 (N_5416,N_5107,N_5231);
nor U5417 (N_5417,N_5026,N_5058);
xor U5418 (N_5418,N_5013,N_5119);
or U5419 (N_5419,N_5234,N_5244);
or U5420 (N_5420,N_5055,N_5176);
and U5421 (N_5421,N_5196,N_5181);
and U5422 (N_5422,N_5013,N_5077);
nor U5423 (N_5423,N_5096,N_5217);
and U5424 (N_5424,N_5208,N_5090);
and U5425 (N_5425,N_5175,N_5088);
or U5426 (N_5426,N_5159,N_5091);
or U5427 (N_5427,N_5045,N_5137);
and U5428 (N_5428,N_5153,N_5244);
nor U5429 (N_5429,N_5126,N_5110);
and U5430 (N_5430,N_5114,N_5102);
or U5431 (N_5431,N_5038,N_5193);
or U5432 (N_5432,N_5117,N_5165);
or U5433 (N_5433,N_5055,N_5086);
or U5434 (N_5434,N_5206,N_5040);
or U5435 (N_5435,N_5010,N_5122);
or U5436 (N_5436,N_5070,N_5023);
nand U5437 (N_5437,N_5175,N_5125);
nor U5438 (N_5438,N_5070,N_5041);
or U5439 (N_5439,N_5243,N_5161);
nand U5440 (N_5440,N_5043,N_5129);
or U5441 (N_5441,N_5033,N_5160);
and U5442 (N_5442,N_5010,N_5191);
nand U5443 (N_5443,N_5005,N_5086);
nand U5444 (N_5444,N_5153,N_5220);
xor U5445 (N_5445,N_5151,N_5021);
and U5446 (N_5446,N_5173,N_5207);
xnor U5447 (N_5447,N_5157,N_5136);
nand U5448 (N_5448,N_5221,N_5151);
nor U5449 (N_5449,N_5159,N_5200);
xor U5450 (N_5450,N_5138,N_5090);
or U5451 (N_5451,N_5082,N_5028);
and U5452 (N_5452,N_5202,N_5152);
and U5453 (N_5453,N_5102,N_5214);
nor U5454 (N_5454,N_5014,N_5248);
nor U5455 (N_5455,N_5156,N_5145);
xor U5456 (N_5456,N_5040,N_5106);
nand U5457 (N_5457,N_5183,N_5119);
nor U5458 (N_5458,N_5078,N_5121);
and U5459 (N_5459,N_5129,N_5110);
and U5460 (N_5460,N_5070,N_5059);
nor U5461 (N_5461,N_5190,N_5109);
or U5462 (N_5462,N_5157,N_5189);
and U5463 (N_5463,N_5219,N_5172);
nand U5464 (N_5464,N_5100,N_5055);
xor U5465 (N_5465,N_5064,N_5191);
xor U5466 (N_5466,N_5177,N_5209);
nand U5467 (N_5467,N_5068,N_5220);
or U5468 (N_5468,N_5013,N_5030);
nand U5469 (N_5469,N_5157,N_5137);
nor U5470 (N_5470,N_5074,N_5240);
and U5471 (N_5471,N_5157,N_5151);
and U5472 (N_5472,N_5242,N_5218);
xor U5473 (N_5473,N_5135,N_5209);
nand U5474 (N_5474,N_5235,N_5035);
nand U5475 (N_5475,N_5008,N_5081);
and U5476 (N_5476,N_5012,N_5168);
nand U5477 (N_5477,N_5248,N_5136);
and U5478 (N_5478,N_5096,N_5184);
nand U5479 (N_5479,N_5242,N_5070);
nor U5480 (N_5480,N_5029,N_5191);
nand U5481 (N_5481,N_5116,N_5064);
nor U5482 (N_5482,N_5208,N_5095);
xor U5483 (N_5483,N_5148,N_5100);
or U5484 (N_5484,N_5219,N_5043);
or U5485 (N_5485,N_5224,N_5002);
and U5486 (N_5486,N_5246,N_5087);
or U5487 (N_5487,N_5052,N_5223);
or U5488 (N_5488,N_5219,N_5115);
nor U5489 (N_5489,N_5111,N_5046);
or U5490 (N_5490,N_5223,N_5141);
nand U5491 (N_5491,N_5046,N_5123);
nand U5492 (N_5492,N_5018,N_5132);
xnor U5493 (N_5493,N_5218,N_5105);
nor U5494 (N_5494,N_5182,N_5208);
or U5495 (N_5495,N_5140,N_5243);
nor U5496 (N_5496,N_5244,N_5098);
and U5497 (N_5497,N_5120,N_5012);
nor U5498 (N_5498,N_5182,N_5216);
xor U5499 (N_5499,N_5159,N_5015);
or U5500 (N_5500,N_5473,N_5326);
and U5501 (N_5501,N_5487,N_5430);
nand U5502 (N_5502,N_5446,N_5359);
or U5503 (N_5503,N_5346,N_5481);
nand U5504 (N_5504,N_5496,N_5490);
or U5505 (N_5505,N_5288,N_5470);
nor U5506 (N_5506,N_5298,N_5493);
or U5507 (N_5507,N_5335,N_5427);
and U5508 (N_5508,N_5349,N_5374);
nor U5509 (N_5509,N_5268,N_5306);
xnor U5510 (N_5510,N_5278,N_5485);
or U5511 (N_5511,N_5403,N_5489);
xnor U5512 (N_5512,N_5469,N_5358);
and U5513 (N_5513,N_5297,N_5448);
and U5514 (N_5514,N_5354,N_5286);
nor U5515 (N_5515,N_5285,N_5364);
xnor U5516 (N_5516,N_5463,N_5416);
or U5517 (N_5517,N_5435,N_5299);
and U5518 (N_5518,N_5425,N_5263);
nor U5519 (N_5519,N_5353,N_5424);
nor U5520 (N_5520,N_5325,N_5480);
nor U5521 (N_5521,N_5375,N_5382);
xor U5522 (N_5522,N_5466,N_5377);
xnor U5523 (N_5523,N_5401,N_5373);
nand U5524 (N_5524,N_5414,N_5344);
xnor U5525 (N_5525,N_5494,N_5476);
or U5526 (N_5526,N_5402,N_5351);
or U5527 (N_5527,N_5292,N_5295);
or U5528 (N_5528,N_5331,N_5317);
and U5529 (N_5529,N_5314,N_5363);
nand U5530 (N_5530,N_5318,N_5337);
nand U5531 (N_5531,N_5275,N_5342);
nor U5532 (N_5532,N_5459,N_5405);
xnor U5533 (N_5533,N_5366,N_5406);
nand U5534 (N_5534,N_5433,N_5483);
nor U5535 (N_5535,N_5413,N_5323);
or U5536 (N_5536,N_5350,N_5251);
xor U5537 (N_5537,N_5332,N_5407);
and U5538 (N_5538,N_5365,N_5289);
xor U5539 (N_5539,N_5301,N_5256);
nand U5540 (N_5540,N_5451,N_5412);
xnor U5541 (N_5541,N_5294,N_5415);
nand U5542 (N_5542,N_5453,N_5432);
and U5543 (N_5543,N_5362,N_5400);
nor U5544 (N_5544,N_5258,N_5368);
and U5545 (N_5545,N_5272,N_5262);
nand U5546 (N_5546,N_5454,N_5360);
nor U5547 (N_5547,N_5369,N_5273);
or U5548 (N_5548,N_5443,N_5334);
or U5549 (N_5549,N_5269,N_5449);
nor U5550 (N_5550,N_5302,N_5252);
nor U5551 (N_5551,N_5274,N_5361);
and U5552 (N_5552,N_5300,N_5441);
nor U5553 (N_5553,N_5431,N_5267);
nor U5554 (N_5554,N_5277,N_5456);
nand U5555 (N_5555,N_5270,N_5253);
nor U5556 (N_5556,N_5305,N_5303);
and U5557 (N_5557,N_5357,N_5339);
nand U5558 (N_5558,N_5265,N_5257);
nor U5559 (N_5559,N_5444,N_5462);
or U5560 (N_5560,N_5276,N_5338);
nand U5561 (N_5561,N_5290,N_5486);
xnor U5562 (N_5562,N_5310,N_5419);
nand U5563 (N_5563,N_5313,N_5452);
or U5564 (N_5564,N_5395,N_5495);
nand U5565 (N_5565,N_5384,N_5468);
nand U5566 (N_5566,N_5399,N_5381);
xnor U5567 (N_5567,N_5386,N_5421);
xnor U5568 (N_5568,N_5343,N_5385);
nor U5569 (N_5569,N_5409,N_5340);
or U5570 (N_5570,N_5308,N_5330);
and U5571 (N_5571,N_5254,N_5304);
nand U5572 (N_5572,N_5376,N_5355);
nand U5573 (N_5573,N_5387,N_5367);
and U5574 (N_5574,N_5478,N_5333);
nand U5575 (N_5575,N_5460,N_5250);
nand U5576 (N_5576,N_5372,N_5284);
and U5577 (N_5577,N_5404,N_5482);
nand U5578 (N_5578,N_5315,N_5309);
and U5579 (N_5579,N_5390,N_5396);
xor U5580 (N_5580,N_5345,N_5442);
or U5581 (N_5581,N_5434,N_5394);
or U5582 (N_5582,N_5464,N_5436);
and U5583 (N_5583,N_5411,N_5423);
and U5584 (N_5584,N_5388,N_5324);
or U5585 (N_5585,N_5266,N_5371);
nand U5586 (N_5586,N_5474,N_5488);
and U5587 (N_5587,N_5260,N_5471);
nand U5588 (N_5588,N_5499,N_5450);
nor U5589 (N_5589,N_5497,N_5370);
and U5590 (N_5590,N_5465,N_5428);
and U5591 (N_5591,N_5417,N_5479);
or U5592 (N_5592,N_5408,N_5279);
and U5593 (N_5593,N_5356,N_5477);
and U5594 (N_5594,N_5312,N_5475);
or U5595 (N_5595,N_5491,N_5282);
nand U5596 (N_5596,N_5319,N_5391);
and U5597 (N_5597,N_5379,N_5341);
nor U5598 (N_5598,N_5445,N_5280);
nor U5599 (N_5599,N_5393,N_5307);
and U5600 (N_5600,N_5422,N_5316);
and U5601 (N_5601,N_5296,N_5392);
and U5602 (N_5602,N_5455,N_5380);
or U5603 (N_5603,N_5458,N_5329);
nand U5604 (N_5604,N_5320,N_5410);
nor U5605 (N_5605,N_5438,N_5281);
and U5606 (N_5606,N_5447,N_5322);
nor U5607 (N_5607,N_5283,N_5264);
xnor U5608 (N_5608,N_5398,N_5327);
nand U5609 (N_5609,N_5347,N_5321);
nand U5610 (N_5610,N_5492,N_5389);
and U5611 (N_5611,N_5418,N_5348);
nand U5612 (N_5612,N_5352,N_5498);
nand U5613 (N_5613,N_5472,N_5328);
and U5614 (N_5614,N_5437,N_5484);
and U5615 (N_5615,N_5439,N_5467);
and U5616 (N_5616,N_5261,N_5426);
nor U5617 (N_5617,N_5429,N_5293);
xnor U5618 (N_5618,N_5457,N_5383);
or U5619 (N_5619,N_5311,N_5397);
nor U5620 (N_5620,N_5287,N_5291);
nor U5621 (N_5621,N_5271,N_5440);
nand U5622 (N_5622,N_5461,N_5259);
and U5623 (N_5623,N_5255,N_5336);
and U5624 (N_5624,N_5378,N_5420);
and U5625 (N_5625,N_5360,N_5430);
or U5626 (N_5626,N_5417,N_5269);
and U5627 (N_5627,N_5469,N_5346);
nand U5628 (N_5628,N_5405,N_5283);
and U5629 (N_5629,N_5320,N_5345);
nor U5630 (N_5630,N_5315,N_5284);
nor U5631 (N_5631,N_5467,N_5266);
nor U5632 (N_5632,N_5490,N_5455);
or U5633 (N_5633,N_5389,N_5262);
or U5634 (N_5634,N_5456,N_5317);
or U5635 (N_5635,N_5376,N_5278);
or U5636 (N_5636,N_5476,N_5357);
nor U5637 (N_5637,N_5402,N_5391);
nor U5638 (N_5638,N_5456,N_5315);
nand U5639 (N_5639,N_5284,N_5309);
nor U5640 (N_5640,N_5337,N_5379);
nand U5641 (N_5641,N_5344,N_5278);
and U5642 (N_5642,N_5387,N_5456);
nand U5643 (N_5643,N_5447,N_5430);
nand U5644 (N_5644,N_5489,N_5397);
nor U5645 (N_5645,N_5251,N_5324);
nand U5646 (N_5646,N_5398,N_5460);
or U5647 (N_5647,N_5473,N_5308);
and U5648 (N_5648,N_5394,N_5385);
nor U5649 (N_5649,N_5277,N_5352);
nand U5650 (N_5650,N_5338,N_5340);
and U5651 (N_5651,N_5300,N_5285);
nand U5652 (N_5652,N_5418,N_5424);
or U5653 (N_5653,N_5400,N_5324);
and U5654 (N_5654,N_5260,N_5477);
and U5655 (N_5655,N_5254,N_5363);
nand U5656 (N_5656,N_5418,N_5334);
nor U5657 (N_5657,N_5339,N_5476);
xor U5658 (N_5658,N_5463,N_5411);
and U5659 (N_5659,N_5276,N_5480);
nand U5660 (N_5660,N_5302,N_5365);
xnor U5661 (N_5661,N_5269,N_5426);
or U5662 (N_5662,N_5481,N_5336);
nor U5663 (N_5663,N_5346,N_5375);
or U5664 (N_5664,N_5365,N_5369);
or U5665 (N_5665,N_5480,N_5495);
nor U5666 (N_5666,N_5414,N_5322);
nand U5667 (N_5667,N_5270,N_5414);
or U5668 (N_5668,N_5425,N_5452);
nand U5669 (N_5669,N_5464,N_5460);
xor U5670 (N_5670,N_5274,N_5464);
or U5671 (N_5671,N_5351,N_5413);
nand U5672 (N_5672,N_5294,N_5448);
nor U5673 (N_5673,N_5294,N_5371);
or U5674 (N_5674,N_5396,N_5442);
or U5675 (N_5675,N_5254,N_5464);
or U5676 (N_5676,N_5297,N_5260);
nand U5677 (N_5677,N_5328,N_5454);
or U5678 (N_5678,N_5347,N_5465);
nor U5679 (N_5679,N_5499,N_5442);
and U5680 (N_5680,N_5493,N_5443);
nor U5681 (N_5681,N_5497,N_5291);
nor U5682 (N_5682,N_5492,N_5277);
nor U5683 (N_5683,N_5356,N_5461);
nand U5684 (N_5684,N_5275,N_5457);
nor U5685 (N_5685,N_5398,N_5294);
nand U5686 (N_5686,N_5379,N_5459);
or U5687 (N_5687,N_5424,N_5408);
xnor U5688 (N_5688,N_5471,N_5328);
xor U5689 (N_5689,N_5372,N_5322);
nor U5690 (N_5690,N_5456,N_5464);
or U5691 (N_5691,N_5273,N_5480);
nand U5692 (N_5692,N_5450,N_5401);
and U5693 (N_5693,N_5427,N_5435);
or U5694 (N_5694,N_5468,N_5434);
nor U5695 (N_5695,N_5347,N_5411);
nor U5696 (N_5696,N_5312,N_5470);
nor U5697 (N_5697,N_5361,N_5359);
nand U5698 (N_5698,N_5306,N_5372);
or U5699 (N_5699,N_5478,N_5499);
nand U5700 (N_5700,N_5401,N_5355);
nor U5701 (N_5701,N_5445,N_5297);
nand U5702 (N_5702,N_5363,N_5306);
nor U5703 (N_5703,N_5276,N_5431);
or U5704 (N_5704,N_5410,N_5289);
nor U5705 (N_5705,N_5382,N_5282);
or U5706 (N_5706,N_5454,N_5456);
nor U5707 (N_5707,N_5460,N_5336);
or U5708 (N_5708,N_5378,N_5439);
or U5709 (N_5709,N_5283,N_5418);
or U5710 (N_5710,N_5481,N_5443);
or U5711 (N_5711,N_5417,N_5491);
and U5712 (N_5712,N_5369,N_5262);
nor U5713 (N_5713,N_5307,N_5256);
and U5714 (N_5714,N_5407,N_5471);
nor U5715 (N_5715,N_5270,N_5326);
xnor U5716 (N_5716,N_5405,N_5422);
nand U5717 (N_5717,N_5494,N_5292);
xor U5718 (N_5718,N_5318,N_5260);
or U5719 (N_5719,N_5482,N_5331);
nand U5720 (N_5720,N_5320,N_5349);
nand U5721 (N_5721,N_5366,N_5479);
or U5722 (N_5722,N_5499,N_5256);
nor U5723 (N_5723,N_5405,N_5268);
or U5724 (N_5724,N_5498,N_5266);
or U5725 (N_5725,N_5489,N_5265);
or U5726 (N_5726,N_5449,N_5283);
xor U5727 (N_5727,N_5436,N_5296);
nor U5728 (N_5728,N_5269,N_5253);
nor U5729 (N_5729,N_5434,N_5412);
or U5730 (N_5730,N_5370,N_5454);
nand U5731 (N_5731,N_5475,N_5455);
and U5732 (N_5732,N_5250,N_5468);
or U5733 (N_5733,N_5304,N_5272);
nand U5734 (N_5734,N_5263,N_5312);
or U5735 (N_5735,N_5429,N_5346);
or U5736 (N_5736,N_5423,N_5485);
nand U5737 (N_5737,N_5319,N_5378);
nor U5738 (N_5738,N_5370,N_5282);
xor U5739 (N_5739,N_5277,N_5288);
or U5740 (N_5740,N_5486,N_5313);
and U5741 (N_5741,N_5484,N_5449);
and U5742 (N_5742,N_5472,N_5378);
nor U5743 (N_5743,N_5298,N_5424);
and U5744 (N_5744,N_5329,N_5280);
nand U5745 (N_5745,N_5491,N_5425);
nand U5746 (N_5746,N_5269,N_5309);
xor U5747 (N_5747,N_5488,N_5499);
or U5748 (N_5748,N_5396,N_5303);
nand U5749 (N_5749,N_5325,N_5413);
nand U5750 (N_5750,N_5702,N_5549);
or U5751 (N_5751,N_5536,N_5643);
or U5752 (N_5752,N_5617,N_5583);
nand U5753 (N_5753,N_5748,N_5649);
nor U5754 (N_5754,N_5656,N_5640);
xnor U5755 (N_5755,N_5634,N_5519);
and U5756 (N_5756,N_5500,N_5689);
nor U5757 (N_5757,N_5540,N_5569);
nor U5758 (N_5758,N_5693,N_5651);
and U5759 (N_5759,N_5511,N_5558);
nor U5760 (N_5760,N_5650,N_5706);
or U5761 (N_5761,N_5683,N_5692);
xnor U5762 (N_5762,N_5703,N_5741);
and U5763 (N_5763,N_5560,N_5588);
nand U5764 (N_5764,N_5523,N_5648);
xnor U5765 (N_5765,N_5553,N_5713);
or U5766 (N_5766,N_5591,N_5631);
or U5767 (N_5767,N_5654,N_5611);
nor U5768 (N_5768,N_5720,N_5691);
and U5769 (N_5769,N_5736,N_5719);
nor U5770 (N_5770,N_5502,N_5635);
xor U5771 (N_5771,N_5724,N_5729);
or U5772 (N_5772,N_5595,N_5512);
and U5773 (N_5773,N_5527,N_5671);
nor U5774 (N_5774,N_5605,N_5644);
or U5775 (N_5775,N_5725,N_5509);
nand U5776 (N_5776,N_5579,N_5515);
or U5777 (N_5777,N_5716,N_5590);
nor U5778 (N_5778,N_5710,N_5593);
nor U5779 (N_5779,N_5701,N_5533);
and U5780 (N_5780,N_5623,N_5526);
nand U5781 (N_5781,N_5534,N_5561);
nor U5782 (N_5782,N_5525,N_5676);
nand U5783 (N_5783,N_5721,N_5615);
or U5784 (N_5784,N_5550,N_5673);
nor U5785 (N_5785,N_5618,N_5520);
xor U5786 (N_5786,N_5598,N_5602);
or U5787 (N_5787,N_5684,N_5685);
nand U5788 (N_5788,N_5687,N_5697);
or U5789 (N_5789,N_5557,N_5711);
xor U5790 (N_5790,N_5597,N_5739);
nand U5791 (N_5791,N_5562,N_5600);
or U5792 (N_5792,N_5504,N_5688);
nand U5793 (N_5793,N_5638,N_5660);
or U5794 (N_5794,N_5606,N_5532);
nand U5795 (N_5795,N_5528,N_5573);
xor U5796 (N_5796,N_5670,N_5581);
and U5797 (N_5797,N_5546,N_5530);
or U5798 (N_5798,N_5543,N_5521);
or U5799 (N_5799,N_5657,N_5744);
and U5800 (N_5800,N_5517,N_5548);
or U5801 (N_5801,N_5636,N_5728);
nand U5802 (N_5802,N_5659,N_5535);
xnor U5803 (N_5803,N_5686,N_5646);
nor U5804 (N_5804,N_5596,N_5503);
or U5805 (N_5805,N_5514,N_5576);
xnor U5806 (N_5806,N_5614,N_5545);
nand U5807 (N_5807,N_5622,N_5608);
nor U5808 (N_5808,N_5531,N_5680);
nand U5809 (N_5809,N_5541,N_5612);
nand U5810 (N_5810,N_5620,N_5538);
nor U5811 (N_5811,N_5506,N_5580);
or U5812 (N_5812,N_5505,N_5658);
xnor U5813 (N_5813,N_5575,N_5507);
nand U5814 (N_5814,N_5664,N_5607);
or U5815 (N_5815,N_5743,N_5542);
or U5816 (N_5816,N_5574,N_5735);
nand U5817 (N_5817,N_5669,N_5699);
and U5818 (N_5818,N_5647,N_5653);
xnor U5819 (N_5819,N_5714,N_5592);
xnor U5820 (N_5820,N_5740,N_5707);
or U5821 (N_5821,N_5529,N_5737);
and U5822 (N_5822,N_5604,N_5621);
or U5823 (N_5823,N_5537,N_5616);
or U5824 (N_5824,N_5566,N_5601);
and U5825 (N_5825,N_5556,N_5572);
nand U5826 (N_5826,N_5747,N_5565);
or U5827 (N_5827,N_5630,N_5722);
and U5828 (N_5828,N_5661,N_5539);
nand U5829 (N_5829,N_5715,N_5682);
and U5830 (N_5830,N_5637,N_5641);
nand U5831 (N_5831,N_5609,N_5555);
nor U5832 (N_5832,N_5742,N_5632);
nor U5833 (N_5833,N_5522,N_5586);
xnor U5834 (N_5834,N_5589,N_5610);
nor U5835 (N_5835,N_5745,N_5749);
and U5836 (N_5836,N_5655,N_5732);
and U5837 (N_5837,N_5627,N_5567);
nand U5838 (N_5838,N_5578,N_5628);
nand U5839 (N_5839,N_5571,N_5564);
nor U5840 (N_5840,N_5624,N_5613);
or U5841 (N_5841,N_5679,N_5662);
or U5842 (N_5842,N_5667,N_5674);
or U5843 (N_5843,N_5551,N_5508);
nand U5844 (N_5844,N_5663,N_5645);
nor U5845 (N_5845,N_5652,N_5585);
nor U5846 (N_5846,N_5570,N_5625);
or U5847 (N_5847,N_5633,N_5516);
or U5848 (N_5848,N_5681,N_5524);
nor U5849 (N_5849,N_5700,N_5594);
or U5850 (N_5850,N_5518,N_5587);
or U5851 (N_5851,N_5709,N_5501);
nor U5852 (N_5852,N_5568,N_5734);
and U5853 (N_5853,N_5727,N_5544);
and U5854 (N_5854,N_5603,N_5712);
nand U5855 (N_5855,N_5723,N_5746);
nor U5856 (N_5856,N_5554,N_5718);
nand U5857 (N_5857,N_5599,N_5690);
and U5858 (N_5858,N_5547,N_5675);
nand U5859 (N_5859,N_5559,N_5629);
and U5860 (N_5860,N_5510,N_5619);
nor U5861 (N_5861,N_5665,N_5696);
nor U5862 (N_5862,N_5705,N_5731);
nor U5863 (N_5863,N_5552,N_5733);
nand U5864 (N_5864,N_5730,N_5695);
and U5865 (N_5865,N_5582,N_5672);
nor U5866 (N_5866,N_5678,N_5698);
nor U5867 (N_5867,N_5563,N_5639);
nor U5868 (N_5868,N_5694,N_5642);
nor U5869 (N_5869,N_5738,N_5717);
or U5870 (N_5870,N_5584,N_5677);
nand U5871 (N_5871,N_5513,N_5666);
and U5872 (N_5872,N_5577,N_5704);
nor U5873 (N_5873,N_5626,N_5708);
and U5874 (N_5874,N_5726,N_5668);
nand U5875 (N_5875,N_5683,N_5745);
and U5876 (N_5876,N_5624,N_5529);
nor U5877 (N_5877,N_5638,N_5742);
xor U5878 (N_5878,N_5539,N_5573);
xnor U5879 (N_5879,N_5653,N_5628);
and U5880 (N_5880,N_5533,N_5690);
nand U5881 (N_5881,N_5616,N_5644);
nor U5882 (N_5882,N_5694,N_5606);
xnor U5883 (N_5883,N_5591,N_5646);
and U5884 (N_5884,N_5582,N_5511);
nand U5885 (N_5885,N_5737,N_5686);
nor U5886 (N_5886,N_5590,N_5597);
or U5887 (N_5887,N_5613,N_5625);
nor U5888 (N_5888,N_5741,N_5642);
nor U5889 (N_5889,N_5715,N_5676);
nand U5890 (N_5890,N_5642,N_5682);
and U5891 (N_5891,N_5570,N_5599);
or U5892 (N_5892,N_5628,N_5531);
nand U5893 (N_5893,N_5578,N_5576);
or U5894 (N_5894,N_5586,N_5631);
xnor U5895 (N_5895,N_5612,N_5565);
nor U5896 (N_5896,N_5542,N_5585);
nand U5897 (N_5897,N_5573,N_5685);
xor U5898 (N_5898,N_5625,N_5623);
nor U5899 (N_5899,N_5714,N_5576);
nor U5900 (N_5900,N_5582,N_5584);
nand U5901 (N_5901,N_5554,N_5612);
or U5902 (N_5902,N_5594,N_5716);
or U5903 (N_5903,N_5572,N_5602);
nor U5904 (N_5904,N_5716,N_5562);
or U5905 (N_5905,N_5597,N_5668);
nand U5906 (N_5906,N_5583,N_5650);
and U5907 (N_5907,N_5670,N_5522);
or U5908 (N_5908,N_5726,N_5532);
and U5909 (N_5909,N_5585,N_5678);
or U5910 (N_5910,N_5601,N_5673);
xor U5911 (N_5911,N_5610,N_5732);
and U5912 (N_5912,N_5733,N_5702);
or U5913 (N_5913,N_5519,N_5539);
nor U5914 (N_5914,N_5517,N_5668);
and U5915 (N_5915,N_5525,N_5654);
or U5916 (N_5916,N_5660,N_5689);
nor U5917 (N_5917,N_5729,N_5602);
and U5918 (N_5918,N_5535,N_5714);
or U5919 (N_5919,N_5660,N_5720);
nand U5920 (N_5920,N_5689,N_5566);
or U5921 (N_5921,N_5682,N_5515);
and U5922 (N_5922,N_5550,N_5729);
nor U5923 (N_5923,N_5625,N_5636);
nor U5924 (N_5924,N_5525,N_5603);
xor U5925 (N_5925,N_5596,N_5598);
and U5926 (N_5926,N_5736,N_5562);
nand U5927 (N_5927,N_5695,N_5529);
nand U5928 (N_5928,N_5587,N_5606);
and U5929 (N_5929,N_5699,N_5628);
and U5930 (N_5930,N_5718,N_5679);
xnor U5931 (N_5931,N_5724,N_5635);
nand U5932 (N_5932,N_5668,N_5682);
nand U5933 (N_5933,N_5617,N_5679);
nor U5934 (N_5934,N_5608,N_5549);
or U5935 (N_5935,N_5712,N_5601);
nand U5936 (N_5936,N_5621,N_5666);
nor U5937 (N_5937,N_5737,N_5679);
xor U5938 (N_5938,N_5564,N_5684);
and U5939 (N_5939,N_5555,N_5696);
and U5940 (N_5940,N_5559,N_5649);
or U5941 (N_5941,N_5579,N_5508);
nand U5942 (N_5942,N_5641,N_5564);
nand U5943 (N_5943,N_5692,N_5661);
nand U5944 (N_5944,N_5675,N_5506);
xnor U5945 (N_5945,N_5572,N_5606);
nand U5946 (N_5946,N_5631,N_5657);
nor U5947 (N_5947,N_5591,N_5511);
or U5948 (N_5948,N_5697,N_5617);
xnor U5949 (N_5949,N_5520,N_5594);
nand U5950 (N_5950,N_5656,N_5627);
or U5951 (N_5951,N_5727,N_5700);
nand U5952 (N_5952,N_5576,N_5659);
and U5953 (N_5953,N_5624,N_5692);
and U5954 (N_5954,N_5684,N_5532);
and U5955 (N_5955,N_5518,N_5628);
and U5956 (N_5956,N_5685,N_5526);
nand U5957 (N_5957,N_5741,N_5663);
or U5958 (N_5958,N_5708,N_5518);
and U5959 (N_5959,N_5603,N_5700);
nor U5960 (N_5960,N_5504,N_5556);
or U5961 (N_5961,N_5719,N_5589);
or U5962 (N_5962,N_5515,N_5529);
xor U5963 (N_5963,N_5627,N_5620);
nand U5964 (N_5964,N_5546,N_5525);
and U5965 (N_5965,N_5715,N_5705);
xor U5966 (N_5966,N_5668,N_5664);
xnor U5967 (N_5967,N_5674,N_5528);
or U5968 (N_5968,N_5602,N_5627);
nand U5969 (N_5969,N_5583,N_5660);
nor U5970 (N_5970,N_5634,N_5627);
nand U5971 (N_5971,N_5703,N_5600);
and U5972 (N_5972,N_5729,N_5643);
nor U5973 (N_5973,N_5557,N_5520);
xnor U5974 (N_5974,N_5633,N_5660);
nor U5975 (N_5975,N_5545,N_5654);
nor U5976 (N_5976,N_5662,N_5513);
and U5977 (N_5977,N_5579,N_5641);
nor U5978 (N_5978,N_5685,N_5687);
nor U5979 (N_5979,N_5664,N_5723);
and U5980 (N_5980,N_5576,N_5532);
and U5981 (N_5981,N_5630,N_5515);
or U5982 (N_5982,N_5644,N_5688);
and U5983 (N_5983,N_5525,N_5549);
nand U5984 (N_5984,N_5554,N_5530);
or U5985 (N_5985,N_5716,N_5596);
or U5986 (N_5986,N_5529,N_5556);
and U5987 (N_5987,N_5613,N_5657);
nand U5988 (N_5988,N_5522,N_5729);
or U5989 (N_5989,N_5582,N_5551);
and U5990 (N_5990,N_5731,N_5720);
nor U5991 (N_5991,N_5528,N_5525);
nand U5992 (N_5992,N_5634,N_5595);
xor U5993 (N_5993,N_5517,N_5520);
nand U5994 (N_5994,N_5688,N_5733);
and U5995 (N_5995,N_5566,N_5596);
or U5996 (N_5996,N_5654,N_5640);
nor U5997 (N_5997,N_5560,N_5687);
xnor U5998 (N_5998,N_5572,N_5726);
nand U5999 (N_5999,N_5623,N_5743);
nand U6000 (N_6000,N_5808,N_5814);
and U6001 (N_6001,N_5932,N_5950);
nor U6002 (N_6002,N_5949,N_5904);
xor U6003 (N_6003,N_5910,N_5793);
and U6004 (N_6004,N_5789,N_5752);
and U6005 (N_6005,N_5943,N_5867);
nand U6006 (N_6006,N_5925,N_5885);
xnor U6007 (N_6007,N_5948,N_5962);
or U6008 (N_6008,N_5770,N_5985);
or U6009 (N_6009,N_5824,N_5795);
nand U6010 (N_6010,N_5807,N_5975);
nor U6011 (N_6011,N_5883,N_5783);
nand U6012 (N_6012,N_5862,N_5777);
nor U6013 (N_6013,N_5798,N_5858);
xor U6014 (N_6014,N_5919,N_5857);
or U6015 (N_6015,N_5846,N_5983);
nand U6016 (N_6016,N_5847,N_5986);
or U6017 (N_6017,N_5960,N_5889);
and U6018 (N_6018,N_5827,N_5923);
xnor U6019 (N_6019,N_5840,N_5816);
and U6020 (N_6020,N_5900,N_5912);
nor U6021 (N_6021,N_5915,N_5757);
nor U6022 (N_6022,N_5895,N_5945);
nor U6023 (N_6023,N_5917,N_5878);
or U6024 (N_6024,N_5781,N_5829);
or U6025 (N_6025,N_5864,N_5787);
xor U6026 (N_6026,N_5812,N_5921);
nand U6027 (N_6027,N_5930,N_5784);
xor U6028 (N_6028,N_5767,N_5868);
and U6029 (N_6029,N_5905,N_5833);
nand U6030 (N_6030,N_5936,N_5791);
or U6031 (N_6031,N_5761,N_5966);
or U6032 (N_6032,N_5974,N_5804);
nor U6033 (N_6033,N_5753,N_5838);
or U6034 (N_6034,N_5815,N_5859);
nand U6035 (N_6035,N_5852,N_5913);
nand U6036 (N_6036,N_5990,N_5995);
nor U6037 (N_6037,N_5882,N_5877);
nand U6038 (N_6038,N_5773,N_5786);
and U6039 (N_6039,N_5794,N_5834);
or U6040 (N_6040,N_5954,N_5965);
nand U6041 (N_6041,N_5785,N_5763);
nand U6042 (N_6042,N_5780,N_5931);
and U6043 (N_6043,N_5832,N_5826);
nand U6044 (N_6044,N_5916,N_5978);
nand U6045 (N_6045,N_5874,N_5750);
nand U6046 (N_6046,N_5902,N_5860);
and U6047 (N_6047,N_5766,N_5853);
xor U6048 (N_6048,N_5825,N_5979);
or U6049 (N_6049,N_5911,N_5881);
xor U6050 (N_6050,N_5891,N_5755);
nor U6051 (N_6051,N_5926,N_5981);
nor U6052 (N_6052,N_5823,N_5813);
and U6053 (N_6053,N_5776,N_5788);
or U6054 (N_6054,N_5946,N_5952);
nand U6055 (N_6055,N_5951,N_5872);
and U6056 (N_6056,N_5959,N_5774);
and U6057 (N_6057,N_5821,N_5903);
nor U6058 (N_6058,N_5969,N_5875);
nand U6059 (N_6059,N_5841,N_5897);
nand U6060 (N_6060,N_5811,N_5848);
or U6061 (N_6061,N_5850,N_5751);
nor U6062 (N_6062,N_5802,N_5797);
and U6063 (N_6063,N_5775,N_5982);
xor U6064 (N_6064,N_5768,N_5764);
nor U6065 (N_6065,N_5844,N_5928);
and U6066 (N_6066,N_5935,N_5842);
xor U6067 (N_6067,N_5855,N_5765);
nand U6068 (N_6068,N_5849,N_5817);
nor U6069 (N_6069,N_5861,N_5898);
or U6070 (N_6070,N_5800,N_5828);
or U6071 (N_6071,N_5984,N_5994);
and U6072 (N_6072,N_5754,N_5933);
nand U6073 (N_6073,N_5956,N_5799);
or U6074 (N_6074,N_5830,N_5908);
nand U6075 (N_6075,N_5820,N_5914);
and U6076 (N_6076,N_5888,N_5958);
nand U6077 (N_6077,N_5760,N_5927);
xor U6078 (N_6078,N_5890,N_5924);
nand U6079 (N_6079,N_5884,N_5992);
and U6080 (N_6080,N_5909,N_5976);
nand U6081 (N_6081,N_5906,N_5866);
or U6082 (N_6082,N_5977,N_5769);
nor U6083 (N_6083,N_5886,N_5971);
and U6084 (N_6084,N_5892,N_5887);
and U6085 (N_6085,N_5873,N_5806);
nor U6086 (N_6086,N_5805,N_5759);
xor U6087 (N_6087,N_5893,N_5792);
and U6088 (N_6088,N_5937,N_5996);
nor U6089 (N_6089,N_5856,N_5854);
nand U6090 (N_6090,N_5993,N_5899);
nand U6091 (N_6091,N_5809,N_5968);
nand U6092 (N_6092,N_5991,N_5967);
xor U6093 (N_6093,N_5970,N_5973);
xor U6094 (N_6094,N_5837,N_5940);
nor U6095 (N_6095,N_5819,N_5879);
nand U6096 (N_6096,N_5782,N_5803);
or U6097 (N_6097,N_5790,N_5934);
nor U6098 (N_6098,N_5869,N_5896);
nand U6099 (N_6099,N_5762,N_5801);
and U6100 (N_6100,N_5988,N_5929);
or U6101 (N_6101,N_5880,N_5772);
nor U6102 (N_6102,N_5818,N_5778);
nor U6103 (N_6103,N_5835,N_5997);
nor U6104 (N_6104,N_5987,N_5947);
nand U6105 (N_6105,N_5822,N_5989);
nand U6106 (N_6106,N_5843,N_5865);
or U6107 (N_6107,N_5980,N_5836);
nand U6108 (N_6108,N_5999,N_5839);
or U6109 (N_6109,N_5963,N_5771);
or U6110 (N_6110,N_5758,N_5810);
or U6111 (N_6111,N_5918,N_5944);
or U6112 (N_6112,N_5894,N_5955);
nand U6113 (N_6113,N_5939,N_5964);
and U6114 (N_6114,N_5942,N_5871);
nor U6115 (N_6115,N_5845,N_5998);
nand U6116 (N_6116,N_5941,N_5863);
or U6117 (N_6117,N_5922,N_5957);
and U6118 (N_6118,N_5851,N_5938);
and U6119 (N_6119,N_5953,N_5901);
and U6120 (N_6120,N_5907,N_5972);
nor U6121 (N_6121,N_5876,N_5756);
nor U6122 (N_6122,N_5796,N_5920);
nor U6123 (N_6123,N_5961,N_5870);
xor U6124 (N_6124,N_5831,N_5779);
and U6125 (N_6125,N_5953,N_5969);
and U6126 (N_6126,N_5891,N_5780);
and U6127 (N_6127,N_5773,N_5849);
and U6128 (N_6128,N_5840,N_5937);
or U6129 (N_6129,N_5845,N_5944);
or U6130 (N_6130,N_5876,N_5939);
xor U6131 (N_6131,N_5858,N_5829);
xor U6132 (N_6132,N_5994,N_5795);
or U6133 (N_6133,N_5872,N_5813);
xor U6134 (N_6134,N_5874,N_5915);
and U6135 (N_6135,N_5963,N_5947);
nand U6136 (N_6136,N_5990,N_5875);
nand U6137 (N_6137,N_5979,N_5856);
xor U6138 (N_6138,N_5954,N_5959);
or U6139 (N_6139,N_5943,N_5879);
or U6140 (N_6140,N_5819,N_5921);
xor U6141 (N_6141,N_5813,N_5992);
xor U6142 (N_6142,N_5927,N_5849);
and U6143 (N_6143,N_5964,N_5924);
and U6144 (N_6144,N_5751,N_5868);
and U6145 (N_6145,N_5949,N_5832);
nor U6146 (N_6146,N_5815,N_5979);
nand U6147 (N_6147,N_5752,N_5908);
xnor U6148 (N_6148,N_5970,N_5760);
or U6149 (N_6149,N_5907,N_5758);
xor U6150 (N_6150,N_5818,N_5905);
and U6151 (N_6151,N_5775,N_5968);
nor U6152 (N_6152,N_5909,N_5816);
nand U6153 (N_6153,N_5793,N_5914);
and U6154 (N_6154,N_5844,N_5972);
and U6155 (N_6155,N_5941,N_5998);
and U6156 (N_6156,N_5900,N_5860);
nand U6157 (N_6157,N_5913,N_5946);
and U6158 (N_6158,N_5908,N_5813);
xor U6159 (N_6159,N_5774,N_5975);
or U6160 (N_6160,N_5782,N_5972);
or U6161 (N_6161,N_5922,N_5988);
and U6162 (N_6162,N_5862,N_5913);
nor U6163 (N_6163,N_5985,N_5958);
nand U6164 (N_6164,N_5940,N_5916);
or U6165 (N_6165,N_5989,N_5985);
and U6166 (N_6166,N_5752,N_5961);
xor U6167 (N_6167,N_5818,N_5886);
nand U6168 (N_6168,N_5887,N_5779);
nand U6169 (N_6169,N_5797,N_5931);
xnor U6170 (N_6170,N_5959,N_5872);
nand U6171 (N_6171,N_5789,N_5885);
nand U6172 (N_6172,N_5970,N_5840);
nor U6173 (N_6173,N_5964,N_5815);
nand U6174 (N_6174,N_5796,N_5989);
nor U6175 (N_6175,N_5821,N_5868);
or U6176 (N_6176,N_5898,N_5930);
nand U6177 (N_6177,N_5876,N_5888);
or U6178 (N_6178,N_5953,N_5897);
or U6179 (N_6179,N_5842,N_5920);
nand U6180 (N_6180,N_5818,N_5947);
or U6181 (N_6181,N_5987,N_5931);
or U6182 (N_6182,N_5911,N_5839);
or U6183 (N_6183,N_5950,N_5968);
nor U6184 (N_6184,N_5855,N_5794);
and U6185 (N_6185,N_5902,N_5861);
nand U6186 (N_6186,N_5882,N_5968);
nand U6187 (N_6187,N_5818,N_5851);
nor U6188 (N_6188,N_5849,N_5898);
or U6189 (N_6189,N_5939,N_5907);
xor U6190 (N_6190,N_5818,N_5917);
nor U6191 (N_6191,N_5820,N_5792);
or U6192 (N_6192,N_5900,N_5895);
nor U6193 (N_6193,N_5820,N_5863);
and U6194 (N_6194,N_5847,N_5843);
nand U6195 (N_6195,N_5954,N_5975);
and U6196 (N_6196,N_5835,N_5904);
and U6197 (N_6197,N_5819,N_5756);
nand U6198 (N_6198,N_5945,N_5904);
or U6199 (N_6199,N_5833,N_5889);
nor U6200 (N_6200,N_5812,N_5873);
and U6201 (N_6201,N_5904,N_5774);
nor U6202 (N_6202,N_5771,N_5758);
or U6203 (N_6203,N_5828,N_5945);
nor U6204 (N_6204,N_5916,N_5762);
nor U6205 (N_6205,N_5764,N_5793);
xnor U6206 (N_6206,N_5767,N_5830);
nand U6207 (N_6207,N_5958,N_5836);
nor U6208 (N_6208,N_5856,N_5944);
nor U6209 (N_6209,N_5772,N_5870);
or U6210 (N_6210,N_5935,N_5908);
and U6211 (N_6211,N_5947,N_5942);
nor U6212 (N_6212,N_5941,N_5861);
nor U6213 (N_6213,N_5977,N_5980);
nand U6214 (N_6214,N_5830,N_5833);
nor U6215 (N_6215,N_5837,N_5873);
xnor U6216 (N_6216,N_5806,N_5957);
and U6217 (N_6217,N_5900,N_5924);
or U6218 (N_6218,N_5752,N_5854);
nand U6219 (N_6219,N_5776,N_5946);
and U6220 (N_6220,N_5937,N_5960);
xor U6221 (N_6221,N_5855,N_5826);
nand U6222 (N_6222,N_5912,N_5781);
or U6223 (N_6223,N_5964,N_5954);
nor U6224 (N_6224,N_5958,N_5946);
nor U6225 (N_6225,N_5752,N_5801);
or U6226 (N_6226,N_5926,N_5879);
and U6227 (N_6227,N_5946,N_5885);
nand U6228 (N_6228,N_5881,N_5800);
nand U6229 (N_6229,N_5757,N_5890);
xnor U6230 (N_6230,N_5896,N_5856);
nand U6231 (N_6231,N_5947,N_5953);
and U6232 (N_6232,N_5964,N_5966);
nor U6233 (N_6233,N_5794,N_5795);
and U6234 (N_6234,N_5806,N_5790);
or U6235 (N_6235,N_5839,N_5866);
nor U6236 (N_6236,N_5901,N_5791);
nor U6237 (N_6237,N_5913,N_5853);
nor U6238 (N_6238,N_5930,N_5796);
and U6239 (N_6239,N_5793,N_5861);
nor U6240 (N_6240,N_5800,N_5887);
or U6241 (N_6241,N_5981,N_5795);
or U6242 (N_6242,N_5843,N_5863);
nor U6243 (N_6243,N_5775,N_5806);
nor U6244 (N_6244,N_5984,N_5968);
nor U6245 (N_6245,N_5942,N_5882);
and U6246 (N_6246,N_5773,N_5862);
nor U6247 (N_6247,N_5752,N_5764);
or U6248 (N_6248,N_5808,N_5792);
and U6249 (N_6249,N_5759,N_5844);
and U6250 (N_6250,N_6110,N_6097);
and U6251 (N_6251,N_6079,N_6232);
or U6252 (N_6252,N_6026,N_6021);
nand U6253 (N_6253,N_6249,N_6091);
or U6254 (N_6254,N_6235,N_6187);
and U6255 (N_6255,N_6063,N_6158);
nand U6256 (N_6256,N_6139,N_6014);
or U6257 (N_6257,N_6041,N_6210);
xor U6258 (N_6258,N_6118,N_6189);
nand U6259 (N_6259,N_6105,N_6168);
nor U6260 (N_6260,N_6046,N_6141);
and U6261 (N_6261,N_6180,N_6129);
nor U6262 (N_6262,N_6179,N_6221);
nand U6263 (N_6263,N_6003,N_6149);
nor U6264 (N_6264,N_6108,N_6011);
and U6265 (N_6265,N_6178,N_6215);
xnor U6266 (N_6266,N_6166,N_6220);
and U6267 (N_6267,N_6237,N_6174);
xnor U6268 (N_6268,N_6078,N_6100);
nand U6269 (N_6269,N_6009,N_6085);
and U6270 (N_6270,N_6116,N_6126);
and U6271 (N_6271,N_6121,N_6095);
nor U6272 (N_6272,N_6114,N_6099);
nor U6273 (N_6273,N_6130,N_6045);
nand U6274 (N_6274,N_6172,N_6248);
nand U6275 (N_6275,N_6096,N_6144);
and U6276 (N_6276,N_6173,N_6195);
or U6277 (N_6277,N_6194,N_6142);
and U6278 (N_6278,N_6034,N_6208);
or U6279 (N_6279,N_6247,N_6070);
xnor U6280 (N_6280,N_6150,N_6015);
nor U6281 (N_6281,N_6036,N_6084);
nor U6282 (N_6282,N_6153,N_6010);
nor U6283 (N_6283,N_6048,N_6101);
or U6284 (N_6284,N_6081,N_6002);
nor U6285 (N_6285,N_6224,N_6109);
nand U6286 (N_6286,N_6171,N_6062);
xor U6287 (N_6287,N_6028,N_6090);
nand U6288 (N_6288,N_6127,N_6152);
nand U6289 (N_6289,N_6004,N_6064);
and U6290 (N_6290,N_6234,N_6076);
xnor U6291 (N_6291,N_6124,N_6163);
nor U6292 (N_6292,N_6056,N_6103);
and U6293 (N_6293,N_6112,N_6167);
nand U6294 (N_6294,N_6106,N_6191);
or U6295 (N_6295,N_6136,N_6007);
and U6296 (N_6296,N_6077,N_6098);
nor U6297 (N_6297,N_6151,N_6053);
or U6298 (N_6298,N_6117,N_6212);
or U6299 (N_6299,N_6027,N_6154);
nand U6300 (N_6300,N_6082,N_6029);
or U6301 (N_6301,N_6075,N_6033);
nand U6302 (N_6302,N_6190,N_6175);
xor U6303 (N_6303,N_6155,N_6233);
and U6304 (N_6304,N_6209,N_6199);
xor U6305 (N_6305,N_6006,N_6069);
nor U6306 (N_6306,N_6111,N_6023);
nor U6307 (N_6307,N_6193,N_6217);
nand U6308 (N_6308,N_6134,N_6222);
or U6309 (N_6309,N_6071,N_6065);
and U6310 (N_6310,N_6185,N_6032);
or U6311 (N_6311,N_6223,N_6244);
nor U6312 (N_6312,N_6113,N_6022);
nor U6313 (N_6313,N_6120,N_6211);
or U6314 (N_6314,N_6236,N_6164);
or U6315 (N_6315,N_6005,N_6241);
nand U6316 (N_6316,N_6133,N_6092);
and U6317 (N_6317,N_6083,N_6102);
and U6318 (N_6318,N_6119,N_6128);
nand U6319 (N_6319,N_6072,N_6165);
nor U6320 (N_6320,N_6067,N_6156);
and U6321 (N_6321,N_6214,N_6051);
nor U6322 (N_6322,N_6170,N_6205);
xor U6323 (N_6323,N_6049,N_6184);
nand U6324 (N_6324,N_6186,N_6219);
or U6325 (N_6325,N_6054,N_6135);
nand U6326 (N_6326,N_6104,N_6204);
nand U6327 (N_6327,N_6012,N_6239);
and U6328 (N_6328,N_6226,N_6035);
and U6329 (N_6329,N_6008,N_6231);
or U6330 (N_6330,N_6060,N_6227);
nand U6331 (N_6331,N_6086,N_6203);
nor U6332 (N_6332,N_6225,N_6157);
and U6333 (N_6333,N_6196,N_6125);
and U6334 (N_6334,N_6206,N_6183);
nand U6335 (N_6335,N_6242,N_6115);
nand U6336 (N_6336,N_6019,N_6093);
and U6337 (N_6337,N_6137,N_6200);
or U6338 (N_6338,N_6073,N_6031);
xor U6339 (N_6339,N_6030,N_6016);
or U6340 (N_6340,N_6087,N_6162);
nor U6341 (N_6341,N_6228,N_6243);
and U6342 (N_6342,N_6143,N_6055);
or U6343 (N_6343,N_6122,N_6024);
nor U6344 (N_6344,N_6001,N_6013);
nand U6345 (N_6345,N_6107,N_6043);
or U6346 (N_6346,N_6230,N_6198);
nand U6347 (N_6347,N_6068,N_6161);
nor U6348 (N_6348,N_6052,N_6039);
xnor U6349 (N_6349,N_6148,N_6025);
and U6350 (N_6350,N_6123,N_6182);
nand U6351 (N_6351,N_6201,N_6197);
nand U6352 (N_6352,N_6074,N_6037);
nand U6353 (N_6353,N_6066,N_6042);
and U6354 (N_6354,N_6020,N_6188);
or U6355 (N_6355,N_6050,N_6047);
nand U6356 (N_6356,N_6088,N_6192);
nor U6357 (N_6357,N_6017,N_6038);
nand U6358 (N_6358,N_6044,N_6246);
or U6359 (N_6359,N_6058,N_6147);
nor U6360 (N_6360,N_6089,N_6213);
and U6361 (N_6361,N_6059,N_6040);
nand U6362 (N_6362,N_6216,N_6061);
or U6363 (N_6363,N_6202,N_6132);
or U6364 (N_6364,N_6146,N_6140);
nor U6365 (N_6365,N_6218,N_6094);
xnor U6366 (N_6366,N_6160,N_6176);
xor U6367 (N_6367,N_6080,N_6229);
xor U6368 (N_6368,N_6057,N_6131);
nand U6369 (N_6369,N_6181,N_6238);
nand U6370 (N_6370,N_6177,N_6245);
and U6371 (N_6371,N_6207,N_6018);
or U6372 (N_6372,N_6138,N_6169);
or U6373 (N_6373,N_6240,N_6145);
or U6374 (N_6374,N_6159,N_6000);
and U6375 (N_6375,N_6008,N_6101);
nor U6376 (N_6376,N_6151,N_6223);
or U6377 (N_6377,N_6183,N_6243);
nor U6378 (N_6378,N_6221,N_6021);
or U6379 (N_6379,N_6143,N_6244);
nand U6380 (N_6380,N_6128,N_6056);
or U6381 (N_6381,N_6016,N_6237);
xor U6382 (N_6382,N_6042,N_6192);
and U6383 (N_6383,N_6122,N_6007);
or U6384 (N_6384,N_6173,N_6087);
or U6385 (N_6385,N_6031,N_6048);
and U6386 (N_6386,N_6001,N_6133);
or U6387 (N_6387,N_6125,N_6157);
nor U6388 (N_6388,N_6056,N_6085);
xor U6389 (N_6389,N_6158,N_6177);
xor U6390 (N_6390,N_6241,N_6242);
nor U6391 (N_6391,N_6138,N_6185);
nand U6392 (N_6392,N_6172,N_6030);
xnor U6393 (N_6393,N_6214,N_6129);
nand U6394 (N_6394,N_6097,N_6154);
nand U6395 (N_6395,N_6062,N_6048);
nor U6396 (N_6396,N_6216,N_6031);
xor U6397 (N_6397,N_6053,N_6059);
xnor U6398 (N_6398,N_6017,N_6099);
xor U6399 (N_6399,N_6064,N_6212);
and U6400 (N_6400,N_6209,N_6091);
nor U6401 (N_6401,N_6171,N_6142);
nand U6402 (N_6402,N_6212,N_6239);
nor U6403 (N_6403,N_6002,N_6211);
or U6404 (N_6404,N_6153,N_6126);
or U6405 (N_6405,N_6240,N_6065);
nor U6406 (N_6406,N_6068,N_6105);
nor U6407 (N_6407,N_6202,N_6088);
or U6408 (N_6408,N_6060,N_6012);
nand U6409 (N_6409,N_6047,N_6120);
or U6410 (N_6410,N_6053,N_6139);
and U6411 (N_6411,N_6213,N_6074);
nor U6412 (N_6412,N_6219,N_6079);
nor U6413 (N_6413,N_6121,N_6005);
and U6414 (N_6414,N_6143,N_6187);
nor U6415 (N_6415,N_6217,N_6168);
nor U6416 (N_6416,N_6105,N_6023);
and U6417 (N_6417,N_6035,N_6149);
xor U6418 (N_6418,N_6204,N_6110);
or U6419 (N_6419,N_6222,N_6168);
nor U6420 (N_6420,N_6026,N_6192);
xor U6421 (N_6421,N_6196,N_6245);
nor U6422 (N_6422,N_6114,N_6023);
nor U6423 (N_6423,N_6222,N_6105);
nand U6424 (N_6424,N_6118,N_6073);
or U6425 (N_6425,N_6055,N_6002);
and U6426 (N_6426,N_6055,N_6024);
nor U6427 (N_6427,N_6056,N_6072);
or U6428 (N_6428,N_6196,N_6229);
and U6429 (N_6429,N_6008,N_6074);
and U6430 (N_6430,N_6237,N_6017);
nor U6431 (N_6431,N_6026,N_6077);
and U6432 (N_6432,N_6174,N_6120);
and U6433 (N_6433,N_6009,N_6237);
xor U6434 (N_6434,N_6002,N_6098);
nand U6435 (N_6435,N_6248,N_6083);
and U6436 (N_6436,N_6177,N_6204);
and U6437 (N_6437,N_6198,N_6022);
nor U6438 (N_6438,N_6122,N_6012);
nor U6439 (N_6439,N_6141,N_6120);
or U6440 (N_6440,N_6121,N_6068);
or U6441 (N_6441,N_6096,N_6066);
xnor U6442 (N_6442,N_6074,N_6221);
xor U6443 (N_6443,N_6200,N_6227);
and U6444 (N_6444,N_6111,N_6048);
and U6445 (N_6445,N_6157,N_6104);
and U6446 (N_6446,N_6220,N_6062);
or U6447 (N_6447,N_6162,N_6091);
nand U6448 (N_6448,N_6161,N_6160);
nand U6449 (N_6449,N_6137,N_6076);
and U6450 (N_6450,N_6181,N_6047);
and U6451 (N_6451,N_6126,N_6103);
nand U6452 (N_6452,N_6175,N_6102);
nor U6453 (N_6453,N_6188,N_6170);
or U6454 (N_6454,N_6235,N_6059);
nand U6455 (N_6455,N_6171,N_6117);
nor U6456 (N_6456,N_6239,N_6238);
xor U6457 (N_6457,N_6106,N_6090);
or U6458 (N_6458,N_6249,N_6085);
nand U6459 (N_6459,N_6152,N_6239);
nor U6460 (N_6460,N_6182,N_6111);
or U6461 (N_6461,N_6031,N_6083);
or U6462 (N_6462,N_6224,N_6071);
or U6463 (N_6463,N_6083,N_6233);
or U6464 (N_6464,N_6016,N_6120);
xor U6465 (N_6465,N_6248,N_6200);
xor U6466 (N_6466,N_6032,N_6125);
nand U6467 (N_6467,N_6203,N_6217);
or U6468 (N_6468,N_6022,N_6078);
nor U6469 (N_6469,N_6138,N_6172);
or U6470 (N_6470,N_6246,N_6249);
nand U6471 (N_6471,N_6074,N_6033);
and U6472 (N_6472,N_6179,N_6188);
nand U6473 (N_6473,N_6054,N_6031);
nand U6474 (N_6474,N_6031,N_6084);
and U6475 (N_6475,N_6221,N_6142);
and U6476 (N_6476,N_6091,N_6071);
nand U6477 (N_6477,N_6123,N_6038);
nand U6478 (N_6478,N_6149,N_6131);
or U6479 (N_6479,N_6122,N_6152);
or U6480 (N_6480,N_6027,N_6163);
nor U6481 (N_6481,N_6160,N_6207);
or U6482 (N_6482,N_6091,N_6140);
nor U6483 (N_6483,N_6095,N_6239);
nor U6484 (N_6484,N_6185,N_6037);
or U6485 (N_6485,N_6239,N_6101);
and U6486 (N_6486,N_6051,N_6090);
xor U6487 (N_6487,N_6196,N_6111);
nand U6488 (N_6488,N_6213,N_6073);
nor U6489 (N_6489,N_6163,N_6080);
nand U6490 (N_6490,N_6115,N_6248);
nor U6491 (N_6491,N_6152,N_6031);
nand U6492 (N_6492,N_6244,N_6128);
and U6493 (N_6493,N_6002,N_6008);
nand U6494 (N_6494,N_6239,N_6244);
nor U6495 (N_6495,N_6213,N_6162);
nor U6496 (N_6496,N_6228,N_6017);
nor U6497 (N_6497,N_6062,N_6144);
and U6498 (N_6498,N_6025,N_6090);
nand U6499 (N_6499,N_6127,N_6185);
or U6500 (N_6500,N_6306,N_6362);
and U6501 (N_6501,N_6370,N_6299);
nor U6502 (N_6502,N_6452,N_6406);
and U6503 (N_6503,N_6459,N_6250);
and U6504 (N_6504,N_6498,N_6387);
nand U6505 (N_6505,N_6258,N_6279);
and U6506 (N_6506,N_6453,N_6294);
nand U6507 (N_6507,N_6487,N_6397);
nor U6508 (N_6508,N_6348,N_6363);
nand U6509 (N_6509,N_6485,N_6484);
or U6510 (N_6510,N_6357,N_6347);
nand U6511 (N_6511,N_6263,N_6376);
nor U6512 (N_6512,N_6283,N_6403);
nand U6513 (N_6513,N_6417,N_6448);
and U6514 (N_6514,N_6367,N_6409);
or U6515 (N_6515,N_6284,N_6456);
nand U6516 (N_6516,N_6253,N_6385);
or U6517 (N_6517,N_6340,N_6424);
nor U6518 (N_6518,N_6413,N_6343);
and U6519 (N_6519,N_6301,N_6489);
nor U6520 (N_6520,N_6359,N_6255);
and U6521 (N_6521,N_6303,N_6304);
or U6522 (N_6522,N_6454,N_6445);
nor U6523 (N_6523,N_6261,N_6346);
nor U6524 (N_6524,N_6285,N_6432);
nor U6525 (N_6525,N_6429,N_6289);
and U6526 (N_6526,N_6380,N_6468);
nand U6527 (N_6527,N_6278,N_6313);
or U6528 (N_6528,N_6321,N_6420);
nand U6529 (N_6529,N_6441,N_6488);
and U6530 (N_6530,N_6312,N_6423);
nand U6531 (N_6531,N_6266,N_6422);
or U6532 (N_6532,N_6315,N_6439);
nor U6533 (N_6533,N_6349,N_6434);
and U6534 (N_6534,N_6351,N_6273);
or U6535 (N_6535,N_6355,N_6444);
nand U6536 (N_6536,N_6337,N_6476);
and U6537 (N_6537,N_6458,N_6341);
nand U6538 (N_6538,N_6475,N_6467);
and U6539 (N_6539,N_6461,N_6252);
and U6540 (N_6540,N_6316,N_6426);
nor U6541 (N_6541,N_6322,N_6386);
nand U6542 (N_6542,N_6272,N_6259);
nor U6543 (N_6543,N_6414,N_6265);
nor U6544 (N_6544,N_6494,N_6282);
nor U6545 (N_6545,N_6437,N_6449);
or U6546 (N_6546,N_6293,N_6411);
nand U6547 (N_6547,N_6329,N_6428);
nand U6548 (N_6548,N_6466,N_6412);
and U6549 (N_6549,N_6277,N_6395);
nor U6550 (N_6550,N_6275,N_6371);
nor U6551 (N_6551,N_6332,N_6495);
nor U6552 (N_6552,N_6496,N_6354);
or U6553 (N_6553,N_6281,N_6430);
or U6554 (N_6554,N_6374,N_6368);
or U6555 (N_6555,N_6296,N_6419);
nor U6556 (N_6556,N_6270,N_6269);
and U6557 (N_6557,N_6256,N_6460);
and U6558 (N_6558,N_6479,N_6440);
or U6559 (N_6559,N_6307,N_6431);
nand U6560 (N_6560,N_6251,N_6310);
nor U6561 (N_6561,N_6290,N_6470);
or U6562 (N_6562,N_6302,N_6398);
nand U6563 (N_6563,N_6268,N_6305);
or U6564 (N_6564,N_6342,N_6328);
nand U6565 (N_6565,N_6391,N_6309);
nor U6566 (N_6566,N_6350,N_6443);
nand U6567 (N_6567,N_6483,N_6474);
and U6568 (N_6568,N_6473,N_6369);
nand U6569 (N_6569,N_6325,N_6298);
nand U6570 (N_6570,N_6388,N_6384);
xnor U6571 (N_6571,N_6356,N_6469);
nand U6572 (N_6572,N_6421,N_6405);
nand U6573 (N_6573,N_6280,N_6499);
and U6574 (N_6574,N_6415,N_6338);
nor U6575 (N_6575,N_6271,N_6317);
and U6576 (N_6576,N_6292,N_6404);
nor U6577 (N_6577,N_6327,N_6345);
nand U6578 (N_6578,N_6274,N_6407);
and U6579 (N_6579,N_6442,N_6364);
and U6580 (N_6580,N_6465,N_6490);
nand U6581 (N_6581,N_6308,N_6288);
nand U6582 (N_6582,N_6254,N_6320);
and U6583 (N_6583,N_6333,N_6326);
or U6584 (N_6584,N_6295,N_6318);
and U6585 (N_6585,N_6464,N_6323);
nor U6586 (N_6586,N_6471,N_6377);
and U6587 (N_6587,N_6389,N_6447);
or U6588 (N_6588,N_6393,N_6383);
and U6589 (N_6589,N_6335,N_6416);
xor U6590 (N_6590,N_6390,N_6446);
nor U6591 (N_6591,N_6334,N_6433);
xor U6592 (N_6592,N_6478,N_6372);
nor U6593 (N_6593,N_6497,N_6400);
nor U6594 (N_6594,N_6291,N_6378);
or U6595 (N_6595,N_6396,N_6300);
and U6596 (N_6596,N_6286,N_6330);
and U6597 (N_6597,N_6392,N_6365);
nand U6598 (N_6598,N_6360,N_6438);
or U6599 (N_6599,N_6491,N_6314);
xor U6600 (N_6600,N_6492,N_6477);
nand U6601 (N_6601,N_6493,N_6480);
and U6602 (N_6602,N_6379,N_6319);
or U6603 (N_6603,N_6399,N_6336);
nor U6604 (N_6604,N_6463,N_6276);
nor U6605 (N_6605,N_6435,N_6451);
nand U6606 (N_6606,N_6401,N_6481);
nand U6607 (N_6607,N_6450,N_6455);
nor U6608 (N_6608,N_6353,N_6486);
xor U6609 (N_6609,N_6311,N_6408);
nand U6610 (N_6610,N_6361,N_6457);
or U6611 (N_6611,N_6375,N_6287);
nor U6612 (N_6612,N_6260,N_6381);
and U6613 (N_6613,N_6482,N_6462);
nor U6614 (N_6614,N_6358,N_6324);
or U6615 (N_6615,N_6427,N_6297);
or U6616 (N_6616,N_6264,N_6402);
and U6617 (N_6617,N_6352,N_6425);
nand U6618 (N_6618,N_6373,N_6394);
and U6619 (N_6619,N_6366,N_6472);
nand U6620 (N_6620,N_6262,N_6257);
nor U6621 (N_6621,N_6267,N_6331);
nand U6622 (N_6622,N_6418,N_6410);
or U6623 (N_6623,N_6382,N_6436);
nor U6624 (N_6624,N_6339,N_6344);
or U6625 (N_6625,N_6489,N_6394);
and U6626 (N_6626,N_6426,N_6346);
or U6627 (N_6627,N_6447,N_6351);
and U6628 (N_6628,N_6282,N_6338);
nand U6629 (N_6629,N_6499,N_6477);
nor U6630 (N_6630,N_6367,N_6298);
or U6631 (N_6631,N_6469,N_6454);
xor U6632 (N_6632,N_6456,N_6328);
nand U6633 (N_6633,N_6255,N_6266);
xnor U6634 (N_6634,N_6435,N_6409);
nor U6635 (N_6635,N_6250,N_6357);
nor U6636 (N_6636,N_6475,N_6446);
nor U6637 (N_6637,N_6424,N_6441);
or U6638 (N_6638,N_6427,N_6479);
or U6639 (N_6639,N_6445,N_6317);
and U6640 (N_6640,N_6304,N_6391);
or U6641 (N_6641,N_6449,N_6495);
and U6642 (N_6642,N_6426,N_6435);
or U6643 (N_6643,N_6368,N_6469);
and U6644 (N_6644,N_6385,N_6428);
or U6645 (N_6645,N_6357,N_6495);
or U6646 (N_6646,N_6397,N_6323);
and U6647 (N_6647,N_6444,N_6283);
or U6648 (N_6648,N_6265,N_6402);
nand U6649 (N_6649,N_6357,N_6471);
xnor U6650 (N_6650,N_6473,N_6379);
and U6651 (N_6651,N_6308,N_6409);
nand U6652 (N_6652,N_6438,N_6488);
nor U6653 (N_6653,N_6389,N_6326);
nor U6654 (N_6654,N_6469,N_6384);
and U6655 (N_6655,N_6276,N_6391);
nor U6656 (N_6656,N_6322,N_6308);
or U6657 (N_6657,N_6486,N_6448);
xor U6658 (N_6658,N_6278,N_6298);
nor U6659 (N_6659,N_6384,N_6250);
and U6660 (N_6660,N_6408,N_6353);
nor U6661 (N_6661,N_6294,N_6258);
and U6662 (N_6662,N_6471,N_6290);
and U6663 (N_6663,N_6277,N_6402);
nor U6664 (N_6664,N_6329,N_6277);
nor U6665 (N_6665,N_6259,N_6403);
nand U6666 (N_6666,N_6356,N_6323);
nand U6667 (N_6667,N_6292,N_6303);
nand U6668 (N_6668,N_6272,N_6347);
nand U6669 (N_6669,N_6259,N_6278);
xor U6670 (N_6670,N_6425,N_6281);
or U6671 (N_6671,N_6278,N_6459);
or U6672 (N_6672,N_6377,N_6302);
nand U6673 (N_6673,N_6399,N_6461);
or U6674 (N_6674,N_6263,N_6256);
nand U6675 (N_6675,N_6455,N_6382);
and U6676 (N_6676,N_6447,N_6470);
nand U6677 (N_6677,N_6308,N_6417);
nand U6678 (N_6678,N_6321,N_6252);
nor U6679 (N_6679,N_6433,N_6308);
or U6680 (N_6680,N_6451,N_6457);
or U6681 (N_6681,N_6496,N_6492);
nand U6682 (N_6682,N_6288,N_6448);
nand U6683 (N_6683,N_6275,N_6304);
and U6684 (N_6684,N_6410,N_6433);
or U6685 (N_6685,N_6327,N_6488);
or U6686 (N_6686,N_6381,N_6268);
and U6687 (N_6687,N_6395,N_6318);
nand U6688 (N_6688,N_6499,N_6354);
nand U6689 (N_6689,N_6312,N_6370);
nand U6690 (N_6690,N_6353,N_6318);
nor U6691 (N_6691,N_6460,N_6357);
nand U6692 (N_6692,N_6456,N_6318);
nor U6693 (N_6693,N_6424,N_6325);
or U6694 (N_6694,N_6349,N_6383);
nor U6695 (N_6695,N_6414,N_6493);
or U6696 (N_6696,N_6407,N_6474);
and U6697 (N_6697,N_6267,N_6290);
and U6698 (N_6698,N_6289,N_6300);
nand U6699 (N_6699,N_6330,N_6452);
nor U6700 (N_6700,N_6295,N_6342);
or U6701 (N_6701,N_6472,N_6263);
nand U6702 (N_6702,N_6298,N_6442);
nand U6703 (N_6703,N_6323,N_6360);
nor U6704 (N_6704,N_6459,N_6336);
nor U6705 (N_6705,N_6250,N_6484);
nor U6706 (N_6706,N_6482,N_6347);
nand U6707 (N_6707,N_6449,N_6277);
xnor U6708 (N_6708,N_6258,N_6374);
nor U6709 (N_6709,N_6349,N_6312);
or U6710 (N_6710,N_6430,N_6254);
nand U6711 (N_6711,N_6285,N_6359);
nand U6712 (N_6712,N_6263,N_6441);
nand U6713 (N_6713,N_6253,N_6430);
nand U6714 (N_6714,N_6256,N_6366);
and U6715 (N_6715,N_6423,N_6251);
or U6716 (N_6716,N_6345,N_6442);
nor U6717 (N_6717,N_6309,N_6399);
xnor U6718 (N_6718,N_6383,N_6468);
nand U6719 (N_6719,N_6464,N_6368);
or U6720 (N_6720,N_6404,N_6473);
or U6721 (N_6721,N_6429,N_6277);
xor U6722 (N_6722,N_6372,N_6256);
nor U6723 (N_6723,N_6395,N_6414);
xor U6724 (N_6724,N_6445,N_6334);
or U6725 (N_6725,N_6463,N_6329);
and U6726 (N_6726,N_6267,N_6411);
and U6727 (N_6727,N_6311,N_6438);
and U6728 (N_6728,N_6260,N_6306);
and U6729 (N_6729,N_6278,N_6370);
nor U6730 (N_6730,N_6298,N_6263);
and U6731 (N_6731,N_6373,N_6291);
or U6732 (N_6732,N_6302,N_6308);
and U6733 (N_6733,N_6460,N_6391);
nor U6734 (N_6734,N_6361,N_6355);
and U6735 (N_6735,N_6489,N_6373);
nand U6736 (N_6736,N_6412,N_6338);
nand U6737 (N_6737,N_6456,N_6435);
or U6738 (N_6738,N_6283,N_6309);
or U6739 (N_6739,N_6445,N_6473);
nor U6740 (N_6740,N_6449,N_6374);
or U6741 (N_6741,N_6390,N_6261);
or U6742 (N_6742,N_6275,N_6341);
nand U6743 (N_6743,N_6340,N_6441);
nor U6744 (N_6744,N_6382,N_6292);
nand U6745 (N_6745,N_6333,N_6361);
or U6746 (N_6746,N_6369,N_6301);
or U6747 (N_6747,N_6251,N_6439);
xor U6748 (N_6748,N_6467,N_6358);
nand U6749 (N_6749,N_6297,N_6424);
and U6750 (N_6750,N_6594,N_6505);
or U6751 (N_6751,N_6542,N_6668);
or U6752 (N_6752,N_6699,N_6558);
nand U6753 (N_6753,N_6693,N_6595);
and U6754 (N_6754,N_6695,N_6718);
nor U6755 (N_6755,N_6611,N_6539);
or U6756 (N_6756,N_6662,N_6655);
or U6757 (N_6757,N_6717,N_6538);
or U6758 (N_6758,N_6522,N_6688);
nand U6759 (N_6759,N_6553,N_6567);
and U6760 (N_6760,N_6703,N_6544);
nand U6761 (N_6761,N_6577,N_6515);
and U6762 (N_6762,N_6689,N_6554);
nor U6763 (N_6763,N_6716,N_6527);
or U6764 (N_6764,N_6671,N_6720);
nand U6765 (N_6765,N_6518,N_6678);
nor U6766 (N_6766,N_6534,N_6549);
and U6767 (N_6767,N_6593,N_6541);
nand U6768 (N_6768,N_6510,N_6643);
or U6769 (N_6769,N_6691,N_6574);
xor U6770 (N_6770,N_6630,N_6638);
or U6771 (N_6771,N_6686,N_6513);
xor U6772 (N_6772,N_6627,N_6568);
or U6773 (N_6773,N_6559,N_6632);
and U6774 (N_6774,N_6569,N_6673);
nand U6775 (N_6775,N_6620,N_6670);
and U6776 (N_6776,N_6659,N_6636);
nand U6777 (N_6777,N_6587,N_6552);
or U6778 (N_6778,N_6692,N_6625);
nand U6779 (N_6779,N_6713,N_6645);
nand U6780 (N_6780,N_6555,N_6584);
nand U6781 (N_6781,N_6640,N_6649);
nor U6782 (N_6782,N_6712,N_6633);
or U6783 (N_6783,N_6747,N_6672);
nand U6784 (N_6784,N_6580,N_6631);
or U6785 (N_6785,N_6512,N_6591);
and U6786 (N_6786,N_6579,N_6637);
nand U6787 (N_6787,N_6621,N_6709);
nor U6788 (N_6788,N_6602,N_6606);
nor U6789 (N_6789,N_6677,N_6694);
nand U6790 (N_6790,N_6743,N_6700);
xnor U6791 (N_6791,N_6710,N_6573);
xor U6792 (N_6792,N_6502,N_6592);
or U6793 (N_6793,N_6639,N_6521);
nor U6794 (N_6794,N_6701,N_6546);
nor U6795 (N_6795,N_6628,N_6690);
nand U6796 (N_6796,N_6605,N_6723);
nand U6797 (N_6797,N_6617,N_6742);
and U6798 (N_6798,N_6660,N_6597);
nand U6799 (N_6799,N_6744,N_6599);
nor U6800 (N_6800,N_6545,N_6565);
nor U6801 (N_6801,N_6618,N_6547);
or U6802 (N_6802,N_6654,N_6681);
nor U6803 (N_6803,N_6726,N_6560);
nand U6804 (N_6804,N_6615,N_6529);
or U6805 (N_6805,N_6586,N_6504);
or U6806 (N_6806,N_6725,N_6629);
nand U6807 (N_6807,N_6731,N_6714);
and U6808 (N_6808,N_6642,N_6697);
and U6809 (N_6809,N_6607,N_6550);
and U6810 (N_6810,N_6740,N_6500);
or U6811 (N_6811,N_6508,N_6656);
or U6812 (N_6812,N_6501,N_6614);
nand U6813 (N_6813,N_6646,N_6582);
xnor U6814 (N_6814,N_6571,N_6590);
nand U6815 (N_6815,N_6526,N_6664);
xnor U6816 (N_6816,N_6531,N_6589);
nand U6817 (N_6817,N_6736,N_6674);
or U6818 (N_6818,N_6684,N_6746);
or U6819 (N_6819,N_6509,N_6657);
nand U6820 (N_6820,N_6634,N_6596);
xnor U6821 (N_6821,N_6506,N_6598);
xor U6822 (N_6822,N_6724,N_6514);
nor U6823 (N_6823,N_6685,N_6581);
nor U6824 (N_6824,N_6698,N_6610);
nor U6825 (N_6825,N_6696,N_6722);
nor U6826 (N_6826,N_6728,N_6738);
xnor U6827 (N_6827,N_6585,N_6663);
and U6828 (N_6828,N_6702,N_6612);
xor U6829 (N_6829,N_6708,N_6675);
or U6830 (N_6830,N_6564,N_6721);
nand U6831 (N_6831,N_6575,N_6706);
nand U6832 (N_6832,N_6519,N_6613);
nor U6833 (N_6833,N_6669,N_6661);
xor U6834 (N_6834,N_6648,N_6619);
and U6835 (N_6835,N_6665,N_6651);
nor U6836 (N_6836,N_6676,N_6540);
and U6837 (N_6837,N_6537,N_6601);
and U6838 (N_6838,N_6516,N_6563);
xor U6839 (N_6839,N_6556,N_6557);
nand U6840 (N_6840,N_6523,N_6745);
or U6841 (N_6841,N_6732,N_6707);
nor U6842 (N_6842,N_6525,N_6562);
or U6843 (N_6843,N_6623,N_6533);
nor U6844 (N_6844,N_6734,N_6737);
nand U6845 (N_6845,N_6524,N_6741);
nand U6846 (N_6846,N_6733,N_6626);
nand U6847 (N_6847,N_6566,N_6604);
or U6848 (N_6848,N_6729,N_6609);
nor U6849 (N_6849,N_6667,N_6551);
or U6850 (N_6850,N_6583,N_6719);
or U6851 (N_6851,N_6715,N_6588);
nor U6852 (N_6852,N_6624,N_6503);
or U6853 (N_6853,N_6517,N_6666);
or U6854 (N_6854,N_6616,N_6711);
nor U6855 (N_6855,N_6727,N_6680);
nor U6856 (N_6856,N_6730,N_6603);
or U6857 (N_6857,N_6687,N_6578);
nor U6858 (N_6858,N_6749,N_6570);
or U6859 (N_6859,N_6530,N_6644);
and U6860 (N_6860,N_6622,N_6528);
and U6861 (N_6861,N_6641,N_6507);
and U6862 (N_6862,N_6650,N_6658);
and U6863 (N_6863,N_6548,N_6705);
nor U6864 (N_6864,N_6576,N_6532);
nand U6865 (N_6865,N_6561,N_6679);
or U6866 (N_6866,N_6572,N_6536);
nand U6867 (N_6867,N_6682,N_6535);
and U6868 (N_6868,N_6652,N_6683);
nor U6869 (N_6869,N_6608,N_6635);
nor U6870 (N_6870,N_6647,N_6520);
and U6871 (N_6871,N_6739,N_6748);
nand U6872 (N_6872,N_6735,N_6511);
nor U6873 (N_6873,N_6543,N_6600);
or U6874 (N_6874,N_6704,N_6653);
or U6875 (N_6875,N_6528,N_6612);
nand U6876 (N_6876,N_6716,N_6505);
nor U6877 (N_6877,N_6729,N_6680);
and U6878 (N_6878,N_6692,N_6551);
and U6879 (N_6879,N_6721,N_6749);
nor U6880 (N_6880,N_6529,N_6591);
nand U6881 (N_6881,N_6545,N_6503);
or U6882 (N_6882,N_6732,N_6596);
and U6883 (N_6883,N_6646,N_6624);
nand U6884 (N_6884,N_6599,N_6679);
and U6885 (N_6885,N_6612,N_6665);
and U6886 (N_6886,N_6619,N_6680);
and U6887 (N_6887,N_6679,N_6636);
or U6888 (N_6888,N_6564,N_6738);
nand U6889 (N_6889,N_6554,N_6633);
nand U6890 (N_6890,N_6648,N_6586);
nand U6891 (N_6891,N_6524,N_6681);
nand U6892 (N_6892,N_6518,N_6738);
nand U6893 (N_6893,N_6716,N_6745);
and U6894 (N_6894,N_6644,N_6559);
nor U6895 (N_6895,N_6524,N_6554);
xor U6896 (N_6896,N_6748,N_6628);
or U6897 (N_6897,N_6525,N_6565);
or U6898 (N_6898,N_6658,N_6519);
nor U6899 (N_6899,N_6503,N_6700);
and U6900 (N_6900,N_6732,N_6568);
and U6901 (N_6901,N_6566,N_6700);
nand U6902 (N_6902,N_6659,N_6734);
nand U6903 (N_6903,N_6655,N_6540);
nor U6904 (N_6904,N_6507,N_6525);
or U6905 (N_6905,N_6704,N_6712);
nor U6906 (N_6906,N_6628,N_6564);
and U6907 (N_6907,N_6651,N_6576);
nor U6908 (N_6908,N_6688,N_6749);
nor U6909 (N_6909,N_6599,N_6669);
and U6910 (N_6910,N_6523,N_6559);
nand U6911 (N_6911,N_6639,N_6652);
nand U6912 (N_6912,N_6601,N_6632);
and U6913 (N_6913,N_6661,N_6686);
or U6914 (N_6914,N_6688,N_6648);
and U6915 (N_6915,N_6602,N_6626);
and U6916 (N_6916,N_6553,N_6732);
nor U6917 (N_6917,N_6667,N_6633);
nand U6918 (N_6918,N_6660,N_6521);
and U6919 (N_6919,N_6520,N_6707);
xnor U6920 (N_6920,N_6749,N_6719);
or U6921 (N_6921,N_6598,N_6504);
nand U6922 (N_6922,N_6730,N_6578);
nor U6923 (N_6923,N_6567,N_6656);
or U6924 (N_6924,N_6526,N_6738);
xnor U6925 (N_6925,N_6586,N_6532);
nand U6926 (N_6926,N_6702,N_6749);
and U6927 (N_6927,N_6719,N_6697);
nor U6928 (N_6928,N_6729,N_6714);
nor U6929 (N_6929,N_6736,N_6543);
nor U6930 (N_6930,N_6672,N_6553);
or U6931 (N_6931,N_6627,N_6748);
and U6932 (N_6932,N_6632,N_6729);
nor U6933 (N_6933,N_6702,N_6624);
or U6934 (N_6934,N_6588,N_6604);
xor U6935 (N_6935,N_6659,N_6564);
nand U6936 (N_6936,N_6620,N_6588);
nor U6937 (N_6937,N_6551,N_6625);
or U6938 (N_6938,N_6738,N_6687);
and U6939 (N_6939,N_6723,N_6710);
nand U6940 (N_6940,N_6601,N_6597);
nand U6941 (N_6941,N_6666,N_6527);
nor U6942 (N_6942,N_6653,N_6587);
nor U6943 (N_6943,N_6721,N_6550);
nor U6944 (N_6944,N_6554,N_6574);
nand U6945 (N_6945,N_6501,N_6620);
or U6946 (N_6946,N_6622,N_6614);
nor U6947 (N_6947,N_6716,N_6568);
xor U6948 (N_6948,N_6696,N_6520);
and U6949 (N_6949,N_6522,N_6620);
nand U6950 (N_6950,N_6656,N_6742);
and U6951 (N_6951,N_6514,N_6744);
and U6952 (N_6952,N_6510,N_6673);
nand U6953 (N_6953,N_6643,N_6566);
xnor U6954 (N_6954,N_6682,N_6501);
nor U6955 (N_6955,N_6559,N_6534);
nand U6956 (N_6956,N_6743,N_6523);
and U6957 (N_6957,N_6619,N_6595);
nor U6958 (N_6958,N_6563,N_6622);
nor U6959 (N_6959,N_6524,N_6706);
and U6960 (N_6960,N_6622,N_6729);
xnor U6961 (N_6961,N_6582,N_6685);
or U6962 (N_6962,N_6683,N_6645);
nor U6963 (N_6963,N_6745,N_6656);
or U6964 (N_6964,N_6588,N_6601);
or U6965 (N_6965,N_6634,N_6748);
or U6966 (N_6966,N_6608,N_6559);
and U6967 (N_6967,N_6610,N_6585);
nand U6968 (N_6968,N_6720,N_6728);
nor U6969 (N_6969,N_6574,N_6662);
or U6970 (N_6970,N_6715,N_6719);
and U6971 (N_6971,N_6656,N_6601);
or U6972 (N_6972,N_6585,N_6578);
nor U6973 (N_6973,N_6501,N_6641);
xnor U6974 (N_6974,N_6678,N_6689);
and U6975 (N_6975,N_6599,N_6676);
or U6976 (N_6976,N_6628,N_6696);
or U6977 (N_6977,N_6605,N_6525);
and U6978 (N_6978,N_6683,N_6695);
and U6979 (N_6979,N_6524,N_6567);
nand U6980 (N_6980,N_6572,N_6645);
nand U6981 (N_6981,N_6653,N_6539);
or U6982 (N_6982,N_6726,N_6707);
xnor U6983 (N_6983,N_6584,N_6690);
nor U6984 (N_6984,N_6602,N_6652);
and U6985 (N_6985,N_6503,N_6593);
or U6986 (N_6986,N_6684,N_6717);
nand U6987 (N_6987,N_6636,N_6516);
nand U6988 (N_6988,N_6749,N_6634);
nand U6989 (N_6989,N_6611,N_6545);
nor U6990 (N_6990,N_6662,N_6625);
nor U6991 (N_6991,N_6537,N_6518);
or U6992 (N_6992,N_6710,N_6650);
or U6993 (N_6993,N_6554,N_6599);
nand U6994 (N_6994,N_6591,N_6587);
and U6995 (N_6995,N_6591,N_6603);
nand U6996 (N_6996,N_6537,N_6556);
nand U6997 (N_6997,N_6713,N_6555);
nor U6998 (N_6998,N_6622,N_6590);
and U6999 (N_6999,N_6520,N_6573);
and U7000 (N_7000,N_6993,N_6933);
nand U7001 (N_7001,N_6994,N_6967);
or U7002 (N_7002,N_6843,N_6830);
or U7003 (N_7003,N_6758,N_6823);
nand U7004 (N_7004,N_6948,N_6975);
nor U7005 (N_7005,N_6884,N_6792);
nand U7006 (N_7006,N_6803,N_6896);
and U7007 (N_7007,N_6946,N_6965);
and U7008 (N_7008,N_6928,N_6868);
nor U7009 (N_7009,N_6937,N_6772);
or U7010 (N_7010,N_6750,N_6938);
and U7011 (N_7011,N_6754,N_6809);
nand U7012 (N_7012,N_6811,N_6831);
or U7013 (N_7013,N_6777,N_6793);
or U7014 (N_7014,N_6880,N_6764);
nor U7015 (N_7015,N_6867,N_6922);
or U7016 (N_7016,N_6924,N_6852);
or U7017 (N_7017,N_6824,N_6783);
xnor U7018 (N_7018,N_6769,N_6818);
and U7019 (N_7019,N_6847,N_6888);
xor U7020 (N_7020,N_6945,N_6817);
nor U7021 (N_7021,N_6905,N_6807);
or U7022 (N_7022,N_6857,N_6826);
and U7023 (N_7023,N_6813,N_6804);
xor U7024 (N_7024,N_6976,N_6844);
nand U7025 (N_7025,N_6856,N_6907);
and U7026 (N_7026,N_6910,N_6909);
xor U7027 (N_7027,N_6768,N_6997);
nand U7028 (N_7028,N_6869,N_6902);
and U7029 (N_7029,N_6920,N_6927);
nand U7030 (N_7030,N_6865,N_6849);
nor U7031 (N_7031,N_6915,N_6767);
and U7032 (N_7032,N_6977,N_6969);
or U7033 (N_7033,N_6763,N_6986);
and U7034 (N_7034,N_6926,N_6753);
nand U7035 (N_7035,N_6752,N_6828);
nand U7036 (N_7036,N_6851,N_6987);
nand U7037 (N_7037,N_6776,N_6839);
nand U7038 (N_7038,N_6755,N_6981);
nand U7039 (N_7039,N_6874,N_6808);
nand U7040 (N_7040,N_6855,N_6913);
or U7041 (N_7041,N_6995,N_6858);
nand U7042 (N_7042,N_6952,N_6848);
nor U7043 (N_7043,N_6889,N_6791);
nor U7044 (N_7044,N_6918,N_6757);
nand U7045 (N_7045,N_6954,N_6797);
nor U7046 (N_7046,N_6985,N_6778);
nor U7047 (N_7047,N_6898,N_6935);
or U7048 (N_7048,N_6879,N_6980);
nand U7049 (N_7049,N_6883,N_6814);
nand U7050 (N_7050,N_6765,N_6882);
or U7051 (N_7051,N_6904,N_6881);
nand U7052 (N_7052,N_6988,N_6953);
nor U7053 (N_7053,N_6895,N_6825);
nor U7054 (N_7054,N_6766,N_6756);
nor U7055 (N_7055,N_6859,N_6875);
nor U7056 (N_7056,N_6822,N_6978);
nor U7057 (N_7057,N_6786,N_6914);
or U7058 (N_7058,N_6762,N_6770);
nand U7059 (N_7059,N_6829,N_6984);
and U7060 (N_7060,N_6827,N_6853);
and U7061 (N_7061,N_6890,N_6941);
and U7062 (N_7062,N_6983,N_6796);
or U7063 (N_7063,N_6960,N_6971);
and U7064 (N_7064,N_6932,N_6854);
and U7065 (N_7065,N_6943,N_6950);
nand U7066 (N_7066,N_6788,N_6892);
nand U7067 (N_7067,N_6801,N_6963);
xor U7068 (N_7068,N_6939,N_6784);
nor U7069 (N_7069,N_6957,N_6773);
xnor U7070 (N_7070,N_6841,N_6805);
or U7071 (N_7071,N_6958,N_6992);
nand U7072 (N_7072,N_6780,N_6897);
nand U7073 (N_7073,N_6774,N_6872);
or U7074 (N_7074,N_6850,N_6789);
nor U7075 (N_7075,N_6956,N_6876);
xor U7076 (N_7076,N_6942,N_6925);
nor U7077 (N_7077,N_6833,N_6917);
nand U7078 (N_7078,N_6919,N_6899);
nor U7079 (N_7079,N_6802,N_6800);
xnor U7080 (N_7080,N_6837,N_6834);
nand U7081 (N_7081,N_6842,N_6799);
or U7082 (N_7082,N_6761,N_6863);
nor U7083 (N_7083,N_6835,N_6785);
or U7084 (N_7084,N_6878,N_6947);
nand U7085 (N_7085,N_6934,N_6979);
nor U7086 (N_7086,N_6893,N_6944);
nor U7087 (N_7087,N_6832,N_6923);
nand U7088 (N_7088,N_6815,N_6996);
and U7089 (N_7089,N_6760,N_6860);
nor U7090 (N_7090,N_6759,N_6775);
and U7091 (N_7091,N_6877,N_6862);
nor U7092 (N_7092,N_6891,N_6887);
or U7093 (N_7093,N_6816,N_6794);
nor U7094 (N_7094,N_6840,N_6871);
nand U7095 (N_7095,N_6779,N_6921);
or U7096 (N_7096,N_6903,N_6991);
nand U7097 (N_7097,N_6886,N_6973);
nand U7098 (N_7098,N_6838,N_6955);
nand U7099 (N_7099,N_6836,N_6810);
nand U7100 (N_7100,N_6821,N_6970);
or U7101 (N_7101,N_6866,N_6845);
nor U7102 (N_7102,N_6787,N_6951);
nor U7103 (N_7103,N_6968,N_6820);
and U7104 (N_7104,N_6782,N_6795);
nand U7105 (N_7105,N_6930,N_6959);
or U7106 (N_7106,N_6790,N_6936);
nand U7107 (N_7107,N_6771,N_6806);
or U7108 (N_7108,N_6929,N_6900);
nand U7109 (N_7109,N_6812,N_6931);
or U7110 (N_7110,N_6974,N_6982);
nand U7111 (N_7111,N_6908,N_6990);
nand U7112 (N_7112,N_6906,N_6916);
nor U7113 (N_7113,N_6964,N_6846);
nor U7114 (N_7114,N_6894,N_6940);
and U7115 (N_7115,N_6873,N_6961);
or U7116 (N_7116,N_6751,N_6912);
nand U7117 (N_7117,N_6781,N_6870);
and U7118 (N_7118,N_6885,N_6962);
xnor U7119 (N_7119,N_6861,N_6901);
xnor U7120 (N_7120,N_6972,N_6999);
and U7121 (N_7121,N_6989,N_6819);
or U7122 (N_7122,N_6966,N_6949);
nor U7123 (N_7123,N_6864,N_6998);
and U7124 (N_7124,N_6798,N_6911);
and U7125 (N_7125,N_6855,N_6870);
and U7126 (N_7126,N_6987,N_6911);
or U7127 (N_7127,N_6961,N_6803);
and U7128 (N_7128,N_6907,N_6825);
or U7129 (N_7129,N_6839,N_6972);
and U7130 (N_7130,N_6911,N_6841);
xnor U7131 (N_7131,N_6985,N_6792);
or U7132 (N_7132,N_6811,N_6772);
or U7133 (N_7133,N_6887,N_6980);
nand U7134 (N_7134,N_6881,N_6800);
and U7135 (N_7135,N_6758,N_6825);
and U7136 (N_7136,N_6974,N_6843);
xor U7137 (N_7137,N_6787,N_6988);
nand U7138 (N_7138,N_6949,N_6753);
nor U7139 (N_7139,N_6878,N_6958);
nor U7140 (N_7140,N_6984,N_6933);
or U7141 (N_7141,N_6861,N_6773);
and U7142 (N_7142,N_6786,N_6960);
nand U7143 (N_7143,N_6951,N_6862);
or U7144 (N_7144,N_6982,N_6894);
and U7145 (N_7145,N_6972,N_6899);
or U7146 (N_7146,N_6954,N_6974);
nor U7147 (N_7147,N_6873,N_6953);
xor U7148 (N_7148,N_6878,N_6873);
and U7149 (N_7149,N_6954,N_6822);
and U7150 (N_7150,N_6783,N_6919);
and U7151 (N_7151,N_6784,N_6754);
nor U7152 (N_7152,N_6762,N_6996);
nand U7153 (N_7153,N_6874,N_6773);
or U7154 (N_7154,N_6828,N_6965);
or U7155 (N_7155,N_6942,N_6766);
nor U7156 (N_7156,N_6822,N_6923);
nand U7157 (N_7157,N_6770,N_6964);
nor U7158 (N_7158,N_6920,N_6962);
xnor U7159 (N_7159,N_6885,N_6947);
or U7160 (N_7160,N_6938,N_6796);
nor U7161 (N_7161,N_6980,N_6894);
or U7162 (N_7162,N_6777,N_6847);
xnor U7163 (N_7163,N_6917,N_6978);
or U7164 (N_7164,N_6792,N_6826);
nor U7165 (N_7165,N_6781,N_6984);
or U7166 (N_7166,N_6869,N_6753);
nor U7167 (N_7167,N_6932,N_6959);
and U7168 (N_7168,N_6912,N_6875);
and U7169 (N_7169,N_6931,N_6756);
xnor U7170 (N_7170,N_6994,N_6888);
and U7171 (N_7171,N_6937,N_6920);
or U7172 (N_7172,N_6994,N_6772);
nor U7173 (N_7173,N_6797,N_6768);
nor U7174 (N_7174,N_6991,N_6767);
or U7175 (N_7175,N_6881,N_6792);
nor U7176 (N_7176,N_6970,N_6936);
or U7177 (N_7177,N_6766,N_6879);
and U7178 (N_7178,N_6815,N_6781);
xor U7179 (N_7179,N_6922,N_6830);
xnor U7180 (N_7180,N_6919,N_6912);
xor U7181 (N_7181,N_6756,N_6966);
and U7182 (N_7182,N_6841,N_6996);
and U7183 (N_7183,N_6763,N_6804);
and U7184 (N_7184,N_6982,N_6869);
xor U7185 (N_7185,N_6921,N_6978);
nand U7186 (N_7186,N_6856,N_6951);
nor U7187 (N_7187,N_6843,N_6774);
xor U7188 (N_7188,N_6970,N_6778);
and U7189 (N_7189,N_6773,N_6867);
nand U7190 (N_7190,N_6970,N_6937);
or U7191 (N_7191,N_6862,N_6843);
xnor U7192 (N_7192,N_6840,N_6993);
nand U7193 (N_7193,N_6777,N_6901);
and U7194 (N_7194,N_6957,N_6781);
nor U7195 (N_7195,N_6977,N_6756);
or U7196 (N_7196,N_6840,N_6911);
and U7197 (N_7197,N_6894,N_6774);
nor U7198 (N_7198,N_6960,N_6907);
and U7199 (N_7199,N_6808,N_6864);
nand U7200 (N_7200,N_6898,N_6767);
and U7201 (N_7201,N_6901,N_6979);
and U7202 (N_7202,N_6909,N_6814);
nor U7203 (N_7203,N_6869,N_6862);
xor U7204 (N_7204,N_6959,N_6973);
and U7205 (N_7205,N_6991,N_6898);
and U7206 (N_7206,N_6995,N_6802);
and U7207 (N_7207,N_6834,N_6751);
nand U7208 (N_7208,N_6909,N_6802);
or U7209 (N_7209,N_6948,N_6898);
nand U7210 (N_7210,N_6840,N_6778);
and U7211 (N_7211,N_6995,N_6962);
xnor U7212 (N_7212,N_6831,N_6969);
xor U7213 (N_7213,N_6847,N_6939);
and U7214 (N_7214,N_6891,N_6759);
nor U7215 (N_7215,N_6768,N_6788);
nand U7216 (N_7216,N_6981,N_6907);
xor U7217 (N_7217,N_6854,N_6907);
nand U7218 (N_7218,N_6898,N_6846);
or U7219 (N_7219,N_6821,N_6869);
or U7220 (N_7220,N_6805,N_6970);
nand U7221 (N_7221,N_6864,N_6898);
nand U7222 (N_7222,N_6815,N_6777);
nor U7223 (N_7223,N_6782,N_6885);
and U7224 (N_7224,N_6832,N_6783);
nor U7225 (N_7225,N_6941,N_6755);
nand U7226 (N_7226,N_6770,N_6956);
or U7227 (N_7227,N_6845,N_6872);
nor U7228 (N_7228,N_6834,N_6881);
nand U7229 (N_7229,N_6926,N_6942);
nor U7230 (N_7230,N_6884,N_6997);
nor U7231 (N_7231,N_6936,N_6985);
nor U7232 (N_7232,N_6917,N_6949);
nor U7233 (N_7233,N_6865,N_6892);
and U7234 (N_7234,N_6760,N_6930);
nor U7235 (N_7235,N_6917,N_6887);
nor U7236 (N_7236,N_6880,N_6783);
or U7237 (N_7237,N_6952,N_6912);
xor U7238 (N_7238,N_6959,N_6811);
and U7239 (N_7239,N_6948,N_6976);
xor U7240 (N_7240,N_6799,N_6914);
nand U7241 (N_7241,N_6996,N_6777);
or U7242 (N_7242,N_6822,N_6973);
nand U7243 (N_7243,N_6861,N_6998);
or U7244 (N_7244,N_6947,N_6857);
xor U7245 (N_7245,N_6884,N_6949);
xor U7246 (N_7246,N_6862,N_6925);
and U7247 (N_7247,N_6837,N_6920);
nand U7248 (N_7248,N_6782,N_6870);
nand U7249 (N_7249,N_6908,N_6766);
nand U7250 (N_7250,N_7089,N_7214);
nand U7251 (N_7251,N_7084,N_7164);
or U7252 (N_7252,N_7226,N_7065);
nand U7253 (N_7253,N_7036,N_7098);
xor U7254 (N_7254,N_7026,N_7019);
nand U7255 (N_7255,N_7160,N_7027);
nor U7256 (N_7256,N_7095,N_7238);
and U7257 (N_7257,N_7047,N_7107);
and U7258 (N_7258,N_7112,N_7038);
and U7259 (N_7259,N_7063,N_7079);
and U7260 (N_7260,N_7074,N_7024);
and U7261 (N_7261,N_7087,N_7240);
or U7262 (N_7262,N_7099,N_7118);
or U7263 (N_7263,N_7013,N_7044);
nor U7264 (N_7264,N_7059,N_7202);
and U7265 (N_7265,N_7097,N_7188);
and U7266 (N_7266,N_7033,N_7200);
nand U7267 (N_7267,N_7113,N_7009);
xor U7268 (N_7268,N_7052,N_7022);
nor U7269 (N_7269,N_7078,N_7204);
and U7270 (N_7270,N_7073,N_7137);
or U7271 (N_7271,N_7215,N_7075);
or U7272 (N_7272,N_7191,N_7181);
or U7273 (N_7273,N_7001,N_7085);
and U7274 (N_7274,N_7157,N_7201);
and U7275 (N_7275,N_7172,N_7245);
nor U7276 (N_7276,N_7124,N_7244);
nor U7277 (N_7277,N_7125,N_7028);
or U7278 (N_7278,N_7086,N_7061);
and U7279 (N_7279,N_7042,N_7170);
and U7280 (N_7280,N_7173,N_7020);
and U7281 (N_7281,N_7011,N_7104);
nand U7282 (N_7282,N_7021,N_7071);
nand U7283 (N_7283,N_7187,N_7182);
or U7284 (N_7284,N_7093,N_7135);
nor U7285 (N_7285,N_7235,N_7212);
and U7286 (N_7286,N_7211,N_7183);
or U7287 (N_7287,N_7231,N_7106);
nor U7288 (N_7288,N_7133,N_7242);
or U7289 (N_7289,N_7067,N_7072);
or U7290 (N_7290,N_7195,N_7165);
nand U7291 (N_7291,N_7248,N_7102);
and U7292 (N_7292,N_7123,N_7139);
and U7293 (N_7293,N_7101,N_7145);
and U7294 (N_7294,N_7144,N_7234);
and U7295 (N_7295,N_7041,N_7008);
and U7296 (N_7296,N_7184,N_7229);
nand U7297 (N_7297,N_7247,N_7222);
nand U7298 (N_7298,N_7228,N_7227);
and U7299 (N_7299,N_7018,N_7151);
and U7300 (N_7300,N_7108,N_7005);
nand U7301 (N_7301,N_7025,N_7190);
or U7302 (N_7302,N_7080,N_7158);
and U7303 (N_7303,N_7014,N_7029);
nor U7304 (N_7304,N_7092,N_7109);
and U7305 (N_7305,N_7000,N_7010);
and U7306 (N_7306,N_7233,N_7006);
or U7307 (N_7307,N_7171,N_7091);
nand U7308 (N_7308,N_7031,N_7239);
and U7309 (N_7309,N_7069,N_7083);
nor U7310 (N_7310,N_7205,N_7115);
or U7311 (N_7311,N_7179,N_7128);
or U7312 (N_7312,N_7156,N_7210);
xor U7313 (N_7313,N_7166,N_7105);
or U7314 (N_7314,N_7155,N_7002);
and U7315 (N_7315,N_7185,N_7132);
xor U7316 (N_7316,N_7060,N_7230);
or U7317 (N_7317,N_7066,N_7237);
or U7318 (N_7318,N_7243,N_7142);
or U7319 (N_7319,N_7134,N_7152);
xor U7320 (N_7320,N_7121,N_7032);
nor U7321 (N_7321,N_7167,N_7154);
and U7322 (N_7322,N_7090,N_7189);
nand U7323 (N_7323,N_7081,N_7140);
or U7324 (N_7324,N_7051,N_7159);
or U7325 (N_7325,N_7034,N_7058);
nor U7326 (N_7326,N_7012,N_7241);
and U7327 (N_7327,N_7054,N_7209);
or U7328 (N_7328,N_7143,N_7117);
and U7329 (N_7329,N_7035,N_7088);
nand U7330 (N_7330,N_7126,N_7207);
xor U7331 (N_7331,N_7127,N_7203);
nor U7332 (N_7332,N_7039,N_7147);
and U7333 (N_7333,N_7040,N_7068);
nor U7334 (N_7334,N_7194,N_7153);
nand U7335 (N_7335,N_7208,N_7064);
nor U7336 (N_7336,N_7216,N_7129);
xnor U7337 (N_7337,N_7103,N_7221);
nand U7338 (N_7338,N_7070,N_7116);
or U7339 (N_7339,N_7053,N_7045);
or U7340 (N_7340,N_7178,N_7246);
nand U7341 (N_7341,N_7138,N_7219);
nor U7342 (N_7342,N_7136,N_7149);
and U7343 (N_7343,N_7023,N_7030);
or U7344 (N_7344,N_7094,N_7082);
and U7345 (N_7345,N_7146,N_7055);
nand U7346 (N_7346,N_7110,N_7003);
xnor U7347 (N_7347,N_7177,N_7223);
nand U7348 (N_7348,N_7225,N_7114);
nand U7349 (N_7349,N_7220,N_7206);
xor U7350 (N_7350,N_7192,N_7180);
or U7351 (N_7351,N_7048,N_7096);
and U7352 (N_7352,N_7249,N_7198);
and U7353 (N_7353,N_7122,N_7049);
nor U7354 (N_7354,N_7050,N_7213);
nand U7355 (N_7355,N_7186,N_7169);
or U7356 (N_7356,N_7176,N_7119);
xnor U7357 (N_7357,N_7196,N_7062);
xor U7358 (N_7358,N_7130,N_7163);
nor U7359 (N_7359,N_7161,N_7037);
and U7360 (N_7360,N_7056,N_7162);
nor U7361 (N_7361,N_7077,N_7004);
nor U7362 (N_7362,N_7232,N_7043);
nor U7363 (N_7363,N_7148,N_7046);
and U7364 (N_7364,N_7150,N_7193);
and U7365 (N_7365,N_7236,N_7015);
nand U7366 (N_7366,N_7217,N_7197);
or U7367 (N_7367,N_7168,N_7007);
and U7368 (N_7368,N_7100,N_7224);
nor U7369 (N_7369,N_7016,N_7076);
nor U7370 (N_7370,N_7131,N_7017);
and U7371 (N_7371,N_7199,N_7218);
nand U7372 (N_7372,N_7111,N_7174);
nor U7373 (N_7373,N_7141,N_7057);
and U7374 (N_7374,N_7175,N_7120);
xnor U7375 (N_7375,N_7006,N_7160);
nand U7376 (N_7376,N_7096,N_7129);
nand U7377 (N_7377,N_7014,N_7063);
nand U7378 (N_7378,N_7006,N_7214);
or U7379 (N_7379,N_7194,N_7112);
nand U7380 (N_7380,N_7127,N_7235);
nor U7381 (N_7381,N_7097,N_7145);
nand U7382 (N_7382,N_7174,N_7232);
and U7383 (N_7383,N_7232,N_7026);
and U7384 (N_7384,N_7238,N_7118);
and U7385 (N_7385,N_7187,N_7019);
or U7386 (N_7386,N_7041,N_7075);
nand U7387 (N_7387,N_7206,N_7037);
nor U7388 (N_7388,N_7149,N_7121);
xnor U7389 (N_7389,N_7079,N_7149);
and U7390 (N_7390,N_7234,N_7152);
and U7391 (N_7391,N_7003,N_7124);
nand U7392 (N_7392,N_7214,N_7174);
xor U7393 (N_7393,N_7152,N_7135);
and U7394 (N_7394,N_7095,N_7146);
nand U7395 (N_7395,N_7155,N_7129);
xnor U7396 (N_7396,N_7249,N_7052);
xnor U7397 (N_7397,N_7010,N_7026);
nand U7398 (N_7398,N_7072,N_7148);
nand U7399 (N_7399,N_7071,N_7234);
nand U7400 (N_7400,N_7069,N_7115);
or U7401 (N_7401,N_7175,N_7227);
and U7402 (N_7402,N_7014,N_7180);
xnor U7403 (N_7403,N_7155,N_7208);
nor U7404 (N_7404,N_7120,N_7173);
nor U7405 (N_7405,N_7028,N_7185);
nor U7406 (N_7406,N_7227,N_7187);
nand U7407 (N_7407,N_7243,N_7182);
or U7408 (N_7408,N_7249,N_7146);
or U7409 (N_7409,N_7056,N_7009);
or U7410 (N_7410,N_7226,N_7233);
nor U7411 (N_7411,N_7083,N_7164);
xor U7412 (N_7412,N_7189,N_7223);
xnor U7413 (N_7413,N_7172,N_7189);
and U7414 (N_7414,N_7030,N_7194);
nor U7415 (N_7415,N_7003,N_7018);
nor U7416 (N_7416,N_7120,N_7021);
nor U7417 (N_7417,N_7127,N_7100);
xnor U7418 (N_7418,N_7116,N_7012);
or U7419 (N_7419,N_7208,N_7179);
or U7420 (N_7420,N_7025,N_7213);
and U7421 (N_7421,N_7006,N_7074);
xor U7422 (N_7422,N_7023,N_7237);
nand U7423 (N_7423,N_7063,N_7242);
or U7424 (N_7424,N_7214,N_7093);
or U7425 (N_7425,N_7130,N_7155);
or U7426 (N_7426,N_7130,N_7178);
or U7427 (N_7427,N_7026,N_7234);
and U7428 (N_7428,N_7246,N_7182);
nand U7429 (N_7429,N_7081,N_7070);
and U7430 (N_7430,N_7032,N_7247);
xnor U7431 (N_7431,N_7239,N_7219);
nor U7432 (N_7432,N_7244,N_7133);
nand U7433 (N_7433,N_7036,N_7185);
nor U7434 (N_7434,N_7011,N_7123);
and U7435 (N_7435,N_7242,N_7209);
nor U7436 (N_7436,N_7163,N_7196);
nand U7437 (N_7437,N_7062,N_7187);
and U7438 (N_7438,N_7045,N_7036);
and U7439 (N_7439,N_7240,N_7011);
nand U7440 (N_7440,N_7138,N_7031);
nand U7441 (N_7441,N_7077,N_7117);
or U7442 (N_7442,N_7035,N_7162);
xnor U7443 (N_7443,N_7202,N_7143);
xnor U7444 (N_7444,N_7050,N_7109);
nand U7445 (N_7445,N_7069,N_7100);
nand U7446 (N_7446,N_7236,N_7059);
nor U7447 (N_7447,N_7110,N_7207);
and U7448 (N_7448,N_7156,N_7024);
nor U7449 (N_7449,N_7212,N_7088);
nor U7450 (N_7450,N_7217,N_7153);
and U7451 (N_7451,N_7246,N_7045);
nor U7452 (N_7452,N_7098,N_7055);
and U7453 (N_7453,N_7196,N_7035);
or U7454 (N_7454,N_7060,N_7104);
nand U7455 (N_7455,N_7193,N_7142);
nor U7456 (N_7456,N_7028,N_7134);
nand U7457 (N_7457,N_7185,N_7122);
and U7458 (N_7458,N_7095,N_7230);
or U7459 (N_7459,N_7176,N_7240);
xnor U7460 (N_7460,N_7238,N_7168);
or U7461 (N_7461,N_7020,N_7229);
and U7462 (N_7462,N_7193,N_7186);
or U7463 (N_7463,N_7121,N_7045);
and U7464 (N_7464,N_7072,N_7139);
or U7465 (N_7465,N_7180,N_7082);
nor U7466 (N_7466,N_7226,N_7244);
xnor U7467 (N_7467,N_7116,N_7026);
xor U7468 (N_7468,N_7158,N_7061);
nand U7469 (N_7469,N_7212,N_7103);
nor U7470 (N_7470,N_7127,N_7085);
nor U7471 (N_7471,N_7168,N_7239);
nand U7472 (N_7472,N_7077,N_7019);
xor U7473 (N_7473,N_7127,N_7036);
nor U7474 (N_7474,N_7142,N_7205);
or U7475 (N_7475,N_7241,N_7109);
xor U7476 (N_7476,N_7096,N_7204);
or U7477 (N_7477,N_7187,N_7032);
nor U7478 (N_7478,N_7033,N_7201);
nand U7479 (N_7479,N_7203,N_7094);
or U7480 (N_7480,N_7019,N_7005);
and U7481 (N_7481,N_7107,N_7128);
nor U7482 (N_7482,N_7206,N_7105);
or U7483 (N_7483,N_7131,N_7166);
or U7484 (N_7484,N_7154,N_7099);
and U7485 (N_7485,N_7244,N_7143);
nand U7486 (N_7486,N_7092,N_7203);
nand U7487 (N_7487,N_7157,N_7132);
nor U7488 (N_7488,N_7044,N_7153);
nor U7489 (N_7489,N_7009,N_7149);
or U7490 (N_7490,N_7199,N_7058);
nand U7491 (N_7491,N_7093,N_7181);
or U7492 (N_7492,N_7187,N_7063);
or U7493 (N_7493,N_7061,N_7125);
or U7494 (N_7494,N_7000,N_7074);
and U7495 (N_7495,N_7216,N_7243);
nand U7496 (N_7496,N_7065,N_7053);
or U7497 (N_7497,N_7092,N_7036);
nand U7498 (N_7498,N_7196,N_7142);
or U7499 (N_7499,N_7144,N_7202);
and U7500 (N_7500,N_7293,N_7437);
nand U7501 (N_7501,N_7332,N_7372);
or U7502 (N_7502,N_7459,N_7285);
and U7503 (N_7503,N_7493,N_7331);
xnor U7504 (N_7504,N_7328,N_7439);
and U7505 (N_7505,N_7391,N_7484);
and U7506 (N_7506,N_7485,N_7448);
xor U7507 (N_7507,N_7295,N_7317);
nor U7508 (N_7508,N_7438,N_7263);
or U7509 (N_7509,N_7407,N_7398);
nor U7510 (N_7510,N_7253,N_7307);
or U7511 (N_7511,N_7381,N_7472);
and U7512 (N_7512,N_7426,N_7498);
xor U7513 (N_7513,N_7443,N_7408);
or U7514 (N_7514,N_7402,N_7454);
nand U7515 (N_7515,N_7283,N_7475);
or U7516 (N_7516,N_7281,N_7414);
nor U7517 (N_7517,N_7250,N_7278);
nor U7518 (N_7518,N_7313,N_7464);
and U7519 (N_7519,N_7320,N_7302);
and U7520 (N_7520,N_7298,N_7413);
and U7521 (N_7521,N_7481,N_7259);
nand U7522 (N_7522,N_7455,N_7430);
nand U7523 (N_7523,N_7482,N_7262);
nor U7524 (N_7524,N_7383,N_7271);
nor U7525 (N_7525,N_7258,N_7277);
nand U7526 (N_7526,N_7396,N_7497);
nand U7527 (N_7527,N_7340,N_7294);
nand U7528 (N_7528,N_7411,N_7375);
nor U7529 (N_7529,N_7456,N_7490);
nand U7530 (N_7530,N_7255,N_7412);
nor U7531 (N_7531,N_7489,N_7296);
xor U7532 (N_7532,N_7462,N_7363);
nand U7533 (N_7533,N_7379,N_7447);
nor U7534 (N_7534,N_7405,N_7432);
or U7535 (N_7535,N_7457,N_7303);
nand U7536 (N_7536,N_7257,N_7395);
nor U7537 (N_7537,N_7324,N_7279);
and U7538 (N_7538,N_7406,N_7306);
nand U7539 (N_7539,N_7460,N_7358);
or U7540 (N_7540,N_7446,N_7282);
xor U7541 (N_7541,N_7483,N_7376);
or U7542 (N_7542,N_7321,N_7287);
and U7543 (N_7543,N_7491,N_7393);
or U7544 (N_7544,N_7327,N_7478);
nor U7545 (N_7545,N_7386,N_7424);
nor U7546 (N_7546,N_7355,N_7444);
xnor U7547 (N_7547,N_7349,N_7449);
or U7548 (N_7548,N_7275,N_7284);
nor U7549 (N_7549,N_7382,N_7465);
nor U7550 (N_7550,N_7356,N_7445);
nand U7551 (N_7551,N_7397,N_7494);
xor U7552 (N_7552,N_7318,N_7374);
and U7553 (N_7553,N_7290,N_7268);
or U7554 (N_7554,N_7336,N_7289);
nor U7555 (N_7555,N_7467,N_7300);
nand U7556 (N_7556,N_7270,N_7390);
xnor U7557 (N_7557,N_7431,N_7461);
and U7558 (N_7558,N_7473,N_7442);
nand U7559 (N_7559,N_7429,N_7333);
nor U7560 (N_7560,N_7341,N_7256);
or U7561 (N_7561,N_7335,N_7435);
or U7562 (N_7562,N_7458,N_7392);
nand U7563 (N_7563,N_7487,N_7347);
or U7564 (N_7564,N_7264,N_7394);
or U7565 (N_7565,N_7301,N_7404);
or U7566 (N_7566,N_7369,N_7418);
nand U7567 (N_7567,N_7365,N_7451);
nand U7568 (N_7568,N_7387,N_7377);
and U7569 (N_7569,N_7343,N_7370);
nor U7570 (N_7570,N_7316,N_7415);
xnor U7571 (N_7571,N_7378,N_7314);
xnor U7572 (N_7572,N_7361,N_7423);
nand U7573 (N_7573,N_7260,N_7338);
and U7574 (N_7574,N_7434,N_7488);
nor U7575 (N_7575,N_7440,N_7311);
nor U7576 (N_7576,N_7466,N_7288);
or U7577 (N_7577,N_7305,N_7471);
or U7578 (N_7578,N_7353,N_7409);
nand U7579 (N_7579,N_7388,N_7267);
nor U7580 (N_7580,N_7419,N_7280);
nand U7581 (N_7581,N_7308,N_7420);
and U7582 (N_7582,N_7499,N_7348);
nand U7583 (N_7583,N_7399,N_7354);
nand U7584 (N_7584,N_7362,N_7359);
or U7585 (N_7585,N_7325,N_7463);
nand U7586 (N_7586,N_7299,N_7479);
nor U7587 (N_7587,N_7428,N_7269);
nand U7588 (N_7588,N_7323,N_7342);
nand U7589 (N_7589,N_7385,N_7367);
or U7590 (N_7590,N_7474,N_7319);
nor U7591 (N_7591,N_7315,N_7329);
nand U7592 (N_7592,N_7425,N_7480);
nor U7593 (N_7593,N_7310,N_7477);
nor U7594 (N_7594,N_7401,N_7273);
or U7595 (N_7595,N_7366,N_7368);
nand U7596 (N_7596,N_7326,N_7252);
xnor U7597 (N_7597,N_7297,N_7357);
nand U7598 (N_7598,N_7496,N_7476);
or U7599 (N_7599,N_7371,N_7261);
nand U7600 (N_7600,N_7330,N_7389);
or U7601 (N_7601,N_7422,N_7400);
or U7602 (N_7602,N_7436,N_7421);
nor U7603 (N_7603,N_7251,N_7384);
xnor U7604 (N_7604,N_7360,N_7322);
nor U7605 (N_7605,N_7495,N_7334);
and U7606 (N_7606,N_7470,N_7304);
or U7607 (N_7607,N_7312,N_7265);
nor U7608 (N_7608,N_7272,N_7346);
nand U7609 (N_7609,N_7468,N_7441);
or U7610 (N_7610,N_7274,N_7452);
nand U7611 (N_7611,N_7453,N_7364);
xor U7612 (N_7612,N_7291,N_7292);
xnor U7613 (N_7613,N_7339,N_7416);
or U7614 (N_7614,N_7286,N_7380);
nor U7615 (N_7615,N_7352,N_7427);
nor U7616 (N_7616,N_7450,N_7433);
or U7617 (N_7617,N_7373,N_7345);
and U7618 (N_7618,N_7350,N_7266);
and U7619 (N_7619,N_7417,N_7486);
and U7620 (N_7620,N_7469,N_7254);
or U7621 (N_7621,N_7276,N_7492);
nand U7622 (N_7622,N_7351,N_7337);
and U7623 (N_7623,N_7403,N_7309);
nor U7624 (N_7624,N_7410,N_7344);
or U7625 (N_7625,N_7439,N_7327);
nand U7626 (N_7626,N_7251,N_7309);
and U7627 (N_7627,N_7397,N_7390);
nand U7628 (N_7628,N_7389,N_7403);
nor U7629 (N_7629,N_7304,N_7427);
nand U7630 (N_7630,N_7469,N_7291);
nand U7631 (N_7631,N_7337,N_7384);
xnor U7632 (N_7632,N_7472,N_7432);
or U7633 (N_7633,N_7261,N_7431);
and U7634 (N_7634,N_7318,N_7272);
xor U7635 (N_7635,N_7252,N_7271);
or U7636 (N_7636,N_7423,N_7394);
or U7637 (N_7637,N_7325,N_7428);
and U7638 (N_7638,N_7406,N_7334);
and U7639 (N_7639,N_7296,N_7298);
xor U7640 (N_7640,N_7330,N_7498);
nand U7641 (N_7641,N_7339,N_7311);
nor U7642 (N_7642,N_7365,N_7302);
nand U7643 (N_7643,N_7282,N_7489);
nand U7644 (N_7644,N_7330,N_7418);
and U7645 (N_7645,N_7336,N_7452);
nand U7646 (N_7646,N_7303,N_7476);
and U7647 (N_7647,N_7492,N_7326);
and U7648 (N_7648,N_7260,N_7323);
nor U7649 (N_7649,N_7420,N_7317);
nand U7650 (N_7650,N_7315,N_7423);
and U7651 (N_7651,N_7343,N_7250);
and U7652 (N_7652,N_7438,N_7417);
and U7653 (N_7653,N_7477,N_7315);
nor U7654 (N_7654,N_7429,N_7440);
and U7655 (N_7655,N_7433,N_7493);
nor U7656 (N_7656,N_7382,N_7251);
nand U7657 (N_7657,N_7452,N_7367);
nand U7658 (N_7658,N_7312,N_7451);
nor U7659 (N_7659,N_7356,N_7417);
nor U7660 (N_7660,N_7441,N_7312);
nand U7661 (N_7661,N_7273,N_7389);
or U7662 (N_7662,N_7425,N_7467);
nand U7663 (N_7663,N_7478,N_7335);
nor U7664 (N_7664,N_7328,N_7294);
and U7665 (N_7665,N_7424,N_7429);
and U7666 (N_7666,N_7303,N_7499);
and U7667 (N_7667,N_7355,N_7405);
and U7668 (N_7668,N_7496,N_7468);
nor U7669 (N_7669,N_7461,N_7441);
and U7670 (N_7670,N_7319,N_7451);
nand U7671 (N_7671,N_7253,N_7449);
nor U7672 (N_7672,N_7495,N_7454);
or U7673 (N_7673,N_7448,N_7284);
nor U7674 (N_7674,N_7480,N_7331);
nand U7675 (N_7675,N_7292,N_7493);
nand U7676 (N_7676,N_7472,N_7333);
nand U7677 (N_7677,N_7388,N_7485);
and U7678 (N_7678,N_7403,N_7421);
or U7679 (N_7679,N_7445,N_7428);
nor U7680 (N_7680,N_7365,N_7257);
nand U7681 (N_7681,N_7353,N_7482);
nor U7682 (N_7682,N_7311,N_7410);
or U7683 (N_7683,N_7368,N_7378);
nand U7684 (N_7684,N_7356,N_7493);
or U7685 (N_7685,N_7417,N_7342);
or U7686 (N_7686,N_7262,N_7452);
or U7687 (N_7687,N_7259,N_7322);
or U7688 (N_7688,N_7433,N_7463);
nand U7689 (N_7689,N_7442,N_7317);
and U7690 (N_7690,N_7349,N_7312);
xor U7691 (N_7691,N_7363,N_7333);
nand U7692 (N_7692,N_7308,N_7253);
nor U7693 (N_7693,N_7252,N_7380);
or U7694 (N_7694,N_7279,N_7326);
nor U7695 (N_7695,N_7363,N_7463);
and U7696 (N_7696,N_7297,N_7314);
and U7697 (N_7697,N_7338,N_7417);
and U7698 (N_7698,N_7336,N_7320);
nor U7699 (N_7699,N_7387,N_7299);
nor U7700 (N_7700,N_7343,N_7401);
nand U7701 (N_7701,N_7422,N_7332);
or U7702 (N_7702,N_7267,N_7491);
and U7703 (N_7703,N_7259,N_7435);
and U7704 (N_7704,N_7251,N_7479);
nand U7705 (N_7705,N_7474,N_7325);
or U7706 (N_7706,N_7441,N_7337);
nor U7707 (N_7707,N_7423,N_7436);
nand U7708 (N_7708,N_7366,N_7438);
xor U7709 (N_7709,N_7359,N_7387);
and U7710 (N_7710,N_7276,N_7412);
and U7711 (N_7711,N_7270,N_7330);
xnor U7712 (N_7712,N_7259,N_7377);
nor U7713 (N_7713,N_7384,N_7355);
nor U7714 (N_7714,N_7395,N_7424);
or U7715 (N_7715,N_7340,N_7385);
xnor U7716 (N_7716,N_7381,N_7376);
or U7717 (N_7717,N_7435,N_7383);
nor U7718 (N_7718,N_7471,N_7328);
nand U7719 (N_7719,N_7460,N_7463);
and U7720 (N_7720,N_7428,N_7494);
nand U7721 (N_7721,N_7412,N_7316);
or U7722 (N_7722,N_7300,N_7414);
nor U7723 (N_7723,N_7303,N_7278);
nor U7724 (N_7724,N_7286,N_7334);
nand U7725 (N_7725,N_7334,N_7288);
or U7726 (N_7726,N_7462,N_7485);
nor U7727 (N_7727,N_7469,N_7486);
nor U7728 (N_7728,N_7264,N_7483);
nand U7729 (N_7729,N_7371,N_7256);
or U7730 (N_7730,N_7416,N_7432);
or U7731 (N_7731,N_7351,N_7393);
nor U7732 (N_7732,N_7444,N_7439);
nor U7733 (N_7733,N_7368,N_7437);
or U7734 (N_7734,N_7371,N_7284);
nand U7735 (N_7735,N_7452,N_7440);
nor U7736 (N_7736,N_7307,N_7310);
nand U7737 (N_7737,N_7280,N_7497);
nor U7738 (N_7738,N_7298,N_7393);
and U7739 (N_7739,N_7356,N_7274);
xor U7740 (N_7740,N_7283,N_7435);
and U7741 (N_7741,N_7420,N_7335);
nor U7742 (N_7742,N_7425,N_7334);
xnor U7743 (N_7743,N_7345,N_7473);
and U7744 (N_7744,N_7289,N_7474);
nor U7745 (N_7745,N_7410,N_7455);
nor U7746 (N_7746,N_7299,N_7476);
nand U7747 (N_7747,N_7281,N_7398);
and U7748 (N_7748,N_7395,N_7354);
nor U7749 (N_7749,N_7403,N_7250);
xor U7750 (N_7750,N_7678,N_7597);
or U7751 (N_7751,N_7592,N_7520);
nor U7752 (N_7752,N_7566,N_7668);
xor U7753 (N_7753,N_7687,N_7624);
xor U7754 (N_7754,N_7543,N_7614);
nor U7755 (N_7755,N_7518,N_7605);
xor U7756 (N_7756,N_7588,N_7527);
nor U7757 (N_7757,N_7729,N_7655);
and U7758 (N_7758,N_7516,N_7573);
nand U7759 (N_7759,N_7617,N_7541);
and U7760 (N_7760,N_7737,N_7623);
or U7761 (N_7761,N_7599,N_7611);
nor U7762 (N_7762,N_7690,N_7734);
xnor U7763 (N_7763,N_7529,N_7533);
nand U7764 (N_7764,N_7702,N_7556);
nor U7765 (N_7765,N_7580,N_7576);
and U7766 (N_7766,N_7583,N_7713);
nor U7767 (N_7767,N_7646,N_7717);
and U7768 (N_7768,N_7513,N_7530);
and U7769 (N_7769,N_7712,N_7552);
or U7770 (N_7770,N_7582,N_7521);
nor U7771 (N_7771,N_7695,N_7720);
nor U7772 (N_7772,N_7616,N_7648);
nand U7773 (N_7773,N_7620,N_7662);
or U7774 (N_7774,N_7600,N_7632);
nand U7775 (N_7775,N_7501,N_7504);
and U7776 (N_7776,N_7524,N_7663);
and U7777 (N_7777,N_7581,N_7650);
nand U7778 (N_7778,N_7571,N_7666);
nor U7779 (N_7779,N_7680,N_7548);
nor U7780 (N_7780,N_7633,N_7686);
or U7781 (N_7781,N_7664,N_7740);
nor U7782 (N_7782,N_7508,N_7682);
and U7783 (N_7783,N_7558,N_7515);
xor U7784 (N_7784,N_7739,N_7715);
nor U7785 (N_7785,N_7550,N_7639);
or U7786 (N_7786,N_7636,N_7511);
or U7787 (N_7787,N_7629,N_7572);
nor U7788 (N_7788,N_7670,N_7679);
and U7789 (N_7789,N_7719,N_7509);
nand U7790 (N_7790,N_7522,N_7743);
nand U7791 (N_7791,N_7728,N_7612);
xnor U7792 (N_7792,N_7747,N_7593);
nor U7793 (N_7793,N_7741,N_7707);
or U7794 (N_7794,N_7708,N_7506);
and U7795 (N_7795,N_7726,N_7642);
nor U7796 (N_7796,N_7718,N_7586);
and U7797 (N_7797,N_7585,N_7652);
or U7798 (N_7798,N_7748,N_7565);
nand U7799 (N_7799,N_7727,N_7602);
nor U7800 (N_7800,N_7570,N_7746);
nor U7801 (N_7801,N_7613,N_7595);
and U7802 (N_7802,N_7535,N_7704);
and U7803 (N_7803,N_7626,N_7667);
and U7804 (N_7804,N_7738,N_7564);
and U7805 (N_7805,N_7507,N_7544);
xor U7806 (N_7806,N_7697,N_7696);
nand U7807 (N_7807,N_7619,N_7536);
nand U7808 (N_7808,N_7540,N_7677);
xor U7809 (N_7809,N_7590,N_7724);
or U7810 (N_7810,N_7731,N_7553);
nand U7811 (N_7811,N_7688,N_7563);
nand U7812 (N_7812,N_7630,N_7512);
or U7813 (N_7813,N_7654,N_7596);
nand U7814 (N_7814,N_7587,N_7574);
nand U7815 (N_7815,N_7594,N_7621);
and U7816 (N_7816,N_7549,N_7672);
nor U7817 (N_7817,N_7510,N_7693);
and U7818 (N_7818,N_7607,N_7584);
and U7819 (N_7819,N_7625,N_7545);
nor U7820 (N_7820,N_7742,N_7730);
or U7821 (N_7821,N_7542,N_7627);
xor U7822 (N_7822,N_7555,N_7560);
and U7823 (N_7823,N_7661,N_7532);
or U7824 (N_7824,N_7559,N_7660);
and U7825 (N_7825,N_7669,N_7526);
nand U7826 (N_7826,N_7637,N_7500);
nand U7827 (N_7827,N_7736,N_7685);
or U7828 (N_7828,N_7554,N_7631);
nand U7829 (N_7829,N_7723,N_7517);
nand U7830 (N_7830,N_7537,N_7575);
nor U7831 (N_7831,N_7606,N_7745);
xor U7832 (N_7832,N_7567,N_7683);
nand U7833 (N_7833,N_7657,N_7681);
or U7834 (N_7834,N_7716,N_7665);
nand U7835 (N_7835,N_7610,N_7505);
nand U7836 (N_7836,N_7722,N_7711);
and U7837 (N_7837,N_7675,N_7538);
nand U7838 (N_7838,N_7603,N_7699);
nor U7839 (N_7839,N_7609,N_7691);
xor U7840 (N_7840,N_7618,N_7644);
nand U7841 (N_7841,N_7604,N_7634);
nand U7842 (N_7842,N_7591,N_7577);
nand U7843 (N_7843,N_7653,N_7598);
and U7844 (N_7844,N_7579,N_7638);
xor U7845 (N_7845,N_7523,N_7735);
nand U7846 (N_7846,N_7689,N_7701);
and U7847 (N_7847,N_7615,N_7698);
nor U7848 (N_7848,N_7561,N_7539);
xor U7849 (N_7849,N_7622,N_7643);
and U7850 (N_7850,N_7601,N_7562);
or U7851 (N_7851,N_7514,N_7503);
or U7852 (N_7852,N_7589,N_7721);
xnor U7853 (N_7853,N_7703,N_7546);
xnor U7854 (N_7854,N_7725,N_7519);
and U7855 (N_7855,N_7706,N_7656);
or U7856 (N_7856,N_7647,N_7525);
or U7857 (N_7857,N_7749,N_7733);
nand U7858 (N_7858,N_7641,N_7692);
nand U7859 (N_7859,N_7534,N_7744);
nand U7860 (N_7860,N_7709,N_7531);
nand U7861 (N_7861,N_7568,N_7732);
nor U7862 (N_7862,N_7714,N_7547);
xnor U7863 (N_7863,N_7569,N_7557);
nor U7864 (N_7864,N_7710,N_7651);
nand U7865 (N_7865,N_7640,N_7700);
and U7866 (N_7866,N_7528,N_7705);
nor U7867 (N_7867,N_7502,N_7649);
nor U7868 (N_7868,N_7658,N_7676);
and U7869 (N_7869,N_7645,N_7608);
nor U7870 (N_7870,N_7671,N_7684);
and U7871 (N_7871,N_7674,N_7628);
or U7872 (N_7872,N_7578,N_7659);
or U7873 (N_7873,N_7635,N_7673);
nand U7874 (N_7874,N_7551,N_7694);
or U7875 (N_7875,N_7654,N_7658);
and U7876 (N_7876,N_7543,N_7553);
nor U7877 (N_7877,N_7733,N_7711);
nand U7878 (N_7878,N_7657,N_7621);
nand U7879 (N_7879,N_7674,N_7651);
nand U7880 (N_7880,N_7645,N_7749);
nor U7881 (N_7881,N_7698,N_7703);
nand U7882 (N_7882,N_7627,N_7749);
xor U7883 (N_7883,N_7623,N_7648);
or U7884 (N_7884,N_7528,N_7707);
nor U7885 (N_7885,N_7730,N_7692);
nor U7886 (N_7886,N_7550,N_7558);
and U7887 (N_7887,N_7560,N_7715);
or U7888 (N_7888,N_7743,N_7512);
and U7889 (N_7889,N_7717,N_7682);
and U7890 (N_7890,N_7666,N_7653);
or U7891 (N_7891,N_7602,N_7656);
and U7892 (N_7892,N_7531,N_7598);
nand U7893 (N_7893,N_7602,N_7582);
and U7894 (N_7894,N_7650,N_7594);
or U7895 (N_7895,N_7619,N_7578);
and U7896 (N_7896,N_7608,N_7730);
xnor U7897 (N_7897,N_7537,N_7663);
or U7898 (N_7898,N_7709,N_7527);
and U7899 (N_7899,N_7678,N_7714);
nand U7900 (N_7900,N_7613,N_7540);
nor U7901 (N_7901,N_7585,N_7595);
nand U7902 (N_7902,N_7537,N_7632);
nor U7903 (N_7903,N_7700,N_7618);
nand U7904 (N_7904,N_7520,N_7669);
xor U7905 (N_7905,N_7671,N_7672);
nand U7906 (N_7906,N_7698,N_7509);
nor U7907 (N_7907,N_7637,N_7547);
xor U7908 (N_7908,N_7744,N_7599);
and U7909 (N_7909,N_7633,N_7559);
and U7910 (N_7910,N_7708,N_7652);
nor U7911 (N_7911,N_7719,N_7510);
or U7912 (N_7912,N_7520,N_7703);
nand U7913 (N_7913,N_7740,N_7645);
or U7914 (N_7914,N_7655,N_7677);
nand U7915 (N_7915,N_7519,N_7724);
nor U7916 (N_7916,N_7631,N_7678);
nand U7917 (N_7917,N_7644,N_7647);
xnor U7918 (N_7918,N_7705,N_7539);
nand U7919 (N_7919,N_7558,N_7571);
and U7920 (N_7920,N_7637,N_7622);
xnor U7921 (N_7921,N_7669,N_7548);
nand U7922 (N_7922,N_7552,N_7588);
or U7923 (N_7923,N_7600,N_7516);
or U7924 (N_7924,N_7722,N_7744);
nand U7925 (N_7925,N_7749,N_7671);
and U7926 (N_7926,N_7650,N_7589);
nand U7927 (N_7927,N_7579,N_7663);
and U7928 (N_7928,N_7555,N_7581);
and U7929 (N_7929,N_7729,N_7580);
nor U7930 (N_7930,N_7507,N_7690);
and U7931 (N_7931,N_7598,N_7589);
nand U7932 (N_7932,N_7743,N_7500);
or U7933 (N_7933,N_7738,N_7652);
or U7934 (N_7934,N_7595,N_7734);
xor U7935 (N_7935,N_7568,N_7609);
or U7936 (N_7936,N_7614,N_7661);
nand U7937 (N_7937,N_7741,N_7532);
nor U7938 (N_7938,N_7647,N_7690);
or U7939 (N_7939,N_7524,N_7581);
nor U7940 (N_7940,N_7744,N_7694);
nor U7941 (N_7941,N_7735,N_7721);
or U7942 (N_7942,N_7650,N_7631);
and U7943 (N_7943,N_7682,N_7569);
or U7944 (N_7944,N_7631,N_7686);
and U7945 (N_7945,N_7619,N_7682);
nand U7946 (N_7946,N_7535,N_7715);
nand U7947 (N_7947,N_7580,N_7584);
nand U7948 (N_7948,N_7698,N_7728);
and U7949 (N_7949,N_7726,N_7651);
nand U7950 (N_7950,N_7709,N_7714);
xnor U7951 (N_7951,N_7609,N_7522);
nor U7952 (N_7952,N_7645,N_7616);
and U7953 (N_7953,N_7641,N_7501);
and U7954 (N_7954,N_7668,N_7674);
or U7955 (N_7955,N_7508,N_7664);
and U7956 (N_7956,N_7578,N_7668);
nor U7957 (N_7957,N_7609,N_7552);
and U7958 (N_7958,N_7618,N_7583);
nand U7959 (N_7959,N_7559,N_7693);
nand U7960 (N_7960,N_7587,N_7606);
nand U7961 (N_7961,N_7528,N_7570);
nor U7962 (N_7962,N_7579,N_7642);
nor U7963 (N_7963,N_7649,N_7624);
or U7964 (N_7964,N_7633,N_7638);
nor U7965 (N_7965,N_7618,N_7686);
and U7966 (N_7966,N_7736,N_7697);
and U7967 (N_7967,N_7620,N_7676);
and U7968 (N_7968,N_7576,N_7617);
nand U7969 (N_7969,N_7688,N_7605);
xnor U7970 (N_7970,N_7528,N_7730);
nor U7971 (N_7971,N_7689,N_7648);
nor U7972 (N_7972,N_7512,N_7670);
nand U7973 (N_7973,N_7565,N_7513);
nor U7974 (N_7974,N_7604,N_7731);
and U7975 (N_7975,N_7521,N_7660);
nor U7976 (N_7976,N_7624,N_7719);
or U7977 (N_7977,N_7674,N_7703);
nand U7978 (N_7978,N_7667,N_7560);
and U7979 (N_7979,N_7577,N_7551);
nor U7980 (N_7980,N_7640,N_7613);
nor U7981 (N_7981,N_7638,N_7503);
and U7982 (N_7982,N_7540,N_7516);
or U7983 (N_7983,N_7643,N_7585);
and U7984 (N_7984,N_7535,N_7672);
nor U7985 (N_7985,N_7725,N_7531);
xor U7986 (N_7986,N_7517,N_7653);
nand U7987 (N_7987,N_7711,N_7527);
nor U7988 (N_7988,N_7712,N_7631);
or U7989 (N_7989,N_7701,N_7565);
and U7990 (N_7990,N_7735,N_7743);
nor U7991 (N_7991,N_7563,N_7607);
or U7992 (N_7992,N_7629,N_7619);
nor U7993 (N_7993,N_7589,N_7635);
xor U7994 (N_7994,N_7726,N_7522);
and U7995 (N_7995,N_7531,N_7561);
nor U7996 (N_7996,N_7733,N_7746);
xor U7997 (N_7997,N_7652,N_7526);
nor U7998 (N_7998,N_7640,N_7638);
and U7999 (N_7999,N_7541,N_7678);
nor U8000 (N_8000,N_7948,N_7995);
and U8001 (N_8001,N_7929,N_7863);
xor U8002 (N_8002,N_7949,N_7869);
nor U8003 (N_8003,N_7844,N_7784);
nor U8004 (N_8004,N_7840,N_7901);
or U8005 (N_8005,N_7881,N_7757);
and U8006 (N_8006,N_7775,N_7825);
or U8007 (N_8007,N_7909,N_7983);
and U8008 (N_8008,N_7846,N_7816);
nor U8009 (N_8009,N_7808,N_7986);
and U8010 (N_8010,N_7865,N_7954);
nor U8011 (N_8011,N_7771,N_7812);
nand U8012 (N_8012,N_7867,N_7820);
nand U8013 (N_8013,N_7829,N_7841);
xor U8014 (N_8014,N_7975,N_7979);
xnor U8015 (N_8015,N_7951,N_7911);
nand U8016 (N_8016,N_7776,N_7802);
nand U8017 (N_8017,N_7786,N_7770);
nand U8018 (N_8018,N_7999,N_7781);
or U8019 (N_8019,N_7896,N_7964);
xnor U8020 (N_8020,N_7800,N_7972);
nor U8021 (N_8021,N_7967,N_7906);
or U8022 (N_8022,N_7918,N_7762);
and U8023 (N_8023,N_7772,N_7847);
nor U8024 (N_8024,N_7871,N_7822);
nor U8025 (N_8025,N_7789,N_7859);
xnor U8026 (N_8026,N_7850,N_7917);
and U8027 (N_8027,N_7882,N_7766);
nor U8028 (N_8028,N_7916,N_7971);
and U8029 (N_8029,N_7893,N_7946);
xor U8030 (N_8030,N_7858,N_7837);
nor U8031 (N_8031,N_7985,N_7980);
xnor U8032 (N_8032,N_7815,N_7994);
nand U8033 (N_8033,N_7814,N_7810);
nand U8034 (N_8034,N_7805,N_7774);
or U8035 (N_8035,N_7934,N_7852);
xor U8036 (N_8036,N_7862,N_7904);
nand U8037 (N_8037,N_7780,N_7883);
nand U8038 (N_8038,N_7941,N_7834);
nor U8039 (N_8039,N_7927,N_7796);
nand U8040 (N_8040,N_7777,N_7799);
xnor U8041 (N_8041,N_7887,N_7750);
nor U8042 (N_8042,N_7760,N_7861);
nor U8043 (N_8043,N_7889,N_7765);
or U8044 (N_8044,N_7895,N_7966);
nand U8045 (N_8045,N_7952,N_7935);
or U8046 (N_8046,N_7940,N_7768);
nor U8047 (N_8047,N_7987,N_7924);
nand U8048 (N_8048,N_7791,N_7913);
or U8049 (N_8049,N_7880,N_7806);
nor U8050 (N_8050,N_7813,N_7794);
or U8051 (N_8051,N_7976,N_7832);
nor U8052 (N_8052,N_7908,N_7845);
and U8053 (N_8053,N_7960,N_7956);
or U8054 (N_8054,N_7892,N_7989);
xor U8055 (N_8055,N_7992,N_7835);
and U8056 (N_8056,N_7752,N_7769);
xnor U8057 (N_8057,N_7782,N_7758);
nand U8058 (N_8058,N_7943,N_7885);
nor U8059 (N_8059,N_7804,N_7756);
or U8060 (N_8060,N_7886,N_7767);
nand U8061 (N_8061,N_7932,N_7945);
nor U8062 (N_8062,N_7902,N_7950);
nand U8063 (N_8063,N_7860,N_7928);
nand U8064 (N_8064,N_7833,N_7849);
nor U8065 (N_8065,N_7915,N_7962);
or U8066 (N_8066,N_7891,N_7821);
or U8067 (N_8067,N_7974,N_7823);
nor U8068 (N_8068,N_7899,N_7857);
or U8069 (N_8069,N_7998,N_7873);
nand U8070 (N_8070,N_7968,N_7991);
nand U8071 (N_8071,N_7783,N_7751);
nor U8072 (N_8072,N_7773,N_7856);
nand U8073 (N_8073,N_7853,N_7926);
nand U8074 (N_8074,N_7939,N_7936);
nand U8075 (N_8075,N_7912,N_7933);
or U8076 (N_8076,N_7763,N_7828);
nor U8077 (N_8077,N_7779,N_7826);
and U8078 (N_8078,N_7836,N_7961);
nor U8079 (N_8079,N_7817,N_7888);
xnor U8080 (N_8080,N_7803,N_7997);
nor U8081 (N_8081,N_7793,N_7955);
nand U8082 (N_8082,N_7996,N_7905);
nand U8083 (N_8083,N_7819,N_7801);
nand U8084 (N_8084,N_7978,N_7843);
or U8085 (N_8085,N_7963,N_7764);
and U8086 (N_8086,N_7855,N_7953);
nor U8087 (N_8087,N_7854,N_7759);
or U8088 (N_8088,N_7942,N_7778);
or U8089 (N_8089,N_7923,N_7795);
and U8090 (N_8090,N_7914,N_7984);
nor U8091 (N_8091,N_7838,N_7761);
or U8092 (N_8092,N_7753,N_7993);
xnor U8093 (N_8093,N_7910,N_7900);
and U8094 (N_8094,N_7754,N_7879);
and U8095 (N_8095,N_7864,N_7930);
nor U8096 (N_8096,N_7809,N_7903);
nor U8097 (N_8097,N_7907,N_7959);
nor U8098 (N_8098,N_7890,N_7969);
or U8099 (N_8099,N_7851,N_7872);
nand U8100 (N_8100,N_7982,N_7874);
nor U8101 (N_8101,N_7897,N_7973);
or U8102 (N_8102,N_7977,N_7925);
nor U8103 (N_8103,N_7990,N_7868);
or U8104 (N_8104,N_7827,N_7830);
nand U8105 (N_8105,N_7839,N_7824);
or U8106 (N_8106,N_7785,N_7988);
nor U8107 (N_8107,N_7919,N_7755);
and U8108 (N_8108,N_7937,N_7877);
xor U8109 (N_8109,N_7957,N_7876);
nand U8110 (N_8110,N_7818,N_7848);
and U8111 (N_8111,N_7798,N_7866);
or U8112 (N_8112,N_7875,N_7831);
or U8113 (N_8113,N_7797,N_7884);
or U8114 (N_8114,N_7922,N_7898);
or U8115 (N_8115,N_7787,N_7981);
nand U8116 (N_8116,N_7792,N_7921);
and U8117 (N_8117,N_7842,N_7894);
nor U8118 (N_8118,N_7938,N_7807);
nor U8119 (N_8119,N_7970,N_7947);
nand U8120 (N_8120,N_7790,N_7944);
nand U8121 (N_8121,N_7878,N_7788);
nand U8122 (N_8122,N_7870,N_7965);
nor U8123 (N_8123,N_7931,N_7958);
nand U8124 (N_8124,N_7920,N_7811);
nor U8125 (N_8125,N_7921,N_7853);
nor U8126 (N_8126,N_7789,N_7830);
and U8127 (N_8127,N_7967,N_7768);
and U8128 (N_8128,N_7913,N_7871);
or U8129 (N_8129,N_7860,N_7997);
or U8130 (N_8130,N_7862,N_7809);
nand U8131 (N_8131,N_7760,N_7883);
nor U8132 (N_8132,N_7893,N_7879);
or U8133 (N_8133,N_7870,N_7757);
or U8134 (N_8134,N_7921,N_7838);
or U8135 (N_8135,N_7951,N_7949);
nor U8136 (N_8136,N_7769,N_7992);
nand U8137 (N_8137,N_7983,N_7767);
and U8138 (N_8138,N_7789,N_7894);
or U8139 (N_8139,N_7898,N_7882);
nand U8140 (N_8140,N_7993,N_7930);
and U8141 (N_8141,N_7766,N_7956);
nand U8142 (N_8142,N_7819,N_7934);
nand U8143 (N_8143,N_7814,N_7855);
nor U8144 (N_8144,N_7833,N_7998);
nor U8145 (N_8145,N_7824,N_7801);
xor U8146 (N_8146,N_7967,N_7793);
and U8147 (N_8147,N_7857,N_7825);
nor U8148 (N_8148,N_7884,N_7882);
nor U8149 (N_8149,N_7784,N_7841);
nor U8150 (N_8150,N_7841,N_7759);
nor U8151 (N_8151,N_7949,N_7957);
or U8152 (N_8152,N_7933,N_7903);
or U8153 (N_8153,N_7949,N_7991);
xnor U8154 (N_8154,N_7878,N_7823);
or U8155 (N_8155,N_7922,N_7762);
nor U8156 (N_8156,N_7981,N_7794);
nor U8157 (N_8157,N_7928,N_7813);
or U8158 (N_8158,N_7977,N_7905);
or U8159 (N_8159,N_7966,N_7991);
xnor U8160 (N_8160,N_7801,N_7841);
nand U8161 (N_8161,N_7866,N_7949);
nor U8162 (N_8162,N_7874,N_7837);
nand U8163 (N_8163,N_7881,N_7961);
nand U8164 (N_8164,N_7814,N_7893);
or U8165 (N_8165,N_7815,N_7935);
xor U8166 (N_8166,N_7999,N_7936);
nor U8167 (N_8167,N_7989,N_7954);
nand U8168 (N_8168,N_7874,N_7914);
and U8169 (N_8169,N_7762,N_7992);
nand U8170 (N_8170,N_7759,N_7767);
or U8171 (N_8171,N_7827,N_7989);
nand U8172 (N_8172,N_7915,N_7862);
nor U8173 (N_8173,N_7882,N_7791);
or U8174 (N_8174,N_7952,N_7864);
nor U8175 (N_8175,N_7996,N_7971);
nand U8176 (N_8176,N_7987,N_7921);
nand U8177 (N_8177,N_7971,N_7877);
or U8178 (N_8178,N_7767,N_7999);
nor U8179 (N_8179,N_7897,N_7839);
or U8180 (N_8180,N_7768,N_7817);
and U8181 (N_8181,N_7781,N_7767);
nand U8182 (N_8182,N_7973,N_7796);
xor U8183 (N_8183,N_7777,N_7916);
or U8184 (N_8184,N_7930,N_7855);
nand U8185 (N_8185,N_7806,N_7754);
nor U8186 (N_8186,N_7756,N_7938);
xnor U8187 (N_8187,N_7856,N_7940);
and U8188 (N_8188,N_7935,N_7890);
or U8189 (N_8189,N_7817,N_7845);
and U8190 (N_8190,N_7828,N_7874);
nor U8191 (N_8191,N_7867,N_7984);
or U8192 (N_8192,N_7890,N_7911);
xnor U8193 (N_8193,N_7920,N_7790);
and U8194 (N_8194,N_7922,N_7984);
and U8195 (N_8195,N_7854,N_7912);
and U8196 (N_8196,N_7812,N_7815);
and U8197 (N_8197,N_7827,N_7999);
and U8198 (N_8198,N_7867,N_7779);
nand U8199 (N_8199,N_7831,N_7805);
or U8200 (N_8200,N_7809,N_7989);
or U8201 (N_8201,N_7774,N_7998);
nand U8202 (N_8202,N_7815,N_7820);
nor U8203 (N_8203,N_7899,N_7824);
and U8204 (N_8204,N_7944,N_7882);
or U8205 (N_8205,N_7933,N_7769);
nor U8206 (N_8206,N_7841,N_7798);
or U8207 (N_8207,N_7882,N_7897);
nor U8208 (N_8208,N_7762,N_7763);
or U8209 (N_8209,N_7996,N_7825);
nor U8210 (N_8210,N_7919,N_7964);
xnor U8211 (N_8211,N_7920,N_7851);
nand U8212 (N_8212,N_7788,N_7773);
nor U8213 (N_8213,N_7870,N_7809);
and U8214 (N_8214,N_7765,N_7843);
nand U8215 (N_8215,N_7910,N_7783);
and U8216 (N_8216,N_7827,N_7954);
and U8217 (N_8217,N_7941,N_7879);
or U8218 (N_8218,N_7791,N_7928);
nand U8219 (N_8219,N_7967,N_7780);
and U8220 (N_8220,N_7873,N_7813);
or U8221 (N_8221,N_7827,N_7844);
or U8222 (N_8222,N_7973,N_7833);
or U8223 (N_8223,N_7926,N_7806);
or U8224 (N_8224,N_7902,N_7984);
nand U8225 (N_8225,N_7912,N_7812);
xor U8226 (N_8226,N_7774,N_7775);
nor U8227 (N_8227,N_7851,N_7849);
nor U8228 (N_8228,N_7955,N_7988);
nor U8229 (N_8229,N_7972,N_7815);
and U8230 (N_8230,N_7901,N_7919);
xnor U8231 (N_8231,N_7938,N_7870);
nor U8232 (N_8232,N_7789,N_7782);
nor U8233 (N_8233,N_7820,N_7910);
or U8234 (N_8234,N_7996,N_7769);
nand U8235 (N_8235,N_7872,N_7875);
nor U8236 (N_8236,N_7970,N_7860);
and U8237 (N_8237,N_7862,N_7766);
xnor U8238 (N_8238,N_7933,N_7860);
or U8239 (N_8239,N_7967,N_7935);
nand U8240 (N_8240,N_7995,N_7994);
nand U8241 (N_8241,N_7750,N_7844);
nand U8242 (N_8242,N_7881,N_7838);
or U8243 (N_8243,N_7804,N_7856);
and U8244 (N_8244,N_7870,N_7819);
nor U8245 (N_8245,N_7920,N_7900);
nor U8246 (N_8246,N_7989,N_7967);
or U8247 (N_8247,N_7829,N_7838);
or U8248 (N_8248,N_7790,N_7874);
and U8249 (N_8249,N_7816,N_7962);
nand U8250 (N_8250,N_8118,N_8241);
nor U8251 (N_8251,N_8036,N_8154);
nand U8252 (N_8252,N_8020,N_8097);
or U8253 (N_8253,N_8018,N_8176);
or U8254 (N_8254,N_8088,N_8231);
and U8255 (N_8255,N_8148,N_8216);
and U8256 (N_8256,N_8081,N_8199);
nor U8257 (N_8257,N_8084,N_8203);
nor U8258 (N_8258,N_8201,N_8169);
nand U8259 (N_8259,N_8219,N_8180);
or U8260 (N_8260,N_8043,N_8016);
or U8261 (N_8261,N_8165,N_8217);
nand U8262 (N_8262,N_8156,N_8242);
or U8263 (N_8263,N_8143,N_8030);
nand U8264 (N_8264,N_8129,N_8008);
and U8265 (N_8265,N_8021,N_8247);
nor U8266 (N_8266,N_8175,N_8170);
and U8267 (N_8267,N_8104,N_8107);
xor U8268 (N_8268,N_8075,N_8208);
nor U8269 (N_8269,N_8130,N_8200);
and U8270 (N_8270,N_8237,N_8089);
nand U8271 (N_8271,N_8019,N_8172);
nand U8272 (N_8272,N_8099,N_8212);
or U8273 (N_8273,N_8090,N_8010);
nand U8274 (N_8274,N_8005,N_8164);
nand U8275 (N_8275,N_8114,N_8057);
nand U8276 (N_8276,N_8179,N_8022);
or U8277 (N_8277,N_8105,N_8235);
or U8278 (N_8278,N_8093,N_8066);
xor U8279 (N_8279,N_8085,N_8220);
nand U8280 (N_8280,N_8198,N_8101);
nand U8281 (N_8281,N_8236,N_8152);
nor U8282 (N_8282,N_8186,N_8136);
or U8283 (N_8283,N_8132,N_8206);
and U8284 (N_8284,N_8222,N_8213);
xnor U8285 (N_8285,N_8183,N_8139);
nand U8286 (N_8286,N_8063,N_8153);
nand U8287 (N_8287,N_8168,N_8048);
nor U8288 (N_8288,N_8207,N_8161);
and U8289 (N_8289,N_8028,N_8192);
nand U8290 (N_8290,N_8230,N_8062);
and U8291 (N_8291,N_8115,N_8080);
nor U8292 (N_8292,N_8195,N_8171);
nand U8293 (N_8293,N_8050,N_8095);
and U8294 (N_8294,N_8045,N_8126);
xor U8295 (N_8295,N_8160,N_8078);
nor U8296 (N_8296,N_8002,N_8127);
nor U8297 (N_8297,N_8042,N_8249);
nor U8298 (N_8298,N_8025,N_8073);
nand U8299 (N_8299,N_8162,N_8158);
and U8300 (N_8300,N_8193,N_8024);
and U8301 (N_8301,N_8121,N_8068);
or U8302 (N_8302,N_8026,N_8091);
nor U8303 (N_8303,N_8226,N_8218);
xor U8304 (N_8304,N_8079,N_8044);
or U8305 (N_8305,N_8058,N_8248);
xnor U8306 (N_8306,N_8145,N_8069);
and U8307 (N_8307,N_8188,N_8037);
and U8308 (N_8308,N_8196,N_8067);
xor U8309 (N_8309,N_8049,N_8119);
nor U8310 (N_8310,N_8125,N_8159);
nand U8311 (N_8311,N_8013,N_8173);
nor U8312 (N_8312,N_8023,N_8181);
and U8313 (N_8313,N_8137,N_8240);
and U8314 (N_8314,N_8000,N_8116);
or U8315 (N_8315,N_8122,N_8046);
and U8316 (N_8316,N_8056,N_8215);
nor U8317 (N_8317,N_8205,N_8033);
nor U8318 (N_8318,N_8191,N_8076);
nor U8319 (N_8319,N_8184,N_8017);
nor U8320 (N_8320,N_8106,N_8047);
nor U8321 (N_8321,N_8166,N_8167);
nor U8322 (N_8322,N_8117,N_8053);
nand U8323 (N_8323,N_8149,N_8006);
nand U8324 (N_8324,N_8003,N_8086);
nor U8325 (N_8325,N_8052,N_8051);
or U8326 (N_8326,N_8015,N_8178);
or U8327 (N_8327,N_8014,N_8009);
nor U8328 (N_8328,N_8054,N_8040);
xnor U8329 (N_8329,N_8072,N_8060);
nand U8330 (N_8330,N_8142,N_8246);
or U8331 (N_8331,N_8100,N_8113);
and U8332 (N_8332,N_8182,N_8098);
nand U8333 (N_8333,N_8038,N_8144);
nand U8334 (N_8334,N_8135,N_8082);
and U8335 (N_8335,N_8083,N_8032);
nor U8336 (N_8336,N_8147,N_8041);
or U8337 (N_8337,N_8110,N_8224);
nor U8338 (N_8338,N_8227,N_8138);
xnor U8339 (N_8339,N_8238,N_8204);
nand U8340 (N_8340,N_8027,N_8232);
nand U8341 (N_8341,N_8189,N_8065);
or U8342 (N_8342,N_8234,N_8112);
nor U8343 (N_8343,N_8035,N_8109);
and U8344 (N_8344,N_8233,N_8239);
nor U8345 (N_8345,N_8133,N_8131);
and U8346 (N_8346,N_8155,N_8197);
nand U8347 (N_8347,N_8209,N_8034);
nor U8348 (N_8348,N_8102,N_8011);
and U8349 (N_8349,N_8120,N_8244);
nand U8350 (N_8350,N_8214,N_8187);
or U8351 (N_8351,N_8064,N_8146);
or U8352 (N_8352,N_8055,N_8087);
or U8353 (N_8353,N_8229,N_8070);
and U8354 (N_8354,N_8108,N_8141);
and U8355 (N_8355,N_8245,N_8140);
nor U8356 (N_8356,N_8174,N_8059);
or U8357 (N_8357,N_8004,N_8243);
nor U8358 (N_8358,N_8094,N_8103);
nor U8359 (N_8359,N_8061,N_8074);
nand U8360 (N_8360,N_8123,N_8128);
or U8361 (N_8361,N_8225,N_8150);
or U8362 (N_8362,N_8039,N_8190);
and U8363 (N_8363,N_8111,N_8194);
xnor U8364 (N_8364,N_8077,N_8096);
xnor U8365 (N_8365,N_8185,N_8031);
nand U8366 (N_8366,N_8001,N_8228);
nor U8367 (N_8367,N_8029,N_8211);
nand U8368 (N_8368,N_8157,N_8223);
nand U8369 (N_8369,N_8221,N_8012);
xor U8370 (N_8370,N_8007,N_8151);
nor U8371 (N_8371,N_8124,N_8071);
nor U8372 (N_8372,N_8134,N_8202);
nand U8373 (N_8373,N_8210,N_8177);
or U8374 (N_8374,N_8092,N_8163);
and U8375 (N_8375,N_8018,N_8055);
nand U8376 (N_8376,N_8022,N_8243);
and U8377 (N_8377,N_8092,N_8239);
nand U8378 (N_8378,N_8083,N_8038);
and U8379 (N_8379,N_8013,N_8194);
and U8380 (N_8380,N_8024,N_8142);
nor U8381 (N_8381,N_8006,N_8159);
nand U8382 (N_8382,N_8205,N_8025);
nand U8383 (N_8383,N_8050,N_8190);
nand U8384 (N_8384,N_8054,N_8031);
and U8385 (N_8385,N_8006,N_8223);
nor U8386 (N_8386,N_8008,N_8035);
nor U8387 (N_8387,N_8061,N_8116);
or U8388 (N_8388,N_8141,N_8008);
or U8389 (N_8389,N_8209,N_8175);
or U8390 (N_8390,N_8199,N_8111);
and U8391 (N_8391,N_8183,N_8000);
and U8392 (N_8392,N_8097,N_8072);
nor U8393 (N_8393,N_8197,N_8105);
and U8394 (N_8394,N_8128,N_8022);
or U8395 (N_8395,N_8012,N_8098);
and U8396 (N_8396,N_8231,N_8210);
nor U8397 (N_8397,N_8059,N_8142);
nand U8398 (N_8398,N_8248,N_8001);
nor U8399 (N_8399,N_8167,N_8087);
nand U8400 (N_8400,N_8099,N_8151);
or U8401 (N_8401,N_8054,N_8062);
nor U8402 (N_8402,N_8146,N_8224);
and U8403 (N_8403,N_8182,N_8185);
or U8404 (N_8404,N_8026,N_8216);
nor U8405 (N_8405,N_8031,N_8131);
nand U8406 (N_8406,N_8000,N_8192);
or U8407 (N_8407,N_8201,N_8193);
xnor U8408 (N_8408,N_8074,N_8175);
nand U8409 (N_8409,N_8049,N_8129);
and U8410 (N_8410,N_8168,N_8011);
nor U8411 (N_8411,N_8105,N_8183);
nor U8412 (N_8412,N_8031,N_8100);
or U8413 (N_8413,N_8179,N_8032);
or U8414 (N_8414,N_8114,N_8229);
or U8415 (N_8415,N_8014,N_8204);
and U8416 (N_8416,N_8134,N_8082);
nand U8417 (N_8417,N_8244,N_8172);
nand U8418 (N_8418,N_8199,N_8018);
nand U8419 (N_8419,N_8046,N_8127);
nand U8420 (N_8420,N_8221,N_8234);
and U8421 (N_8421,N_8010,N_8208);
nand U8422 (N_8422,N_8106,N_8186);
nand U8423 (N_8423,N_8128,N_8221);
nand U8424 (N_8424,N_8224,N_8047);
nor U8425 (N_8425,N_8097,N_8235);
nor U8426 (N_8426,N_8208,N_8246);
nor U8427 (N_8427,N_8047,N_8020);
and U8428 (N_8428,N_8235,N_8209);
nand U8429 (N_8429,N_8039,N_8177);
nor U8430 (N_8430,N_8103,N_8057);
and U8431 (N_8431,N_8149,N_8087);
nand U8432 (N_8432,N_8029,N_8223);
and U8433 (N_8433,N_8183,N_8243);
nand U8434 (N_8434,N_8118,N_8182);
nand U8435 (N_8435,N_8035,N_8019);
and U8436 (N_8436,N_8011,N_8070);
nor U8437 (N_8437,N_8236,N_8199);
nor U8438 (N_8438,N_8089,N_8245);
and U8439 (N_8439,N_8005,N_8134);
or U8440 (N_8440,N_8189,N_8139);
nand U8441 (N_8441,N_8108,N_8057);
and U8442 (N_8442,N_8220,N_8011);
nand U8443 (N_8443,N_8095,N_8239);
nor U8444 (N_8444,N_8176,N_8212);
nor U8445 (N_8445,N_8135,N_8180);
or U8446 (N_8446,N_8082,N_8233);
nand U8447 (N_8447,N_8133,N_8093);
nand U8448 (N_8448,N_8173,N_8207);
and U8449 (N_8449,N_8006,N_8158);
and U8450 (N_8450,N_8000,N_8154);
or U8451 (N_8451,N_8152,N_8201);
nor U8452 (N_8452,N_8153,N_8242);
xor U8453 (N_8453,N_8082,N_8037);
nor U8454 (N_8454,N_8173,N_8095);
and U8455 (N_8455,N_8090,N_8198);
nand U8456 (N_8456,N_8160,N_8096);
nand U8457 (N_8457,N_8116,N_8128);
and U8458 (N_8458,N_8014,N_8135);
and U8459 (N_8459,N_8210,N_8208);
or U8460 (N_8460,N_8248,N_8073);
xnor U8461 (N_8461,N_8097,N_8111);
nor U8462 (N_8462,N_8003,N_8207);
nor U8463 (N_8463,N_8233,N_8086);
or U8464 (N_8464,N_8104,N_8121);
xor U8465 (N_8465,N_8132,N_8004);
nand U8466 (N_8466,N_8201,N_8100);
nand U8467 (N_8467,N_8032,N_8128);
nor U8468 (N_8468,N_8004,N_8165);
nand U8469 (N_8469,N_8026,N_8078);
and U8470 (N_8470,N_8118,N_8084);
xnor U8471 (N_8471,N_8149,N_8068);
or U8472 (N_8472,N_8167,N_8013);
and U8473 (N_8473,N_8192,N_8127);
or U8474 (N_8474,N_8121,N_8101);
nand U8475 (N_8475,N_8067,N_8058);
or U8476 (N_8476,N_8138,N_8219);
nand U8477 (N_8477,N_8194,N_8177);
xor U8478 (N_8478,N_8103,N_8213);
nand U8479 (N_8479,N_8162,N_8104);
or U8480 (N_8480,N_8199,N_8225);
nand U8481 (N_8481,N_8204,N_8088);
and U8482 (N_8482,N_8107,N_8027);
or U8483 (N_8483,N_8004,N_8139);
or U8484 (N_8484,N_8173,N_8012);
or U8485 (N_8485,N_8076,N_8081);
nor U8486 (N_8486,N_8194,N_8130);
nand U8487 (N_8487,N_8123,N_8011);
or U8488 (N_8488,N_8016,N_8190);
and U8489 (N_8489,N_8130,N_8140);
or U8490 (N_8490,N_8009,N_8115);
nor U8491 (N_8491,N_8006,N_8032);
or U8492 (N_8492,N_8067,N_8235);
and U8493 (N_8493,N_8038,N_8183);
or U8494 (N_8494,N_8018,N_8060);
nand U8495 (N_8495,N_8214,N_8235);
and U8496 (N_8496,N_8015,N_8122);
nor U8497 (N_8497,N_8100,N_8004);
nor U8498 (N_8498,N_8219,N_8207);
nor U8499 (N_8499,N_8036,N_8233);
nand U8500 (N_8500,N_8364,N_8273);
nor U8501 (N_8501,N_8295,N_8386);
xnor U8502 (N_8502,N_8382,N_8255);
nand U8503 (N_8503,N_8272,N_8318);
and U8504 (N_8504,N_8487,N_8279);
nor U8505 (N_8505,N_8323,N_8427);
or U8506 (N_8506,N_8300,N_8443);
nor U8507 (N_8507,N_8349,N_8311);
nor U8508 (N_8508,N_8458,N_8337);
and U8509 (N_8509,N_8481,N_8282);
nor U8510 (N_8510,N_8438,N_8319);
and U8511 (N_8511,N_8355,N_8285);
and U8512 (N_8512,N_8309,N_8470);
xor U8513 (N_8513,N_8302,N_8440);
nor U8514 (N_8514,N_8299,N_8499);
or U8515 (N_8515,N_8368,N_8340);
or U8516 (N_8516,N_8320,N_8265);
nand U8517 (N_8517,N_8287,N_8415);
nor U8518 (N_8518,N_8426,N_8419);
or U8519 (N_8519,N_8479,N_8322);
nand U8520 (N_8520,N_8478,N_8348);
nand U8521 (N_8521,N_8377,N_8448);
nor U8522 (N_8522,N_8412,N_8310);
nor U8523 (N_8523,N_8293,N_8359);
and U8524 (N_8524,N_8421,N_8476);
or U8525 (N_8525,N_8338,N_8290);
or U8526 (N_8526,N_8334,N_8308);
or U8527 (N_8527,N_8395,N_8417);
nand U8528 (N_8528,N_8473,N_8294);
nor U8529 (N_8529,N_8370,N_8406);
xor U8530 (N_8530,N_8456,N_8469);
nand U8531 (N_8531,N_8393,N_8463);
or U8532 (N_8532,N_8498,N_8266);
or U8533 (N_8533,N_8327,N_8388);
nor U8534 (N_8534,N_8490,N_8314);
and U8535 (N_8535,N_8392,N_8271);
nor U8536 (N_8536,N_8489,N_8468);
or U8537 (N_8537,N_8485,N_8466);
nor U8538 (N_8538,N_8374,N_8332);
nor U8539 (N_8539,N_8464,N_8398);
and U8540 (N_8540,N_8407,N_8424);
and U8541 (N_8541,N_8445,N_8253);
nand U8542 (N_8542,N_8455,N_8250);
nand U8543 (N_8543,N_8353,N_8409);
and U8544 (N_8544,N_8436,N_8371);
nor U8545 (N_8545,N_8408,N_8281);
nor U8546 (N_8546,N_8423,N_8467);
nor U8547 (N_8547,N_8321,N_8275);
nor U8548 (N_8548,N_8383,N_8335);
xor U8549 (N_8549,N_8399,N_8343);
nand U8550 (N_8550,N_8461,N_8416);
nand U8551 (N_8551,N_8256,N_8429);
nor U8552 (N_8552,N_8397,N_8339);
nor U8553 (N_8553,N_8475,N_8284);
xnor U8554 (N_8554,N_8330,N_8352);
nor U8555 (N_8555,N_8252,N_8439);
nand U8556 (N_8556,N_8306,N_8486);
nor U8557 (N_8557,N_8431,N_8373);
or U8558 (N_8558,N_8301,N_8432);
and U8559 (N_8559,N_8278,N_8303);
and U8560 (N_8560,N_8442,N_8345);
or U8561 (N_8561,N_8283,N_8401);
nand U8562 (N_8562,N_8292,N_8454);
nor U8563 (N_8563,N_8262,N_8474);
xnor U8564 (N_8564,N_8304,N_8385);
nor U8565 (N_8565,N_8280,N_8405);
nor U8566 (N_8566,N_8402,N_8488);
or U8567 (N_8567,N_8333,N_8298);
and U8568 (N_8568,N_8259,N_8324);
and U8569 (N_8569,N_8483,N_8325);
nand U8570 (N_8570,N_8369,N_8434);
nor U8571 (N_8571,N_8261,N_8257);
nand U8572 (N_8572,N_8270,N_8317);
or U8573 (N_8573,N_8471,N_8346);
xnor U8574 (N_8574,N_8449,N_8496);
nor U8575 (N_8575,N_8307,N_8326);
nand U8576 (N_8576,N_8495,N_8372);
or U8577 (N_8577,N_8267,N_8404);
and U8578 (N_8578,N_8376,N_8358);
nor U8579 (N_8579,N_8493,N_8251);
or U8580 (N_8580,N_8465,N_8389);
nor U8581 (N_8581,N_8258,N_8492);
or U8582 (N_8582,N_8296,N_8384);
or U8583 (N_8583,N_8363,N_8460);
nor U8584 (N_8584,N_8354,N_8452);
and U8585 (N_8585,N_8396,N_8297);
and U8586 (N_8586,N_8457,N_8313);
nand U8587 (N_8587,N_8269,N_8291);
nand U8588 (N_8588,N_8444,N_8263);
xnor U8589 (N_8589,N_8472,N_8453);
or U8590 (N_8590,N_8380,N_8450);
nand U8591 (N_8591,N_8400,N_8446);
nand U8592 (N_8592,N_8441,N_8276);
or U8593 (N_8593,N_8379,N_8433);
nor U8594 (N_8594,N_8361,N_8347);
or U8595 (N_8595,N_8418,N_8288);
or U8596 (N_8596,N_8328,N_8494);
nand U8597 (N_8597,N_8430,N_8437);
nor U8598 (N_8598,N_8362,N_8435);
nand U8599 (N_8599,N_8484,N_8316);
nand U8600 (N_8600,N_8286,N_8447);
nor U8601 (N_8601,N_8274,N_8420);
nor U8602 (N_8602,N_8381,N_8342);
nand U8603 (N_8603,N_8366,N_8480);
and U8604 (N_8604,N_8289,N_8350);
nor U8605 (N_8605,N_8344,N_8390);
and U8606 (N_8606,N_8315,N_8365);
nor U8607 (N_8607,N_8387,N_8428);
and U8608 (N_8608,N_8394,N_8391);
nand U8609 (N_8609,N_8477,N_8367);
or U8610 (N_8610,N_8268,N_8360);
nand U8611 (N_8611,N_8497,N_8277);
and U8612 (N_8612,N_8425,N_8336);
nor U8613 (N_8613,N_8254,N_8329);
and U8614 (N_8614,N_8410,N_8357);
nand U8615 (N_8615,N_8331,N_8403);
nor U8616 (N_8616,N_8378,N_8413);
and U8617 (N_8617,N_8414,N_8351);
and U8618 (N_8618,N_8356,N_8305);
nand U8619 (N_8619,N_8451,N_8462);
or U8620 (N_8620,N_8312,N_8411);
xnor U8621 (N_8621,N_8341,N_8491);
nor U8622 (N_8622,N_8375,N_8459);
nand U8623 (N_8623,N_8260,N_8264);
nand U8624 (N_8624,N_8422,N_8482);
or U8625 (N_8625,N_8321,N_8313);
and U8626 (N_8626,N_8251,N_8255);
or U8627 (N_8627,N_8369,N_8295);
or U8628 (N_8628,N_8356,N_8307);
or U8629 (N_8629,N_8307,N_8281);
nor U8630 (N_8630,N_8445,N_8497);
nor U8631 (N_8631,N_8465,N_8365);
and U8632 (N_8632,N_8293,N_8445);
or U8633 (N_8633,N_8429,N_8485);
nor U8634 (N_8634,N_8448,N_8499);
nand U8635 (N_8635,N_8429,N_8455);
nand U8636 (N_8636,N_8470,N_8448);
and U8637 (N_8637,N_8307,N_8304);
xor U8638 (N_8638,N_8486,N_8484);
nand U8639 (N_8639,N_8368,N_8456);
nand U8640 (N_8640,N_8347,N_8376);
or U8641 (N_8641,N_8448,N_8351);
nand U8642 (N_8642,N_8489,N_8417);
nor U8643 (N_8643,N_8445,N_8465);
nand U8644 (N_8644,N_8315,N_8386);
or U8645 (N_8645,N_8250,N_8275);
or U8646 (N_8646,N_8495,N_8361);
nand U8647 (N_8647,N_8498,N_8497);
nor U8648 (N_8648,N_8406,N_8439);
and U8649 (N_8649,N_8368,N_8337);
nor U8650 (N_8650,N_8466,N_8293);
nor U8651 (N_8651,N_8406,N_8317);
or U8652 (N_8652,N_8303,N_8446);
xor U8653 (N_8653,N_8404,N_8393);
nor U8654 (N_8654,N_8435,N_8265);
and U8655 (N_8655,N_8349,N_8292);
and U8656 (N_8656,N_8314,N_8376);
and U8657 (N_8657,N_8492,N_8332);
nor U8658 (N_8658,N_8338,N_8431);
nand U8659 (N_8659,N_8430,N_8326);
nand U8660 (N_8660,N_8358,N_8374);
nand U8661 (N_8661,N_8473,N_8382);
nand U8662 (N_8662,N_8420,N_8409);
and U8663 (N_8663,N_8405,N_8266);
nor U8664 (N_8664,N_8460,N_8324);
nand U8665 (N_8665,N_8400,N_8454);
and U8666 (N_8666,N_8342,N_8334);
xor U8667 (N_8667,N_8294,N_8477);
nor U8668 (N_8668,N_8445,N_8480);
and U8669 (N_8669,N_8406,N_8473);
or U8670 (N_8670,N_8254,N_8430);
or U8671 (N_8671,N_8268,N_8321);
or U8672 (N_8672,N_8314,N_8469);
nand U8673 (N_8673,N_8302,N_8265);
and U8674 (N_8674,N_8431,N_8415);
and U8675 (N_8675,N_8403,N_8361);
nor U8676 (N_8676,N_8286,N_8275);
nand U8677 (N_8677,N_8323,N_8258);
nand U8678 (N_8678,N_8376,N_8355);
xnor U8679 (N_8679,N_8434,N_8413);
nor U8680 (N_8680,N_8468,N_8311);
and U8681 (N_8681,N_8466,N_8358);
or U8682 (N_8682,N_8261,N_8390);
and U8683 (N_8683,N_8372,N_8310);
and U8684 (N_8684,N_8475,N_8461);
nor U8685 (N_8685,N_8312,N_8306);
nor U8686 (N_8686,N_8372,N_8323);
and U8687 (N_8687,N_8373,N_8366);
or U8688 (N_8688,N_8310,N_8370);
nand U8689 (N_8689,N_8411,N_8433);
nor U8690 (N_8690,N_8269,N_8261);
nand U8691 (N_8691,N_8435,N_8406);
nor U8692 (N_8692,N_8346,N_8408);
and U8693 (N_8693,N_8411,N_8322);
and U8694 (N_8694,N_8384,N_8276);
nor U8695 (N_8695,N_8255,N_8306);
nor U8696 (N_8696,N_8321,N_8395);
and U8697 (N_8697,N_8266,N_8494);
nor U8698 (N_8698,N_8358,N_8441);
nand U8699 (N_8699,N_8427,N_8485);
and U8700 (N_8700,N_8402,N_8336);
nor U8701 (N_8701,N_8415,N_8450);
and U8702 (N_8702,N_8381,N_8258);
nand U8703 (N_8703,N_8467,N_8293);
and U8704 (N_8704,N_8411,N_8329);
or U8705 (N_8705,N_8286,N_8418);
nand U8706 (N_8706,N_8401,N_8477);
nand U8707 (N_8707,N_8250,N_8251);
or U8708 (N_8708,N_8355,N_8490);
or U8709 (N_8709,N_8416,N_8356);
nor U8710 (N_8710,N_8427,N_8307);
nor U8711 (N_8711,N_8479,N_8452);
nand U8712 (N_8712,N_8393,N_8277);
nand U8713 (N_8713,N_8419,N_8260);
and U8714 (N_8714,N_8251,N_8468);
nand U8715 (N_8715,N_8415,N_8262);
or U8716 (N_8716,N_8363,N_8391);
xnor U8717 (N_8717,N_8406,N_8485);
and U8718 (N_8718,N_8467,N_8299);
and U8719 (N_8719,N_8358,N_8316);
nor U8720 (N_8720,N_8335,N_8450);
nand U8721 (N_8721,N_8385,N_8325);
and U8722 (N_8722,N_8360,N_8438);
xnor U8723 (N_8723,N_8273,N_8480);
or U8724 (N_8724,N_8433,N_8294);
nor U8725 (N_8725,N_8464,N_8293);
nand U8726 (N_8726,N_8354,N_8417);
and U8727 (N_8727,N_8321,N_8369);
nand U8728 (N_8728,N_8450,N_8403);
or U8729 (N_8729,N_8434,N_8366);
nand U8730 (N_8730,N_8308,N_8408);
nor U8731 (N_8731,N_8420,N_8445);
or U8732 (N_8732,N_8474,N_8269);
xor U8733 (N_8733,N_8455,N_8289);
nand U8734 (N_8734,N_8434,N_8339);
nand U8735 (N_8735,N_8324,N_8439);
xor U8736 (N_8736,N_8277,N_8320);
and U8737 (N_8737,N_8282,N_8287);
nand U8738 (N_8738,N_8497,N_8258);
nand U8739 (N_8739,N_8269,N_8317);
and U8740 (N_8740,N_8273,N_8430);
nand U8741 (N_8741,N_8406,N_8267);
or U8742 (N_8742,N_8473,N_8495);
nor U8743 (N_8743,N_8253,N_8263);
and U8744 (N_8744,N_8498,N_8434);
and U8745 (N_8745,N_8402,N_8399);
xnor U8746 (N_8746,N_8479,N_8459);
nor U8747 (N_8747,N_8371,N_8349);
nor U8748 (N_8748,N_8441,N_8345);
or U8749 (N_8749,N_8388,N_8322);
nor U8750 (N_8750,N_8712,N_8544);
or U8751 (N_8751,N_8651,N_8565);
xnor U8752 (N_8752,N_8692,N_8566);
xor U8753 (N_8753,N_8625,N_8581);
and U8754 (N_8754,N_8593,N_8556);
and U8755 (N_8755,N_8693,N_8512);
xor U8756 (N_8756,N_8539,N_8570);
nand U8757 (N_8757,N_8584,N_8740);
and U8758 (N_8758,N_8647,N_8618);
nor U8759 (N_8759,N_8559,N_8578);
nand U8760 (N_8760,N_8634,N_8612);
nor U8761 (N_8761,N_8610,N_8645);
nand U8762 (N_8762,N_8734,N_8710);
and U8763 (N_8763,N_8600,N_8542);
nor U8764 (N_8764,N_8528,N_8719);
or U8765 (N_8765,N_8702,N_8705);
nor U8766 (N_8766,N_8553,N_8687);
or U8767 (N_8767,N_8621,N_8525);
nand U8768 (N_8768,N_8518,N_8511);
nor U8769 (N_8769,N_8502,N_8686);
nor U8770 (N_8770,N_8604,N_8738);
nor U8771 (N_8771,N_8530,N_8603);
or U8772 (N_8772,N_8642,N_8620);
nand U8773 (N_8773,N_8709,N_8665);
or U8774 (N_8774,N_8688,N_8713);
or U8775 (N_8775,N_8558,N_8737);
or U8776 (N_8776,N_8636,N_8663);
and U8777 (N_8777,N_8729,N_8562);
nand U8778 (N_8778,N_8617,N_8653);
nor U8779 (N_8779,N_8522,N_8633);
or U8780 (N_8780,N_8624,N_8704);
nor U8781 (N_8781,N_8657,N_8671);
nor U8782 (N_8782,N_8601,N_8700);
nand U8783 (N_8783,N_8561,N_8668);
and U8784 (N_8784,N_8715,N_8635);
nand U8785 (N_8785,N_8745,N_8598);
or U8786 (N_8786,N_8726,N_8546);
or U8787 (N_8787,N_8507,N_8649);
or U8788 (N_8788,N_8652,N_8718);
xor U8789 (N_8789,N_8732,N_8733);
nor U8790 (N_8790,N_8520,N_8646);
nor U8791 (N_8791,N_8523,N_8536);
and U8792 (N_8792,N_8670,N_8516);
xor U8793 (N_8793,N_8676,N_8583);
or U8794 (N_8794,N_8680,N_8567);
and U8795 (N_8795,N_8748,N_8637);
xor U8796 (N_8796,N_8622,N_8648);
and U8797 (N_8797,N_8557,N_8747);
or U8798 (N_8798,N_8678,N_8717);
nor U8799 (N_8799,N_8681,N_8563);
nand U8800 (N_8800,N_8661,N_8723);
and U8801 (N_8801,N_8694,N_8576);
and U8802 (N_8802,N_8607,N_8725);
nor U8803 (N_8803,N_8508,N_8735);
nand U8804 (N_8804,N_8742,N_8540);
nand U8805 (N_8805,N_8632,N_8714);
nand U8806 (N_8806,N_8506,N_8672);
and U8807 (N_8807,N_8741,N_8724);
nor U8808 (N_8808,N_8691,N_8585);
or U8809 (N_8809,N_8572,N_8675);
and U8810 (N_8810,N_8743,N_8664);
or U8811 (N_8811,N_8623,N_8543);
or U8812 (N_8812,N_8510,N_8527);
or U8813 (N_8813,N_8500,N_8613);
nand U8814 (N_8814,N_8602,N_8673);
xor U8815 (N_8815,N_8614,N_8596);
and U8816 (N_8816,N_8524,N_8669);
and U8817 (N_8817,N_8504,N_8739);
and U8818 (N_8818,N_8655,N_8582);
nand U8819 (N_8819,N_8533,N_8722);
or U8820 (N_8820,N_8644,N_8609);
nand U8821 (N_8821,N_8611,N_8592);
or U8822 (N_8822,N_8594,N_8608);
or U8823 (N_8823,N_8656,N_8552);
nand U8824 (N_8824,N_8630,N_8716);
or U8825 (N_8825,N_8616,N_8654);
and U8826 (N_8826,N_8514,N_8677);
nand U8827 (N_8827,N_8509,N_8550);
nand U8828 (N_8828,N_8631,N_8545);
nand U8829 (N_8829,N_8568,N_8515);
nand U8830 (N_8830,N_8554,N_8549);
or U8831 (N_8831,N_8564,N_8590);
nor U8832 (N_8832,N_8721,N_8685);
and U8833 (N_8833,N_8501,N_8683);
or U8834 (N_8834,N_8597,N_8736);
or U8835 (N_8835,N_8503,N_8587);
and U8836 (N_8836,N_8571,N_8526);
or U8837 (N_8837,N_8706,N_8577);
and U8838 (N_8838,N_8701,N_8684);
and U8839 (N_8839,N_8679,N_8555);
xor U8840 (N_8840,N_8708,N_8731);
nor U8841 (N_8841,N_8696,N_8730);
or U8842 (N_8842,N_8605,N_8746);
nand U8843 (N_8843,N_8575,N_8643);
nand U8844 (N_8844,N_8529,N_8521);
or U8845 (N_8845,N_8551,N_8660);
xnor U8846 (N_8846,N_8547,N_8727);
nor U8847 (N_8847,N_8695,N_8586);
or U8848 (N_8848,N_8619,N_8707);
and U8849 (N_8849,N_8532,N_8749);
nand U8850 (N_8850,N_8667,N_8599);
nand U8851 (N_8851,N_8689,N_8541);
nor U8852 (N_8852,N_8690,N_8534);
nand U8853 (N_8853,N_8535,N_8574);
or U8854 (N_8854,N_8641,N_8560);
and U8855 (N_8855,N_8519,N_8531);
xnor U8856 (N_8856,N_8711,N_8674);
xor U8857 (N_8857,N_8517,N_8629);
nor U8858 (N_8858,N_8589,N_8666);
xor U8859 (N_8859,N_8628,N_8569);
or U8860 (N_8860,N_8638,N_8697);
nand U8861 (N_8861,N_8595,N_8699);
and U8862 (N_8862,N_8580,N_8744);
nor U8863 (N_8863,N_8573,N_8682);
nor U8864 (N_8864,N_8591,N_8658);
nand U8865 (N_8865,N_8627,N_8537);
and U8866 (N_8866,N_8639,N_8588);
nor U8867 (N_8867,N_8640,N_8615);
nand U8868 (N_8868,N_8720,N_8548);
and U8869 (N_8869,N_8606,N_8662);
and U8870 (N_8870,N_8659,N_8728);
and U8871 (N_8871,N_8538,N_8698);
or U8872 (N_8872,N_8505,N_8703);
and U8873 (N_8873,N_8513,N_8626);
and U8874 (N_8874,N_8579,N_8650);
and U8875 (N_8875,N_8668,N_8655);
nor U8876 (N_8876,N_8540,N_8571);
nand U8877 (N_8877,N_8562,N_8680);
nor U8878 (N_8878,N_8724,N_8700);
nor U8879 (N_8879,N_8665,N_8625);
xnor U8880 (N_8880,N_8622,N_8663);
or U8881 (N_8881,N_8597,N_8556);
xnor U8882 (N_8882,N_8607,N_8717);
or U8883 (N_8883,N_8678,N_8550);
nand U8884 (N_8884,N_8604,N_8535);
or U8885 (N_8885,N_8572,N_8729);
or U8886 (N_8886,N_8636,N_8513);
and U8887 (N_8887,N_8631,N_8715);
or U8888 (N_8888,N_8748,N_8633);
nand U8889 (N_8889,N_8630,N_8664);
and U8890 (N_8890,N_8565,N_8500);
or U8891 (N_8891,N_8685,N_8694);
or U8892 (N_8892,N_8541,N_8634);
nand U8893 (N_8893,N_8527,N_8592);
xor U8894 (N_8894,N_8514,N_8696);
xnor U8895 (N_8895,N_8665,N_8635);
and U8896 (N_8896,N_8562,N_8535);
nand U8897 (N_8897,N_8722,N_8598);
and U8898 (N_8898,N_8518,N_8525);
nand U8899 (N_8899,N_8591,N_8661);
or U8900 (N_8900,N_8550,N_8567);
nand U8901 (N_8901,N_8620,N_8526);
nor U8902 (N_8902,N_8570,N_8699);
and U8903 (N_8903,N_8698,N_8562);
or U8904 (N_8904,N_8603,N_8536);
nor U8905 (N_8905,N_8734,N_8612);
xnor U8906 (N_8906,N_8714,N_8687);
nor U8907 (N_8907,N_8623,N_8524);
or U8908 (N_8908,N_8574,N_8637);
nand U8909 (N_8909,N_8535,N_8634);
nor U8910 (N_8910,N_8514,N_8527);
nor U8911 (N_8911,N_8552,N_8745);
nor U8912 (N_8912,N_8731,N_8606);
nor U8913 (N_8913,N_8639,N_8607);
and U8914 (N_8914,N_8682,N_8641);
xnor U8915 (N_8915,N_8547,N_8604);
and U8916 (N_8916,N_8679,N_8514);
or U8917 (N_8917,N_8608,N_8528);
nand U8918 (N_8918,N_8514,N_8572);
nand U8919 (N_8919,N_8722,N_8727);
nor U8920 (N_8920,N_8561,N_8672);
nor U8921 (N_8921,N_8520,N_8509);
or U8922 (N_8922,N_8692,N_8567);
nand U8923 (N_8923,N_8526,N_8527);
or U8924 (N_8924,N_8594,N_8553);
and U8925 (N_8925,N_8683,N_8642);
nor U8926 (N_8926,N_8711,N_8740);
or U8927 (N_8927,N_8611,N_8502);
or U8928 (N_8928,N_8584,N_8557);
nand U8929 (N_8929,N_8539,N_8701);
and U8930 (N_8930,N_8629,N_8612);
and U8931 (N_8931,N_8602,N_8601);
nor U8932 (N_8932,N_8608,N_8705);
nand U8933 (N_8933,N_8583,N_8514);
xnor U8934 (N_8934,N_8615,N_8716);
nand U8935 (N_8935,N_8596,N_8705);
and U8936 (N_8936,N_8574,N_8689);
and U8937 (N_8937,N_8598,N_8560);
nor U8938 (N_8938,N_8702,N_8621);
and U8939 (N_8939,N_8694,N_8615);
nor U8940 (N_8940,N_8610,N_8562);
and U8941 (N_8941,N_8724,N_8656);
or U8942 (N_8942,N_8656,N_8517);
nor U8943 (N_8943,N_8657,N_8749);
xnor U8944 (N_8944,N_8507,N_8622);
and U8945 (N_8945,N_8632,N_8607);
nor U8946 (N_8946,N_8565,N_8645);
nand U8947 (N_8947,N_8702,N_8597);
xnor U8948 (N_8948,N_8698,N_8513);
nand U8949 (N_8949,N_8749,N_8586);
and U8950 (N_8950,N_8518,N_8575);
nand U8951 (N_8951,N_8715,N_8588);
or U8952 (N_8952,N_8636,N_8628);
nor U8953 (N_8953,N_8651,N_8691);
nand U8954 (N_8954,N_8582,N_8669);
or U8955 (N_8955,N_8558,N_8665);
and U8956 (N_8956,N_8706,N_8734);
nand U8957 (N_8957,N_8618,N_8581);
nor U8958 (N_8958,N_8629,N_8627);
nor U8959 (N_8959,N_8737,N_8684);
and U8960 (N_8960,N_8552,N_8586);
or U8961 (N_8961,N_8582,N_8574);
nor U8962 (N_8962,N_8620,N_8579);
or U8963 (N_8963,N_8749,N_8703);
xnor U8964 (N_8964,N_8718,N_8548);
and U8965 (N_8965,N_8565,N_8637);
nor U8966 (N_8966,N_8711,N_8533);
nor U8967 (N_8967,N_8561,N_8602);
or U8968 (N_8968,N_8510,N_8719);
or U8969 (N_8969,N_8510,N_8558);
and U8970 (N_8970,N_8694,N_8628);
nor U8971 (N_8971,N_8684,N_8550);
or U8972 (N_8972,N_8574,N_8703);
and U8973 (N_8973,N_8682,N_8686);
nor U8974 (N_8974,N_8642,N_8530);
nand U8975 (N_8975,N_8672,N_8705);
xnor U8976 (N_8976,N_8706,N_8521);
and U8977 (N_8977,N_8649,N_8746);
or U8978 (N_8978,N_8660,N_8714);
nor U8979 (N_8979,N_8602,N_8699);
nor U8980 (N_8980,N_8554,N_8737);
nor U8981 (N_8981,N_8723,N_8553);
nand U8982 (N_8982,N_8677,N_8504);
or U8983 (N_8983,N_8685,N_8676);
xor U8984 (N_8984,N_8723,N_8527);
nand U8985 (N_8985,N_8680,N_8595);
and U8986 (N_8986,N_8508,N_8603);
nor U8987 (N_8987,N_8748,N_8630);
xor U8988 (N_8988,N_8678,N_8628);
xor U8989 (N_8989,N_8649,N_8713);
and U8990 (N_8990,N_8628,N_8713);
nor U8991 (N_8991,N_8701,N_8594);
xnor U8992 (N_8992,N_8530,N_8677);
nand U8993 (N_8993,N_8511,N_8598);
nand U8994 (N_8994,N_8709,N_8646);
nand U8995 (N_8995,N_8675,N_8548);
nand U8996 (N_8996,N_8640,N_8638);
nor U8997 (N_8997,N_8639,N_8670);
or U8998 (N_8998,N_8615,N_8515);
and U8999 (N_8999,N_8701,N_8622);
nor U9000 (N_9000,N_8966,N_8878);
nand U9001 (N_9001,N_8852,N_8882);
or U9002 (N_9002,N_8861,N_8762);
or U9003 (N_9003,N_8783,N_8890);
or U9004 (N_9004,N_8960,N_8871);
or U9005 (N_9005,N_8795,N_8886);
nand U9006 (N_9006,N_8989,N_8856);
xor U9007 (N_9007,N_8912,N_8991);
and U9008 (N_9008,N_8793,N_8962);
or U9009 (N_9009,N_8864,N_8953);
nand U9010 (N_9010,N_8946,N_8927);
or U9011 (N_9011,N_8846,N_8821);
xor U9012 (N_9012,N_8870,N_8829);
and U9013 (N_9013,N_8761,N_8893);
or U9014 (N_9014,N_8913,N_8948);
nand U9015 (N_9015,N_8844,N_8802);
and U9016 (N_9016,N_8947,N_8919);
and U9017 (N_9017,N_8756,N_8869);
and U9018 (N_9018,N_8961,N_8866);
or U9019 (N_9019,N_8796,N_8797);
nand U9020 (N_9020,N_8954,N_8930);
nand U9021 (N_9021,N_8977,N_8895);
nand U9022 (N_9022,N_8828,N_8941);
or U9023 (N_9023,N_8790,N_8775);
nand U9024 (N_9024,N_8767,N_8901);
and U9025 (N_9025,N_8957,N_8759);
nand U9026 (N_9026,N_8970,N_8965);
nand U9027 (N_9027,N_8809,N_8786);
nor U9028 (N_9028,N_8938,N_8838);
xor U9029 (N_9029,N_8815,N_8848);
nor U9030 (N_9030,N_8928,N_8891);
and U9031 (N_9031,N_8751,N_8936);
nand U9032 (N_9032,N_8900,N_8906);
or U9033 (N_9033,N_8776,N_8841);
nand U9034 (N_9034,N_8868,N_8950);
and U9035 (N_9035,N_8914,N_8998);
and U9036 (N_9036,N_8874,N_8972);
nand U9037 (N_9037,N_8757,N_8984);
nand U9038 (N_9038,N_8782,N_8896);
or U9039 (N_9039,N_8842,N_8955);
xnor U9040 (N_9040,N_8839,N_8902);
nor U9041 (N_9041,N_8899,N_8820);
or U9042 (N_9042,N_8787,N_8911);
nand U9043 (N_9043,N_8804,N_8924);
nor U9044 (N_9044,N_8781,N_8840);
nor U9045 (N_9045,N_8898,N_8826);
or U9046 (N_9046,N_8794,N_8929);
nand U9047 (N_9047,N_8812,N_8753);
and U9048 (N_9048,N_8905,N_8925);
xor U9049 (N_9049,N_8758,N_8850);
and U9050 (N_9050,N_8872,N_8892);
nand U9051 (N_9051,N_8923,N_8752);
and U9052 (N_9052,N_8884,N_8830);
xor U9053 (N_9053,N_8897,N_8979);
nor U9054 (N_9054,N_8949,N_8849);
nor U9055 (N_9055,N_8785,N_8771);
or U9056 (N_9056,N_8940,N_8888);
and U9057 (N_9057,N_8769,N_8855);
or U9058 (N_9058,N_8932,N_8779);
or U9059 (N_9059,N_8833,N_8974);
and U9060 (N_9060,N_8880,N_8944);
nor U9061 (N_9061,N_8875,N_8881);
and U9062 (N_9062,N_8780,N_8937);
nor U9063 (N_9063,N_8860,N_8964);
xnor U9064 (N_9064,N_8766,N_8836);
nand U9065 (N_9065,N_8920,N_8770);
or U9066 (N_9066,N_8777,N_8963);
nor U9067 (N_9067,N_8877,N_8784);
or U9068 (N_9068,N_8969,N_8847);
nor U9069 (N_9069,N_8917,N_8851);
and U9070 (N_9070,N_8992,N_8800);
nor U9071 (N_9071,N_8813,N_8943);
or U9072 (N_9072,N_8831,N_8889);
and U9073 (N_9073,N_8755,N_8824);
nand U9074 (N_9074,N_8985,N_8987);
and U9075 (N_9075,N_8993,N_8810);
or U9076 (N_9076,N_8816,N_8971);
nand U9077 (N_9077,N_8980,N_8910);
or U9078 (N_9078,N_8825,N_8883);
and U9079 (N_9079,N_8933,N_8894);
nor U9080 (N_9080,N_8967,N_8837);
xor U9081 (N_9081,N_8959,N_8976);
nand U9082 (N_9082,N_8981,N_8939);
or U9083 (N_9083,N_8773,N_8935);
and U9084 (N_9084,N_8922,N_8999);
and U9085 (N_9085,N_8931,N_8863);
and U9086 (N_9086,N_8982,N_8885);
xnor U9087 (N_9087,N_8834,N_8791);
or U9088 (N_9088,N_8952,N_8801);
or U9089 (N_9089,N_8814,N_8988);
nand U9090 (N_9090,N_8975,N_8857);
nor U9091 (N_9091,N_8843,N_8990);
nor U9092 (N_9092,N_8763,N_8835);
or U9093 (N_9093,N_8956,N_8807);
nand U9094 (N_9094,N_8754,N_8978);
nand U9095 (N_9095,N_8853,N_8798);
or U9096 (N_9096,N_8926,N_8865);
and U9097 (N_9097,N_8958,N_8750);
xor U9098 (N_9098,N_8803,N_8778);
or U9099 (N_9099,N_8879,N_8768);
or U9100 (N_9100,N_8873,N_8887);
xor U9101 (N_9101,N_8818,N_8921);
nand U9102 (N_9102,N_8942,N_8792);
and U9103 (N_9103,N_8845,N_8822);
nand U9104 (N_9104,N_8907,N_8934);
xor U9105 (N_9105,N_8823,N_8862);
and U9106 (N_9106,N_8983,N_8774);
or U9107 (N_9107,N_8916,N_8817);
and U9108 (N_9108,N_8806,N_8908);
and U9109 (N_9109,N_8997,N_8772);
nand U9110 (N_9110,N_8765,N_8789);
or U9111 (N_9111,N_8805,N_8996);
nand U9112 (N_9112,N_8968,N_8904);
or U9113 (N_9113,N_8827,N_8951);
nor U9114 (N_9114,N_8808,N_8915);
xor U9115 (N_9115,N_8858,N_8945);
or U9116 (N_9116,N_8986,N_8764);
and U9117 (N_9117,N_8867,N_8918);
nand U9118 (N_9118,N_8859,N_8819);
or U9119 (N_9119,N_8854,N_8876);
and U9120 (N_9120,N_8832,N_8994);
nand U9121 (N_9121,N_8760,N_8811);
nor U9122 (N_9122,N_8909,N_8903);
nand U9123 (N_9123,N_8995,N_8799);
and U9124 (N_9124,N_8973,N_8788);
nor U9125 (N_9125,N_8923,N_8849);
nor U9126 (N_9126,N_8848,N_8757);
nand U9127 (N_9127,N_8903,N_8860);
or U9128 (N_9128,N_8758,N_8796);
xor U9129 (N_9129,N_8923,N_8945);
or U9130 (N_9130,N_8979,N_8820);
nand U9131 (N_9131,N_8877,N_8840);
nand U9132 (N_9132,N_8974,N_8814);
and U9133 (N_9133,N_8813,N_8773);
or U9134 (N_9134,N_8838,N_8952);
and U9135 (N_9135,N_8889,N_8782);
and U9136 (N_9136,N_8931,N_8836);
nand U9137 (N_9137,N_8937,N_8963);
xnor U9138 (N_9138,N_8843,N_8893);
nand U9139 (N_9139,N_8849,N_8761);
nor U9140 (N_9140,N_8936,N_8799);
and U9141 (N_9141,N_8940,N_8923);
or U9142 (N_9142,N_8781,N_8933);
and U9143 (N_9143,N_8766,N_8803);
or U9144 (N_9144,N_8960,N_8956);
nand U9145 (N_9145,N_8784,N_8896);
nand U9146 (N_9146,N_8791,N_8997);
and U9147 (N_9147,N_8929,N_8797);
nand U9148 (N_9148,N_8785,N_8930);
and U9149 (N_9149,N_8821,N_8763);
or U9150 (N_9150,N_8894,N_8795);
or U9151 (N_9151,N_8988,N_8927);
and U9152 (N_9152,N_8805,N_8882);
or U9153 (N_9153,N_8886,N_8763);
and U9154 (N_9154,N_8973,N_8772);
nand U9155 (N_9155,N_8835,N_8841);
or U9156 (N_9156,N_8776,N_8910);
and U9157 (N_9157,N_8944,N_8963);
nand U9158 (N_9158,N_8906,N_8804);
and U9159 (N_9159,N_8785,N_8855);
nand U9160 (N_9160,N_8784,N_8797);
nor U9161 (N_9161,N_8906,N_8887);
nand U9162 (N_9162,N_8920,N_8945);
and U9163 (N_9163,N_8871,N_8938);
and U9164 (N_9164,N_8908,N_8798);
nor U9165 (N_9165,N_8936,N_8803);
and U9166 (N_9166,N_8983,N_8956);
xor U9167 (N_9167,N_8898,N_8780);
nor U9168 (N_9168,N_8807,N_8883);
xnor U9169 (N_9169,N_8929,N_8815);
nand U9170 (N_9170,N_8829,N_8942);
or U9171 (N_9171,N_8887,N_8942);
nor U9172 (N_9172,N_8879,N_8858);
or U9173 (N_9173,N_8791,N_8953);
and U9174 (N_9174,N_8905,N_8783);
and U9175 (N_9175,N_8773,N_8889);
xor U9176 (N_9176,N_8907,N_8752);
and U9177 (N_9177,N_8820,N_8909);
and U9178 (N_9178,N_8907,N_8915);
nor U9179 (N_9179,N_8869,N_8960);
nor U9180 (N_9180,N_8987,N_8799);
nor U9181 (N_9181,N_8889,N_8937);
or U9182 (N_9182,N_8957,N_8813);
and U9183 (N_9183,N_8772,N_8800);
xnor U9184 (N_9184,N_8801,N_8848);
nor U9185 (N_9185,N_8862,N_8876);
nor U9186 (N_9186,N_8899,N_8839);
or U9187 (N_9187,N_8829,N_8834);
nand U9188 (N_9188,N_8792,N_8910);
or U9189 (N_9189,N_8848,N_8865);
and U9190 (N_9190,N_8984,N_8752);
xor U9191 (N_9191,N_8929,N_8859);
nand U9192 (N_9192,N_8954,N_8901);
nand U9193 (N_9193,N_8844,N_8834);
and U9194 (N_9194,N_8812,N_8872);
or U9195 (N_9195,N_8969,N_8961);
and U9196 (N_9196,N_8962,N_8956);
xor U9197 (N_9197,N_8996,N_8883);
nand U9198 (N_9198,N_8840,N_8832);
nor U9199 (N_9199,N_8765,N_8817);
or U9200 (N_9200,N_8956,N_8845);
and U9201 (N_9201,N_8839,N_8961);
and U9202 (N_9202,N_8984,N_8779);
nand U9203 (N_9203,N_8828,N_8862);
nor U9204 (N_9204,N_8950,N_8889);
or U9205 (N_9205,N_8907,N_8758);
nor U9206 (N_9206,N_8859,N_8801);
and U9207 (N_9207,N_8782,N_8891);
or U9208 (N_9208,N_8795,N_8941);
or U9209 (N_9209,N_8936,N_8885);
xor U9210 (N_9210,N_8803,N_8970);
or U9211 (N_9211,N_8881,N_8855);
and U9212 (N_9212,N_8991,N_8862);
or U9213 (N_9213,N_8880,N_8788);
xor U9214 (N_9214,N_8953,N_8785);
or U9215 (N_9215,N_8850,N_8973);
nand U9216 (N_9216,N_8795,N_8991);
and U9217 (N_9217,N_8890,N_8996);
or U9218 (N_9218,N_8996,N_8843);
nor U9219 (N_9219,N_8859,N_8992);
and U9220 (N_9220,N_8961,N_8783);
xor U9221 (N_9221,N_8779,N_8822);
xnor U9222 (N_9222,N_8959,N_8788);
or U9223 (N_9223,N_8912,N_8791);
xnor U9224 (N_9224,N_8910,N_8956);
nand U9225 (N_9225,N_8956,N_8833);
nand U9226 (N_9226,N_8913,N_8989);
or U9227 (N_9227,N_8923,N_8997);
or U9228 (N_9228,N_8786,N_8896);
and U9229 (N_9229,N_8856,N_8919);
and U9230 (N_9230,N_8924,N_8921);
nor U9231 (N_9231,N_8928,N_8954);
nand U9232 (N_9232,N_8761,N_8809);
nor U9233 (N_9233,N_8787,N_8897);
and U9234 (N_9234,N_8925,N_8980);
nor U9235 (N_9235,N_8946,N_8964);
nand U9236 (N_9236,N_8909,N_8758);
and U9237 (N_9237,N_8876,N_8836);
nand U9238 (N_9238,N_8957,N_8905);
and U9239 (N_9239,N_8785,N_8891);
nand U9240 (N_9240,N_8863,N_8871);
and U9241 (N_9241,N_8902,N_8954);
nor U9242 (N_9242,N_8855,N_8959);
nor U9243 (N_9243,N_8886,N_8921);
nor U9244 (N_9244,N_8782,N_8933);
or U9245 (N_9245,N_8996,N_8887);
nand U9246 (N_9246,N_8830,N_8939);
nand U9247 (N_9247,N_8786,N_8768);
or U9248 (N_9248,N_8936,N_8984);
or U9249 (N_9249,N_8940,N_8769);
nor U9250 (N_9250,N_9173,N_9023);
nor U9251 (N_9251,N_9075,N_9131);
and U9252 (N_9252,N_9241,N_9222);
nor U9253 (N_9253,N_9074,N_9120);
and U9254 (N_9254,N_9190,N_9051);
nand U9255 (N_9255,N_9133,N_9101);
or U9256 (N_9256,N_9172,N_9117);
or U9257 (N_9257,N_9056,N_9020);
or U9258 (N_9258,N_9239,N_9076);
and U9259 (N_9259,N_9149,N_9165);
and U9260 (N_9260,N_9046,N_9061);
nor U9261 (N_9261,N_9093,N_9016);
or U9262 (N_9262,N_9179,N_9195);
or U9263 (N_9263,N_9155,N_9066);
nand U9264 (N_9264,N_9216,N_9132);
nor U9265 (N_9265,N_9105,N_9090);
and U9266 (N_9266,N_9049,N_9236);
nor U9267 (N_9267,N_9048,N_9007);
nor U9268 (N_9268,N_9013,N_9204);
nor U9269 (N_9269,N_9189,N_9191);
nand U9270 (N_9270,N_9002,N_9147);
and U9271 (N_9271,N_9010,N_9006);
and U9272 (N_9272,N_9121,N_9040);
nor U9273 (N_9273,N_9087,N_9035);
nand U9274 (N_9274,N_9161,N_9055);
nor U9275 (N_9275,N_9152,N_9018);
nand U9276 (N_9276,N_9178,N_9208);
nor U9277 (N_9277,N_9118,N_9140);
nand U9278 (N_9278,N_9205,N_9188);
or U9279 (N_9279,N_9242,N_9041);
nor U9280 (N_9280,N_9124,N_9108);
or U9281 (N_9281,N_9114,N_9111);
nand U9282 (N_9282,N_9158,N_9171);
nand U9283 (N_9283,N_9135,N_9017);
nor U9284 (N_9284,N_9065,N_9160);
nand U9285 (N_9285,N_9156,N_9110);
nand U9286 (N_9286,N_9166,N_9092);
and U9287 (N_9287,N_9116,N_9215);
nand U9288 (N_9288,N_9005,N_9247);
and U9289 (N_9289,N_9115,N_9176);
nor U9290 (N_9290,N_9070,N_9200);
nor U9291 (N_9291,N_9138,N_9083);
nand U9292 (N_9292,N_9032,N_9159);
or U9293 (N_9293,N_9003,N_9184);
xor U9294 (N_9294,N_9021,N_9063);
nand U9295 (N_9295,N_9091,N_9211);
xnor U9296 (N_9296,N_9054,N_9145);
or U9297 (N_9297,N_9246,N_9226);
nand U9298 (N_9298,N_9099,N_9085);
or U9299 (N_9299,N_9137,N_9029);
and U9300 (N_9300,N_9014,N_9037);
nand U9301 (N_9301,N_9059,N_9001);
nand U9302 (N_9302,N_9198,N_9106);
xnor U9303 (N_9303,N_9045,N_9095);
nor U9304 (N_9304,N_9047,N_9139);
and U9305 (N_9305,N_9201,N_9043);
nand U9306 (N_9306,N_9019,N_9126);
or U9307 (N_9307,N_9183,N_9067);
xnor U9308 (N_9308,N_9207,N_9213);
nand U9309 (N_9309,N_9233,N_9234);
nor U9310 (N_9310,N_9096,N_9097);
or U9311 (N_9311,N_9125,N_9206);
nand U9312 (N_9312,N_9080,N_9248);
and U9313 (N_9313,N_9202,N_9244);
and U9314 (N_9314,N_9119,N_9130);
nand U9315 (N_9315,N_9199,N_9079);
nor U9316 (N_9316,N_9238,N_9036);
nand U9317 (N_9317,N_9000,N_9192);
or U9318 (N_9318,N_9237,N_9069);
nor U9319 (N_9319,N_9086,N_9068);
xnor U9320 (N_9320,N_9098,N_9012);
nor U9321 (N_9321,N_9058,N_9136);
or U9322 (N_9322,N_9185,N_9122);
or U9323 (N_9323,N_9245,N_9225);
nand U9324 (N_9324,N_9243,N_9217);
or U9325 (N_9325,N_9218,N_9170);
nand U9326 (N_9326,N_9009,N_9194);
nand U9327 (N_9327,N_9052,N_9077);
nor U9328 (N_9328,N_9011,N_9025);
and U9329 (N_9329,N_9187,N_9231);
and U9330 (N_9330,N_9064,N_9157);
xnor U9331 (N_9331,N_9078,N_9109);
and U9332 (N_9332,N_9232,N_9146);
or U9333 (N_9333,N_9031,N_9151);
nor U9334 (N_9334,N_9028,N_9154);
xor U9335 (N_9335,N_9150,N_9210);
and U9336 (N_9336,N_9103,N_9107);
or U9337 (N_9337,N_9113,N_9081);
or U9338 (N_9338,N_9039,N_9220);
or U9339 (N_9339,N_9134,N_9062);
nand U9340 (N_9340,N_9094,N_9181);
or U9341 (N_9341,N_9162,N_9203);
or U9342 (N_9342,N_9084,N_9167);
or U9343 (N_9343,N_9044,N_9240);
nor U9344 (N_9344,N_9144,N_9142);
xnor U9345 (N_9345,N_9228,N_9030);
xnor U9346 (N_9346,N_9008,N_9141);
nand U9347 (N_9347,N_9024,N_9219);
and U9348 (N_9348,N_9175,N_9112);
nand U9349 (N_9349,N_9128,N_9027);
nand U9350 (N_9350,N_9197,N_9163);
nand U9351 (N_9351,N_9224,N_9129);
nor U9352 (N_9352,N_9057,N_9033);
nand U9353 (N_9353,N_9169,N_9223);
or U9354 (N_9354,N_9235,N_9182);
or U9355 (N_9355,N_9015,N_9148);
or U9356 (N_9356,N_9153,N_9229);
and U9357 (N_9357,N_9221,N_9082);
or U9358 (N_9358,N_9212,N_9089);
or U9359 (N_9359,N_9073,N_9214);
or U9360 (N_9360,N_9227,N_9193);
xnor U9361 (N_9361,N_9072,N_9168);
or U9362 (N_9362,N_9004,N_9104);
and U9363 (N_9363,N_9164,N_9196);
nand U9364 (N_9364,N_9230,N_9177);
or U9365 (N_9365,N_9249,N_9050);
or U9366 (N_9366,N_9071,N_9100);
nor U9367 (N_9367,N_9127,N_9180);
nand U9368 (N_9368,N_9174,N_9042);
nand U9369 (N_9369,N_9123,N_9209);
and U9370 (N_9370,N_9186,N_9038);
xor U9371 (N_9371,N_9034,N_9022);
and U9372 (N_9372,N_9088,N_9053);
and U9373 (N_9373,N_9102,N_9060);
nand U9374 (N_9374,N_9026,N_9143);
and U9375 (N_9375,N_9205,N_9169);
xor U9376 (N_9376,N_9050,N_9213);
xnor U9377 (N_9377,N_9041,N_9141);
nand U9378 (N_9378,N_9059,N_9176);
nand U9379 (N_9379,N_9050,N_9112);
and U9380 (N_9380,N_9221,N_9092);
and U9381 (N_9381,N_9042,N_9163);
or U9382 (N_9382,N_9227,N_9017);
nor U9383 (N_9383,N_9052,N_9078);
and U9384 (N_9384,N_9043,N_9204);
or U9385 (N_9385,N_9101,N_9031);
and U9386 (N_9386,N_9218,N_9040);
xor U9387 (N_9387,N_9055,N_9198);
nor U9388 (N_9388,N_9146,N_9054);
nor U9389 (N_9389,N_9238,N_9248);
or U9390 (N_9390,N_9239,N_9181);
nor U9391 (N_9391,N_9199,N_9236);
nand U9392 (N_9392,N_9003,N_9048);
or U9393 (N_9393,N_9044,N_9129);
xor U9394 (N_9394,N_9079,N_9167);
nor U9395 (N_9395,N_9188,N_9051);
and U9396 (N_9396,N_9248,N_9212);
or U9397 (N_9397,N_9216,N_9042);
and U9398 (N_9398,N_9080,N_9115);
nand U9399 (N_9399,N_9110,N_9167);
or U9400 (N_9400,N_9131,N_9182);
and U9401 (N_9401,N_9103,N_9206);
nand U9402 (N_9402,N_9085,N_9176);
xnor U9403 (N_9403,N_9082,N_9028);
or U9404 (N_9404,N_9004,N_9053);
or U9405 (N_9405,N_9078,N_9139);
nand U9406 (N_9406,N_9115,N_9054);
nor U9407 (N_9407,N_9053,N_9058);
nand U9408 (N_9408,N_9121,N_9239);
nand U9409 (N_9409,N_9002,N_9112);
nand U9410 (N_9410,N_9098,N_9172);
and U9411 (N_9411,N_9038,N_9025);
or U9412 (N_9412,N_9213,N_9125);
nor U9413 (N_9413,N_9129,N_9176);
or U9414 (N_9414,N_9132,N_9102);
and U9415 (N_9415,N_9124,N_9113);
nor U9416 (N_9416,N_9240,N_9201);
nor U9417 (N_9417,N_9040,N_9203);
and U9418 (N_9418,N_9144,N_9187);
nand U9419 (N_9419,N_9072,N_9038);
or U9420 (N_9420,N_9201,N_9133);
or U9421 (N_9421,N_9012,N_9061);
and U9422 (N_9422,N_9095,N_9148);
and U9423 (N_9423,N_9230,N_9006);
or U9424 (N_9424,N_9187,N_9043);
and U9425 (N_9425,N_9162,N_9215);
nor U9426 (N_9426,N_9197,N_9206);
nand U9427 (N_9427,N_9068,N_9247);
and U9428 (N_9428,N_9073,N_9151);
nor U9429 (N_9429,N_9103,N_9053);
and U9430 (N_9430,N_9192,N_9209);
nand U9431 (N_9431,N_9022,N_9180);
and U9432 (N_9432,N_9190,N_9123);
nand U9433 (N_9433,N_9206,N_9166);
and U9434 (N_9434,N_9156,N_9038);
nor U9435 (N_9435,N_9061,N_9151);
or U9436 (N_9436,N_9095,N_9143);
nor U9437 (N_9437,N_9140,N_9207);
nor U9438 (N_9438,N_9228,N_9049);
and U9439 (N_9439,N_9080,N_9098);
nor U9440 (N_9440,N_9000,N_9151);
and U9441 (N_9441,N_9048,N_9112);
and U9442 (N_9442,N_9186,N_9011);
and U9443 (N_9443,N_9020,N_9209);
nand U9444 (N_9444,N_9219,N_9062);
or U9445 (N_9445,N_9206,N_9235);
nand U9446 (N_9446,N_9231,N_9137);
and U9447 (N_9447,N_9038,N_9228);
and U9448 (N_9448,N_9228,N_9073);
xor U9449 (N_9449,N_9235,N_9215);
and U9450 (N_9450,N_9099,N_9186);
nor U9451 (N_9451,N_9107,N_9165);
or U9452 (N_9452,N_9229,N_9101);
and U9453 (N_9453,N_9015,N_9177);
or U9454 (N_9454,N_9174,N_9198);
nor U9455 (N_9455,N_9116,N_9144);
and U9456 (N_9456,N_9018,N_9045);
nand U9457 (N_9457,N_9096,N_9170);
xor U9458 (N_9458,N_9065,N_9018);
xor U9459 (N_9459,N_9063,N_9222);
nor U9460 (N_9460,N_9030,N_9147);
nor U9461 (N_9461,N_9190,N_9137);
or U9462 (N_9462,N_9069,N_9169);
xor U9463 (N_9463,N_9198,N_9150);
nand U9464 (N_9464,N_9200,N_9164);
nand U9465 (N_9465,N_9091,N_9083);
and U9466 (N_9466,N_9181,N_9089);
and U9467 (N_9467,N_9117,N_9173);
or U9468 (N_9468,N_9212,N_9125);
nand U9469 (N_9469,N_9170,N_9145);
xor U9470 (N_9470,N_9013,N_9058);
or U9471 (N_9471,N_9123,N_9009);
nand U9472 (N_9472,N_9186,N_9059);
nor U9473 (N_9473,N_9065,N_9100);
and U9474 (N_9474,N_9074,N_9181);
nand U9475 (N_9475,N_9089,N_9036);
nor U9476 (N_9476,N_9009,N_9016);
xor U9477 (N_9477,N_9184,N_9170);
nor U9478 (N_9478,N_9231,N_9052);
and U9479 (N_9479,N_9063,N_9000);
nand U9480 (N_9480,N_9249,N_9139);
and U9481 (N_9481,N_9096,N_9108);
and U9482 (N_9482,N_9152,N_9074);
or U9483 (N_9483,N_9190,N_9114);
nor U9484 (N_9484,N_9108,N_9112);
and U9485 (N_9485,N_9171,N_9128);
or U9486 (N_9486,N_9188,N_9184);
or U9487 (N_9487,N_9058,N_9009);
and U9488 (N_9488,N_9039,N_9112);
and U9489 (N_9489,N_9091,N_9173);
nor U9490 (N_9490,N_9108,N_9072);
nand U9491 (N_9491,N_9052,N_9164);
nand U9492 (N_9492,N_9039,N_9237);
and U9493 (N_9493,N_9022,N_9091);
and U9494 (N_9494,N_9094,N_9243);
or U9495 (N_9495,N_9135,N_9169);
or U9496 (N_9496,N_9160,N_9067);
xnor U9497 (N_9497,N_9221,N_9109);
and U9498 (N_9498,N_9234,N_9207);
nor U9499 (N_9499,N_9248,N_9146);
and U9500 (N_9500,N_9407,N_9448);
xor U9501 (N_9501,N_9253,N_9330);
xnor U9502 (N_9502,N_9318,N_9365);
nor U9503 (N_9503,N_9285,N_9466);
or U9504 (N_9504,N_9492,N_9334);
nor U9505 (N_9505,N_9412,N_9396);
nand U9506 (N_9506,N_9320,N_9474);
or U9507 (N_9507,N_9265,N_9374);
xnor U9508 (N_9508,N_9279,N_9468);
nor U9509 (N_9509,N_9389,N_9333);
or U9510 (N_9510,N_9347,N_9331);
nor U9511 (N_9511,N_9312,N_9354);
nor U9512 (N_9512,N_9344,N_9256);
and U9513 (N_9513,N_9300,N_9410);
nand U9514 (N_9514,N_9342,N_9337);
and U9515 (N_9515,N_9499,N_9328);
and U9516 (N_9516,N_9455,N_9440);
nor U9517 (N_9517,N_9377,N_9379);
nor U9518 (N_9518,N_9489,N_9481);
and U9519 (N_9519,N_9280,N_9409);
nand U9520 (N_9520,N_9414,N_9338);
and U9521 (N_9521,N_9370,N_9319);
or U9522 (N_9522,N_9433,N_9257);
and U9523 (N_9523,N_9498,N_9335);
or U9524 (N_9524,N_9266,N_9294);
or U9525 (N_9525,N_9443,N_9281);
and U9526 (N_9526,N_9416,N_9491);
and U9527 (N_9527,N_9306,N_9252);
or U9528 (N_9528,N_9329,N_9479);
and U9529 (N_9529,N_9355,N_9322);
xnor U9530 (N_9530,N_9385,N_9388);
nand U9531 (N_9531,N_9386,N_9434);
and U9532 (N_9532,N_9324,N_9418);
xnor U9533 (N_9533,N_9399,N_9454);
nor U9534 (N_9534,N_9462,N_9356);
and U9535 (N_9535,N_9393,N_9382);
and U9536 (N_9536,N_9442,N_9264);
or U9537 (N_9537,N_9371,N_9341);
nand U9538 (N_9538,N_9268,N_9406);
nor U9539 (N_9539,N_9295,N_9470);
xnor U9540 (N_9540,N_9284,N_9384);
nor U9541 (N_9541,N_9304,N_9287);
and U9542 (N_9542,N_9436,N_9378);
nor U9543 (N_9543,N_9428,N_9313);
nor U9544 (N_9544,N_9293,N_9340);
nand U9545 (N_9545,N_9387,N_9361);
nor U9546 (N_9546,N_9269,N_9299);
and U9547 (N_9547,N_9472,N_9453);
and U9548 (N_9548,N_9450,N_9263);
xor U9549 (N_9549,N_9480,N_9345);
nand U9550 (N_9550,N_9458,N_9497);
xnor U9551 (N_9551,N_9292,N_9441);
and U9552 (N_9552,N_9309,N_9346);
or U9553 (N_9553,N_9426,N_9251);
nor U9554 (N_9554,N_9302,N_9425);
nor U9555 (N_9555,N_9296,N_9459);
nand U9556 (N_9556,N_9259,N_9272);
nor U9557 (N_9557,N_9368,N_9317);
nor U9558 (N_9558,N_9392,N_9349);
or U9559 (N_9559,N_9339,N_9314);
or U9560 (N_9560,N_9326,N_9430);
nor U9561 (N_9561,N_9276,N_9278);
nand U9562 (N_9562,N_9478,N_9417);
or U9563 (N_9563,N_9283,N_9362);
nor U9564 (N_9564,N_9363,N_9273);
or U9565 (N_9565,N_9488,N_9424);
nor U9566 (N_9566,N_9250,N_9432);
or U9567 (N_9567,N_9282,N_9277);
xnor U9568 (N_9568,N_9305,N_9381);
or U9569 (N_9569,N_9469,N_9311);
or U9570 (N_9570,N_9380,N_9485);
nor U9571 (N_9571,N_9288,N_9486);
or U9572 (N_9572,N_9400,N_9332);
or U9573 (N_9573,N_9286,N_9401);
and U9574 (N_9574,N_9353,N_9415);
nand U9575 (N_9575,N_9348,N_9402);
nand U9576 (N_9576,N_9270,N_9445);
nand U9577 (N_9577,N_9427,N_9411);
nand U9578 (N_9578,N_9383,N_9366);
nand U9579 (N_9579,N_9420,N_9460);
nor U9580 (N_9580,N_9289,N_9303);
or U9581 (N_9581,N_9301,N_9315);
and U9582 (N_9582,N_9423,N_9465);
xor U9583 (N_9583,N_9260,N_9463);
nor U9584 (N_9584,N_9372,N_9464);
and U9585 (N_9585,N_9290,N_9394);
nor U9586 (N_9586,N_9487,N_9467);
or U9587 (N_9587,N_9369,N_9473);
nor U9588 (N_9588,N_9360,N_9475);
and U9589 (N_9589,N_9404,N_9439);
or U9590 (N_9590,N_9456,N_9391);
and U9591 (N_9591,N_9395,N_9350);
nand U9592 (N_9592,N_9352,N_9477);
or U9593 (N_9593,N_9490,N_9496);
nor U9594 (N_9594,N_9343,N_9449);
and U9595 (N_9595,N_9494,N_9398);
and U9596 (N_9596,N_9451,N_9403);
nor U9597 (N_9597,N_9262,N_9321);
or U9598 (N_9598,N_9359,N_9307);
nand U9599 (N_9599,N_9316,N_9327);
nand U9600 (N_9600,N_9375,N_9255);
or U9601 (N_9601,N_9471,N_9438);
or U9602 (N_9602,N_9483,N_9431);
nor U9603 (N_9603,N_9297,N_9493);
nand U9604 (N_9604,N_9336,N_9267);
or U9605 (N_9605,N_9429,N_9325);
xnor U9606 (N_9606,N_9408,N_9275);
nor U9607 (N_9607,N_9373,N_9364);
or U9608 (N_9608,N_9444,N_9419);
nand U9609 (N_9609,N_9435,N_9367);
or U9610 (N_9610,N_9495,N_9291);
nor U9611 (N_9611,N_9261,N_9421);
or U9612 (N_9612,N_9397,N_9447);
and U9613 (N_9613,N_9357,N_9413);
nand U9614 (N_9614,N_9254,N_9258);
or U9615 (N_9615,N_9274,N_9351);
and U9616 (N_9616,N_9323,N_9358);
xor U9617 (N_9617,N_9308,N_9376);
nand U9618 (N_9618,N_9446,N_9457);
and U9619 (N_9619,N_9482,N_9298);
and U9620 (N_9620,N_9452,N_9390);
nor U9621 (N_9621,N_9461,N_9422);
and U9622 (N_9622,N_9476,N_9271);
or U9623 (N_9623,N_9437,N_9405);
xnor U9624 (N_9624,N_9310,N_9484);
xor U9625 (N_9625,N_9422,N_9273);
nor U9626 (N_9626,N_9420,N_9317);
and U9627 (N_9627,N_9323,N_9377);
xor U9628 (N_9628,N_9270,N_9454);
nand U9629 (N_9629,N_9395,N_9341);
nor U9630 (N_9630,N_9282,N_9285);
and U9631 (N_9631,N_9326,N_9401);
or U9632 (N_9632,N_9462,N_9363);
or U9633 (N_9633,N_9432,N_9459);
and U9634 (N_9634,N_9359,N_9352);
nand U9635 (N_9635,N_9369,N_9323);
or U9636 (N_9636,N_9465,N_9343);
nor U9637 (N_9637,N_9480,N_9273);
nand U9638 (N_9638,N_9403,N_9472);
nand U9639 (N_9639,N_9327,N_9417);
or U9640 (N_9640,N_9356,N_9405);
nor U9641 (N_9641,N_9428,N_9305);
xnor U9642 (N_9642,N_9324,N_9441);
nor U9643 (N_9643,N_9308,N_9331);
nand U9644 (N_9644,N_9277,N_9256);
nor U9645 (N_9645,N_9294,N_9274);
or U9646 (N_9646,N_9336,N_9289);
xnor U9647 (N_9647,N_9409,N_9345);
nor U9648 (N_9648,N_9277,N_9369);
and U9649 (N_9649,N_9375,N_9299);
and U9650 (N_9650,N_9354,N_9497);
nand U9651 (N_9651,N_9429,N_9301);
or U9652 (N_9652,N_9288,N_9468);
nor U9653 (N_9653,N_9305,N_9304);
and U9654 (N_9654,N_9352,N_9442);
nand U9655 (N_9655,N_9473,N_9378);
or U9656 (N_9656,N_9308,N_9272);
or U9657 (N_9657,N_9455,N_9253);
nand U9658 (N_9658,N_9331,N_9480);
or U9659 (N_9659,N_9384,N_9370);
nor U9660 (N_9660,N_9280,N_9392);
or U9661 (N_9661,N_9474,N_9457);
and U9662 (N_9662,N_9309,N_9296);
nand U9663 (N_9663,N_9399,N_9403);
or U9664 (N_9664,N_9417,N_9402);
nand U9665 (N_9665,N_9306,N_9348);
xor U9666 (N_9666,N_9322,N_9477);
nand U9667 (N_9667,N_9350,N_9307);
and U9668 (N_9668,N_9443,N_9464);
or U9669 (N_9669,N_9374,N_9414);
nand U9670 (N_9670,N_9299,N_9288);
nor U9671 (N_9671,N_9341,N_9264);
nand U9672 (N_9672,N_9407,N_9486);
and U9673 (N_9673,N_9324,N_9490);
or U9674 (N_9674,N_9417,N_9464);
xor U9675 (N_9675,N_9303,N_9284);
nand U9676 (N_9676,N_9393,N_9284);
nand U9677 (N_9677,N_9492,N_9392);
and U9678 (N_9678,N_9440,N_9447);
nor U9679 (N_9679,N_9369,N_9471);
and U9680 (N_9680,N_9368,N_9324);
or U9681 (N_9681,N_9382,N_9304);
nor U9682 (N_9682,N_9428,N_9336);
nand U9683 (N_9683,N_9445,N_9279);
or U9684 (N_9684,N_9384,N_9448);
or U9685 (N_9685,N_9261,N_9372);
xor U9686 (N_9686,N_9475,N_9285);
nand U9687 (N_9687,N_9425,N_9295);
xnor U9688 (N_9688,N_9277,N_9495);
nor U9689 (N_9689,N_9410,N_9376);
nor U9690 (N_9690,N_9493,N_9314);
nand U9691 (N_9691,N_9423,N_9420);
or U9692 (N_9692,N_9381,N_9366);
or U9693 (N_9693,N_9358,N_9446);
nand U9694 (N_9694,N_9498,N_9436);
nor U9695 (N_9695,N_9354,N_9437);
and U9696 (N_9696,N_9261,N_9279);
and U9697 (N_9697,N_9287,N_9339);
and U9698 (N_9698,N_9354,N_9402);
or U9699 (N_9699,N_9355,N_9314);
or U9700 (N_9700,N_9390,N_9297);
nor U9701 (N_9701,N_9404,N_9438);
nand U9702 (N_9702,N_9396,N_9384);
nor U9703 (N_9703,N_9479,N_9269);
nand U9704 (N_9704,N_9399,N_9336);
nor U9705 (N_9705,N_9348,N_9269);
or U9706 (N_9706,N_9292,N_9271);
nor U9707 (N_9707,N_9297,N_9320);
and U9708 (N_9708,N_9486,N_9255);
nand U9709 (N_9709,N_9445,N_9432);
nor U9710 (N_9710,N_9323,N_9492);
nand U9711 (N_9711,N_9465,N_9376);
or U9712 (N_9712,N_9340,N_9263);
and U9713 (N_9713,N_9331,N_9300);
and U9714 (N_9714,N_9381,N_9484);
and U9715 (N_9715,N_9315,N_9485);
nand U9716 (N_9716,N_9326,N_9253);
nand U9717 (N_9717,N_9288,N_9284);
and U9718 (N_9718,N_9291,N_9313);
xor U9719 (N_9719,N_9417,N_9485);
xor U9720 (N_9720,N_9314,N_9470);
and U9721 (N_9721,N_9350,N_9372);
xor U9722 (N_9722,N_9298,N_9478);
nand U9723 (N_9723,N_9325,N_9423);
nand U9724 (N_9724,N_9498,N_9403);
nor U9725 (N_9725,N_9467,N_9438);
nand U9726 (N_9726,N_9287,N_9350);
and U9727 (N_9727,N_9458,N_9377);
and U9728 (N_9728,N_9252,N_9315);
and U9729 (N_9729,N_9446,N_9387);
nand U9730 (N_9730,N_9289,N_9319);
or U9731 (N_9731,N_9391,N_9274);
or U9732 (N_9732,N_9372,N_9263);
and U9733 (N_9733,N_9349,N_9391);
nor U9734 (N_9734,N_9408,N_9350);
and U9735 (N_9735,N_9342,N_9350);
and U9736 (N_9736,N_9434,N_9362);
or U9737 (N_9737,N_9480,N_9429);
nor U9738 (N_9738,N_9434,N_9361);
and U9739 (N_9739,N_9258,N_9345);
nand U9740 (N_9740,N_9279,N_9309);
nor U9741 (N_9741,N_9341,N_9271);
nor U9742 (N_9742,N_9330,N_9440);
xor U9743 (N_9743,N_9448,N_9330);
or U9744 (N_9744,N_9417,N_9254);
nand U9745 (N_9745,N_9331,N_9418);
or U9746 (N_9746,N_9499,N_9324);
and U9747 (N_9747,N_9252,N_9389);
nor U9748 (N_9748,N_9431,N_9420);
nand U9749 (N_9749,N_9484,N_9356);
nor U9750 (N_9750,N_9532,N_9625);
nor U9751 (N_9751,N_9703,N_9747);
or U9752 (N_9752,N_9666,N_9620);
and U9753 (N_9753,N_9590,N_9578);
nor U9754 (N_9754,N_9698,N_9573);
xor U9755 (N_9755,N_9543,N_9581);
and U9756 (N_9756,N_9694,N_9742);
nor U9757 (N_9757,N_9651,N_9525);
nor U9758 (N_9758,N_9601,N_9583);
or U9759 (N_9759,N_9561,N_9732);
nor U9760 (N_9760,N_9604,N_9683);
nor U9761 (N_9761,N_9609,N_9591);
and U9762 (N_9762,N_9551,N_9664);
nor U9763 (N_9763,N_9663,N_9520);
and U9764 (N_9764,N_9595,N_9706);
or U9765 (N_9765,N_9546,N_9647);
and U9766 (N_9766,N_9711,N_9531);
or U9767 (N_9767,N_9717,N_9735);
and U9768 (N_9768,N_9524,N_9748);
nand U9769 (N_9769,N_9512,N_9724);
or U9770 (N_9770,N_9745,N_9648);
nand U9771 (N_9771,N_9576,N_9707);
and U9772 (N_9772,N_9712,N_9656);
nand U9773 (N_9773,N_9582,N_9746);
xor U9774 (N_9774,N_9642,N_9741);
xor U9775 (N_9775,N_9572,N_9644);
or U9776 (N_9776,N_9661,N_9552);
nand U9777 (N_9777,N_9692,N_9618);
or U9778 (N_9778,N_9569,N_9677);
or U9779 (N_9779,N_9702,N_9550);
nor U9780 (N_9780,N_9743,N_9521);
and U9781 (N_9781,N_9701,N_9669);
or U9782 (N_9782,N_9719,N_9507);
or U9783 (N_9783,N_9690,N_9697);
and U9784 (N_9784,N_9622,N_9641);
and U9785 (N_9785,N_9553,N_9508);
nand U9786 (N_9786,N_9584,N_9602);
nand U9787 (N_9787,N_9660,N_9639);
or U9788 (N_9788,N_9659,N_9614);
and U9789 (N_9789,N_9675,N_9646);
and U9790 (N_9790,N_9668,N_9594);
or U9791 (N_9791,N_9509,N_9565);
nand U9792 (N_9792,N_9617,N_9638);
and U9793 (N_9793,N_9580,N_9676);
nor U9794 (N_9794,N_9517,N_9678);
and U9795 (N_9795,N_9559,N_9686);
and U9796 (N_9796,N_9672,N_9731);
or U9797 (N_9797,N_9548,N_9700);
nand U9798 (N_9798,N_9739,N_9516);
nor U9799 (N_9799,N_9563,N_9611);
or U9800 (N_9800,N_9527,N_9518);
nor U9801 (N_9801,N_9721,N_9574);
and U9802 (N_9802,N_9522,N_9515);
and U9803 (N_9803,N_9635,N_9506);
nand U9804 (N_9804,N_9654,N_9722);
and U9805 (N_9805,N_9681,N_9534);
nor U9806 (N_9806,N_9730,N_9530);
nor U9807 (N_9807,N_9556,N_9529);
and U9808 (N_9808,N_9504,N_9579);
nor U9809 (N_9809,N_9519,N_9673);
or U9810 (N_9810,N_9560,N_9636);
or U9811 (N_9811,N_9631,N_9523);
or U9812 (N_9812,N_9744,N_9691);
nor U9813 (N_9813,N_9586,N_9645);
and U9814 (N_9814,N_9526,N_9542);
or U9815 (N_9815,N_9615,N_9650);
or U9816 (N_9816,N_9699,N_9723);
or U9817 (N_9817,N_9679,N_9536);
nand U9818 (N_9818,N_9557,N_9740);
and U9819 (N_9819,N_9575,N_9599);
nor U9820 (N_9820,N_9674,N_9670);
nand U9821 (N_9821,N_9728,N_9640);
or U9822 (N_9822,N_9685,N_9667);
and U9823 (N_9823,N_9680,N_9535);
and U9824 (N_9824,N_9671,N_9605);
nor U9825 (N_9825,N_9716,N_9577);
nand U9826 (N_9826,N_9738,N_9657);
nand U9827 (N_9827,N_9510,N_9637);
xor U9828 (N_9828,N_9749,N_9727);
or U9829 (N_9829,N_9705,N_9547);
xor U9830 (N_9830,N_9539,N_9693);
and U9831 (N_9831,N_9607,N_9585);
nor U9832 (N_9832,N_9684,N_9729);
nand U9833 (N_9833,N_9649,N_9558);
or U9834 (N_9834,N_9567,N_9513);
xnor U9835 (N_9835,N_9630,N_9709);
nor U9836 (N_9836,N_9733,N_9528);
or U9837 (N_9837,N_9533,N_9715);
or U9838 (N_9838,N_9514,N_9545);
nor U9839 (N_9839,N_9624,N_9562);
or U9840 (N_9840,N_9734,N_9665);
or U9841 (N_9841,N_9689,N_9708);
or U9842 (N_9842,N_9598,N_9633);
or U9843 (N_9843,N_9658,N_9629);
nand U9844 (N_9844,N_9714,N_9710);
xnor U9845 (N_9845,N_9596,N_9549);
or U9846 (N_9846,N_9544,N_9589);
nand U9847 (N_9847,N_9720,N_9632);
xnor U9848 (N_9848,N_9626,N_9718);
and U9849 (N_9849,N_9503,N_9613);
nand U9850 (N_9850,N_9587,N_9662);
nand U9851 (N_9851,N_9566,N_9695);
nand U9852 (N_9852,N_9592,N_9696);
and U9853 (N_9853,N_9726,N_9682);
nor U9854 (N_9854,N_9610,N_9501);
or U9855 (N_9855,N_9612,N_9652);
or U9856 (N_9856,N_9511,N_9541);
nor U9857 (N_9857,N_9568,N_9634);
or U9858 (N_9858,N_9627,N_9623);
and U9859 (N_9859,N_9608,N_9606);
and U9860 (N_9860,N_9643,N_9619);
nand U9861 (N_9861,N_9621,N_9603);
and U9862 (N_9862,N_9737,N_9616);
nand U9863 (N_9863,N_9540,N_9688);
nor U9864 (N_9864,N_9687,N_9597);
nor U9865 (N_9865,N_9505,N_9537);
nand U9866 (N_9866,N_9554,N_9564);
and U9867 (N_9867,N_9538,N_9593);
and U9868 (N_9868,N_9725,N_9570);
nand U9869 (N_9869,N_9628,N_9588);
nor U9870 (N_9870,N_9655,N_9736);
and U9871 (N_9871,N_9502,N_9704);
or U9872 (N_9872,N_9600,N_9713);
and U9873 (N_9873,N_9500,N_9571);
and U9874 (N_9874,N_9653,N_9555);
nand U9875 (N_9875,N_9559,N_9690);
and U9876 (N_9876,N_9667,N_9674);
or U9877 (N_9877,N_9514,N_9707);
and U9878 (N_9878,N_9549,N_9590);
or U9879 (N_9879,N_9516,N_9505);
and U9880 (N_9880,N_9552,N_9666);
nand U9881 (N_9881,N_9531,N_9588);
nand U9882 (N_9882,N_9604,N_9641);
or U9883 (N_9883,N_9632,N_9713);
nor U9884 (N_9884,N_9689,N_9512);
nor U9885 (N_9885,N_9706,N_9742);
nand U9886 (N_9886,N_9685,N_9635);
nand U9887 (N_9887,N_9662,N_9517);
or U9888 (N_9888,N_9665,N_9736);
nor U9889 (N_9889,N_9607,N_9503);
xor U9890 (N_9890,N_9749,N_9613);
or U9891 (N_9891,N_9522,N_9613);
and U9892 (N_9892,N_9518,N_9736);
or U9893 (N_9893,N_9731,N_9691);
nor U9894 (N_9894,N_9618,N_9720);
nand U9895 (N_9895,N_9621,N_9588);
and U9896 (N_9896,N_9643,N_9602);
and U9897 (N_9897,N_9631,N_9543);
nand U9898 (N_9898,N_9597,N_9662);
and U9899 (N_9899,N_9601,N_9509);
nand U9900 (N_9900,N_9522,N_9670);
xor U9901 (N_9901,N_9533,N_9614);
and U9902 (N_9902,N_9500,N_9722);
nand U9903 (N_9903,N_9732,N_9571);
and U9904 (N_9904,N_9705,N_9595);
nand U9905 (N_9905,N_9672,N_9620);
and U9906 (N_9906,N_9572,N_9726);
and U9907 (N_9907,N_9645,N_9729);
or U9908 (N_9908,N_9585,N_9519);
nand U9909 (N_9909,N_9524,N_9732);
nand U9910 (N_9910,N_9659,N_9697);
nand U9911 (N_9911,N_9636,N_9708);
and U9912 (N_9912,N_9662,N_9554);
xnor U9913 (N_9913,N_9506,N_9502);
nand U9914 (N_9914,N_9521,N_9664);
or U9915 (N_9915,N_9685,N_9681);
or U9916 (N_9916,N_9713,N_9658);
nand U9917 (N_9917,N_9743,N_9730);
or U9918 (N_9918,N_9671,N_9729);
nor U9919 (N_9919,N_9572,N_9658);
nand U9920 (N_9920,N_9572,N_9535);
and U9921 (N_9921,N_9693,N_9613);
nand U9922 (N_9922,N_9718,N_9689);
xor U9923 (N_9923,N_9532,N_9591);
nor U9924 (N_9924,N_9722,N_9504);
nor U9925 (N_9925,N_9737,N_9744);
and U9926 (N_9926,N_9714,N_9733);
or U9927 (N_9927,N_9575,N_9605);
nand U9928 (N_9928,N_9709,N_9500);
nor U9929 (N_9929,N_9560,N_9596);
and U9930 (N_9930,N_9599,N_9715);
and U9931 (N_9931,N_9729,N_9578);
or U9932 (N_9932,N_9579,N_9536);
and U9933 (N_9933,N_9749,N_9536);
nand U9934 (N_9934,N_9583,N_9610);
or U9935 (N_9935,N_9657,N_9594);
nand U9936 (N_9936,N_9531,N_9527);
and U9937 (N_9937,N_9576,N_9675);
nor U9938 (N_9938,N_9743,N_9551);
xnor U9939 (N_9939,N_9603,N_9534);
xnor U9940 (N_9940,N_9522,N_9679);
xor U9941 (N_9941,N_9527,N_9733);
or U9942 (N_9942,N_9635,N_9644);
nor U9943 (N_9943,N_9643,N_9573);
or U9944 (N_9944,N_9748,N_9686);
and U9945 (N_9945,N_9730,N_9544);
and U9946 (N_9946,N_9546,N_9644);
or U9947 (N_9947,N_9604,N_9551);
xnor U9948 (N_9948,N_9535,N_9742);
or U9949 (N_9949,N_9734,N_9618);
or U9950 (N_9950,N_9554,N_9547);
and U9951 (N_9951,N_9591,N_9509);
nand U9952 (N_9952,N_9688,N_9502);
nand U9953 (N_9953,N_9510,N_9544);
nand U9954 (N_9954,N_9565,N_9715);
nand U9955 (N_9955,N_9694,N_9692);
and U9956 (N_9956,N_9595,N_9609);
nand U9957 (N_9957,N_9592,N_9725);
or U9958 (N_9958,N_9724,N_9539);
xnor U9959 (N_9959,N_9503,N_9552);
and U9960 (N_9960,N_9566,N_9532);
nand U9961 (N_9961,N_9580,N_9542);
or U9962 (N_9962,N_9631,N_9717);
nor U9963 (N_9963,N_9543,N_9564);
xnor U9964 (N_9964,N_9587,N_9728);
and U9965 (N_9965,N_9673,N_9660);
or U9966 (N_9966,N_9677,N_9712);
nand U9967 (N_9967,N_9514,N_9614);
xnor U9968 (N_9968,N_9682,N_9518);
and U9969 (N_9969,N_9708,N_9739);
nand U9970 (N_9970,N_9517,N_9597);
or U9971 (N_9971,N_9571,N_9508);
or U9972 (N_9972,N_9676,N_9543);
or U9973 (N_9973,N_9670,N_9630);
or U9974 (N_9974,N_9522,N_9518);
nor U9975 (N_9975,N_9712,N_9714);
xnor U9976 (N_9976,N_9649,N_9561);
nand U9977 (N_9977,N_9554,N_9621);
and U9978 (N_9978,N_9618,N_9543);
nand U9979 (N_9979,N_9579,N_9666);
nor U9980 (N_9980,N_9562,N_9687);
nand U9981 (N_9981,N_9604,N_9526);
xor U9982 (N_9982,N_9644,N_9633);
and U9983 (N_9983,N_9716,N_9627);
and U9984 (N_9984,N_9689,N_9539);
xnor U9985 (N_9985,N_9574,N_9580);
or U9986 (N_9986,N_9536,N_9648);
nand U9987 (N_9987,N_9666,N_9553);
nor U9988 (N_9988,N_9647,N_9539);
xor U9989 (N_9989,N_9728,N_9713);
nand U9990 (N_9990,N_9672,N_9606);
or U9991 (N_9991,N_9693,N_9563);
nand U9992 (N_9992,N_9605,N_9529);
nor U9993 (N_9993,N_9538,N_9613);
xnor U9994 (N_9994,N_9672,N_9594);
or U9995 (N_9995,N_9747,N_9510);
xnor U9996 (N_9996,N_9666,N_9656);
or U9997 (N_9997,N_9669,N_9517);
nor U9998 (N_9998,N_9739,N_9748);
and U9999 (N_9999,N_9637,N_9743);
and U10000 (N_10000,N_9868,N_9957);
and U10001 (N_10001,N_9790,N_9910);
and U10002 (N_10002,N_9937,N_9890);
nor U10003 (N_10003,N_9860,N_9752);
or U10004 (N_10004,N_9961,N_9980);
xnor U10005 (N_10005,N_9884,N_9901);
and U10006 (N_10006,N_9875,N_9784);
nor U10007 (N_10007,N_9763,N_9753);
nor U10008 (N_10008,N_9789,N_9944);
nor U10009 (N_10009,N_9807,N_9833);
and U10010 (N_10010,N_9840,N_9935);
or U10011 (N_10011,N_9906,N_9873);
and U10012 (N_10012,N_9851,N_9776);
or U10013 (N_10013,N_9800,N_9773);
and U10014 (N_10014,N_9778,N_9854);
and U10015 (N_10015,N_9962,N_9923);
nand U10016 (N_10016,N_9915,N_9925);
and U10017 (N_10017,N_9827,N_9859);
and U10018 (N_10018,N_9803,N_9788);
or U10019 (N_10019,N_9755,N_9876);
and U10020 (N_10020,N_9902,N_9774);
nand U10021 (N_10021,N_9810,N_9888);
or U10022 (N_10022,N_9954,N_9899);
or U10023 (N_10023,N_9959,N_9832);
and U10024 (N_10024,N_9974,N_9964);
or U10025 (N_10025,N_9870,N_9814);
xnor U10026 (N_10026,N_9936,N_9947);
or U10027 (N_10027,N_9817,N_9751);
nand U10028 (N_10028,N_9858,N_9893);
or U10029 (N_10029,N_9783,N_9965);
or U10030 (N_10030,N_9942,N_9879);
nand U10031 (N_10031,N_9885,N_9762);
and U10032 (N_10032,N_9966,N_9927);
xnor U10033 (N_10033,N_9838,N_9819);
nor U10034 (N_10034,N_9834,N_9904);
or U10035 (N_10035,N_9795,N_9869);
or U10036 (N_10036,N_9798,N_9836);
nor U10037 (N_10037,N_9806,N_9975);
or U10038 (N_10038,N_9891,N_9772);
and U10039 (N_10039,N_9978,N_9920);
xor U10040 (N_10040,N_9958,N_9767);
or U10041 (N_10041,N_9993,N_9951);
or U10042 (N_10042,N_9837,N_9845);
and U10043 (N_10043,N_9887,N_9757);
and U10044 (N_10044,N_9995,N_9907);
nand U10045 (N_10045,N_9843,N_9997);
nor U10046 (N_10046,N_9883,N_9911);
nor U10047 (N_10047,N_9825,N_9956);
xor U10048 (N_10048,N_9897,N_9913);
or U10049 (N_10049,N_9779,N_9846);
and U10050 (N_10050,N_9786,N_9877);
or U10051 (N_10051,N_9990,N_9931);
nand U10052 (N_10052,N_9802,N_9844);
or U10053 (N_10053,N_9841,N_9945);
or U10054 (N_10054,N_9770,N_9754);
nor U10055 (N_10055,N_9797,N_9852);
nand U10056 (N_10056,N_9759,N_9792);
nand U10057 (N_10057,N_9828,N_9898);
nand U10058 (N_10058,N_9862,N_9894);
or U10059 (N_10059,N_9867,N_9924);
and U10060 (N_10060,N_9988,N_9811);
and U10061 (N_10061,N_9805,N_9801);
nor U10062 (N_10062,N_9861,N_9824);
or U10063 (N_10063,N_9874,N_9780);
xnor U10064 (N_10064,N_9812,N_9934);
nand U10065 (N_10065,N_9955,N_9967);
nand U10066 (N_10066,N_9816,N_9808);
xor U10067 (N_10067,N_9787,N_9777);
or U10068 (N_10068,N_9815,N_9865);
nor U10069 (N_10069,N_9758,N_9970);
xnor U10070 (N_10070,N_9881,N_9796);
nand U10071 (N_10071,N_9764,N_9848);
nand U10072 (N_10072,N_9820,N_9863);
nor U10073 (N_10073,N_9892,N_9775);
nor U10074 (N_10074,N_9864,N_9998);
nor U10075 (N_10075,N_9981,N_9856);
xnor U10076 (N_10076,N_9994,N_9919);
or U10077 (N_10077,N_9761,N_9765);
or U10078 (N_10078,N_9850,N_9853);
nor U10079 (N_10079,N_9982,N_9878);
nor U10080 (N_10080,N_9989,N_9791);
and U10081 (N_10081,N_9750,N_9835);
and U10082 (N_10082,N_9932,N_9922);
or U10083 (N_10083,N_9905,N_9768);
nand U10084 (N_10084,N_9909,N_9849);
xor U10085 (N_10085,N_9826,N_9926);
nor U10086 (N_10086,N_9781,N_9963);
nor U10087 (N_10087,N_9760,N_9756);
nor U10088 (N_10088,N_9979,N_9912);
or U10089 (N_10089,N_9908,N_9823);
and U10090 (N_10090,N_9950,N_9799);
and U10091 (N_10091,N_9771,N_9928);
and U10092 (N_10092,N_9992,N_9785);
or U10093 (N_10093,N_9882,N_9903);
and U10094 (N_10094,N_9896,N_9766);
nor U10095 (N_10095,N_9914,N_9933);
or U10096 (N_10096,N_9946,N_9793);
nor U10097 (N_10097,N_9822,N_9769);
and U10098 (N_10098,N_9830,N_9886);
nor U10099 (N_10099,N_9813,N_9818);
xnor U10100 (N_10100,N_9918,N_9889);
nand U10101 (N_10101,N_9999,N_9782);
nand U10102 (N_10102,N_9996,N_9917);
nand U10103 (N_10103,N_9986,N_9938);
and U10104 (N_10104,N_9976,N_9900);
and U10105 (N_10105,N_9939,N_9794);
or U10106 (N_10106,N_9977,N_9960);
or U10107 (N_10107,N_9871,N_9916);
and U10108 (N_10108,N_9949,N_9857);
and U10109 (N_10109,N_9987,N_9872);
nor U10110 (N_10110,N_9866,N_9921);
nor U10111 (N_10111,N_9831,N_9880);
nor U10112 (N_10112,N_9953,N_9985);
or U10113 (N_10113,N_9809,N_9984);
nand U10114 (N_10114,N_9971,N_9983);
or U10115 (N_10115,N_9969,N_9804);
nor U10116 (N_10116,N_9829,N_9952);
or U10117 (N_10117,N_9973,N_9842);
xnor U10118 (N_10118,N_9821,N_9895);
nor U10119 (N_10119,N_9940,N_9948);
and U10120 (N_10120,N_9941,N_9972);
or U10121 (N_10121,N_9943,N_9930);
or U10122 (N_10122,N_9929,N_9991);
or U10123 (N_10123,N_9968,N_9847);
and U10124 (N_10124,N_9855,N_9839);
and U10125 (N_10125,N_9883,N_9936);
nand U10126 (N_10126,N_9981,N_9887);
or U10127 (N_10127,N_9889,N_9963);
or U10128 (N_10128,N_9794,N_9903);
xor U10129 (N_10129,N_9794,N_9822);
nand U10130 (N_10130,N_9926,N_9781);
nand U10131 (N_10131,N_9918,N_9788);
and U10132 (N_10132,N_9992,N_9825);
or U10133 (N_10133,N_9898,N_9969);
nor U10134 (N_10134,N_9924,N_9944);
or U10135 (N_10135,N_9809,N_9822);
nand U10136 (N_10136,N_9777,N_9975);
or U10137 (N_10137,N_9992,N_9967);
or U10138 (N_10138,N_9813,N_9964);
or U10139 (N_10139,N_9850,N_9949);
nand U10140 (N_10140,N_9882,N_9906);
or U10141 (N_10141,N_9929,N_9909);
nor U10142 (N_10142,N_9863,N_9869);
nand U10143 (N_10143,N_9816,N_9751);
or U10144 (N_10144,N_9847,N_9752);
xor U10145 (N_10145,N_9985,N_9949);
nand U10146 (N_10146,N_9816,N_9934);
xnor U10147 (N_10147,N_9953,N_9947);
and U10148 (N_10148,N_9869,N_9898);
or U10149 (N_10149,N_9778,N_9795);
nor U10150 (N_10150,N_9876,N_9975);
nand U10151 (N_10151,N_9754,N_9930);
or U10152 (N_10152,N_9821,N_9919);
nor U10153 (N_10153,N_9908,N_9754);
or U10154 (N_10154,N_9998,N_9986);
or U10155 (N_10155,N_9883,N_9920);
and U10156 (N_10156,N_9808,N_9803);
or U10157 (N_10157,N_9981,N_9936);
and U10158 (N_10158,N_9972,N_9914);
and U10159 (N_10159,N_9826,N_9965);
and U10160 (N_10160,N_9811,N_9897);
xor U10161 (N_10161,N_9841,N_9802);
nand U10162 (N_10162,N_9775,N_9881);
nand U10163 (N_10163,N_9865,N_9940);
nor U10164 (N_10164,N_9892,N_9783);
or U10165 (N_10165,N_9853,N_9924);
nand U10166 (N_10166,N_9873,N_9879);
nor U10167 (N_10167,N_9947,N_9990);
nand U10168 (N_10168,N_9885,N_9773);
nor U10169 (N_10169,N_9900,N_9946);
nand U10170 (N_10170,N_9872,N_9998);
and U10171 (N_10171,N_9988,N_9926);
xnor U10172 (N_10172,N_9892,N_9877);
and U10173 (N_10173,N_9791,N_9956);
nor U10174 (N_10174,N_9924,N_9773);
and U10175 (N_10175,N_9918,N_9775);
nand U10176 (N_10176,N_9814,N_9823);
nor U10177 (N_10177,N_9912,N_9845);
and U10178 (N_10178,N_9882,N_9940);
nor U10179 (N_10179,N_9875,N_9987);
or U10180 (N_10180,N_9930,N_9794);
or U10181 (N_10181,N_9999,N_9980);
and U10182 (N_10182,N_9909,N_9993);
nor U10183 (N_10183,N_9916,N_9812);
nor U10184 (N_10184,N_9885,N_9938);
nand U10185 (N_10185,N_9841,N_9788);
and U10186 (N_10186,N_9955,N_9752);
nand U10187 (N_10187,N_9850,N_9957);
nand U10188 (N_10188,N_9860,N_9983);
nand U10189 (N_10189,N_9961,N_9793);
nor U10190 (N_10190,N_9834,N_9766);
nor U10191 (N_10191,N_9838,N_9837);
and U10192 (N_10192,N_9871,N_9944);
and U10193 (N_10193,N_9913,N_9974);
and U10194 (N_10194,N_9987,N_9922);
and U10195 (N_10195,N_9945,N_9854);
nand U10196 (N_10196,N_9869,N_9778);
nand U10197 (N_10197,N_9912,N_9806);
nor U10198 (N_10198,N_9866,N_9915);
or U10199 (N_10199,N_9765,N_9777);
nor U10200 (N_10200,N_9784,N_9907);
nand U10201 (N_10201,N_9818,N_9980);
or U10202 (N_10202,N_9827,N_9983);
or U10203 (N_10203,N_9817,N_9896);
nand U10204 (N_10204,N_9841,N_9823);
nand U10205 (N_10205,N_9929,N_9932);
nand U10206 (N_10206,N_9891,N_9810);
or U10207 (N_10207,N_9887,N_9825);
or U10208 (N_10208,N_9929,N_9806);
and U10209 (N_10209,N_9859,N_9856);
nor U10210 (N_10210,N_9870,N_9778);
nand U10211 (N_10211,N_9788,N_9845);
nand U10212 (N_10212,N_9824,N_9771);
nand U10213 (N_10213,N_9846,N_9836);
nor U10214 (N_10214,N_9773,N_9890);
nor U10215 (N_10215,N_9784,N_9873);
nand U10216 (N_10216,N_9885,N_9845);
and U10217 (N_10217,N_9906,N_9796);
and U10218 (N_10218,N_9900,N_9845);
or U10219 (N_10219,N_9816,N_9757);
or U10220 (N_10220,N_9979,N_9753);
nor U10221 (N_10221,N_9797,N_9851);
nor U10222 (N_10222,N_9953,N_9760);
nand U10223 (N_10223,N_9869,N_9756);
or U10224 (N_10224,N_9957,N_9955);
or U10225 (N_10225,N_9831,N_9866);
nor U10226 (N_10226,N_9825,N_9978);
nor U10227 (N_10227,N_9752,N_9776);
or U10228 (N_10228,N_9887,N_9882);
nor U10229 (N_10229,N_9960,N_9895);
and U10230 (N_10230,N_9788,N_9864);
nand U10231 (N_10231,N_9966,N_9874);
nand U10232 (N_10232,N_9807,N_9835);
or U10233 (N_10233,N_9826,N_9980);
nand U10234 (N_10234,N_9868,N_9813);
and U10235 (N_10235,N_9783,N_9776);
xnor U10236 (N_10236,N_9799,N_9796);
nor U10237 (N_10237,N_9930,N_9985);
and U10238 (N_10238,N_9817,N_9796);
nand U10239 (N_10239,N_9961,N_9903);
and U10240 (N_10240,N_9920,N_9874);
and U10241 (N_10241,N_9840,N_9801);
nor U10242 (N_10242,N_9864,N_9881);
nand U10243 (N_10243,N_9784,N_9930);
or U10244 (N_10244,N_9913,N_9904);
nand U10245 (N_10245,N_9938,N_9931);
and U10246 (N_10246,N_9932,N_9833);
nand U10247 (N_10247,N_9800,N_9876);
or U10248 (N_10248,N_9997,N_9886);
nor U10249 (N_10249,N_9876,N_9753);
nand U10250 (N_10250,N_10094,N_10072);
nand U10251 (N_10251,N_10240,N_10249);
nor U10252 (N_10252,N_10031,N_10160);
nor U10253 (N_10253,N_10174,N_10211);
nor U10254 (N_10254,N_10025,N_10044);
or U10255 (N_10255,N_10047,N_10048);
nand U10256 (N_10256,N_10041,N_10117);
xnor U10257 (N_10257,N_10054,N_10177);
nor U10258 (N_10258,N_10104,N_10149);
and U10259 (N_10259,N_10195,N_10120);
or U10260 (N_10260,N_10126,N_10171);
or U10261 (N_10261,N_10096,N_10034);
or U10262 (N_10262,N_10085,N_10119);
or U10263 (N_10263,N_10227,N_10093);
nand U10264 (N_10264,N_10183,N_10038);
nor U10265 (N_10265,N_10087,N_10156);
and U10266 (N_10266,N_10222,N_10193);
nor U10267 (N_10267,N_10151,N_10216);
nand U10268 (N_10268,N_10073,N_10059);
nand U10269 (N_10269,N_10238,N_10144);
and U10270 (N_10270,N_10112,N_10239);
nand U10271 (N_10271,N_10192,N_10131);
nand U10272 (N_10272,N_10134,N_10065);
or U10273 (N_10273,N_10001,N_10109);
nand U10274 (N_10274,N_10116,N_10184);
or U10275 (N_10275,N_10063,N_10080);
nand U10276 (N_10276,N_10046,N_10143);
and U10277 (N_10277,N_10005,N_10033);
nor U10278 (N_10278,N_10217,N_10178);
or U10279 (N_10279,N_10081,N_10092);
nand U10280 (N_10280,N_10146,N_10215);
nand U10281 (N_10281,N_10245,N_10152);
nand U10282 (N_10282,N_10069,N_10039);
or U10283 (N_10283,N_10032,N_10235);
nor U10284 (N_10284,N_10064,N_10020);
xor U10285 (N_10285,N_10051,N_10074);
or U10286 (N_10286,N_10127,N_10075);
nand U10287 (N_10287,N_10004,N_10084);
nor U10288 (N_10288,N_10237,N_10050);
nor U10289 (N_10289,N_10002,N_10141);
or U10290 (N_10290,N_10228,N_10089);
or U10291 (N_10291,N_10107,N_10016);
nor U10292 (N_10292,N_10169,N_10187);
nor U10293 (N_10293,N_10147,N_10088);
and U10294 (N_10294,N_10091,N_10139);
nand U10295 (N_10295,N_10021,N_10132);
nor U10296 (N_10296,N_10148,N_10138);
nand U10297 (N_10297,N_10199,N_10225);
nand U10298 (N_10298,N_10142,N_10057);
nand U10299 (N_10299,N_10202,N_10076);
nand U10300 (N_10300,N_10018,N_10232);
or U10301 (N_10301,N_10231,N_10121);
or U10302 (N_10302,N_10223,N_10035);
nand U10303 (N_10303,N_10155,N_10200);
nand U10304 (N_10304,N_10026,N_10172);
xnor U10305 (N_10305,N_10095,N_10077);
nor U10306 (N_10306,N_10067,N_10168);
nand U10307 (N_10307,N_10060,N_10029);
xor U10308 (N_10308,N_10049,N_10037);
xor U10309 (N_10309,N_10179,N_10164);
or U10310 (N_10310,N_10158,N_10090);
xor U10311 (N_10311,N_10201,N_10111);
xor U10312 (N_10312,N_10175,N_10115);
or U10313 (N_10313,N_10113,N_10097);
and U10314 (N_10314,N_10180,N_10043);
and U10315 (N_10315,N_10166,N_10203);
or U10316 (N_10316,N_10230,N_10040);
nand U10317 (N_10317,N_10189,N_10086);
nand U10318 (N_10318,N_10123,N_10098);
or U10319 (N_10319,N_10246,N_10224);
nor U10320 (N_10320,N_10102,N_10182);
nor U10321 (N_10321,N_10150,N_10114);
and U10322 (N_10322,N_10003,N_10011);
nand U10323 (N_10323,N_10130,N_10161);
nor U10324 (N_10324,N_10083,N_10024);
and U10325 (N_10325,N_10218,N_10071);
and U10326 (N_10326,N_10030,N_10068);
nand U10327 (N_10327,N_10248,N_10214);
nand U10328 (N_10328,N_10197,N_10145);
or U10329 (N_10329,N_10101,N_10106);
xnor U10330 (N_10330,N_10221,N_10219);
and U10331 (N_10331,N_10122,N_10000);
nor U10332 (N_10332,N_10017,N_10165);
xor U10333 (N_10333,N_10052,N_10194);
nor U10334 (N_10334,N_10061,N_10108);
and U10335 (N_10335,N_10066,N_10153);
or U10336 (N_10336,N_10007,N_10170);
nor U10337 (N_10337,N_10208,N_10236);
and U10338 (N_10338,N_10210,N_10062);
xnor U10339 (N_10339,N_10055,N_10176);
or U10340 (N_10340,N_10206,N_10118);
or U10341 (N_10341,N_10205,N_10014);
or U10342 (N_10342,N_10188,N_10078);
xor U10343 (N_10343,N_10053,N_10128);
xor U10344 (N_10344,N_10162,N_10082);
nand U10345 (N_10345,N_10181,N_10100);
and U10346 (N_10346,N_10209,N_10042);
or U10347 (N_10347,N_10213,N_10009);
nor U10348 (N_10348,N_10028,N_10137);
nand U10349 (N_10349,N_10015,N_10207);
xor U10350 (N_10350,N_10212,N_10022);
xnor U10351 (N_10351,N_10110,N_10159);
or U10352 (N_10352,N_10129,N_10190);
xor U10353 (N_10353,N_10079,N_10105);
or U10354 (N_10354,N_10241,N_10185);
nand U10355 (N_10355,N_10135,N_10229);
or U10356 (N_10356,N_10013,N_10019);
nor U10357 (N_10357,N_10244,N_10186);
xor U10358 (N_10358,N_10233,N_10234);
and U10359 (N_10359,N_10196,N_10242);
nor U10360 (N_10360,N_10226,N_10220);
nand U10361 (N_10361,N_10012,N_10103);
nor U10362 (N_10362,N_10247,N_10133);
nor U10363 (N_10363,N_10204,N_10140);
or U10364 (N_10364,N_10006,N_10023);
xor U10365 (N_10365,N_10027,N_10125);
and U10366 (N_10366,N_10163,N_10198);
nand U10367 (N_10367,N_10056,N_10036);
and U10368 (N_10368,N_10154,N_10243);
nor U10369 (N_10369,N_10045,N_10010);
xor U10370 (N_10370,N_10191,N_10058);
or U10371 (N_10371,N_10157,N_10136);
nand U10372 (N_10372,N_10070,N_10099);
or U10373 (N_10373,N_10008,N_10167);
xor U10374 (N_10374,N_10124,N_10173);
and U10375 (N_10375,N_10245,N_10019);
nor U10376 (N_10376,N_10222,N_10014);
nand U10377 (N_10377,N_10033,N_10133);
nor U10378 (N_10378,N_10124,N_10233);
nor U10379 (N_10379,N_10044,N_10037);
and U10380 (N_10380,N_10114,N_10243);
nor U10381 (N_10381,N_10051,N_10123);
nand U10382 (N_10382,N_10066,N_10240);
nor U10383 (N_10383,N_10200,N_10009);
and U10384 (N_10384,N_10021,N_10057);
or U10385 (N_10385,N_10128,N_10134);
or U10386 (N_10386,N_10188,N_10126);
and U10387 (N_10387,N_10068,N_10057);
or U10388 (N_10388,N_10094,N_10235);
or U10389 (N_10389,N_10010,N_10211);
xnor U10390 (N_10390,N_10061,N_10019);
and U10391 (N_10391,N_10097,N_10143);
xnor U10392 (N_10392,N_10185,N_10207);
or U10393 (N_10393,N_10134,N_10215);
nand U10394 (N_10394,N_10172,N_10011);
nand U10395 (N_10395,N_10166,N_10094);
nand U10396 (N_10396,N_10072,N_10122);
nor U10397 (N_10397,N_10008,N_10186);
or U10398 (N_10398,N_10190,N_10035);
nor U10399 (N_10399,N_10115,N_10024);
or U10400 (N_10400,N_10120,N_10122);
nand U10401 (N_10401,N_10158,N_10241);
nor U10402 (N_10402,N_10039,N_10000);
or U10403 (N_10403,N_10158,N_10215);
xnor U10404 (N_10404,N_10025,N_10162);
and U10405 (N_10405,N_10038,N_10130);
or U10406 (N_10406,N_10016,N_10114);
nor U10407 (N_10407,N_10069,N_10073);
xor U10408 (N_10408,N_10243,N_10019);
nor U10409 (N_10409,N_10159,N_10096);
nor U10410 (N_10410,N_10019,N_10133);
nand U10411 (N_10411,N_10142,N_10127);
or U10412 (N_10412,N_10114,N_10013);
and U10413 (N_10413,N_10229,N_10176);
nand U10414 (N_10414,N_10075,N_10072);
nand U10415 (N_10415,N_10061,N_10075);
nand U10416 (N_10416,N_10061,N_10030);
and U10417 (N_10417,N_10179,N_10177);
or U10418 (N_10418,N_10013,N_10159);
xor U10419 (N_10419,N_10201,N_10099);
nand U10420 (N_10420,N_10032,N_10089);
nand U10421 (N_10421,N_10225,N_10162);
and U10422 (N_10422,N_10058,N_10227);
or U10423 (N_10423,N_10093,N_10139);
nor U10424 (N_10424,N_10015,N_10095);
or U10425 (N_10425,N_10224,N_10105);
nor U10426 (N_10426,N_10097,N_10099);
xor U10427 (N_10427,N_10249,N_10087);
nor U10428 (N_10428,N_10038,N_10057);
nand U10429 (N_10429,N_10018,N_10230);
nor U10430 (N_10430,N_10216,N_10121);
or U10431 (N_10431,N_10129,N_10109);
or U10432 (N_10432,N_10045,N_10033);
or U10433 (N_10433,N_10202,N_10012);
and U10434 (N_10434,N_10142,N_10172);
nor U10435 (N_10435,N_10242,N_10162);
or U10436 (N_10436,N_10166,N_10232);
xor U10437 (N_10437,N_10123,N_10172);
xor U10438 (N_10438,N_10051,N_10217);
and U10439 (N_10439,N_10111,N_10218);
nand U10440 (N_10440,N_10242,N_10062);
and U10441 (N_10441,N_10194,N_10030);
nand U10442 (N_10442,N_10118,N_10031);
nor U10443 (N_10443,N_10232,N_10019);
or U10444 (N_10444,N_10101,N_10130);
nor U10445 (N_10445,N_10217,N_10235);
or U10446 (N_10446,N_10031,N_10028);
nand U10447 (N_10447,N_10126,N_10128);
nor U10448 (N_10448,N_10030,N_10118);
or U10449 (N_10449,N_10220,N_10206);
and U10450 (N_10450,N_10016,N_10105);
nor U10451 (N_10451,N_10059,N_10149);
nor U10452 (N_10452,N_10193,N_10019);
nor U10453 (N_10453,N_10004,N_10083);
and U10454 (N_10454,N_10160,N_10111);
nand U10455 (N_10455,N_10089,N_10065);
and U10456 (N_10456,N_10035,N_10174);
nor U10457 (N_10457,N_10129,N_10231);
nor U10458 (N_10458,N_10229,N_10139);
and U10459 (N_10459,N_10204,N_10208);
xnor U10460 (N_10460,N_10038,N_10007);
or U10461 (N_10461,N_10019,N_10157);
and U10462 (N_10462,N_10155,N_10107);
nand U10463 (N_10463,N_10189,N_10070);
or U10464 (N_10464,N_10099,N_10040);
and U10465 (N_10465,N_10046,N_10162);
and U10466 (N_10466,N_10051,N_10198);
or U10467 (N_10467,N_10176,N_10230);
and U10468 (N_10468,N_10084,N_10221);
and U10469 (N_10469,N_10146,N_10221);
nor U10470 (N_10470,N_10145,N_10059);
or U10471 (N_10471,N_10049,N_10222);
xor U10472 (N_10472,N_10168,N_10015);
nor U10473 (N_10473,N_10001,N_10152);
and U10474 (N_10474,N_10241,N_10144);
or U10475 (N_10475,N_10186,N_10090);
nand U10476 (N_10476,N_10106,N_10159);
and U10477 (N_10477,N_10100,N_10237);
xor U10478 (N_10478,N_10228,N_10245);
nand U10479 (N_10479,N_10204,N_10143);
nand U10480 (N_10480,N_10148,N_10219);
and U10481 (N_10481,N_10200,N_10003);
nor U10482 (N_10482,N_10127,N_10198);
and U10483 (N_10483,N_10208,N_10247);
or U10484 (N_10484,N_10152,N_10122);
nand U10485 (N_10485,N_10146,N_10123);
or U10486 (N_10486,N_10011,N_10237);
and U10487 (N_10487,N_10236,N_10240);
nand U10488 (N_10488,N_10080,N_10246);
or U10489 (N_10489,N_10046,N_10097);
nand U10490 (N_10490,N_10124,N_10009);
nand U10491 (N_10491,N_10032,N_10009);
or U10492 (N_10492,N_10164,N_10104);
nand U10493 (N_10493,N_10222,N_10008);
and U10494 (N_10494,N_10228,N_10068);
nor U10495 (N_10495,N_10093,N_10071);
and U10496 (N_10496,N_10170,N_10152);
nor U10497 (N_10497,N_10221,N_10108);
or U10498 (N_10498,N_10150,N_10043);
nor U10499 (N_10499,N_10187,N_10076);
nor U10500 (N_10500,N_10489,N_10411);
or U10501 (N_10501,N_10342,N_10335);
nand U10502 (N_10502,N_10377,N_10472);
nand U10503 (N_10503,N_10430,N_10418);
and U10504 (N_10504,N_10269,N_10436);
or U10505 (N_10505,N_10390,N_10284);
nor U10506 (N_10506,N_10258,N_10408);
nor U10507 (N_10507,N_10406,N_10289);
xnor U10508 (N_10508,N_10362,N_10355);
and U10509 (N_10509,N_10407,N_10415);
or U10510 (N_10510,N_10348,N_10290);
or U10511 (N_10511,N_10426,N_10403);
nor U10512 (N_10512,N_10275,N_10378);
nor U10513 (N_10513,N_10404,N_10419);
xnor U10514 (N_10514,N_10259,N_10320);
nor U10515 (N_10515,N_10280,N_10402);
and U10516 (N_10516,N_10484,N_10324);
or U10517 (N_10517,N_10424,N_10434);
or U10518 (N_10518,N_10340,N_10344);
nand U10519 (N_10519,N_10497,N_10343);
or U10520 (N_10520,N_10447,N_10360);
and U10521 (N_10521,N_10492,N_10277);
and U10522 (N_10522,N_10416,N_10410);
nor U10523 (N_10523,N_10391,N_10261);
and U10524 (N_10524,N_10483,N_10444);
and U10525 (N_10525,N_10322,N_10413);
nand U10526 (N_10526,N_10262,N_10253);
xnor U10527 (N_10527,N_10471,N_10432);
nand U10528 (N_10528,N_10329,N_10414);
nand U10529 (N_10529,N_10487,N_10482);
or U10530 (N_10530,N_10496,N_10442);
xor U10531 (N_10531,N_10385,N_10481);
or U10532 (N_10532,N_10267,N_10372);
nand U10533 (N_10533,N_10450,N_10417);
or U10534 (N_10534,N_10465,N_10468);
nor U10535 (N_10535,N_10271,N_10421);
nand U10536 (N_10536,N_10431,N_10333);
nor U10537 (N_10537,N_10376,N_10396);
nor U10538 (N_10538,N_10452,N_10293);
nor U10539 (N_10539,N_10374,N_10282);
or U10540 (N_10540,N_10494,N_10316);
nand U10541 (N_10541,N_10351,N_10347);
xnor U10542 (N_10542,N_10443,N_10306);
or U10543 (N_10543,N_10332,N_10327);
nand U10544 (N_10544,N_10281,N_10254);
nand U10545 (N_10545,N_10305,N_10429);
and U10546 (N_10546,N_10462,N_10346);
and U10547 (N_10547,N_10479,N_10476);
nand U10548 (N_10548,N_10457,N_10321);
or U10549 (N_10549,N_10455,N_10393);
and U10550 (N_10550,N_10400,N_10279);
nor U10551 (N_10551,N_10345,N_10394);
or U10552 (N_10552,N_10311,N_10485);
and U10553 (N_10553,N_10260,N_10428);
nand U10554 (N_10554,N_10466,N_10353);
nand U10555 (N_10555,N_10359,N_10383);
xor U10556 (N_10556,N_10312,N_10274);
and U10557 (N_10557,N_10272,N_10463);
and U10558 (N_10558,N_10338,N_10257);
nand U10559 (N_10559,N_10326,N_10368);
or U10560 (N_10560,N_10303,N_10300);
or U10561 (N_10561,N_10422,N_10364);
or U10562 (N_10562,N_10296,N_10265);
nand U10563 (N_10563,N_10409,N_10352);
and U10564 (N_10564,N_10297,N_10461);
nor U10565 (N_10565,N_10401,N_10298);
and U10566 (N_10566,N_10323,N_10474);
nor U10567 (N_10567,N_10314,N_10301);
and U10568 (N_10568,N_10273,N_10367);
xnor U10569 (N_10569,N_10365,N_10435);
xnor U10570 (N_10570,N_10423,N_10308);
nand U10571 (N_10571,N_10339,N_10325);
nand U10572 (N_10572,N_10349,N_10315);
or U10573 (N_10573,N_10366,N_10491);
nor U10574 (N_10574,N_10486,N_10460);
nand U10575 (N_10575,N_10439,N_10412);
or U10576 (N_10576,N_10251,N_10373);
xor U10577 (N_10577,N_10310,N_10469);
nor U10578 (N_10578,N_10398,N_10445);
nand U10579 (N_10579,N_10456,N_10295);
or U10580 (N_10580,N_10294,N_10341);
nor U10581 (N_10581,N_10438,N_10490);
nand U10582 (N_10582,N_10256,N_10255);
nor U10583 (N_10583,N_10382,N_10287);
and U10584 (N_10584,N_10464,N_10381);
and U10585 (N_10585,N_10425,N_10337);
nand U10586 (N_10586,N_10328,N_10473);
and U10587 (N_10587,N_10389,N_10285);
and U10588 (N_10588,N_10299,N_10331);
nor U10589 (N_10589,N_10356,N_10369);
or U10590 (N_10590,N_10470,N_10350);
or U10591 (N_10591,N_10371,N_10270);
nand U10592 (N_10592,N_10375,N_10475);
or U10593 (N_10593,N_10453,N_10252);
nor U10594 (N_10594,N_10478,N_10399);
nor U10595 (N_10595,N_10334,N_10358);
or U10596 (N_10596,N_10397,N_10427);
xor U10597 (N_10597,N_10441,N_10307);
and U10598 (N_10598,N_10467,N_10302);
or U10599 (N_10599,N_10458,N_10488);
nand U10600 (N_10600,N_10283,N_10264);
xnor U10601 (N_10601,N_10268,N_10379);
xnor U10602 (N_10602,N_10354,N_10493);
nor U10603 (N_10603,N_10370,N_10313);
nor U10604 (N_10604,N_10437,N_10459);
or U10605 (N_10605,N_10357,N_10336);
xor U10606 (N_10606,N_10392,N_10405);
or U10607 (N_10607,N_10250,N_10449);
or U10608 (N_10608,N_10361,N_10498);
nor U10609 (N_10609,N_10278,N_10451);
or U10610 (N_10610,N_10477,N_10387);
and U10611 (N_10611,N_10319,N_10495);
nor U10612 (N_10612,N_10395,N_10433);
and U10613 (N_10613,N_10292,N_10263);
or U10614 (N_10614,N_10420,N_10291);
nand U10615 (N_10615,N_10386,N_10499);
nand U10616 (N_10616,N_10318,N_10286);
nand U10617 (N_10617,N_10304,N_10330);
xor U10618 (N_10618,N_10317,N_10480);
nor U10619 (N_10619,N_10363,N_10454);
and U10620 (N_10620,N_10309,N_10288);
and U10621 (N_10621,N_10276,N_10388);
xnor U10622 (N_10622,N_10380,N_10266);
nand U10623 (N_10623,N_10446,N_10384);
nand U10624 (N_10624,N_10440,N_10448);
or U10625 (N_10625,N_10311,N_10318);
or U10626 (N_10626,N_10329,N_10292);
and U10627 (N_10627,N_10372,N_10391);
or U10628 (N_10628,N_10301,N_10277);
nor U10629 (N_10629,N_10287,N_10270);
nor U10630 (N_10630,N_10261,N_10392);
or U10631 (N_10631,N_10407,N_10350);
or U10632 (N_10632,N_10329,N_10478);
nor U10633 (N_10633,N_10439,N_10471);
nand U10634 (N_10634,N_10490,N_10318);
nor U10635 (N_10635,N_10355,N_10438);
nand U10636 (N_10636,N_10435,N_10326);
xor U10637 (N_10637,N_10364,N_10332);
nand U10638 (N_10638,N_10360,N_10435);
or U10639 (N_10639,N_10454,N_10350);
nand U10640 (N_10640,N_10398,N_10472);
nor U10641 (N_10641,N_10377,N_10420);
or U10642 (N_10642,N_10364,N_10495);
and U10643 (N_10643,N_10359,N_10328);
or U10644 (N_10644,N_10319,N_10437);
nand U10645 (N_10645,N_10274,N_10347);
xor U10646 (N_10646,N_10372,N_10407);
nand U10647 (N_10647,N_10499,N_10282);
or U10648 (N_10648,N_10258,N_10495);
and U10649 (N_10649,N_10385,N_10364);
nor U10650 (N_10650,N_10345,N_10379);
nor U10651 (N_10651,N_10400,N_10282);
and U10652 (N_10652,N_10281,N_10291);
nor U10653 (N_10653,N_10274,N_10437);
nor U10654 (N_10654,N_10427,N_10408);
and U10655 (N_10655,N_10270,N_10310);
xnor U10656 (N_10656,N_10354,N_10454);
and U10657 (N_10657,N_10360,N_10436);
or U10658 (N_10658,N_10479,N_10460);
or U10659 (N_10659,N_10336,N_10377);
or U10660 (N_10660,N_10364,N_10383);
or U10661 (N_10661,N_10415,N_10281);
nand U10662 (N_10662,N_10324,N_10486);
and U10663 (N_10663,N_10476,N_10279);
nor U10664 (N_10664,N_10482,N_10328);
and U10665 (N_10665,N_10479,N_10466);
nor U10666 (N_10666,N_10398,N_10382);
or U10667 (N_10667,N_10302,N_10427);
xor U10668 (N_10668,N_10399,N_10279);
nor U10669 (N_10669,N_10293,N_10385);
and U10670 (N_10670,N_10380,N_10475);
nor U10671 (N_10671,N_10356,N_10269);
or U10672 (N_10672,N_10431,N_10336);
nand U10673 (N_10673,N_10486,N_10493);
nor U10674 (N_10674,N_10420,N_10491);
nor U10675 (N_10675,N_10313,N_10430);
and U10676 (N_10676,N_10299,N_10367);
nor U10677 (N_10677,N_10356,N_10489);
and U10678 (N_10678,N_10387,N_10463);
nand U10679 (N_10679,N_10404,N_10286);
nor U10680 (N_10680,N_10444,N_10283);
and U10681 (N_10681,N_10491,N_10360);
xor U10682 (N_10682,N_10388,N_10269);
nand U10683 (N_10683,N_10393,N_10408);
nor U10684 (N_10684,N_10338,N_10309);
xnor U10685 (N_10685,N_10315,N_10401);
or U10686 (N_10686,N_10395,N_10479);
or U10687 (N_10687,N_10379,N_10397);
or U10688 (N_10688,N_10324,N_10352);
or U10689 (N_10689,N_10435,N_10281);
nor U10690 (N_10690,N_10350,N_10348);
xor U10691 (N_10691,N_10351,N_10498);
xnor U10692 (N_10692,N_10268,N_10377);
nor U10693 (N_10693,N_10408,N_10308);
nand U10694 (N_10694,N_10253,N_10402);
nor U10695 (N_10695,N_10412,N_10440);
nor U10696 (N_10696,N_10348,N_10297);
nor U10697 (N_10697,N_10289,N_10337);
nor U10698 (N_10698,N_10451,N_10293);
nor U10699 (N_10699,N_10314,N_10331);
and U10700 (N_10700,N_10257,N_10360);
xor U10701 (N_10701,N_10359,N_10338);
nand U10702 (N_10702,N_10360,N_10426);
nor U10703 (N_10703,N_10250,N_10486);
xnor U10704 (N_10704,N_10437,N_10360);
nand U10705 (N_10705,N_10364,N_10251);
nor U10706 (N_10706,N_10334,N_10310);
or U10707 (N_10707,N_10479,N_10488);
and U10708 (N_10708,N_10347,N_10325);
or U10709 (N_10709,N_10324,N_10448);
and U10710 (N_10710,N_10465,N_10377);
nor U10711 (N_10711,N_10250,N_10403);
or U10712 (N_10712,N_10294,N_10383);
xnor U10713 (N_10713,N_10394,N_10327);
nand U10714 (N_10714,N_10495,N_10480);
or U10715 (N_10715,N_10358,N_10443);
xor U10716 (N_10716,N_10347,N_10436);
and U10717 (N_10717,N_10348,N_10498);
xnor U10718 (N_10718,N_10409,N_10468);
and U10719 (N_10719,N_10481,N_10305);
nand U10720 (N_10720,N_10420,N_10461);
or U10721 (N_10721,N_10288,N_10290);
and U10722 (N_10722,N_10491,N_10469);
and U10723 (N_10723,N_10385,N_10429);
and U10724 (N_10724,N_10376,N_10285);
and U10725 (N_10725,N_10401,N_10254);
or U10726 (N_10726,N_10290,N_10399);
or U10727 (N_10727,N_10317,N_10283);
nor U10728 (N_10728,N_10490,N_10388);
nor U10729 (N_10729,N_10410,N_10401);
or U10730 (N_10730,N_10252,N_10302);
nor U10731 (N_10731,N_10301,N_10384);
and U10732 (N_10732,N_10358,N_10491);
xor U10733 (N_10733,N_10434,N_10375);
and U10734 (N_10734,N_10447,N_10277);
and U10735 (N_10735,N_10462,N_10345);
and U10736 (N_10736,N_10266,N_10406);
nor U10737 (N_10737,N_10286,N_10490);
nor U10738 (N_10738,N_10491,N_10365);
xnor U10739 (N_10739,N_10394,N_10354);
or U10740 (N_10740,N_10361,N_10445);
nor U10741 (N_10741,N_10324,N_10464);
or U10742 (N_10742,N_10287,N_10445);
nor U10743 (N_10743,N_10413,N_10258);
or U10744 (N_10744,N_10467,N_10329);
xor U10745 (N_10745,N_10409,N_10262);
xnor U10746 (N_10746,N_10485,N_10433);
and U10747 (N_10747,N_10405,N_10498);
or U10748 (N_10748,N_10434,N_10251);
and U10749 (N_10749,N_10360,N_10355);
and U10750 (N_10750,N_10610,N_10629);
and U10751 (N_10751,N_10500,N_10740);
and U10752 (N_10752,N_10552,N_10683);
xor U10753 (N_10753,N_10592,N_10524);
and U10754 (N_10754,N_10677,N_10518);
and U10755 (N_10755,N_10727,N_10655);
nor U10756 (N_10756,N_10643,N_10719);
nand U10757 (N_10757,N_10598,N_10690);
nor U10758 (N_10758,N_10634,N_10558);
nor U10759 (N_10759,N_10584,N_10517);
nand U10760 (N_10760,N_10545,N_10611);
or U10761 (N_10761,N_10506,N_10580);
nor U10762 (N_10762,N_10691,N_10746);
or U10763 (N_10763,N_10652,N_10637);
or U10764 (N_10764,N_10623,N_10555);
xnor U10765 (N_10765,N_10734,N_10559);
and U10766 (N_10766,N_10653,N_10508);
and U10767 (N_10767,N_10704,N_10705);
or U10768 (N_10768,N_10701,N_10586);
or U10769 (N_10769,N_10659,N_10603);
nand U10770 (N_10770,N_10697,N_10692);
and U10771 (N_10771,N_10729,N_10671);
nor U10772 (N_10772,N_10614,N_10544);
nor U10773 (N_10773,N_10503,N_10560);
nand U10774 (N_10774,N_10654,N_10732);
nor U10775 (N_10775,N_10522,N_10672);
nor U10776 (N_10776,N_10514,N_10718);
nor U10777 (N_10777,N_10636,N_10622);
nor U10778 (N_10778,N_10561,N_10707);
and U10779 (N_10779,N_10700,N_10681);
xor U10780 (N_10780,N_10717,N_10650);
nor U10781 (N_10781,N_10733,N_10702);
nand U10782 (N_10782,N_10585,N_10670);
nor U10783 (N_10783,N_10535,N_10641);
nand U10784 (N_10784,N_10696,N_10533);
xnor U10785 (N_10785,N_10620,N_10512);
nand U10786 (N_10786,N_10538,N_10649);
nand U10787 (N_10787,N_10712,N_10599);
xnor U10788 (N_10788,N_10617,N_10627);
nand U10789 (N_10789,N_10534,N_10630);
and U10790 (N_10790,N_10651,N_10725);
or U10791 (N_10791,N_10747,N_10541);
nand U10792 (N_10792,N_10529,N_10749);
and U10793 (N_10793,N_10742,N_10549);
xnor U10794 (N_10794,N_10674,N_10721);
and U10795 (N_10795,N_10590,N_10642);
or U10796 (N_10796,N_10745,N_10602);
nand U10797 (N_10797,N_10635,N_10633);
nand U10798 (N_10798,N_10527,N_10539);
and U10799 (N_10799,N_10647,N_10507);
nand U10800 (N_10800,N_10713,N_10684);
nor U10801 (N_10801,N_10574,N_10588);
nor U10802 (N_10802,N_10613,N_10525);
xnor U10803 (N_10803,N_10710,N_10581);
nor U10804 (N_10804,N_10577,N_10660);
nor U10805 (N_10805,N_10743,N_10706);
nand U10806 (N_10806,N_10669,N_10516);
nand U10807 (N_10807,N_10736,N_10587);
or U10808 (N_10808,N_10509,N_10606);
or U10809 (N_10809,N_10521,N_10565);
or U10810 (N_10810,N_10703,N_10553);
nor U10811 (N_10811,N_10626,N_10644);
or U10812 (N_10812,N_10738,N_10505);
nand U10813 (N_10813,N_10724,N_10609);
and U10814 (N_10814,N_10576,N_10739);
nand U10815 (N_10815,N_10638,N_10583);
or U10816 (N_10816,N_10694,N_10531);
and U10817 (N_10817,N_10511,N_10663);
and U10818 (N_10818,N_10666,N_10667);
nor U10819 (N_10819,N_10612,N_10688);
or U10820 (N_10820,N_10564,N_10720);
and U10821 (N_10821,N_10673,N_10708);
nor U10822 (N_10822,N_10591,N_10569);
nand U10823 (N_10823,N_10748,N_10556);
nand U10824 (N_10824,N_10693,N_10658);
and U10825 (N_10825,N_10741,N_10520);
xor U10826 (N_10826,N_10526,N_10571);
and U10827 (N_10827,N_10657,N_10523);
xnor U10828 (N_10828,N_10711,N_10709);
or U10829 (N_10829,N_10595,N_10607);
or U10830 (N_10830,N_10605,N_10536);
and U10831 (N_10831,N_10624,N_10664);
and U10832 (N_10832,N_10735,N_10625);
nor U10833 (N_10833,N_10715,N_10716);
nor U10834 (N_10834,N_10578,N_10679);
nor U10835 (N_10835,N_10668,N_10730);
or U10836 (N_10836,N_10563,N_10550);
nor U10837 (N_10837,N_10551,N_10618);
xor U10838 (N_10838,N_10723,N_10615);
nor U10839 (N_10839,N_10737,N_10695);
or U10840 (N_10840,N_10680,N_10686);
nor U10841 (N_10841,N_10665,N_10597);
or U10842 (N_10842,N_10582,N_10596);
nor U10843 (N_10843,N_10601,N_10604);
or U10844 (N_10844,N_10519,N_10510);
xor U10845 (N_10845,N_10744,N_10513);
nand U10846 (N_10846,N_10573,N_10567);
and U10847 (N_10847,N_10502,N_10554);
nand U10848 (N_10848,N_10540,N_10648);
nor U10849 (N_10849,N_10728,N_10714);
and U10850 (N_10850,N_10557,N_10656);
nor U10851 (N_10851,N_10528,N_10676);
xor U10852 (N_10852,N_10621,N_10646);
nor U10853 (N_10853,N_10678,N_10542);
nor U10854 (N_10854,N_10532,N_10568);
or U10855 (N_10855,N_10530,N_10628);
or U10856 (N_10856,N_10661,N_10639);
nand U10857 (N_10857,N_10537,N_10698);
nor U10858 (N_10858,N_10546,N_10731);
nand U10859 (N_10859,N_10685,N_10675);
and U10860 (N_10860,N_10589,N_10547);
nand U10861 (N_10861,N_10699,N_10570);
nand U10862 (N_10862,N_10631,N_10501);
and U10863 (N_10863,N_10645,N_10515);
and U10864 (N_10864,N_10600,N_10662);
nor U10865 (N_10865,N_10566,N_10593);
nand U10866 (N_10866,N_10543,N_10572);
or U10867 (N_10867,N_10579,N_10619);
and U10868 (N_10868,N_10722,N_10687);
nor U10869 (N_10869,N_10682,N_10689);
nor U10870 (N_10870,N_10562,N_10548);
or U10871 (N_10871,N_10594,N_10640);
or U10872 (N_10872,N_10632,N_10575);
xor U10873 (N_10873,N_10616,N_10726);
nor U10874 (N_10874,N_10608,N_10504);
xnor U10875 (N_10875,N_10508,N_10627);
nand U10876 (N_10876,N_10679,N_10705);
and U10877 (N_10877,N_10525,N_10547);
xor U10878 (N_10878,N_10740,N_10688);
nand U10879 (N_10879,N_10731,N_10719);
or U10880 (N_10880,N_10725,N_10717);
and U10881 (N_10881,N_10644,N_10512);
and U10882 (N_10882,N_10686,N_10538);
xnor U10883 (N_10883,N_10737,N_10667);
nor U10884 (N_10884,N_10556,N_10592);
xnor U10885 (N_10885,N_10619,N_10716);
or U10886 (N_10886,N_10719,N_10603);
or U10887 (N_10887,N_10681,N_10619);
nor U10888 (N_10888,N_10620,N_10542);
or U10889 (N_10889,N_10569,N_10667);
and U10890 (N_10890,N_10691,N_10707);
nor U10891 (N_10891,N_10509,N_10520);
or U10892 (N_10892,N_10588,N_10611);
or U10893 (N_10893,N_10699,N_10605);
and U10894 (N_10894,N_10623,N_10562);
nor U10895 (N_10895,N_10599,N_10590);
and U10896 (N_10896,N_10553,N_10733);
or U10897 (N_10897,N_10632,N_10733);
nor U10898 (N_10898,N_10731,N_10684);
nand U10899 (N_10899,N_10551,N_10534);
or U10900 (N_10900,N_10743,N_10685);
and U10901 (N_10901,N_10519,N_10655);
and U10902 (N_10902,N_10576,N_10619);
or U10903 (N_10903,N_10698,N_10650);
and U10904 (N_10904,N_10679,N_10687);
nor U10905 (N_10905,N_10572,N_10722);
or U10906 (N_10906,N_10528,N_10541);
xnor U10907 (N_10907,N_10585,N_10576);
and U10908 (N_10908,N_10727,N_10649);
nand U10909 (N_10909,N_10539,N_10685);
nor U10910 (N_10910,N_10590,N_10720);
nand U10911 (N_10911,N_10713,N_10552);
or U10912 (N_10912,N_10563,N_10620);
or U10913 (N_10913,N_10691,N_10537);
nor U10914 (N_10914,N_10715,N_10621);
nand U10915 (N_10915,N_10636,N_10623);
nor U10916 (N_10916,N_10682,N_10510);
and U10917 (N_10917,N_10540,N_10643);
nor U10918 (N_10918,N_10575,N_10549);
xor U10919 (N_10919,N_10747,N_10573);
nor U10920 (N_10920,N_10748,N_10738);
nor U10921 (N_10921,N_10678,N_10521);
and U10922 (N_10922,N_10675,N_10706);
nor U10923 (N_10923,N_10514,N_10707);
nand U10924 (N_10924,N_10678,N_10688);
nand U10925 (N_10925,N_10534,N_10587);
or U10926 (N_10926,N_10739,N_10601);
nor U10927 (N_10927,N_10560,N_10562);
or U10928 (N_10928,N_10562,N_10558);
nor U10929 (N_10929,N_10504,N_10706);
or U10930 (N_10930,N_10617,N_10744);
or U10931 (N_10931,N_10595,N_10709);
or U10932 (N_10932,N_10517,N_10569);
and U10933 (N_10933,N_10598,N_10672);
and U10934 (N_10934,N_10593,N_10628);
and U10935 (N_10935,N_10700,N_10510);
nor U10936 (N_10936,N_10674,N_10626);
nor U10937 (N_10937,N_10645,N_10566);
nand U10938 (N_10938,N_10637,N_10570);
nand U10939 (N_10939,N_10529,N_10618);
nor U10940 (N_10940,N_10643,N_10714);
or U10941 (N_10941,N_10726,N_10641);
and U10942 (N_10942,N_10552,N_10508);
and U10943 (N_10943,N_10732,N_10657);
and U10944 (N_10944,N_10740,N_10528);
and U10945 (N_10945,N_10714,N_10617);
nor U10946 (N_10946,N_10706,N_10542);
nand U10947 (N_10947,N_10586,N_10698);
and U10948 (N_10948,N_10722,N_10620);
nor U10949 (N_10949,N_10564,N_10687);
nor U10950 (N_10950,N_10542,N_10631);
and U10951 (N_10951,N_10748,N_10587);
nor U10952 (N_10952,N_10667,N_10693);
or U10953 (N_10953,N_10545,N_10737);
nor U10954 (N_10954,N_10715,N_10694);
and U10955 (N_10955,N_10716,N_10672);
nand U10956 (N_10956,N_10740,N_10677);
and U10957 (N_10957,N_10553,N_10693);
nand U10958 (N_10958,N_10610,N_10671);
xor U10959 (N_10959,N_10715,N_10511);
xnor U10960 (N_10960,N_10724,N_10602);
xnor U10961 (N_10961,N_10576,N_10609);
nand U10962 (N_10962,N_10719,N_10602);
and U10963 (N_10963,N_10714,N_10649);
nor U10964 (N_10964,N_10659,N_10683);
and U10965 (N_10965,N_10623,N_10643);
or U10966 (N_10966,N_10609,N_10747);
nand U10967 (N_10967,N_10585,N_10537);
or U10968 (N_10968,N_10715,N_10641);
or U10969 (N_10969,N_10538,N_10638);
nand U10970 (N_10970,N_10639,N_10503);
nor U10971 (N_10971,N_10517,N_10556);
nand U10972 (N_10972,N_10738,N_10556);
or U10973 (N_10973,N_10716,N_10556);
nand U10974 (N_10974,N_10610,N_10639);
or U10975 (N_10975,N_10650,N_10714);
or U10976 (N_10976,N_10554,N_10593);
and U10977 (N_10977,N_10645,N_10740);
and U10978 (N_10978,N_10686,N_10569);
nand U10979 (N_10979,N_10696,N_10593);
and U10980 (N_10980,N_10594,N_10631);
and U10981 (N_10981,N_10610,N_10748);
and U10982 (N_10982,N_10671,N_10529);
or U10983 (N_10983,N_10555,N_10506);
and U10984 (N_10984,N_10531,N_10591);
and U10985 (N_10985,N_10526,N_10569);
or U10986 (N_10986,N_10597,N_10595);
or U10987 (N_10987,N_10741,N_10710);
or U10988 (N_10988,N_10577,N_10641);
nor U10989 (N_10989,N_10654,N_10537);
nand U10990 (N_10990,N_10740,N_10531);
and U10991 (N_10991,N_10711,N_10670);
and U10992 (N_10992,N_10579,N_10628);
nor U10993 (N_10993,N_10597,N_10592);
xor U10994 (N_10994,N_10532,N_10731);
nor U10995 (N_10995,N_10657,N_10658);
nor U10996 (N_10996,N_10715,N_10571);
xnor U10997 (N_10997,N_10653,N_10744);
nand U10998 (N_10998,N_10614,N_10613);
nand U10999 (N_10999,N_10571,N_10688);
or U11000 (N_11000,N_10839,N_10912);
nand U11001 (N_11001,N_10790,N_10872);
and U11002 (N_11002,N_10764,N_10988);
nand U11003 (N_11003,N_10935,N_10897);
or U11004 (N_11004,N_10880,N_10850);
and U11005 (N_11005,N_10983,N_10782);
nand U11006 (N_11006,N_10853,N_10902);
and U11007 (N_11007,N_10804,N_10758);
nand U11008 (N_11008,N_10791,N_10963);
and U11009 (N_11009,N_10836,N_10766);
or U11010 (N_11010,N_10827,N_10783);
xor U11011 (N_11011,N_10913,N_10869);
nor U11012 (N_11012,N_10970,N_10977);
xnor U11013 (N_11013,N_10920,N_10968);
and U11014 (N_11014,N_10937,N_10807);
nand U11015 (N_11015,N_10794,N_10773);
nor U11016 (N_11016,N_10991,N_10788);
and U11017 (N_11017,N_10754,N_10847);
and U11018 (N_11018,N_10763,N_10751);
and U11019 (N_11019,N_10928,N_10786);
and U11020 (N_11020,N_10762,N_10958);
and U11021 (N_11021,N_10967,N_10899);
nand U11022 (N_11022,N_10784,N_10965);
nand U11023 (N_11023,N_10802,N_10818);
or U11024 (N_11024,N_10882,N_10881);
nand U11025 (N_11025,N_10856,N_10940);
nand U11026 (N_11026,N_10816,N_10893);
or U11027 (N_11027,N_10757,N_10917);
nor U11028 (N_11028,N_10830,N_10931);
xnor U11029 (N_11029,N_10998,N_10960);
nand U11030 (N_11030,N_10950,N_10769);
or U11031 (N_11031,N_10870,N_10943);
and U11032 (N_11032,N_10889,N_10907);
and U11033 (N_11033,N_10819,N_10808);
nor U11034 (N_11034,N_10979,N_10844);
nor U11035 (N_11035,N_10756,N_10864);
and U11036 (N_11036,N_10813,N_10858);
nand U11037 (N_11037,N_10895,N_10948);
nand U11038 (N_11038,N_10852,N_10849);
or U11039 (N_11039,N_10959,N_10760);
and U11040 (N_11040,N_10837,N_10910);
nand U11041 (N_11041,N_10956,N_10780);
and U11042 (N_11042,N_10774,N_10999);
xnor U11043 (N_11043,N_10946,N_10831);
nand U11044 (N_11044,N_10927,N_10971);
or U11045 (N_11045,N_10771,N_10750);
nand U11046 (N_11046,N_10995,N_10814);
and U11047 (N_11047,N_10996,N_10855);
nor U11048 (N_11048,N_10835,N_10915);
or U11049 (N_11049,N_10871,N_10812);
nor U11050 (N_11050,N_10973,N_10755);
or U11051 (N_11051,N_10976,N_10953);
nor U11052 (N_11052,N_10823,N_10781);
or U11053 (N_11053,N_10944,N_10957);
nand U11054 (N_11054,N_10792,N_10890);
nand U11055 (N_11055,N_10862,N_10777);
or U11056 (N_11056,N_10874,N_10993);
xor U11057 (N_11057,N_10964,N_10972);
and U11058 (N_11058,N_10767,N_10992);
or U11059 (N_11059,N_10942,N_10824);
or U11060 (N_11060,N_10952,N_10798);
or U11061 (N_11061,N_10945,N_10975);
nor U11062 (N_11062,N_10908,N_10949);
and U11063 (N_11063,N_10987,N_10822);
nor U11064 (N_11064,N_10936,N_10803);
and U11065 (N_11065,N_10921,N_10994);
nor U11066 (N_11066,N_10860,N_10974);
or U11067 (N_11067,N_10896,N_10828);
and U11068 (N_11068,N_10955,N_10923);
and U11069 (N_11069,N_10875,N_10752);
xnor U11070 (N_11070,N_10787,N_10984);
and U11071 (N_11071,N_10857,N_10905);
and U11072 (N_11072,N_10768,N_10906);
nand U11073 (N_11073,N_10868,N_10879);
or U11074 (N_11074,N_10938,N_10775);
nand U11075 (N_11075,N_10990,N_10854);
nor U11076 (N_11076,N_10981,N_10900);
and U11077 (N_11077,N_10778,N_10918);
or U11078 (N_11078,N_10911,N_10851);
or U11079 (N_11079,N_10832,N_10817);
nand U11080 (N_11080,N_10922,N_10753);
and U11081 (N_11081,N_10772,N_10962);
nand U11082 (N_11082,N_10891,N_10840);
and U11083 (N_11083,N_10821,N_10888);
nor U11084 (N_11084,N_10863,N_10843);
and U11085 (N_11085,N_10825,N_10932);
nor U11086 (N_11086,N_10809,N_10901);
nor U11087 (N_11087,N_10826,N_10876);
or U11088 (N_11088,N_10796,N_10842);
and U11089 (N_11089,N_10966,N_10969);
nor U11090 (N_11090,N_10815,N_10834);
nor U11091 (N_11091,N_10980,N_10833);
xnor U11092 (N_11092,N_10789,N_10867);
nor U11093 (N_11093,N_10811,N_10894);
nand U11094 (N_11094,N_10898,N_10861);
and U11095 (N_11095,N_10846,N_10793);
nand U11096 (N_11096,N_10797,N_10785);
or U11097 (N_11097,N_10884,N_10904);
or U11098 (N_11098,N_10878,N_10865);
or U11099 (N_11099,N_10810,N_10914);
nor U11100 (N_11100,N_10885,N_10841);
xnor U11101 (N_11101,N_10845,N_10765);
or U11102 (N_11102,N_10829,N_10805);
or U11103 (N_11103,N_10978,N_10933);
xnor U11104 (N_11104,N_10887,N_10909);
and U11105 (N_11105,N_10925,N_10770);
xor U11106 (N_11106,N_10985,N_10941);
and U11107 (N_11107,N_10903,N_10954);
or U11108 (N_11108,N_10820,N_10848);
and U11109 (N_11109,N_10916,N_10926);
nand U11110 (N_11110,N_10838,N_10986);
or U11111 (N_11111,N_10930,N_10883);
nand U11112 (N_11112,N_10892,N_10859);
and U11113 (N_11113,N_10939,N_10886);
and U11114 (N_11114,N_10866,N_10795);
nand U11115 (N_11115,N_10806,N_10800);
nor U11116 (N_11116,N_10799,N_10779);
and U11117 (N_11117,N_10761,N_10934);
or U11118 (N_11118,N_10776,N_10997);
or U11119 (N_11119,N_10929,N_10801);
nand U11120 (N_11120,N_10947,N_10759);
and U11121 (N_11121,N_10989,N_10877);
nand U11122 (N_11122,N_10919,N_10961);
and U11123 (N_11123,N_10924,N_10873);
or U11124 (N_11124,N_10951,N_10982);
nor U11125 (N_11125,N_10812,N_10805);
nor U11126 (N_11126,N_10791,N_10985);
or U11127 (N_11127,N_10873,N_10800);
nor U11128 (N_11128,N_10758,N_10991);
nor U11129 (N_11129,N_10957,N_10782);
or U11130 (N_11130,N_10844,N_10769);
or U11131 (N_11131,N_10937,N_10788);
and U11132 (N_11132,N_10898,N_10860);
or U11133 (N_11133,N_10868,N_10776);
nand U11134 (N_11134,N_10938,N_10954);
or U11135 (N_11135,N_10960,N_10828);
or U11136 (N_11136,N_10865,N_10943);
nand U11137 (N_11137,N_10837,N_10862);
or U11138 (N_11138,N_10996,N_10784);
and U11139 (N_11139,N_10965,N_10859);
nand U11140 (N_11140,N_10913,N_10763);
xnor U11141 (N_11141,N_10954,N_10826);
and U11142 (N_11142,N_10796,N_10950);
or U11143 (N_11143,N_10753,N_10870);
and U11144 (N_11144,N_10902,N_10984);
nor U11145 (N_11145,N_10929,N_10834);
nand U11146 (N_11146,N_10846,N_10783);
and U11147 (N_11147,N_10974,N_10886);
nand U11148 (N_11148,N_10872,N_10831);
or U11149 (N_11149,N_10889,N_10830);
nand U11150 (N_11150,N_10759,N_10814);
or U11151 (N_11151,N_10905,N_10854);
and U11152 (N_11152,N_10874,N_10872);
nand U11153 (N_11153,N_10851,N_10861);
and U11154 (N_11154,N_10780,N_10764);
and U11155 (N_11155,N_10798,N_10962);
nor U11156 (N_11156,N_10796,N_10876);
and U11157 (N_11157,N_10766,N_10947);
nand U11158 (N_11158,N_10966,N_10827);
and U11159 (N_11159,N_10852,N_10761);
and U11160 (N_11160,N_10981,N_10796);
or U11161 (N_11161,N_10781,N_10916);
nand U11162 (N_11162,N_10993,N_10787);
nand U11163 (N_11163,N_10961,N_10999);
nand U11164 (N_11164,N_10943,N_10904);
xor U11165 (N_11165,N_10952,N_10866);
xor U11166 (N_11166,N_10978,N_10815);
xor U11167 (N_11167,N_10856,N_10774);
or U11168 (N_11168,N_10763,N_10966);
nand U11169 (N_11169,N_10829,N_10767);
or U11170 (N_11170,N_10812,N_10948);
xnor U11171 (N_11171,N_10993,N_10848);
nand U11172 (N_11172,N_10950,N_10810);
nand U11173 (N_11173,N_10779,N_10977);
nor U11174 (N_11174,N_10932,N_10770);
or U11175 (N_11175,N_10955,N_10837);
nand U11176 (N_11176,N_10998,N_10763);
nand U11177 (N_11177,N_10810,N_10768);
nor U11178 (N_11178,N_10795,N_10781);
or U11179 (N_11179,N_10883,N_10875);
nand U11180 (N_11180,N_10959,N_10810);
nand U11181 (N_11181,N_10805,N_10758);
xnor U11182 (N_11182,N_10970,N_10814);
and U11183 (N_11183,N_10800,N_10811);
and U11184 (N_11184,N_10827,N_10836);
or U11185 (N_11185,N_10788,N_10836);
nor U11186 (N_11186,N_10780,N_10773);
nor U11187 (N_11187,N_10768,N_10822);
xor U11188 (N_11188,N_10788,N_10964);
or U11189 (N_11189,N_10788,N_10848);
xnor U11190 (N_11190,N_10873,N_10811);
or U11191 (N_11191,N_10868,N_10951);
or U11192 (N_11192,N_10987,N_10855);
and U11193 (N_11193,N_10913,N_10942);
nor U11194 (N_11194,N_10971,N_10855);
and U11195 (N_11195,N_10917,N_10947);
and U11196 (N_11196,N_10855,N_10828);
xor U11197 (N_11197,N_10867,N_10821);
xnor U11198 (N_11198,N_10796,N_10921);
and U11199 (N_11199,N_10761,N_10877);
nand U11200 (N_11200,N_10757,N_10787);
or U11201 (N_11201,N_10772,N_10802);
or U11202 (N_11202,N_10943,N_10858);
and U11203 (N_11203,N_10883,N_10877);
and U11204 (N_11204,N_10753,N_10975);
nand U11205 (N_11205,N_10980,N_10917);
nand U11206 (N_11206,N_10898,N_10760);
and U11207 (N_11207,N_10922,N_10854);
or U11208 (N_11208,N_10754,N_10957);
or U11209 (N_11209,N_10962,N_10762);
or U11210 (N_11210,N_10909,N_10932);
or U11211 (N_11211,N_10916,N_10831);
nor U11212 (N_11212,N_10813,N_10846);
and U11213 (N_11213,N_10773,N_10953);
and U11214 (N_11214,N_10931,N_10777);
nor U11215 (N_11215,N_10947,N_10895);
nor U11216 (N_11216,N_10772,N_10883);
nor U11217 (N_11217,N_10794,N_10907);
nand U11218 (N_11218,N_10962,N_10912);
nand U11219 (N_11219,N_10846,N_10792);
and U11220 (N_11220,N_10756,N_10982);
nor U11221 (N_11221,N_10861,N_10842);
xor U11222 (N_11222,N_10853,N_10976);
and U11223 (N_11223,N_10923,N_10790);
or U11224 (N_11224,N_10845,N_10779);
and U11225 (N_11225,N_10956,N_10775);
xnor U11226 (N_11226,N_10946,N_10915);
nand U11227 (N_11227,N_10811,N_10864);
nor U11228 (N_11228,N_10790,N_10977);
and U11229 (N_11229,N_10950,N_10951);
nor U11230 (N_11230,N_10865,N_10832);
nand U11231 (N_11231,N_10755,N_10991);
or U11232 (N_11232,N_10991,N_10777);
nand U11233 (N_11233,N_10803,N_10775);
xor U11234 (N_11234,N_10782,N_10885);
and U11235 (N_11235,N_10845,N_10889);
or U11236 (N_11236,N_10953,N_10895);
nor U11237 (N_11237,N_10920,N_10946);
nor U11238 (N_11238,N_10814,N_10755);
or U11239 (N_11239,N_10944,N_10964);
xnor U11240 (N_11240,N_10855,N_10894);
nor U11241 (N_11241,N_10761,N_10996);
nor U11242 (N_11242,N_10882,N_10994);
nor U11243 (N_11243,N_10841,N_10834);
and U11244 (N_11244,N_10972,N_10865);
or U11245 (N_11245,N_10857,N_10981);
nor U11246 (N_11246,N_10817,N_10970);
xor U11247 (N_11247,N_10962,N_10989);
and U11248 (N_11248,N_10969,N_10814);
or U11249 (N_11249,N_10986,N_10990);
or U11250 (N_11250,N_11026,N_11084);
nor U11251 (N_11251,N_11219,N_11136);
or U11252 (N_11252,N_11059,N_11038);
nor U11253 (N_11253,N_11137,N_11129);
xnor U11254 (N_11254,N_11027,N_11139);
and U11255 (N_11255,N_11199,N_11039);
and U11256 (N_11256,N_11036,N_11020);
nor U11257 (N_11257,N_11009,N_11078);
nor U11258 (N_11258,N_11110,N_11130);
nand U11259 (N_11259,N_11135,N_11047);
or U11260 (N_11260,N_11091,N_11180);
nor U11261 (N_11261,N_11205,N_11032);
or U11262 (N_11262,N_11150,N_11143);
and U11263 (N_11263,N_11112,N_11007);
nor U11264 (N_11264,N_11092,N_11114);
or U11265 (N_11265,N_11173,N_11045);
or U11266 (N_11266,N_11127,N_11238);
nand U11267 (N_11267,N_11072,N_11156);
and U11268 (N_11268,N_11005,N_11062);
nor U11269 (N_11269,N_11030,N_11165);
nand U11270 (N_11270,N_11017,N_11120);
xor U11271 (N_11271,N_11145,N_11201);
nand U11272 (N_11272,N_11100,N_11119);
or U11273 (N_11273,N_11159,N_11087);
and U11274 (N_11274,N_11211,N_11177);
and U11275 (N_11275,N_11064,N_11086);
or U11276 (N_11276,N_11224,N_11198);
or U11277 (N_11277,N_11021,N_11158);
and U11278 (N_11278,N_11182,N_11171);
nor U11279 (N_11279,N_11022,N_11034);
and U11280 (N_11280,N_11105,N_11181);
or U11281 (N_11281,N_11157,N_11214);
xnor U11282 (N_11282,N_11098,N_11172);
nor U11283 (N_11283,N_11154,N_11204);
or U11284 (N_11284,N_11178,N_11018);
nand U11285 (N_11285,N_11108,N_11044);
and U11286 (N_11286,N_11203,N_11208);
or U11287 (N_11287,N_11174,N_11024);
and U11288 (N_11288,N_11207,N_11161);
nand U11289 (N_11289,N_11115,N_11230);
nand U11290 (N_11290,N_11011,N_11142);
and U11291 (N_11291,N_11057,N_11082);
nand U11292 (N_11292,N_11099,N_11243);
nand U11293 (N_11293,N_11240,N_11235);
or U11294 (N_11294,N_11215,N_11228);
and U11295 (N_11295,N_11233,N_11225);
and U11296 (N_11296,N_11094,N_11186);
xor U11297 (N_11297,N_11152,N_11242);
nand U11298 (N_11298,N_11000,N_11069);
nor U11299 (N_11299,N_11179,N_11241);
nor U11300 (N_11300,N_11080,N_11213);
and U11301 (N_11301,N_11122,N_11079);
nor U11302 (N_11302,N_11169,N_11132);
and U11303 (N_11303,N_11232,N_11209);
nand U11304 (N_11304,N_11226,N_11187);
and U11305 (N_11305,N_11128,N_11245);
nand U11306 (N_11306,N_11088,N_11192);
and U11307 (N_11307,N_11194,N_11055);
or U11308 (N_11308,N_11140,N_11176);
or U11309 (N_11309,N_11247,N_11067);
nor U11310 (N_11310,N_11151,N_11001);
and U11311 (N_11311,N_11166,N_11050);
nand U11312 (N_11312,N_11090,N_11109);
nor U11313 (N_11313,N_11093,N_11025);
nor U11314 (N_11314,N_11004,N_11246);
or U11315 (N_11315,N_11175,N_11075);
nor U11316 (N_11316,N_11141,N_11249);
xnor U11317 (N_11317,N_11239,N_11113);
and U11318 (N_11318,N_11037,N_11218);
and U11319 (N_11319,N_11031,N_11164);
or U11320 (N_11320,N_11125,N_11043);
nor U11321 (N_11321,N_11046,N_11190);
or U11322 (N_11322,N_11051,N_11148);
nor U11323 (N_11323,N_11081,N_11124);
xnor U11324 (N_11324,N_11196,N_11016);
nor U11325 (N_11325,N_11040,N_11210);
nor U11326 (N_11326,N_11063,N_11168);
or U11327 (N_11327,N_11162,N_11073);
nor U11328 (N_11328,N_11227,N_11008);
nor U11329 (N_11329,N_11131,N_11106);
nor U11330 (N_11330,N_11111,N_11134);
nor U11331 (N_11331,N_11085,N_11160);
nor U11332 (N_11332,N_11170,N_11006);
and U11333 (N_11333,N_11155,N_11014);
nand U11334 (N_11334,N_11096,N_11167);
or U11335 (N_11335,N_11195,N_11049);
and U11336 (N_11336,N_11023,N_11189);
nand U11337 (N_11337,N_11133,N_11185);
nand U11338 (N_11338,N_11248,N_11216);
nand U11339 (N_11339,N_11217,N_11102);
nand U11340 (N_11340,N_11074,N_11188);
or U11341 (N_11341,N_11191,N_11065);
nor U11342 (N_11342,N_11116,N_11071);
nand U11343 (N_11343,N_11138,N_11041);
and U11344 (N_11344,N_11048,N_11149);
or U11345 (N_11345,N_11070,N_11035);
nand U11346 (N_11346,N_11076,N_11222);
nand U11347 (N_11347,N_11095,N_11104);
nand U11348 (N_11348,N_11231,N_11234);
nor U11349 (N_11349,N_11123,N_11012);
or U11350 (N_11350,N_11058,N_11206);
nor U11351 (N_11351,N_11056,N_11042);
or U11352 (N_11352,N_11146,N_11101);
or U11353 (N_11353,N_11223,N_11053);
nor U11354 (N_11354,N_11244,N_11060);
xor U11355 (N_11355,N_11015,N_11197);
nand U11356 (N_11356,N_11118,N_11033);
and U11357 (N_11357,N_11153,N_11066);
nand U11358 (N_11358,N_11202,N_11212);
nor U11359 (N_11359,N_11103,N_11077);
or U11360 (N_11360,N_11221,N_11083);
nand U11361 (N_11361,N_11089,N_11193);
xnor U11362 (N_11362,N_11200,N_11010);
or U11363 (N_11363,N_11220,N_11126);
or U11364 (N_11364,N_11117,N_11147);
and U11365 (N_11365,N_11121,N_11184);
nor U11366 (N_11366,N_11003,N_11237);
nand U11367 (N_11367,N_11097,N_11236);
or U11368 (N_11368,N_11028,N_11163);
or U11369 (N_11369,N_11061,N_11068);
nand U11370 (N_11370,N_11019,N_11229);
and U11371 (N_11371,N_11052,N_11002);
nand U11372 (N_11372,N_11013,N_11183);
xor U11373 (N_11373,N_11054,N_11144);
nor U11374 (N_11374,N_11107,N_11029);
nand U11375 (N_11375,N_11141,N_11215);
nor U11376 (N_11376,N_11043,N_11123);
or U11377 (N_11377,N_11132,N_11014);
nor U11378 (N_11378,N_11138,N_11244);
and U11379 (N_11379,N_11187,N_11068);
or U11380 (N_11380,N_11168,N_11167);
nor U11381 (N_11381,N_11196,N_11136);
or U11382 (N_11382,N_11023,N_11064);
nor U11383 (N_11383,N_11003,N_11140);
xor U11384 (N_11384,N_11147,N_11148);
nand U11385 (N_11385,N_11248,N_11136);
nor U11386 (N_11386,N_11150,N_11211);
or U11387 (N_11387,N_11203,N_11099);
nand U11388 (N_11388,N_11009,N_11044);
nand U11389 (N_11389,N_11080,N_11130);
or U11390 (N_11390,N_11040,N_11076);
xnor U11391 (N_11391,N_11163,N_11102);
and U11392 (N_11392,N_11150,N_11137);
xnor U11393 (N_11393,N_11045,N_11054);
and U11394 (N_11394,N_11012,N_11109);
nor U11395 (N_11395,N_11069,N_11196);
nor U11396 (N_11396,N_11082,N_11016);
and U11397 (N_11397,N_11120,N_11138);
xor U11398 (N_11398,N_11222,N_11150);
nor U11399 (N_11399,N_11028,N_11214);
nor U11400 (N_11400,N_11110,N_11058);
and U11401 (N_11401,N_11032,N_11061);
nor U11402 (N_11402,N_11111,N_11064);
nor U11403 (N_11403,N_11004,N_11059);
xnor U11404 (N_11404,N_11091,N_11185);
or U11405 (N_11405,N_11001,N_11056);
and U11406 (N_11406,N_11213,N_11174);
and U11407 (N_11407,N_11087,N_11160);
nand U11408 (N_11408,N_11221,N_11166);
or U11409 (N_11409,N_11206,N_11055);
nand U11410 (N_11410,N_11181,N_11186);
or U11411 (N_11411,N_11106,N_11216);
and U11412 (N_11412,N_11016,N_11142);
and U11413 (N_11413,N_11064,N_11021);
or U11414 (N_11414,N_11192,N_11140);
nor U11415 (N_11415,N_11094,N_11213);
nand U11416 (N_11416,N_11046,N_11180);
nand U11417 (N_11417,N_11170,N_11054);
xor U11418 (N_11418,N_11125,N_11097);
nor U11419 (N_11419,N_11124,N_11216);
nand U11420 (N_11420,N_11131,N_11201);
nand U11421 (N_11421,N_11098,N_11216);
or U11422 (N_11422,N_11051,N_11147);
and U11423 (N_11423,N_11027,N_11086);
and U11424 (N_11424,N_11105,N_11162);
nor U11425 (N_11425,N_11026,N_11123);
and U11426 (N_11426,N_11233,N_11211);
nor U11427 (N_11427,N_11105,N_11094);
nor U11428 (N_11428,N_11130,N_11192);
and U11429 (N_11429,N_11239,N_11196);
and U11430 (N_11430,N_11222,N_11041);
and U11431 (N_11431,N_11170,N_11043);
or U11432 (N_11432,N_11044,N_11075);
nor U11433 (N_11433,N_11120,N_11199);
nor U11434 (N_11434,N_11054,N_11202);
and U11435 (N_11435,N_11127,N_11104);
nand U11436 (N_11436,N_11238,N_11111);
and U11437 (N_11437,N_11054,N_11225);
nand U11438 (N_11438,N_11133,N_11068);
nand U11439 (N_11439,N_11205,N_11023);
nand U11440 (N_11440,N_11075,N_11042);
nand U11441 (N_11441,N_11178,N_11082);
nand U11442 (N_11442,N_11058,N_11195);
nand U11443 (N_11443,N_11069,N_11063);
nand U11444 (N_11444,N_11175,N_11083);
and U11445 (N_11445,N_11053,N_11154);
nor U11446 (N_11446,N_11076,N_11135);
and U11447 (N_11447,N_11022,N_11016);
and U11448 (N_11448,N_11154,N_11219);
nor U11449 (N_11449,N_11191,N_11114);
nand U11450 (N_11450,N_11129,N_11078);
and U11451 (N_11451,N_11022,N_11070);
and U11452 (N_11452,N_11010,N_11063);
nor U11453 (N_11453,N_11139,N_11230);
and U11454 (N_11454,N_11040,N_11055);
nand U11455 (N_11455,N_11181,N_11037);
nor U11456 (N_11456,N_11087,N_11152);
nand U11457 (N_11457,N_11118,N_11207);
nand U11458 (N_11458,N_11087,N_11203);
xnor U11459 (N_11459,N_11152,N_11025);
nand U11460 (N_11460,N_11009,N_11133);
or U11461 (N_11461,N_11175,N_11137);
xnor U11462 (N_11462,N_11037,N_11232);
xor U11463 (N_11463,N_11109,N_11001);
nor U11464 (N_11464,N_11110,N_11069);
nand U11465 (N_11465,N_11181,N_11074);
nor U11466 (N_11466,N_11062,N_11059);
nand U11467 (N_11467,N_11034,N_11158);
and U11468 (N_11468,N_11167,N_11005);
nand U11469 (N_11469,N_11178,N_11179);
or U11470 (N_11470,N_11070,N_11072);
nand U11471 (N_11471,N_11248,N_11211);
and U11472 (N_11472,N_11233,N_11197);
or U11473 (N_11473,N_11046,N_11177);
nand U11474 (N_11474,N_11175,N_11208);
nand U11475 (N_11475,N_11121,N_11215);
and U11476 (N_11476,N_11224,N_11028);
xor U11477 (N_11477,N_11105,N_11165);
and U11478 (N_11478,N_11038,N_11101);
nand U11479 (N_11479,N_11009,N_11089);
nand U11480 (N_11480,N_11150,N_11165);
nand U11481 (N_11481,N_11132,N_11195);
nor U11482 (N_11482,N_11172,N_11168);
or U11483 (N_11483,N_11218,N_11042);
and U11484 (N_11484,N_11192,N_11000);
nand U11485 (N_11485,N_11121,N_11084);
xnor U11486 (N_11486,N_11024,N_11178);
nand U11487 (N_11487,N_11140,N_11119);
or U11488 (N_11488,N_11178,N_11020);
or U11489 (N_11489,N_11139,N_11189);
and U11490 (N_11490,N_11187,N_11179);
nor U11491 (N_11491,N_11085,N_11212);
xor U11492 (N_11492,N_11142,N_11125);
nor U11493 (N_11493,N_11072,N_11098);
nand U11494 (N_11494,N_11033,N_11237);
and U11495 (N_11495,N_11117,N_11129);
and U11496 (N_11496,N_11164,N_11009);
or U11497 (N_11497,N_11127,N_11109);
or U11498 (N_11498,N_11033,N_11096);
nor U11499 (N_11499,N_11174,N_11235);
xnor U11500 (N_11500,N_11373,N_11310);
or U11501 (N_11501,N_11366,N_11266);
nand U11502 (N_11502,N_11476,N_11311);
nor U11503 (N_11503,N_11370,N_11272);
or U11504 (N_11504,N_11323,N_11394);
nand U11505 (N_11505,N_11427,N_11363);
nand U11506 (N_11506,N_11338,N_11441);
nor U11507 (N_11507,N_11492,N_11488);
xor U11508 (N_11508,N_11491,N_11282);
and U11509 (N_11509,N_11430,N_11278);
and U11510 (N_11510,N_11493,N_11390);
or U11511 (N_11511,N_11456,N_11381);
xnor U11512 (N_11512,N_11479,N_11379);
and U11513 (N_11513,N_11314,N_11400);
nand U11514 (N_11514,N_11374,N_11485);
and U11515 (N_11515,N_11481,N_11432);
nand U11516 (N_11516,N_11267,N_11307);
or U11517 (N_11517,N_11384,N_11355);
and U11518 (N_11518,N_11471,N_11306);
nor U11519 (N_11519,N_11412,N_11302);
and U11520 (N_11520,N_11421,N_11459);
and U11521 (N_11521,N_11414,N_11262);
nand U11522 (N_11522,N_11297,N_11340);
and U11523 (N_11523,N_11419,N_11321);
nand U11524 (N_11524,N_11359,N_11475);
nand U11525 (N_11525,N_11404,N_11499);
nor U11526 (N_11526,N_11261,N_11496);
nand U11527 (N_11527,N_11478,N_11446);
and U11528 (N_11528,N_11251,N_11294);
nor U11529 (N_11529,N_11342,N_11292);
nand U11530 (N_11530,N_11354,N_11410);
nand U11531 (N_11531,N_11283,N_11448);
or U11532 (N_11532,N_11250,N_11439);
or U11533 (N_11533,N_11273,N_11423);
and U11534 (N_11534,N_11325,N_11411);
or U11535 (N_11535,N_11489,N_11328);
nand U11536 (N_11536,N_11413,N_11389);
and U11537 (N_11537,N_11405,N_11332);
and U11538 (N_11538,N_11437,N_11349);
and U11539 (N_11539,N_11472,N_11388);
nor U11540 (N_11540,N_11315,N_11377);
nor U11541 (N_11541,N_11433,N_11444);
and U11542 (N_11542,N_11452,N_11317);
or U11543 (N_11543,N_11322,N_11256);
nand U11544 (N_11544,N_11265,N_11420);
and U11545 (N_11545,N_11258,N_11320);
or U11546 (N_11546,N_11350,N_11290);
nor U11547 (N_11547,N_11270,N_11417);
nor U11548 (N_11548,N_11442,N_11276);
nor U11549 (N_11549,N_11333,N_11434);
nor U11550 (N_11550,N_11316,N_11449);
nor U11551 (N_11551,N_11299,N_11467);
nand U11552 (N_11552,N_11406,N_11369);
nor U11553 (N_11553,N_11331,N_11477);
nor U11554 (N_11554,N_11367,N_11398);
nand U11555 (N_11555,N_11457,N_11422);
or U11556 (N_11556,N_11329,N_11454);
and U11557 (N_11557,N_11431,N_11280);
and U11558 (N_11558,N_11259,N_11380);
nand U11559 (N_11559,N_11498,N_11296);
nor U11560 (N_11560,N_11382,N_11426);
nand U11561 (N_11561,N_11344,N_11252);
and U11562 (N_11562,N_11348,N_11371);
or U11563 (N_11563,N_11424,N_11330);
nor U11564 (N_11564,N_11480,N_11428);
or U11565 (N_11565,N_11490,N_11495);
nor U11566 (N_11566,N_11401,N_11466);
nor U11567 (N_11567,N_11260,N_11318);
and U11568 (N_11568,N_11438,N_11284);
nor U11569 (N_11569,N_11253,N_11462);
nor U11570 (N_11570,N_11387,N_11347);
or U11571 (N_11571,N_11268,N_11396);
xor U11572 (N_11572,N_11376,N_11418);
xor U11573 (N_11573,N_11312,N_11407);
or U11574 (N_11574,N_11291,N_11360);
nor U11575 (N_11575,N_11416,N_11443);
nor U11576 (N_11576,N_11327,N_11300);
nor U11577 (N_11577,N_11425,N_11460);
and U11578 (N_11578,N_11453,N_11337);
xnor U11579 (N_11579,N_11346,N_11295);
nor U11580 (N_11580,N_11339,N_11361);
or U11581 (N_11581,N_11458,N_11378);
nand U11582 (N_11582,N_11450,N_11386);
nand U11583 (N_11583,N_11469,N_11362);
or U11584 (N_11584,N_11397,N_11372);
or U11585 (N_11585,N_11356,N_11409);
nor U11586 (N_11586,N_11274,N_11319);
or U11587 (N_11587,N_11463,N_11264);
nand U11588 (N_11588,N_11343,N_11383);
nand U11589 (N_11589,N_11461,N_11468);
or U11590 (N_11590,N_11275,N_11473);
nor U11591 (N_11591,N_11365,N_11385);
nor U11592 (N_11592,N_11482,N_11336);
xor U11593 (N_11593,N_11352,N_11326);
or U11594 (N_11594,N_11357,N_11341);
or U11595 (N_11595,N_11313,N_11415);
nand U11596 (N_11596,N_11353,N_11486);
nand U11597 (N_11597,N_11470,N_11303);
nand U11598 (N_11598,N_11308,N_11403);
xnor U11599 (N_11599,N_11257,N_11334);
nand U11600 (N_11600,N_11484,N_11435);
nand U11601 (N_11601,N_11408,N_11402);
nor U11602 (N_11602,N_11345,N_11436);
nand U11603 (N_11603,N_11474,N_11293);
nand U11604 (N_11604,N_11455,N_11288);
or U11605 (N_11605,N_11375,N_11497);
and U11606 (N_11606,N_11464,N_11301);
nand U11607 (N_11607,N_11465,N_11395);
nor U11608 (N_11608,N_11255,N_11287);
and U11609 (N_11609,N_11309,N_11263);
or U11610 (N_11610,N_11451,N_11391);
or U11611 (N_11611,N_11286,N_11279);
nand U11612 (N_11612,N_11393,N_11392);
and U11613 (N_11613,N_11277,N_11445);
nand U11614 (N_11614,N_11298,N_11304);
or U11615 (N_11615,N_11305,N_11483);
nor U11616 (N_11616,N_11358,N_11281);
nor U11617 (N_11617,N_11324,N_11254);
or U11618 (N_11618,N_11429,N_11368);
and U11619 (N_11619,N_11487,N_11364);
nand U11620 (N_11620,N_11447,N_11494);
nor U11621 (N_11621,N_11440,N_11335);
nor U11622 (N_11622,N_11399,N_11351);
nor U11623 (N_11623,N_11271,N_11289);
or U11624 (N_11624,N_11269,N_11285);
and U11625 (N_11625,N_11422,N_11404);
or U11626 (N_11626,N_11445,N_11418);
nand U11627 (N_11627,N_11474,N_11435);
and U11628 (N_11628,N_11315,N_11338);
nand U11629 (N_11629,N_11348,N_11369);
and U11630 (N_11630,N_11315,N_11402);
or U11631 (N_11631,N_11350,N_11259);
or U11632 (N_11632,N_11306,N_11255);
nor U11633 (N_11633,N_11316,N_11348);
nor U11634 (N_11634,N_11446,N_11403);
and U11635 (N_11635,N_11499,N_11303);
nor U11636 (N_11636,N_11364,N_11414);
and U11637 (N_11637,N_11252,N_11452);
or U11638 (N_11638,N_11277,N_11297);
xor U11639 (N_11639,N_11286,N_11394);
xor U11640 (N_11640,N_11337,N_11422);
and U11641 (N_11641,N_11490,N_11451);
and U11642 (N_11642,N_11486,N_11377);
and U11643 (N_11643,N_11404,N_11300);
or U11644 (N_11644,N_11477,N_11378);
and U11645 (N_11645,N_11464,N_11288);
nand U11646 (N_11646,N_11272,N_11276);
nand U11647 (N_11647,N_11264,N_11380);
xor U11648 (N_11648,N_11406,N_11298);
or U11649 (N_11649,N_11410,N_11347);
and U11650 (N_11650,N_11341,N_11436);
or U11651 (N_11651,N_11398,N_11340);
and U11652 (N_11652,N_11297,N_11257);
xor U11653 (N_11653,N_11428,N_11364);
or U11654 (N_11654,N_11393,N_11469);
nor U11655 (N_11655,N_11357,N_11466);
and U11656 (N_11656,N_11454,N_11429);
and U11657 (N_11657,N_11488,N_11359);
nand U11658 (N_11658,N_11354,N_11342);
nor U11659 (N_11659,N_11404,N_11258);
nor U11660 (N_11660,N_11346,N_11364);
or U11661 (N_11661,N_11497,N_11400);
or U11662 (N_11662,N_11301,N_11362);
nor U11663 (N_11663,N_11393,N_11418);
or U11664 (N_11664,N_11452,N_11483);
nand U11665 (N_11665,N_11387,N_11408);
nand U11666 (N_11666,N_11266,N_11283);
or U11667 (N_11667,N_11410,N_11257);
nand U11668 (N_11668,N_11440,N_11340);
nor U11669 (N_11669,N_11456,N_11383);
nand U11670 (N_11670,N_11401,N_11473);
nor U11671 (N_11671,N_11373,N_11402);
or U11672 (N_11672,N_11479,N_11427);
nand U11673 (N_11673,N_11312,N_11385);
nand U11674 (N_11674,N_11318,N_11272);
nand U11675 (N_11675,N_11351,N_11269);
nand U11676 (N_11676,N_11316,N_11447);
or U11677 (N_11677,N_11360,N_11283);
xnor U11678 (N_11678,N_11371,N_11256);
nor U11679 (N_11679,N_11311,N_11384);
xnor U11680 (N_11680,N_11299,N_11263);
and U11681 (N_11681,N_11268,N_11292);
nand U11682 (N_11682,N_11407,N_11479);
or U11683 (N_11683,N_11349,N_11294);
nor U11684 (N_11684,N_11430,N_11491);
xor U11685 (N_11685,N_11252,N_11336);
nor U11686 (N_11686,N_11276,N_11465);
or U11687 (N_11687,N_11333,N_11287);
nor U11688 (N_11688,N_11454,N_11286);
nand U11689 (N_11689,N_11252,N_11403);
xnor U11690 (N_11690,N_11418,N_11320);
and U11691 (N_11691,N_11355,N_11357);
nor U11692 (N_11692,N_11481,N_11448);
nor U11693 (N_11693,N_11273,N_11430);
nand U11694 (N_11694,N_11434,N_11294);
nand U11695 (N_11695,N_11398,N_11470);
xnor U11696 (N_11696,N_11274,N_11276);
and U11697 (N_11697,N_11384,N_11363);
xnor U11698 (N_11698,N_11278,N_11493);
nand U11699 (N_11699,N_11253,N_11448);
nor U11700 (N_11700,N_11305,N_11371);
nand U11701 (N_11701,N_11431,N_11385);
nor U11702 (N_11702,N_11396,N_11434);
and U11703 (N_11703,N_11447,N_11275);
and U11704 (N_11704,N_11351,N_11296);
or U11705 (N_11705,N_11364,N_11475);
or U11706 (N_11706,N_11258,N_11491);
and U11707 (N_11707,N_11441,N_11339);
nand U11708 (N_11708,N_11443,N_11287);
nand U11709 (N_11709,N_11401,N_11316);
nor U11710 (N_11710,N_11437,N_11361);
xnor U11711 (N_11711,N_11279,N_11465);
or U11712 (N_11712,N_11494,N_11437);
nor U11713 (N_11713,N_11485,N_11353);
nand U11714 (N_11714,N_11494,N_11362);
nand U11715 (N_11715,N_11382,N_11307);
or U11716 (N_11716,N_11359,N_11459);
and U11717 (N_11717,N_11463,N_11296);
or U11718 (N_11718,N_11479,N_11311);
nor U11719 (N_11719,N_11487,N_11363);
and U11720 (N_11720,N_11446,N_11439);
and U11721 (N_11721,N_11348,N_11332);
and U11722 (N_11722,N_11325,N_11382);
and U11723 (N_11723,N_11284,N_11361);
nor U11724 (N_11724,N_11258,N_11310);
and U11725 (N_11725,N_11406,N_11478);
or U11726 (N_11726,N_11497,N_11402);
nand U11727 (N_11727,N_11394,N_11345);
or U11728 (N_11728,N_11442,N_11287);
and U11729 (N_11729,N_11308,N_11322);
and U11730 (N_11730,N_11298,N_11336);
and U11731 (N_11731,N_11423,N_11446);
and U11732 (N_11732,N_11484,N_11268);
or U11733 (N_11733,N_11305,N_11313);
and U11734 (N_11734,N_11475,N_11422);
or U11735 (N_11735,N_11464,N_11498);
nand U11736 (N_11736,N_11377,N_11303);
or U11737 (N_11737,N_11294,N_11478);
or U11738 (N_11738,N_11331,N_11499);
and U11739 (N_11739,N_11276,N_11351);
xor U11740 (N_11740,N_11477,N_11309);
xor U11741 (N_11741,N_11412,N_11330);
or U11742 (N_11742,N_11354,N_11315);
and U11743 (N_11743,N_11302,N_11320);
and U11744 (N_11744,N_11377,N_11439);
nor U11745 (N_11745,N_11398,N_11492);
nor U11746 (N_11746,N_11459,N_11381);
nor U11747 (N_11747,N_11418,N_11454);
nor U11748 (N_11748,N_11345,N_11276);
or U11749 (N_11749,N_11293,N_11304);
and U11750 (N_11750,N_11664,N_11577);
and U11751 (N_11751,N_11536,N_11705);
nor U11752 (N_11752,N_11623,N_11678);
nor U11753 (N_11753,N_11691,N_11519);
nor U11754 (N_11754,N_11745,N_11548);
and U11755 (N_11755,N_11600,N_11570);
or U11756 (N_11756,N_11598,N_11684);
or U11757 (N_11757,N_11746,N_11500);
or U11758 (N_11758,N_11749,N_11516);
nand U11759 (N_11759,N_11680,N_11734);
nor U11760 (N_11760,N_11586,N_11532);
nand U11761 (N_11761,N_11510,N_11544);
and U11762 (N_11762,N_11742,N_11579);
or U11763 (N_11763,N_11662,N_11638);
or U11764 (N_11764,N_11744,N_11661);
and U11765 (N_11765,N_11730,N_11550);
and U11766 (N_11766,N_11640,N_11655);
nor U11767 (N_11767,N_11563,N_11694);
or U11768 (N_11768,N_11549,N_11551);
nor U11769 (N_11769,N_11525,N_11528);
xnor U11770 (N_11770,N_11634,N_11722);
nand U11771 (N_11771,N_11572,N_11505);
or U11772 (N_11772,N_11587,N_11567);
or U11773 (N_11773,N_11670,N_11689);
nor U11774 (N_11774,N_11732,N_11725);
nand U11775 (N_11775,N_11679,N_11574);
and U11776 (N_11776,N_11639,N_11612);
nand U11777 (N_11777,N_11568,N_11696);
or U11778 (N_11778,N_11513,N_11697);
or U11779 (N_11779,N_11533,N_11613);
nor U11780 (N_11780,N_11594,N_11537);
nor U11781 (N_11781,N_11521,N_11520);
or U11782 (N_11782,N_11699,N_11658);
nand U11783 (N_11783,N_11713,N_11740);
nand U11784 (N_11784,N_11667,N_11704);
nor U11785 (N_11785,N_11663,N_11523);
and U11786 (N_11786,N_11605,N_11685);
xor U11787 (N_11787,N_11714,N_11649);
nand U11788 (N_11788,N_11580,N_11674);
and U11789 (N_11789,N_11614,N_11712);
nor U11790 (N_11790,N_11524,N_11522);
nand U11791 (N_11791,N_11619,N_11592);
nor U11792 (N_11792,N_11671,N_11615);
nor U11793 (N_11793,N_11683,N_11687);
nor U11794 (N_11794,N_11602,N_11535);
or U11795 (N_11795,N_11653,N_11622);
and U11796 (N_11796,N_11660,N_11541);
nand U11797 (N_11797,N_11644,N_11737);
or U11798 (N_11798,N_11741,N_11628);
and U11799 (N_11799,N_11665,N_11647);
or U11800 (N_11800,N_11569,N_11502);
or U11801 (N_11801,N_11603,N_11616);
nor U11802 (N_11802,N_11727,N_11554);
and U11803 (N_11803,N_11641,N_11573);
and U11804 (N_11804,N_11666,N_11534);
or U11805 (N_11805,N_11627,N_11546);
or U11806 (N_11806,N_11717,N_11538);
and U11807 (N_11807,N_11632,N_11575);
and U11808 (N_11808,N_11723,N_11631);
or U11809 (N_11809,N_11669,N_11625);
nand U11810 (N_11810,N_11511,N_11552);
xor U11811 (N_11811,N_11564,N_11698);
nor U11812 (N_11812,N_11743,N_11581);
and U11813 (N_11813,N_11630,N_11606);
and U11814 (N_11814,N_11709,N_11618);
nand U11815 (N_11815,N_11748,N_11692);
or U11816 (N_11816,N_11620,N_11635);
nor U11817 (N_11817,N_11518,N_11643);
or U11818 (N_11818,N_11553,N_11590);
nor U11819 (N_11819,N_11738,N_11576);
nor U11820 (N_11820,N_11585,N_11729);
nand U11821 (N_11821,N_11584,N_11539);
or U11822 (N_11822,N_11506,N_11545);
and U11823 (N_11823,N_11675,N_11503);
nand U11824 (N_11824,N_11621,N_11591);
or U11825 (N_11825,N_11626,N_11595);
nand U11826 (N_11826,N_11645,N_11693);
and U11827 (N_11827,N_11646,N_11700);
and U11828 (N_11828,N_11558,N_11681);
or U11829 (N_11829,N_11596,N_11716);
or U11830 (N_11830,N_11512,N_11711);
and U11831 (N_11831,N_11526,N_11710);
nor U11832 (N_11832,N_11637,N_11707);
xor U11833 (N_11833,N_11610,N_11629);
and U11834 (N_11834,N_11560,N_11571);
nand U11835 (N_11835,N_11686,N_11677);
nor U11836 (N_11836,N_11715,N_11611);
xor U11837 (N_11837,N_11731,N_11648);
nand U11838 (N_11838,N_11657,N_11682);
xor U11839 (N_11839,N_11515,N_11739);
and U11840 (N_11840,N_11589,N_11708);
nand U11841 (N_11841,N_11650,N_11726);
or U11842 (N_11842,N_11668,N_11633);
xor U11843 (N_11843,N_11597,N_11651);
nand U11844 (N_11844,N_11509,N_11703);
or U11845 (N_11845,N_11608,N_11556);
nand U11846 (N_11846,N_11593,N_11652);
nor U11847 (N_11847,N_11642,N_11721);
nor U11848 (N_11848,N_11540,N_11688);
and U11849 (N_11849,N_11702,N_11604);
and U11850 (N_11850,N_11517,N_11501);
or U11851 (N_11851,N_11659,N_11529);
and U11852 (N_11852,N_11547,N_11559);
nand U11853 (N_11853,N_11531,N_11530);
xnor U11854 (N_11854,N_11557,N_11527);
nand U11855 (N_11855,N_11701,N_11656);
or U11856 (N_11856,N_11543,N_11565);
or U11857 (N_11857,N_11673,N_11583);
nand U11858 (N_11858,N_11695,N_11507);
nand U11859 (N_11859,N_11607,N_11508);
nor U11860 (N_11860,N_11720,N_11578);
nor U11861 (N_11861,N_11718,N_11636);
and U11862 (N_11862,N_11566,N_11676);
or U11863 (N_11863,N_11672,N_11617);
or U11864 (N_11864,N_11735,N_11733);
nand U11865 (N_11865,N_11588,N_11724);
nor U11866 (N_11866,N_11706,N_11555);
and U11867 (N_11867,N_11582,N_11601);
and U11868 (N_11868,N_11514,N_11747);
nor U11869 (N_11869,N_11561,N_11562);
nand U11870 (N_11870,N_11690,N_11654);
nor U11871 (N_11871,N_11504,N_11736);
or U11872 (N_11872,N_11728,N_11609);
or U11873 (N_11873,N_11599,N_11624);
and U11874 (N_11874,N_11542,N_11719);
nor U11875 (N_11875,N_11560,N_11649);
or U11876 (N_11876,N_11505,N_11720);
and U11877 (N_11877,N_11574,N_11601);
nand U11878 (N_11878,N_11595,N_11685);
nor U11879 (N_11879,N_11624,N_11697);
nand U11880 (N_11880,N_11660,N_11672);
nand U11881 (N_11881,N_11640,N_11691);
nand U11882 (N_11882,N_11626,N_11732);
nand U11883 (N_11883,N_11533,N_11532);
and U11884 (N_11884,N_11682,N_11603);
nand U11885 (N_11885,N_11669,N_11667);
and U11886 (N_11886,N_11614,N_11618);
or U11887 (N_11887,N_11738,N_11714);
nor U11888 (N_11888,N_11567,N_11542);
nand U11889 (N_11889,N_11688,N_11572);
and U11890 (N_11890,N_11523,N_11664);
nand U11891 (N_11891,N_11660,N_11724);
nor U11892 (N_11892,N_11633,N_11661);
and U11893 (N_11893,N_11694,N_11635);
nor U11894 (N_11894,N_11504,N_11617);
nor U11895 (N_11895,N_11556,N_11679);
and U11896 (N_11896,N_11570,N_11723);
or U11897 (N_11897,N_11583,N_11666);
and U11898 (N_11898,N_11637,N_11681);
or U11899 (N_11899,N_11535,N_11618);
or U11900 (N_11900,N_11570,N_11544);
nand U11901 (N_11901,N_11622,N_11561);
or U11902 (N_11902,N_11502,N_11721);
nand U11903 (N_11903,N_11708,N_11649);
nor U11904 (N_11904,N_11539,N_11603);
nor U11905 (N_11905,N_11525,N_11531);
and U11906 (N_11906,N_11667,N_11738);
nand U11907 (N_11907,N_11528,N_11672);
nand U11908 (N_11908,N_11560,N_11536);
nor U11909 (N_11909,N_11648,N_11558);
xor U11910 (N_11910,N_11540,N_11651);
nor U11911 (N_11911,N_11707,N_11590);
nor U11912 (N_11912,N_11595,N_11668);
or U11913 (N_11913,N_11504,N_11505);
and U11914 (N_11914,N_11551,N_11524);
nand U11915 (N_11915,N_11569,N_11626);
xnor U11916 (N_11916,N_11554,N_11522);
nor U11917 (N_11917,N_11506,N_11560);
nand U11918 (N_11918,N_11640,N_11707);
nor U11919 (N_11919,N_11618,N_11666);
nand U11920 (N_11920,N_11528,N_11712);
or U11921 (N_11921,N_11572,N_11730);
and U11922 (N_11922,N_11633,N_11653);
nor U11923 (N_11923,N_11636,N_11601);
or U11924 (N_11924,N_11705,N_11636);
nor U11925 (N_11925,N_11717,N_11566);
xor U11926 (N_11926,N_11579,N_11563);
xor U11927 (N_11927,N_11582,N_11600);
nand U11928 (N_11928,N_11655,N_11708);
nand U11929 (N_11929,N_11543,N_11582);
nor U11930 (N_11930,N_11511,N_11689);
or U11931 (N_11931,N_11617,N_11510);
nand U11932 (N_11932,N_11703,N_11579);
nand U11933 (N_11933,N_11524,N_11521);
or U11934 (N_11934,N_11561,N_11505);
nand U11935 (N_11935,N_11535,N_11605);
nand U11936 (N_11936,N_11621,N_11647);
nand U11937 (N_11937,N_11651,N_11745);
and U11938 (N_11938,N_11582,N_11679);
or U11939 (N_11939,N_11540,N_11666);
or U11940 (N_11940,N_11541,N_11589);
nand U11941 (N_11941,N_11741,N_11633);
or U11942 (N_11942,N_11610,N_11518);
nand U11943 (N_11943,N_11652,N_11745);
nor U11944 (N_11944,N_11621,N_11691);
nand U11945 (N_11945,N_11528,N_11513);
nor U11946 (N_11946,N_11687,N_11681);
and U11947 (N_11947,N_11590,N_11721);
or U11948 (N_11948,N_11522,N_11697);
and U11949 (N_11949,N_11581,N_11631);
nor U11950 (N_11950,N_11657,N_11738);
or U11951 (N_11951,N_11637,N_11702);
nor U11952 (N_11952,N_11544,N_11645);
or U11953 (N_11953,N_11661,N_11700);
and U11954 (N_11954,N_11586,N_11548);
and U11955 (N_11955,N_11622,N_11525);
nand U11956 (N_11956,N_11720,N_11679);
and U11957 (N_11957,N_11620,N_11599);
nor U11958 (N_11958,N_11725,N_11599);
nor U11959 (N_11959,N_11605,N_11516);
xnor U11960 (N_11960,N_11721,N_11696);
nand U11961 (N_11961,N_11633,N_11609);
nor U11962 (N_11962,N_11733,N_11532);
or U11963 (N_11963,N_11713,N_11586);
and U11964 (N_11964,N_11644,N_11589);
and U11965 (N_11965,N_11656,N_11717);
or U11966 (N_11966,N_11671,N_11518);
xor U11967 (N_11967,N_11672,N_11709);
nor U11968 (N_11968,N_11511,N_11576);
nand U11969 (N_11969,N_11542,N_11679);
nor U11970 (N_11970,N_11540,N_11582);
or U11971 (N_11971,N_11660,N_11641);
nor U11972 (N_11972,N_11557,N_11605);
or U11973 (N_11973,N_11598,N_11555);
and U11974 (N_11974,N_11527,N_11596);
and U11975 (N_11975,N_11610,N_11600);
nor U11976 (N_11976,N_11535,N_11546);
nand U11977 (N_11977,N_11727,N_11620);
nor U11978 (N_11978,N_11740,N_11651);
nand U11979 (N_11979,N_11689,N_11608);
nor U11980 (N_11980,N_11656,N_11713);
nand U11981 (N_11981,N_11590,N_11725);
nor U11982 (N_11982,N_11524,N_11704);
or U11983 (N_11983,N_11558,N_11701);
or U11984 (N_11984,N_11675,N_11616);
nand U11985 (N_11985,N_11654,N_11598);
or U11986 (N_11986,N_11694,N_11538);
or U11987 (N_11987,N_11714,N_11700);
nor U11988 (N_11988,N_11698,N_11638);
and U11989 (N_11989,N_11700,N_11711);
nor U11990 (N_11990,N_11646,N_11540);
nand U11991 (N_11991,N_11514,N_11681);
and U11992 (N_11992,N_11684,N_11690);
nor U11993 (N_11993,N_11722,N_11628);
and U11994 (N_11994,N_11621,N_11728);
or U11995 (N_11995,N_11651,N_11708);
xor U11996 (N_11996,N_11632,N_11732);
or U11997 (N_11997,N_11601,N_11650);
or U11998 (N_11998,N_11500,N_11658);
nor U11999 (N_11999,N_11546,N_11688);
nand U12000 (N_12000,N_11798,N_11958);
and U12001 (N_12001,N_11860,N_11903);
or U12002 (N_12002,N_11941,N_11771);
nor U12003 (N_12003,N_11775,N_11761);
and U12004 (N_12004,N_11897,N_11780);
nand U12005 (N_12005,N_11964,N_11874);
nand U12006 (N_12006,N_11859,N_11823);
or U12007 (N_12007,N_11993,N_11949);
or U12008 (N_12008,N_11869,N_11953);
nor U12009 (N_12009,N_11801,N_11822);
and U12010 (N_12010,N_11977,N_11789);
xor U12011 (N_12011,N_11765,N_11882);
nand U12012 (N_12012,N_11804,N_11991);
and U12013 (N_12013,N_11936,N_11965);
nand U12014 (N_12014,N_11792,N_11939);
and U12015 (N_12015,N_11986,N_11898);
nand U12016 (N_12016,N_11797,N_11750);
nand U12017 (N_12017,N_11870,N_11945);
nand U12018 (N_12018,N_11995,N_11967);
nand U12019 (N_12019,N_11819,N_11842);
nor U12020 (N_12020,N_11934,N_11907);
and U12021 (N_12021,N_11767,N_11794);
or U12022 (N_12022,N_11937,N_11932);
and U12023 (N_12023,N_11800,N_11880);
and U12024 (N_12024,N_11807,N_11774);
and U12025 (N_12025,N_11994,N_11997);
or U12026 (N_12026,N_11865,N_11835);
or U12027 (N_12027,N_11996,N_11830);
nand U12028 (N_12028,N_11918,N_11754);
nand U12029 (N_12029,N_11920,N_11884);
nand U12030 (N_12030,N_11809,N_11979);
nand U12031 (N_12031,N_11879,N_11838);
and U12032 (N_12032,N_11887,N_11817);
or U12033 (N_12033,N_11843,N_11970);
or U12034 (N_12034,N_11966,N_11814);
or U12035 (N_12035,N_11832,N_11772);
nand U12036 (N_12036,N_11781,N_11873);
nand U12037 (N_12037,N_11975,N_11872);
xnor U12038 (N_12038,N_11763,N_11971);
nand U12039 (N_12039,N_11866,N_11960);
nor U12040 (N_12040,N_11899,N_11854);
nor U12041 (N_12041,N_11755,N_11885);
nor U12042 (N_12042,N_11776,N_11974);
nor U12043 (N_12043,N_11824,N_11955);
and U12044 (N_12044,N_11791,N_11943);
and U12045 (N_12045,N_11779,N_11930);
or U12046 (N_12046,N_11891,N_11923);
nor U12047 (N_12047,N_11987,N_11957);
and U12048 (N_12048,N_11810,N_11983);
and U12049 (N_12049,N_11850,N_11803);
nor U12050 (N_12050,N_11788,N_11961);
and U12051 (N_12051,N_11826,N_11881);
or U12052 (N_12052,N_11856,N_11922);
nand U12053 (N_12053,N_11827,N_11844);
or U12054 (N_12054,N_11831,N_11852);
xnor U12055 (N_12055,N_11906,N_11752);
nor U12056 (N_12056,N_11841,N_11851);
nand U12057 (N_12057,N_11821,N_11892);
and U12058 (N_12058,N_11799,N_11768);
nand U12059 (N_12059,N_11905,N_11806);
or U12060 (N_12060,N_11929,N_11786);
xor U12061 (N_12061,N_11998,N_11858);
nand U12062 (N_12062,N_11783,N_11895);
xnor U12063 (N_12063,N_11904,N_11762);
xor U12064 (N_12064,N_11982,N_11833);
and U12065 (N_12065,N_11886,N_11769);
nand U12066 (N_12066,N_11978,N_11909);
nand U12067 (N_12067,N_11883,N_11942);
nor U12068 (N_12068,N_11840,N_11926);
xor U12069 (N_12069,N_11976,N_11901);
and U12070 (N_12070,N_11861,N_11900);
nand U12071 (N_12071,N_11816,N_11751);
nand U12072 (N_12072,N_11921,N_11848);
nor U12073 (N_12073,N_11876,N_11847);
nand U12074 (N_12074,N_11888,N_11924);
nor U12075 (N_12075,N_11917,N_11893);
xnor U12076 (N_12076,N_11862,N_11950);
nor U12077 (N_12077,N_11868,N_11948);
xor U12078 (N_12078,N_11871,N_11959);
nor U12079 (N_12079,N_11829,N_11855);
nor U12080 (N_12080,N_11952,N_11787);
and U12081 (N_12081,N_11812,N_11928);
nand U12082 (N_12082,N_11825,N_11815);
and U12083 (N_12083,N_11912,N_11805);
xor U12084 (N_12084,N_11980,N_11875);
xor U12085 (N_12085,N_11818,N_11947);
or U12086 (N_12086,N_11839,N_11968);
or U12087 (N_12087,N_11889,N_11784);
or U12088 (N_12088,N_11972,N_11944);
or U12089 (N_12089,N_11896,N_11785);
nor U12090 (N_12090,N_11914,N_11846);
nand U12091 (N_12091,N_11890,N_11931);
nand U12092 (N_12092,N_11770,N_11756);
xnor U12093 (N_12093,N_11894,N_11778);
nor U12094 (N_12094,N_11782,N_11940);
and U12095 (N_12095,N_11954,N_11802);
xnor U12096 (N_12096,N_11933,N_11867);
nand U12097 (N_12097,N_11915,N_11911);
or U12098 (N_12098,N_11793,N_11969);
xor U12099 (N_12099,N_11913,N_11935);
nor U12100 (N_12100,N_11956,N_11984);
nand U12101 (N_12101,N_11938,N_11760);
or U12102 (N_12102,N_11795,N_11981);
nor U12103 (N_12103,N_11853,N_11864);
nor U12104 (N_12104,N_11857,N_11820);
or U12105 (N_12105,N_11808,N_11919);
xor U12106 (N_12106,N_11849,N_11992);
and U12107 (N_12107,N_11796,N_11837);
or U12108 (N_12108,N_11925,N_11863);
xor U12109 (N_12109,N_11927,N_11828);
or U12110 (N_12110,N_11946,N_11764);
xor U12111 (N_12111,N_11902,N_11962);
nor U12112 (N_12112,N_11790,N_11999);
xnor U12113 (N_12113,N_11951,N_11878);
nor U12114 (N_12114,N_11766,N_11989);
nand U12115 (N_12115,N_11845,N_11773);
nand U12116 (N_12116,N_11777,N_11811);
or U12117 (N_12117,N_11910,N_11758);
and U12118 (N_12118,N_11988,N_11759);
nor U12119 (N_12119,N_11813,N_11963);
and U12120 (N_12120,N_11753,N_11836);
nand U12121 (N_12121,N_11877,N_11908);
nor U12122 (N_12122,N_11973,N_11990);
and U12123 (N_12123,N_11757,N_11916);
and U12124 (N_12124,N_11985,N_11834);
nand U12125 (N_12125,N_11983,N_11959);
or U12126 (N_12126,N_11959,N_11904);
nor U12127 (N_12127,N_11917,N_11973);
and U12128 (N_12128,N_11805,N_11833);
or U12129 (N_12129,N_11876,N_11875);
nand U12130 (N_12130,N_11925,N_11935);
and U12131 (N_12131,N_11794,N_11955);
and U12132 (N_12132,N_11985,N_11909);
or U12133 (N_12133,N_11994,N_11779);
or U12134 (N_12134,N_11862,N_11804);
nand U12135 (N_12135,N_11884,N_11854);
or U12136 (N_12136,N_11977,N_11782);
or U12137 (N_12137,N_11757,N_11933);
nor U12138 (N_12138,N_11906,N_11911);
and U12139 (N_12139,N_11754,N_11874);
and U12140 (N_12140,N_11867,N_11863);
nand U12141 (N_12141,N_11797,N_11941);
nor U12142 (N_12142,N_11932,N_11853);
or U12143 (N_12143,N_11863,N_11855);
xnor U12144 (N_12144,N_11798,N_11852);
nor U12145 (N_12145,N_11802,N_11859);
and U12146 (N_12146,N_11991,N_11770);
and U12147 (N_12147,N_11946,N_11834);
nor U12148 (N_12148,N_11818,N_11938);
and U12149 (N_12149,N_11793,N_11782);
and U12150 (N_12150,N_11855,N_11940);
nand U12151 (N_12151,N_11901,N_11871);
and U12152 (N_12152,N_11959,N_11970);
or U12153 (N_12153,N_11793,N_11951);
and U12154 (N_12154,N_11936,N_11751);
nor U12155 (N_12155,N_11899,N_11839);
nand U12156 (N_12156,N_11925,N_11907);
xnor U12157 (N_12157,N_11939,N_11940);
and U12158 (N_12158,N_11770,N_11820);
or U12159 (N_12159,N_11982,N_11858);
or U12160 (N_12160,N_11790,N_11777);
nand U12161 (N_12161,N_11903,N_11857);
nand U12162 (N_12162,N_11932,N_11836);
nor U12163 (N_12163,N_11915,N_11881);
nand U12164 (N_12164,N_11946,N_11760);
nor U12165 (N_12165,N_11838,N_11756);
nor U12166 (N_12166,N_11820,N_11883);
and U12167 (N_12167,N_11796,N_11922);
and U12168 (N_12168,N_11989,N_11757);
xor U12169 (N_12169,N_11817,N_11766);
nand U12170 (N_12170,N_11993,N_11841);
nand U12171 (N_12171,N_11795,N_11999);
or U12172 (N_12172,N_11807,N_11923);
xor U12173 (N_12173,N_11979,N_11881);
and U12174 (N_12174,N_11904,N_11917);
nand U12175 (N_12175,N_11858,N_11811);
and U12176 (N_12176,N_11853,N_11760);
and U12177 (N_12177,N_11845,N_11931);
or U12178 (N_12178,N_11942,N_11856);
nor U12179 (N_12179,N_11875,N_11759);
and U12180 (N_12180,N_11814,N_11938);
or U12181 (N_12181,N_11887,N_11842);
nand U12182 (N_12182,N_11769,N_11864);
nand U12183 (N_12183,N_11844,N_11928);
and U12184 (N_12184,N_11799,N_11815);
or U12185 (N_12185,N_11956,N_11986);
nor U12186 (N_12186,N_11839,N_11911);
nor U12187 (N_12187,N_11832,N_11997);
nand U12188 (N_12188,N_11861,N_11761);
and U12189 (N_12189,N_11777,N_11975);
nor U12190 (N_12190,N_11977,N_11917);
nand U12191 (N_12191,N_11767,N_11837);
nand U12192 (N_12192,N_11890,N_11968);
and U12193 (N_12193,N_11981,N_11817);
nor U12194 (N_12194,N_11790,N_11778);
nand U12195 (N_12195,N_11832,N_11972);
nor U12196 (N_12196,N_11903,N_11754);
nor U12197 (N_12197,N_11766,N_11975);
and U12198 (N_12198,N_11815,N_11814);
or U12199 (N_12199,N_11770,N_11817);
and U12200 (N_12200,N_11942,N_11823);
and U12201 (N_12201,N_11866,N_11879);
nand U12202 (N_12202,N_11991,N_11981);
nor U12203 (N_12203,N_11888,N_11764);
nor U12204 (N_12204,N_11988,N_11840);
nor U12205 (N_12205,N_11935,N_11948);
nor U12206 (N_12206,N_11966,N_11992);
or U12207 (N_12207,N_11892,N_11833);
xor U12208 (N_12208,N_11920,N_11995);
nand U12209 (N_12209,N_11784,N_11798);
nand U12210 (N_12210,N_11965,N_11959);
or U12211 (N_12211,N_11989,N_11880);
or U12212 (N_12212,N_11825,N_11793);
nor U12213 (N_12213,N_11997,N_11851);
or U12214 (N_12214,N_11858,N_11845);
nand U12215 (N_12215,N_11775,N_11758);
nand U12216 (N_12216,N_11875,N_11788);
nand U12217 (N_12217,N_11877,N_11794);
or U12218 (N_12218,N_11958,N_11944);
and U12219 (N_12219,N_11831,N_11981);
and U12220 (N_12220,N_11959,N_11843);
or U12221 (N_12221,N_11954,N_11931);
and U12222 (N_12222,N_11933,N_11764);
xor U12223 (N_12223,N_11963,N_11926);
nand U12224 (N_12224,N_11865,N_11952);
nor U12225 (N_12225,N_11845,N_11955);
or U12226 (N_12226,N_11916,N_11842);
and U12227 (N_12227,N_11873,N_11934);
nand U12228 (N_12228,N_11919,N_11796);
or U12229 (N_12229,N_11950,N_11824);
xnor U12230 (N_12230,N_11946,N_11952);
nor U12231 (N_12231,N_11852,N_11899);
nor U12232 (N_12232,N_11800,N_11848);
nor U12233 (N_12233,N_11895,N_11900);
nor U12234 (N_12234,N_11786,N_11797);
and U12235 (N_12235,N_11812,N_11779);
nand U12236 (N_12236,N_11885,N_11787);
and U12237 (N_12237,N_11953,N_11858);
xor U12238 (N_12238,N_11999,N_11823);
and U12239 (N_12239,N_11862,N_11756);
and U12240 (N_12240,N_11983,N_11752);
and U12241 (N_12241,N_11998,N_11903);
nor U12242 (N_12242,N_11941,N_11957);
nor U12243 (N_12243,N_11915,N_11844);
nand U12244 (N_12244,N_11818,N_11978);
and U12245 (N_12245,N_11868,N_11912);
nor U12246 (N_12246,N_11951,N_11909);
nor U12247 (N_12247,N_11780,N_11989);
nor U12248 (N_12248,N_11992,N_11815);
or U12249 (N_12249,N_11962,N_11923);
nand U12250 (N_12250,N_12187,N_12182);
nand U12251 (N_12251,N_12152,N_12243);
or U12252 (N_12252,N_12203,N_12193);
xor U12253 (N_12253,N_12127,N_12037);
and U12254 (N_12254,N_12188,N_12020);
and U12255 (N_12255,N_12007,N_12247);
and U12256 (N_12256,N_12015,N_12008);
xor U12257 (N_12257,N_12110,N_12028);
nand U12258 (N_12258,N_12150,N_12240);
xor U12259 (N_12259,N_12124,N_12135);
nor U12260 (N_12260,N_12225,N_12047);
and U12261 (N_12261,N_12083,N_12231);
and U12262 (N_12262,N_12016,N_12222);
nor U12263 (N_12263,N_12035,N_12245);
xnor U12264 (N_12264,N_12244,N_12073);
nand U12265 (N_12265,N_12079,N_12153);
nand U12266 (N_12266,N_12197,N_12145);
and U12267 (N_12267,N_12022,N_12040);
nor U12268 (N_12268,N_12216,N_12185);
and U12269 (N_12269,N_12012,N_12190);
and U12270 (N_12270,N_12043,N_12238);
nor U12271 (N_12271,N_12180,N_12075);
nand U12272 (N_12272,N_12181,N_12171);
nor U12273 (N_12273,N_12018,N_12233);
and U12274 (N_12274,N_12101,N_12228);
and U12275 (N_12275,N_12239,N_12144);
nor U12276 (N_12276,N_12177,N_12086);
nor U12277 (N_12277,N_12207,N_12049);
nand U12278 (N_12278,N_12092,N_12024);
and U12279 (N_12279,N_12149,N_12192);
or U12280 (N_12280,N_12045,N_12178);
nand U12281 (N_12281,N_12036,N_12089);
or U12282 (N_12282,N_12057,N_12219);
and U12283 (N_12283,N_12074,N_12235);
xnor U12284 (N_12284,N_12082,N_12196);
nor U12285 (N_12285,N_12179,N_12053);
or U12286 (N_12286,N_12170,N_12148);
nand U12287 (N_12287,N_12199,N_12044);
xnor U12288 (N_12288,N_12098,N_12194);
and U12289 (N_12289,N_12224,N_12003);
nor U12290 (N_12290,N_12106,N_12102);
nor U12291 (N_12291,N_12195,N_12121);
nor U12292 (N_12292,N_12052,N_12155);
and U12293 (N_12293,N_12031,N_12010);
nand U12294 (N_12294,N_12234,N_12019);
nand U12295 (N_12295,N_12107,N_12054);
or U12296 (N_12296,N_12087,N_12151);
nand U12297 (N_12297,N_12004,N_12061);
or U12298 (N_12298,N_12162,N_12189);
nand U12299 (N_12299,N_12038,N_12223);
nand U12300 (N_12300,N_12030,N_12058);
nand U12301 (N_12301,N_12112,N_12117);
nand U12302 (N_12302,N_12129,N_12146);
or U12303 (N_12303,N_12227,N_12116);
nand U12304 (N_12304,N_12120,N_12130);
nor U12305 (N_12305,N_12159,N_12081);
or U12306 (N_12306,N_12248,N_12023);
or U12307 (N_12307,N_12201,N_12209);
or U12308 (N_12308,N_12068,N_12137);
xor U12309 (N_12309,N_12128,N_12033);
or U12310 (N_12310,N_12034,N_12100);
xor U12311 (N_12311,N_12039,N_12021);
xnor U12312 (N_12312,N_12183,N_12133);
nand U12313 (N_12313,N_12080,N_12096);
or U12314 (N_12314,N_12208,N_12164);
and U12315 (N_12315,N_12184,N_12090);
xor U12316 (N_12316,N_12191,N_12095);
and U12317 (N_12317,N_12161,N_12204);
nor U12318 (N_12318,N_12111,N_12168);
nand U12319 (N_12319,N_12006,N_12026);
nand U12320 (N_12320,N_12115,N_12143);
nand U12321 (N_12321,N_12139,N_12114);
xnor U12322 (N_12322,N_12085,N_12217);
or U12323 (N_12323,N_12041,N_12202);
nor U12324 (N_12324,N_12165,N_12205);
and U12325 (N_12325,N_12241,N_12025);
nand U12326 (N_12326,N_12062,N_12104);
and U12327 (N_12327,N_12136,N_12051);
nand U12328 (N_12328,N_12002,N_12186);
nor U12329 (N_12329,N_12131,N_12154);
nor U12330 (N_12330,N_12071,N_12230);
or U12331 (N_12331,N_12229,N_12105);
and U12332 (N_12332,N_12066,N_12046);
nand U12333 (N_12333,N_12138,N_12059);
nand U12334 (N_12334,N_12005,N_12042);
nand U12335 (N_12335,N_12220,N_12174);
nand U12336 (N_12336,N_12166,N_12147);
or U12337 (N_12337,N_12122,N_12014);
or U12338 (N_12338,N_12076,N_12027);
and U12339 (N_12339,N_12064,N_12176);
and U12340 (N_12340,N_12063,N_12132);
and U12341 (N_12341,N_12212,N_12001);
nand U12342 (N_12342,N_12211,N_12077);
or U12343 (N_12343,N_12125,N_12242);
nand U12344 (N_12344,N_12175,N_12070);
and U12345 (N_12345,N_12097,N_12091);
nand U12346 (N_12346,N_12093,N_12032);
xor U12347 (N_12347,N_12246,N_12213);
nand U12348 (N_12348,N_12249,N_12078);
nand U12349 (N_12349,N_12119,N_12067);
nand U12350 (N_12350,N_12055,N_12134);
nor U12351 (N_12351,N_12167,N_12226);
nor U12352 (N_12352,N_12084,N_12017);
xnor U12353 (N_12353,N_12065,N_12232);
or U12354 (N_12354,N_12156,N_12237);
and U12355 (N_12355,N_12013,N_12088);
nor U12356 (N_12356,N_12123,N_12103);
nand U12357 (N_12357,N_12158,N_12140);
and U12358 (N_12358,N_12160,N_12126);
xnor U12359 (N_12359,N_12029,N_12214);
and U12360 (N_12360,N_12218,N_12236);
or U12361 (N_12361,N_12157,N_12173);
nor U12362 (N_12362,N_12048,N_12009);
and U12363 (N_12363,N_12050,N_12215);
nor U12364 (N_12364,N_12069,N_12200);
or U12365 (N_12365,N_12206,N_12169);
and U12366 (N_12366,N_12060,N_12000);
nand U12367 (N_12367,N_12142,N_12099);
nand U12368 (N_12368,N_12113,N_12072);
or U12369 (N_12369,N_12163,N_12141);
or U12370 (N_12370,N_12210,N_12198);
xnor U12371 (N_12371,N_12056,N_12221);
and U12372 (N_12372,N_12109,N_12108);
nand U12373 (N_12373,N_12094,N_12118);
or U12374 (N_12374,N_12172,N_12011);
and U12375 (N_12375,N_12069,N_12010);
nand U12376 (N_12376,N_12191,N_12154);
and U12377 (N_12377,N_12122,N_12040);
or U12378 (N_12378,N_12195,N_12079);
or U12379 (N_12379,N_12239,N_12054);
or U12380 (N_12380,N_12197,N_12056);
or U12381 (N_12381,N_12068,N_12008);
xnor U12382 (N_12382,N_12078,N_12130);
and U12383 (N_12383,N_12089,N_12159);
and U12384 (N_12384,N_12240,N_12173);
nand U12385 (N_12385,N_12131,N_12165);
nand U12386 (N_12386,N_12210,N_12141);
nand U12387 (N_12387,N_12097,N_12159);
nand U12388 (N_12388,N_12182,N_12217);
xor U12389 (N_12389,N_12153,N_12120);
xnor U12390 (N_12390,N_12224,N_12084);
and U12391 (N_12391,N_12043,N_12088);
and U12392 (N_12392,N_12045,N_12234);
nand U12393 (N_12393,N_12212,N_12042);
nand U12394 (N_12394,N_12053,N_12135);
nor U12395 (N_12395,N_12078,N_12171);
or U12396 (N_12396,N_12192,N_12044);
or U12397 (N_12397,N_12137,N_12039);
nand U12398 (N_12398,N_12147,N_12109);
xor U12399 (N_12399,N_12219,N_12174);
or U12400 (N_12400,N_12129,N_12242);
nand U12401 (N_12401,N_12184,N_12029);
nor U12402 (N_12402,N_12202,N_12174);
or U12403 (N_12403,N_12033,N_12210);
or U12404 (N_12404,N_12219,N_12157);
and U12405 (N_12405,N_12175,N_12076);
and U12406 (N_12406,N_12182,N_12199);
and U12407 (N_12407,N_12198,N_12036);
nand U12408 (N_12408,N_12130,N_12246);
nand U12409 (N_12409,N_12076,N_12099);
nand U12410 (N_12410,N_12033,N_12029);
nor U12411 (N_12411,N_12215,N_12177);
nor U12412 (N_12412,N_12073,N_12066);
or U12413 (N_12413,N_12023,N_12204);
nand U12414 (N_12414,N_12094,N_12107);
nor U12415 (N_12415,N_12216,N_12125);
and U12416 (N_12416,N_12106,N_12154);
and U12417 (N_12417,N_12096,N_12062);
nand U12418 (N_12418,N_12100,N_12131);
nor U12419 (N_12419,N_12089,N_12247);
nand U12420 (N_12420,N_12047,N_12041);
nor U12421 (N_12421,N_12121,N_12247);
or U12422 (N_12422,N_12144,N_12132);
nand U12423 (N_12423,N_12161,N_12024);
nand U12424 (N_12424,N_12132,N_12149);
and U12425 (N_12425,N_12249,N_12107);
xor U12426 (N_12426,N_12005,N_12212);
or U12427 (N_12427,N_12233,N_12080);
and U12428 (N_12428,N_12158,N_12149);
xnor U12429 (N_12429,N_12038,N_12080);
nand U12430 (N_12430,N_12156,N_12094);
and U12431 (N_12431,N_12059,N_12171);
xor U12432 (N_12432,N_12013,N_12048);
or U12433 (N_12433,N_12129,N_12213);
nand U12434 (N_12434,N_12165,N_12187);
and U12435 (N_12435,N_12144,N_12158);
or U12436 (N_12436,N_12123,N_12025);
xnor U12437 (N_12437,N_12158,N_12142);
nor U12438 (N_12438,N_12055,N_12029);
and U12439 (N_12439,N_12041,N_12246);
nor U12440 (N_12440,N_12132,N_12022);
and U12441 (N_12441,N_12152,N_12186);
nand U12442 (N_12442,N_12131,N_12044);
nand U12443 (N_12443,N_12088,N_12087);
nor U12444 (N_12444,N_12126,N_12117);
or U12445 (N_12445,N_12048,N_12063);
or U12446 (N_12446,N_12195,N_12169);
nor U12447 (N_12447,N_12199,N_12029);
or U12448 (N_12448,N_12244,N_12164);
or U12449 (N_12449,N_12068,N_12027);
and U12450 (N_12450,N_12183,N_12072);
or U12451 (N_12451,N_12204,N_12123);
and U12452 (N_12452,N_12016,N_12021);
or U12453 (N_12453,N_12119,N_12052);
and U12454 (N_12454,N_12169,N_12213);
and U12455 (N_12455,N_12212,N_12097);
nand U12456 (N_12456,N_12044,N_12224);
nand U12457 (N_12457,N_12188,N_12133);
or U12458 (N_12458,N_12020,N_12155);
nor U12459 (N_12459,N_12006,N_12204);
nand U12460 (N_12460,N_12070,N_12045);
xor U12461 (N_12461,N_12116,N_12043);
nor U12462 (N_12462,N_12014,N_12083);
xor U12463 (N_12463,N_12210,N_12034);
nand U12464 (N_12464,N_12142,N_12094);
or U12465 (N_12465,N_12018,N_12079);
nor U12466 (N_12466,N_12212,N_12076);
or U12467 (N_12467,N_12180,N_12143);
xor U12468 (N_12468,N_12241,N_12243);
nor U12469 (N_12469,N_12078,N_12057);
or U12470 (N_12470,N_12048,N_12001);
nand U12471 (N_12471,N_12137,N_12243);
or U12472 (N_12472,N_12124,N_12213);
and U12473 (N_12473,N_12173,N_12029);
nor U12474 (N_12474,N_12080,N_12144);
nor U12475 (N_12475,N_12169,N_12200);
nand U12476 (N_12476,N_12220,N_12134);
nor U12477 (N_12477,N_12122,N_12009);
or U12478 (N_12478,N_12148,N_12085);
xnor U12479 (N_12479,N_12200,N_12029);
nand U12480 (N_12480,N_12076,N_12176);
nand U12481 (N_12481,N_12067,N_12029);
and U12482 (N_12482,N_12112,N_12158);
or U12483 (N_12483,N_12080,N_12159);
and U12484 (N_12484,N_12107,N_12160);
xor U12485 (N_12485,N_12192,N_12167);
or U12486 (N_12486,N_12216,N_12190);
or U12487 (N_12487,N_12082,N_12214);
or U12488 (N_12488,N_12129,N_12014);
and U12489 (N_12489,N_12146,N_12009);
nor U12490 (N_12490,N_12098,N_12064);
nand U12491 (N_12491,N_12088,N_12218);
nand U12492 (N_12492,N_12243,N_12107);
nor U12493 (N_12493,N_12113,N_12244);
nand U12494 (N_12494,N_12160,N_12001);
xnor U12495 (N_12495,N_12016,N_12122);
nand U12496 (N_12496,N_12198,N_12241);
and U12497 (N_12497,N_12112,N_12186);
and U12498 (N_12498,N_12084,N_12007);
xnor U12499 (N_12499,N_12224,N_12057);
and U12500 (N_12500,N_12330,N_12458);
nand U12501 (N_12501,N_12311,N_12377);
or U12502 (N_12502,N_12362,N_12485);
or U12503 (N_12503,N_12290,N_12279);
nor U12504 (N_12504,N_12402,N_12304);
nor U12505 (N_12505,N_12379,N_12498);
and U12506 (N_12506,N_12338,N_12334);
or U12507 (N_12507,N_12324,N_12447);
nand U12508 (N_12508,N_12488,N_12360);
xor U12509 (N_12509,N_12481,N_12435);
and U12510 (N_12510,N_12348,N_12342);
xnor U12511 (N_12511,N_12388,N_12321);
and U12512 (N_12512,N_12349,N_12415);
nor U12513 (N_12513,N_12476,N_12448);
nor U12514 (N_12514,N_12474,N_12264);
or U12515 (N_12515,N_12392,N_12370);
and U12516 (N_12516,N_12433,N_12440);
or U12517 (N_12517,N_12420,N_12390);
nand U12518 (N_12518,N_12254,N_12442);
or U12519 (N_12519,N_12278,N_12315);
and U12520 (N_12520,N_12371,N_12261);
nor U12521 (N_12521,N_12364,N_12475);
nand U12522 (N_12522,N_12367,N_12266);
or U12523 (N_12523,N_12387,N_12359);
and U12524 (N_12524,N_12332,N_12470);
and U12525 (N_12525,N_12312,N_12272);
and U12526 (N_12526,N_12375,N_12283);
nor U12527 (N_12527,N_12428,N_12309);
or U12528 (N_12528,N_12449,N_12437);
or U12529 (N_12529,N_12483,N_12352);
nor U12530 (N_12530,N_12372,N_12471);
and U12531 (N_12531,N_12412,N_12275);
and U12532 (N_12532,N_12429,N_12457);
nand U12533 (N_12533,N_12368,N_12282);
nand U12534 (N_12534,N_12381,N_12285);
and U12535 (N_12535,N_12487,N_12284);
nor U12536 (N_12536,N_12306,N_12409);
or U12537 (N_12537,N_12413,N_12462);
or U12538 (N_12538,N_12453,N_12408);
nand U12539 (N_12539,N_12347,N_12373);
or U12540 (N_12540,N_12451,N_12329);
and U12541 (N_12541,N_12361,N_12291);
or U12542 (N_12542,N_12477,N_12496);
and U12543 (N_12543,N_12494,N_12469);
and U12544 (N_12544,N_12489,N_12386);
nand U12545 (N_12545,N_12465,N_12389);
nor U12546 (N_12546,N_12490,N_12380);
xor U12547 (N_12547,N_12436,N_12473);
and U12548 (N_12548,N_12400,N_12423);
or U12549 (N_12549,N_12450,N_12363);
nand U12550 (N_12550,N_12317,N_12397);
xor U12551 (N_12551,N_12406,N_12365);
or U12552 (N_12552,N_12350,N_12425);
nand U12553 (N_12553,N_12461,N_12258);
xor U12554 (N_12554,N_12288,N_12444);
or U12555 (N_12555,N_12314,N_12382);
nor U12556 (N_12556,N_12289,N_12274);
nor U12557 (N_12557,N_12252,N_12426);
or U12558 (N_12558,N_12346,N_12286);
or U12559 (N_12559,N_12486,N_12333);
nand U12560 (N_12560,N_12293,N_12260);
nor U12561 (N_12561,N_12398,N_12302);
nor U12562 (N_12562,N_12335,N_12292);
nand U12563 (N_12563,N_12299,N_12401);
nand U12564 (N_12564,N_12438,N_12434);
or U12565 (N_12565,N_12493,N_12280);
nand U12566 (N_12566,N_12472,N_12424);
and U12567 (N_12567,N_12456,N_12326);
nand U12568 (N_12568,N_12405,N_12296);
nor U12569 (N_12569,N_12267,N_12439);
and U12570 (N_12570,N_12407,N_12259);
or U12571 (N_12571,N_12336,N_12313);
nor U12572 (N_12572,N_12298,N_12403);
or U12573 (N_12573,N_12432,N_12301);
and U12574 (N_12574,N_12480,N_12418);
or U12575 (N_12575,N_12263,N_12353);
nand U12576 (N_12576,N_12253,N_12460);
nand U12577 (N_12577,N_12297,N_12499);
and U12578 (N_12578,N_12325,N_12497);
nand U12579 (N_12579,N_12351,N_12310);
nor U12580 (N_12580,N_12356,N_12300);
or U12581 (N_12581,N_12273,N_12337);
nor U12582 (N_12582,N_12467,N_12416);
nor U12583 (N_12583,N_12340,N_12294);
and U12584 (N_12584,N_12250,N_12445);
nand U12585 (N_12585,N_12464,N_12478);
or U12586 (N_12586,N_12251,N_12354);
nor U12587 (N_12587,N_12305,N_12417);
or U12588 (N_12588,N_12410,N_12441);
xor U12589 (N_12589,N_12262,N_12399);
nand U12590 (N_12590,N_12421,N_12318);
or U12591 (N_12591,N_12358,N_12307);
nor U12592 (N_12592,N_12265,N_12303);
nand U12593 (N_12593,N_12277,N_12491);
or U12594 (N_12594,N_12446,N_12308);
nor U12595 (N_12595,N_12404,N_12454);
nand U12596 (N_12596,N_12270,N_12414);
or U12597 (N_12597,N_12331,N_12452);
or U12598 (N_12598,N_12427,N_12484);
or U12599 (N_12599,N_12355,N_12271);
nor U12600 (N_12600,N_12256,N_12411);
nor U12601 (N_12601,N_12327,N_12492);
or U12602 (N_12602,N_12495,N_12395);
nand U12603 (N_12603,N_12384,N_12369);
nand U12604 (N_12604,N_12466,N_12393);
or U12605 (N_12605,N_12455,N_12383);
or U12606 (N_12606,N_12479,N_12339);
nand U12607 (N_12607,N_12468,N_12255);
or U12608 (N_12608,N_12385,N_12268);
or U12609 (N_12609,N_12394,N_12443);
nand U12610 (N_12610,N_12463,N_12343);
nand U12611 (N_12611,N_12482,N_12345);
and U12612 (N_12612,N_12459,N_12276);
or U12613 (N_12613,N_12328,N_12419);
nor U12614 (N_12614,N_12391,N_12269);
nand U12615 (N_12615,N_12430,N_12422);
nand U12616 (N_12616,N_12322,N_12281);
xor U12617 (N_12617,N_12316,N_12378);
or U12618 (N_12618,N_12366,N_12374);
xor U12619 (N_12619,N_12344,N_12319);
xor U12620 (N_12620,N_12357,N_12323);
xor U12621 (N_12621,N_12431,N_12376);
nor U12622 (N_12622,N_12257,N_12295);
or U12623 (N_12623,N_12341,N_12287);
and U12624 (N_12624,N_12396,N_12320);
nand U12625 (N_12625,N_12345,N_12460);
and U12626 (N_12626,N_12417,N_12316);
or U12627 (N_12627,N_12346,N_12257);
nand U12628 (N_12628,N_12441,N_12330);
nand U12629 (N_12629,N_12305,N_12473);
and U12630 (N_12630,N_12440,N_12437);
or U12631 (N_12631,N_12425,N_12264);
nand U12632 (N_12632,N_12419,N_12475);
or U12633 (N_12633,N_12438,N_12454);
nor U12634 (N_12634,N_12480,N_12394);
or U12635 (N_12635,N_12389,N_12359);
xor U12636 (N_12636,N_12302,N_12445);
and U12637 (N_12637,N_12316,N_12390);
and U12638 (N_12638,N_12313,N_12356);
and U12639 (N_12639,N_12418,N_12328);
nand U12640 (N_12640,N_12398,N_12429);
nor U12641 (N_12641,N_12295,N_12261);
or U12642 (N_12642,N_12358,N_12413);
and U12643 (N_12643,N_12445,N_12475);
nand U12644 (N_12644,N_12328,N_12261);
or U12645 (N_12645,N_12494,N_12386);
and U12646 (N_12646,N_12417,N_12403);
nor U12647 (N_12647,N_12291,N_12443);
nor U12648 (N_12648,N_12327,N_12384);
and U12649 (N_12649,N_12274,N_12252);
and U12650 (N_12650,N_12456,N_12435);
or U12651 (N_12651,N_12305,N_12468);
or U12652 (N_12652,N_12269,N_12451);
nand U12653 (N_12653,N_12308,N_12489);
and U12654 (N_12654,N_12446,N_12494);
nor U12655 (N_12655,N_12257,N_12481);
or U12656 (N_12656,N_12420,N_12319);
and U12657 (N_12657,N_12417,N_12433);
nand U12658 (N_12658,N_12304,N_12461);
or U12659 (N_12659,N_12426,N_12251);
or U12660 (N_12660,N_12431,N_12396);
and U12661 (N_12661,N_12415,N_12492);
nor U12662 (N_12662,N_12469,N_12374);
nor U12663 (N_12663,N_12412,N_12408);
or U12664 (N_12664,N_12408,N_12388);
nor U12665 (N_12665,N_12397,N_12440);
or U12666 (N_12666,N_12357,N_12467);
nand U12667 (N_12667,N_12474,N_12437);
and U12668 (N_12668,N_12482,N_12264);
nor U12669 (N_12669,N_12316,N_12335);
xnor U12670 (N_12670,N_12306,N_12452);
and U12671 (N_12671,N_12489,N_12366);
and U12672 (N_12672,N_12454,N_12334);
nor U12673 (N_12673,N_12336,N_12455);
and U12674 (N_12674,N_12278,N_12479);
and U12675 (N_12675,N_12431,N_12498);
nand U12676 (N_12676,N_12419,N_12458);
and U12677 (N_12677,N_12361,N_12480);
and U12678 (N_12678,N_12296,N_12445);
and U12679 (N_12679,N_12454,N_12391);
nand U12680 (N_12680,N_12413,N_12488);
nor U12681 (N_12681,N_12394,N_12321);
nor U12682 (N_12682,N_12393,N_12416);
nand U12683 (N_12683,N_12316,N_12452);
nor U12684 (N_12684,N_12332,N_12483);
and U12685 (N_12685,N_12320,N_12258);
nor U12686 (N_12686,N_12367,N_12330);
nor U12687 (N_12687,N_12355,N_12452);
nor U12688 (N_12688,N_12330,N_12321);
nand U12689 (N_12689,N_12353,N_12369);
nand U12690 (N_12690,N_12490,N_12456);
or U12691 (N_12691,N_12366,N_12400);
nand U12692 (N_12692,N_12255,N_12478);
and U12693 (N_12693,N_12293,N_12271);
and U12694 (N_12694,N_12423,N_12421);
and U12695 (N_12695,N_12356,N_12315);
nand U12696 (N_12696,N_12481,N_12321);
or U12697 (N_12697,N_12331,N_12382);
nand U12698 (N_12698,N_12417,N_12325);
and U12699 (N_12699,N_12465,N_12317);
and U12700 (N_12700,N_12380,N_12294);
and U12701 (N_12701,N_12300,N_12359);
nand U12702 (N_12702,N_12305,N_12379);
or U12703 (N_12703,N_12362,N_12399);
or U12704 (N_12704,N_12450,N_12456);
or U12705 (N_12705,N_12377,N_12407);
xor U12706 (N_12706,N_12416,N_12304);
or U12707 (N_12707,N_12424,N_12402);
nor U12708 (N_12708,N_12381,N_12281);
xnor U12709 (N_12709,N_12347,N_12340);
nand U12710 (N_12710,N_12286,N_12482);
nand U12711 (N_12711,N_12394,N_12267);
nor U12712 (N_12712,N_12467,N_12280);
or U12713 (N_12713,N_12490,N_12384);
nand U12714 (N_12714,N_12255,N_12360);
xor U12715 (N_12715,N_12330,N_12284);
nand U12716 (N_12716,N_12471,N_12409);
nor U12717 (N_12717,N_12341,N_12402);
nor U12718 (N_12718,N_12260,N_12258);
or U12719 (N_12719,N_12434,N_12451);
or U12720 (N_12720,N_12487,N_12485);
or U12721 (N_12721,N_12357,N_12458);
nand U12722 (N_12722,N_12439,N_12292);
and U12723 (N_12723,N_12380,N_12297);
nand U12724 (N_12724,N_12280,N_12343);
and U12725 (N_12725,N_12328,N_12467);
nand U12726 (N_12726,N_12251,N_12317);
nor U12727 (N_12727,N_12426,N_12337);
xor U12728 (N_12728,N_12430,N_12457);
and U12729 (N_12729,N_12452,N_12432);
or U12730 (N_12730,N_12345,N_12310);
nand U12731 (N_12731,N_12494,N_12322);
and U12732 (N_12732,N_12414,N_12493);
and U12733 (N_12733,N_12445,N_12349);
or U12734 (N_12734,N_12301,N_12410);
and U12735 (N_12735,N_12433,N_12366);
nand U12736 (N_12736,N_12296,N_12334);
nor U12737 (N_12737,N_12298,N_12276);
nor U12738 (N_12738,N_12254,N_12295);
and U12739 (N_12739,N_12443,N_12455);
nand U12740 (N_12740,N_12445,N_12342);
and U12741 (N_12741,N_12352,N_12420);
xnor U12742 (N_12742,N_12472,N_12355);
or U12743 (N_12743,N_12325,N_12314);
and U12744 (N_12744,N_12286,N_12493);
nand U12745 (N_12745,N_12281,N_12300);
or U12746 (N_12746,N_12258,N_12490);
nor U12747 (N_12747,N_12442,N_12407);
xnor U12748 (N_12748,N_12387,N_12485);
nor U12749 (N_12749,N_12269,N_12360);
or U12750 (N_12750,N_12559,N_12728);
nor U12751 (N_12751,N_12741,N_12658);
and U12752 (N_12752,N_12568,N_12727);
nand U12753 (N_12753,N_12512,N_12744);
nand U12754 (N_12754,N_12607,N_12710);
or U12755 (N_12755,N_12694,N_12587);
nand U12756 (N_12756,N_12716,N_12505);
or U12757 (N_12757,N_12507,N_12611);
nor U12758 (N_12758,N_12628,N_12686);
or U12759 (N_12759,N_12519,N_12683);
or U12760 (N_12760,N_12502,N_12506);
or U12761 (N_12761,N_12558,N_12583);
nor U12762 (N_12762,N_12682,N_12678);
nand U12763 (N_12763,N_12580,N_12545);
nor U12764 (N_12764,N_12712,N_12711);
and U12765 (N_12765,N_12622,N_12567);
nor U12766 (N_12766,N_12717,N_12597);
and U12767 (N_12767,N_12518,N_12608);
or U12768 (N_12768,N_12586,N_12569);
xor U12769 (N_12769,N_12614,N_12644);
or U12770 (N_12770,N_12613,N_12537);
or U12771 (N_12771,N_12721,N_12737);
and U12772 (N_12772,N_12630,N_12731);
nand U12773 (N_12773,N_12536,N_12632);
xnor U12774 (N_12774,N_12531,N_12603);
and U12775 (N_12775,N_12680,N_12570);
nor U12776 (N_12776,N_12525,N_12604);
or U12777 (N_12777,N_12551,N_12688);
or U12778 (N_12778,N_12701,N_12708);
and U12779 (N_12779,N_12585,N_12535);
and U12780 (N_12780,N_12692,N_12740);
nor U12781 (N_12781,N_12641,N_12655);
and U12782 (N_12782,N_12696,N_12500);
nand U12783 (N_12783,N_12550,N_12543);
and U12784 (N_12784,N_12511,N_12725);
or U12785 (N_12785,N_12730,N_12625);
and U12786 (N_12786,N_12733,N_12662);
and U12787 (N_12787,N_12602,N_12668);
and U12788 (N_12788,N_12629,N_12726);
nand U12789 (N_12789,N_12561,N_12738);
xnor U12790 (N_12790,N_12690,N_12685);
nor U12791 (N_12791,N_12574,N_12554);
or U12792 (N_12792,N_12745,N_12749);
or U12793 (N_12793,N_12566,N_12647);
xnor U12794 (N_12794,N_12703,N_12687);
xor U12795 (N_12795,N_12547,N_12532);
and U12796 (N_12796,N_12538,N_12544);
nor U12797 (N_12797,N_12578,N_12513);
or U12798 (N_12798,N_12573,N_12705);
or U12799 (N_12799,N_12526,N_12504);
nor U12800 (N_12800,N_12640,N_12510);
nand U12801 (N_12801,N_12645,N_12508);
xor U12802 (N_12802,N_12673,N_12563);
and U12803 (N_12803,N_12528,N_12706);
nand U12804 (N_12804,N_12530,N_12605);
nand U12805 (N_12805,N_12557,N_12575);
xnor U12806 (N_12806,N_12729,N_12619);
nand U12807 (N_12807,N_12634,N_12656);
nor U12808 (N_12808,N_12572,N_12618);
xor U12809 (N_12809,N_12514,N_12631);
nor U12810 (N_12810,N_12612,N_12719);
nand U12811 (N_12811,N_12732,N_12643);
or U12812 (N_12812,N_12679,N_12691);
nor U12813 (N_12813,N_12689,N_12649);
or U12814 (N_12814,N_12665,N_12577);
or U12815 (N_12815,N_12589,N_12722);
nor U12816 (N_12816,N_12675,N_12609);
nand U12817 (N_12817,N_12592,N_12661);
or U12818 (N_12818,N_12638,N_12642);
nand U12819 (N_12819,N_12534,N_12540);
nor U12820 (N_12820,N_12714,N_12624);
xnor U12821 (N_12821,N_12746,N_12501);
and U12822 (N_12822,N_12677,N_12527);
and U12823 (N_12823,N_12659,N_12582);
or U12824 (N_12824,N_12523,N_12562);
nand U12825 (N_12825,N_12541,N_12684);
and U12826 (N_12826,N_12529,N_12657);
nand U12827 (N_12827,N_12584,N_12713);
or U12828 (N_12828,N_12588,N_12595);
or U12829 (N_12829,N_12698,N_12593);
nand U12830 (N_12830,N_12555,N_12548);
and U12831 (N_12831,N_12702,N_12669);
nand U12832 (N_12832,N_12620,N_12697);
and U12833 (N_12833,N_12546,N_12533);
nand U12834 (N_12834,N_12742,N_12598);
and U12835 (N_12835,N_12650,N_12503);
nand U12836 (N_12836,N_12633,N_12664);
nor U12837 (N_12837,N_12600,N_12542);
nor U12838 (N_12838,N_12700,N_12581);
or U12839 (N_12839,N_12695,N_12672);
xnor U12840 (N_12840,N_12709,N_12539);
nand U12841 (N_12841,N_12648,N_12653);
nor U12842 (N_12842,N_12670,N_12623);
or U12843 (N_12843,N_12724,N_12590);
xnor U12844 (N_12844,N_12639,N_12704);
nor U12845 (N_12845,N_12553,N_12734);
nand U12846 (N_12846,N_12606,N_12594);
or U12847 (N_12847,N_12616,N_12636);
nand U12848 (N_12848,N_12681,N_12720);
and U12849 (N_12849,N_12646,N_12517);
and U12850 (N_12850,N_12674,N_12651);
or U12851 (N_12851,N_12635,N_12564);
or U12852 (N_12852,N_12591,N_12660);
xnor U12853 (N_12853,N_12718,N_12516);
and U12854 (N_12854,N_12601,N_12747);
and U12855 (N_12855,N_12739,N_12599);
or U12856 (N_12856,N_12723,N_12515);
nand U12857 (N_12857,N_12556,N_12663);
xor U12858 (N_12858,N_12552,N_12549);
and U12859 (N_12859,N_12524,N_12576);
nor U12860 (N_12860,N_12667,N_12520);
or U12861 (N_12861,N_12666,N_12571);
nand U12862 (N_12862,N_12654,N_12596);
xnor U12863 (N_12863,N_12743,N_12621);
nand U12864 (N_12864,N_12693,N_12735);
nand U12865 (N_12865,N_12671,N_12748);
or U12866 (N_12866,N_12610,N_12627);
and U12867 (N_12867,N_12521,N_12676);
nand U12868 (N_12868,N_12626,N_12715);
or U12869 (N_12869,N_12707,N_12579);
or U12870 (N_12870,N_12615,N_12522);
nor U12871 (N_12871,N_12509,N_12699);
nand U12872 (N_12872,N_12736,N_12565);
and U12873 (N_12873,N_12617,N_12652);
nand U12874 (N_12874,N_12560,N_12637);
nand U12875 (N_12875,N_12643,N_12662);
nand U12876 (N_12876,N_12643,N_12519);
or U12877 (N_12877,N_12513,N_12541);
nand U12878 (N_12878,N_12540,N_12503);
or U12879 (N_12879,N_12651,N_12536);
nor U12880 (N_12880,N_12651,N_12518);
nor U12881 (N_12881,N_12547,N_12724);
or U12882 (N_12882,N_12736,N_12503);
xnor U12883 (N_12883,N_12635,N_12672);
or U12884 (N_12884,N_12661,N_12692);
nor U12885 (N_12885,N_12738,N_12521);
nor U12886 (N_12886,N_12688,N_12637);
and U12887 (N_12887,N_12564,N_12731);
nand U12888 (N_12888,N_12734,N_12629);
nand U12889 (N_12889,N_12555,N_12521);
nand U12890 (N_12890,N_12716,N_12705);
nand U12891 (N_12891,N_12600,N_12512);
nor U12892 (N_12892,N_12742,N_12721);
and U12893 (N_12893,N_12573,N_12697);
xor U12894 (N_12894,N_12631,N_12593);
or U12895 (N_12895,N_12692,N_12545);
nor U12896 (N_12896,N_12502,N_12536);
or U12897 (N_12897,N_12602,N_12721);
or U12898 (N_12898,N_12539,N_12545);
nor U12899 (N_12899,N_12656,N_12646);
or U12900 (N_12900,N_12635,N_12671);
and U12901 (N_12901,N_12733,N_12666);
xor U12902 (N_12902,N_12656,N_12673);
nor U12903 (N_12903,N_12650,N_12742);
nor U12904 (N_12904,N_12624,N_12707);
or U12905 (N_12905,N_12555,N_12680);
nand U12906 (N_12906,N_12704,N_12619);
or U12907 (N_12907,N_12707,N_12721);
or U12908 (N_12908,N_12535,N_12639);
and U12909 (N_12909,N_12742,N_12581);
or U12910 (N_12910,N_12657,N_12680);
and U12911 (N_12911,N_12726,N_12625);
nor U12912 (N_12912,N_12577,N_12560);
or U12913 (N_12913,N_12737,N_12641);
nand U12914 (N_12914,N_12672,N_12655);
or U12915 (N_12915,N_12615,N_12631);
nand U12916 (N_12916,N_12595,N_12718);
and U12917 (N_12917,N_12534,N_12543);
and U12918 (N_12918,N_12572,N_12617);
or U12919 (N_12919,N_12558,N_12722);
nor U12920 (N_12920,N_12632,N_12624);
and U12921 (N_12921,N_12688,N_12740);
and U12922 (N_12922,N_12564,N_12674);
and U12923 (N_12923,N_12733,N_12718);
nand U12924 (N_12924,N_12520,N_12731);
and U12925 (N_12925,N_12546,N_12607);
nand U12926 (N_12926,N_12715,N_12749);
nor U12927 (N_12927,N_12524,N_12657);
or U12928 (N_12928,N_12527,N_12546);
and U12929 (N_12929,N_12580,N_12663);
and U12930 (N_12930,N_12734,N_12645);
or U12931 (N_12931,N_12705,N_12596);
and U12932 (N_12932,N_12733,N_12740);
or U12933 (N_12933,N_12655,N_12605);
nand U12934 (N_12934,N_12552,N_12691);
or U12935 (N_12935,N_12602,N_12665);
nor U12936 (N_12936,N_12627,N_12585);
and U12937 (N_12937,N_12687,N_12606);
nand U12938 (N_12938,N_12699,N_12669);
nor U12939 (N_12939,N_12578,N_12736);
xnor U12940 (N_12940,N_12553,N_12545);
or U12941 (N_12941,N_12521,N_12662);
nand U12942 (N_12942,N_12658,N_12513);
nor U12943 (N_12943,N_12668,N_12511);
nor U12944 (N_12944,N_12609,N_12670);
nor U12945 (N_12945,N_12669,N_12585);
and U12946 (N_12946,N_12696,N_12608);
nand U12947 (N_12947,N_12558,N_12601);
or U12948 (N_12948,N_12715,N_12638);
nor U12949 (N_12949,N_12640,N_12692);
nor U12950 (N_12950,N_12683,N_12696);
or U12951 (N_12951,N_12740,N_12704);
or U12952 (N_12952,N_12705,N_12641);
and U12953 (N_12953,N_12673,N_12508);
and U12954 (N_12954,N_12712,N_12741);
nor U12955 (N_12955,N_12600,N_12670);
or U12956 (N_12956,N_12649,N_12567);
xnor U12957 (N_12957,N_12567,N_12610);
nand U12958 (N_12958,N_12707,N_12606);
nand U12959 (N_12959,N_12704,N_12587);
and U12960 (N_12960,N_12583,N_12701);
nor U12961 (N_12961,N_12502,N_12678);
or U12962 (N_12962,N_12701,N_12570);
nor U12963 (N_12963,N_12743,N_12558);
or U12964 (N_12964,N_12625,N_12545);
nand U12965 (N_12965,N_12558,N_12553);
nand U12966 (N_12966,N_12646,N_12527);
and U12967 (N_12967,N_12731,N_12515);
nor U12968 (N_12968,N_12550,N_12603);
xnor U12969 (N_12969,N_12727,N_12680);
or U12970 (N_12970,N_12559,N_12720);
nand U12971 (N_12971,N_12743,N_12613);
or U12972 (N_12972,N_12531,N_12576);
or U12973 (N_12973,N_12650,N_12701);
and U12974 (N_12974,N_12656,N_12545);
or U12975 (N_12975,N_12620,N_12562);
and U12976 (N_12976,N_12648,N_12543);
and U12977 (N_12977,N_12522,N_12681);
or U12978 (N_12978,N_12550,N_12636);
nand U12979 (N_12979,N_12647,N_12507);
xor U12980 (N_12980,N_12692,N_12557);
and U12981 (N_12981,N_12574,N_12700);
and U12982 (N_12982,N_12573,N_12643);
or U12983 (N_12983,N_12654,N_12653);
nor U12984 (N_12984,N_12589,N_12642);
and U12985 (N_12985,N_12692,N_12674);
nand U12986 (N_12986,N_12735,N_12694);
and U12987 (N_12987,N_12656,N_12563);
nor U12988 (N_12988,N_12584,N_12749);
nand U12989 (N_12989,N_12524,N_12541);
nand U12990 (N_12990,N_12723,N_12680);
or U12991 (N_12991,N_12739,N_12616);
nor U12992 (N_12992,N_12521,N_12731);
nor U12993 (N_12993,N_12554,N_12718);
and U12994 (N_12994,N_12725,N_12517);
xnor U12995 (N_12995,N_12681,N_12742);
and U12996 (N_12996,N_12543,N_12502);
xor U12997 (N_12997,N_12592,N_12738);
or U12998 (N_12998,N_12543,N_12569);
xor U12999 (N_12999,N_12712,N_12665);
and U13000 (N_13000,N_12776,N_12910);
or U13001 (N_13001,N_12969,N_12835);
and U13002 (N_13002,N_12811,N_12925);
and U13003 (N_13003,N_12764,N_12853);
nand U13004 (N_13004,N_12894,N_12859);
and U13005 (N_13005,N_12887,N_12826);
nor U13006 (N_13006,N_12768,N_12911);
nor U13007 (N_13007,N_12822,N_12815);
or U13008 (N_13008,N_12947,N_12921);
xnor U13009 (N_13009,N_12818,N_12990);
nor U13010 (N_13010,N_12861,N_12760);
nand U13011 (N_13011,N_12769,N_12888);
and U13012 (N_13012,N_12812,N_12903);
nand U13013 (N_13013,N_12880,N_12941);
xnor U13014 (N_13014,N_12908,N_12875);
xnor U13015 (N_13015,N_12985,N_12851);
nor U13016 (N_13016,N_12895,N_12789);
xor U13017 (N_13017,N_12898,N_12839);
or U13018 (N_13018,N_12899,N_12936);
and U13019 (N_13019,N_12977,N_12772);
or U13020 (N_13020,N_12750,N_12961);
nor U13021 (N_13021,N_12962,N_12943);
nor U13022 (N_13022,N_12945,N_12785);
xnor U13023 (N_13023,N_12967,N_12868);
nand U13024 (N_13024,N_12890,N_12916);
and U13025 (N_13025,N_12753,N_12993);
nand U13026 (N_13026,N_12992,N_12968);
nand U13027 (N_13027,N_12850,N_12854);
or U13028 (N_13028,N_12855,N_12847);
nor U13029 (N_13029,N_12809,N_12821);
nand U13030 (N_13030,N_12758,N_12844);
and U13031 (N_13031,N_12950,N_12877);
and U13032 (N_13032,N_12796,N_12782);
nand U13033 (N_13033,N_12765,N_12838);
or U13034 (N_13034,N_12814,N_12960);
nand U13035 (N_13035,N_12884,N_12813);
or U13036 (N_13036,N_12841,N_12865);
nand U13037 (N_13037,N_12801,N_12878);
nand U13038 (N_13038,N_12879,N_12805);
nand U13039 (N_13039,N_12933,N_12923);
and U13040 (N_13040,N_12998,N_12840);
nor U13041 (N_13041,N_12790,N_12931);
and U13042 (N_13042,N_12832,N_12901);
or U13043 (N_13043,N_12792,N_12966);
or U13044 (N_13044,N_12797,N_12869);
nor U13045 (N_13045,N_12775,N_12779);
nand U13046 (N_13046,N_12783,N_12852);
or U13047 (N_13047,N_12824,N_12981);
nor U13048 (N_13048,N_12795,N_12873);
nor U13049 (N_13049,N_12843,N_12994);
nand U13050 (N_13050,N_12807,N_12808);
nor U13051 (N_13051,N_12823,N_12800);
or U13052 (N_13052,N_12949,N_12924);
or U13053 (N_13053,N_12876,N_12829);
or U13054 (N_13054,N_12964,N_12781);
or U13055 (N_13055,N_12846,N_12928);
and U13056 (N_13056,N_12777,N_12870);
nor U13057 (N_13057,N_12897,N_12940);
and U13058 (N_13058,N_12885,N_12918);
nand U13059 (N_13059,N_12794,N_12778);
nand U13060 (N_13060,N_12770,N_12944);
nand U13061 (N_13061,N_12893,N_12817);
xor U13062 (N_13062,N_12751,N_12984);
nand U13063 (N_13063,N_12942,N_12787);
nor U13064 (N_13064,N_12939,N_12988);
nor U13065 (N_13065,N_12834,N_12881);
nor U13066 (N_13066,N_12905,N_12827);
nor U13067 (N_13067,N_12935,N_12799);
and U13068 (N_13068,N_12788,N_12804);
and U13069 (N_13069,N_12874,N_12973);
nand U13070 (N_13070,N_12803,N_12934);
nor U13071 (N_13071,N_12991,N_12932);
or U13072 (N_13072,N_12957,N_12970);
or U13073 (N_13073,N_12983,N_12907);
xor U13074 (N_13074,N_12997,N_12915);
nor U13075 (N_13075,N_12909,N_12784);
or U13076 (N_13076,N_12906,N_12856);
nand U13077 (N_13077,N_12857,N_12989);
or U13078 (N_13078,N_12946,N_12761);
and U13079 (N_13079,N_12948,N_12980);
or U13080 (N_13080,N_12987,N_12974);
nand U13081 (N_13081,N_12902,N_12979);
nor U13082 (N_13082,N_12871,N_12848);
and U13083 (N_13083,N_12978,N_12845);
xnor U13084 (N_13084,N_12842,N_12767);
or U13085 (N_13085,N_12922,N_12959);
nand U13086 (N_13086,N_12972,N_12791);
nor U13087 (N_13087,N_12867,N_12900);
nor U13088 (N_13088,N_12927,N_12913);
nand U13089 (N_13089,N_12820,N_12786);
and U13090 (N_13090,N_12830,N_12810);
nand U13091 (N_13091,N_12938,N_12862);
nand U13092 (N_13092,N_12866,N_12951);
xnor U13093 (N_13093,N_12889,N_12757);
or U13094 (N_13094,N_12917,N_12763);
nand U13095 (N_13095,N_12920,N_12860);
and U13096 (N_13096,N_12774,N_12955);
or U13097 (N_13097,N_12912,N_12816);
or U13098 (N_13098,N_12971,N_12752);
nand U13099 (N_13099,N_12793,N_12996);
and U13100 (N_13100,N_12836,N_12891);
nand U13101 (N_13101,N_12864,N_12780);
xnor U13102 (N_13102,N_12937,N_12956);
or U13103 (N_13103,N_12802,N_12896);
xor U13104 (N_13104,N_12766,N_12952);
nand U13105 (N_13105,N_12849,N_12883);
and U13106 (N_13106,N_12958,N_12754);
nand U13107 (N_13107,N_12919,N_12954);
or U13108 (N_13108,N_12975,N_12756);
nand U13109 (N_13109,N_12882,N_12771);
nor U13110 (N_13110,N_12819,N_12762);
or U13111 (N_13111,N_12892,N_12837);
xor U13112 (N_13112,N_12825,N_12953);
xor U13113 (N_13113,N_12904,N_12963);
or U13114 (N_13114,N_12986,N_12798);
nand U13115 (N_13115,N_12930,N_12858);
and U13116 (N_13116,N_12886,N_12759);
nand U13117 (N_13117,N_12806,N_12926);
nor U13118 (N_13118,N_12982,N_12872);
and U13119 (N_13119,N_12773,N_12965);
nor U13120 (N_13120,N_12833,N_12999);
and U13121 (N_13121,N_12828,N_12863);
nor U13122 (N_13122,N_12755,N_12929);
or U13123 (N_13123,N_12914,N_12831);
and U13124 (N_13124,N_12976,N_12995);
nand U13125 (N_13125,N_12900,N_12766);
nand U13126 (N_13126,N_12820,N_12769);
or U13127 (N_13127,N_12755,N_12771);
and U13128 (N_13128,N_12775,N_12871);
xor U13129 (N_13129,N_12935,N_12947);
or U13130 (N_13130,N_12922,N_12810);
nand U13131 (N_13131,N_12804,N_12819);
or U13132 (N_13132,N_12977,N_12995);
and U13133 (N_13133,N_12759,N_12807);
nand U13134 (N_13134,N_12788,N_12935);
and U13135 (N_13135,N_12835,N_12820);
or U13136 (N_13136,N_12851,N_12961);
nor U13137 (N_13137,N_12885,N_12974);
or U13138 (N_13138,N_12764,N_12977);
xnor U13139 (N_13139,N_12842,N_12952);
and U13140 (N_13140,N_12930,N_12937);
nor U13141 (N_13141,N_12959,N_12967);
nand U13142 (N_13142,N_12788,N_12876);
nor U13143 (N_13143,N_12907,N_12942);
nor U13144 (N_13144,N_12803,N_12988);
or U13145 (N_13145,N_12836,N_12757);
and U13146 (N_13146,N_12900,N_12998);
nand U13147 (N_13147,N_12905,N_12856);
or U13148 (N_13148,N_12890,N_12983);
nor U13149 (N_13149,N_12958,N_12826);
or U13150 (N_13150,N_12907,N_12812);
nor U13151 (N_13151,N_12841,N_12839);
or U13152 (N_13152,N_12940,N_12955);
and U13153 (N_13153,N_12883,N_12886);
nand U13154 (N_13154,N_12995,N_12982);
or U13155 (N_13155,N_12971,N_12952);
nand U13156 (N_13156,N_12867,N_12909);
nand U13157 (N_13157,N_12903,N_12932);
or U13158 (N_13158,N_12921,N_12899);
or U13159 (N_13159,N_12797,N_12987);
nand U13160 (N_13160,N_12897,N_12853);
nor U13161 (N_13161,N_12899,N_12783);
or U13162 (N_13162,N_12895,N_12941);
and U13163 (N_13163,N_12815,N_12881);
and U13164 (N_13164,N_12849,N_12894);
nor U13165 (N_13165,N_12911,N_12904);
or U13166 (N_13166,N_12839,N_12884);
nor U13167 (N_13167,N_12828,N_12879);
nand U13168 (N_13168,N_12981,N_12949);
or U13169 (N_13169,N_12927,N_12876);
or U13170 (N_13170,N_12905,N_12765);
or U13171 (N_13171,N_12814,N_12926);
and U13172 (N_13172,N_12858,N_12789);
or U13173 (N_13173,N_12912,N_12937);
or U13174 (N_13174,N_12809,N_12991);
nand U13175 (N_13175,N_12814,N_12923);
and U13176 (N_13176,N_12828,N_12860);
nor U13177 (N_13177,N_12769,N_12761);
or U13178 (N_13178,N_12936,N_12874);
or U13179 (N_13179,N_12853,N_12797);
nand U13180 (N_13180,N_12861,N_12944);
and U13181 (N_13181,N_12868,N_12851);
nor U13182 (N_13182,N_12881,N_12922);
and U13183 (N_13183,N_12829,N_12796);
or U13184 (N_13184,N_12798,N_12865);
nand U13185 (N_13185,N_12822,N_12817);
nor U13186 (N_13186,N_12829,N_12793);
and U13187 (N_13187,N_12898,N_12998);
or U13188 (N_13188,N_12949,N_12790);
nand U13189 (N_13189,N_12929,N_12840);
nand U13190 (N_13190,N_12893,N_12825);
nor U13191 (N_13191,N_12857,N_12933);
nor U13192 (N_13192,N_12905,N_12926);
and U13193 (N_13193,N_12920,N_12955);
nor U13194 (N_13194,N_12926,N_12767);
xnor U13195 (N_13195,N_12864,N_12869);
or U13196 (N_13196,N_12989,N_12921);
and U13197 (N_13197,N_12905,N_12833);
nor U13198 (N_13198,N_12941,N_12772);
nor U13199 (N_13199,N_12808,N_12754);
xor U13200 (N_13200,N_12861,N_12899);
or U13201 (N_13201,N_12850,N_12768);
nand U13202 (N_13202,N_12841,N_12858);
nor U13203 (N_13203,N_12803,N_12946);
or U13204 (N_13204,N_12964,N_12896);
or U13205 (N_13205,N_12896,N_12918);
xor U13206 (N_13206,N_12890,N_12860);
xor U13207 (N_13207,N_12809,N_12945);
nand U13208 (N_13208,N_12984,N_12762);
nor U13209 (N_13209,N_12972,N_12954);
and U13210 (N_13210,N_12884,N_12988);
nand U13211 (N_13211,N_12784,N_12875);
or U13212 (N_13212,N_12866,N_12898);
nand U13213 (N_13213,N_12862,N_12934);
nor U13214 (N_13214,N_12824,N_12994);
and U13215 (N_13215,N_12750,N_12966);
or U13216 (N_13216,N_12899,N_12805);
and U13217 (N_13217,N_12997,N_12903);
or U13218 (N_13218,N_12995,N_12974);
or U13219 (N_13219,N_12878,N_12960);
nand U13220 (N_13220,N_12799,N_12987);
nor U13221 (N_13221,N_12809,N_12953);
and U13222 (N_13222,N_12901,N_12857);
and U13223 (N_13223,N_12939,N_12825);
nor U13224 (N_13224,N_12875,N_12939);
xor U13225 (N_13225,N_12767,N_12850);
nor U13226 (N_13226,N_12892,N_12753);
and U13227 (N_13227,N_12810,N_12822);
and U13228 (N_13228,N_12869,N_12872);
or U13229 (N_13229,N_12843,N_12906);
nor U13230 (N_13230,N_12973,N_12862);
nor U13231 (N_13231,N_12796,N_12895);
or U13232 (N_13232,N_12979,N_12930);
nor U13233 (N_13233,N_12886,N_12979);
nand U13234 (N_13234,N_12975,N_12871);
or U13235 (N_13235,N_12963,N_12792);
and U13236 (N_13236,N_12805,N_12814);
and U13237 (N_13237,N_12975,N_12773);
nor U13238 (N_13238,N_12989,N_12907);
and U13239 (N_13239,N_12819,N_12922);
nand U13240 (N_13240,N_12830,N_12993);
and U13241 (N_13241,N_12979,N_12919);
or U13242 (N_13242,N_12900,N_12966);
nand U13243 (N_13243,N_12813,N_12756);
nor U13244 (N_13244,N_12753,N_12821);
nor U13245 (N_13245,N_12925,N_12877);
and U13246 (N_13246,N_12929,N_12827);
and U13247 (N_13247,N_12903,N_12794);
or U13248 (N_13248,N_12790,N_12832);
or U13249 (N_13249,N_12906,N_12822);
nor U13250 (N_13250,N_13012,N_13022);
nor U13251 (N_13251,N_13061,N_13093);
nor U13252 (N_13252,N_13241,N_13117);
nor U13253 (N_13253,N_13208,N_13226);
nor U13254 (N_13254,N_13115,N_13206);
nand U13255 (N_13255,N_13196,N_13045);
nor U13256 (N_13256,N_13192,N_13182);
nor U13257 (N_13257,N_13205,N_13167);
and U13258 (N_13258,N_13214,N_13216);
and U13259 (N_13259,N_13212,N_13028);
or U13260 (N_13260,N_13126,N_13018);
nand U13261 (N_13261,N_13002,N_13131);
nor U13262 (N_13262,N_13148,N_13005);
nor U13263 (N_13263,N_13073,N_13238);
or U13264 (N_13264,N_13137,N_13118);
and U13265 (N_13265,N_13019,N_13043);
xor U13266 (N_13266,N_13079,N_13114);
nand U13267 (N_13267,N_13049,N_13047);
nand U13268 (N_13268,N_13020,N_13229);
and U13269 (N_13269,N_13149,N_13199);
and U13270 (N_13270,N_13165,N_13158);
or U13271 (N_13271,N_13111,N_13071);
and U13272 (N_13272,N_13039,N_13136);
xor U13273 (N_13273,N_13072,N_13219);
xor U13274 (N_13274,N_13036,N_13188);
or U13275 (N_13275,N_13105,N_13098);
xnor U13276 (N_13276,N_13135,N_13198);
and U13277 (N_13277,N_13184,N_13175);
and U13278 (N_13278,N_13017,N_13203);
and U13279 (N_13279,N_13178,N_13223);
or U13280 (N_13280,N_13001,N_13121);
or U13281 (N_13281,N_13142,N_13101);
nor U13282 (N_13282,N_13075,N_13247);
and U13283 (N_13283,N_13202,N_13038);
nor U13284 (N_13284,N_13180,N_13228);
nand U13285 (N_13285,N_13147,N_13130);
or U13286 (N_13286,N_13164,N_13086);
nand U13287 (N_13287,N_13236,N_13094);
and U13288 (N_13288,N_13222,N_13050);
and U13289 (N_13289,N_13032,N_13225);
nand U13290 (N_13290,N_13194,N_13024);
nor U13291 (N_13291,N_13051,N_13080);
or U13292 (N_13292,N_13227,N_13240);
or U13293 (N_13293,N_13059,N_13161);
nand U13294 (N_13294,N_13186,N_13044);
and U13295 (N_13295,N_13144,N_13189);
nor U13296 (N_13296,N_13168,N_13084);
and U13297 (N_13297,N_13100,N_13204);
nor U13298 (N_13298,N_13154,N_13174);
or U13299 (N_13299,N_13119,N_13006);
or U13300 (N_13300,N_13244,N_13143);
and U13301 (N_13301,N_13155,N_13081);
or U13302 (N_13302,N_13058,N_13245);
nor U13303 (N_13303,N_13095,N_13070);
xor U13304 (N_13304,N_13000,N_13063);
nand U13305 (N_13305,N_13069,N_13067);
and U13306 (N_13306,N_13140,N_13060);
and U13307 (N_13307,N_13097,N_13128);
xnor U13308 (N_13308,N_13132,N_13087);
xor U13309 (N_13309,N_13220,N_13108);
and U13310 (N_13310,N_13150,N_13023);
nand U13311 (N_13311,N_13146,N_13190);
and U13312 (N_13312,N_13195,N_13153);
or U13313 (N_13313,N_13052,N_13089);
nor U13314 (N_13314,N_13215,N_13109);
nor U13315 (N_13315,N_13177,N_13056);
nand U13316 (N_13316,N_13159,N_13090);
nand U13317 (N_13317,N_13003,N_13179);
and U13318 (N_13318,N_13207,N_13242);
nor U13319 (N_13319,N_13096,N_13091);
xor U13320 (N_13320,N_13173,N_13152);
and U13321 (N_13321,N_13011,N_13110);
and U13322 (N_13322,N_13124,N_13027);
or U13323 (N_13323,N_13112,N_13014);
nor U13324 (N_13324,N_13104,N_13004);
nand U13325 (N_13325,N_13123,N_13034);
nand U13326 (N_13326,N_13145,N_13120);
and U13327 (N_13327,N_13221,N_13016);
nand U13328 (N_13328,N_13193,N_13156);
nor U13329 (N_13329,N_13054,N_13026);
nand U13330 (N_13330,N_13127,N_13107);
nor U13331 (N_13331,N_13055,N_13138);
or U13332 (N_13332,N_13009,N_13239);
or U13333 (N_13333,N_13064,N_13134);
nand U13334 (N_13334,N_13077,N_13106);
nor U13335 (N_13335,N_13197,N_13224);
and U13336 (N_13336,N_13187,N_13243);
and U13337 (N_13337,N_13041,N_13213);
nor U13338 (N_13338,N_13113,N_13170);
nor U13339 (N_13339,N_13157,N_13230);
nor U13340 (N_13340,N_13025,N_13076);
and U13341 (N_13341,N_13040,N_13141);
or U13342 (N_13342,N_13037,N_13169);
nand U13343 (N_13343,N_13068,N_13013);
nor U13344 (N_13344,N_13234,N_13172);
nor U13345 (N_13345,N_13035,N_13066);
nand U13346 (N_13346,N_13031,N_13092);
and U13347 (N_13347,N_13166,N_13085);
nor U13348 (N_13348,N_13176,N_13053);
and U13349 (N_13349,N_13209,N_13102);
nand U13350 (N_13350,N_13122,N_13232);
or U13351 (N_13351,N_13181,N_13218);
or U13352 (N_13352,N_13249,N_13160);
or U13353 (N_13353,N_13030,N_13033);
nor U13354 (N_13354,N_13008,N_13231);
nor U13355 (N_13355,N_13103,N_13201);
and U13356 (N_13356,N_13099,N_13139);
and U13357 (N_13357,N_13183,N_13133);
nor U13358 (N_13358,N_13083,N_13233);
or U13359 (N_13359,N_13129,N_13074);
or U13360 (N_13360,N_13057,N_13235);
nand U13361 (N_13361,N_13151,N_13042);
nor U13362 (N_13362,N_13210,N_13237);
nor U13363 (N_13363,N_13211,N_13163);
nor U13364 (N_13364,N_13046,N_13116);
nand U13365 (N_13365,N_13021,N_13065);
nand U13366 (N_13366,N_13246,N_13171);
and U13367 (N_13367,N_13015,N_13029);
xnor U13368 (N_13368,N_13185,N_13088);
nand U13369 (N_13369,N_13082,N_13062);
and U13370 (N_13370,N_13078,N_13217);
or U13371 (N_13371,N_13191,N_13125);
nor U13372 (N_13372,N_13248,N_13162);
nor U13373 (N_13373,N_13200,N_13048);
nor U13374 (N_13374,N_13010,N_13007);
nor U13375 (N_13375,N_13080,N_13058);
and U13376 (N_13376,N_13064,N_13244);
and U13377 (N_13377,N_13087,N_13029);
xor U13378 (N_13378,N_13034,N_13074);
and U13379 (N_13379,N_13132,N_13114);
and U13380 (N_13380,N_13014,N_13000);
nand U13381 (N_13381,N_13055,N_13040);
or U13382 (N_13382,N_13239,N_13005);
xor U13383 (N_13383,N_13065,N_13081);
nand U13384 (N_13384,N_13120,N_13038);
or U13385 (N_13385,N_13229,N_13022);
nand U13386 (N_13386,N_13089,N_13137);
xnor U13387 (N_13387,N_13181,N_13135);
or U13388 (N_13388,N_13058,N_13011);
nand U13389 (N_13389,N_13228,N_13076);
nand U13390 (N_13390,N_13077,N_13083);
nor U13391 (N_13391,N_13057,N_13062);
nor U13392 (N_13392,N_13049,N_13019);
nor U13393 (N_13393,N_13191,N_13176);
and U13394 (N_13394,N_13147,N_13206);
or U13395 (N_13395,N_13043,N_13187);
nand U13396 (N_13396,N_13137,N_13106);
nand U13397 (N_13397,N_13137,N_13156);
and U13398 (N_13398,N_13248,N_13136);
and U13399 (N_13399,N_13087,N_13092);
nor U13400 (N_13400,N_13161,N_13112);
nor U13401 (N_13401,N_13097,N_13244);
and U13402 (N_13402,N_13205,N_13233);
nor U13403 (N_13403,N_13240,N_13036);
and U13404 (N_13404,N_13132,N_13017);
or U13405 (N_13405,N_13110,N_13159);
or U13406 (N_13406,N_13209,N_13110);
or U13407 (N_13407,N_13048,N_13234);
and U13408 (N_13408,N_13071,N_13196);
and U13409 (N_13409,N_13031,N_13185);
and U13410 (N_13410,N_13240,N_13082);
xnor U13411 (N_13411,N_13206,N_13065);
or U13412 (N_13412,N_13148,N_13004);
nand U13413 (N_13413,N_13021,N_13198);
nand U13414 (N_13414,N_13207,N_13133);
and U13415 (N_13415,N_13197,N_13179);
and U13416 (N_13416,N_13059,N_13234);
nor U13417 (N_13417,N_13068,N_13153);
and U13418 (N_13418,N_13072,N_13129);
or U13419 (N_13419,N_13069,N_13092);
nand U13420 (N_13420,N_13011,N_13017);
nor U13421 (N_13421,N_13129,N_13037);
nor U13422 (N_13422,N_13212,N_13050);
nor U13423 (N_13423,N_13011,N_13160);
and U13424 (N_13424,N_13079,N_13186);
or U13425 (N_13425,N_13043,N_13227);
and U13426 (N_13426,N_13010,N_13116);
nand U13427 (N_13427,N_13233,N_13012);
nand U13428 (N_13428,N_13117,N_13160);
xnor U13429 (N_13429,N_13160,N_13015);
and U13430 (N_13430,N_13115,N_13089);
and U13431 (N_13431,N_13141,N_13204);
xnor U13432 (N_13432,N_13100,N_13195);
xor U13433 (N_13433,N_13239,N_13102);
nand U13434 (N_13434,N_13054,N_13044);
nor U13435 (N_13435,N_13210,N_13155);
or U13436 (N_13436,N_13129,N_13184);
and U13437 (N_13437,N_13017,N_13040);
nand U13438 (N_13438,N_13208,N_13136);
or U13439 (N_13439,N_13095,N_13127);
and U13440 (N_13440,N_13138,N_13146);
nand U13441 (N_13441,N_13143,N_13243);
or U13442 (N_13442,N_13084,N_13093);
or U13443 (N_13443,N_13201,N_13007);
nand U13444 (N_13444,N_13202,N_13163);
nand U13445 (N_13445,N_13232,N_13091);
or U13446 (N_13446,N_13087,N_13188);
nand U13447 (N_13447,N_13143,N_13148);
nand U13448 (N_13448,N_13127,N_13152);
or U13449 (N_13449,N_13128,N_13063);
nand U13450 (N_13450,N_13143,N_13242);
xnor U13451 (N_13451,N_13045,N_13131);
nor U13452 (N_13452,N_13172,N_13027);
nand U13453 (N_13453,N_13108,N_13206);
and U13454 (N_13454,N_13054,N_13063);
xor U13455 (N_13455,N_13225,N_13050);
and U13456 (N_13456,N_13009,N_13246);
or U13457 (N_13457,N_13007,N_13159);
nand U13458 (N_13458,N_13124,N_13079);
nand U13459 (N_13459,N_13011,N_13153);
nor U13460 (N_13460,N_13103,N_13165);
nor U13461 (N_13461,N_13018,N_13174);
nor U13462 (N_13462,N_13102,N_13226);
or U13463 (N_13463,N_13187,N_13091);
or U13464 (N_13464,N_13095,N_13040);
or U13465 (N_13465,N_13023,N_13224);
nor U13466 (N_13466,N_13212,N_13033);
and U13467 (N_13467,N_13240,N_13160);
and U13468 (N_13468,N_13053,N_13064);
nand U13469 (N_13469,N_13107,N_13070);
or U13470 (N_13470,N_13015,N_13040);
nand U13471 (N_13471,N_13144,N_13187);
and U13472 (N_13472,N_13147,N_13020);
or U13473 (N_13473,N_13213,N_13110);
nor U13474 (N_13474,N_13062,N_13118);
or U13475 (N_13475,N_13206,N_13157);
nand U13476 (N_13476,N_13239,N_13190);
nand U13477 (N_13477,N_13243,N_13000);
nor U13478 (N_13478,N_13011,N_13027);
nor U13479 (N_13479,N_13194,N_13014);
or U13480 (N_13480,N_13170,N_13242);
nor U13481 (N_13481,N_13068,N_13239);
or U13482 (N_13482,N_13195,N_13048);
nand U13483 (N_13483,N_13111,N_13035);
nor U13484 (N_13484,N_13064,N_13160);
and U13485 (N_13485,N_13122,N_13024);
nand U13486 (N_13486,N_13005,N_13164);
nand U13487 (N_13487,N_13241,N_13193);
nor U13488 (N_13488,N_13211,N_13147);
nor U13489 (N_13489,N_13228,N_13241);
xor U13490 (N_13490,N_13140,N_13184);
and U13491 (N_13491,N_13049,N_13121);
nor U13492 (N_13492,N_13031,N_13117);
xor U13493 (N_13493,N_13243,N_13207);
and U13494 (N_13494,N_13131,N_13146);
and U13495 (N_13495,N_13069,N_13103);
nand U13496 (N_13496,N_13191,N_13198);
nand U13497 (N_13497,N_13145,N_13112);
or U13498 (N_13498,N_13223,N_13150);
and U13499 (N_13499,N_13157,N_13190);
or U13500 (N_13500,N_13439,N_13350);
nand U13501 (N_13501,N_13295,N_13473);
or U13502 (N_13502,N_13395,N_13352);
and U13503 (N_13503,N_13337,N_13406);
nor U13504 (N_13504,N_13388,N_13267);
and U13505 (N_13505,N_13289,N_13357);
nand U13506 (N_13506,N_13292,N_13476);
nor U13507 (N_13507,N_13447,N_13259);
and U13508 (N_13508,N_13396,N_13417);
xnor U13509 (N_13509,N_13260,N_13347);
or U13510 (N_13510,N_13392,N_13252);
or U13511 (N_13511,N_13302,N_13270);
nor U13512 (N_13512,N_13366,N_13264);
or U13513 (N_13513,N_13485,N_13311);
or U13514 (N_13514,N_13462,N_13477);
or U13515 (N_13515,N_13428,N_13420);
and U13516 (N_13516,N_13414,N_13367);
xnor U13517 (N_13517,N_13467,N_13436);
or U13518 (N_13518,N_13387,N_13391);
and U13519 (N_13519,N_13271,N_13361);
and U13520 (N_13520,N_13360,N_13442);
or U13521 (N_13521,N_13374,N_13318);
or U13522 (N_13522,N_13268,N_13433);
xnor U13523 (N_13523,N_13489,N_13445);
and U13524 (N_13524,N_13272,N_13369);
xor U13525 (N_13525,N_13384,N_13338);
or U13526 (N_13526,N_13342,N_13487);
nor U13527 (N_13527,N_13326,N_13349);
and U13528 (N_13528,N_13483,N_13315);
nor U13529 (N_13529,N_13362,N_13278);
nand U13530 (N_13530,N_13498,N_13423);
and U13531 (N_13531,N_13339,N_13340);
nand U13532 (N_13532,N_13280,N_13474);
nor U13533 (N_13533,N_13364,N_13418);
or U13534 (N_13534,N_13377,N_13261);
or U13535 (N_13535,N_13307,N_13468);
nor U13536 (N_13536,N_13408,N_13425);
nand U13537 (N_13537,N_13312,N_13263);
and U13538 (N_13538,N_13275,N_13372);
nand U13539 (N_13539,N_13375,N_13328);
or U13540 (N_13540,N_13457,N_13290);
nand U13541 (N_13541,N_13276,N_13293);
and U13542 (N_13542,N_13303,N_13454);
or U13543 (N_13543,N_13257,N_13285);
nand U13544 (N_13544,N_13426,N_13334);
nor U13545 (N_13545,N_13385,N_13415);
and U13546 (N_13546,N_13421,N_13472);
nor U13547 (N_13547,N_13262,N_13465);
nor U13548 (N_13548,N_13443,N_13282);
or U13549 (N_13549,N_13363,N_13281);
and U13550 (N_13550,N_13359,N_13351);
xor U13551 (N_13551,N_13284,N_13441);
or U13552 (N_13552,N_13298,N_13460);
nand U13553 (N_13553,N_13410,N_13258);
xor U13554 (N_13554,N_13304,N_13386);
and U13555 (N_13555,N_13399,N_13481);
or U13556 (N_13556,N_13383,N_13305);
nor U13557 (N_13557,N_13435,N_13355);
or U13558 (N_13558,N_13309,N_13286);
nor U13559 (N_13559,N_13389,N_13480);
nor U13560 (N_13560,N_13308,N_13354);
or U13561 (N_13561,N_13493,N_13291);
nand U13562 (N_13562,N_13411,N_13409);
or U13563 (N_13563,N_13310,N_13331);
or U13564 (N_13564,N_13440,N_13373);
xnor U13565 (N_13565,N_13322,N_13346);
nand U13566 (N_13566,N_13356,N_13496);
nand U13567 (N_13567,N_13491,N_13412);
xor U13568 (N_13568,N_13466,N_13452);
nand U13569 (N_13569,N_13314,N_13313);
nand U13570 (N_13570,N_13279,N_13269);
nor U13571 (N_13571,N_13431,N_13494);
or U13572 (N_13572,N_13378,N_13422);
nor U13573 (N_13573,N_13427,N_13458);
nor U13574 (N_13574,N_13482,N_13424);
nor U13575 (N_13575,N_13450,N_13444);
nor U13576 (N_13576,N_13419,N_13459);
and U13577 (N_13577,N_13390,N_13319);
and U13578 (N_13578,N_13393,N_13397);
nor U13579 (N_13579,N_13461,N_13253);
nand U13580 (N_13580,N_13429,N_13353);
xor U13581 (N_13581,N_13336,N_13273);
nand U13582 (N_13582,N_13376,N_13297);
nand U13583 (N_13583,N_13438,N_13495);
or U13584 (N_13584,N_13432,N_13330);
nor U13585 (N_13585,N_13325,N_13402);
xnor U13586 (N_13586,N_13329,N_13327);
and U13587 (N_13587,N_13478,N_13251);
or U13588 (N_13588,N_13451,N_13449);
and U13589 (N_13589,N_13499,N_13324);
nor U13590 (N_13590,N_13341,N_13469);
and U13591 (N_13591,N_13484,N_13437);
and U13592 (N_13592,N_13463,N_13475);
or U13593 (N_13593,N_13358,N_13368);
nand U13594 (N_13594,N_13416,N_13407);
and U13595 (N_13595,N_13323,N_13401);
or U13596 (N_13596,N_13446,N_13371);
xor U13597 (N_13597,N_13380,N_13455);
or U13598 (N_13598,N_13254,N_13497);
or U13599 (N_13599,N_13413,N_13343);
or U13600 (N_13600,N_13296,N_13403);
and U13601 (N_13601,N_13317,N_13382);
and U13602 (N_13602,N_13430,N_13255);
xor U13603 (N_13603,N_13434,N_13488);
nand U13604 (N_13604,N_13365,N_13448);
and U13605 (N_13605,N_13348,N_13277);
and U13606 (N_13606,N_13287,N_13492);
and U13607 (N_13607,N_13266,N_13381);
and U13608 (N_13608,N_13379,N_13265);
xnor U13609 (N_13609,N_13345,N_13394);
or U13610 (N_13610,N_13486,N_13470);
nand U13611 (N_13611,N_13453,N_13274);
xor U13612 (N_13612,N_13344,N_13283);
nor U13613 (N_13613,N_13256,N_13288);
or U13614 (N_13614,N_13335,N_13332);
and U13615 (N_13615,N_13321,N_13316);
nand U13616 (N_13616,N_13301,N_13306);
xor U13617 (N_13617,N_13299,N_13456);
and U13618 (N_13618,N_13490,N_13400);
nor U13619 (N_13619,N_13464,N_13479);
nand U13620 (N_13620,N_13294,N_13250);
xnor U13621 (N_13621,N_13471,N_13320);
nand U13622 (N_13622,N_13333,N_13398);
or U13623 (N_13623,N_13404,N_13370);
and U13624 (N_13624,N_13300,N_13405);
or U13625 (N_13625,N_13417,N_13333);
nor U13626 (N_13626,N_13498,N_13427);
nor U13627 (N_13627,N_13283,N_13497);
or U13628 (N_13628,N_13286,N_13250);
nor U13629 (N_13629,N_13446,N_13409);
nor U13630 (N_13630,N_13291,N_13494);
or U13631 (N_13631,N_13480,N_13447);
nand U13632 (N_13632,N_13387,N_13280);
and U13633 (N_13633,N_13271,N_13442);
nand U13634 (N_13634,N_13276,N_13306);
and U13635 (N_13635,N_13440,N_13313);
and U13636 (N_13636,N_13398,N_13431);
xnor U13637 (N_13637,N_13465,N_13266);
nand U13638 (N_13638,N_13344,N_13336);
or U13639 (N_13639,N_13438,N_13272);
nand U13640 (N_13640,N_13318,N_13358);
and U13641 (N_13641,N_13455,N_13348);
or U13642 (N_13642,N_13281,N_13423);
or U13643 (N_13643,N_13358,N_13392);
nor U13644 (N_13644,N_13429,N_13465);
nor U13645 (N_13645,N_13305,N_13467);
nand U13646 (N_13646,N_13352,N_13279);
and U13647 (N_13647,N_13488,N_13451);
nor U13648 (N_13648,N_13439,N_13291);
nand U13649 (N_13649,N_13282,N_13264);
and U13650 (N_13650,N_13275,N_13365);
xnor U13651 (N_13651,N_13311,N_13375);
nand U13652 (N_13652,N_13327,N_13267);
nand U13653 (N_13653,N_13477,N_13369);
nor U13654 (N_13654,N_13315,N_13378);
xor U13655 (N_13655,N_13307,N_13457);
and U13656 (N_13656,N_13482,N_13383);
xor U13657 (N_13657,N_13379,N_13299);
nand U13658 (N_13658,N_13436,N_13423);
nor U13659 (N_13659,N_13288,N_13275);
or U13660 (N_13660,N_13456,N_13420);
or U13661 (N_13661,N_13317,N_13466);
or U13662 (N_13662,N_13273,N_13407);
and U13663 (N_13663,N_13368,N_13402);
xor U13664 (N_13664,N_13344,N_13368);
xor U13665 (N_13665,N_13462,N_13470);
nand U13666 (N_13666,N_13320,N_13300);
or U13667 (N_13667,N_13425,N_13401);
and U13668 (N_13668,N_13273,N_13305);
nor U13669 (N_13669,N_13265,N_13491);
xnor U13670 (N_13670,N_13390,N_13465);
or U13671 (N_13671,N_13269,N_13409);
or U13672 (N_13672,N_13378,N_13354);
nor U13673 (N_13673,N_13443,N_13392);
and U13674 (N_13674,N_13444,N_13363);
xnor U13675 (N_13675,N_13300,N_13431);
and U13676 (N_13676,N_13265,N_13453);
nor U13677 (N_13677,N_13449,N_13272);
nor U13678 (N_13678,N_13384,N_13322);
and U13679 (N_13679,N_13488,N_13301);
xor U13680 (N_13680,N_13406,N_13484);
or U13681 (N_13681,N_13357,N_13412);
nand U13682 (N_13682,N_13309,N_13388);
nor U13683 (N_13683,N_13493,N_13441);
nor U13684 (N_13684,N_13279,N_13331);
nand U13685 (N_13685,N_13378,N_13294);
or U13686 (N_13686,N_13378,N_13473);
nand U13687 (N_13687,N_13382,N_13295);
nor U13688 (N_13688,N_13282,N_13281);
nand U13689 (N_13689,N_13285,N_13266);
or U13690 (N_13690,N_13461,N_13480);
nor U13691 (N_13691,N_13318,N_13443);
nand U13692 (N_13692,N_13380,N_13383);
and U13693 (N_13693,N_13416,N_13335);
or U13694 (N_13694,N_13324,N_13486);
nand U13695 (N_13695,N_13409,N_13367);
nor U13696 (N_13696,N_13271,N_13334);
xor U13697 (N_13697,N_13351,N_13438);
nor U13698 (N_13698,N_13341,N_13362);
and U13699 (N_13699,N_13388,N_13459);
nand U13700 (N_13700,N_13256,N_13397);
or U13701 (N_13701,N_13259,N_13495);
nor U13702 (N_13702,N_13385,N_13344);
and U13703 (N_13703,N_13468,N_13254);
nand U13704 (N_13704,N_13498,N_13282);
nand U13705 (N_13705,N_13273,N_13347);
nor U13706 (N_13706,N_13270,N_13263);
or U13707 (N_13707,N_13485,N_13359);
xor U13708 (N_13708,N_13387,N_13453);
or U13709 (N_13709,N_13330,N_13402);
or U13710 (N_13710,N_13485,N_13406);
nand U13711 (N_13711,N_13488,N_13269);
or U13712 (N_13712,N_13481,N_13478);
nand U13713 (N_13713,N_13285,N_13271);
nor U13714 (N_13714,N_13315,N_13388);
or U13715 (N_13715,N_13263,N_13388);
nand U13716 (N_13716,N_13445,N_13428);
nand U13717 (N_13717,N_13336,N_13462);
or U13718 (N_13718,N_13472,N_13488);
nand U13719 (N_13719,N_13364,N_13329);
nor U13720 (N_13720,N_13366,N_13337);
nor U13721 (N_13721,N_13458,N_13340);
or U13722 (N_13722,N_13418,N_13432);
nand U13723 (N_13723,N_13403,N_13384);
or U13724 (N_13724,N_13394,N_13315);
and U13725 (N_13725,N_13263,N_13300);
nor U13726 (N_13726,N_13473,N_13369);
and U13727 (N_13727,N_13273,N_13341);
nor U13728 (N_13728,N_13449,N_13408);
nor U13729 (N_13729,N_13425,N_13405);
and U13730 (N_13730,N_13266,N_13313);
nand U13731 (N_13731,N_13317,N_13490);
nor U13732 (N_13732,N_13420,N_13286);
and U13733 (N_13733,N_13250,N_13371);
nand U13734 (N_13734,N_13283,N_13342);
nor U13735 (N_13735,N_13330,N_13410);
nor U13736 (N_13736,N_13326,N_13290);
xnor U13737 (N_13737,N_13267,N_13396);
or U13738 (N_13738,N_13269,N_13357);
xor U13739 (N_13739,N_13328,N_13313);
nor U13740 (N_13740,N_13337,N_13484);
nand U13741 (N_13741,N_13383,N_13362);
or U13742 (N_13742,N_13375,N_13256);
or U13743 (N_13743,N_13319,N_13347);
or U13744 (N_13744,N_13277,N_13473);
nor U13745 (N_13745,N_13250,N_13386);
nand U13746 (N_13746,N_13283,N_13345);
and U13747 (N_13747,N_13479,N_13468);
nor U13748 (N_13748,N_13275,N_13305);
nand U13749 (N_13749,N_13316,N_13440);
xor U13750 (N_13750,N_13504,N_13630);
nand U13751 (N_13751,N_13540,N_13616);
xor U13752 (N_13752,N_13749,N_13727);
nand U13753 (N_13753,N_13605,N_13519);
nor U13754 (N_13754,N_13639,N_13674);
or U13755 (N_13755,N_13649,N_13570);
nor U13756 (N_13756,N_13672,N_13596);
and U13757 (N_13757,N_13664,N_13723);
and U13758 (N_13758,N_13697,N_13594);
nand U13759 (N_13759,N_13642,N_13647);
and U13760 (N_13760,N_13502,N_13693);
or U13761 (N_13761,N_13509,N_13620);
nand U13762 (N_13762,N_13617,N_13656);
nor U13763 (N_13763,N_13583,N_13548);
or U13764 (N_13764,N_13748,N_13621);
nor U13765 (N_13765,N_13562,N_13590);
or U13766 (N_13766,N_13625,N_13588);
nand U13767 (N_13767,N_13657,N_13582);
or U13768 (N_13768,N_13730,N_13613);
or U13769 (N_13769,N_13640,N_13618);
nor U13770 (N_13770,N_13709,N_13506);
nand U13771 (N_13771,N_13595,N_13729);
nor U13772 (N_13772,N_13566,N_13603);
and U13773 (N_13773,N_13623,N_13682);
nor U13774 (N_13774,N_13573,N_13563);
xnor U13775 (N_13775,N_13626,N_13556);
and U13776 (N_13776,N_13578,N_13526);
nand U13777 (N_13777,N_13670,N_13745);
xnor U13778 (N_13778,N_13634,N_13706);
nor U13779 (N_13779,N_13591,N_13511);
or U13780 (N_13780,N_13731,N_13718);
and U13781 (N_13781,N_13669,N_13736);
nor U13782 (N_13782,N_13662,N_13539);
xor U13783 (N_13783,N_13606,N_13505);
or U13784 (N_13784,N_13632,N_13546);
and U13785 (N_13785,N_13512,N_13728);
nand U13786 (N_13786,N_13516,N_13658);
xor U13787 (N_13787,N_13660,N_13587);
nand U13788 (N_13788,N_13576,N_13501);
and U13789 (N_13789,N_13691,N_13712);
and U13790 (N_13790,N_13523,N_13653);
or U13791 (N_13791,N_13609,N_13619);
xor U13792 (N_13792,N_13654,N_13611);
nand U13793 (N_13793,N_13571,N_13503);
or U13794 (N_13794,N_13694,N_13535);
nor U13795 (N_13795,N_13740,N_13637);
nor U13796 (N_13796,N_13724,N_13671);
nor U13797 (N_13797,N_13685,N_13585);
nor U13798 (N_13798,N_13610,N_13560);
and U13799 (N_13799,N_13507,N_13627);
or U13800 (N_13800,N_13710,N_13557);
nor U13801 (N_13801,N_13746,N_13542);
nor U13802 (N_13802,N_13677,N_13711);
nor U13803 (N_13803,N_13581,N_13598);
or U13804 (N_13804,N_13707,N_13584);
xor U13805 (N_13805,N_13579,N_13513);
and U13806 (N_13806,N_13741,N_13600);
and U13807 (N_13807,N_13518,N_13555);
nand U13808 (N_13808,N_13679,N_13597);
nor U13809 (N_13809,N_13565,N_13551);
and U13810 (N_13810,N_13702,N_13726);
nor U13811 (N_13811,N_13547,N_13527);
nor U13812 (N_13812,N_13692,N_13524);
and U13813 (N_13813,N_13529,N_13738);
nor U13814 (N_13814,N_13725,N_13715);
or U13815 (N_13815,N_13686,N_13577);
xor U13816 (N_13816,N_13646,N_13569);
nor U13817 (N_13817,N_13699,N_13586);
nor U13818 (N_13818,N_13567,N_13716);
nor U13819 (N_13819,N_13622,N_13667);
nor U13820 (N_13820,N_13521,N_13528);
nor U13821 (N_13821,N_13676,N_13681);
and U13822 (N_13822,N_13572,N_13631);
nand U13823 (N_13823,N_13544,N_13739);
and U13824 (N_13824,N_13744,N_13604);
and U13825 (N_13825,N_13638,N_13589);
nor U13826 (N_13826,N_13633,N_13703);
nand U13827 (N_13827,N_13648,N_13678);
xnor U13828 (N_13828,N_13517,N_13698);
nand U13829 (N_13829,N_13675,N_13665);
and U13830 (N_13830,N_13515,N_13614);
nor U13831 (N_13831,N_13574,N_13700);
nor U13832 (N_13832,N_13629,N_13680);
nor U13833 (N_13833,N_13538,N_13559);
nor U13834 (N_13834,N_13532,N_13722);
nor U13835 (N_13835,N_13545,N_13690);
or U13836 (N_13836,N_13732,N_13659);
or U13837 (N_13837,N_13534,N_13673);
or U13838 (N_13838,N_13708,N_13561);
and U13839 (N_13839,N_13593,N_13599);
and U13840 (N_13840,N_13701,N_13689);
nor U13841 (N_13841,N_13525,N_13636);
and U13842 (N_13842,N_13522,N_13721);
xor U13843 (N_13843,N_13735,N_13550);
and U13844 (N_13844,N_13608,N_13549);
nor U13845 (N_13845,N_13531,N_13543);
nor U13846 (N_13846,N_13541,N_13553);
or U13847 (N_13847,N_13601,N_13602);
or U13848 (N_13848,N_13592,N_13624);
and U13849 (N_13849,N_13644,N_13533);
nor U13850 (N_13850,N_13530,N_13514);
xnor U13851 (N_13851,N_13695,N_13663);
and U13852 (N_13852,N_13510,N_13734);
or U13853 (N_13853,N_13554,N_13737);
and U13854 (N_13854,N_13645,N_13719);
and U13855 (N_13855,N_13643,N_13733);
nand U13856 (N_13856,N_13500,N_13628);
or U13857 (N_13857,N_13717,N_13705);
and U13858 (N_13858,N_13704,N_13580);
nand U13859 (N_13859,N_13650,N_13641);
and U13860 (N_13860,N_13537,N_13635);
and U13861 (N_13861,N_13661,N_13747);
nor U13862 (N_13862,N_13720,N_13668);
nor U13863 (N_13863,N_13508,N_13568);
or U13864 (N_13864,N_13552,N_13575);
or U13865 (N_13865,N_13607,N_13615);
xor U13866 (N_13866,N_13612,N_13666);
nor U13867 (N_13867,N_13536,N_13696);
nor U13868 (N_13868,N_13714,N_13520);
or U13869 (N_13869,N_13684,N_13743);
or U13870 (N_13870,N_13558,N_13655);
nand U13871 (N_13871,N_13713,N_13742);
or U13872 (N_13872,N_13683,N_13651);
and U13873 (N_13873,N_13564,N_13687);
and U13874 (N_13874,N_13652,N_13688);
nor U13875 (N_13875,N_13572,N_13675);
nor U13876 (N_13876,N_13634,N_13624);
or U13877 (N_13877,N_13685,N_13626);
and U13878 (N_13878,N_13630,N_13633);
or U13879 (N_13879,N_13640,N_13716);
and U13880 (N_13880,N_13708,N_13722);
nor U13881 (N_13881,N_13655,N_13725);
and U13882 (N_13882,N_13667,N_13645);
nor U13883 (N_13883,N_13655,N_13694);
nor U13884 (N_13884,N_13676,N_13519);
nand U13885 (N_13885,N_13714,N_13590);
xor U13886 (N_13886,N_13581,N_13539);
nand U13887 (N_13887,N_13701,N_13737);
nor U13888 (N_13888,N_13676,N_13707);
nor U13889 (N_13889,N_13587,N_13626);
or U13890 (N_13890,N_13691,N_13650);
or U13891 (N_13891,N_13656,N_13669);
nand U13892 (N_13892,N_13708,N_13661);
nand U13893 (N_13893,N_13600,N_13640);
and U13894 (N_13894,N_13715,N_13534);
and U13895 (N_13895,N_13701,N_13544);
and U13896 (N_13896,N_13507,N_13586);
or U13897 (N_13897,N_13645,N_13736);
or U13898 (N_13898,N_13692,N_13655);
nor U13899 (N_13899,N_13704,N_13548);
or U13900 (N_13900,N_13571,N_13741);
nor U13901 (N_13901,N_13535,N_13565);
nor U13902 (N_13902,N_13548,N_13617);
or U13903 (N_13903,N_13740,N_13554);
nor U13904 (N_13904,N_13643,N_13522);
nor U13905 (N_13905,N_13546,N_13677);
or U13906 (N_13906,N_13741,N_13714);
nor U13907 (N_13907,N_13621,N_13710);
nand U13908 (N_13908,N_13541,N_13594);
xor U13909 (N_13909,N_13531,N_13616);
nand U13910 (N_13910,N_13568,N_13654);
or U13911 (N_13911,N_13625,N_13503);
nor U13912 (N_13912,N_13596,N_13665);
and U13913 (N_13913,N_13538,N_13675);
or U13914 (N_13914,N_13653,N_13546);
nand U13915 (N_13915,N_13694,N_13540);
or U13916 (N_13916,N_13620,N_13664);
nor U13917 (N_13917,N_13645,N_13552);
and U13918 (N_13918,N_13718,N_13562);
or U13919 (N_13919,N_13580,N_13571);
nor U13920 (N_13920,N_13730,N_13710);
and U13921 (N_13921,N_13740,N_13583);
or U13922 (N_13922,N_13657,N_13548);
and U13923 (N_13923,N_13739,N_13662);
nor U13924 (N_13924,N_13548,N_13559);
xnor U13925 (N_13925,N_13608,N_13585);
nand U13926 (N_13926,N_13654,N_13609);
nor U13927 (N_13927,N_13505,N_13580);
and U13928 (N_13928,N_13668,N_13723);
nor U13929 (N_13929,N_13512,N_13717);
nor U13930 (N_13930,N_13522,N_13706);
nor U13931 (N_13931,N_13681,N_13665);
nand U13932 (N_13932,N_13578,N_13522);
and U13933 (N_13933,N_13610,N_13689);
nor U13934 (N_13934,N_13747,N_13542);
nand U13935 (N_13935,N_13519,N_13716);
nor U13936 (N_13936,N_13709,N_13645);
or U13937 (N_13937,N_13509,N_13732);
nor U13938 (N_13938,N_13698,N_13649);
nor U13939 (N_13939,N_13631,N_13668);
nand U13940 (N_13940,N_13540,N_13627);
nor U13941 (N_13941,N_13691,N_13591);
xnor U13942 (N_13942,N_13609,N_13642);
nand U13943 (N_13943,N_13579,N_13598);
and U13944 (N_13944,N_13593,N_13743);
nor U13945 (N_13945,N_13604,N_13622);
nor U13946 (N_13946,N_13718,N_13724);
or U13947 (N_13947,N_13641,N_13687);
nor U13948 (N_13948,N_13522,N_13617);
or U13949 (N_13949,N_13567,N_13687);
nor U13950 (N_13950,N_13556,N_13630);
nand U13951 (N_13951,N_13646,N_13635);
nor U13952 (N_13952,N_13593,N_13649);
or U13953 (N_13953,N_13680,N_13715);
or U13954 (N_13954,N_13548,N_13650);
and U13955 (N_13955,N_13642,N_13568);
nor U13956 (N_13956,N_13615,N_13618);
or U13957 (N_13957,N_13717,N_13566);
and U13958 (N_13958,N_13732,N_13541);
or U13959 (N_13959,N_13714,N_13669);
and U13960 (N_13960,N_13570,N_13596);
xnor U13961 (N_13961,N_13668,N_13564);
or U13962 (N_13962,N_13643,N_13542);
or U13963 (N_13963,N_13586,N_13533);
nor U13964 (N_13964,N_13688,N_13732);
and U13965 (N_13965,N_13578,N_13506);
and U13966 (N_13966,N_13727,N_13630);
nor U13967 (N_13967,N_13594,N_13670);
and U13968 (N_13968,N_13612,N_13634);
and U13969 (N_13969,N_13690,N_13556);
or U13970 (N_13970,N_13532,N_13504);
nor U13971 (N_13971,N_13741,N_13637);
nor U13972 (N_13972,N_13602,N_13693);
nor U13973 (N_13973,N_13512,N_13519);
nor U13974 (N_13974,N_13688,N_13532);
nor U13975 (N_13975,N_13676,N_13515);
xnor U13976 (N_13976,N_13674,N_13566);
nor U13977 (N_13977,N_13576,N_13520);
nand U13978 (N_13978,N_13710,N_13661);
nand U13979 (N_13979,N_13671,N_13584);
and U13980 (N_13980,N_13691,N_13655);
or U13981 (N_13981,N_13678,N_13661);
xnor U13982 (N_13982,N_13658,N_13647);
nand U13983 (N_13983,N_13730,N_13602);
nand U13984 (N_13984,N_13544,N_13633);
nand U13985 (N_13985,N_13609,N_13590);
and U13986 (N_13986,N_13607,N_13642);
nand U13987 (N_13987,N_13530,N_13702);
xor U13988 (N_13988,N_13725,N_13660);
or U13989 (N_13989,N_13579,N_13567);
and U13990 (N_13990,N_13678,N_13601);
or U13991 (N_13991,N_13614,N_13744);
or U13992 (N_13992,N_13515,N_13720);
and U13993 (N_13993,N_13672,N_13534);
and U13994 (N_13994,N_13508,N_13737);
or U13995 (N_13995,N_13573,N_13614);
nor U13996 (N_13996,N_13627,N_13700);
nand U13997 (N_13997,N_13600,N_13579);
or U13998 (N_13998,N_13597,N_13703);
nand U13999 (N_13999,N_13556,N_13560);
xnor U14000 (N_14000,N_13827,N_13942);
or U14001 (N_14001,N_13786,N_13814);
and U14002 (N_14002,N_13899,N_13758);
nor U14003 (N_14003,N_13900,N_13916);
nand U14004 (N_14004,N_13773,N_13926);
nand U14005 (N_14005,N_13909,N_13794);
nor U14006 (N_14006,N_13845,N_13933);
nand U14007 (N_14007,N_13980,N_13997);
nand U14008 (N_14008,N_13917,N_13903);
nand U14009 (N_14009,N_13863,N_13800);
xor U14010 (N_14010,N_13757,N_13763);
or U14011 (N_14011,N_13948,N_13904);
or U14012 (N_14012,N_13878,N_13868);
nor U14013 (N_14013,N_13759,N_13831);
nand U14014 (N_14014,N_13879,N_13880);
or U14015 (N_14015,N_13789,N_13784);
xnor U14016 (N_14016,N_13776,N_13986);
or U14017 (N_14017,N_13881,N_13824);
nor U14018 (N_14018,N_13820,N_13849);
or U14019 (N_14019,N_13848,N_13844);
or U14020 (N_14020,N_13927,N_13852);
xnor U14021 (N_14021,N_13872,N_13887);
nand U14022 (N_14022,N_13974,N_13842);
xor U14023 (N_14023,N_13825,N_13817);
nor U14024 (N_14024,N_13875,N_13764);
or U14025 (N_14025,N_13965,N_13962);
and U14026 (N_14026,N_13939,N_13898);
or U14027 (N_14027,N_13755,N_13992);
nor U14028 (N_14028,N_13777,N_13853);
nor U14029 (N_14029,N_13782,N_13778);
and U14030 (N_14030,N_13840,N_13905);
nor U14031 (N_14031,N_13843,N_13988);
xor U14032 (N_14032,N_13972,N_13791);
nand U14033 (N_14033,N_13932,N_13792);
and U14034 (N_14034,N_13924,N_13876);
or U14035 (N_14035,N_13947,N_13799);
nor U14036 (N_14036,N_13921,N_13923);
or U14037 (N_14037,N_13866,N_13877);
or U14038 (N_14038,N_13954,N_13781);
and U14039 (N_14039,N_13772,N_13979);
and U14040 (N_14040,N_13833,N_13841);
and U14041 (N_14041,N_13983,N_13906);
or U14042 (N_14042,N_13822,N_13811);
or U14043 (N_14043,N_13834,N_13801);
and U14044 (N_14044,N_13861,N_13832);
and U14045 (N_14045,N_13934,N_13754);
or U14046 (N_14046,N_13936,N_13808);
or U14047 (N_14047,N_13892,N_13991);
nor U14048 (N_14048,N_13860,N_13810);
nor U14049 (N_14049,N_13989,N_13796);
nor U14050 (N_14050,N_13978,N_13961);
xor U14051 (N_14051,N_13813,N_13968);
or U14052 (N_14052,N_13804,N_13809);
nand U14053 (N_14053,N_13915,N_13886);
and U14054 (N_14054,N_13910,N_13751);
or U14055 (N_14055,N_13768,N_13793);
and U14056 (N_14056,N_13785,N_13753);
and U14057 (N_14057,N_13857,N_13869);
and U14058 (N_14058,N_13984,N_13953);
nor U14059 (N_14059,N_13815,N_13874);
nand U14060 (N_14060,N_13993,N_13994);
or U14061 (N_14061,N_13836,N_13952);
and U14062 (N_14062,N_13889,N_13945);
and U14063 (N_14063,N_13966,N_13911);
or U14064 (N_14064,N_13788,N_13771);
or U14065 (N_14065,N_13920,N_13929);
nor U14066 (N_14066,N_13885,N_13851);
nand U14067 (N_14067,N_13779,N_13805);
or U14068 (N_14068,N_13816,N_13882);
nor U14069 (N_14069,N_13865,N_13873);
nand U14070 (N_14070,N_13985,N_13914);
xnor U14071 (N_14071,N_13750,N_13957);
nor U14072 (N_14072,N_13893,N_13901);
nand U14073 (N_14073,N_13982,N_13996);
and U14074 (N_14074,N_13862,N_13756);
xor U14075 (N_14075,N_13798,N_13821);
nand U14076 (N_14076,N_13956,N_13990);
nor U14077 (N_14077,N_13761,N_13976);
and U14078 (N_14078,N_13971,N_13802);
nand U14079 (N_14079,N_13967,N_13987);
nor U14080 (N_14080,N_13912,N_13839);
or U14081 (N_14081,N_13846,N_13855);
or U14082 (N_14082,N_13891,N_13894);
xnor U14083 (N_14083,N_13977,N_13818);
or U14084 (N_14084,N_13963,N_13871);
or U14085 (N_14085,N_13931,N_13895);
nand U14086 (N_14086,N_13850,N_13765);
and U14087 (N_14087,N_13795,N_13838);
or U14088 (N_14088,N_13925,N_13973);
xnor U14089 (N_14089,N_13888,N_13883);
nor U14090 (N_14090,N_13918,N_13790);
nand U14091 (N_14091,N_13830,N_13870);
or U14092 (N_14092,N_13981,N_13775);
xnor U14093 (N_14093,N_13958,N_13944);
and U14094 (N_14094,N_13950,N_13955);
and U14095 (N_14095,N_13919,N_13884);
or U14096 (N_14096,N_13752,N_13907);
nand U14097 (N_14097,N_13770,N_13995);
or U14098 (N_14098,N_13856,N_13847);
or U14099 (N_14099,N_13959,N_13797);
nand U14100 (N_14100,N_13807,N_13928);
xnor U14101 (N_14101,N_13819,N_13951);
or U14102 (N_14102,N_13999,N_13812);
or U14103 (N_14103,N_13937,N_13837);
nor U14104 (N_14104,N_13829,N_13890);
and U14105 (N_14105,N_13760,N_13835);
or U14106 (N_14106,N_13769,N_13864);
nand U14107 (N_14107,N_13896,N_13908);
nand U14108 (N_14108,N_13766,N_13941);
nor U14109 (N_14109,N_13859,N_13858);
nor U14110 (N_14110,N_13826,N_13975);
nand U14111 (N_14111,N_13762,N_13902);
and U14112 (N_14112,N_13922,N_13823);
or U14113 (N_14113,N_13913,N_13828);
nor U14114 (N_14114,N_13897,N_13867);
and U14115 (N_14115,N_13998,N_13780);
and U14116 (N_14116,N_13787,N_13943);
nand U14117 (N_14117,N_13970,N_13949);
nor U14118 (N_14118,N_13960,N_13938);
or U14119 (N_14119,N_13854,N_13969);
nand U14120 (N_14120,N_13964,N_13806);
nand U14121 (N_14121,N_13774,N_13803);
and U14122 (N_14122,N_13767,N_13783);
nor U14123 (N_14123,N_13946,N_13940);
or U14124 (N_14124,N_13935,N_13930);
nor U14125 (N_14125,N_13815,N_13785);
nor U14126 (N_14126,N_13809,N_13881);
nand U14127 (N_14127,N_13848,N_13785);
nand U14128 (N_14128,N_13788,N_13993);
nand U14129 (N_14129,N_13879,N_13884);
or U14130 (N_14130,N_13757,N_13840);
and U14131 (N_14131,N_13929,N_13973);
and U14132 (N_14132,N_13879,N_13912);
and U14133 (N_14133,N_13941,N_13757);
nor U14134 (N_14134,N_13925,N_13903);
xor U14135 (N_14135,N_13914,N_13974);
and U14136 (N_14136,N_13772,N_13998);
xnor U14137 (N_14137,N_13954,N_13836);
nor U14138 (N_14138,N_13926,N_13885);
or U14139 (N_14139,N_13775,N_13995);
nor U14140 (N_14140,N_13755,N_13777);
and U14141 (N_14141,N_13919,N_13844);
and U14142 (N_14142,N_13824,N_13764);
and U14143 (N_14143,N_13902,N_13925);
nand U14144 (N_14144,N_13797,N_13773);
and U14145 (N_14145,N_13831,N_13789);
nor U14146 (N_14146,N_13942,N_13822);
and U14147 (N_14147,N_13896,N_13750);
and U14148 (N_14148,N_13779,N_13759);
nand U14149 (N_14149,N_13878,N_13957);
or U14150 (N_14150,N_13949,N_13940);
and U14151 (N_14151,N_13920,N_13846);
nor U14152 (N_14152,N_13833,N_13904);
and U14153 (N_14153,N_13826,N_13939);
or U14154 (N_14154,N_13914,N_13771);
nand U14155 (N_14155,N_13954,N_13893);
or U14156 (N_14156,N_13797,N_13832);
or U14157 (N_14157,N_13999,N_13787);
nand U14158 (N_14158,N_13803,N_13760);
nor U14159 (N_14159,N_13807,N_13842);
nand U14160 (N_14160,N_13807,N_13917);
nor U14161 (N_14161,N_13907,N_13864);
nor U14162 (N_14162,N_13795,N_13836);
and U14163 (N_14163,N_13827,N_13881);
and U14164 (N_14164,N_13891,N_13831);
nor U14165 (N_14165,N_13977,N_13984);
nand U14166 (N_14166,N_13787,N_13885);
nand U14167 (N_14167,N_13802,N_13793);
nand U14168 (N_14168,N_13998,N_13815);
nand U14169 (N_14169,N_13829,N_13909);
and U14170 (N_14170,N_13929,N_13900);
nand U14171 (N_14171,N_13861,N_13892);
and U14172 (N_14172,N_13897,N_13766);
and U14173 (N_14173,N_13947,N_13839);
nor U14174 (N_14174,N_13959,N_13785);
nor U14175 (N_14175,N_13876,N_13949);
or U14176 (N_14176,N_13976,N_13856);
and U14177 (N_14177,N_13852,N_13875);
xnor U14178 (N_14178,N_13994,N_13852);
nor U14179 (N_14179,N_13872,N_13785);
nand U14180 (N_14180,N_13812,N_13761);
nand U14181 (N_14181,N_13773,N_13975);
nor U14182 (N_14182,N_13987,N_13834);
and U14183 (N_14183,N_13968,N_13863);
or U14184 (N_14184,N_13888,N_13978);
nor U14185 (N_14185,N_13822,N_13975);
nor U14186 (N_14186,N_13761,N_13931);
and U14187 (N_14187,N_13919,N_13784);
nor U14188 (N_14188,N_13985,N_13979);
or U14189 (N_14189,N_13997,N_13926);
xnor U14190 (N_14190,N_13846,N_13797);
nor U14191 (N_14191,N_13901,N_13832);
xor U14192 (N_14192,N_13792,N_13976);
or U14193 (N_14193,N_13886,N_13977);
nand U14194 (N_14194,N_13825,N_13979);
nand U14195 (N_14195,N_13806,N_13928);
nand U14196 (N_14196,N_13983,N_13773);
nand U14197 (N_14197,N_13922,N_13941);
and U14198 (N_14198,N_13843,N_13877);
or U14199 (N_14199,N_13950,N_13908);
and U14200 (N_14200,N_13782,N_13912);
nand U14201 (N_14201,N_13966,N_13751);
or U14202 (N_14202,N_13991,N_13973);
nor U14203 (N_14203,N_13760,N_13929);
nand U14204 (N_14204,N_13779,N_13870);
and U14205 (N_14205,N_13956,N_13934);
or U14206 (N_14206,N_13821,N_13839);
or U14207 (N_14207,N_13863,N_13959);
or U14208 (N_14208,N_13877,N_13873);
and U14209 (N_14209,N_13974,N_13848);
nand U14210 (N_14210,N_13807,N_13811);
or U14211 (N_14211,N_13777,N_13837);
xor U14212 (N_14212,N_13763,N_13808);
nand U14213 (N_14213,N_13783,N_13803);
or U14214 (N_14214,N_13953,N_13854);
xnor U14215 (N_14215,N_13828,N_13766);
nand U14216 (N_14216,N_13762,N_13961);
nand U14217 (N_14217,N_13962,N_13861);
nand U14218 (N_14218,N_13848,N_13985);
nand U14219 (N_14219,N_13850,N_13842);
nor U14220 (N_14220,N_13812,N_13750);
nand U14221 (N_14221,N_13766,N_13764);
and U14222 (N_14222,N_13941,N_13897);
or U14223 (N_14223,N_13908,N_13877);
or U14224 (N_14224,N_13979,N_13935);
nand U14225 (N_14225,N_13879,N_13917);
and U14226 (N_14226,N_13993,N_13908);
nand U14227 (N_14227,N_13946,N_13779);
nand U14228 (N_14228,N_13967,N_13859);
nor U14229 (N_14229,N_13920,N_13983);
or U14230 (N_14230,N_13910,N_13886);
nor U14231 (N_14231,N_13803,N_13902);
nor U14232 (N_14232,N_13906,N_13818);
and U14233 (N_14233,N_13891,N_13842);
or U14234 (N_14234,N_13859,N_13751);
nand U14235 (N_14235,N_13767,N_13816);
nand U14236 (N_14236,N_13882,N_13899);
and U14237 (N_14237,N_13980,N_13824);
nand U14238 (N_14238,N_13912,N_13841);
or U14239 (N_14239,N_13957,N_13838);
nand U14240 (N_14240,N_13824,N_13768);
or U14241 (N_14241,N_13771,N_13892);
and U14242 (N_14242,N_13965,N_13877);
nand U14243 (N_14243,N_13947,N_13835);
nor U14244 (N_14244,N_13879,N_13819);
nor U14245 (N_14245,N_13960,N_13921);
and U14246 (N_14246,N_13811,N_13956);
and U14247 (N_14247,N_13753,N_13789);
or U14248 (N_14248,N_13972,N_13919);
xor U14249 (N_14249,N_13906,N_13790);
xor U14250 (N_14250,N_14027,N_14071);
nor U14251 (N_14251,N_14019,N_14119);
and U14252 (N_14252,N_14125,N_14033);
or U14253 (N_14253,N_14200,N_14085);
nand U14254 (N_14254,N_14065,N_14234);
nand U14255 (N_14255,N_14205,N_14016);
nand U14256 (N_14256,N_14068,N_14081);
and U14257 (N_14257,N_14003,N_14172);
or U14258 (N_14258,N_14020,N_14182);
nor U14259 (N_14259,N_14127,N_14115);
nor U14260 (N_14260,N_14195,N_14135);
nand U14261 (N_14261,N_14140,N_14201);
nor U14262 (N_14262,N_14225,N_14228);
or U14263 (N_14263,N_14030,N_14211);
nor U14264 (N_14264,N_14209,N_14112);
nor U14265 (N_14265,N_14212,N_14208);
nor U14266 (N_14266,N_14083,N_14248);
nand U14267 (N_14267,N_14072,N_14063);
or U14268 (N_14268,N_14196,N_14165);
or U14269 (N_14269,N_14224,N_14036);
and U14270 (N_14270,N_14064,N_14107);
nor U14271 (N_14271,N_14075,N_14077);
nand U14272 (N_14272,N_14168,N_14181);
nand U14273 (N_14273,N_14050,N_14220);
or U14274 (N_14274,N_14169,N_14149);
xor U14275 (N_14275,N_14092,N_14244);
and U14276 (N_14276,N_14154,N_14150);
or U14277 (N_14277,N_14034,N_14194);
nor U14278 (N_14278,N_14192,N_14162);
nor U14279 (N_14279,N_14018,N_14185);
xnor U14280 (N_14280,N_14067,N_14137);
nor U14281 (N_14281,N_14025,N_14114);
or U14282 (N_14282,N_14032,N_14179);
or U14283 (N_14283,N_14005,N_14221);
or U14284 (N_14284,N_14245,N_14229);
and U14285 (N_14285,N_14111,N_14055);
or U14286 (N_14286,N_14106,N_14082);
nand U14287 (N_14287,N_14101,N_14223);
nand U14288 (N_14288,N_14084,N_14163);
and U14289 (N_14289,N_14045,N_14178);
nor U14290 (N_14290,N_14053,N_14131);
and U14291 (N_14291,N_14061,N_14096);
and U14292 (N_14292,N_14060,N_14059);
nand U14293 (N_14293,N_14120,N_14191);
or U14294 (N_14294,N_14143,N_14100);
or U14295 (N_14295,N_14177,N_14237);
nand U14296 (N_14296,N_14159,N_14066);
nand U14297 (N_14297,N_14156,N_14022);
nand U14298 (N_14298,N_14117,N_14186);
and U14299 (N_14299,N_14011,N_14146);
nand U14300 (N_14300,N_14057,N_14029);
nand U14301 (N_14301,N_14031,N_14189);
nand U14302 (N_14302,N_14128,N_14051);
nor U14303 (N_14303,N_14086,N_14008);
nand U14304 (N_14304,N_14080,N_14023);
nand U14305 (N_14305,N_14009,N_14171);
xnor U14306 (N_14306,N_14142,N_14139);
nand U14307 (N_14307,N_14166,N_14155);
nand U14308 (N_14308,N_14144,N_14052);
xnor U14309 (N_14309,N_14090,N_14222);
nand U14310 (N_14310,N_14152,N_14199);
nor U14311 (N_14311,N_14094,N_14048);
nor U14312 (N_14312,N_14037,N_14238);
and U14313 (N_14313,N_14188,N_14054);
nor U14314 (N_14314,N_14180,N_14113);
and U14315 (N_14315,N_14078,N_14138);
and U14316 (N_14316,N_14157,N_14073);
and U14317 (N_14317,N_14001,N_14058);
nor U14318 (N_14318,N_14148,N_14242);
or U14319 (N_14319,N_14176,N_14207);
nand U14320 (N_14320,N_14004,N_14197);
nor U14321 (N_14321,N_14006,N_14151);
and U14322 (N_14322,N_14217,N_14216);
and U14323 (N_14323,N_14183,N_14091);
nor U14324 (N_14324,N_14193,N_14088);
nand U14325 (N_14325,N_14133,N_14028);
nor U14326 (N_14326,N_14041,N_14102);
or U14327 (N_14327,N_14012,N_14121);
or U14328 (N_14328,N_14239,N_14235);
xnor U14329 (N_14329,N_14219,N_14035);
xor U14330 (N_14330,N_14206,N_14056);
or U14331 (N_14331,N_14174,N_14203);
nand U14332 (N_14332,N_14110,N_14026);
nand U14333 (N_14333,N_14069,N_14126);
or U14334 (N_14334,N_14187,N_14062);
and U14335 (N_14335,N_14099,N_14095);
nor U14336 (N_14336,N_14214,N_14087);
and U14337 (N_14337,N_14098,N_14044);
or U14338 (N_14338,N_14042,N_14000);
nor U14339 (N_14339,N_14132,N_14202);
or U14340 (N_14340,N_14118,N_14007);
nand U14341 (N_14341,N_14164,N_14122);
nand U14342 (N_14342,N_14230,N_14184);
or U14343 (N_14343,N_14145,N_14215);
nand U14344 (N_14344,N_14014,N_14213);
nor U14345 (N_14345,N_14038,N_14103);
and U14346 (N_14346,N_14232,N_14240);
and U14347 (N_14347,N_14043,N_14013);
nand U14348 (N_14348,N_14141,N_14097);
and U14349 (N_14349,N_14116,N_14231);
xnor U14350 (N_14350,N_14161,N_14175);
or U14351 (N_14351,N_14198,N_14070);
nand U14352 (N_14352,N_14249,N_14093);
or U14353 (N_14353,N_14190,N_14109);
or U14354 (N_14354,N_14124,N_14024);
nand U14355 (N_14355,N_14104,N_14241);
nand U14356 (N_14356,N_14233,N_14015);
nor U14357 (N_14357,N_14079,N_14153);
nand U14358 (N_14358,N_14089,N_14002);
nor U14359 (N_14359,N_14218,N_14170);
nor U14360 (N_14360,N_14236,N_14123);
nor U14361 (N_14361,N_14134,N_14021);
and U14362 (N_14362,N_14173,N_14227);
nand U14363 (N_14363,N_14010,N_14129);
and U14364 (N_14364,N_14136,N_14074);
nand U14365 (N_14365,N_14160,N_14039);
or U14366 (N_14366,N_14204,N_14017);
or U14367 (N_14367,N_14105,N_14247);
or U14368 (N_14368,N_14046,N_14147);
nor U14369 (N_14369,N_14246,N_14226);
nand U14370 (N_14370,N_14158,N_14076);
and U14371 (N_14371,N_14130,N_14243);
xnor U14372 (N_14372,N_14108,N_14040);
nand U14373 (N_14373,N_14047,N_14210);
and U14374 (N_14374,N_14049,N_14167);
xor U14375 (N_14375,N_14123,N_14010);
nand U14376 (N_14376,N_14127,N_14058);
or U14377 (N_14377,N_14213,N_14239);
nand U14378 (N_14378,N_14182,N_14030);
xor U14379 (N_14379,N_14024,N_14244);
and U14380 (N_14380,N_14246,N_14132);
nand U14381 (N_14381,N_14152,N_14209);
or U14382 (N_14382,N_14073,N_14137);
or U14383 (N_14383,N_14024,N_14232);
and U14384 (N_14384,N_14169,N_14136);
or U14385 (N_14385,N_14023,N_14183);
nand U14386 (N_14386,N_14238,N_14189);
or U14387 (N_14387,N_14206,N_14077);
or U14388 (N_14388,N_14088,N_14222);
nand U14389 (N_14389,N_14223,N_14181);
and U14390 (N_14390,N_14224,N_14120);
and U14391 (N_14391,N_14042,N_14078);
nor U14392 (N_14392,N_14017,N_14111);
and U14393 (N_14393,N_14154,N_14241);
and U14394 (N_14394,N_14100,N_14216);
and U14395 (N_14395,N_14112,N_14005);
or U14396 (N_14396,N_14061,N_14127);
nand U14397 (N_14397,N_14128,N_14133);
and U14398 (N_14398,N_14241,N_14080);
or U14399 (N_14399,N_14077,N_14012);
nand U14400 (N_14400,N_14076,N_14040);
xnor U14401 (N_14401,N_14105,N_14042);
and U14402 (N_14402,N_14082,N_14116);
nor U14403 (N_14403,N_14057,N_14154);
nor U14404 (N_14404,N_14203,N_14121);
or U14405 (N_14405,N_14110,N_14108);
or U14406 (N_14406,N_14134,N_14096);
nand U14407 (N_14407,N_14123,N_14025);
or U14408 (N_14408,N_14004,N_14138);
nand U14409 (N_14409,N_14066,N_14048);
or U14410 (N_14410,N_14101,N_14131);
nand U14411 (N_14411,N_14176,N_14230);
nor U14412 (N_14412,N_14207,N_14246);
nand U14413 (N_14413,N_14132,N_14228);
or U14414 (N_14414,N_14081,N_14143);
or U14415 (N_14415,N_14082,N_14016);
nor U14416 (N_14416,N_14016,N_14052);
and U14417 (N_14417,N_14124,N_14234);
nor U14418 (N_14418,N_14064,N_14047);
and U14419 (N_14419,N_14236,N_14000);
and U14420 (N_14420,N_14117,N_14015);
or U14421 (N_14421,N_14160,N_14209);
and U14422 (N_14422,N_14210,N_14213);
and U14423 (N_14423,N_14025,N_14077);
nor U14424 (N_14424,N_14025,N_14239);
or U14425 (N_14425,N_14093,N_14190);
nand U14426 (N_14426,N_14149,N_14029);
or U14427 (N_14427,N_14132,N_14010);
nand U14428 (N_14428,N_14216,N_14248);
nand U14429 (N_14429,N_14196,N_14068);
nor U14430 (N_14430,N_14217,N_14124);
and U14431 (N_14431,N_14168,N_14248);
nand U14432 (N_14432,N_14123,N_14008);
xnor U14433 (N_14433,N_14121,N_14165);
nor U14434 (N_14434,N_14018,N_14110);
or U14435 (N_14435,N_14151,N_14079);
or U14436 (N_14436,N_14205,N_14209);
and U14437 (N_14437,N_14158,N_14137);
and U14438 (N_14438,N_14086,N_14034);
nand U14439 (N_14439,N_14200,N_14028);
xnor U14440 (N_14440,N_14198,N_14154);
nand U14441 (N_14441,N_14125,N_14002);
nand U14442 (N_14442,N_14210,N_14127);
nor U14443 (N_14443,N_14090,N_14011);
nand U14444 (N_14444,N_14188,N_14217);
nand U14445 (N_14445,N_14028,N_14087);
nor U14446 (N_14446,N_14078,N_14184);
and U14447 (N_14447,N_14247,N_14092);
and U14448 (N_14448,N_14005,N_14076);
or U14449 (N_14449,N_14021,N_14227);
nor U14450 (N_14450,N_14100,N_14186);
xnor U14451 (N_14451,N_14121,N_14236);
or U14452 (N_14452,N_14237,N_14057);
and U14453 (N_14453,N_14187,N_14024);
and U14454 (N_14454,N_14075,N_14057);
nand U14455 (N_14455,N_14178,N_14198);
nor U14456 (N_14456,N_14225,N_14015);
or U14457 (N_14457,N_14001,N_14168);
and U14458 (N_14458,N_14143,N_14090);
nor U14459 (N_14459,N_14135,N_14148);
or U14460 (N_14460,N_14174,N_14079);
nand U14461 (N_14461,N_14007,N_14012);
nand U14462 (N_14462,N_14167,N_14215);
nor U14463 (N_14463,N_14156,N_14164);
and U14464 (N_14464,N_14085,N_14084);
or U14465 (N_14465,N_14056,N_14028);
nor U14466 (N_14466,N_14033,N_14184);
xor U14467 (N_14467,N_14170,N_14174);
or U14468 (N_14468,N_14020,N_14047);
and U14469 (N_14469,N_14119,N_14081);
and U14470 (N_14470,N_14131,N_14144);
xnor U14471 (N_14471,N_14222,N_14137);
and U14472 (N_14472,N_14149,N_14109);
nor U14473 (N_14473,N_14047,N_14022);
nor U14474 (N_14474,N_14046,N_14139);
or U14475 (N_14475,N_14241,N_14034);
and U14476 (N_14476,N_14071,N_14233);
nand U14477 (N_14477,N_14069,N_14002);
and U14478 (N_14478,N_14191,N_14065);
nor U14479 (N_14479,N_14179,N_14241);
nand U14480 (N_14480,N_14226,N_14040);
nand U14481 (N_14481,N_14006,N_14166);
nor U14482 (N_14482,N_14017,N_14160);
nand U14483 (N_14483,N_14239,N_14212);
nor U14484 (N_14484,N_14205,N_14027);
and U14485 (N_14485,N_14192,N_14229);
nor U14486 (N_14486,N_14199,N_14204);
and U14487 (N_14487,N_14179,N_14195);
or U14488 (N_14488,N_14200,N_14191);
nand U14489 (N_14489,N_14012,N_14134);
nor U14490 (N_14490,N_14136,N_14176);
nand U14491 (N_14491,N_14034,N_14109);
nor U14492 (N_14492,N_14038,N_14018);
nand U14493 (N_14493,N_14100,N_14047);
nand U14494 (N_14494,N_14247,N_14013);
nor U14495 (N_14495,N_14248,N_14128);
nand U14496 (N_14496,N_14210,N_14248);
or U14497 (N_14497,N_14246,N_14249);
nor U14498 (N_14498,N_14032,N_14053);
nor U14499 (N_14499,N_14005,N_14231);
or U14500 (N_14500,N_14307,N_14299);
or U14501 (N_14501,N_14374,N_14303);
nand U14502 (N_14502,N_14274,N_14305);
nor U14503 (N_14503,N_14285,N_14356);
or U14504 (N_14504,N_14316,N_14369);
or U14505 (N_14505,N_14329,N_14338);
or U14506 (N_14506,N_14460,N_14428);
xor U14507 (N_14507,N_14270,N_14280);
xor U14508 (N_14508,N_14416,N_14392);
and U14509 (N_14509,N_14425,N_14447);
or U14510 (N_14510,N_14282,N_14423);
nor U14511 (N_14511,N_14490,N_14441);
and U14512 (N_14512,N_14367,N_14343);
nor U14513 (N_14513,N_14276,N_14284);
and U14514 (N_14514,N_14375,N_14349);
and U14515 (N_14515,N_14334,N_14293);
or U14516 (N_14516,N_14308,N_14250);
and U14517 (N_14517,N_14398,N_14278);
and U14518 (N_14518,N_14409,N_14326);
nand U14519 (N_14519,N_14281,N_14333);
or U14520 (N_14520,N_14489,N_14471);
and U14521 (N_14521,N_14472,N_14484);
and U14522 (N_14522,N_14351,N_14426);
or U14523 (N_14523,N_14394,N_14256);
or U14524 (N_14524,N_14380,N_14422);
nand U14525 (N_14525,N_14314,N_14434);
xor U14526 (N_14526,N_14451,N_14306);
or U14527 (N_14527,N_14266,N_14468);
and U14528 (N_14528,N_14442,N_14264);
nand U14529 (N_14529,N_14494,N_14353);
or U14530 (N_14530,N_14404,N_14363);
nand U14531 (N_14531,N_14301,N_14342);
nor U14532 (N_14532,N_14435,N_14432);
nand U14533 (N_14533,N_14324,N_14372);
nand U14534 (N_14534,N_14357,N_14302);
and U14535 (N_14535,N_14393,N_14295);
and U14536 (N_14536,N_14262,N_14366);
or U14537 (N_14537,N_14355,N_14354);
nand U14538 (N_14538,N_14454,N_14457);
and U14539 (N_14539,N_14257,N_14352);
nand U14540 (N_14540,N_14283,N_14419);
xnor U14541 (N_14541,N_14481,N_14347);
nor U14542 (N_14542,N_14474,N_14444);
or U14543 (N_14543,N_14414,N_14410);
xnor U14544 (N_14544,N_14327,N_14325);
or U14545 (N_14545,N_14383,N_14368);
and U14546 (N_14546,N_14438,N_14406);
nand U14547 (N_14547,N_14261,N_14498);
nor U14548 (N_14548,N_14408,N_14331);
or U14549 (N_14549,N_14317,N_14297);
and U14550 (N_14550,N_14350,N_14479);
or U14551 (N_14551,N_14470,N_14411);
nand U14552 (N_14552,N_14493,N_14277);
nand U14553 (N_14553,N_14449,N_14311);
nand U14554 (N_14554,N_14415,N_14348);
and U14555 (N_14555,N_14332,N_14461);
or U14556 (N_14556,N_14495,N_14260);
xnor U14557 (N_14557,N_14464,N_14429);
and U14558 (N_14558,N_14336,N_14279);
or U14559 (N_14559,N_14358,N_14251);
and U14560 (N_14560,N_14466,N_14364);
nor U14561 (N_14561,N_14335,N_14252);
nor U14562 (N_14562,N_14390,N_14319);
or U14563 (N_14563,N_14405,N_14321);
and U14564 (N_14564,N_14318,N_14371);
nand U14565 (N_14565,N_14439,N_14340);
or U14566 (N_14566,N_14476,N_14480);
or U14567 (N_14567,N_14491,N_14482);
xnor U14568 (N_14568,N_14492,N_14395);
and U14569 (N_14569,N_14269,N_14310);
xnor U14570 (N_14570,N_14463,N_14437);
nand U14571 (N_14571,N_14268,N_14487);
nand U14572 (N_14572,N_14385,N_14328);
nand U14573 (N_14573,N_14396,N_14477);
and U14574 (N_14574,N_14388,N_14397);
nand U14575 (N_14575,N_14499,N_14465);
and U14576 (N_14576,N_14259,N_14373);
xor U14577 (N_14577,N_14475,N_14272);
nand U14578 (N_14578,N_14407,N_14453);
or U14579 (N_14579,N_14273,N_14459);
nor U14580 (N_14580,N_14300,N_14433);
xnor U14581 (N_14581,N_14417,N_14399);
or U14582 (N_14582,N_14362,N_14483);
nand U14583 (N_14583,N_14253,N_14309);
xor U14584 (N_14584,N_14298,N_14421);
or U14585 (N_14585,N_14486,N_14275);
nor U14586 (N_14586,N_14361,N_14296);
and U14587 (N_14587,N_14455,N_14391);
nor U14588 (N_14588,N_14462,N_14267);
and U14589 (N_14589,N_14401,N_14379);
xor U14590 (N_14590,N_14389,N_14381);
nor U14591 (N_14591,N_14452,N_14387);
nand U14592 (N_14592,N_14400,N_14344);
nand U14593 (N_14593,N_14478,N_14377);
or U14594 (N_14594,N_14496,N_14420);
and U14595 (N_14595,N_14445,N_14263);
nand U14596 (N_14596,N_14485,N_14291);
and U14597 (N_14597,N_14431,N_14418);
and U14598 (N_14598,N_14488,N_14255);
and U14599 (N_14599,N_14430,N_14287);
nand U14600 (N_14600,N_14382,N_14378);
xnor U14601 (N_14601,N_14446,N_14286);
and U14602 (N_14602,N_14473,N_14288);
or U14603 (N_14603,N_14312,N_14467);
and U14604 (N_14604,N_14376,N_14386);
nand U14605 (N_14605,N_14402,N_14427);
and U14606 (N_14606,N_14313,N_14271);
nand U14607 (N_14607,N_14359,N_14450);
nand U14608 (N_14608,N_14370,N_14384);
or U14609 (N_14609,N_14304,N_14289);
and U14610 (N_14610,N_14341,N_14458);
nand U14611 (N_14611,N_14254,N_14436);
or U14612 (N_14612,N_14448,N_14294);
or U14613 (N_14613,N_14323,N_14456);
and U14614 (N_14614,N_14443,N_14346);
nand U14615 (N_14615,N_14360,N_14403);
nor U14616 (N_14616,N_14258,N_14412);
or U14617 (N_14617,N_14292,N_14469);
nand U14618 (N_14618,N_14322,N_14345);
xnor U14619 (N_14619,N_14290,N_14337);
nor U14620 (N_14620,N_14320,N_14265);
or U14621 (N_14621,N_14440,N_14497);
xnor U14622 (N_14622,N_14413,N_14424);
or U14623 (N_14623,N_14315,N_14365);
or U14624 (N_14624,N_14339,N_14330);
or U14625 (N_14625,N_14484,N_14326);
xnor U14626 (N_14626,N_14447,N_14344);
or U14627 (N_14627,N_14498,N_14393);
and U14628 (N_14628,N_14355,N_14388);
and U14629 (N_14629,N_14484,N_14417);
nor U14630 (N_14630,N_14330,N_14294);
and U14631 (N_14631,N_14485,N_14438);
and U14632 (N_14632,N_14344,N_14373);
nand U14633 (N_14633,N_14392,N_14353);
or U14634 (N_14634,N_14413,N_14335);
and U14635 (N_14635,N_14377,N_14434);
nand U14636 (N_14636,N_14457,N_14253);
nand U14637 (N_14637,N_14293,N_14272);
xnor U14638 (N_14638,N_14266,N_14435);
nor U14639 (N_14639,N_14425,N_14293);
or U14640 (N_14640,N_14466,N_14457);
nand U14641 (N_14641,N_14430,N_14378);
or U14642 (N_14642,N_14324,N_14413);
or U14643 (N_14643,N_14450,N_14443);
nor U14644 (N_14644,N_14457,N_14425);
or U14645 (N_14645,N_14394,N_14318);
and U14646 (N_14646,N_14346,N_14447);
and U14647 (N_14647,N_14276,N_14321);
and U14648 (N_14648,N_14333,N_14314);
nand U14649 (N_14649,N_14463,N_14325);
or U14650 (N_14650,N_14261,N_14467);
and U14651 (N_14651,N_14307,N_14341);
nand U14652 (N_14652,N_14299,N_14285);
nor U14653 (N_14653,N_14482,N_14354);
nor U14654 (N_14654,N_14329,N_14397);
xnor U14655 (N_14655,N_14337,N_14468);
xnor U14656 (N_14656,N_14490,N_14361);
nor U14657 (N_14657,N_14268,N_14383);
and U14658 (N_14658,N_14352,N_14435);
xnor U14659 (N_14659,N_14371,N_14280);
or U14660 (N_14660,N_14280,N_14305);
nor U14661 (N_14661,N_14290,N_14353);
and U14662 (N_14662,N_14392,N_14253);
or U14663 (N_14663,N_14405,N_14379);
nor U14664 (N_14664,N_14315,N_14347);
and U14665 (N_14665,N_14259,N_14348);
or U14666 (N_14666,N_14447,N_14450);
nand U14667 (N_14667,N_14372,N_14359);
nor U14668 (N_14668,N_14293,N_14325);
or U14669 (N_14669,N_14448,N_14410);
or U14670 (N_14670,N_14412,N_14372);
nand U14671 (N_14671,N_14369,N_14254);
or U14672 (N_14672,N_14342,N_14487);
nand U14673 (N_14673,N_14284,N_14433);
nor U14674 (N_14674,N_14420,N_14395);
nand U14675 (N_14675,N_14462,N_14265);
xor U14676 (N_14676,N_14485,N_14360);
nor U14677 (N_14677,N_14473,N_14429);
nor U14678 (N_14678,N_14277,N_14299);
or U14679 (N_14679,N_14479,N_14461);
or U14680 (N_14680,N_14498,N_14276);
and U14681 (N_14681,N_14444,N_14473);
nor U14682 (N_14682,N_14269,N_14366);
nor U14683 (N_14683,N_14448,N_14407);
nor U14684 (N_14684,N_14429,N_14463);
or U14685 (N_14685,N_14311,N_14373);
nand U14686 (N_14686,N_14284,N_14333);
and U14687 (N_14687,N_14302,N_14385);
nor U14688 (N_14688,N_14403,N_14491);
nand U14689 (N_14689,N_14496,N_14273);
or U14690 (N_14690,N_14352,N_14259);
xor U14691 (N_14691,N_14354,N_14330);
nand U14692 (N_14692,N_14478,N_14301);
or U14693 (N_14693,N_14377,N_14250);
or U14694 (N_14694,N_14385,N_14252);
nor U14695 (N_14695,N_14474,N_14400);
and U14696 (N_14696,N_14439,N_14434);
xor U14697 (N_14697,N_14314,N_14390);
and U14698 (N_14698,N_14491,N_14497);
or U14699 (N_14699,N_14449,N_14267);
or U14700 (N_14700,N_14350,N_14492);
nor U14701 (N_14701,N_14373,N_14287);
nor U14702 (N_14702,N_14390,N_14364);
or U14703 (N_14703,N_14255,N_14400);
nor U14704 (N_14704,N_14476,N_14251);
nor U14705 (N_14705,N_14307,N_14351);
nand U14706 (N_14706,N_14421,N_14319);
nand U14707 (N_14707,N_14311,N_14284);
or U14708 (N_14708,N_14440,N_14281);
nand U14709 (N_14709,N_14413,N_14471);
and U14710 (N_14710,N_14289,N_14285);
or U14711 (N_14711,N_14288,N_14338);
or U14712 (N_14712,N_14497,N_14431);
and U14713 (N_14713,N_14345,N_14261);
nor U14714 (N_14714,N_14398,N_14330);
nand U14715 (N_14715,N_14491,N_14419);
or U14716 (N_14716,N_14434,N_14473);
or U14717 (N_14717,N_14256,N_14446);
nor U14718 (N_14718,N_14312,N_14405);
or U14719 (N_14719,N_14328,N_14295);
nand U14720 (N_14720,N_14484,N_14468);
nor U14721 (N_14721,N_14295,N_14345);
nand U14722 (N_14722,N_14318,N_14376);
or U14723 (N_14723,N_14449,N_14251);
and U14724 (N_14724,N_14428,N_14421);
or U14725 (N_14725,N_14330,N_14426);
nor U14726 (N_14726,N_14456,N_14304);
and U14727 (N_14727,N_14313,N_14438);
nor U14728 (N_14728,N_14263,N_14458);
or U14729 (N_14729,N_14326,N_14441);
and U14730 (N_14730,N_14250,N_14444);
xor U14731 (N_14731,N_14399,N_14312);
xor U14732 (N_14732,N_14290,N_14392);
or U14733 (N_14733,N_14328,N_14298);
and U14734 (N_14734,N_14431,N_14485);
and U14735 (N_14735,N_14452,N_14440);
and U14736 (N_14736,N_14253,N_14329);
and U14737 (N_14737,N_14415,N_14262);
nor U14738 (N_14738,N_14289,N_14401);
nand U14739 (N_14739,N_14310,N_14456);
nor U14740 (N_14740,N_14420,N_14331);
xnor U14741 (N_14741,N_14304,N_14438);
nor U14742 (N_14742,N_14379,N_14406);
and U14743 (N_14743,N_14442,N_14308);
nand U14744 (N_14744,N_14461,N_14324);
nand U14745 (N_14745,N_14447,N_14302);
xnor U14746 (N_14746,N_14445,N_14320);
and U14747 (N_14747,N_14299,N_14259);
nand U14748 (N_14748,N_14260,N_14290);
nor U14749 (N_14749,N_14333,N_14425);
or U14750 (N_14750,N_14729,N_14564);
or U14751 (N_14751,N_14594,N_14681);
and U14752 (N_14752,N_14561,N_14513);
nand U14753 (N_14753,N_14745,N_14726);
nand U14754 (N_14754,N_14610,N_14715);
or U14755 (N_14755,N_14504,N_14735);
or U14756 (N_14756,N_14728,N_14690);
and U14757 (N_14757,N_14687,N_14623);
nand U14758 (N_14758,N_14702,N_14721);
nor U14759 (N_14759,N_14588,N_14636);
or U14760 (N_14760,N_14551,N_14746);
or U14761 (N_14761,N_14549,N_14632);
or U14762 (N_14762,N_14619,N_14615);
and U14763 (N_14763,N_14696,N_14624);
or U14764 (N_14764,N_14714,N_14741);
or U14765 (N_14765,N_14628,N_14571);
nand U14766 (N_14766,N_14502,N_14575);
nor U14767 (N_14767,N_14531,N_14693);
and U14768 (N_14768,N_14734,N_14583);
xor U14769 (N_14769,N_14650,N_14676);
nand U14770 (N_14770,N_14621,N_14671);
or U14771 (N_14771,N_14568,N_14518);
and U14772 (N_14772,N_14592,N_14521);
nor U14773 (N_14773,N_14709,N_14700);
xnor U14774 (N_14774,N_14566,N_14530);
and U14775 (N_14775,N_14581,N_14540);
and U14776 (N_14776,N_14682,N_14578);
nand U14777 (N_14777,N_14717,N_14607);
or U14778 (N_14778,N_14556,N_14674);
nor U14779 (N_14779,N_14668,N_14543);
or U14780 (N_14780,N_14641,N_14582);
nand U14781 (N_14781,N_14595,N_14579);
nand U14782 (N_14782,N_14562,N_14697);
nor U14783 (N_14783,N_14644,N_14679);
nor U14784 (N_14784,N_14605,N_14684);
nand U14785 (N_14785,N_14538,N_14550);
nor U14786 (N_14786,N_14629,N_14638);
nand U14787 (N_14787,N_14665,N_14639);
or U14788 (N_14788,N_14739,N_14585);
xnor U14789 (N_14789,N_14706,N_14612);
or U14790 (N_14790,N_14507,N_14692);
nand U14791 (N_14791,N_14705,N_14733);
nand U14792 (N_14792,N_14618,N_14673);
nand U14793 (N_14793,N_14635,N_14569);
nand U14794 (N_14794,N_14511,N_14565);
or U14795 (N_14795,N_14694,N_14500);
nor U14796 (N_14796,N_14512,N_14663);
and U14797 (N_14797,N_14652,N_14712);
nor U14798 (N_14798,N_14608,N_14600);
nor U14799 (N_14799,N_14601,N_14554);
nor U14800 (N_14800,N_14630,N_14670);
nand U14801 (N_14801,N_14738,N_14730);
or U14802 (N_14802,N_14688,N_14508);
nand U14803 (N_14803,N_14748,N_14537);
nor U14804 (N_14804,N_14517,N_14699);
or U14805 (N_14805,N_14707,N_14660);
nor U14806 (N_14806,N_14558,N_14541);
xor U14807 (N_14807,N_14719,N_14553);
xor U14808 (N_14808,N_14529,N_14576);
nor U14809 (N_14809,N_14614,N_14666);
nor U14810 (N_14810,N_14677,N_14524);
or U14811 (N_14811,N_14573,N_14503);
nor U14812 (N_14812,N_14539,N_14593);
and U14813 (N_14813,N_14557,N_14604);
nor U14814 (N_14814,N_14742,N_14722);
nand U14815 (N_14815,N_14546,N_14545);
nand U14816 (N_14816,N_14625,N_14747);
or U14817 (N_14817,N_14515,N_14662);
nand U14818 (N_14818,N_14737,N_14648);
nand U14819 (N_14819,N_14678,N_14590);
and U14820 (N_14820,N_14643,N_14613);
and U14821 (N_14821,N_14544,N_14718);
or U14822 (N_14822,N_14528,N_14520);
nand U14823 (N_14823,N_14727,N_14523);
nand U14824 (N_14824,N_14620,N_14708);
nor U14825 (N_14825,N_14559,N_14563);
or U14826 (N_14826,N_14640,N_14606);
or U14827 (N_14827,N_14580,N_14634);
nor U14828 (N_14828,N_14647,N_14536);
nor U14829 (N_14829,N_14587,N_14514);
or U14830 (N_14830,N_14725,N_14586);
and U14831 (N_14831,N_14691,N_14599);
and U14832 (N_14832,N_14532,N_14589);
nand U14833 (N_14833,N_14616,N_14720);
nand U14834 (N_14834,N_14637,N_14659);
and U14835 (N_14835,N_14732,N_14667);
xnor U14836 (N_14836,N_14574,N_14710);
or U14837 (N_14837,N_14649,N_14555);
or U14838 (N_14838,N_14617,N_14533);
and U14839 (N_14839,N_14716,N_14548);
or U14840 (N_14840,N_14685,N_14547);
xor U14841 (N_14841,N_14611,N_14552);
nor U14842 (N_14842,N_14686,N_14598);
or U14843 (N_14843,N_14658,N_14519);
nor U14844 (N_14844,N_14645,N_14669);
nand U14845 (N_14845,N_14522,N_14653);
nor U14846 (N_14846,N_14744,N_14560);
nor U14847 (N_14847,N_14654,N_14633);
nor U14848 (N_14848,N_14631,N_14743);
nor U14849 (N_14849,N_14534,N_14596);
xnor U14850 (N_14850,N_14506,N_14661);
and U14851 (N_14851,N_14703,N_14570);
nor U14852 (N_14852,N_14651,N_14704);
or U14853 (N_14853,N_14510,N_14591);
nand U14854 (N_14854,N_14642,N_14572);
nor U14855 (N_14855,N_14683,N_14736);
nor U14856 (N_14856,N_14698,N_14622);
and U14857 (N_14857,N_14603,N_14680);
or U14858 (N_14858,N_14501,N_14609);
and U14859 (N_14859,N_14731,N_14602);
nor U14860 (N_14860,N_14509,N_14542);
nor U14861 (N_14861,N_14646,N_14657);
xnor U14862 (N_14862,N_14526,N_14689);
or U14863 (N_14863,N_14656,N_14505);
nor U14864 (N_14864,N_14701,N_14713);
nand U14865 (N_14865,N_14597,N_14672);
or U14866 (N_14866,N_14664,N_14655);
nor U14867 (N_14867,N_14627,N_14723);
nor U14868 (N_14868,N_14675,N_14711);
or U14869 (N_14869,N_14525,N_14740);
nand U14870 (N_14870,N_14577,N_14516);
nand U14871 (N_14871,N_14567,N_14749);
nor U14872 (N_14872,N_14626,N_14584);
or U14873 (N_14873,N_14535,N_14527);
nor U14874 (N_14874,N_14724,N_14695);
or U14875 (N_14875,N_14634,N_14522);
or U14876 (N_14876,N_14672,N_14725);
nand U14877 (N_14877,N_14501,N_14560);
or U14878 (N_14878,N_14705,N_14698);
or U14879 (N_14879,N_14561,N_14627);
nor U14880 (N_14880,N_14569,N_14621);
nor U14881 (N_14881,N_14518,N_14557);
nor U14882 (N_14882,N_14549,N_14602);
nand U14883 (N_14883,N_14724,N_14700);
nor U14884 (N_14884,N_14507,N_14626);
nor U14885 (N_14885,N_14627,N_14529);
and U14886 (N_14886,N_14673,N_14554);
nand U14887 (N_14887,N_14524,N_14601);
nand U14888 (N_14888,N_14516,N_14624);
or U14889 (N_14889,N_14713,N_14704);
nand U14890 (N_14890,N_14572,N_14680);
nor U14891 (N_14891,N_14671,N_14630);
and U14892 (N_14892,N_14564,N_14673);
and U14893 (N_14893,N_14574,N_14647);
and U14894 (N_14894,N_14668,N_14590);
nand U14895 (N_14895,N_14688,N_14586);
nor U14896 (N_14896,N_14548,N_14745);
and U14897 (N_14897,N_14591,N_14548);
nor U14898 (N_14898,N_14667,N_14721);
and U14899 (N_14899,N_14590,N_14564);
or U14900 (N_14900,N_14674,N_14555);
xnor U14901 (N_14901,N_14704,N_14694);
and U14902 (N_14902,N_14668,N_14509);
nand U14903 (N_14903,N_14556,N_14731);
or U14904 (N_14904,N_14734,N_14652);
nand U14905 (N_14905,N_14660,N_14678);
nor U14906 (N_14906,N_14500,N_14693);
xor U14907 (N_14907,N_14540,N_14708);
or U14908 (N_14908,N_14679,N_14719);
and U14909 (N_14909,N_14726,N_14669);
xnor U14910 (N_14910,N_14661,N_14653);
or U14911 (N_14911,N_14508,N_14652);
and U14912 (N_14912,N_14736,N_14533);
and U14913 (N_14913,N_14551,N_14684);
or U14914 (N_14914,N_14606,N_14507);
nor U14915 (N_14915,N_14625,N_14722);
and U14916 (N_14916,N_14618,N_14610);
nand U14917 (N_14917,N_14697,N_14680);
nand U14918 (N_14918,N_14649,N_14621);
or U14919 (N_14919,N_14518,N_14567);
or U14920 (N_14920,N_14620,N_14577);
or U14921 (N_14921,N_14630,N_14625);
or U14922 (N_14922,N_14582,N_14578);
and U14923 (N_14923,N_14574,N_14635);
nor U14924 (N_14924,N_14676,N_14596);
nand U14925 (N_14925,N_14502,N_14656);
nor U14926 (N_14926,N_14668,N_14635);
or U14927 (N_14927,N_14616,N_14614);
and U14928 (N_14928,N_14650,N_14746);
nand U14929 (N_14929,N_14625,N_14683);
xor U14930 (N_14930,N_14567,N_14561);
and U14931 (N_14931,N_14668,N_14707);
or U14932 (N_14932,N_14623,N_14697);
nor U14933 (N_14933,N_14738,N_14626);
nor U14934 (N_14934,N_14597,N_14682);
nor U14935 (N_14935,N_14593,N_14717);
and U14936 (N_14936,N_14717,N_14589);
and U14937 (N_14937,N_14571,N_14551);
nor U14938 (N_14938,N_14673,N_14643);
nand U14939 (N_14939,N_14706,N_14733);
and U14940 (N_14940,N_14641,N_14665);
nor U14941 (N_14941,N_14744,N_14679);
and U14942 (N_14942,N_14541,N_14706);
xor U14943 (N_14943,N_14505,N_14612);
or U14944 (N_14944,N_14555,N_14700);
nor U14945 (N_14945,N_14526,N_14566);
and U14946 (N_14946,N_14670,N_14673);
nand U14947 (N_14947,N_14526,N_14624);
nor U14948 (N_14948,N_14583,N_14630);
nor U14949 (N_14949,N_14545,N_14725);
nand U14950 (N_14950,N_14715,N_14595);
nand U14951 (N_14951,N_14622,N_14706);
and U14952 (N_14952,N_14602,N_14550);
nand U14953 (N_14953,N_14740,N_14716);
or U14954 (N_14954,N_14732,N_14556);
xor U14955 (N_14955,N_14727,N_14547);
and U14956 (N_14956,N_14662,N_14682);
and U14957 (N_14957,N_14558,N_14577);
nor U14958 (N_14958,N_14718,N_14621);
nor U14959 (N_14959,N_14679,N_14702);
and U14960 (N_14960,N_14502,N_14653);
xor U14961 (N_14961,N_14559,N_14640);
or U14962 (N_14962,N_14725,N_14575);
nand U14963 (N_14963,N_14528,N_14717);
xnor U14964 (N_14964,N_14695,N_14625);
or U14965 (N_14965,N_14656,N_14653);
or U14966 (N_14966,N_14567,N_14621);
nor U14967 (N_14967,N_14674,N_14568);
or U14968 (N_14968,N_14705,N_14613);
nor U14969 (N_14969,N_14527,N_14555);
nor U14970 (N_14970,N_14589,N_14520);
nand U14971 (N_14971,N_14721,N_14617);
nor U14972 (N_14972,N_14576,N_14559);
nor U14973 (N_14973,N_14722,N_14506);
xnor U14974 (N_14974,N_14534,N_14529);
nor U14975 (N_14975,N_14534,N_14516);
nor U14976 (N_14976,N_14617,N_14679);
nand U14977 (N_14977,N_14677,N_14725);
or U14978 (N_14978,N_14658,N_14651);
nor U14979 (N_14979,N_14523,N_14535);
nor U14980 (N_14980,N_14644,N_14643);
and U14981 (N_14981,N_14551,N_14654);
nor U14982 (N_14982,N_14746,N_14501);
nor U14983 (N_14983,N_14743,N_14547);
and U14984 (N_14984,N_14706,N_14593);
or U14985 (N_14985,N_14570,N_14506);
xnor U14986 (N_14986,N_14620,N_14593);
nand U14987 (N_14987,N_14721,N_14671);
nand U14988 (N_14988,N_14661,N_14523);
and U14989 (N_14989,N_14689,N_14666);
xor U14990 (N_14990,N_14520,N_14649);
or U14991 (N_14991,N_14662,N_14570);
nor U14992 (N_14992,N_14611,N_14555);
nor U14993 (N_14993,N_14569,N_14545);
nand U14994 (N_14994,N_14596,N_14633);
nor U14995 (N_14995,N_14742,N_14743);
nand U14996 (N_14996,N_14567,N_14549);
nand U14997 (N_14997,N_14743,N_14558);
nor U14998 (N_14998,N_14712,N_14739);
nand U14999 (N_14999,N_14707,N_14583);
or UO_0 (O_0,N_14807,N_14823);
and UO_1 (O_1,N_14850,N_14934);
xor UO_2 (O_2,N_14930,N_14861);
or UO_3 (O_3,N_14775,N_14926);
nand UO_4 (O_4,N_14827,N_14868);
nor UO_5 (O_5,N_14858,N_14853);
nor UO_6 (O_6,N_14952,N_14776);
and UO_7 (O_7,N_14997,N_14919);
and UO_8 (O_8,N_14855,N_14838);
nand UO_9 (O_9,N_14943,N_14866);
and UO_10 (O_10,N_14797,N_14785);
nand UO_11 (O_11,N_14802,N_14774);
nand UO_12 (O_12,N_14801,N_14949);
or UO_13 (O_13,N_14968,N_14900);
and UO_14 (O_14,N_14769,N_14878);
xor UO_15 (O_15,N_14799,N_14892);
nand UO_16 (O_16,N_14831,N_14989);
xor UO_17 (O_17,N_14933,N_14773);
nand UO_18 (O_18,N_14996,N_14864);
nand UO_19 (O_19,N_14800,N_14992);
and UO_20 (O_20,N_14795,N_14834);
nor UO_21 (O_21,N_14925,N_14995);
nand UO_22 (O_22,N_14862,N_14915);
xor UO_23 (O_23,N_14879,N_14907);
nor UO_24 (O_24,N_14824,N_14993);
nor UO_25 (O_25,N_14828,N_14813);
or UO_26 (O_26,N_14948,N_14890);
or UO_27 (O_27,N_14778,N_14811);
and UO_28 (O_28,N_14984,N_14896);
nor UO_29 (O_29,N_14931,N_14897);
nor UO_30 (O_30,N_14846,N_14825);
and UO_31 (O_31,N_14793,N_14920);
and UO_32 (O_32,N_14945,N_14760);
xnor UO_33 (O_33,N_14967,N_14912);
nor UO_34 (O_34,N_14821,N_14937);
and UO_35 (O_35,N_14780,N_14901);
nor UO_36 (O_36,N_14922,N_14941);
and UO_37 (O_37,N_14911,N_14960);
xnor UO_38 (O_38,N_14833,N_14979);
and UO_39 (O_39,N_14781,N_14765);
and UO_40 (O_40,N_14750,N_14805);
nand UO_41 (O_41,N_14990,N_14756);
or UO_42 (O_42,N_14779,N_14757);
nor UO_43 (O_43,N_14875,N_14786);
xor UO_44 (O_44,N_14763,N_14998);
nor UO_45 (O_45,N_14830,N_14815);
and UO_46 (O_46,N_14857,N_14905);
nor UO_47 (O_47,N_14891,N_14810);
and UO_48 (O_48,N_14856,N_14782);
xnor UO_49 (O_49,N_14955,N_14944);
nand UO_50 (O_50,N_14964,N_14963);
nor UO_51 (O_51,N_14942,N_14822);
and UO_52 (O_52,N_14909,N_14953);
or UO_53 (O_53,N_14806,N_14788);
xor UO_54 (O_54,N_14870,N_14991);
xnor UO_55 (O_55,N_14917,N_14804);
nand UO_56 (O_56,N_14983,N_14816);
and UO_57 (O_57,N_14938,N_14843);
xor UO_58 (O_58,N_14887,N_14839);
or UO_59 (O_59,N_14777,N_14819);
or UO_60 (O_60,N_14874,N_14977);
and UO_61 (O_61,N_14969,N_14783);
and UO_62 (O_62,N_14910,N_14986);
nand UO_63 (O_63,N_14794,N_14761);
or UO_64 (O_64,N_14842,N_14840);
nand UO_65 (O_65,N_14921,N_14913);
nor UO_66 (O_66,N_14904,N_14906);
nor UO_67 (O_67,N_14882,N_14981);
or UO_68 (O_68,N_14994,N_14884);
or UO_69 (O_69,N_14820,N_14865);
nand UO_70 (O_70,N_14764,N_14927);
xnor UO_71 (O_71,N_14852,N_14766);
nor UO_72 (O_72,N_14872,N_14835);
and UO_73 (O_73,N_14869,N_14950);
and UO_74 (O_74,N_14908,N_14784);
xnor UO_75 (O_75,N_14768,N_14848);
and UO_76 (O_76,N_14854,N_14947);
nand UO_77 (O_77,N_14936,N_14894);
or UO_78 (O_78,N_14791,N_14787);
and UO_79 (O_79,N_14898,N_14972);
and UO_80 (O_80,N_14836,N_14974);
xor UO_81 (O_81,N_14889,N_14899);
nand UO_82 (O_82,N_14754,N_14863);
nor UO_83 (O_83,N_14770,N_14888);
nor UO_84 (O_84,N_14867,N_14790);
and UO_85 (O_85,N_14812,N_14946);
nand UO_86 (O_86,N_14847,N_14923);
or UO_87 (O_87,N_14829,N_14767);
nand UO_88 (O_88,N_14924,N_14753);
and UO_89 (O_89,N_14959,N_14832);
and UO_90 (O_90,N_14956,N_14814);
xor UO_91 (O_91,N_14849,N_14916);
nand UO_92 (O_92,N_14975,N_14962);
and UO_93 (O_93,N_14928,N_14859);
nor UO_94 (O_94,N_14803,N_14751);
and UO_95 (O_95,N_14957,N_14885);
nor UO_96 (O_96,N_14762,N_14789);
nor UO_97 (O_97,N_14893,N_14973);
nor UO_98 (O_98,N_14903,N_14954);
nor UO_99 (O_99,N_14966,N_14980);
and UO_100 (O_100,N_14932,N_14965);
or UO_101 (O_101,N_14841,N_14873);
xnor UO_102 (O_102,N_14939,N_14771);
nor UO_103 (O_103,N_14877,N_14798);
nor UO_104 (O_104,N_14987,N_14940);
nand UO_105 (O_105,N_14971,N_14837);
xnor UO_106 (O_106,N_14918,N_14929);
nor UO_107 (O_107,N_14759,N_14758);
nor UO_108 (O_108,N_14961,N_14792);
and UO_109 (O_109,N_14880,N_14755);
and UO_110 (O_110,N_14976,N_14876);
nand UO_111 (O_111,N_14985,N_14982);
nor UO_112 (O_112,N_14844,N_14845);
nor UO_113 (O_113,N_14817,N_14752);
and UO_114 (O_114,N_14818,N_14772);
nor UO_115 (O_115,N_14978,N_14826);
xnor UO_116 (O_116,N_14871,N_14914);
and UO_117 (O_117,N_14951,N_14970);
and UO_118 (O_118,N_14796,N_14881);
xor UO_119 (O_119,N_14883,N_14809);
nor UO_120 (O_120,N_14851,N_14935);
nand UO_121 (O_121,N_14988,N_14902);
and UO_122 (O_122,N_14999,N_14808);
and UO_123 (O_123,N_14958,N_14860);
nor UO_124 (O_124,N_14895,N_14886);
and UO_125 (O_125,N_14767,N_14990);
or UO_126 (O_126,N_14838,N_14928);
and UO_127 (O_127,N_14865,N_14756);
xnor UO_128 (O_128,N_14867,N_14847);
nand UO_129 (O_129,N_14971,N_14995);
and UO_130 (O_130,N_14814,N_14998);
nand UO_131 (O_131,N_14760,N_14904);
or UO_132 (O_132,N_14957,N_14851);
and UO_133 (O_133,N_14852,N_14997);
or UO_134 (O_134,N_14815,N_14970);
xor UO_135 (O_135,N_14804,N_14805);
or UO_136 (O_136,N_14946,N_14887);
nor UO_137 (O_137,N_14883,N_14811);
and UO_138 (O_138,N_14975,N_14815);
nand UO_139 (O_139,N_14821,N_14784);
and UO_140 (O_140,N_14840,N_14781);
and UO_141 (O_141,N_14852,N_14787);
and UO_142 (O_142,N_14818,N_14941);
or UO_143 (O_143,N_14936,N_14960);
and UO_144 (O_144,N_14827,N_14898);
and UO_145 (O_145,N_14809,N_14781);
and UO_146 (O_146,N_14826,N_14939);
xor UO_147 (O_147,N_14973,N_14920);
and UO_148 (O_148,N_14941,N_14983);
nor UO_149 (O_149,N_14811,N_14823);
nand UO_150 (O_150,N_14865,N_14844);
xor UO_151 (O_151,N_14769,N_14858);
nor UO_152 (O_152,N_14824,N_14866);
or UO_153 (O_153,N_14977,N_14763);
and UO_154 (O_154,N_14938,N_14772);
xnor UO_155 (O_155,N_14905,N_14922);
and UO_156 (O_156,N_14792,N_14968);
nand UO_157 (O_157,N_14796,N_14934);
nor UO_158 (O_158,N_14836,N_14959);
or UO_159 (O_159,N_14959,N_14750);
and UO_160 (O_160,N_14933,N_14924);
or UO_161 (O_161,N_14990,N_14988);
and UO_162 (O_162,N_14902,N_14867);
or UO_163 (O_163,N_14835,N_14935);
nor UO_164 (O_164,N_14882,N_14874);
or UO_165 (O_165,N_14882,N_14869);
nand UO_166 (O_166,N_14977,N_14836);
and UO_167 (O_167,N_14862,N_14917);
nor UO_168 (O_168,N_14839,N_14840);
nand UO_169 (O_169,N_14948,N_14930);
nand UO_170 (O_170,N_14800,N_14761);
xnor UO_171 (O_171,N_14771,N_14843);
nand UO_172 (O_172,N_14890,N_14928);
or UO_173 (O_173,N_14767,N_14855);
nor UO_174 (O_174,N_14948,N_14831);
nand UO_175 (O_175,N_14981,N_14953);
xor UO_176 (O_176,N_14907,N_14945);
nand UO_177 (O_177,N_14930,N_14834);
and UO_178 (O_178,N_14872,N_14828);
nor UO_179 (O_179,N_14901,N_14772);
and UO_180 (O_180,N_14825,N_14802);
xnor UO_181 (O_181,N_14917,N_14913);
or UO_182 (O_182,N_14837,N_14874);
or UO_183 (O_183,N_14816,N_14845);
nor UO_184 (O_184,N_14809,N_14821);
nor UO_185 (O_185,N_14978,N_14848);
nand UO_186 (O_186,N_14958,N_14816);
nor UO_187 (O_187,N_14877,N_14998);
xor UO_188 (O_188,N_14790,N_14753);
nand UO_189 (O_189,N_14806,N_14999);
nand UO_190 (O_190,N_14789,N_14830);
nand UO_191 (O_191,N_14974,N_14803);
nand UO_192 (O_192,N_14800,N_14935);
or UO_193 (O_193,N_14784,N_14859);
nor UO_194 (O_194,N_14973,N_14932);
xor UO_195 (O_195,N_14923,N_14839);
nor UO_196 (O_196,N_14920,N_14864);
or UO_197 (O_197,N_14873,N_14883);
or UO_198 (O_198,N_14923,N_14902);
nand UO_199 (O_199,N_14975,N_14770);
nand UO_200 (O_200,N_14832,N_14753);
nor UO_201 (O_201,N_14955,N_14954);
or UO_202 (O_202,N_14972,N_14822);
and UO_203 (O_203,N_14857,N_14919);
and UO_204 (O_204,N_14993,N_14983);
or UO_205 (O_205,N_14971,N_14917);
nor UO_206 (O_206,N_14874,N_14893);
nand UO_207 (O_207,N_14905,N_14923);
nor UO_208 (O_208,N_14924,N_14758);
nor UO_209 (O_209,N_14858,N_14865);
or UO_210 (O_210,N_14784,N_14959);
and UO_211 (O_211,N_14938,N_14863);
or UO_212 (O_212,N_14825,N_14768);
nor UO_213 (O_213,N_14967,N_14818);
or UO_214 (O_214,N_14914,N_14805);
and UO_215 (O_215,N_14811,N_14976);
xor UO_216 (O_216,N_14923,N_14981);
and UO_217 (O_217,N_14920,N_14788);
and UO_218 (O_218,N_14950,N_14966);
or UO_219 (O_219,N_14807,N_14805);
and UO_220 (O_220,N_14945,N_14811);
xnor UO_221 (O_221,N_14906,N_14840);
and UO_222 (O_222,N_14968,N_14925);
nor UO_223 (O_223,N_14826,N_14782);
nand UO_224 (O_224,N_14756,N_14937);
nand UO_225 (O_225,N_14963,N_14928);
nor UO_226 (O_226,N_14765,N_14800);
nor UO_227 (O_227,N_14790,N_14961);
or UO_228 (O_228,N_14890,N_14994);
and UO_229 (O_229,N_14852,N_14834);
or UO_230 (O_230,N_14961,N_14903);
and UO_231 (O_231,N_14777,N_14861);
nand UO_232 (O_232,N_14804,N_14897);
nor UO_233 (O_233,N_14775,N_14972);
nand UO_234 (O_234,N_14893,N_14872);
or UO_235 (O_235,N_14905,N_14827);
and UO_236 (O_236,N_14923,N_14990);
nand UO_237 (O_237,N_14959,N_14909);
or UO_238 (O_238,N_14824,N_14784);
xor UO_239 (O_239,N_14953,N_14911);
nand UO_240 (O_240,N_14907,N_14987);
nand UO_241 (O_241,N_14806,N_14885);
or UO_242 (O_242,N_14778,N_14927);
nor UO_243 (O_243,N_14962,N_14973);
nand UO_244 (O_244,N_14784,N_14883);
nand UO_245 (O_245,N_14890,N_14844);
and UO_246 (O_246,N_14909,N_14995);
nor UO_247 (O_247,N_14777,N_14892);
or UO_248 (O_248,N_14761,N_14818);
nand UO_249 (O_249,N_14864,N_14874);
nor UO_250 (O_250,N_14806,N_14784);
and UO_251 (O_251,N_14839,N_14924);
nor UO_252 (O_252,N_14940,N_14892);
nand UO_253 (O_253,N_14812,N_14847);
or UO_254 (O_254,N_14906,N_14778);
xnor UO_255 (O_255,N_14947,N_14805);
or UO_256 (O_256,N_14872,N_14915);
nor UO_257 (O_257,N_14898,N_14938);
xor UO_258 (O_258,N_14913,N_14762);
nor UO_259 (O_259,N_14838,N_14982);
nand UO_260 (O_260,N_14825,N_14898);
or UO_261 (O_261,N_14793,N_14750);
and UO_262 (O_262,N_14756,N_14787);
nand UO_263 (O_263,N_14811,N_14953);
nor UO_264 (O_264,N_14843,N_14891);
nand UO_265 (O_265,N_14990,N_14779);
and UO_266 (O_266,N_14922,N_14768);
and UO_267 (O_267,N_14911,N_14933);
or UO_268 (O_268,N_14983,N_14761);
nand UO_269 (O_269,N_14919,N_14864);
xor UO_270 (O_270,N_14999,N_14924);
or UO_271 (O_271,N_14857,N_14775);
nand UO_272 (O_272,N_14839,N_14834);
nand UO_273 (O_273,N_14902,N_14750);
nand UO_274 (O_274,N_14778,N_14963);
or UO_275 (O_275,N_14906,N_14917);
or UO_276 (O_276,N_14992,N_14873);
nand UO_277 (O_277,N_14837,N_14919);
nand UO_278 (O_278,N_14782,N_14974);
nor UO_279 (O_279,N_14918,N_14870);
nor UO_280 (O_280,N_14899,N_14855);
xor UO_281 (O_281,N_14762,N_14963);
and UO_282 (O_282,N_14838,N_14947);
nor UO_283 (O_283,N_14828,N_14926);
nand UO_284 (O_284,N_14993,N_14882);
and UO_285 (O_285,N_14998,N_14759);
nand UO_286 (O_286,N_14964,N_14886);
and UO_287 (O_287,N_14762,N_14927);
nand UO_288 (O_288,N_14946,N_14917);
and UO_289 (O_289,N_14930,N_14887);
nor UO_290 (O_290,N_14902,N_14948);
and UO_291 (O_291,N_14930,N_14949);
nor UO_292 (O_292,N_14829,N_14887);
nand UO_293 (O_293,N_14752,N_14835);
nand UO_294 (O_294,N_14908,N_14969);
and UO_295 (O_295,N_14942,N_14989);
nor UO_296 (O_296,N_14971,N_14885);
or UO_297 (O_297,N_14782,N_14825);
and UO_298 (O_298,N_14846,N_14864);
and UO_299 (O_299,N_14809,N_14832);
and UO_300 (O_300,N_14836,N_14759);
xor UO_301 (O_301,N_14881,N_14845);
xnor UO_302 (O_302,N_14835,N_14838);
or UO_303 (O_303,N_14941,N_14974);
and UO_304 (O_304,N_14838,N_14939);
and UO_305 (O_305,N_14781,N_14913);
nor UO_306 (O_306,N_14961,N_14751);
and UO_307 (O_307,N_14908,N_14971);
xnor UO_308 (O_308,N_14972,N_14940);
nor UO_309 (O_309,N_14837,N_14877);
xnor UO_310 (O_310,N_14916,N_14831);
and UO_311 (O_311,N_14855,N_14882);
nor UO_312 (O_312,N_14813,N_14838);
and UO_313 (O_313,N_14880,N_14813);
and UO_314 (O_314,N_14889,N_14853);
xor UO_315 (O_315,N_14784,N_14944);
nand UO_316 (O_316,N_14798,N_14860);
nand UO_317 (O_317,N_14942,N_14930);
xnor UO_318 (O_318,N_14886,N_14917);
and UO_319 (O_319,N_14752,N_14945);
nor UO_320 (O_320,N_14822,N_14873);
nand UO_321 (O_321,N_14927,N_14934);
and UO_322 (O_322,N_14893,N_14821);
nor UO_323 (O_323,N_14900,N_14948);
or UO_324 (O_324,N_14764,N_14956);
and UO_325 (O_325,N_14796,N_14879);
or UO_326 (O_326,N_14802,N_14875);
nor UO_327 (O_327,N_14780,N_14796);
or UO_328 (O_328,N_14899,N_14904);
nor UO_329 (O_329,N_14756,N_14907);
xor UO_330 (O_330,N_14769,N_14935);
and UO_331 (O_331,N_14827,N_14775);
and UO_332 (O_332,N_14801,N_14902);
nand UO_333 (O_333,N_14989,N_14779);
nor UO_334 (O_334,N_14957,N_14784);
xor UO_335 (O_335,N_14951,N_14998);
nor UO_336 (O_336,N_14862,N_14976);
nand UO_337 (O_337,N_14987,N_14889);
xnor UO_338 (O_338,N_14937,N_14773);
and UO_339 (O_339,N_14856,N_14959);
xnor UO_340 (O_340,N_14981,N_14751);
nor UO_341 (O_341,N_14774,N_14948);
nand UO_342 (O_342,N_14958,N_14791);
and UO_343 (O_343,N_14951,N_14923);
xnor UO_344 (O_344,N_14948,N_14856);
xor UO_345 (O_345,N_14950,N_14927);
nor UO_346 (O_346,N_14780,N_14903);
or UO_347 (O_347,N_14866,N_14962);
nand UO_348 (O_348,N_14841,N_14981);
nand UO_349 (O_349,N_14787,N_14817);
nor UO_350 (O_350,N_14953,N_14946);
xnor UO_351 (O_351,N_14931,N_14782);
nand UO_352 (O_352,N_14787,N_14895);
xnor UO_353 (O_353,N_14919,N_14826);
nor UO_354 (O_354,N_14888,N_14808);
nor UO_355 (O_355,N_14847,N_14897);
and UO_356 (O_356,N_14893,N_14772);
and UO_357 (O_357,N_14822,N_14839);
nor UO_358 (O_358,N_14779,N_14796);
and UO_359 (O_359,N_14776,N_14821);
nor UO_360 (O_360,N_14775,N_14820);
and UO_361 (O_361,N_14997,N_14827);
nand UO_362 (O_362,N_14870,N_14932);
and UO_363 (O_363,N_14862,N_14965);
and UO_364 (O_364,N_14758,N_14751);
and UO_365 (O_365,N_14930,N_14917);
nand UO_366 (O_366,N_14991,N_14913);
nand UO_367 (O_367,N_14923,N_14948);
and UO_368 (O_368,N_14864,N_14924);
nor UO_369 (O_369,N_14939,N_14985);
nand UO_370 (O_370,N_14894,N_14766);
xor UO_371 (O_371,N_14844,N_14828);
nand UO_372 (O_372,N_14866,N_14897);
nor UO_373 (O_373,N_14883,N_14978);
nand UO_374 (O_374,N_14955,N_14846);
xnor UO_375 (O_375,N_14941,N_14886);
and UO_376 (O_376,N_14765,N_14758);
nand UO_377 (O_377,N_14996,N_14909);
nor UO_378 (O_378,N_14805,N_14840);
or UO_379 (O_379,N_14876,N_14750);
nand UO_380 (O_380,N_14925,N_14967);
and UO_381 (O_381,N_14785,N_14990);
and UO_382 (O_382,N_14963,N_14879);
and UO_383 (O_383,N_14972,N_14939);
and UO_384 (O_384,N_14779,N_14750);
nand UO_385 (O_385,N_14868,N_14956);
and UO_386 (O_386,N_14842,N_14948);
and UO_387 (O_387,N_14757,N_14992);
xor UO_388 (O_388,N_14841,N_14814);
and UO_389 (O_389,N_14822,N_14831);
or UO_390 (O_390,N_14947,N_14787);
nand UO_391 (O_391,N_14932,N_14776);
and UO_392 (O_392,N_14884,N_14827);
and UO_393 (O_393,N_14876,N_14828);
and UO_394 (O_394,N_14777,N_14833);
and UO_395 (O_395,N_14907,N_14894);
nand UO_396 (O_396,N_14818,N_14954);
or UO_397 (O_397,N_14779,N_14857);
or UO_398 (O_398,N_14756,N_14982);
nand UO_399 (O_399,N_14770,N_14943);
nand UO_400 (O_400,N_14975,N_14894);
or UO_401 (O_401,N_14995,N_14956);
and UO_402 (O_402,N_14848,N_14754);
nor UO_403 (O_403,N_14942,N_14859);
or UO_404 (O_404,N_14984,N_14844);
nor UO_405 (O_405,N_14867,N_14805);
and UO_406 (O_406,N_14921,N_14763);
and UO_407 (O_407,N_14953,N_14914);
and UO_408 (O_408,N_14800,N_14802);
and UO_409 (O_409,N_14774,N_14854);
nor UO_410 (O_410,N_14834,N_14810);
xor UO_411 (O_411,N_14755,N_14783);
and UO_412 (O_412,N_14946,N_14888);
nand UO_413 (O_413,N_14899,N_14992);
xnor UO_414 (O_414,N_14958,N_14903);
nand UO_415 (O_415,N_14854,N_14876);
and UO_416 (O_416,N_14777,N_14883);
and UO_417 (O_417,N_14803,N_14938);
and UO_418 (O_418,N_14961,N_14989);
nor UO_419 (O_419,N_14891,N_14836);
or UO_420 (O_420,N_14852,N_14871);
nand UO_421 (O_421,N_14789,N_14900);
or UO_422 (O_422,N_14830,N_14868);
or UO_423 (O_423,N_14854,N_14949);
nand UO_424 (O_424,N_14822,N_14963);
nand UO_425 (O_425,N_14899,N_14769);
and UO_426 (O_426,N_14801,N_14893);
nand UO_427 (O_427,N_14896,N_14795);
nor UO_428 (O_428,N_14791,N_14911);
xnor UO_429 (O_429,N_14982,N_14899);
nor UO_430 (O_430,N_14993,N_14767);
or UO_431 (O_431,N_14885,N_14974);
or UO_432 (O_432,N_14825,N_14961);
and UO_433 (O_433,N_14922,N_14802);
xor UO_434 (O_434,N_14754,N_14955);
nor UO_435 (O_435,N_14855,N_14869);
nor UO_436 (O_436,N_14884,N_14778);
nand UO_437 (O_437,N_14775,N_14998);
nand UO_438 (O_438,N_14776,N_14877);
xnor UO_439 (O_439,N_14769,N_14865);
nand UO_440 (O_440,N_14825,N_14943);
or UO_441 (O_441,N_14755,N_14832);
or UO_442 (O_442,N_14849,N_14992);
xnor UO_443 (O_443,N_14831,N_14961);
and UO_444 (O_444,N_14895,N_14891);
nand UO_445 (O_445,N_14771,N_14965);
or UO_446 (O_446,N_14832,N_14817);
nor UO_447 (O_447,N_14903,N_14813);
and UO_448 (O_448,N_14804,N_14857);
nand UO_449 (O_449,N_14937,N_14762);
or UO_450 (O_450,N_14913,N_14969);
and UO_451 (O_451,N_14752,N_14972);
nor UO_452 (O_452,N_14893,N_14890);
and UO_453 (O_453,N_14793,N_14783);
or UO_454 (O_454,N_14925,N_14778);
and UO_455 (O_455,N_14785,N_14772);
and UO_456 (O_456,N_14765,N_14836);
nand UO_457 (O_457,N_14973,N_14850);
nor UO_458 (O_458,N_14787,N_14930);
and UO_459 (O_459,N_14803,N_14950);
nand UO_460 (O_460,N_14873,N_14756);
nand UO_461 (O_461,N_14764,N_14878);
and UO_462 (O_462,N_14757,N_14962);
xor UO_463 (O_463,N_14923,N_14854);
or UO_464 (O_464,N_14975,N_14969);
nor UO_465 (O_465,N_14939,N_14943);
and UO_466 (O_466,N_14858,N_14915);
nor UO_467 (O_467,N_14995,N_14804);
nand UO_468 (O_468,N_14848,N_14795);
or UO_469 (O_469,N_14819,N_14991);
nor UO_470 (O_470,N_14840,N_14831);
xor UO_471 (O_471,N_14986,N_14940);
nand UO_472 (O_472,N_14756,N_14969);
or UO_473 (O_473,N_14924,N_14879);
and UO_474 (O_474,N_14958,N_14761);
and UO_475 (O_475,N_14804,N_14757);
nand UO_476 (O_476,N_14945,N_14842);
or UO_477 (O_477,N_14779,N_14944);
nor UO_478 (O_478,N_14966,N_14762);
or UO_479 (O_479,N_14753,N_14928);
and UO_480 (O_480,N_14780,N_14867);
xnor UO_481 (O_481,N_14942,N_14780);
nand UO_482 (O_482,N_14885,N_14789);
or UO_483 (O_483,N_14795,N_14760);
or UO_484 (O_484,N_14965,N_14925);
xor UO_485 (O_485,N_14894,N_14913);
and UO_486 (O_486,N_14861,N_14878);
nor UO_487 (O_487,N_14826,N_14772);
nand UO_488 (O_488,N_14911,N_14857);
nand UO_489 (O_489,N_14980,N_14897);
nand UO_490 (O_490,N_14780,N_14940);
nor UO_491 (O_491,N_14810,N_14938);
or UO_492 (O_492,N_14941,N_14945);
and UO_493 (O_493,N_14960,N_14789);
nor UO_494 (O_494,N_14994,N_14818);
nand UO_495 (O_495,N_14756,N_14939);
xor UO_496 (O_496,N_14814,N_14933);
nor UO_497 (O_497,N_14793,N_14854);
nor UO_498 (O_498,N_14931,N_14945);
nand UO_499 (O_499,N_14839,N_14855);
xnor UO_500 (O_500,N_14768,N_14751);
nand UO_501 (O_501,N_14901,N_14797);
nand UO_502 (O_502,N_14983,N_14970);
and UO_503 (O_503,N_14975,N_14964);
and UO_504 (O_504,N_14851,N_14925);
nor UO_505 (O_505,N_14992,N_14775);
xor UO_506 (O_506,N_14958,N_14949);
nor UO_507 (O_507,N_14874,N_14796);
nor UO_508 (O_508,N_14822,N_14905);
or UO_509 (O_509,N_14882,N_14913);
and UO_510 (O_510,N_14761,N_14972);
nand UO_511 (O_511,N_14932,N_14802);
xnor UO_512 (O_512,N_14754,N_14924);
nor UO_513 (O_513,N_14979,N_14753);
xnor UO_514 (O_514,N_14884,N_14791);
or UO_515 (O_515,N_14913,N_14979);
xnor UO_516 (O_516,N_14826,N_14890);
nand UO_517 (O_517,N_14887,N_14775);
nor UO_518 (O_518,N_14992,N_14833);
and UO_519 (O_519,N_14782,N_14821);
nand UO_520 (O_520,N_14978,N_14965);
nor UO_521 (O_521,N_14969,N_14843);
and UO_522 (O_522,N_14820,N_14918);
xnor UO_523 (O_523,N_14931,N_14920);
and UO_524 (O_524,N_14908,N_14859);
or UO_525 (O_525,N_14978,N_14957);
and UO_526 (O_526,N_14851,N_14850);
nand UO_527 (O_527,N_14870,N_14905);
xor UO_528 (O_528,N_14938,N_14935);
nand UO_529 (O_529,N_14796,N_14790);
and UO_530 (O_530,N_14878,N_14840);
or UO_531 (O_531,N_14938,N_14834);
xnor UO_532 (O_532,N_14931,N_14844);
nand UO_533 (O_533,N_14974,N_14899);
nor UO_534 (O_534,N_14971,N_14782);
and UO_535 (O_535,N_14902,N_14918);
and UO_536 (O_536,N_14801,N_14948);
nand UO_537 (O_537,N_14892,N_14780);
nor UO_538 (O_538,N_14934,N_14907);
and UO_539 (O_539,N_14884,N_14765);
and UO_540 (O_540,N_14958,N_14822);
and UO_541 (O_541,N_14780,N_14794);
nand UO_542 (O_542,N_14791,N_14821);
nand UO_543 (O_543,N_14834,N_14961);
nor UO_544 (O_544,N_14924,N_14874);
nand UO_545 (O_545,N_14823,N_14853);
and UO_546 (O_546,N_14786,N_14985);
nand UO_547 (O_547,N_14942,N_14751);
nand UO_548 (O_548,N_14928,N_14912);
nand UO_549 (O_549,N_14801,N_14797);
xor UO_550 (O_550,N_14752,N_14922);
nand UO_551 (O_551,N_14962,N_14928);
nand UO_552 (O_552,N_14756,N_14981);
and UO_553 (O_553,N_14805,N_14787);
nor UO_554 (O_554,N_14970,N_14817);
or UO_555 (O_555,N_14967,N_14814);
or UO_556 (O_556,N_14954,N_14833);
or UO_557 (O_557,N_14761,N_14883);
nand UO_558 (O_558,N_14902,N_14950);
nor UO_559 (O_559,N_14834,N_14945);
or UO_560 (O_560,N_14965,N_14816);
nand UO_561 (O_561,N_14792,N_14984);
xor UO_562 (O_562,N_14819,N_14962);
nor UO_563 (O_563,N_14903,N_14937);
xor UO_564 (O_564,N_14992,N_14943);
nor UO_565 (O_565,N_14753,N_14996);
nor UO_566 (O_566,N_14799,N_14807);
nor UO_567 (O_567,N_14992,N_14930);
or UO_568 (O_568,N_14777,N_14937);
or UO_569 (O_569,N_14892,N_14802);
or UO_570 (O_570,N_14961,N_14906);
or UO_571 (O_571,N_14927,N_14830);
nor UO_572 (O_572,N_14759,N_14750);
xor UO_573 (O_573,N_14759,N_14989);
nand UO_574 (O_574,N_14906,N_14989);
nor UO_575 (O_575,N_14843,N_14993);
or UO_576 (O_576,N_14932,N_14888);
nand UO_577 (O_577,N_14776,N_14888);
or UO_578 (O_578,N_14913,N_14784);
nand UO_579 (O_579,N_14803,N_14783);
or UO_580 (O_580,N_14841,N_14996);
nor UO_581 (O_581,N_14795,N_14766);
nor UO_582 (O_582,N_14831,N_14862);
or UO_583 (O_583,N_14833,N_14924);
nand UO_584 (O_584,N_14955,N_14761);
or UO_585 (O_585,N_14756,N_14988);
nor UO_586 (O_586,N_14861,N_14789);
and UO_587 (O_587,N_14856,N_14790);
or UO_588 (O_588,N_14975,N_14955);
xor UO_589 (O_589,N_14883,N_14832);
or UO_590 (O_590,N_14764,N_14787);
nand UO_591 (O_591,N_14798,N_14937);
or UO_592 (O_592,N_14940,N_14763);
nand UO_593 (O_593,N_14875,N_14904);
nand UO_594 (O_594,N_14838,N_14798);
or UO_595 (O_595,N_14891,N_14942);
and UO_596 (O_596,N_14847,N_14766);
nand UO_597 (O_597,N_14862,N_14912);
and UO_598 (O_598,N_14999,N_14949);
nand UO_599 (O_599,N_14881,N_14925);
nand UO_600 (O_600,N_14883,N_14807);
nand UO_601 (O_601,N_14904,N_14876);
nand UO_602 (O_602,N_14964,N_14833);
nand UO_603 (O_603,N_14990,N_14894);
nor UO_604 (O_604,N_14785,N_14953);
or UO_605 (O_605,N_14828,N_14989);
nor UO_606 (O_606,N_14870,N_14864);
nand UO_607 (O_607,N_14956,N_14813);
xnor UO_608 (O_608,N_14980,N_14875);
nor UO_609 (O_609,N_14751,N_14772);
nor UO_610 (O_610,N_14797,N_14879);
nor UO_611 (O_611,N_14856,N_14895);
and UO_612 (O_612,N_14868,N_14892);
nand UO_613 (O_613,N_14772,N_14872);
xor UO_614 (O_614,N_14973,N_14846);
xnor UO_615 (O_615,N_14988,N_14996);
nor UO_616 (O_616,N_14926,N_14774);
nand UO_617 (O_617,N_14774,N_14915);
and UO_618 (O_618,N_14783,N_14766);
or UO_619 (O_619,N_14956,N_14819);
and UO_620 (O_620,N_14895,N_14883);
nand UO_621 (O_621,N_14895,N_14919);
xnor UO_622 (O_622,N_14859,N_14884);
xor UO_623 (O_623,N_14798,N_14828);
or UO_624 (O_624,N_14961,N_14770);
nand UO_625 (O_625,N_14850,N_14982);
nor UO_626 (O_626,N_14988,N_14989);
and UO_627 (O_627,N_14870,N_14928);
and UO_628 (O_628,N_14909,N_14791);
and UO_629 (O_629,N_14907,N_14992);
and UO_630 (O_630,N_14855,N_14859);
and UO_631 (O_631,N_14800,N_14996);
nor UO_632 (O_632,N_14915,N_14947);
nand UO_633 (O_633,N_14774,N_14763);
nand UO_634 (O_634,N_14991,N_14871);
and UO_635 (O_635,N_14868,N_14907);
and UO_636 (O_636,N_14883,N_14886);
or UO_637 (O_637,N_14836,N_14990);
nand UO_638 (O_638,N_14912,N_14811);
xnor UO_639 (O_639,N_14843,N_14810);
nor UO_640 (O_640,N_14954,N_14814);
nand UO_641 (O_641,N_14934,N_14916);
nor UO_642 (O_642,N_14943,N_14801);
or UO_643 (O_643,N_14951,N_14815);
nor UO_644 (O_644,N_14995,N_14927);
nor UO_645 (O_645,N_14839,N_14948);
and UO_646 (O_646,N_14783,N_14837);
nand UO_647 (O_647,N_14959,N_14966);
and UO_648 (O_648,N_14808,N_14843);
nor UO_649 (O_649,N_14932,N_14914);
or UO_650 (O_650,N_14796,N_14750);
xnor UO_651 (O_651,N_14830,N_14979);
or UO_652 (O_652,N_14777,N_14869);
nor UO_653 (O_653,N_14792,N_14858);
xor UO_654 (O_654,N_14826,N_14827);
and UO_655 (O_655,N_14899,N_14783);
and UO_656 (O_656,N_14859,N_14854);
nand UO_657 (O_657,N_14839,N_14982);
or UO_658 (O_658,N_14841,N_14879);
and UO_659 (O_659,N_14792,N_14877);
and UO_660 (O_660,N_14777,N_14781);
and UO_661 (O_661,N_14826,N_14947);
or UO_662 (O_662,N_14815,N_14789);
or UO_663 (O_663,N_14885,N_14933);
nor UO_664 (O_664,N_14874,N_14916);
nand UO_665 (O_665,N_14897,N_14953);
and UO_666 (O_666,N_14892,N_14964);
nor UO_667 (O_667,N_14773,N_14983);
or UO_668 (O_668,N_14933,N_14995);
nor UO_669 (O_669,N_14908,N_14842);
nor UO_670 (O_670,N_14830,N_14974);
nand UO_671 (O_671,N_14864,N_14787);
or UO_672 (O_672,N_14797,N_14991);
or UO_673 (O_673,N_14939,N_14862);
nand UO_674 (O_674,N_14957,N_14880);
or UO_675 (O_675,N_14924,N_14824);
nand UO_676 (O_676,N_14855,N_14863);
xnor UO_677 (O_677,N_14800,N_14776);
and UO_678 (O_678,N_14757,N_14760);
or UO_679 (O_679,N_14907,N_14834);
or UO_680 (O_680,N_14833,N_14857);
nor UO_681 (O_681,N_14919,N_14854);
or UO_682 (O_682,N_14790,N_14910);
nor UO_683 (O_683,N_14863,N_14784);
and UO_684 (O_684,N_14990,N_14777);
or UO_685 (O_685,N_14932,N_14899);
nand UO_686 (O_686,N_14894,N_14984);
and UO_687 (O_687,N_14808,N_14818);
nand UO_688 (O_688,N_14949,N_14765);
nand UO_689 (O_689,N_14990,N_14753);
or UO_690 (O_690,N_14768,N_14759);
xnor UO_691 (O_691,N_14970,N_14777);
and UO_692 (O_692,N_14986,N_14819);
nand UO_693 (O_693,N_14775,N_14907);
nor UO_694 (O_694,N_14840,N_14923);
xor UO_695 (O_695,N_14923,N_14920);
and UO_696 (O_696,N_14766,N_14844);
nand UO_697 (O_697,N_14871,N_14940);
and UO_698 (O_698,N_14882,N_14927);
nand UO_699 (O_699,N_14885,N_14954);
or UO_700 (O_700,N_14898,N_14840);
or UO_701 (O_701,N_14765,N_14915);
nor UO_702 (O_702,N_14824,N_14885);
nand UO_703 (O_703,N_14768,N_14761);
nor UO_704 (O_704,N_14969,N_14976);
nand UO_705 (O_705,N_14921,N_14894);
nor UO_706 (O_706,N_14974,N_14770);
nand UO_707 (O_707,N_14932,N_14904);
nand UO_708 (O_708,N_14857,N_14898);
and UO_709 (O_709,N_14887,N_14779);
and UO_710 (O_710,N_14985,N_14948);
nor UO_711 (O_711,N_14892,N_14905);
nor UO_712 (O_712,N_14785,N_14876);
nand UO_713 (O_713,N_14883,N_14868);
or UO_714 (O_714,N_14764,N_14875);
and UO_715 (O_715,N_14771,N_14784);
nand UO_716 (O_716,N_14840,N_14877);
nor UO_717 (O_717,N_14816,N_14935);
nand UO_718 (O_718,N_14993,N_14794);
and UO_719 (O_719,N_14872,N_14806);
nand UO_720 (O_720,N_14796,N_14794);
or UO_721 (O_721,N_14827,N_14962);
and UO_722 (O_722,N_14966,N_14933);
nand UO_723 (O_723,N_14885,N_14893);
or UO_724 (O_724,N_14814,N_14819);
nand UO_725 (O_725,N_14913,N_14766);
nor UO_726 (O_726,N_14887,N_14795);
nand UO_727 (O_727,N_14880,N_14829);
nor UO_728 (O_728,N_14834,N_14753);
and UO_729 (O_729,N_14934,N_14861);
and UO_730 (O_730,N_14770,N_14973);
and UO_731 (O_731,N_14800,N_14898);
or UO_732 (O_732,N_14910,N_14801);
or UO_733 (O_733,N_14765,N_14975);
and UO_734 (O_734,N_14972,N_14845);
nor UO_735 (O_735,N_14836,N_14815);
xor UO_736 (O_736,N_14834,N_14979);
nor UO_737 (O_737,N_14822,N_14891);
or UO_738 (O_738,N_14788,N_14786);
or UO_739 (O_739,N_14958,N_14808);
and UO_740 (O_740,N_14752,N_14845);
or UO_741 (O_741,N_14918,N_14851);
or UO_742 (O_742,N_14969,N_14773);
nor UO_743 (O_743,N_14873,N_14770);
and UO_744 (O_744,N_14939,N_14919);
or UO_745 (O_745,N_14912,N_14831);
and UO_746 (O_746,N_14900,N_14764);
or UO_747 (O_747,N_14962,N_14790);
xnor UO_748 (O_748,N_14805,N_14779);
and UO_749 (O_749,N_14824,N_14777);
nor UO_750 (O_750,N_14869,N_14824);
nor UO_751 (O_751,N_14830,N_14763);
nor UO_752 (O_752,N_14801,N_14759);
xor UO_753 (O_753,N_14832,N_14852);
nand UO_754 (O_754,N_14771,N_14793);
nand UO_755 (O_755,N_14757,N_14996);
nor UO_756 (O_756,N_14797,N_14822);
or UO_757 (O_757,N_14754,N_14853);
or UO_758 (O_758,N_14967,N_14755);
or UO_759 (O_759,N_14865,N_14971);
or UO_760 (O_760,N_14857,N_14780);
and UO_761 (O_761,N_14789,N_14915);
xor UO_762 (O_762,N_14948,N_14876);
nor UO_763 (O_763,N_14944,N_14915);
nor UO_764 (O_764,N_14760,N_14766);
or UO_765 (O_765,N_14958,N_14902);
or UO_766 (O_766,N_14819,N_14912);
nand UO_767 (O_767,N_14929,N_14947);
nand UO_768 (O_768,N_14937,N_14909);
nor UO_769 (O_769,N_14960,N_14937);
nand UO_770 (O_770,N_14774,N_14940);
or UO_771 (O_771,N_14798,N_14804);
nor UO_772 (O_772,N_14760,N_14780);
nor UO_773 (O_773,N_14865,N_14832);
nor UO_774 (O_774,N_14754,N_14772);
and UO_775 (O_775,N_14767,N_14810);
nand UO_776 (O_776,N_14855,N_14857);
and UO_777 (O_777,N_14887,N_14830);
or UO_778 (O_778,N_14852,N_14781);
and UO_779 (O_779,N_14782,N_14889);
nand UO_780 (O_780,N_14822,N_14898);
or UO_781 (O_781,N_14769,N_14816);
xnor UO_782 (O_782,N_14945,N_14848);
or UO_783 (O_783,N_14996,N_14830);
and UO_784 (O_784,N_14795,N_14996);
or UO_785 (O_785,N_14956,N_14776);
nand UO_786 (O_786,N_14909,N_14941);
nand UO_787 (O_787,N_14881,N_14903);
or UO_788 (O_788,N_14790,N_14792);
and UO_789 (O_789,N_14782,N_14886);
nor UO_790 (O_790,N_14835,N_14793);
nor UO_791 (O_791,N_14788,N_14895);
nand UO_792 (O_792,N_14993,N_14864);
xor UO_793 (O_793,N_14959,N_14932);
or UO_794 (O_794,N_14756,N_14888);
or UO_795 (O_795,N_14883,N_14995);
or UO_796 (O_796,N_14999,N_14811);
or UO_797 (O_797,N_14788,N_14912);
and UO_798 (O_798,N_14984,N_14830);
nor UO_799 (O_799,N_14901,N_14917);
and UO_800 (O_800,N_14883,N_14882);
nor UO_801 (O_801,N_14853,N_14846);
and UO_802 (O_802,N_14918,N_14986);
nand UO_803 (O_803,N_14800,N_14995);
nor UO_804 (O_804,N_14970,N_14801);
and UO_805 (O_805,N_14978,N_14802);
and UO_806 (O_806,N_14878,N_14876);
xnor UO_807 (O_807,N_14972,N_14847);
nand UO_808 (O_808,N_14799,N_14775);
or UO_809 (O_809,N_14815,N_14832);
and UO_810 (O_810,N_14916,N_14816);
or UO_811 (O_811,N_14759,N_14755);
and UO_812 (O_812,N_14950,N_14988);
and UO_813 (O_813,N_14822,N_14924);
and UO_814 (O_814,N_14960,N_14951);
or UO_815 (O_815,N_14819,N_14786);
nand UO_816 (O_816,N_14911,N_14783);
or UO_817 (O_817,N_14775,N_14924);
xnor UO_818 (O_818,N_14766,N_14952);
xnor UO_819 (O_819,N_14934,N_14847);
nand UO_820 (O_820,N_14817,N_14986);
nor UO_821 (O_821,N_14757,N_14929);
nand UO_822 (O_822,N_14895,N_14819);
nor UO_823 (O_823,N_14892,N_14822);
nor UO_824 (O_824,N_14761,N_14984);
or UO_825 (O_825,N_14856,N_14842);
xnor UO_826 (O_826,N_14939,N_14847);
nor UO_827 (O_827,N_14865,N_14774);
xnor UO_828 (O_828,N_14980,N_14788);
or UO_829 (O_829,N_14827,N_14955);
or UO_830 (O_830,N_14852,N_14967);
and UO_831 (O_831,N_14851,N_14961);
nor UO_832 (O_832,N_14750,N_14856);
nand UO_833 (O_833,N_14827,N_14782);
nor UO_834 (O_834,N_14890,N_14878);
nor UO_835 (O_835,N_14841,N_14813);
or UO_836 (O_836,N_14808,N_14864);
or UO_837 (O_837,N_14810,N_14896);
nand UO_838 (O_838,N_14871,N_14832);
xnor UO_839 (O_839,N_14940,N_14929);
and UO_840 (O_840,N_14823,N_14979);
or UO_841 (O_841,N_14928,N_14936);
and UO_842 (O_842,N_14792,N_14919);
or UO_843 (O_843,N_14947,N_14982);
xor UO_844 (O_844,N_14841,N_14945);
and UO_845 (O_845,N_14926,N_14873);
nand UO_846 (O_846,N_14860,N_14830);
and UO_847 (O_847,N_14774,N_14871);
and UO_848 (O_848,N_14804,N_14771);
nor UO_849 (O_849,N_14898,N_14949);
and UO_850 (O_850,N_14960,N_14881);
xnor UO_851 (O_851,N_14893,N_14753);
nor UO_852 (O_852,N_14960,N_14861);
nand UO_853 (O_853,N_14993,N_14778);
and UO_854 (O_854,N_14817,N_14875);
and UO_855 (O_855,N_14899,N_14915);
nor UO_856 (O_856,N_14799,N_14808);
nor UO_857 (O_857,N_14913,N_14945);
xnor UO_858 (O_858,N_14991,N_14843);
nor UO_859 (O_859,N_14868,N_14974);
nor UO_860 (O_860,N_14771,N_14951);
xor UO_861 (O_861,N_14901,N_14808);
nor UO_862 (O_862,N_14929,N_14848);
nor UO_863 (O_863,N_14994,N_14829);
and UO_864 (O_864,N_14917,N_14863);
or UO_865 (O_865,N_14957,N_14781);
nand UO_866 (O_866,N_14966,N_14799);
nor UO_867 (O_867,N_14944,N_14921);
nor UO_868 (O_868,N_14786,N_14995);
xor UO_869 (O_869,N_14839,N_14975);
nor UO_870 (O_870,N_14868,N_14988);
nand UO_871 (O_871,N_14788,N_14929);
nand UO_872 (O_872,N_14784,N_14758);
or UO_873 (O_873,N_14963,N_14877);
and UO_874 (O_874,N_14825,N_14830);
and UO_875 (O_875,N_14937,N_14832);
nand UO_876 (O_876,N_14755,N_14921);
nor UO_877 (O_877,N_14880,N_14939);
nand UO_878 (O_878,N_14976,N_14890);
nor UO_879 (O_879,N_14977,N_14812);
nand UO_880 (O_880,N_14812,N_14982);
nor UO_881 (O_881,N_14751,N_14886);
and UO_882 (O_882,N_14922,N_14968);
and UO_883 (O_883,N_14835,N_14940);
nor UO_884 (O_884,N_14872,N_14978);
or UO_885 (O_885,N_14848,N_14864);
nand UO_886 (O_886,N_14854,N_14760);
nand UO_887 (O_887,N_14787,N_14983);
nand UO_888 (O_888,N_14836,N_14805);
and UO_889 (O_889,N_14938,N_14986);
or UO_890 (O_890,N_14929,N_14780);
nor UO_891 (O_891,N_14758,N_14863);
nand UO_892 (O_892,N_14951,N_14765);
nor UO_893 (O_893,N_14892,N_14769);
or UO_894 (O_894,N_14854,N_14980);
nand UO_895 (O_895,N_14921,N_14940);
xor UO_896 (O_896,N_14761,N_14902);
xnor UO_897 (O_897,N_14870,N_14873);
or UO_898 (O_898,N_14884,N_14872);
or UO_899 (O_899,N_14877,N_14861);
nand UO_900 (O_900,N_14985,N_14937);
and UO_901 (O_901,N_14848,N_14832);
nor UO_902 (O_902,N_14860,N_14910);
nand UO_903 (O_903,N_14837,N_14993);
nand UO_904 (O_904,N_14918,N_14841);
and UO_905 (O_905,N_14920,N_14795);
nor UO_906 (O_906,N_14910,N_14817);
and UO_907 (O_907,N_14907,N_14909);
and UO_908 (O_908,N_14987,N_14849);
and UO_909 (O_909,N_14760,N_14869);
and UO_910 (O_910,N_14785,N_14902);
nor UO_911 (O_911,N_14896,N_14864);
xor UO_912 (O_912,N_14951,N_14831);
or UO_913 (O_913,N_14771,N_14967);
nand UO_914 (O_914,N_14926,N_14846);
nor UO_915 (O_915,N_14932,N_14900);
and UO_916 (O_916,N_14944,N_14792);
nand UO_917 (O_917,N_14856,N_14993);
or UO_918 (O_918,N_14994,N_14831);
and UO_919 (O_919,N_14764,N_14912);
and UO_920 (O_920,N_14959,N_14795);
or UO_921 (O_921,N_14807,N_14915);
and UO_922 (O_922,N_14971,N_14816);
nand UO_923 (O_923,N_14998,N_14878);
and UO_924 (O_924,N_14756,N_14862);
nor UO_925 (O_925,N_14957,N_14947);
nor UO_926 (O_926,N_14806,N_14958);
xor UO_927 (O_927,N_14945,N_14921);
or UO_928 (O_928,N_14937,N_14788);
xnor UO_929 (O_929,N_14759,N_14821);
or UO_930 (O_930,N_14971,N_14861);
nand UO_931 (O_931,N_14959,N_14940);
or UO_932 (O_932,N_14798,N_14805);
or UO_933 (O_933,N_14864,N_14817);
nand UO_934 (O_934,N_14934,N_14778);
nor UO_935 (O_935,N_14988,N_14987);
or UO_936 (O_936,N_14952,N_14931);
or UO_937 (O_937,N_14868,N_14783);
nor UO_938 (O_938,N_14869,N_14817);
and UO_939 (O_939,N_14930,N_14848);
nor UO_940 (O_940,N_14809,N_14977);
or UO_941 (O_941,N_14755,N_14792);
or UO_942 (O_942,N_14941,N_14927);
or UO_943 (O_943,N_14805,N_14769);
nand UO_944 (O_944,N_14763,N_14980);
or UO_945 (O_945,N_14756,N_14973);
and UO_946 (O_946,N_14825,N_14804);
nand UO_947 (O_947,N_14838,N_14986);
xnor UO_948 (O_948,N_14965,N_14885);
nor UO_949 (O_949,N_14921,N_14777);
nand UO_950 (O_950,N_14848,N_14905);
nand UO_951 (O_951,N_14999,N_14815);
nor UO_952 (O_952,N_14928,N_14995);
nor UO_953 (O_953,N_14976,N_14986);
or UO_954 (O_954,N_14929,N_14751);
nor UO_955 (O_955,N_14921,N_14922);
xor UO_956 (O_956,N_14955,N_14783);
nor UO_957 (O_957,N_14867,N_14837);
and UO_958 (O_958,N_14843,N_14992);
and UO_959 (O_959,N_14755,N_14886);
nand UO_960 (O_960,N_14814,N_14965);
nand UO_961 (O_961,N_14758,N_14830);
or UO_962 (O_962,N_14978,N_14887);
and UO_963 (O_963,N_14939,N_14802);
nor UO_964 (O_964,N_14951,N_14807);
or UO_965 (O_965,N_14769,N_14857);
nor UO_966 (O_966,N_14755,N_14987);
or UO_967 (O_967,N_14926,N_14984);
nor UO_968 (O_968,N_14854,N_14757);
or UO_969 (O_969,N_14992,N_14959);
or UO_970 (O_970,N_14953,N_14805);
xor UO_971 (O_971,N_14866,N_14990);
nor UO_972 (O_972,N_14967,N_14863);
or UO_973 (O_973,N_14923,N_14830);
xor UO_974 (O_974,N_14953,N_14944);
and UO_975 (O_975,N_14891,N_14888);
nor UO_976 (O_976,N_14871,N_14952);
and UO_977 (O_977,N_14772,N_14840);
and UO_978 (O_978,N_14946,N_14826);
and UO_979 (O_979,N_14810,N_14762);
nor UO_980 (O_980,N_14983,N_14833);
or UO_981 (O_981,N_14899,N_14778);
nor UO_982 (O_982,N_14976,N_14903);
or UO_983 (O_983,N_14802,N_14988);
xnor UO_984 (O_984,N_14779,N_14972);
nand UO_985 (O_985,N_14795,N_14787);
or UO_986 (O_986,N_14789,N_14805);
nand UO_987 (O_987,N_14830,N_14869);
nand UO_988 (O_988,N_14990,N_14887);
and UO_989 (O_989,N_14812,N_14777);
nand UO_990 (O_990,N_14971,N_14902);
and UO_991 (O_991,N_14949,N_14858);
nand UO_992 (O_992,N_14985,N_14917);
nand UO_993 (O_993,N_14873,N_14937);
and UO_994 (O_994,N_14859,N_14830);
nor UO_995 (O_995,N_14836,N_14753);
or UO_996 (O_996,N_14875,N_14967);
or UO_997 (O_997,N_14822,N_14802);
and UO_998 (O_998,N_14866,N_14907);
or UO_999 (O_999,N_14787,N_14956);
nand UO_1000 (O_1000,N_14753,N_14917);
xor UO_1001 (O_1001,N_14806,N_14860);
and UO_1002 (O_1002,N_14782,N_14818);
or UO_1003 (O_1003,N_14959,N_14972);
xnor UO_1004 (O_1004,N_14796,N_14876);
and UO_1005 (O_1005,N_14855,N_14901);
and UO_1006 (O_1006,N_14796,N_14903);
nand UO_1007 (O_1007,N_14909,N_14969);
nor UO_1008 (O_1008,N_14911,N_14792);
xor UO_1009 (O_1009,N_14868,N_14814);
nand UO_1010 (O_1010,N_14797,N_14936);
or UO_1011 (O_1011,N_14819,N_14835);
or UO_1012 (O_1012,N_14929,N_14785);
nor UO_1013 (O_1013,N_14780,N_14773);
and UO_1014 (O_1014,N_14779,N_14788);
or UO_1015 (O_1015,N_14865,N_14998);
xor UO_1016 (O_1016,N_14957,N_14834);
or UO_1017 (O_1017,N_14847,N_14997);
or UO_1018 (O_1018,N_14764,N_14819);
nor UO_1019 (O_1019,N_14787,N_14850);
xor UO_1020 (O_1020,N_14975,N_14852);
or UO_1021 (O_1021,N_14887,N_14994);
nor UO_1022 (O_1022,N_14903,N_14995);
and UO_1023 (O_1023,N_14999,N_14843);
nand UO_1024 (O_1024,N_14752,N_14814);
nor UO_1025 (O_1025,N_14870,N_14835);
or UO_1026 (O_1026,N_14824,N_14950);
xor UO_1027 (O_1027,N_14804,N_14762);
nand UO_1028 (O_1028,N_14863,N_14999);
and UO_1029 (O_1029,N_14903,N_14779);
nand UO_1030 (O_1030,N_14792,N_14781);
or UO_1031 (O_1031,N_14924,N_14836);
or UO_1032 (O_1032,N_14975,N_14788);
or UO_1033 (O_1033,N_14794,N_14984);
and UO_1034 (O_1034,N_14935,N_14909);
and UO_1035 (O_1035,N_14929,N_14814);
or UO_1036 (O_1036,N_14853,N_14751);
nand UO_1037 (O_1037,N_14813,N_14862);
or UO_1038 (O_1038,N_14821,N_14964);
nand UO_1039 (O_1039,N_14823,N_14876);
nand UO_1040 (O_1040,N_14771,N_14915);
and UO_1041 (O_1041,N_14893,N_14923);
nand UO_1042 (O_1042,N_14972,N_14987);
nor UO_1043 (O_1043,N_14994,N_14979);
nand UO_1044 (O_1044,N_14980,N_14953);
nand UO_1045 (O_1045,N_14752,N_14753);
nor UO_1046 (O_1046,N_14900,N_14899);
or UO_1047 (O_1047,N_14960,N_14888);
or UO_1048 (O_1048,N_14988,N_14844);
or UO_1049 (O_1049,N_14943,N_14819);
nor UO_1050 (O_1050,N_14878,N_14853);
xnor UO_1051 (O_1051,N_14953,N_14955);
and UO_1052 (O_1052,N_14775,N_14791);
nand UO_1053 (O_1053,N_14799,N_14809);
or UO_1054 (O_1054,N_14900,N_14978);
xor UO_1055 (O_1055,N_14860,N_14841);
nand UO_1056 (O_1056,N_14922,N_14995);
nor UO_1057 (O_1057,N_14818,N_14864);
and UO_1058 (O_1058,N_14889,N_14921);
nand UO_1059 (O_1059,N_14812,N_14963);
or UO_1060 (O_1060,N_14797,N_14964);
or UO_1061 (O_1061,N_14983,N_14820);
or UO_1062 (O_1062,N_14802,N_14779);
and UO_1063 (O_1063,N_14891,N_14998);
and UO_1064 (O_1064,N_14825,N_14954);
nor UO_1065 (O_1065,N_14968,N_14840);
nand UO_1066 (O_1066,N_14855,N_14774);
nand UO_1067 (O_1067,N_14904,N_14991);
or UO_1068 (O_1068,N_14975,N_14796);
or UO_1069 (O_1069,N_14765,N_14829);
and UO_1070 (O_1070,N_14823,N_14974);
nand UO_1071 (O_1071,N_14763,N_14917);
or UO_1072 (O_1072,N_14855,N_14932);
or UO_1073 (O_1073,N_14851,N_14936);
nand UO_1074 (O_1074,N_14985,N_14942);
nand UO_1075 (O_1075,N_14786,N_14911);
and UO_1076 (O_1076,N_14950,N_14808);
xor UO_1077 (O_1077,N_14828,N_14918);
and UO_1078 (O_1078,N_14814,N_14788);
nand UO_1079 (O_1079,N_14895,N_14912);
xnor UO_1080 (O_1080,N_14900,N_14909);
and UO_1081 (O_1081,N_14764,N_14981);
and UO_1082 (O_1082,N_14835,N_14989);
nand UO_1083 (O_1083,N_14819,N_14797);
and UO_1084 (O_1084,N_14852,N_14844);
or UO_1085 (O_1085,N_14766,N_14924);
nor UO_1086 (O_1086,N_14798,N_14852);
nor UO_1087 (O_1087,N_14772,N_14848);
and UO_1088 (O_1088,N_14966,N_14865);
or UO_1089 (O_1089,N_14795,N_14968);
nor UO_1090 (O_1090,N_14932,N_14885);
or UO_1091 (O_1091,N_14753,N_14930);
nand UO_1092 (O_1092,N_14850,N_14821);
or UO_1093 (O_1093,N_14905,N_14998);
nor UO_1094 (O_1094,N_14913,N_14861);
or UO_1095 (O_1095,N_14809,N_14992);
nor UO_1096 (O_1096,N_14817,N_14975);
nand UO_1097 (O_1097,N_14996,N_14925);
and UO_1098 (O_1098,N_14929,N_14988);
nor UO_1099 (O_1099,N_14882,N_14755);
xor UO_1100 (O_1100,N_14813,N_14957);
nor UO_1101 (O_1101,N_14983,N_14829);
xnor UO_1102 (O_1102,N_14918,N_14944);
nand UO_1103 (O_1103,N_14991,N_14820);
xnor UO_1104 (O_1104,N_14894,N_14777);
xnor UO_1105 (O_1105,N_14765,N_14889);
or UO_1106 (O_1106,N_14841,N_14849);
or UO_1107 (O_1107,N_14908,N_14849);
and UO_1108 (O_1108,N_14817,N_14916);
nand UO_1109 (O_1109,N_14872,N_14800);
or UO_1110 (O_1110,N_14759,N_14905);
nand UO_1111 (O_1111,N_14774,N_14929);
nand UO_1112 (O_1112,N_14860,N_14939);
nand UO_1113 (O_1113,N_14758,N_14927);
and UO_1114 (O_1114,N_14859,N_14916);
nand UO_1115 (O_1115,N_14914,N_14801);
xor UO_1116 (O_1116,N_14911,N_14921);
nand UO_1117 (O_1117,N_14954,N_14866);
and UO_1118 (O_1118,N_14805,N_14841);
nor UO_1119 (O_1119,N_14978,N_14811);
nor UO_1120 (O_1120,N_14978,N_14936);
or UO_1121 (O_1121,N_14799,N_14981);
or UO_1122 (O_1122,N_14791,N_14863);
and UO_1123 (O_1123,N_14933,N_14757);
xnor UO_1124 (O_1124,N_14982,N_14956);
nand UO_1125 (O_1125,N_14799,N_14803);
nor UO_1126 (O_1126,N_14774,N_14881);
nor UO_1127 (O_1127,N_14988,N_14787);
nand UO_1128 (O_1128,N_14755,N_14876);
nand UO_1129 (O_1129,N_14790,N_14773);
nand UO_1130 (O_1130,N_14878,N_14893);
nand UO_1131 (O_1131,N_14921,N_14891);
nand UO_1132 (O_1132,N_14836,N_14750);
or UO_1133 (O_1133,N_14942,N_14769);
and UO_1134 (O_1134,N_14888,N_14780);
or UO_1135 (O_1135,N_14813,N_14887);
or UO_1136 (O_1136,N_14933,N_14818);
xor UO_1137 (O_1137,N_14870,N_14934);
nor UO_1138 (O_1138,N_14832,N_14982);
nor UO_1139 (O_1139,N_14860,N_14896);
nor UO_1140 (O_1140,N_14832,N_14949);
or UO_1141 (O_1141,N_14831,N_14802);
nand UO_1142 (O_1142,N_14913,N_14846);
or UO_1143 (O_1143,N_14808,N_14810);
nand UO_1144 (O_1144,N_14924,N_14921);
nor UO_1145 (O_1145,N_14791,N_14806);
xnor UO_1146 (O_1146,N_14813,N_14837);
nand UO_1147 (O_1147,N_14811,N_14800);
xnor UO_1148 (O_1148,N_14894,N_14807);
nand UO_1149 (O_1149,N_14817,N_14833);
and UO_1150 (O_1150,N_14775,N_14935);
or UO_1151 (O_1151,N_14836,N_14848);
nor UO_1152 (O_1152,N_14897,N_14904);
xnor UO_1153 (O_1153,N_14997,N_14755);
nor UO_1154 (O_1154,N_14816,N_14806);
nand UO_1155 (O_1155,N_14903,N_14755);
and UO_1156 (O_1156,N_14944,N_14855);
and UO_1157 (O_1157,N_14890,N_14974);
nor UO_1158 (O_1158,N_14966,N_14763);
or UO_1159 (O_1159,N_14788,N_14860);
and UO_1160 (O_1160,N_14916,N_14882);
or UO_1161 (O_1161,N_14877,N_14805);
or UO_1162 (O_1162,N_14866,N_14931);
nand UO_1163 (O_1163,N_14858,N_14859);
or UO_1164 (O_1164,N_14830,N_14946);
nor UO_1165 (O_1165,N_14868,N_14873);
and UO_1166 (O_1166,N_14902,N_14966);
and UO_1167 (O_1167,N_14970,N_14882);
nand UO_1168 (O_1168,N_14780,N_14806);
and UO_1169 (O_1169,N_14874,N_14830);
or UO_1170 (O_1170,N_14992,N_14990);
nor UO_1171 (O_1171,N_14821,N_14820);
and UO_1172 (O_1172,N_14870,N_14933);
nand UO_1173 (O_1173,N_14991,N_14883);
nand UO_1174 (O_1174,N_14800,N_14982);
nand UO_1175 (O_1175,N_14927,N_14945);
nand UO_1176 (O_1176,N_14993,N_14803);
and UO_1177 (O_1177,N_14755,N_14862);
and UO_1178 (O_1178,N_14966,N_14894);
or UO_1179 (O_1179,N_14779,N_14873);
nand UO_1180 (O_1180,N_14809,N_14880);
nor UO_1181 (O_1181,N_14964,N_14915);
nor UO_1182 (O_1182,N_14834,N_14820);
nand UO_1183 (O_1183,N_14843,N_14927);
or UO_1184 (O_1184,N_14897,N_14954);
or UO_1185 (O_1185,N_14776,N_14972);
or UO_1186 (O_1186,N_14912,N_14962);
nand UO_1187 (O_1187,N_14869,N_14995);
nor UO_1188 (O_1188,N_14962,N_14956);
nor UO_1189 (O_1189,N_14961,N_14974);
nor UO_1190 (O_1190,N_14896,N_14790);
or UO_1191 (O_1191,N_14977,N_14999);
nor UO_1192 (O_1192,N_14832,N_14768);
nor UO_1193 (O_1193,N_14886,N_14869);
nand UO_1194 (O_1194,N_14821,N_14915);
nand UO_1195 (O_1195,N_14797,N_14780);
and UO_1196 (O_1196,N_14835,N_14886);
nor UO_1197 (O_1197,N_14942,N_14814);
or UO_1198 (O_1198,N_14964,N_14777);
or UO_1199 (O_1199,N_14922,N_14908);
nand UO_1200 (O_1200,N_14922,N_14755);
and UO_1201 (O_1201,N_14893,N_14883);
or UO_1202 (O_1202,N_14910,N_14991);
nor UO_1203 (O_1203,N_14767,N_14837);
xor UO_1204 (O_1204,N_14991,N_14824);
nor UO_1205 (O_1205,N_14947,N_14844);
nand UO_1206 (O_1206,N_14870,N_14753);
or UO_1207 (O_1207,N_14769,N_14976);
nor UO_1208 (O_1208,N_14812,N_14921);
or UO_1209 (O_1209,N_14946,N_14754);
or UO_1210 (O_1210,N_14928,N_14888);
nor UO_1211 (O_1211,N_14903,N_14838);
and UO_1212 (O_1212,N_14942,N_14875);
and UO_1213 (O_1213,N_14957,N_14827);
nand UO_1214 (O_1214,N_14851,N_14907);
and UO_1215 (O_1215,N_14794,N_14771);
nor UO_1216 (O_1216,N_14856,N_14762);
or UO_1217 (O_1217,N_14904,N_14909);
or UO_1218 (O_1218,N_14760,N_14981);
and UO_1219 (O_1219,N_14792,N_14800);
xor UO_1220 (O_1220,N_14805,N_14903);
and UO_1221 (O_1221,N_14843,N_14920);
nand UO_1222 (O_1222,N_14993,N_14791);
and UO_1223 (O_1223,N_14923,N_14917);
nor UO_1224 (O_1224,N_14887,N_14967);
and UO_1225 (O_1225,N_14937,N_14973);
and UO_1226 (O_1226,N_14882,N_14931);
nor UO_1227 (O_1227,N_14783,N_14757);
xor UO_1228 (O_1228,N_14818,N_14830);
nor UO_1229 (O_1229,N_14845,N_14878);
and UO_1230 (O_1230,N_14784,N_14905);
nor UO_1231 (O_1231,N_14884,N_14815);
or UO_1232 (O_1232,N_14894,N_14767);
and UO_1233 (O_1233,N_14821,N_14857);
xor UO_1234 (O_1234,N_14842,N_14778);
nor UO_1235 (O_1235,N_14880,N_14899);
nand UO_1236 (O_1236,N_14792,N_14834);
nor UO_1237 (O_1237,N_14763,N_14965);
and UO_1238 (O_1238,N_14800,N_14750);
and UO_1239 (O_1239,N_14833,N_14802);
or UO_1240 (O_1240,N_14845,N_14953);
nand UO_1241 (O_1241,N_14994,N_14827);
nand UO_1242 (O_1242,N_14766,N_14851);
nor UO_1243 (O_1243,N_14916,N_14870);
and UO_1244 (O_1244,N_14989,N_14776);
or UO_1245 (O_1245,N_14903,N_14883);
nand UO_1246 (O_1246,N_14926,N_14839);
or UO_1247 (O_1247,N_14966,N_14825);
or UO_1248 (O_1248,N_14818,N_14844);
nor UO_1249 (O_1249,N_14853,N_14841);
nor UO_1250 (O_1250,N_14825,N_14837);
nor UO_1251 (O_1251,N_14957,N_14935);
or UO_1252 (O_1252,N_14957,N_14954);
and UO_1253 (O_1253,N_14782,N_14831);
and UO_1254 (O_1254,N_14969,N_14752);
and UO_1255 (O_1255,N_14757,N_14778);
or UO_1256 (O_1256,N_14952,N_14851);
or UO_1257 (O_1257,N_14959,N_14973);
nand UO_1258 (O_1258,N_14955,N_14789);
and UO_1259 (O_1259,N_14876,N_14867);
and UO_1260 (O_1260,N_14816,N_14979);
and UO_1261 (O_1261,N_14946,N_14828);
nor UO_1262 (O_1262,N_14995,N_14851);
nand UO_1263 (O_1263,N_14850,N_14801);
and UO_1264 (O_1264,N_14979,N_14891);
nor UO_1265 (O_1265,N_14937,N_14824);
nor UO_1266 (O_1266,N_14852,N_14977);
nand UO_1267 (O_1267,N_14759,N_14828);
and UO_1268 (O_1268,N_14894,N_14828);
nor UO_1269 (O_1269,N_14792,N_14913);
and UO_1270 (O_1270,N_14819,N_14862);
nand UO_1271 (O_1271,N_14869,N_14982);
xor UO_1272 (O_1272,N_14960,N_14837);
nand UO_1273 (O_1273,N_14885,N_14845);
nor UO_1274 (O_1274,N_14960,N_14889);
nand UO_1275 (O_1275,N_14830,N_14752);
or UO_1276 (O_1276,N_14979,N_14980);
and UO_1277 (O_1277,N_14816,N_14819);
xor UO_1278 (O_1278,N_14881,N_14828);
nand UO_1279 (O_1279,N_14757,N_14874);
nand UO_1280 (O_1280,N_14879,N_14794);
and UO_1281 (O_1281,N_14823,N_14793);
or UO_1282 (O_1282,N_14924,N_14984);
xnor UO_1283 (O_1283,N_14813,N_14771);
and UO_1284 (O_1284,N_14942,N_14812);
or UO_1285 (O_1285,N_14932,N_14970);
and UO_1286 (O_1286,N_14778,N_14983);
or UO_1287 (O_1287,N_14876,N_14956);
nor UO_1288 (O_1288,N_14782,N_14869);
and UO_1289 (O_1289,N_14787,N_14828);
and UO_1290 (O_1290,N_14883,N_14821);
xnor UO_1291 (O_1291,N_14908,N_14972);
nor UO_1292 (O_1292,N_14952,N_14963);
nor UO_1293 (O_1293,N_14865,N_14920);
nor UO_1294 (O_1294,N_14773,N_14979);
xor UO_1295 (O_1295,N_14766,N_14812);
nor UO_1296 (O_1296,N_14899,N_14895);
nor UO_1297 (O_1297,N_14965,N_14924);
nand UO_1298 (O_1298,N_14924,N_14865);
nand UO_1299 (O_1299,N_14960,N_14794);
nor UO_1300 (O_1300,N_14835,N_14972);
or UO_1301 (O_1301,N_14843,N_14831);
nand UO_1302 (O_1302,N_14888,N_14779);
nand UO_1303 (O_1303,N_14789,N_14853);
nand UO_1304 (O_1304,N_14822,N_14918);
xnor UO_1305 (O_1305,N_14999,N_14900);
nand UO_1306 (O_1306,N_14795,N_14803);
xor UO_1307 (O_1307,N_14875,N_14831);
nor UO_1308 (O_1308,N_14833,N_14831);
nand UO_1309 (O_1309,N_14809,N_14751);
nand UO_1310 (O_1310,N_14847,N_14836);
nand UO_1311 (O_1311,N_14890,N_14792);
xnor UO_1312 (O_1312,N_14929,N_14938);
and UO_1313 (O_1313,N_14901,N_14994);
or UO_1314 (O_1314,N_14873,N_14925);
and UO_1315 (O_1315,N_14849,N_14957);
xnor UO_1316 (O_1316,N_14916,N_14993);
and UO_1317 (O_1317,N_14926,N_14845);
or UO_1318 (O_1318,N_14809,N_14778);
or UO_1319 (O_1319,N_14837,N_14979);
nand UO_1320 (O_1320,N_14889,N_14985);
nor UO_1321 (O_1321,N_14956,N_14831);
or UO_1322 (O_1322,N_14996,N_14759);
xnor UO_1323 (O_1323,N_14922,N_14873);
nor UO_1324 (O_1324,N_14791,N_14854);
nand UO_1325 (O_1325,N_14867,N_14859);
and UO_1326 (O_1326,N_14808,N_14929);
nor UO_1327 (O_1327,N_14776,N_14856);
or UO_1328 (O_1328,N_14776,N_14878);
or UO_1329 (O_1329,N_14849,N_14861);
nand UO_1330 (O_1330,N_14841,N_14831);
and UO_1331 (O_1331,N_14808,N_14814);
or UO_1332 (O_1332,N_14942,N_14766);
nand UO_1333 (O_1333,N_14933,N_14957);
nor UO_1334 (O_1334,N_14916,N_14774);
nor UO_1335 (O_1335,N_14959,N_14965);
or UO_1336 (O_1336,N_14985,N_14919);
xor UO_1337 (O_1337,N_14887,N_14989);
nor UO_1338 (O_1338,N_14854,N_14964);
or UO_1339 (O_1339,N_14935,N_14896);
and UO_1340 (O_1340,N_14813,N_14800);
or UO_1341 (O_1341,N_14784,N_14755);
or UO_1342 (O_1342,N_14894,N_14847);
nor UO_1343 (O_1343,N_14795,N_14994);
nor UO_1344 (O_1344,N_14777,N_14853);
nand UO_1345 (O_1345,N_14797,N_14860);
or UO_1346 (O_1346,N_14904,N_14848);
nor UO_1347 (O_1347,N_14991,N_14982);
nand UO_1348 (O_1348,N_14829,N_14875);
and UO_1349 (O_1349,N_14904,N_14942);
nor UO_1350 (O_1350,N_14839,N_14767);
nand UO_1351 (O_1351,N_14951,N_14904);
and UO_1352 (O_1352,N_14765,N_14864);
xor UO_1353 (O_1353,N_14896,N_14771);
nor UO_1354 (O_1354,N_14976,N_14863);
nand UO_1355 (O_1355,N_14982,N_14883);
nor UO_1356 (O_1356,N_14840,N_14919);
xnor UO_1357 (O_1357,N_14847,N_14805);
and UO_1358 (O_1358,N_14802,N_14896);
or UO_1359 (O_1359,N_14913,N_14785);
or UO_1360 (O_1360,N_14937,N_14859);
nand UO_1361 (O_1361,N_14942,N_14791);
or UO_1362 (O_1362,N_14775,N_14957);
or UO_1363 (O_1363,N_14921,N_14759);
or UO_1364 (O_1364,N_14919,N_14902);
or UO_1365 (O_1365,N_14860,N_14855);
nand UO_1366 (O_1366,N_14843,N_14823);
or UO_1367 (O_1367,N_14917,N_14787);
and UO_1368 (O_1368,N_14921,N_14771);
nand UO_1369 (O_1369,N_14758,N_14862);
nand UO_1370 (O_1370,N_14776,N_14969);
and UO_1371 (O_1371,N_14911,N_14900);
xor UO_1372 (O_1372,N_14810,N_14803);
xnor UO_1373 (O_1373,N_14810,N_14924);
nand UO_1374 (O_1374,N_14907,N_14790);
nor UO_1375 (O_1375,N_14930,N_14927);
nand UO_1376 (O_1376,N_14893,N_14879);
and UO_1377 (O_1377,N_14999,N_14951);
and UO_1378 (O_1378,N_14929,N_14886);
and UO_1379 (O_1379,N_14761,N_14839);
nor UO_1380 (O_1380,N_14941,N_14972);
and UO_1381 (O_1381,N_14865,N_14826);
nand UO_1382 (O_1382,N_14799,N_14831);
or UO_1383 (O_1383,N_14943,N_14822);
nor UO_1384 (O_1384,N_14865,N_14981);
or UO_1385 (O_1385,N_14883,N_14948);
nor UO_1386 (O_1386,N_14846,N_14993);
and UO_1387 (O_1387,N_14891,N_14817);
or UO_1388 (O_1388,N_14870,N_14857);
nor UO_1389 (O_1389,N_14785,N_14930);
nor UO_1390 (O_1390,N_14756,N_14960);
or UO_1391 (O_1391,N_14959,N_14850);
nor UO_1392 (O_1392,N_14876,N_14789);
or UO_1393 (O_1393,N_14860,N_14804);
nor UO_1394 (O_1394,N_14890,N_14980);
or UO_1395 (O_1395,N_14920,N_14753);
nor UO_1396 (O_1396,N_14763,N_14986);
and UO_1397 (O_1397,N_14784,N_14918);
and UO_1398 (O_1398,N_14851,N_14754);
nand UO_1399 (O_1399,N_14964,N_14900);
nand UO_1400 (O_1400,N_14903,N_14860);
nor UO_1401 (O_1401,N_14827,N_14870);
and UO_1402 (O_1402,N_14753,N_14800);
nor UO_1403 (O_1403,N_14784,N_14966);
nor UO_1404 (O_1404,N_14774,N_14781);
nor UO_1405 (O_1405,N_14950,N_14891);
xnor UO_1406 (O_1406,N_14773,N_14985);
or UO_1407 (O_1407,N_14825,N_14772);
xor UO_1408 (O_1408,N_14763,N_14820);
nand UO_1409 (O_1409,N_14963,N_14957);
nor UO_1410 (O_1410,N_14899,N_14898);
or UO_1411 (O_1411,N_14928,N_14996);
nand UO_1412 (O_1412,N_14774,N_14899);
xor UO_1413 (O_1413,N_14982,N_14825);
nor UO_1414 (O_1414,N_14886,N_14807);
nand UO_1415 (O_1415,N_14857,N_14954);
or UO_1416 (O_1416,N_14804,N_14811);
or UO_1417 (O_1417,N_14922,N_14933);
xor UO_1418 (O_1418,N_14859,N_14888);
nand UO_1419 (O_1419,N_14761,N_14886);
and UO_1420 (O_1420,N_14887,N_14848);
xor UO_1421 (O_1421,N_14954,N_14935);
nor UO_1422 (O_1422,N_14980,N_14964);
and UO_1423 (O_1423,N_14993,N_14847);
nand UO_1424 (O_1424,N_14951,N_14918);
and UO_1425 (O_1425,N_14778,N_14941);
or UO_1426 (O_1426,N_14874,N_14878);
nor UO_1427 (O_1427,N_14995,N_14757);
nand UO_1428 (O_1428,N_14830,N_14826);
nor UO_1429 (O_1429,N_14982,N_14856);
or UO_1430 (O_1430,N_14769,N_14882);
or UO_1431 (O_1431,N_14894,N_14770);
and UO_1432 (O_1432,N_14890,N_14879);
and UO_1433 (O_1433,N_14893,N_14897);
and UO_1434 (O_1434,N_14916,N_14903);
and UO_1435 (O_1435,N_14870,N_14869);
xnor UO_1436 (O_1436,N_14830,N_14899);
or UO_1437 (O_1437,N_14901,N_14858);
nand UO_1438 (O_1438,N_14938,N_14960);
xnor UO_1439 (O_1439,N_14996,N_14821);
and UO_1440 (O_1440,N_14814,N_14980);
nor UO_1441 (O_1441,N_14765,N_14787);
nand UO_1442 (O_1442,N_14974,N_14842);
or UO_1443 (O_1443,N_14771,N_14957);
nand UO_1444 (O_1444,N_14790,N_14882);
xnor UO_1445 (O_1445,N_14784,N_14768);
or UO_1446 (O_1446,N_14792,N_14949);
nand UO_1447 (O_1447,N_14811,N_14768);
and UO_1448 (O_1448,N_14991,N_14969);
and UO_1449 (O_1449,N_14887,N_14793);
nor UO_1450 (O_1450,N_14987,N_14991);
and UO_1451 (O_1451,N_14873,N_14954);
nor UO_1452 (O_1452,N_14903,N_14877);
and UO_1453 (O_1453,N_14852,N_14795);
or UO_1454 (O_1454,N_14916,N_14944);
nor UO_1455 (O_1455,N_14937,N_14843);
and UO_1456 (O_1456,N_14916,N_14991);
or UO_1457 (O_1457,N_14766,N_14880);
nand UO_1458 (O_1458,N_14794,N_14760);
and UO_1459 (O_1459,N_14937,N_14839);
nor UO_1460 (O_1460,N_14765,N_14796);
xnor UO_1461 (O_1461,N_14902,N_14842);
nand UO_1462 (O_1462,N_14773,N_14791);
nand UO_1463 (O_1463,N_14919,N_14953);
and UO_1464 (O_1464,N_14984,N_14843);
nor UO_1465 (O_1465,N_14755,N_14981);
nand UO_1466 (O_1466,N_14854,N_14933);
and UO_1467 (O_1467,N_14992,N_14904);
nor UO_1468 (O_1468,N_14794,N_14873);
nor UO_1469 (O_1469,N_14785,N_14874);
and UO_1470 (O_1470,N_14879,N_14932);
and UO_1471 (O_1471,N_14750,N_14973);
nand UO_1472 (O_1472,N_14753,N_14982);
nor UO_1473 (O_1473,N_14814,N_14858);
or UO_1474 (O_1474,N_14874,N_14947);
and UO_1475 (O_1475,N_14909,N_14844);
xnor UO_1476 (O_1476,N_14944,N_14905);
nand UO_1477 (O_1477,N_14941,N_14953);
or UO_1478 (O_1478,N_14915,N_14942);
and UO_1479 (O_1479,N_14969,N_14855);
xor UO_1480 (O_1480,N_14892,N_14965);
nor UO_1481 (O_1481,N_14761,N_14762);
nor UO_1482 (O_1482,N_14803,N_14769);
or UO_1483 (O_1483,N_14816,N_14877);
nand UO_1484 (O_1484,N_14931,N_14770);
and UO_1485 (O_1485,N_14923,N_14815);
nand UO_1486 (O_1486,N_14766,N_14932);
nor UO_1487 (O_1487,N_14900,N_14804);
or UO_1488 (O_1488,N_14793,N_14830);
nand UO_1489 (O_1489,N_14820,N_14789);
or UO_1490 (O_1490,N_14858,N_14911);
and UO_1491 (O_1491,N_14849,N_14990);
nor UO_1492 (O_1492,N_14924,N_14818);
or UO_1493 (O_1493,N_14916,N_14864);
nand UO_1494 (O_1494,N_14803,N_14901);
nor UO_1495 (O_1495,N_14796,N_14926);
or UO_1496 (O_1496,N_14856,N_14980);
nand UO_1497 (O_1497,N_14945,N_14953);
xnor UO_1498 (O_1498,N_14953,N_14863);
and UO_1499 (O_1499,N_14973,N_14878);
nand UO_1500 (O_1500,N_14869,N_14944);
xor UO_1501 (O_1501,N_14808,N_14917);
xnor UO_1502 (O_1502,N_14789,N_14799);
or UO_1503 (O_1503,N_14826,N_14886);
or UO_1504 (O_1504,N_14782,N_14834);
or UO_1505 (O_1505,N_14870,N_14957);
nor UO_1506 (O_1506,N_14927,N_14990);
and UO_1507 (O_1507,N_14936,N_14929);
or UO_1508 (O_1508,N_14892,N_14841);
and UO_1509 (O_1509,N_14764,N_14843);
and UO_1510 (O_1510,N_14905,N_14887);
or UO_1511 (O_1511,N_14940,N_14854);
and UO_1512 (O_1512,N_14978,N_14796);
or UO_1513 (O_1513,N_14908,N_14831);
and UO_1514 (O_1514,N_14985,N_14766);
or UO_1515 (O_1515,N_14844,N_14846);
or UO_1516 (O_1516,N_14778,N_14981);
or UO_1517 (O_1517,N_14971,N_14993);
or UO_1518 (O_1518,N_14869,N_14948);
nand UO_1519 (O_1519,N_14994,N_14992);
or UO_1520 (O_1520,N_14751,N_14820);
nor UO_1521 (O_1521,N_14865,N_14915);
nand UO_1522 (O_1522,N_14950,N_14843);
nand UO_1523 (O_1523,N_14992,N_14929);
nand UO_1524 (O_1524,N_14974,N_14910);
nor UO_1525 (O_1525,N_14995,N_14889);
nor UO_1526 (O_1526,N_14858,N_14815);
and UO_1527 (O_1527,N_14989,N_14914);
nand UO_1528 (O_1528,N_14948,N_14901);
nand UO_1529 (O_1529,N_14779,N_14792);
nor UO_1530 (O_1530,N_14904,N_14948);
or UO_1531 (O_1531,N_14989,N_14944);
nand UO_1532 (O_1532,N_14797,N_14841);
nor UO_1533 (O_1533,N_14970,N_14884);
xor UO_1534 (O_1534,N_14796,N_14882);
and UO_1535 (O_1535,N_14785,N_14827);
or UO_1536 (O_1536,N_14964,N_14979);
and UO_1537 (O_1537,N_14818,N_14775);
and UO_1538 (O_1538,N_14865,N_14989);
and UO_1539 (O_1539,N_14838,N_14871);
and UO_1540 (O_1540,N_14981,N_14779);
nor UO_1541 (O_1541,N_14889,N_14931);
nor UO_1542 (O_1542,N_14756,N_14959);
nand UO_1543 (O_1543,N_14779,N_14889);
nor UO_1544 (O_1544,N_14923,N_14910);
nand UO_1545 (O_1545,N_14901,N_14929);
or UO_1546 (O_1546,N_14956,N_14977);
nand UO_1547 (O_1547,N_14814,N_14779);
nand UO_1548 (O_1548,N_14832,N_14780);
nand UO_1549 (O_1549,N_14893,N_14780);
nor UO_1550 (O_1550,N_14882,N_14995);
nor UO_1551 (O_1551,N_14966,N_14765);
nor UO_1552 (O_1552,N_14811,N_14812);
or UO_1553 (O_1553,N_14969,N_14770);
and UO_1554 (O_1554,N_14833,N_14970);
or UO_1555 (O_1555,N_14959,N_14859);
nor UO_1556 (O_1556,N_14932,N_14822);
xor UO_1557 (O_1557,N_14956,N_14901);
nor UO_1558 (O_1558,N_14914,N_14838);
or UO_1559 (O_1559,N_14843,N_14828);
and UO_1560 (O_1560,N_14920,N_14782);
nor UO_1561 (O_1561,N_14942,N_14830);
or UO_1562 (O_1562,N_14982,N_14961);
xor UO_1563 (O_1563,N_14963,N_14783);
nor UO_1564 (O_1564,N_14866,N_14762);
and UO_1565 (O_1565,N_14940,N_14886);
or UO_1566 (O_1566,N_14999,N_14998);
nand UO_1567 (O_1567,N_14940,N_14833);
or UO_1568 (O_1568,N_14934,N_14957);
or UO_1569 (O_1569,N_14821,N_14769);
nand UO_1570 (O_1570,N_14908,N_14977);
nor UO_1571 (O_1571,N_14908,N_14973);
nand UO_1572 (O_1572,N_14839,N_14980);
xnor UO_1573 (O_1573,N_14849,N_14972);
xor UO_1574 (O_1574,N_14985,N_14959);
nor UO_1575 (O_1575,N_14928,N_14908);
nand UO_1576 (O_1576,N_14996,N_14755);
nand UO_1577 (O_1577,N_14924,N_14906);
nand UO_1578 (O_1578,N_14870,N_14904);
nand UO_1579 (O_1579,N_14780,N_14936);
nand UO_1580 (O_1580,N_14917,N_14980);
or UO_1581 (O_1581,N_14852,N_14947);
nand UO_1582 (O_1582,N_14781,N_14817);
nand UO_1583 (O_1583,N_14976,N_14914);
nand UO_1584 (O_1584,N_14832,N_14972);
nand UO_1585 (O_1585,N_14840,N_14879);
and UO_1586 (O_1586,N_14912,N_14845);
or UO_1587 (O_1587,N_14889,N_14862);
nor UO_1588 (O_1588,N_14913,N_14925);
and UO_1589 (O_1589,N_14753,N_14987);
xor UO_1590 (O_1590,N_14822,N_14979);
nor UO_1591 (O_1591,N_14983,N_14926);
nand UO_1592 (O_1592,N_14846,N_14992);
or UO_1593 (O_1593,N_14888,N_14944);
or UO_1594 (O_1594,N_14935,N_14814);
nand UO_1595 (O_1595,N_14779,N_14773);
nor UO_1596 (O_1596,N_14882,N_14968);
or UO_1597 (O_1597,N_14948,N_14921);
nand UO_1598 (O_1598,N_14770,N_14942);
and UO_1599 (O_1599,N_14925,N_14946);
or UO_1600 (O_1600,N_14931,N_14754);
nand UO_1601 (O_1601,N_14947,N_14759);
or UO_1602 (O_1602,N_14998,N_14798);
nand UO_1603 (O_1603,N_14991,N_14933);
nand UO_1604 (O_1604,N_14968,N_14997);
nor UO_1605 (O_1605,N_14823,N_14977);
nor UO_1606 (O_1606,N_14918,N_14829);
nor UO_1607 (O_1607,N_14873,N_14766);
nand UO_1608 (O_1608,N_14917,N_14897);
nand UO_1609 (O_1609,N_14887,N_14961);
nand UO_1610 (O_1610,N_14964,N_14936);
nor UO_1611 (O_1611,N_14902,N_14929);
nand UO_1612 (O_1612,N_14827,N_14829);
and UO_1613 (O_1613,N_14997,N_14821);
and UO_1614 (O_1614,N_14995,N_14874);
or UO_1615 (O_1615,N_14975,N_14941);
nor UO_1616 (O_1616,N_14862,N_14789);
and UO_1617 (O_1617,N_14771,N_14982);
xor UO_1618 (O_1618,N_14773,N_14903);
or UO_1619 (O_1619,N_14855,N_14989);
and UO_1620 (O_1620,N_14929,N_14887);
nand UO_1621 (O_1621,N_14809,N_14875);
and UO_1622 (O_1622,N_14892,N_14845);
nor UO_1623 (O_1623,N_14976,N_14974);
and UO_1624 (O_1624,N_14806,N_14825);
nor UO_1625 (O_1625,N_14973,N_14833);
or UO_1626 (O_1626,N_14781,N_14786);
nor UO_1627 (O_1627,N_14997,N_14918);
and UO_1628 (O_1628,N_14894,N_14970);
or UO_1629 (O_1629,N_14984,N_14760);
nor UO_1630 (O_1630,N_14970,N_14766);
and UO_1631 (O_1631,N_14915,N_14795);
xnor UO_1632 (O_1632,N_14797,N_14842);
nor UO_1633 (O_1633,N_14775,N_14870);
or UO_1634 (O_1634,N_14762,N_14974);
nor UO_1635 (O_1635,N_14865,N_14921);
or UO_1636 (O_1636,N_14828,N_14833);
or UO_1637 (O_1637,N_14819,N_14992);
nand UO_1638 (O_1638,N_14760,N_14819);
and UO_1639 (O_1639,N_14763,N_14778);
or UO_1640 (O_1640,N_14838,N_14996);
nand UO_1641 (O_1641,N_14875,N_14937);
or UO_1642 (O_1642,N_14968,N_14797);
and UO_1643 (O_1643,N_14981,N_14884);
nor UO_1644 (O_1644,N_14776,N_14754);
nand UO_1645 (O_1645,N_14961,N_14971);
nand UO_1646 (O_1646,N_14987,N_14816);
or UO_1647 (O_1647,N_14995,N_14970);
and UO_1648 (O_1648,N_14959,N_14758);
nand UO_1649 (O_1649,N_14827,N_14885);
nand UO_1650 (O_1650,N_14942,N_14753);
nor UO_1651 (O_1651,N_14919,N_14816);
nand UO_1652 (O_1652,N_14772,N_14878);
nand UO_1653 (O_1653,N_14803,N_14832);
nand UO_1654 (O_1654,N_14935,N_14787);
nor UO_1655 (O_1655,N_14786,N_14932);
or UO_1656 (O_1656,N_14855,N_14929);
nor UO_1657 (O_1657,N_14994,N_14843);
and UO_1658 (O_1658,N_14861,N_14774);
and UO_1659 (O_1659,N_14772,N_14766);
or UO_1660 (O_1660,N_14834,N_14983);
nand UO_1661 (O_1661,N_14991,N_14946);
and UO_1662 (O_1662,N_14769,N_14943);
or UO_1663 (O_1663,N_14801,N_14942);
nand UO_1664 (O_1664,N_14837,N_14800);
or UO_1665 (O_1665,N_14843,N_14996);
and UO_1666 (O_1666,N_14771,N_14750);
and UO_1667 (O_1667,N_14878,N_14852);
nor UO_1668 (O_1668,N_14902,N_14793);
and UO_1669 (O_1669,N_14795,N_14790);
and UO_1670 (O_1670,N_14995,N_14957);
or UO_1671 (O_1671,N_14926,N_14951);
and UO_1672 (O_1672,N_14872,N_14986);
or UO_1673 (O_1673,N_14916,N_14967);
and UO_1674 (O_1674,N_14913,N_14929);
and UO_1675 (O_1675,N_14841,N_14992);
and UO_1676 (O_1676,N_14765,N_14992);
and UO_1677 (O_1677,N_14767,N_14916);
nand UO_1678 (O_1678,N_14884,N_14837);
and UO_1679 (O_1679,N_14813,N_14891);
nand UO_1680 (O_1680,N_14802,N_14889);
nand UO_1681 (O_1681,N_14948,N_14903);
nand UO_1682 (O_1682,N_14838,N_14966);
nor UO_1683 (O_1683,N_14840,N_14894);
nand UO_1684 (O_1684,N_14952,N_14840);
or UO_1685 (O_1685,N_14974,N_14792);
or UO_1686 (O_1686,N_14992,N_14852);
nand UO_1687 (O_1687,N_14871,N_14795);
xor UO_1688 (O_1688,N_14913,N_14850);
nor UO_1689 (O_1689,N_14930,N_14857);
nand UO_1690 (O_1690,N_14885,N_14775);
nor UO_1691 (O_1691,N_14860,N_14913);
xnor UO_1692 (O_1692,N_14846,N_14781);
or UO_1693 (O_1693,N_14941,N_14977);
nand UO_1694 (O_1694,N_14933,N_14961);
or UO_1695 (O_1695,N_14904,N_14887);
nand UO_1696 (O_1696,N_14939,N_14770);
and UO_1697 (O_1697,N_14979,N_14900);
nor UO_1698 (O_1698,N_14850,N_14760);
or UO_1699 (O_1699,N_14858,N_14760);
nand UO_1700 (O_1700,N_14750,N_14804);
and UO_1701 (O_1701,N_14839,N_14755);
xor UO_1702 (O_1702,N_14819,N_14832);
and UO_1703 (O_1703,N_14752,N_14837);
or UO_1704 (O_1704,N_14820,N_14856);
xor UO_1705 (O_1705,N_14925,N_14768);
and UO_1706 (O_1706,N_14873,N_14768);
nor UO_1707 (O_1707,N_14949,N_14927);
or UO_1708 (O_1708,N_14879,N_14949);
and UO_1709 (O_1709,N_14885,N_14876);
nand UO_1710 (O_1710,N_14913,N_14994);
nand UO_1711 (O_1711,N_14924,N_14750);
nor UO_1712 (O_1712,N_14760,N_14959);
and UO_1713 (O_1713,N_14862,N_14996);
xor UO_1714 (O_1714,N_14852,N_14825);
xnor UO_1715 (O_1715,N_14890,N_14843);
or UO_1716 (O_1716,N_14974,N_14861);
nand UO_1717 (O_1717,N_14906,N_14863);
xnor UO_1718 (O_1718,N_14921,N_14961);
nor UO_1719 (O_1719,N_14764,N_14957);
nand UO_1720 (O_1720,N_14827,N_14866);
and UO_1721 (O_1721,N_14836,N_14995);
nor UO_1722 (O_1722,N_14943,N_14861);
and UO_1723 (O_1723,N_14953,N_14932);
nor UO_1724 (O_1724,N_14950,N_14753);
nand UO_1725 (O_1725,N_14845,N_14913);
nor UO_1726 (O_1726,N_14778,N_14919);
and UO_1727 (O_1727,N_14992,N_14987);
and UO_1728 (O_1728,N_14992,N_14895);
nand UO_1729 (O_1729,N_14871,N_14878);
nor UO_1730 (O_1730,N_14855,N_14966);
nand UO_1731 (O_1731,N_14849,N_14754);
nor UO_1732 (O_1732,N_14815,N_14861);
nand UO_1733 (O_1733,N_14887,N_14985);
nor UO_1734 (O_1734,N_14765,N_14825);
or UO_1735 (O_1735,N_14823,N_14776);
or UO_1736 (O_1736,N_14796,N_14956);
nand UO_1737 (O_1737,N_14754,N_14839);
nor UO_1738 (O_1738,N_14783,N_14873);
and UO_1739 (O_1739,N_14885,N_14947);
and UO_1740 (O_1740,N_14834,N_14926);
and UO_1741 (O_1741,N_14874,N_14790);
nand UO_1742 (O_1742,N_14967,N_14806);
and UO_1743 (O_1743,N_14861,N_14795);
nor UO_1744 (O_1744,N_14963,N_14787);
or UO_1745 (O_1745,N_14788,N_14924);
nor UO_1746 (O_1746,N_14874,N_14948);
nand UO_1747 (O_1747,N_14872,N_14860);
or UO_1748 (O_1748,N_14808,N_14973);
and UO_1749 (O_1749,N_14935,N_14980);
and UO_1750 (O_1750,N_14961,N_14926);
or UO_1751 (O_1751,N_14980,N_14912);
nor UO_1752 (O_1752,N_14940,N_14989);
nand UO_1753 (O_1753,N_14984,N_14771);
and UO_1754 (O_1754,N_14803,N_14786);
nor UO_1755 (O_1755,N_14940,N_14796);
or UO_1756 (O_1756,N_14944,N_14980);
and UO_1757 (O_1757,N_14965,N_14758);
and UO_1758 (O_1758,N_14773,N_14940);
nor UO_1759 (O_1759,N_14938,N_14879);
nand UO_1760 (O_1760,N_14994,N_14773);
nand UO_1761 (O_1761,N_14959,N_14820);
and UO_1762 (O_1762,N_14915,N_14772);
xnor UO_1763 (O_1763,N_14869,N_14839);
xnor UO_1764 (O_1764,N_14794,N_14894);
nand UO_1765 (O_1765,N_14940,N_14755);
nor UO_1766 (O_1766,N_14755,N_14884);
xnor UO_1767 (O_1767,N_14763,N_14999);
nand UO_1768 (O_1768,N_14928,N_14967);
and UO_1769 (O_1769,N_14844,N_14868);
and UO_1770 (O_1770,N_14815,N_14802);
or UO_1771 (O_1771,N_14765,N_14925);
nor UO_1772 (O_1772,N_14825,N_14927);
nor UO_1773 (O_1773,N_14946,N_14984);
or UO_1774 (O_1774,N_14892,N_14766);
or UO_1775 (O_1775,N_14816,N_14754);
xnor UO_1776 (O_1776,N_14927,N_14936);
nand UO_1777 (O_1777,N_14900,N_14980);
nand UO_1778 (O_1778,N_14796,N_14883);
or UO_1779 (O_1779,N_14876,N_14916);
or UO_1780 (O_1780,N_14954,N_14894);
or UO_1781 (O_1781,N_14866,N_14849);
nand UO_1782 (O_1782,N_14885,N_14849);
nand UO_1783 (O_1783,N_14815,N_14775);
or UO_1784 (O_1784,N_14758,N_14752);
xnor UO_1785 (O_1785,N_14935,N_14912);
or UO_1786 (O_1786,N_14961,N_14810);
or UO_1787 (O_1787,N_14838,N_14750);
nor UO_1788 (O_1788,N_14880,N_14830);
and UO_1789 (O_1789,N_14984,N_14974);
nor UO_1790 (O_1790,N_14884,N_14899);
nand UO_1791 (O_1791,N_14919,N_14758);
nor UO_1792 (O_1792,N_14768,N_14888);
or UO_1793 (O_1793,N_14987,N_14759);
nand UO_1794 (O_1794,N_14837,N_14939);
nor UO_1795 (O_1795,N_14866,N_14956);
nand UO_1796 (O_1796,N_14969,N_14899);
and UO_1797 (O_1797,N_14882,N_14818);
nor UO_1798 (O_1798,N_14996,N_14994);
nor UO_1799 (O_1799,N_14858,N_14854);
xnor UO_1800 (O_1800,N_14857,N_14953);
nand UO_1801 (O_1801,N_14819,N_14868);
nand UO_1802 (O_1802,N_14883,N_14828);
and UO_1803 (O_1803,N_14754,N_14793);
xnor UO_1804 (O_1804,N_14792,N_14805);
and UO_1805 (O_1805,N_14884,N_14769);
nor UO_1806 (O_1806,N_14840,N_14814);
or UO_1807 (O_1807,N_14962,N_14982);
xor UO_1808 (O_1808,N_14992,N_14792);
nor UO_1809 (O_1809,N_14921,N_14840);
nor UO_1810 (O_1810,N_14802,N_14794);
nand UO_1811 (O_1811,N_14905,N_14793);
or UO_1812 (O_1812,N_14837,N_14897);
or UO_1813 (O_1813,N_14976,N_14954);
nor UO_1814 (O_1814,N_14882,N_14975);
and UO_1815 (O_1815,N_14871,N_14911);
nand UO_1816 (O_1816,N_14891,N_14868);
nor UO_1817 (O_1817,N_14848,N_14899);
nor UO_1818 (O_1818,N_14759,N_14936);
and UO_1819 (O_1819,N_14915,N_14775);
nor UO_1820 (O_1820,N_14782,N_14932);
xnor UO_1821 (O_1821,N_14968,N_14904);
or UO_1822 (O_1822,N_14814,N_14838);
nand UO_1823 (O_1823,N_14906,N_14991);
and UO_1824 (O_1824,N_14801,N_14779);
nand UO_1825 (O_1825,N_14871,N_14963);
nor UO_1826 (O_1826,N_14879,N_14809);
nor UO_1827 (O_1827,N_14844,N_14930);
nand UO_1828 (O_1828,N_14774,N_14908);
and UO_1829 (O_1829,N_14834,N_14991);
and UO_1830 (O_1830,N_14915,N_14847);
nand UO_1831 (O_1831,N_14866,N_14752);
and UO_1832 (O_1832,N_14785,N_14986);
nor UO_1833 (O_1833,N_14976,N_14851);
or UO_1834 (O_1834,N_14831,N_14792);
nor UO_1835 (O_1835,N_14911,N_14812);
or UO_1836 (O_1836,N_14823,N_14842);
nor UO_1837 (O_1837,N_14943,N_14982);
or UO_1838 (O_1838,N_14791,N_14818);
nand UO_1839 (O_1839,N_14786,N_14759);
and UO_1840 (O_1840,N_14820,N_14860);
or UO_1841 (O_1841,N_14798,N_14750);
and UO_1842 (O_1842,N_14987,N_14838);
nand UO_1843 (O_1843,N_14774,N_14963);
nor UO_1844 (O_1844,N_14875,N_14848);
or UO_1845 (O_1845,N_14923,N_14909);
or UO_1846 (O_1846,N_14802,N_14903);
and UO_1847 (O_1847,N_14918,N_14890);
nor UO_1848 (O_1848,N_14815,N_14826);
nor UO_1849 (O_1849,N_14958,N_14758);
nand UO_1850 (O_1850,N_14892,N_14911);
nand UO_1851 (O_1851,N_14857,N_14801);
nand UO_1852 (O_1852,N_14975,N_14887);
xnor UO_1853 (O_1853,N_14966,N_14760);
xor UO_1854 (O_1854,N_14946,N_14873);
nor UO_1855 (O_1855,N_14922,N_14893);
or UO_1856 (O_1856,N_14930,N_14756);
or UO_1857 (O_1857,N_14929,N_14846);
nand UO_1858 (O_1858,N_14787,N_14953);
nor UO_1859 (O_1859,N_14850,N_14782);
and UO_1860 (O_1860,N_14777,N_14943);
nor UO_1861 (O_1861,N_14760,N_14823);
or UO_1862 (O_1862,N_14946,N_14885);
xnor UO_1863 (O_1863,N_14890,N_14782);
or UO_1864 (O_1864,N_14844,N_14806);
nor UO_1865 (O_1865,N_14843,N_14910);
or UO_1866 (O_1866,N_14808,N_14802);
or UO_1867 (O_1867,N_14938,N_14925);
and UO_1868 (O_1868,N_14773,N_14761);
and UO_1869 (O_1869,N_14983,N_14883);
nand UO_1870 (O_1870,N_14839,N_14771);
and UO_1871 (O_1871,N_14878,N_14891);
or UO_1872 (O_1872,N_14910,N_14750);
nand UO_1873 (O_1873,N_14933,N_14976);
and UO_1874 (O_1874,N_14955,N_14817);
and UO_1875 (O_1875,N_14947,N_14869);
xor UO_1876 (O_1876,N_14864,N_14883);
nand UO_1877 (O_1877,N_14966,N_14755);
nor UO_1878 (O_1878,N_14969,N_14992);
xor UO_1879 (O_1879,N_14874,N_14946);
or UO_1880 (O_1880,N_14873,N_14891);
and UO_1881 (O_1881,N_14760,N_14999);
or UO_1882 (O_1882,N_14940,N_14977);
or UO_1883 (O_1883,N_14904,N_14753);
or UO_1884 (O_1884,N_14967,N_14906);
nand UO_1885 (O_1885,N_14904,N_14842);
xnor UO_1886 (O_1886,N_14780,N_14878);
and UO_1887 (O_1887,N_14795,N_14853);
xor UO_1888 (O_1888,N_14925,N_14912);
xor UO_1889 (O_1889,N_14890,N_14986);
nor UO_1890 (O_1890,N_14789,N_14780);
nor UO_1891 (O_1891,N_14878,N_14916);
or UO_1892 (O_1892,N_14985,N_14848);
nor UO_1893 (O_1893,N_14954,N_14878);
xor UO_1894 (O_1894,N_14795,N_14929);
nor UO_1895 (O_1895,N_14932,N_14976);
nand UO_1896 (O_1896,N_14875,N_14836);
nand UO_1897 (O_1897,N_14899,N_14781);
nor UO_1898 (O_1898,N_14925,N_14752);
and UO_1899 (O_1899,N_14896,N_14997);
or UO_1900 (O_1900,N_14906,N_14790);
xnor UO_1901 (O_1901,N_14755,N_14879);
or UO_1902 (O_1902,N_14813,N_14763);
and UO_1903 (O_1903,N_14807,N_14763);
or UO_1904 (O_1904,N_14825,N_14827);
nand UO_1905 (O_1905,N_14968,N_14971);
xnor UO_1906 (O_1906,N_14943,N_14851);
nor UO_1907 (O_1907,N_14929,N_14949);
nand UO_1908 (O_1908,N_14853,N_14750);
xnor UO_1909 (O_1909,N_14906,N_14848);
nand UO_1910 (O_1910,N_14859,N_14900);
and UO_1911 (O_1911,N_14890,N_14766);
nor UO_1912 (O_1912,N_14900,N_14838);
and UO_1913 (O_1913,N_14967,N_14848);
nor UO_1914 (O_1914,N_14755,N_14855);
nor UO_1915 (O_1915,N_14941,N_14921);
xnor UO_1916 (O_1916,N_14834,N_14808);
or UO_1917 (O_1917,N_14774,N_14973);
nor UO_1918 (O_1918,N_14959,N_14839);
nor UO_1919 (O_1919,N_14758,N_14983);
xor UO_1920 (O_1920,N_14911,N_14803);
nand UO_1921 (O_1921,N_14823,N_14984);
nor UO_1922 (O_1922,N_14882,N_14771);
nor UO_1923 (O_1923,N_14969,N_14793);
xnor UO_1924 (O_1924,N_14979,N_14859);
nand UO_1925 (O_1925,N_14894,N_14752);
nand UO_1926 (O_1926,N_14987,N_14750);
nand UO_1927 (O_1927,N_14769,N_14864);
nor UO_1928 (O_1928,N_14952,N_14921);
nor UO_1929 (O_1929,N_14825,N_14828);
nand UO_1930 (O_1930,N_14873,N_14980);
nor UO_1931 (O_1931,N_14827,N_14944);
or UO_1932 (O_1932,N_14825,N_14998);
and UO_1933 (O_1933,N_14962,N_14917);
nor UO_1934 (O_1934,N_14784,N_14811);
nor UO_1935 (O_1935,N_14869,N_14860);
nor UO_1936 (O_1936,N_14977,N_14998);
or UO_1937 (O_1937,N_14861,N_14828);
nand UO_1938 (O_1938,N_14950,N_14798);
nor UO_1939 (O_1939,N_14898,N_14928);
nor UO_1940 (O_1940,N_14803,N_14969);
or UO_1941 (O_1941,N_14875,N_14814);
nor UO_1942 (O_1942,N_14760,N_14774);
and UO_1943 (O_1943,N_14939,N_14980);
or UO_1944 (O_1944,N_14794,N_14753);
nand UO_1945 (O_1945,N_14779,N_14874);
nand UO_1946 (O_1946,N_14952,N_14792);
or UO_1947 (O_1947,N_14935,N_14767);
or UO_1948 (O_1948,N_14915,N_14950);
nor UO_1949 (O_1949,N_14960,N_14891);
or UO_1950 (O_1950,N_14908,N_14761);
and UO_1951 (O_1951,N_14887,N_14934);
nor UO_1952 (O_1952,N_14886,N_14892);
nand UO_1953 (O_1953,N_14996,N_14974);
or UO_1954 (O_1954,N_14831,N_14939);
nand UO_1955 (O_1955,N_14839,N_14781);
xor UO_1956 (O_1956,N_14810,N_14877);
nor UO_1957 (O_1957,N_14894,N_14851);
or UO_1958 (O_1958,N_14922,N_14902);
or UO_1959 (O_1959,N_14857,N_14810);
and UO_1960 (O_1960,N_14812,N_14930);
or UO_1961 (O_1961,N_14805,N_14921);
nor UO_1962 (O_1962,N_14775,N_14997);
and UO_1963 (O_1963,N_14902,N_14979);
xor UO_1964 (O_1964,N_14802,N_14935);
and UO_1965 (O_1965,N_14952,N_14850);
and UO_1966 (O_1966,N_14795,N_14752);
and UO_1967 (O_1967,N_14865,N_14917);
or UO_1968 (O_1968,N_14868,N_14825);
and UO_1969 (O_1969,N_14980,N_14806);
or UO_1970 (O_1970,N_14785,N_14841);
nand UO_1971 (O_1971,N_14793,N_14790);
and UO_1972 (O_1972,N_14934,N_14876);
nand UO_1973 (O_1973,N_14894,N_14838);
nand UO_1974 (O_1974,N_14983,N_14909);
nand UO_1975 (O_1975,N_14976,N_14834);
nor UO_1976 (O_1976,N_14946,N_14972);
or UO_1977 (O_1977,N_14763,N_14776);
or UO_1978 (O_1978,N_14983,N_14844);
or UO_1979 (O_1979,N_14965,N_14967);
xor UO_1980 (O_1980,N_14848,N_14950);
nor UO_1981 (O_1981,N_14761,N_14834);
and UO_1982 (O_1982,N_14924,N_14998);
or UO_1983 (O_1983,N_14893,N_14982);
nand UO_1984 (O_1984,N_14753,N_14993);
and UO_1985 (O_1985,N_14946,N_14767);
or UO_1986 (O_1986,N_14899,N_14908);
and UO_1987 (O_1987,N_14758,N_14874);
nor UO_1988 (O_1988,N_14916,N_14926);
nand UO_1989 (O_1989,N_14877,N_14826);
nand UO_1990 (O_1990,N_14882,N_14858);
and UO_1991 (O_1991,N_14954,N_14781);
or UO_1992 (O_1992,N_14979,N_14985);
or UO_1993 (O_1993,N_14767,N_14856);
nor UO_1994 (O_1994,N_14953,N_14826);
xor UO_1995 (O_1995,N_14869,N_14987);
nor UO_1996 (O_1996,N_14955,N_14769);
or UO_1997 (O_1997,N_14846,N_14778);
xnor UO_1998 (O_1998,N_14928,N_14846);
and UO_1999 (O_1999,N_14965,N_14946);
endmodule